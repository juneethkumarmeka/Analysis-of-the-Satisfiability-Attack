module basic_5000_50000_5000_25_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_668,In_2964);
and U1 (N_1,In_714,In_4103);
and U2 (N_2,In_146,In_623);
and U3 (N_3,In_1037,In_1220);
nor U4 (N_4,In_4680,In_2974);
nor U5 (N_5,In_4065,In_91);
nand U6 (N_6,In_1129,In_1515);
nor U7 (N_7,In_3621,In_2044);
nor U8 (N_8,In_2553,In_4972);
and U9 (N_9,In_1552,In_4049);
or U10 (N_10,In_2942,In_4189);
and U11 (N_11,In_4342,In_890);
or U12 (N_12,In_4806,In_1463);
or U13 (N_13,In_4528,In_1286);
or U14 (N_14,In_533,In_1748);
xor U15 (N_15,In_3701,In_4419);
nand U16 (N_16,In_4783,In_1284);
xnor U17 (N_17,In_296,In_2811);
and U18 (N_18,In_4709,In_2101);
xnor U19 (N_19,In_410,In_1900);
nor U20 (N_20,In_4693,In_2732);
and U21 (N_21,In_2304,In_2057);
and U22 (N_22,In_4984,In_900);
nand U23 (N_23,In_3528,In_4212);
xor U24 (N_24,In_966,In_4928);
xor U25 (N_25,In_1789,In_970);
nand U26 (N_26,In_1446,In_4257);
nor U27 (N_27,In_3113,In_984);
xor U28 (N_28,In_3912,In_2865);
nor U29 (N_29,In_581,In_4341);
nand U30 (N_30,In_3221,In_4601);
nand U31 (N_31,In_2658,In_1066);
and U32 (N_32,In_1973,In_4399);
or U33 (N_33,In_4921,In_3204);
nand U34 (N_34,In_2456,In_342);
nor U35 (N_35,In_3860,In_1353);
or U36 (N_36,In_4112,In_1257);
nor U37 (N_37,In_2807,In_854);
xor U38 (N_38,In_3906,In_1662);
or U39 (N_39,In_4454,In_1450);
nor U40 (N_40,In_2370,In_2579);
and U41 (N_41,In_2440,In_1548);
xor U42 (N_42,In_1094,In_525);
nand U43 (N_43,In_1486,In_3542);
xor U44 (N_44,In_2709,In_1691);
nand U45 (N_45,In_246,In_4417);
nand U46 (N_46,In_978,In_3414);
nor U47 (N_47,In_4588,In_4871);
or U48 (N_48,In_3579,In_1798);
nand U49 (N_49,In_3781,In_645);
and U50 (N_50,In_3729,In_4164);
xor U51 (N_51,In_2688,In_2405);
and U52 (N_52,In_85,In_3180);
nand U53 (N_53,In_618,In_317);
nand U54 (N_54,In_3532,In_4523);
and U55 (N_55,In_3474,In_1437);
xnor U56 (N_56,In_2008,In_2866);
nand U57 (N_57,In_2661,In_4444);
nand U58 (N_58,In_3775,In_3144);
xor U59 (N_59,In_365,In_4014);
nand U60 (N_60,In_1641,In_2346);
or U61 (N_61,In_4083,In_1851);
nand U62 (N_62,In_251,In_2186);
nand U63 (N_63,In_1524,In_1895);
and U64 (N_64,In_2045,In_281);
and U65 (N_65,In_1656,In_4824);
xnor U66 (N_66,In_823,In_1199);
and U67 (N_67,In_1022,In_4916);
or U68 (N_68,In_2264,In_53);
nor U69 (N_69,In_4079,In_4794);
nor U70 (N_70,In_467,In_1473);
nor U71 (N_71,In_4911,In_3615);
and U72 (N_72,In_4954,In_3009);
nand U73 (N_73,In_1146,In_4532);
and U74 (N_74,In_4231,In_2891);
and U75 (N_75,In_695,In_3027);
nor U76 (N_76,In_2544,In_1593);
nand U77 (N_77,In_2261,In_3051);
xor U78 (N_78,In_2337,In_2576);
nor U79 (N_79,In_3226,In_3718);
xnor U80 (N_80,In_1665,In_1152);
nor U81 (N_81,In_2495,In_3963);
xor U82 (N_82,In_1669,In_4360);
nand U83 (N_83,In_4271,In_248);
xnor U84 (N_84,In_1390,In_4756);
nand U85 (N_85,In_4787,In_1890);
nand U86 (N_86,In_1738,In_3823);
xnor U87 (N_87,In_4622,In_3698);
nand U88 (N_88,In_3185,In_3451);
xor U89 (N_89,In_547,In_130);
or U90 (N_90,In_4799,In_4747);
nor U91 (N_91,In_812,In_4701);
or U92 (N_92,In_4283,In_4035);
xor U93 (N_93,In_958,In_1767);
xor U94 (N_94,In_1521,In_3037);
nand U95 (N_95,In_2721,In_1763);
nor U96 (N_96,In_3067,In_273);
nor U97 (N_97,In_876,In_711);
or U98 (N_98,In_4643,In_1931);
and U99 (N_99,In_1359,In_767);
or U100 (N_100,In_3398,In_2616);
nand U101 (N_101,In_670,In_4941);
or U102 (N_102,In_4520,In_4834);
nand U103 (N_103,In_308,In_2394);
xnor U104 (N_104,In_537,In_1779);
nand U105 (N_105,In_1154,In_1417);
xnor U106 (N_106,In_4619,In_2284);
or U107 (N_107,In_3952,In_49);
xnor U108 (N_108,In_3564,In_3863);
and U109 (N_109,In_381,In_4133);
nand U110 (N_110,In_4544,In_1468);
nor U111 (N_111,In_4440,In_1025);
nand U112 (N_112,In_4255,In_4561);
nand U113 (N_113,In_1668,In_2242);
xnor U114 (N_114,In_2682,In_4056);
nor U115 (N_115,In_2859,In_4980);
nand U116 (N_116,In_1855,In_2410);
nor U117 (N_117,In_1651,In_3201);
or U118 (N_118,In_2398,In_797);
and U119 (N_119,In_2366,In_2283);
or U120 (N_120,In_156,In_3272);
nor U121 (N_121,In_1397,In_4117);
and U122 (N_122,In_124,In_2637);
xnor U123 (N_123,In_4839,In_3846);
or U124 (N_124,In_3991,In_1938);
nand U125 (N_125,In_1781,In_2787);
nor U126 (N_126,In_451,In_3352);
and U127 (N_127,In_2670,In_2292);
xor U128 (N_128,In_2023,In_4404);
nand U129 (N_129,In_1331,In_4141);
or U130 (N_130,In_2607,In_2014);
or U131 (N_131,In_1635,In_2236);
nand U132 (N_132,In_3752,In_3102);
and U133 (N_133,In_2977,In_1147);
nand U134 (N_134,In_1646,In_4529);
or U135 (N_135,In_3560,In_3138);
nor U136 (N_136,In_2493,In_4193);
or U137 (N_137,In_408,In_834);
xnor U138 (N_138,In_931,In_4307);
and U139 (N_139,In_107,In_2517);
or U140 (N_140,In_3047,In_3189);
nand U141 (N_141,In_1113,In_2208);
nand U142 (N_142,In_1160,In_4940);
nor U143 (N_143,In_3114,In_535);
or U144 (N_144,In_538,In_2981);
nand U145 (N_145,In_968,In_4067);
nor U146 (N_146,In_4265,In_2263);
nor U147 (N_147,In_153,In_3499);
nand U148 (N_148,In_3676,In_1616);
nor U149 (N_149,In_932,In_3919);
nor U150 (N_150,In_4568,In_4856);
nand U151 (N_151,In_4971,In_3458);
or U152 (N_152,In_3750,In_2600);
or U153 (N_153,In_3192,In_3657);
nor U154 (N_154,In_440,In_2021);
nand U155 (N_155,In_4483,In_2880);
xnor U156 (N_156,In_1716,In_4229);
xnor U157 (N_157,In_364,In_496);
and U158 (N_158,In_2274,In_1126);
xnor U159 (N_159,In_64,In_4763);
nand U160 (N_160,In_1679,In_2796);
and U161 (N_161,In_4986,In_1339);
xor U162 (N_162,In_1686,In_1557);
nand U163 (N_163,In_4884,In_1989);
or U164 (N_164,In_889,In_2597);
nand U165 (N_165,In_2349,In_2334);
or U166 (N_166,In_1513,In_898);
or U167 (N_167,In_3257,In_3531);
or U168 (N_168,In_2845,In_3374);
xnor U169 (N_169,In_716,In_2673);
xor U170 (N_170,In_24,In_2590);
nor U171 (N_171,In_4861,In_2126);
and U172 (N_172,In_4654,In_2190);
nor U173 (N_173,In_4573,In_222);
or U174 (N_174,In_4198,In_956);
nand U175 (N_175,In_4148,In_1768);
and U176 (N_176,In_2698,In_974);
nor U177 (N_177,In_3856,In_1831);
nand U178 (N_178,In_3042,In_4685);
xnor U179 (N_179,In_4280,In_151);
or U180 (N_180,In_1326,In_2238);
xnor U181 (N_181,In_2257,In_2804);
xnor U182 (N_182,In_2656,In_1754);
nand U183 (N_183,In_3259,In_2737);
nor U184 (N_184,In_2327,In_1366);
nand U185 (N_185,In_1806,In_875);
nor U186 (N_186,In_4492,In_3332);
or U187 (N_187,In_3251,In_295);
nand U188 (N_188,In_516,In_4114);
and U189 (N_189,In_3101,In_388);
xnor U190 (N_190,In_4807,In_3538);
nand U191 (N_191,In_3589,In_2062);
xor U192 (N_192,In_475,In_1912);
and U193 (N_193,In_2736,In_1687);
nand U194 (N_194,In_4062,In_1300);
nor U195 (N_195,In_4479,In_4167);
nor U196 (N_196,In_1902,In_701);
nor U197 (N_197,In_1554,In_4119);
or U198 (N_198,In_710,In_2149);
nand U199 (N_199,In_3566,In_4223);
and U200 (N_200,In_1345,In_4534);
xor U201 (N_201,In_4660,In_3696);
nand U202 (N_202,In_3899,In_3525);
or U203 (N_203,In_92,In_4462);
xor U204 (N_204,In_461,In_3671);
and U205 (N_205,In_3040,In_2157);
nor U206 (N_206,In_3596,In_1528);
or U207 (N_207,In_3078,In_933);
xor U208 (N_208,In_1215,In_340);
or U209 (N_209,In_3306,In_4388);
and U210 (N_210,In_2901,In_1231);
xor U211 (N_211,In_2183,In_1360);
nor U212 (N_212,In_4951,In_550);
or U213 (N_213,In_989,In_3502);
or U214 (N_214,In_3409,In_1292);
nand U215 (N_215,In_916,In_4927);
and U216 (N_216,In_393,In_1044);
and U217 (N_217,In_3521,In_2154);
xor U218 (N_218,In_4368,In_913);
or U219 (N_219,In_1032,In_600);
or U220 (N_220,In_4249,In_565);
and U221 (N_221,In_644,In_1774);
nor U222 (N_222,In_1550,In_2067);
nand U223 (N_223,In_4599,In_4098);
nor U224 (N_224,In_83,In_4590);
nand U225 (N_225,In_4298,In_4044);
nand U226 (N_226,In_87,In_2818);
or U227 (N_227,In_2547,In_3291);
nand U228 (N_228,In_790,In_1074);
nor U229 (N_229,In_3449,In_4057);
nor U230 (N_230,In_4381,In_2623);
xor U231 (N_231,In_4731,In_2055);
and U232 (N_232,In_1277,In_4330);
nor U233 (N_233,In_2330,In_2114);
nor U234 (N_234,In_1853,In_3748);
and U235 (N_235,In_3762,In_2123);
nor U236 (N_236,In_1186,In_2924);
or U237 (N_237,In_655,In_2505);
xnor U238 (N_238,In_3650,In_2543);
nor U239 (N_239,In_2396,In_753);
xnor U240 (N_240,In_4109,In_2674);
nor U241 (N_241,In_4463,In_1881);
nor U242 (N_242,In_1703,In_563);
and U243 (N_243,In_2905,In_3982);
nand U244 (N_244,In_1083,In_4585);
or U245 (N_245,In_4482,In_4220);
or U246 (N_246,In_3642,In_3243);
xor U247 (N_247,In_1375,In_4400);
xnor U248 (N_248,In_3703,In_1442);
xor U249 (N_249,In_2426,In_948);
nand U250 (N_250,In_2163,In_522);
nand U251 (N_251,In_3710,In_4749);
nand U252 (N_252,In_2446,In_3129);
and U253 (N_253,In_4459,In_333);
nand U254 (N_254,In_835,In_2357);
xnor U255 (N_255,In_2680,In_1761);
or U256 (N_256,In_4879,In_3280);
xor U257 (N_257,In_3225,In_975);
xor U258 (N_258,In_4161,In_4153);
xnor U259 (N_259,In_397,In_1002);
nor U260 (N_260,In_3063,In_2249);
xnor U261 (N_261,In_2423,In_4843);
nand U262 (N_262,In_2235,In_3784);
nor U263 (N_263,In_386,In_2816);
xnor U264 (N_264,In_720,In_2138);
nor U265 (N_265,In_3307,In_2244);
xor U266 (N_266,In_1033,In_1648);
nand U267 (N_267,In_576,In_532);
and U268 (N_268,In_4258,In_3723);
xor U269 (N_269,In_3337,In_1117);
or U270 (N_270,In_3890,In_424);
or U271 (N_271,In_1050,In_3794);
nor U272 (N_272,In_4346,In_3686);
nand U273 (N_273,In_1079,In_189);
xnor U274 (N_274,In_2609,In_1261);
and U275 (N_275,In_1183,In_558);
nor U276 (N_276,In_4810,In_2795);
nor U277 (N_277,In_3377,In_2004);
nor U278 (N_278,In_73,In_3881);
nand U279 (N_279,In_4210,In_2710);
nor U280 (N_280,In_4636,In_4581);
nor U281 (N_281,In_1886,In_1492);
nor U282 (N_282,In_4978,In_93);
nor U283 (N_283,In_2742,In_2910);
and U284 (N_284,In_1872,In_3660);
xor U285 (N_285,In_2518,In_4465);
nand U286 (N_286,In_3341,In_4647);
and U287 (N_287,In_990,In_3817);
and U288 (N_288,In_2417,In_731);
xor U289 (N_289,In_1356,In_3746);
or U290 (N_290,In_432,In_3446);
xnor U291 (N_291,In_1475,In_2936);
nor U292 (N_292,In_2539,In_1801);
nand U293 (N_293,In_4005,In_2326);
and U294 (N_294,In_1553,In_3223);
and U295 (N_295,In_4841,In_1047);
nand U296 (N_296,In_3420,In_1558);
nand U297 (N_297,In_2428,In_3049);
and U298 (N_298,In_3619,In_1631);
nand U299 (N_299,In_477,In_4548);
nand U300 (N_300,In_3549,In_169);
nor U301 (N_301,In_908,In_4142);
nor U302 (N_302,In_689,In_4719);
and U303 (N_303,In_3187,In_2512);
xnor U304 (N_304,In_4769,In_1052);
nor U305 (N_305,In_3422,In_1135);
nor U306 (N_306,In_3391,In_2900);
nor U307 (N_307,In_4269,In_3406);
nor U308 (N_308,In_896,In_3680);
nor U309 (N_309,In_1734,In_2010);
and U310 (N_310,In_4698,In_4696);
or U311 (N_311,In_1311,In_3069);
or U312 (N_312,In_4274,In_936);
and U313 (N_313,In_1522,In_765);
or U314 (N_314,In_658,In_4738);
xor U315 (N_315,In_831,In_2016);
xnor U316 (N_316,In_3007,In_3440);
and U317 (N_317,In_3764,In_3957);
and U318 (N_318,In_3289,In_2174);
nand U319 (N_319,In_4100,In_1663);
or U320 (N_320,In_2684,In_4620);
nor U321 (N_321,In_2206,In_4352);
nand U322 (N_322,In_771,In_4754);
nand U323 (N_323,In_3845,In_1670);
xor U324 (N_324,In_906,In_266);
xor U325 (N_325,In_4953,In_1019);
and U326 (N_326,In_3554,In_339);
or U327 (N_327,In_2514,In_3568);
nor U328 (N_328,In_607,In_3778);
and U329 (N_329,In_369,In_3541);
xor U330 (N_330,In_2983,In_1170);
nor U331 (N_331,In_3501,In_4616);
nor U332 (N_332,In_775,In_3324);
nand U333 (N_333,In_887,In_2689);
or U334 (N_334,In_3507,In_971);
xnor U335 (N_335,In_777,In_1472);
and U336 (N_336,In_4942,In_2935);
nand U337 (N_337,In_1263,In_55);
nor U338 (N_338,In_2888,In_3662);
or U339 (N_339,In_1488,In_415);
nand U340 (N_340,In_1601,In_969);
xnor U341 (N_341,In_4550,In_3519);
nor U342 (N_342,In_999,In_4932);
nand U343 (N_343,In_2077,In_821);
xor U344 (N_344,In_669,In_3600);
or U345 (N_345,In_2827,In_2681);
nand U346 (N_346,In_4335,In_1351);
or U347 (N_347,In_2963,In_1151);
nand U348 (N_348,In_242,In_1792);
or U349 (N_349,In_726,In_3236);
nor U350 (N_350,In_257,In_4134);
and U351 (N_351,In_991,In_4868);
or U352 (N_352,In_1958,In_4318);
xnor U353 (N_353,In_713,In_3924);
or U354 (N_354,In_2666,In_1934);
nand U355 (N_355,In_4786,In_1706);
nand U356 (N_356,In_4429,In_1992);
nor U357 (N_357,In_370,In_3512);
nand U358 (N_358,In_1308,In_676);
xnor U359 (N_359,In_4725,In_1101);
or U360 (N_360,In_518,In_4502);
or U361 (N_361,In_4895,In_4516);
xor U362 (N_362,In_1184,In_4642);
xor U363 (N_363,In_789,In_2105);
or U364 (N_364,In_1963,In_832);
and U365 (N_365,In_1699,In_3682);
nor U366 (N_366,In_4245,In_1585);
xnor U367 (N_367,In_2202,In_2619);
xnor U368 (N_368,In_4686,In_367);
xor U369 (N_369,In_2228,In_447);
and U370 (N_370,In_1636,In_4096);
or U371 (N_371,In_960,In_316);
nand U372 (N_372,In_3346,In_4517);
and U373 (N_373,In_2817,In_2205);
nor U374 (N_374,In_4877,In_3136);
or U375 (N_375,In_311,In_411);
and U376 (N_376,In_1112,In_1385);
or U377 (N_377,In_1659,In_1690);
and U378 (N_378,In_4692,In_4339);
and U379 (N_379,In_4387,In_3885);
nand U380 (N_380,In_2716,In_1494);
or U381 (N_381,In_4301,In_4624);
and U382 (N_382,In_2167,In_363);
and U383 (N_383,In_557,In_2175);
or U384 (N_384,In_4991,In_837);
or U385 (N_385,In_4905,In_443);
xnor U386 (N_386,In_155,In_926);
and U387 (N_387,In_2497,In_1325);
nand U388 (N_388,In_2707,In_3168);
xnor U389 (N_389,In_4498,In_548);
nand U390 (N_390,In_3454,In_2280);
nor U391 (N_391,In_852,In_2266);
nor U392 (N_392,In_3811,In_2295);
xor U393 (N_393,In_1911,In_1658);
nand U394 (N_394,In_285,In_2692);
or U395 (N_395,In_4358,In_3652);
xor U396 (N_396,In_2041,In_4332);
xnor U397 (N_397,In_4321,In_3064);
xor U398 (N_398,In_3767,In_2482);
nand U399 (N_399,In_882,In_4170);
or U400 (N_400,In_3843,In_774);
or U401 (N_401,In_1649,In_1588);
xor U402 (N_402,In_1192,In_4415);
and U403 (N_403,In_4540,In_4397);
nor U404 (N_404,In_3693,In_211);
nand U405 (N_405,In_1814,In_4575);
xor U406 (N_406,In_3882,In_2335);
and U407 (N_407,In_1723,In_703);
xnor U408 (N_408,In_2082,In_1667);
nand U409 (N_409,In_2513,In_885);
and U410 (N_410,In_1193,In_2465);
or U411 (N_411,In_2618,In_1371);
nor U412 (N_412,In_1626,In_904);
nand U413 (N_413,In_2533,In_4425);
nand U414 (N_414,In_145,In_3791);
xnor U415 (N_415,In_1408,In_985);
nand U416 (N_416,In_4551,In_1982);
and U417 (N_417,In_46,In_4542);
or U418 (N_418,In_769,In_1919);
and U419 (N_419,In_3770,In_728);
or U420 (N_420,In_2463,In_4094);
and U421 (N_421,In_3107,In_3066);
xor U422 (N_422,In_2146,In_858);
nand U423 (N_423,In_2191,In_1424);
and U424 (N_424,In_2402,In_3490);
nor U425 (N_425,In_4968,In_840);
and U426 (N_426,In_2837,In_1563);
and U427 (N_427,In_2291,In_4536);
or U428 (N_428,In_1861,In_3649);
nor U429 (N_429,In_1158,In_983);
and U430 (N_430,In_1544,In_292);
nor U431 (N_431,In_2120,In_360);
nor U432 (N_432,In_2856,In_1948);
nor U433 (N_433,In_2270,In_32);
xnor U434 (N_434,In_2654,In_2665);
nor U435 (N_435,In_1090,In_2662);
or U436 (N_436,In_78,In_3287);
xnor U437 (N_437,In_4537,In_458);
nand U438 (N_438,In_629,In_2971);
or U439 (N_439,In_392,In_3635);
xor U440 (N_440,In_907,In_825);
nand U441 (N_441,In_2430,In_1453);
nor U442 (N_442,In_592,In_1570);
and U443 (N_443,In_1114,In_770);
or U444 (N_444,In_3981,In_4236);
xnor U445 (N_445,In_1834,In_4595);
and U446 (N_446,In_800,In_4663);
and U447 (N_447,In_2229,In_2121);
or U448 (N_448,In_195,In_4037);
and U449 (N_449,In_2051,In_2520);
xor U450 (N_450,In_788,In_2777);
and U451 (N_451,In_3433,In_4937);
xnor U452 (N_452,In_1423,In_2649);
nand U453 (N_453,In_4836,In_3237);
or U454 (N_454,In_2005,In_2009);
nor U455 (N_455,In_4481,In_1946);
and U456 (N_456,In_1305,In_1055);
and U457 (N_457,In_338,In_33);
xor U458 (N_458,In_3343,In_2250);
nor U459 (N_459,In_1684,In_2902);
nor U460 (N_460,In_4402,In_921);
xnor U461 (N_461,In_4262,In_3712);
and U462 (N_462,In_1237,In_4204);
and U463 (N_463,In_2281,In_2080);
and U464 (N_464,In_3720,In_2371);
xnor U465 (N_465,In_2298,In_1248);
xor U466 (N_466,In_1014,In_2652);
xor U467 (N_467,In_4450,In_4466);
or U468 (N_468,In_1727,In_3252);
and U469 (N_469,In_735,In_3603);
nand U470 (N_470,In_1695,In_3363);
xor U471 (N_471,In_4602,In_4804);
nor U472 (N_472,In_2227,In_2610);
nor U473 (N_473,In_3432,In_1745);
nor U474 (N_474,In_681,In_1046);
nand U475 (N_475,In_1732,In_915);
and U476 (N_476,In_154,In_2347);
xnor U477 (N_477,In_757,In_540);
and U478 (N_478,In_2510,In_665);
nor U479 (N_479,In_3705,In_1377);
or U480 (N_480,In_699,In_2892);
or U481 (N_481,In_1270,In_2847);
nor U482 (N_482,In_2825,In_4263);
nand U483 (N_483,In_4088,In_3366);
xnor U484 (N_484,In_1759,In_3574);
or U485 (N_485,In_1045,In_4811);
and U486 (N_486,In_2245,In_773);
nand U487 (N_487,In_1559,In_2108);
nor U488 (N_488,In_3820,In_3232);
nand U489 (N_489,In_3371,In_1202);
nand U490 (N_490,In_842,In_2642);
and U491 (N_491,In_1015,In_233);
xor U492 (N_492,In_1478,In_42);
nand U493 (N_493,In_2842,In_2694);
xor U494 (N_494,In_3203,In_1384);
xor U495 (N_495,In_168,In_3484);
nor U496 (N_496,In_964,In_2925);
or U497 (N_497,In_802,In_3290);
xor U498 (N_498,In_1060,In_2199);
and U499 (N_499,In_4264,In_4190);
xor U500 (N_500,In_435,In_2869);
nor U501 (N_501,In_4784,In_1354);
nand U502 (N_502,In_321,In_4281);
and U503 (N_503,In_1245,In_2267);
or U504 (N_504,In_416,In_3916);
xnor U505 (N_505,In_4552,In_529);
xor U506 (N_506,In_2608,In_3877);
nor U507 (N_507,In_2061,In_43);
xnor U508 (N_508,In_3514,In_2955);
xnor U509 (N_509,In_2611,In_2714);
nand U510 (N_510,In_3293,In_1505);
nor U511 (N_511,In_2068,In_4722);
xor U512 (N_512,In_4063,In_3878);
nand U513 (N_513,In_3424,In_2303);
or U514 (N_514,In_715,In_694);
and U515 (N_515,In_814,In_3585);
nor U516 (N_516,In_4697,In_1637);
nand U517 (N_517,In_3831,In_1869);
nand U518 (N_518,In_1730,In_15);
nor U519 (N_519,In_575,In_4582);
or U520 (N_520,In_610,In_4753);
nor U521 (N_521,In_4159,In_4726);
xnor U522 (N_522,In_3935,In_1476);
nor U523 (N_523,In_979,In_3212);
nand U524 (N_524,In_3553,In_1336);
nor U525 (N_525,In_2207,In_3467);
nor U526 (N_526,In_4011,In_2166);
nor U527 (N_527,In_1089,In_402);
and U528 (N_528,In_3179,In_2630);
nand U529 (N_529,In_1185,In_488);
nor U530 (N_530,In_4902,In_4788);
xor U531 (N_531,In_4187,In_925);
nor U532 (N_532,In_389,In_3628);
or U533 (N_533,In_319,In_744);
nand U534 (N_534,In_2494,In_1671);
xnor U535 (N_535,In_4797,In_3441);
and U536 (N_536,In_2889,In_1837);
nand U537 (N_537,In_4237,In_1343);
nor U538 (N_538,In_4934,In_1721);
and U539 (N_539,In_3169,In_3523);
xnor U540 (N_540,In_138,In_1443);
xnor U541 (N_541,In_739,In_3959);
xor U542 (N_542,In_4860,In_4508);
nor U543 (N_543,In_4120,In_3612);
and U544 (N_544,In_2956,In_4064);
or U545 (N_545,In_2354,In_1477);
xor U546 (N_546,In_4909,In_4896);
nor U547 (N_547,In_2328,In_686);
nand U548 (N_548,In_4471,In_2243);
and U549 (N_549,In_4745,In_2271);
nor U550 (N_550,In_3572,In_3897);
and U551 (N_551,In_1746,In_1415);
xor U552 (N_552,In_3898,In_3522);
and U553 (N_553,In_335,In_3996);
nor U554 (N_554,In_1341,In_4093);
nor U555 (N_555,In_2833,In_4132);
nor U556 (N_556,In_177,In_353);
or U557 (N_557,In_1736,In_2233);
and U558 (N_558,In_128,In_4261);
and U559 (N_559,In_4186,In_1969);
nor U560 (N_560,In_309,In_2124);
or U561 (N_561,In_2594,In_3140);
nor U562 (N_562,In_506,In_3655);
nor U563 (N_563,In_4043,In_4369);
nand U564 (N_564,In_4665,In_3271);
or U565 (N_565,In_3402,In_1751);
or U566 (N_566,In_315,In_4543);
and U567 (N_567,In_3111,In_4514);
and U568 (N_568,In_3095,In_2568);
or U569 (N_569,In_3806,In_4610);
nand U570 (N_570,In_1276,In_1865);
xor U571 (N_571,In_2403,In_2184);
nand U572 (N_572,In_1538,In_4814);
nor U573 (N_573,In_3689,In_2416);
or U574 (N_574,In_1283,In_826);
xor U575 (N_575,In_4611,In_2957);
nand U576 (N_576,In_2744,In_4333);
nor U577 (N_577,In_1799,In_2785);
or U578 (N_578,In_1533,In_1097);
nor U579 (N_579,In_859,In_1951);
or U580 (N_580,In_4614,In_4729);
nand U581 (N_581,In_4250,In_2534);
or U582 (N_582,In_3024,In_4870);
xor U583 (N_583,In_144,In_593);
or U584 (N_584,In_4104,In_4331);
or U585 (N_585,In_3588,In_724);
and U586 (N_586,In_746,In_1974);
xnor U587 (N_587,In_3086,In_208);
or U588 (N_588,In_2294,In_725);
nor U589 (N_589,In_1864,In_1116);
nor U590 (N_590,In_3810,In_3215);
xnor U591 (N_591,In_2085,In_1312);
nor U592 (N_592,In_500,In_2315);
or U593 (N_593,In_4604,In_212);
and U594 (N_594,In_819,In_1595);
or U595 (N_595,In_3970,In_223);
xnor U596 (N_596,In_1769,In_188);
or U597 (N_597,In_2598,In_3943);
or U598 (N_598,In_4714,In_1181);
and U599 (N_599,In_4091,In_973);
or U600 (N_600,In_3739,In_856);
or U601 (N_601,In_2990,In_1504);
and U602 (N_602,In_1030,In_3728);
or U603 (N_603,In_2194,In_3428);
and U604 (N_604,In_2784,In_3247);
nor U605 (N_605,In_4718,In_441);
nand U606 (N_606,In_1306,In_3319);
nand U607 (N_607,In_591,In_2726);
and U608 (N_608,In_578,In_3904);
nor U609 (N_609,In_3172,In_1889);
nand U610 (N_610,In_4716,In_3457);
or U611 (N_611,In_4129,In_3685);
nand U612 (N_612,In_1209,In_3435);
or U613 (N_613,In_1262,In_627);
nor U614 (N_614,In_4832,In_1747);
and U615 (N_615,In_2217,In_3617);
or U616 (N_616,In_1971,In_4033);
or U617 (N_617,In_1105,In_229);
and U618 (N_618,In_2959,In_2141);
xnor U619 (N_619,In_2380,In_4290);
or U620 (N_620,In_4757,In_806);
nand U621 (N_621,In_2498,In_698);
nand U622 (N_622,In_1597,In_2523);
xnor U623 (N_623,In_4969,In_493);
nor U624 (N_624,In_2143,In_3031);
xnor U625 (N_625,In_3866,In_3076);
nor U626 (N_626,In_1464,In_1717);
or U627 (N_627,In_4865,In_2765);
and U628 (N_628,In_1786,In_4950);
nand U629 (N_629,In_650,In_3880);
xor U630 (N_630,In_1288,In_4664);
xor U631 (N_631,In_4110,In_1947);
xor U632 (N_632,In_1575,In_122);
nor U633 (N_633,In_2624,In_1512);
nor U634 (N_634,In_3353,In_293);
nand U635 (N_635,In_3464,In_2162);
nor U636 (N_636,In_3798,In_3150);
and U637 (N_637,In_2741,In_4173);
nor U638 (N_638,In_2723,In_3869);
or U639 (N_639,In_4771,In_2029);
nor U640 (N_640,In_1579,In_3944);
nor U641 (N_641,In_4485,In_3840);
xor U642 (N_642,In_4571,In_833);
nor U643 (N_643,In_2074,In_1395);
and U644 (N_644,In_4422,In_4819);
nor U645 (N_645,In_3852,In_4446);
and U646 (N_646,In_267,In_2125);
or U647 (N_647,In_844,In_4556);
nand U648 (N_648,In_3665,In_4506);
and U649 (N_649,In_3176,In_2397);
or U650 (N_650,In_4070,In_1268);
nor U651 (N_651,In_261,In_3083);
nor U652 (N_652,In_504,In_3950);
xor U653 (N_653,In_619,In_4966);
nor U654 (N_654,In_2711,In_1427);
nand U655 (N_655,In_2017,In_2110);
or U656 (N_656,In_3838,In_1672);
xnor U657 (N_657,In_2164,In_3166);
and U658 (N_658,In_4166,In_1139);
and U659 (N_659,In_4743,In_3216);
xnor U660 (N_660,In_2188,In_594);
or U661 (N_661,In_240,In_2923);
nand U662 (N_662,In_439,In_1489);
xor U663 (N_663,In_2675,In_1187);
or U664 (N_664,In_1027,In_3627);
or U665 (N_665,In_1501,In_2251);
nor U666 (N_666,In_4026,In_1772);
and U667 (N_667,In_656,In_4470);
nor U668 (N_668,In_2958,In_922);
nor U669 (N_669,In_4728,In_3551);
or U670 (N_670,In_4646,In_1099);
nand U671 (N_671,In_2415,In_1029);
nand U672 (N_672,In_3565,In_1368);
nor U673 (N_673,In_382,In_4957);
and U674 (N_674,In_1955,In_957);
xnor U675 (N_675,In_3121,In_944);
nor U676 (N_676,In_387,In_3046);
and U677 (N_677,In_4039,In_1071);
and U678 (N_678,In_4640,In_1643);
or U679 (N_679,In_4500,In_1537);
and U680 (N_680,In_1564,In_4597);
nor U681 (N_681,In_1190,In_453);
and U682 (N_682,In_4406,In_1657);
and U683 (N_683,In_2996,In_510);
nor U684 (N_684,In_630,In_1560);
nor U685 (N_685,In_4442,In_4046);
nand U686 (N_686,In_4427,In_3938);
nand U687 (N_687,In_1711,In_3931);
or U688 (N_688,In_98,In_2321);
or U689 (N_689,In_320,In_4320);
xnor U690 (N_690,In_3903,In_190);
and U691 (N_691,In_3980,In_2040);
and U692 (N_692,In_4505,In_329);
nor U693 (N_693,In_4710,In_4366);
nor U694 (N_694,In_2700,In_684);
or U695 (N_695,In_2820,In_993);
nor U696 (N_696,In_2161,In_4195);
xor U697 (N_697,In_620,In_3581);
or U698 (N_698,In_371,In_567);
nor U699 (N_699,In_4917,In_301);
nor U700 (N_700,In_1701,In_2739);
nor U701 (N_701,In_1925,In_2445);
xor U702 (N_702,In_1796,In_4393);
or U703 (N_703,In_3595,In_4881);
xor U704 (N_704,In_517,In_290);
nor U705 (N_705,In_507,In_3928);
xor U706 (N_706,In_1457,In_4293);
nor U707 (N_707,In_1918,In_4848);
nor U708 (N_708,In_1766,In_692);
nand U709 (N_709,In_4507,In_2254);
xor U710 (N_710,In_114,In_102);
xor U711 (N_711,In_3607,In_2504);
nand U712 (N_712,In_4107,In_1121);
or U713 (N_713,In_2156,In_2180);
xor U714 (N_714,In_3870,In_3308);
nand U715 (N_715,In_4503,In_2308);
nand U716 (N_716,In_3797,In_2117);
nand U717 (N_717,In_4036,In_38);
nand U718 (N_718,In_3555,In_4650);
nor U719 (N_719,In_707,In_3438);
or U720 (N_720,In_3951,In_1363);
or U721 (N_721,In_9,In_2365);
nor U722 (N_722,In_3369,In_76);
or U723 (N_723,In_845,In_1720);
nor U724 (N_724,In_2986,In_1580);
nor U725 (N_725,In_1979,In_1212);
xnor U726 (N_726,In_2492,In_312);
or U727 (N_727,In_4246,In_1358);
nand U728 (N_728,In_2092,In_4915);
and U729 (N_729,In_2962,In_4287);
nand U730 (N_730,In_1434,In_3128);
or U731 (N_731,In_3188,In_4024);
nor U732 (N_732,In_4509,In_1210);
or U733 (N_733,In_4914,In_793);
and U734 (N_734,In_1607,In_4032);
nor U735 (N_735,In_3018,In_4068);
nand U736 (N_736,In_2890,In_252);
nor U737 (N_737,In_865,In_183);
xnor U738 (N_738,In_3664,In_2189);
nand U739 (N_739,In_4078,In_3154);
nor U740 (N_740,In_704,In_2436);
nand U741 (N_741,In_1755,In_847);
and U742 (N_742,In_1076,In_3699);
and U743 (N_743,In_331,In_3757);
nand U744 (N_744,In_1987,In_4750);
nand U745 (N_745,In_48,In_2645);
nand U746 (N_746,In_755,In_2390);
and U747 (N_747,In_2148,In_3857);
xnor U748 (N_748,In_1059,In_555);
or U749 (N_749,In_4185,In_1021);
nand U750 (N_750,In_3989,In_4538);
xnor U751 (N_751,In_498,In_3043);
xor U752 (N_752,In_358,In_798);
nor U753 (N_753,In_2224,In_2476);
xor U754 (N_754,In_2948,In_1518);
xnor U755 (N_755,In_4631,In_841);
nand U756 (N_756,In_2951,In_4922);
xnor U757 (N_757,In_946,In_4874);
nor U758 (N_758,In_1213,In_167);
and U759 (N_759,In_1229,In_4215);
nand U760 (N_760,In_1274,In_4303);
nor U761 (N_761,In_917,In_1758);
or U762 (N_762,In_227,In_2733);
or U763 (N_763,In_1998,In_1396);
xor U764 (N_764,In_417,In_4244);
xor U765 (N_765,In_799,In_198);
and U766 (N_766,In_3224,In_1961);
and U767 (N_767,In_3331,In_4338);
or U768 (N_768,In_3073,In_2871);
or U769 (N_769,In_67,In_3632);
or U770 (N_770,In_2982,In_4759);
xnor U771 (N_771,In_1884,In_4644);
xor U772 (N_772,In_2503,In_401);
or U773 (N_773,In_1361,In_1571);
nand U774 (N_774,In_3965,In_481);
or U775 (N_775,In_3001,In_4038);
nor U776 (N_776,In_3582,In_3275);
xor U777 (N_777,In_1618,In_3248);
xor U778 (N_778,In_2461,In_603);
and U779 (N_779,In_215,In_1269);
xor U780 (N_780,In_3506,In_4408);
xnor U781 (N_781,In_4648,In_1115);
nor U782 (N_782,In_2556,In_456);
xnor U783 (N_783,In_3819,In_479);
and U784 (N_784,In_4999,In_125);
and U785 (N_785,In_4515,In_2305);
or U786 (N_786,In_1770,In_4150);
or U787 (N_787,In_3990,In_4008);
or U788 (N_788,In_2095,In_4910);
or U789 (N_789,In_4935,In_191);
nor U790 (N_790,In_4821,In_3941);
nor U791 (N_791,In_1520,In_4894);
xor U792 (N_792,In_2708,In_1809);
nor U793 (N_793,In_2122,In_1198);
nand U794 (N_794,In_4939,In_3622);
or U795 (N_795,In_1735,In_412);
nor U796 (N_796,In_4657,In_104);
xor U797 (N_797,In_2639,In_3022);
xor U798 (N_798,In_2060,In_3392);
xor U799 (N_799,In_4102,In_4407);
xnor U800 (N_800,In_2241,In_2425);
and U801 (N_801,In_1870,In_4480);
nor U802 (N_802,In_2039,In_2858);
nor U803 (N_803,In_2950,In_4398);
or U804 (N_804,In_3719,In_30);
and U805 (N_805,In_224,In_238);
or U806 (N_806,In_2567,In_4003);
or U807 (N_807,In_459,In_3302);
or U808 (N_808,In_383,In_1655);
xnor U809 (N_809,In_181,In_3074);
xor U810 (N_810,In_3813,In_3126);
or U811 (N_811,In_1335,In_3751);
nor U812 (N_812,In_3325,In_3774);
nor U813 (N_813,In_3161,In_2914);
nand U814 (N_814,In_1416,In_2586);
nor U815 (N_815,In_636,In_3100);
and U816 (N_816,In_3687,In_1719);
xnor U817 (N_817,In_2359,In_3075);
and U818 (N_818,In_1847,In_3217);
and U819 (N_819,In_941,In_4933);
and U820 (N_820,In_2127,In_492);
nand U821 (N_821,In_2992,In_2918);
nor U822 (N_822,In_4059,In_836);
and U823 (N_823,In_4042,In_2756);
xor U824 (N_824,In_549,In_4854);
or U825 (N_825,In_1355,In_1244);
or U826 (N_826,In_3526,In_4837);
and U827 (N_827,In_4216,In_822);
or U828 (N_828,In_407,In_3876);
and U829 (N_829,In_3210,In_1056);
nand U830 (N_830,In_1956,In_2922);
and U831 (N_831,In_1431,In_4943);
nand U832 (N_832,In_4831,In_1815);
and U833 (N_833,In_1959,In_3170);
and U834 (N_834,In_1950,In_4791);
nor U835 (N_835,In_1320,In_3021);
or U836 (N_836,In_3839,In_884);
or U837 (N_837,In_2863,In_2715);
xor U838 (N_838,In_4286,In_4234);
nor U839 (N_839,In_71,In_1057);
and U840 (N_840,In_2945,In_2132);
or U841 (N_841,In_3142,In_3961);
xnor U842 (N_842,In_3481,In_660);
xor U843 (N_843,In_4439,In_4923);
or U844 (N_844,In_919,In_3357);
nand U845 (N_845,In_3974,In_1805);
or U846 (N_846,In_3338,In_2633);
xnor U847 (N_847,In_218,In_3246);
and U848 (N_848,In_1342,In_4460);
and U849 (N_849,In_86,In_1705);
xnor U850 (N_850,In_2677,In_304);
nor U851 (N_851,In_4591,In_2604);
or U852 (N_852,In_2808,In_2444);
xnor U853 (N_853,In_4883,In_3985);
xor U854 (N_854,In_2596,In_1791);
nand U855 (N_855,In_3456,In_1818);
nor U856 (N_856,In_2540,In_4328);
and U857 (N_857,In_2460,In_3861);
xor U858 (N_858,In_326,In_307);
and U859 (N_859,In_4477,In_3381);
xor U860 (N_860,In_4072,In_3887);
nand U861 (N_861,In_3893,In_413);
or U862 (N_862,In_4676,In_2605);
xor U863 (N_863,In_2282,In_3907);
or U864 (N_864,In_2671,In_3883);
xnor U865 (N_865,In_3068,In_3795);
nand U866 (N_866,In_3058,In_3659);
nor U867 (N_867,In_117,In_909);
or U868 (N_868,In_2939,In_3814);
or U869 (N_869,In_2526,In_4732);
and U870 (N_870,In_3533,In_1945);
or U871 (N_871,In_546,In_4578);
nor U872 (N_872,In_341,In_2096);
xor U873 (N_873,In_103,In_2933);
nor U874 (N_874,In_3087,In_3430);
xor U875 (N_875,In_552,In_3380);
nand U876 (N_876,In_4899,In_1348);
xnor U877 (N_877,In_918,In_3884);
and U878 (N_878,In_4958,In_4690);
and U879 (N_879,In_4484,In_2522);
nor U880 (N_880,In_1892,In_2669);
nand U881 (N_881,In_2089,In_4613);
nand U882 (N_882,In_2260,In_1623);
nand U883 (N_883,In_4084,In_3630);
xor U884 (N_884,In_4947,In_2524);
nand U885 (N_885,In_1638,In_2153);
nor U886 (N_886,In_2582,In_3491);
nand U887 (N_887,In_1640,In_996);
or U888 (N_888,In_2400,In_3336);
nand U889 (N_889,In_2511,In_4765);
nor U890 (N_890,In_1386,In_2247);
xnor U891 (N_891,In_2985,In_2448);
nor U892 (N_892,In_404,In_2187);
nand U893 (N_893,In_4829,In_2248);
or U894 (N_894,In_531,In_1708);
nand U895 (N_895,In_2102,In_992);
nor U896 (N_896,In_3743,In_2176);
nor U897 (N_897,In_1822,In_2574);
nor U898 (N_898,In_2532,In_1525);
or U899 (N_899,In_4001,In_1908);
xor U900 (N_900,In_1016,In_1846);
or U901 (N_901,In_3020,In_642);
nor U902 (N_902,In_888,In_4925);
and U903 (N_903,In_583,In_4362);
xnor U904 (N_904,In_2659,In_325);
or U905 (N_905,In_1906,In_3300);
or U906 (N_906,In_283,In_3930);
and U907 (N_907,In_4977,In_2160);
and U908 (N_908,In_10,In_1433);
and U909 (N_909,In_1500,In_419);
and U910 (N_910,In_1582,In_1860);
or U911 (N_911,In_3997,In_3028);
or U912 (N_912,In_2393,In_795);
or U913 (N_913,In_173,In_3644);
nor U914 (N_914,In_2967,In_3785);
xor U915 (N_915,In_1227,In_199);
xor U916 (N_916,In_3763,In_471);
and U917 (N_917,In_3808,In_4717);
nand U918 (N_918,In_2766,In_324);
or U919 (N_919,In_4151,In_489);
xnor U920 (N_920,In_4,In_2500);
nand U921 (N_921,In_3771,In_3242);
or U922 (N_922,In_1347,In_2519);
and U923 (N_923,In_1321,In_2548);
nand U924 (N_924,In_3503,In_1968);
nor U925 (N_925,In_637,In_1615);
nand U926 (N_926,In_2879,In_1965);
or U927 (N_927,In_1782,In_3311);
or U928 (N_928,In_178,In_2660);
xor U929 (N_929,In_106,In_3439);
nor U930 (N_930,In_536,In_4006);
or U931 (N_931,In_4655,In_1221);
xor U932 (N_932,In_2213,In_3370);
and U933 (N_933,In_1997,In_2793);
nor U934 (N_934,In_332,In_2776);
nand U935 (N_935,In_3220,In_2803);
nand U936 (N_936,In_4074,In_1040);
nand U937 (N_937,In_4594,In_586);
xnor U938 (N_938,In_79,In_362);
nor U939 (N_939,In_1685,In_1172);
nand U940 (N_940,In_1328,In_2750);
and U941 (N_941,In_4535,In_3855);
or U942 (N_942,In_2762,In_2868);
and U943 (N_943,In_2727,In_4146);
nand U944 (N_944,In_2852,In_3416);
nand U945 (N_945,In_2364,In_1038);
and U946 (N_946,In_465,In_2455);
xor U947 (N_947,In_2472,In_1785);
nor U948 (N_948,In_1259,In_2088);
or U949 (N_949,In_879,In_2584);
or U950 (N_950,In_3954,In_2007);
nand U951 (N_951,In_1290,In_1191);
nor U952 (N_952,In_1254,In_2706);
nand U953 (N_953,In_2059,In_1495);
xnor U954 (N_954,In_4343,In_3695);
or U955 (N_955,In_1077,In_1);
xnor U956 (N_956,In_2730,In_3638);
nand U957 (N_957,In_2066,In_219);
and U958 (N_958,In_1709,In_3362);
xnor U959 (N_959,In_70,In_1529);
nor U960 (N_960,In_2262,In_1365);
nor U961 (N_961,In_3610,In_3504);
nand U962 (N_962,In_3721,In_2065);
and U963 (N_963,In_3697,In_3986);
nand U964 (N_964,In_2142,In_2897);
and U965 (N_965,In_63,In_4684);
nor U966 (N_966,In_2558,In_351);
and U967 (N_967,In_1994,In_3139);
or U968 (N_968,In_3397,In_2323);
nand U969 (N_969,In_3056,In_763);
xor U970 (N_970,In_4606,In_1924);
and U971 (N_971,In_2617,In_3732);
nor U972 (N_972,In_4579,In_4421);
and U973 (N_973,In_1370,In_680);
nand U974 (N_974,In_1756,In_1402);
nor U975 (N_975,In_1078,In_3296);
and U976 (N_976,In_3837,In_2631);
nor U977 (N_977,In_2771,In_1120);
and U978 (N_978,In_4111,In_820);
xor U979 (N_979,In_2477,In_4420);
nor U980 (N_980,In_3418,In_1652);
nand U981 (N_981,In_4034,In_2064);
nand U982 (N_982,In_4090,In_509);
xnor U983 (N_983,In_2705,In_3376);
or U984 (N_984,In_3871,In_4278);
nand U985 (N_985,In_3334,In_693);
or U986 (N_986,In_318,In_4577);
or U987 (N_987,In_4071,In_616);
xor U988 (N_988,In_2854,In_1775);
and U989 (N_989,In_3368,In_237);
nor U990 (N_990,In_4209,In_1683);
nand U991 (N_991,In_4031,In_1527);
nor U992 (N_992,In_254,In_3030);
nand U993 (N_993,In_1546,In_4987);
xor U994 (N_994,In_1260,In_4617);
nor U995 (N_995,In_1608,In_2782);
or U996 (N_996,In_3408,In_4539);
or U997 (N_997,In_3977,In_3080);
nor U998 (N_998,In_62,In_4645);
nor U999 (N_999,In_162,In_721);
and U1000 (N_1000,In_1704,In_4478);
or U1001 (N_1001,In_228,In_1299);
xnor U1002 (N_1002,In_1373,In_1885);
nand U1003 (N_1003,In_4961,In_4123);
or U1004 (N_1004,In_31,In_3090);
nand U1005 (N_1005,In_45,In_1243);
nand U1006 (N_1006,In_4880,In_4475);
or U1007 (N_1007,In_4089,In_69);
xnor U1008 (N_1008,In_3477,In_200);
nand U1009 (N_1009,In_3328,In_1750);
nor U1010 (N_1010,In_3896,In_1188);
nand U1011 (N_1011,In_4491,In_521);
nor U1012 (N_1012,In_1317,In_2779);
nor U1013 (N_1013,In_3900,In_2620);
xnor U1014 (N_1014,In_997,In_1962);
and U1015 (N_1015,In_4455,In_400);
or U1016 (N_1016,In_4260,In_1155);
xor U1017 (N_1017,In_2179,In_3053);
and U1018 (N_1018,In_1073,In_463);
nor U1019 (N_1019,In_2486,In_2790);
or U1020 (N_1020,In_2887,In_2575);
nor U1021 (N_1021,In_873,In_1617);
and U1022 (N_1022,In_1203,In_2411);
and U1023 (N_1023,In_163,In_2159);
nand U1024 (N_1024,In_3301,In_1983);
nand U1025 (N_1025,In_3265,In_1379);
nor U1026 (N_1026,In_1603,In_1485);
or U1027 (N_1027,In_3395,In_1168);
xor U1028 (N_1028,In_1310,In_3517);
nor U1029 (N_1029,In_2385,In_2442);
or U1030 (N_1030,In_4122,In_4228);
nand U1031 (N_1031,In_1630,In_2541);
xnor U1032 (N_1032,In_4181,In_2297);
or U1033 (N_1033,In_204,In_1048);
and U1034 (N_1034,In_2792,In_4576);
or U1035 (N_1035,In_3065,In_1854);
or U1036 (N_1036,In_4428,In_1586);
or U1037 (N_1037,In_1642,In_2336);
xor U1038 (N_1038,In_3691,In_3156);
nand U1039 (N_1039,In_4411,In_1882);
and U1040 (N_1040,In_4469,In_3492);
nor U1041 (N_1041,In_4144,In_3844);
or U1042 (N_1042,In_2489,In_3914);
or U1043 (N_1043,In_687,In_220);
xor U1044 (N_1044,In_786,In_2894);
nor U1045 (N_1045,In_372,In_4898);
and U1046 (N_1046,In_484,In_34);
nor U1047 (N_1047,In_4344,In_2849);
and U1048 (N_1048,In_149,In_1986);
and U1049 (N_1049,In_1859,In_2000);
xnor U1050 (N_1050,In_3423,In_2937);
xnor U1051 (N_1051,In_2860,In_1783);
xor U1052 (N_1052,In_2028,In_4196);
nand U1053 (N_1053,In_2697,In_1700);
nor U1054 (N_1054,In_2404,In_3276);
xor U1055 (N_1055,In_2995,In_2198);
nand U1056 (N_1056,In_1393,In_860);
xnor U1057 (N_1057,In_1914,In_4687);
or U1058 (N_1058,In_8,In_495);
and U1059 (N_1059,In_2479,In_1737);
nor U1060 (N_1060,In_2054,In_1376);
nand U1061 (N_1061,In_4095,In_4519);
nand U1062 (N_1062,In_3597,In_398);
nor U1063 (N_1063,In_3511,In_3886);
or U1064 (N_1064,In_3274,In_472);
xor U1065 (N_1065,In_3143,In_3599);
or U1066 (N_1066,In_1372,In_96);
nor U1067 (N_1067,In_1091,In_3062);
xor U1068 (N_1068,In_628,In_359);
xnor U1069 (N_1069,In_1422,In_1419);
or U1070 (N_1070,In_2767,In_2546);
and U1071 (N_1071,In_1070,In_84);
and U1072 (N_1072,In_3364,In_105);
nand U1073 (N_1073,In_3614,In_4372);
or U1074 (N_1074,In_4768,In_310);
or U1075 (N_1075,In_4700,In_3039);
nand U1076 (N_1076,In_664,In_3487);
and U1077 (N_1077,In_1063,In_3918);
nand U1078 (N_1078,In_4705,In_3459);
xor U1079 (N_1079,In_288,In_3672);
or U1080 (N_1080,In_3208,In_235);
nand U1081 (N_1081,In_2602,In_866);
nor U1082 (N_1082,In_4887,In_3921);
nand U1083 (N_1083,In_4377,In_4323);
nor U1084 (N_1084,In_3834,In_1250);
nand U1085 (N_1085,In_1003,In_3173);
xor U1086 (N_1086,In_4202,In_2220);
xnor U1087 (N_1087,In_3266,In_1136);
and U1088 (N_1088,In_3580,In_3322);
nand U1089 (N_1089,In_197,In_1825);
or U1090 (N_1090,In_4628,In_3450);
nand U1091 (N_1091,In_2286,In_1196);
nor U1092 (N_1092,In_1095,In_2799);
nand U1093 (N_1093,In_1173,In_3577);
nand U1094 (N_1094,In_1578,In_3476);
xnor U1095 (N_1095,In_4605,In_4827);
or U1096 (N_1096,In_4412,In_1780);
nand U1097 (N_1097,In_4998,In_742);
nand U1098 (N_1098,In_1179,In_758);
or U1099 (N_1099,In_409,In_3545);
nand U1100 (N_1100,In_2753,In_3163);
or U1101 (N_1101,In_1156,In_4240);
xor U1102 (N_1102,In_4174,In_3092);
and U1103 (N_1103,In_4448,In_962);
and U1104 (N_1104,In_1258,In_2111);
xor U1105 (N_1105,In_2268,In_3983);
and U1106 (N_1106,In_2968,In_385);
nor U1107 (N_1107,In_951,In_2566);
or U1108 (N_1108,In_3645,In_4267);
and U1109 (N_1109,In_4379,In_3199);
and U1110 (N_1110,In_3105,In_476);
xnor U1111 (N_1111,In_959,In_2031);
or U1112 (N_1112,In_3740,In_4097);
and U1113 (N_1113,In_2898,In_3735);
xnor U1114 (N_1114,In_1327,In_1909);
nand U1115 (N_1115,In_4997,In_1634);
xor U1116 (N_1116,In_1676,In_4524);
or U1117 (N_1117,In_2376,In_1403);
nand U1118 (N_1118,In_1692,In_748);
nand U1119 (N_1119,In_3901,In_4053);
and U1120 (N_1120,In_3256,In_3827);
nand U1121 (N_1121,In_894,In_808);
or U1122 (N_1122,In_4900,In_652);
and U1123 (N_1123,In_903,In_892);
or U1124 (N_1124,In_347,In_4995);
or U1125 (N_1125,In_1874,In_2026);
and U1126 (N_1126,In_874,In_57);
or U1127 (N_1127,In_657,In_2988);
nand U1128 (N_1128,In_3608,In_3194);
and U1129 (N_1129,In_1096,In_4441);
xor U1130 (N_1130,In_1599,In_1904);
or U1131 (N_1131,In_4276,In_61);
xor U1132 (N_1132,In_1410,In_2509);
nand U1133 (N_1133,In_4279,In_4553);
nand U1134 (N_1134,In_16,In_1344);
xnor U1135 (N_1135,In_4353,In_3350);
and U1136 (N_1136,In_3473,In_1977);
and U1137 (N_1137,In_545,In_1828);
nand U1138 (N_1138,In_2830,In_972);
nor U1139 (N_1139,In_3875,In_1910);
nand U1140 (N_1140,In_4760,In_2555);
nand U1141 (N_1141,In_2678,In_3513);
xor U1142 (N_1142,In_977,In_4213);
and U1143 (N_1143,In_3663,In_851);
or U1144 (N_1144,In_4367,In_4028);
and U1145 (N_1145,In_1086,In_2106);
xor U1146 (N_1146,In_3340,In_3724);
xor U1147 (N_1147,In_2137,In_4259);
nand U1148 (N_1148,In_1967,In_3234);
or U1149 (N_1149,In_749,In_643);
nor U1150 (N_1150,In_1871,In_2084);
or U1151 (N_1151,In_1389,In_1879);
or U1152 (N_1152,In_3908,In_2701);
xor U1153 (N_1153,In_1087,In_2834);
nand U1154 (N_1154,In_2136,In_3181);
nor U1155 (N_1155,In_44,In_961);
nor U1156 (N_1156,In_2258,In_3315);
or U1157 (N_1157,In_4545,In_1519);
xor U1158 (N_1158,In_1182,In_158);
nand U1159 (N_1159,In_1688,In_4054);
nor U1160 (N_1160,In_22,In_4081);
xnor U1161 (N_1161,In_639,In_1594);
or U1162 (N_1162,In_3648,In_2810);
xor U1163 (N_1163,In_176,In_1439);
nor U1164 (N_1164,In_1264,In_1315);
nor U1165 (N_1165,In_3152,In_1689);
xnor U1166 (N_1166,In_3850,In_929);
nand U1167 (N_1167,In_2672,In_2052);
nand U1168 (N_1168,In_2018,In_2831);
and U1169 (N_1169,In_4121,In_4678);
or U1170 (N_1170,In_1163,In_3934);
or U1171 (N_1171,In_4194,In_2181);
and U1172 (N_1172,In_4681,In_3495);
xnor U1173 (N_1173,In_3104,In_3123);
or U1174 (N_1174,In_3889,In_1984);
and U1175 (N_1175,In_1104,In_4809);
xnor U1176 (N_1176,In_1189,In_1561);
xor U1177 (N_1177,In_2839,In_4143);
or U1178 (N_1178,In_998,In_2885);
nor U1179 (N_1179,In_4252,In_4327);
and U1180 (N_1180,In_196,In_4975);
nor U1181 (N_1181,In_954,In_803);
nand U1182 (N_1182,In_1843,In_4557);
and U1183 (N_1183,In_914,In_3260);
and U1184 (N_1184,In_217,In_2545);
nand U1185 (N_1185,In_99,In_4405);
nand U1186 (N_1186,In_3186,In_4706);
and U1187 (N_1187,In_1108,In_4504);
and U1188 (N_1188,In_807,In_4560);
nand U1189 (N_1189,In_1821,In_4563);
and U1190 (N_1190,In_647,In_2447);
or U1191 (N_1191,In_2087,In_3415);
or U1192 (N_1192,In_1204,In_3399);
or U1193 (N_1193,In_2920,In_2150);
or U1194 (N_1194,In_4867,In_2070);
and U1195 (N_1195,In_2109,In_3469);
nor U1196 (N_1196,In_4183,In_2071);
or U1197 (N_1197,In_278,In_4840);
and U1198 (N_1198,In_120,In_3417);
or U1199 (N_1199,In_2306,In_2140);
or U1200 (N_1200,In_4592,In_3158);
and U1201 (N_1201,In_4739,In_28);
or U1202 (N_1202,In_2050,In_1661);
xor U1203 (N_1203,In_3853,In_1367);
and U1204 (N_1204,In_2097,In_65);
and U1205 (N_1205,In_3948,In_4688);
xnor U1206 (N_1206,In_4833,In_4295);
xor U1207 (N_1207,In_2368,In_4434);
nand U1208 (N_1208,In_4790,In_4823);
xnor U1209 (N_1209,In_2812,In_2844);
and U1210 (N_1210,In_4587,In_3978);
nand U1211 (N_1211,In_1829,In_1441);
and U1212 (N_1212,In_3048,In_1133);
or U1213 (N_1213,In_1810,In_1764);
nand U1214 (N_1214,In_2433,In_2320);
xnor U1215 (N_1215,In_1285,In_3761);
and U1216 (N_1216,In_3282,In_4890);
nor U1217 (N_1217,In_3227,In_4126);
nor U1218 (N_1218,In_1928,In_3445);
nor U1219 (N_1219,In_2083,In_3081);
xor U1220 (N_1220,In_667,In_3003);
and U1221 (N_1221,In_4288,In_4780);
xnor U1222 (N_1222,In_1232,In_762);
or U1223 (N_1223,In_1085,In_4558);
and U1224 (N_1224,In_4447,In_1901);
and U1225 (N_1225,In_3826,In_3836);
or U1226 (N_1226,In_418,In_3320);
nor U1227 (N_1227,In_4702,In_1137);
nor U1228 (N_1228,In_1226,In_3643);
nor U1229 (N_1229,In_2975,In_1011);
nor U1230 (N_1230,In_1707,In_3576);
or U1231 (N_1231,In_4512,In_3255);
nand U1232 (N_1232,In_2193,In_1549);
nor U1233 (N_1233,In_3631,In_910);
xor U1234 (N_1234,In_920,In_3816);
and U1235 (N_1235,In_3925,In_4849);
xor U1236 (N_1236,In_4467,In_221);
nor U1237 (N_1237,In_4302,In_1392);
and U1238 (N_1238,In_3032,In_2751);
nor U1239 (N_1239,In_4774,In_2867);
or U1240 (N_1240,In_2949,In_3443);
nand U1241 (N_1241,In_4740,In_3874);
xor U1242 (N_1242,In_4099,In_1093);
or U1243 (N_1243,In_4525,In_4919);
nor U1244 (N_1244,In_469,In_2480);
nor U1245 (N_1245,In_2944,In_1715);
nand U1246 (N_1246,In_2388,In_142);
nor U1247 (N_1247,In_3002,In_1174);
nor U1248 (N_1248,In_4671,In_2453);
and U1249 (N_1249,In_3998,In_2128);
nor U1250 (N_1250,In_4023,In_2794);
nand U1251 (N_1251,In_2931,In_4770);
xnor U1252 (N_1252,In_1013,In_2772);
xor U1253 (N_1253,In_4566,In_855);
and U1254 (N_1254,In_754,In_3633);
nor U1255 (N_1255,In_2169,In_2075);
nand U1256 (N_1256,In_3412,In_3651);
and U1257 (N_1257,In_2056,In_2316);
and U1258 (N_1258,In_260,In_1697);
and U1259 (N_1259,In_1930,In_112);
nor U1260 (N_1260,In_1496,In_1677);
nor U1261 (N_1261,In_3707,In_1444);
nor U1262 (N_1262,In_4580,In_3773);
xor U1263 (N_1263,In_3624,In_3769);
xnor U1264 (N_1264,In_1065,In_1031);
or U1265 (N_1265,In_4222,In_1207);
nand U1266 (N_1266,In_3004,In_2027);
and U1267 (N_1267,In_141,In_1178);
and U1268 (N_1268,In_4364,In_4695);
nand U1269 (N_1269,In_1596,In_3571);
and U1270 (N_1270,In_2342,In_601);
or U1271 (N_1271,In_3284,In_611);
and U1272 (N_1272,In_2738,In_1161);
or U1273 (N_1273,In_3879,In_589);
and U1274 (N_1274,In_3444,In_3094);
nor U1275 (N_1275,In_3011,In_1583);
xnor U1276 (N_1276,In_1625,In_468);
nor U1277 (N_1277,In_491,In_4145);
nand U1278 (N_1278,In_2725,In_164);
or U1279 (N_1279,In_912,In_988);
nand U1280 (N_1280,In_1621,In_850);
and U1281 (N_1281,In_3147,In_2802);
nor U1282 (N_1282,In_2020,In_4891);
or U1283 (N_1283,In_895,In_2360);
xor U1284 (N_1284,In_4962,In_216);
or U1285 (N_1285,In_2130,In_1915);
or U1286 (N_1286,In_1724,In_2536);
xor U1287 (N_1287,In_394,In_2022);
nor U1288 (N_1288,In_564,In_1629);
or U1289 (N_1289,In_2091,In_4682);
xor U1290 (N_1290,In_3196,In_1481);
and U1291 (N_1291,In_4607,In_1445);
nand U1292 (N_1292,In_4996,In_4251);
or U1293 (N_1293,In_691,In_4000);
nand U1294 (N_1294,In_17,In_2651);
nand U1295 (N_1295,In_2319,In_2301);
nor U1296 (N_1296,In_2435,In_1200);
xnor U1297 (N_1297,In_1482,In_1993);
xor U1298 (N_1298,In_1600,In_1110);
nor U1299 (N_1299,In_1614,In_1722);
xnor U1300 (N_1300,In_118,In_4656);
and U1301 (N_1301,In_2781,In_3734);
xnor U1302 (N_1302,In_863,In_743);
nand U1303 (N_1303,In_4574,In_4864);
or U1304 (N_1304,In_345,In_4779);
or U1305 (N_1305,In_126,In_1051);
nor U1306 (N_1306,In_1790,In_3706);
nor U1307 (N_1307,In_2668,In_3543);
xnor U1308 (N_1308,In_1543,In_2113);
nand U1309 (N_1309,In_406,In_1411);
nor U1310 (N_1310,In_1252,In_2821);
xor U1311 (N_1311,In_2490,In_2119);
xnor U1312 (N_1312,In_1225,In_4683);
nor U1313 (N_1313,In_2643,In_4828);
xnor U1314 (N_1314,In_3518,In_1797);
xnor U1315 (N_1315,In_2583,In_853);
and U1316 (N_1316,In_1374,In_2991);
or U1317 (N_1317,In_641,In_3786);
or U1318 (N_1318,In_4818,In_2984);
nand U1319 (N_1319,In_2909,In_2381);
or U1320 (N_1320,In_1338,In_2961);
nand U1321 (N_1321,In_4675,In_3149);
nor U1322 (N_1322,In_4055,In_1833);
or U1323 (N_1323,In_2325,In_4017);
or U1324 (N_1324,In_4742,In_1632);
nand U1325 (N_1325,In_723,In_3745);
and U1326 (N_1326,In_4629,In_4370);
xor U1327 (N_1327,In_1069,In_1944);
nor U1328 (N_1328,In_3231,In_376);
and U1329 (N_1329,In_1205,In_3198);
nor U1330 (N_1330,In_2952,In_4802);
xnor U1331 (N_1331,In_4748,In_3285);
xnor U1332 (N_1332,In_4669,In_1545);
nor U1333 (N_1333,In_4127,In_3552);
xnor U1334 (N_1334,In_3304,In_4983);
or U1335 (N_1335,In_3347,In_1921);
nand U1336 (N_1336,In_2030,In_3153);
nand U1337 (N_1337,In_4974,In_3493);
or U1338 (N_1338,In_1429,In_3945);
or U1339 (N_1339,In_1435,In_3859);
nor U1340 (N_1340,In_792,In_245);
nand U1341 (N_1341,In_4241,In_3833);
nor U1342 (N_1342,In_1819,In_949);
or U1343 (N_1343,In_1017,In_501);
xnor U1344 (N_1344,In_2466,In_206);
nand U1345 (N_1345,In_1952,In_512);
and U1346 (N_1346,In_4382,In_3520);
or U1347 (N_1347,In_4315,In_2655);
nor U1348 (N_1348,In_3263,In_1880);
or U1349 (N_1349,In_1043,In_3590);
and U1350 (N_1350,In_303,In_734);
xor U1351 (N_1351,In_4456,In_530);
or U1352 (N_1352,In_4336,In_502);
and U1353 (N_1353,In_3262,In_3570);
or U1354 (N_1354,In_1157,In_3130);
and U1355 (N_1355,In_4612,In_1943);
xnor U1356 (N_1356,In_1214,In_4495);
nand U1357 (N_1357,In_712,In_3569);
nand U1358 (N_1358,In_1241,In_2757);
and U1359 (N_1359,In_74,In_1295);
nand U1360 (N_1360,In_391,In_4473);
nand U1361 (N_1361,In_1407,In_3780);
or U1362 (N_1362,In_838,In_1145);
or U1363 (N_1363,In_1957,In_423);
and U1364 (N_1364,In_1447,In_4291);
or U1365 (N_1365,In_3471,In_2769);
or U1366 (N_1366,In_2569,In_2424);
nand U1367 (N_1367,In_1169,In_945);
xnor U1368 (N_1368,In_4873,In_207);
xor U1369 (N_1369,In_1171,In_4546);
or U1370 (N_1370,In_4727,In_499);
and U1371 (N_1371,In_2165,In_738);
or U1372 (N_1372,In_596,In_3807);
xnor U1373 (N_1373,In_1827,In_4137);
xor U1374 (N_1374,In_3546,In_3524);
nor U1375 (N_1375,In_4882,In_4162);
and U1376 (N_1376,In_4242,In_3298);
and U1377 (N_1377,In_3175,In_1903);
xnor U1378 (N_1378,In_2838,In_4876);
or U1379 (N_1379,In_4365,In_3436);
xor U1380 (N_1380,In_4010,In_1273);
and U1381 (N_1381,In_1954,In_602);
nor U1382 (N_1382,In_2340,In_4355);
nand U1383 (N_1383,In_2683,In_450);
and U1384 (N_1384,In_3245,In_2090);
nand U1385 (N_1385,In_66,In_2815);
xor U1386 (N_1386,In_4157,In_608);
nor U1387 (N_1387,In_4497,In_132);
and U1388 (N_1388,In_3754,In_4735);
nor U1389 (N_1389,In_3872,In_588);
xor U1390 (N_1390,In_1134,In_3618);
nor U1391 (N_1391,In_2353,In_511);
nor U1392 (N_1392,In_4853,In_3228);
nand U1393 (N_1393,In_520,In_1510);
and U1394 (N_1394,In_4029,In_4908);
xnor U1395 (N_1395,In_136,In_334);
nor U1396 (N_1396,In_3137,In_4168);
or U1397 (N_1397,In_1267,In_2976);
nor U1398 (N_1398,In_4699,In_1159);
nor U1399 (N_1399,In_2542,In_1857);
or U1400 (N_1400,In_3972,In_202);
xnor U1401 (N_1401,In_2745,In_2919);
xor U1402 (N_1402,In_3591,In_562);
nor U1403 (N_1403,In_4857,In_3992);
xor U1404 (N_1404,In_4075,In_4993);
and U1405 (N_1405,In_3818,In_429);
or U1406 (N_1406,In_2913,In_674);
or U1407 (N_1407,In_4175,In_2592);
xor U1408 (N_1408,In_911,In_1042);
xnor U1409 (N_1409,In_2209,In_3401);
nor U1410 (N_1410,In_1633,In_3061);
or U1411 (N_1411,In_3716,In_2927);
or U1412 (N_1412,In_1551,In_327);
xor U1413 (N_1413,In_718,In_868);
or U1414 (N_1414,In_3958,In_3383);
nor U1415 (N_1415,In_2024,In_3488);
and U1416 (N_1416,In_4061,In_2001);
xnor U1417 (N_1417,In_870,In_1905);
nor U1418 (N_1418,In_113,In_4443);
and U1419 (N_1419,In_4058,In_1949);
nor U1420 (N_1420,In_425,In_1555);
and U1421 (N_1421,In_1298,In_1491);
nand U1422 (N_1422,In_1409,In_2438);
or U1423 (N_1423,In_4820,In_761);
nor U1424 (N_1424,In_3267,In_3288);
nand U1425 (N_1425,In_828,In_3821);
and U1426 (N_1426,In_1740,In_4087);
nand U1427 (N_1427,In_2550,In_3174);
xor U1428 (N_1428,In_2042,In_1138);
xor U1429 (N_1429,In_2599,In_150);
nand U1430 (N_1430,In_1581,In_4907);
nand U1431 (N_1431,In_2943,In_3586);
xnor U1432 (N_1432,In_3323,In_2259);
nand U1433 (N_1433,In_604,In_2911);
xor U1434 (N_1434,In_2318,In_2135);
or U1435 (N_1435,In_3382,In_1026);
nand U1436 (N_1436,In_3854,In_437);
and U1437 (N_1437,In_2998,In_3427);
nor U1438 (N_1438,In_3393,In_673);
nor U1439 (N_1439,In_551,In_2559);
or U1440 (N_1440,In_2735,In_1530);
nor U1441 (N_1441,In_161,In_3803);
or U1442 (N_1442,In_2036,In_3313);
nand U1443 (N_1443,In_449,In_4452);
or U1444 (N_1444,In_1142,In_3999);
nor U1445 (N_1445,In_928,In_3540);
nand U1446 (N_1446,In_4959,In_2912);
or U1447 (N_1447,In_1400,In_1867);
nor U1448 (N_1448,In_1966,In_1399);
or U1449 (N_1449,In_1049,In_1565);
xor U1450 (N_1450,In_2628,In_3731);
nand U1451 (N_1451,In_1024,In_4638);
nor U1452 (N_1452,In_1436,In_2780);
xor U1453 (N_1453,In_729,In_1438);
or U1454 (N_1454,In_675,In_4830);
and U1455 (N_1455,In_877,In_2773);
or U1456 (N_1456,In_1523,In_2805);
xnor U1457 (N_1457,In_4413,In_3268);
xnor U1458 (N_1458,In_2713,In_542);
nor U1459 (N_1459,In_2147,In_3472);
nor U1460 (N_1460,In_2895,In_3264);
or U1461 (N_1461,In_1936,In_3431);
nor U1462 (N_1462,In_4200,In_298);
nand U1463 (N_1463,In_1462,In_3920);
xor U1464 (N_1464,In_1023,In_3016);
and U1465 (N_1465,In_3125,In_1592);
or U1466 (N_1466,In_4639,In_3442);
nand U1467 (N_1467,In_3926,In_3587);
nor U1468 (N_1468,In_2980,In_4929);
nand U1469 (N_1469,In_1271,In_4285);
and U1470 (N_1470,In_4207,In_346);
nand U1471 (N_1471,In_4310,In_4979);
nor U1472 (N_1472,In_390,In_3044);
or U1473 (N_1473,In_2277,In_3132);
nor U1474 (N_1474,In_2226,In_2214);
and U1475 (N_1475,In_3613,In_23);
xor U1476 (N_1476,In_2876,In_1541);
nand U1477 (N_1477,In_2873,In_4603);
nor U1478 (N_1478,In_2749,In_4967);
nand U1479 (N_1479,In_986,In_1678);
or U1480 (N_1480,In_131,In_2530);
nor U1481 (N_1481,In_1118,In_3968);
xnor U1482 (N_1482,In_2386,In_1610);
nor U1483 (N_1483,In_275,In_4125);
or U1484 (N_1484,In_4711,In_3802);
nor U1485 (N_1485,In_3361,In_677);
xnor U1486 (N_1486,In_3133,In_264);
nand U1487 (N_1487,In_4225,In_3942);
xor U1488 (N_1488,In_2640,In_3233);
or U1489 (N_1489,In_3321,In_140);
and U1490 (N_1490,In_37,In_4282);
and U1491 (N_1491,In_965,In_4521);
nand U1492 (N_1492,In_1627,In_705);
or U1493 (N_1493,In_2934,In_1605);
xor U1494 (N_1494,In_662,In_4486);
or U1495 (N_1495,In_1839,In_4378);
and U1496 (N_1496,In_2502,In_963);
or U1497 (N_1497,In_1484,In_59);
and U1498 (N_1498,In_3768,In_784);
xor U1499 (N_1499,In_1451,In_262);
nor U1500 (N_1500,In_2929,In_2806);
or U1501 (N_1501,In_3749,In_3261);
or U1502 (N_1502,In_4275,In_772);
nor U1503 (N_1503,In_1680,In_3403);
or U1504 (N_1504,In_1508,In_1802);
and U1505 (N_1505,In_1235,In_3394);
nor U1506 (N_1506,In_3116,In_4721);
and U1507 (N_1507,In_1153,In_165);
nor U1508 (N_1508,In_4177,In_2002);
or U1509 (N_1509,In_2798,In_3335);
xnor U1510 (N_1510,In_571,In_4050);
or U1511 (N_1511,In_3815,In_3015);
and U1512 (N_1512,In_1535,In_3164);
and U1513 (N_1513,In_519,In_598);
nand U1514 (N_1514,In_2966,In_2470);
and U1515 (N_1515,In_2926,In_280);
xnor U1516 (N_1516,In_4822,In_4374);
nor U1517 (N_1517,In_2786,In_375);
nand U1518 (N_1518,In_4518,In_434);
nand U1519 (N_1519,In_3971,In_4608);
or U1520 (N_1520,In_1452,In_2118);
nor U1521 (N_1521,In_3758,In_955);
or U1522 (N_1522,In_2561,In_236);
and U1523 (N_1523,In_3654,In_2761);
xor U1524 (N_1524,In_2313,In_291);
and U1525 (N_1525,In_244,In_3911);
nand U1526 (N_1526,In_3200,In_778);
nor U1527 (N_1527,In_2361,In_700);
or U1528 (N_1528,In_1293,In_97);
nor U1529 (N_1529,In_1562,In_2379);
nand U1530 (N_1530,In_3936,In_2231);
and U1531 (N_1531,In_1793,In_1346);
and U1532 (N_1532,In_4273,In_3437);
nand U1533 (N_1533,In_1349,In_3421);
and U1534 (N_1534,In_1875,In_4158);
nand U1535 (N_1535,In_1028,In_1710);
nor U1536 (N_1536,In_2369,In_709);
nor U1537 (N_1537,In_2554,In_380);
nor U1538 (N_1538,In_2232,In_3825);
nand U1539 (N_1539,In_2468,In_482);
nand U1540 (N_1540,In_776,In_587);
nand U1541 (N_1541,In_1333,In_4025);
nand U1542 (N_1542,In_41,In_4499);
and U1543 (N_1543,In_1165,In_4179);
nand U1544 (N_1544,In_4334,In_1357);
xnor U1545 (N_1545,In_135,In_697);
nor U1546 (N_1546,In_861,In_2158);
xor U1547 (N_1547,In_3281,In_843);
xor U1548 (N_1548,In_848,In_3790);
nand U1549 (N_1549,In_3688,In_4012);
xnor U1550 (N_1550,In_2478,In_3700);
nand U1551 (N_1551,In_3312,In_1304);
nand U1552 (N_1552,In_1666,In_2634);
nor U1553 (N_1553,In_4826,In_1613);
xnor U1554 (N_1554,In_1352,In_2537);
or U1555 (N_1555,In_3182,In_4389);
nor U1556 (N_1556,In_4363,In_1811);
or U1557 (N_1557,In_433,In_405);
xor U1558 (N_1558,In_3547,In_4449);
nor U1559 (N_1559,In_947,In_1107);
nand U1560 (N_1560,In_3070,In_2287);
xor U1561 (N_1561,In_2636,In_514);
or U1562 (N_1562,In_3756,In_4764);
or U1563 (N_1563,In_2626,In_1449);
nor U1564 (N_1564,In_3385,In_3270);
nand U1565 (N_1565,In_1787,In_4247);
xnor U1566 (N_1566,In_1929,In_2904);
xnor U1567 (N_1567,In_4782,In_1266);
nor U1568 (N_1568,In_666,In_3358);
nor U1569 (N_1569,In_1456,In_4569);
nand U1570 (N_1570,In_4436,In_313);
and U1571 (N_1571,In_2999,In_3634);
and U1572 (N_1572,In_3167,In_4386);
or U1573 (N_1573,In_1222,In_4130);
and U1574 (N_1574,In_3678,In_214);
nor U1575 (N_1575,In_804,In_2629);
nor U1576 (N_1576,In_1234,In_205);
nor U1577 (N_1577,In_3611,In_1887);
xor U1578 (N_1578,In_2832,In_2427);
or U1579 (N_1579,In_3799,In_752);
nand U1580 (N_1580,In_4666,In_166);
nand U1581 (N_1581,In_3240,In_4796);
or U1582 (N_1582,In_1823,In_862);
nor U1583 (N_1583,In_256,In_2557);
or U1584 (N_1584,In_4453,In_1569);
nand U1585 (N_1585,In_3909,In_1206);
or U1586 (N_1586,In_3867,In_3796);
nor U1587 (N_1587,In_2033,In_3329);
and U1588 (N_1588,In_4633,In_300);
or U1589 (N_1589,In_3059,In_4199);
or U1590 (N_1590,In_4651,In_3106);
and U1591 (N_1591,In_4913,In_867);
nor U1592 (N_1592,In_2037,In_2870);
or U1593 (N_1593,In_4632,In_3733);
nor U1594 (N_1594,In_2212,In_2145);
xnor U1595 (N_1595,In_4458,In_1064);
xnor U1596 (N_1596,In_1845,In_3940);
or U1597 (N_1597,In_2591,In_3804);
and U1598 (N_1598,In_2099,In_3658);
or U1599 (N_1599,In_2508,In_4570);
xnor U1600 (N_1600,In_378,In_4785);
and U1601 (N_1601,In_2200,In_2151);
and U1602 (N_1602,In_3953,In_4048);
xor U1603 (N_1603,In_2389,In_1006);
or U1604 (N_1604,In_2747,In_1726);
and U1605 (N_1605,In_1836,In_609);
nor U1606 (N_1606,In_4667,In_3994);
and U1607 (N_1607,In_741,In_1009);
xor U1608 (N_1608,In_1800,In_561);
or U1609 (N_1609,In_4359,In_1907);
nand U1610 (N_1610,In_3593,In_2481);
nand U1611 (N_1611,In_1432,In_3333);
nor U1612 (N_1612,In_1001,In_4758);
nand U1613 (N_1613,In_3832,In_3932);
nand U1614 (N_1614,In_3629,In_1053);
nor U1615 (N_1615,In_2801,In_2358);
nand U1616 (N_1616,In_1842,In_4931);
or U1617 (N_1617,In_51,In_4658);
and U1618 (N_1618,In_3014,In_3411);
nor U1619 (N_1619,In_2930,In_4384);
nor U1620 (N_1620,In_4674,In_3922);
or U1621 (N_1621,In_210,In_4924);
xor U1622 (N_1622,In_2861,In_1628);
and U1623 (N_1623,In_3515,In_4383);
xnor U1624 (N_1624,In_3993,In_3558);
nand U1625 (N_1625,In_4304,In_3470);
or U1626 (N_1626,In_50,In_3093);
xnor U1627 (N_1627,In_3326,In_4737);
and U1628 (N_1628,In_3598,In_732);
and U1629 (N_1629,In_1807,In_457);
nor U1630 (N_1630,In_3783,In_2841);
and U1631 (N_1631,In_11,In_573);
nand U1632 (N_1632,In_3753,In_2098);
xor U1633 (N_1633,In_1143,In_2965);
xor U1634 (N_1634,In_3303,In_3213);
and U1635 (N_1635,In_1075,In_384);
and U1636 (N_1636,In_1130,In_1897);
or U1637 (N_1637,In_3052,In_4430);
nor U1638 (N_1638,In_722,In_2252);
xnor U1639 (N_1639,In_1223,In_2412);
nor U1640 (N_1640,In_632,In_4755);
nand U1641 (N_1641,In_357,In_4511);
and U1642 (N_1642,In_4652,In_1404);
or U1643 (N_1643,In_1141,In_824);
xnor U1644 (N_1644,In_1995,In_399);
or U1645 (N_1645,In_2387,In_2578);
xor U1646 (N_1646,In_2829,In_1287);
or U1647 (N_1647,In_4746,In_322);
nand U1648 (N_1648,In_3054,In_209);
xor U1649 (N_1649,In_1917,In_180);
xor U1650 (N_1650,In_4461,In_3483);
and U1651 (N_1651,In_539,In_1088);
or U1652 (N_1652,In_952,In_1479);
and U1653 (N_1653,In_3010,In_3830);
nand U1654 (N_1654,In_1542,In_3060);
xor U1655 (N_1655,In_109,In_4329);
nand U1656 (N_1656,In_4296,In_1771);
and U1657 (N_1657,In_3805,In_2439);
nor U1658 (N_1658,In_2053,In_1067);
nor U1659 (N_1659,In_1125,In_2246);
nor U1660 (N_1660,In_1140,In_4800);
or U1661 (N_1661,In_366,In_2458);
nor U1662 (N_1662,In_3191,In_3000);
nor U1663 (N_1663,In_4562,In_3386);
xnor U1664 (N_1664,In_226,In_4944);
xor U1665 (N_1665,In_3962,In_1534);
or U1666 (N_1666,In_4180,In_1978);
nand U1667 (N_1667,In_4808,In_4217);
or U1668 (N_1668,In_2046,In_4903);
xor U1669 (N_1669,In_2035,In_736);
nand U1670 (N_1670,In_2954,In_2278);
nand U1671 (N_1671,In_3434,In_3360);
and U1672 (N_1672,In_1144,In_2612);
xnor U1673 (N_1673,In_2814,In_4253);
nor U1674 (N_1674,In_4741,In_3527);
xor U1675 (N_1675,In_1920,In_2272);
and U1676 (N_1676,In_1119,In_2333);
xor U1677 (N_1677,In_3776,In_323);
xnor U1678 (N_1678,In_4694,In_1832);
or U1679 (N_1679,In_4392,In_379);
and U1680 (N_1680,In_2703,In_4847);
nor U1681 (N_1681,In_646,In_1777);
nor U1682 (N_1682,In_1020,In_1824);
and U1683 (N_1683,In_3112,In_2797);
nor U1684 (N_1684,In_624,In_4609);
and U1685 (N_1685,In_3452,In_4589);
nor U1686 (N_1686,In_813,In_4041);
nor U1687 (N_1687,In_987,In_4464);
xor U1688 (N_1688,In_1835,In_1878);
and U1689 (N_1689,In_1531,In_3057);
and U1690 (N_1690,In_1788,In_2528);
or U1691 (N_1691,In_871,In_2638);
nand U1692 (N_1692,In_2223,In_613);
nand U1693 (N_1693,In_3035,In_1942);
or U1694 (N_1694,In_1729,In_1547);
xnor U1695 (N_1695,In_3131,In_585);
and U1696 (N_1696,In_3118,In_1981);
xnor U1697 (N_1697,In_3973,In_455);
nor U1698 (N_1698,In_883,In_1493);
xnor U1699 (N_1699,In_3616,In_3314);
xor U1700 (N_1700,In_1413,In_1813);
nor U1701 (N_1701,In_2908,In_1382);
and U1702 (N_1702,In_497,In_3160);
xor U1703 (N_1703,In_4156,In_3205);
or U1704 (N_1704,In_2414,In_473);
nand U1705 (N_1705,In_2195,In_3148);
xor U1706 (N_1706,In_3351,In_2538);
nor U1707 (N_1707,In_3766,In_3667);
or U1708 (N_1708,In_1128,In_1004);
and U1709 (N_1709,In_3646,In_2452);
xor U1710 (N_1710,In_3103,In_192);
nor U1711 (N_1711,In_2382,In_4918);
and U1712 (N_1712,In_1664,In_119);
xnor U1713 (N_1713,In_185,In_4047);
xor U1714 (N_1714,In_4219,In_2237);
nor U1715 (N_1715,In_2755,In_2431);
nor U1716 (N_1716,In_1406,In_1175);
nand U1717 (N_1717,In_2647,In_4313);
or U1718 (N_1718,In_4912,In_4211);
xnor U1719 (N_1719,In_3079,In_4920);
nand U1720 (N_1720,In_2329,In_4679);
or U1721 (N_1721,In_2595,In_94);
xnor U1722 (N_1722,In_3653,In_934);
or U1723 (N_1723,In_3505,In_3283);
nand U1724 (N_1724,In_4472,In_1808);
nand U1725 (N_1725,In_2653,In_3292);
or U1726 (N_1726,In_2094,In_3847);
nand U1727 (N_1727,In_234,In_2003);
xor U1728 (N_1728,In_115,In_3447);
xnor U1729 (N_1729,In_3387,In_3946);
nor U1730 (N_1730,In_2129,In_556);
or U1731 (N_1731,In_4960,In_3717);
nand U1732 (N_1732,In_4154,In_1852);
nand U1733 (N_1733,In_2172,In_1972);
nor U1734 (N_1734,In_4863,In_3567);
nor U1735 (N_1735,In_1177,In_719);
or U1736 (N_1736,In_3091,In_4988);
xor U1737 (N_1737,In_1251,In_4311);
nand U1738 (N_1738,In_1731,In_2696);
and U1739 (N_1739,In_3071,In_1278);
xor U1740 (N_1740,In_1694,In_4713);
nand U1741 (N_1741,In_3330,In_791);
nor U1742 (N_1742,In_1742,In_3690);
nand U1743 (N_1743,In_1891,In_2375);
or U1744 (N_1744,In_426,In_2855);
xor U1745 (N_1745,In_3354,In_430);
nand U1746 (N_1746,In_2302,In_3466);
and U1747 (N_1747,In_2383,In_4949);
or U1748 (N_1748,In_4815,In_420);
or U1749 (N_1749,In_787,In_4850);
and U1750 (N_1750,In_2116,In_4192);
and U1751 (N_1751,In_1622,In_2441);
nor U1752 (N_1752,In_1167,In_3310);
or U1753 (N_1753,In_4326,In_1197);
or U1754 (N_1754,In_2464,In_2422);
nor U1755 (N_1755,In_3209,In_3666);
and U1756 (N_1756,In_3019,In_508);
nand U1757 (N_1757,In_1164,In_2973);
nand U1758 (N_1758,In_4206,In_3461);
nor U1759 (N_1759,In_3741,In_4641);
or U1760 (N_1760,In_1765,In_2572);
or U1761 (N_1761,In_4862,In_3738);
nand U1762 (N_1762,In_1194,In_4069);
nand U1763 (N_1763,In_448,In_3675);
or U1764 (N_1764,In_1131,In_2667);
nor U1765 (N_1765,In_4526,In_4858);
or U1766 (N_1766,In_1812,In_2835);
or U1767 (N_1767,In_994,In_4135);
nor U1768 (N_1768,In_1309,In_54);
xor U1769 (N_1769,In_4227,In_2312);
nor U1770 (N_1770,In_2218,In_2589);
nand U1771 (N_1771,In_1820,In_901);
and U1772 (N_1772,In_1816,In_3917);
xor U1773 (N_1773,In_18,In_3097);
xnor U1774 (N_1774,In_659,In_2850);
and U1775 (N_1775,In_4952,In_2310);
or U1776 (N_1776,In_3375,In_902);
or U1777 (N_1777,In_82,In_4555);
and U1778 (N_1778,In_1612,In_4789);
or U1779 (N_1779,In_4812,In_4869);
nor U1780 (N_1780,In_3647,In_3888);
nor U1781 (N_1781,In_4325,In_1216);
or U1782 (N_1782,In_4101,In_462);
and U1783 (N_1783,In_605,In_2429);
nand U1784 (N_1784,In_101,In_2115);
nor U1785 (N_1785,In_1899,In_3956);
xnor U1786 (N_1786,In_3556,In_1201);
and U1787 (N_1787,In_3902,In_4118);
or U1788 (N_1788,In_2752,In_3498);
or U1789 (N_1789,In_1391,In_626);
or U1790 (N_1790,In_4138,In_4708);
or U1791 (N_1791,In_1247,In_2691);
and U1792 (N_1792,In_1602,In_4414);
nand U1793 (N_1793,In_751,In_2025);
or U1794 (N_1794,In_444,In_4635);
nor U1795 (N_1795,In_3849,In_3536);
xor U1796 (N_1796,In_3508,In_625);
nor U1797 (N_1797,In_2144,In_2432);
nand U1798 (N_1798,In_3510,In_4266);
nor U1799 (N_1799,In_526,In_485);
xor U1800 (N_1800,In_2391,In_373);
nor U1801 (N_1801,In_809,In_554);
xnor U1802 (N_1802,In_638,In_2112);
or U1803 (N_1803,In_4956,In_3910);
nand U1804 (N_1804,In_534,In_4457);
and U1805 (N_1805,In_3583,In_147);
nor U1806 (N_1806,In_1698,In_3800);
and U1807 (N_1807,In_1162,In_1988);
xnor U1808 (N_1808,In_1084,In_330);
or U1809 (N_1809,In_3197,In_953);
nor U1810 (N_1810,In_4030,In_2269);
nor U1811 (N_1811,In_4451,In_577);
nor U1812 (N_1812,In_3575,In_3969);
and U1813 (N_1813,In_1275,In_1976);
nand U1814 (N_1814,In_3279,In_2256);
nand U1815 (N_1815,In_1894,In_1034);
and U1816 (N_1816,In_1122,In_3829);
nor U1817 (N_1817,In_2525,In_967);
or U1818 (N_1818,In_110,In_1572);
or U1819 (N_1819,In_768,In_1673);
and U1820 (N_1820,In_213,In_3135);
xor U1821 (N_1821,In_328,In_4416);
and U1822 (N_1822,In_2822,In_2644);
nand U1823 (N_1823,In_950,In_3297);
xor U1824 (N_1824,In_1866,In_231);
nand U1825 (N_1825,In_1587,In_137);
nand U1826 (N_1826,In_1893,In_1940);
nor U1827 (N_1827,In_4626,In_2527);
xor U1828 (N_1828,In_1127,In_4308);
nand U1829 (N_1829,In_2588,In_1744);
nand U1830 (N_1830,In_4659,In_3548);
and U1831 (N_1831,In_4618,In_3683);
and U1832 (N_1832,In_90,In_1991);
or U1833 (N_1833,In_1253,In_88);
xnor U1834 (N_1834,In_1567,In_172);
or U1835 (N_1835,In_1923,In_1180);
xor U1836 (N_1836,In_1591,In_4775);
or U1837 (N_1837,In_4964,In_3711);
nand U1838 (N_1838,In_2344,In_3636);
or U1839 (N_1839,In_2734,In_4813);
and U1840 (N_1840,In_4892,In_1896);
or U1841 (N_1841,In_1035,In_4348);
or U1842 (N_1842,In_1307,In_2170);
nor U1843 (N_1843,In_3788,In_2034);
nor U1844 (N_1844,In_4139,In_2499);
or U1845 (N_1845,In_4350,In_374);
and U1846 (N_1846,In_3082,In_276);
nand U1847 (N_1847,In_230,In_4052);
nor U1848 (N_1848,In_2314,In_782);
or U1849 (N_1849,In_3115,In_1246);
and U1850 (N_1850,In_3124,In_4584);
nor U1851 (N_1851,In_2459,In_980);
or U1852 (N_1852,In_3828,In_3085);
nand U1853 (N_1853,In_2311,In_2712);
nand U1854 (N_1854,In_942,In_4792);
xnor U1855 (N_1855,In_829,In_3661);
xnor U1856 (N_1856,In_1935,In_612);
or U1857 (N_1857,In_2367,In_513);
xnor U1858 (N_1858,In_1776,In_2171);
xor U1859 (N_1859,In_3389,In_442);
nand U1860 (N_1860,In_2809,In_1294);
or U1861 (N_1861,In_1506,In_259);
nor U1862 (N_1862,In_2133,In_4361);
nor U1863 (N_1863,In_2076,In_3295);
nor U1864 (N_1864,In_414,In_75);
nand U1865 (N_1865,In_3309,In_2690);
or U1866 (N_1866,In_1573,In_3141);
and U1867 (N_1867,In_817,In_2285);
and U1868 (N_1868,In_599,In_4668);
xor U1869 (N_1869,In_1329,In_976);
nand U1870 (N_1870,In_1609,In_1000);
nand U1871 (N_1871,In_1556,In_19);
nor U1872 (N_1872,In_3684,In_544);
nand U1873 (N_1873,In_4677,In_1461);
nor U1874 (N_1874,In_2946,In_4889);
xnor U1875 (N_1875,In_3801,In_2107);
or U1876 (N_1876,In_1474,In_2878);
xor U1877 (N_1877,In_4842,In_750);
nand U1878 (N_1878,In_4715,In_3178);
or U1879 (N_1879,In_2279,In_4989);
and U1880 (N_1880,In_2650,In_2240);
nor U1881 (N_1881,In_2168,In_733);
and U1882 (N_1882,In_4946,In_805);
xor U1883 (N_1883,In_2355,In_247);
or U1884 (N_1884,In_708,In_3760);
and U1885 (N_1885,In_1279,In_95);
nand U1886 (N_1886,In_740,In_1693);
and U1887 (N_1887,In_4340,In_1913);
and U1888 (N_1888,In_422,In_696);
nand U1889 (N_1889,In_2940,In_3084);
and U1890 (N_1890,In_3465,In_4394);
and U1891 (N_1891,In_4375,In_1848);
nand U1892 (N_1892,In_3316,In_1149);
or U1893 (N_1893,In_1281,In_3479);
nor U1894 (N_1894,In_2693,In_4926);
xor U1895 (N_1895,In_3578,In_4781);
nand U1896 (N_1896,In_839,In_1639);
and U1897 (N_1897,In_2989,In_3489);
or U1898 (N_1898,In_781,In_683);
xnor U1899 (N_1899,In_4490,In_672);
nor U1900 (N_1900,In_2641,In_3984);
or U1901 (N_1901,In_255,In_4178);
nor U1902 (N_1902,In_4316,In_671);
xnor U1903 (N_1903,In_4201,In_2775);
xnor U1904 (N_1904,In_3356,In_2770);
or U1905 (N_1905,In_654,In_4945);
or U1906 (N_1906,In_4131,In_2299);
and U1907 (N_1907,In_2407,In_2086);
nand U1908 (N_1908,In_3235,In_3812);
nand U1909 (N_1909,In_4904,In_1316);
or U1910 (N_1910,In_4373,In_3367);
nand U1911 (N_1911,In_3218,In_2462);
nor U1912 (N_1912,In_3939,In_3747);
and U1913 (N_1913,In_2401,In_3960);
nor U1914 (N_1914,In_4418,In_2488);
xor U1915 (N_1915,In_20,In_2729);
nor U1916 (N_1916,In_1102,In_2420);
and U1917 (N_1917,In_3305,In_4300);
and U1918 (N_1918,In_1224,In_4893);
nand U1919 (N_1919,In_1098,In_2276);
or U1920 (N_1920,In_864,In_2882);
nand U1921 (N_1921,In_3964,In_348);
nor U1922 (N_1922,In_3425,In_225);
and U1923 (N_1923,In_4437,In_2899);
xnor U1924 (N_1924,In_3050,In_274);
xnor U1925 (N_1925,In_4051,In_2836);
nand U1926 (N_1926,In_3407,In_1650);
xnor U1927 (N_1927,In_3008,In_4319);
xnor U1928 (N_1928,In_2011,In_2748);
xor U1929 (N_1929,In_4878,In_2300);
nor U1930 (N_1930,In_747,In_1516);
and U1931 (N_1931,In_2622,In_2679);
and U1932 (N_1932,In_923,In_1598);
and U1933 (N_1933,In_194,In_2731);
or U1934 (N_1934,In_3026,In_4147);
xnor U1935 (N_1935,In_1081,In_1817);
xnor U1936 (N_1936,In_569,In_3641);
nand U1937 (N_1937,In_2676,In_3033);
and U1938 (N_1938,In_3355,In_4188);
or U1939 (N_1939,In_2728,In_4985);
or U1940 (N_1940,In_3534,In_3668);
or U1941 (N_1941,In_1883,In_1873);
or U1942 (N_1942,In_897,In_193);
nand U1943 (N_1943,In_1762,In_3709);
nor U1944 (N_1944,In_4662,In_243);
nor U1945 (N_1945,In_1490,In_635);
xnor U1946 (N_1946,In_4347,In_3012);
nor U1947 (N_1947,In_2687,In_368);
and U1948 (N_1948,In_14,In_4689);
nor U1949 (N_1949,In_2019,In_129);
xor U1950 (N_1950,In_2800,In_2356);
xnor U1951 (N_1951,In_2960,In_1364);
nor U1952 (N_1952,In_344,In_2201);
nand U1953 (N_1953,In_3537,In_3318);
xnor U1954 (N_1954,In_4040,In_108);
xor U1955 (N_1955,In_2072,In_3453);
nand U1956 (N_1956,In_249,In_830);
and U1957 (N_1957,In_2471,In_1856);
nor U1958 (N_1958,In_4777,In_857);
nand U1959 (N_1959,In_2928,In_1526);
or U1960 (N_1960,In_4076,In_2392);
xnor U1961 (N_1961,In_4248,In_4885);
or U1962 (N_1962,In_1058,In_4226);
nand U1963 (N_1963,In_4376,In_1106);
nand U1964 (N_1964,In_2699,In_3561);
or U1965 (N_1965,In_2047,In_270);
and U1966 (N_1966,In_3462,In_3145);
and U1967 (N_1967,In_4992,In_1725);
and U1968 (N_1968,In_4583,In_2886);
xor U1969 (N_1969,In_4776,In_796);
and U1970 (N_1970,In_4844,In_1517);
nand U1971 (N_1971,In_4243,In_3250);
nor U1972 (N_1972,In_265,In_4009);
nor U1973 (N_1973,In_2491,In_1487);
or U1974 (N_1974,In_4494,In_3365);
and U1975 (N_1975,In_3146,In_4224);
xor U1976 (N_1976,In_528,In_1753);
nor U1977 (N_1977,In_690,In_263);
nand U1978 (N_1978,In_4172,In_438);
xnor U1979 (N_1979,In_1394,In_446);
nand U1980 (N_1980,In_2921,In_2399);
and U1981 (N_1981,In_349,In_4845);
nor U1982 (N_1982,In_4564,In_1718);
nand U1983 (N_1983,In_3929,In_3915);
nand U1984 (N_1984,In_2139,In_2255);
nand U1985 (N_1985,In_4435,In_584);
and U1986 (N_1986,In_2862,In_232);
nand U1987 (N_1987,In_3873,In_160);
nand U1988 (N_1988,In_26,In_1509);
xnor U1989 (N_1989,In_3891,In_3737);
xnor U1990 (N_1990,In_869,In_3979);
nand U1991 (N_1991,In_1645,In_4356);
or U1992 (N_1992,In_2562,In_1455);
nor U1993 (N_1993,In_4092,In_2564);
xnor U1994 (N_1994,In_1611,In_1132);
or U1995 (N_1995,In_4208,In_1996);
nand U1996 (N_1996,In_3894,In_2516);
nor U1997 (N_1997,In_3765,In_3013);
nor U1998 (N_1998,In_1568,In_2529);
nor U1999 (N_1999,In_3835,In_4272);
nor U2000 (N_2000,N_771,In_2152);
xor U2001 (N_2001,N_1027,N_720);
and U2002 (N_2002,N_509,In_4277);
or U2003 (N_2003,In_1208,N_970);
nor U2004 (N_2004,In_3244,In_4403);
or U2005 (N_2005,In_4752,In_2916);
or U2006 (N_2006,In_3413,N_123);
and U2007 (N_2007,N_192,In_1868);
and U2008 (N_2008,N_790,N_84);
nor U2009 (N_2009,In_1383,N_608);
xnor U2010 (N_2010,In_1061,N_45);
or U2011 (N_2011,N_598,In_4345);
nor U2012 (N_2012,N_796,N_1951);
xnor U2013 (N_2013,N_1556,In_3544);
nand U2014 (N_2014,In_3109,N_1389);
nor U2015 (N_2015,N_1119,In_1862);
nand U2016 (N_2016,N_128,In_1584);
xor U2017 (N_2017,N_993,In_4019);
or U2018 (N_2018,In_21,N_378);
nor U2019 (N_2019,N_404,N_565);
and U2020 (N_2020,N_1272,N_1235);
or U2021 (N_2021,In_2969,In_4077);
or U2022 (N_2022,In_816,In_2896);
or U2023 (N_2023,In_480,In_1195);
and U2024 (N_2024,In_483,In_3);
or U2025 (N_2025,In_3088,In_2351);
or U2026 (N_2026,N_804,N_1464);
nand U2027 (N_2027,N_1686,N_309);
or U2028 (N_2028,N_1010,N_1325);
nand U2029 (N_2029,N_1392,In_3165);
nor U2030 (N_2030,N_1913,In_3550);
and U2031 (N_2031,In_6,N_1538);
nand U2032 (N_2032,N_1608,In_706);
nor U2033 (N_2033,N_1393,N_1061);
nand U2034 (N_2034,N_1720,In_3127);
xnor U2035 (N_2035,In_1660,N_60);
nand U2036 (N_2036,N_1160,N_581);
nor U2037 (N_2037,N_1104,N_924);
nand U2038 (N_2038,N_942,N_748);
or U2039 (N_2039,N_1165,N_353);
and U2040 (N_2040,In_4445,In_4661);
nor U2041 (N_2041,In_3339,In_1863);
and U2042 (N_2042,N_1803,N_1172);
nor U2043 (N_2043,N_171,In_143);
nand U2044 (N_2044,N_97,N_213);
or U2045 (N_2045,N_27,N_1046);
nand U2046 (N_2046,N_613,In_3373);
and U2047 (N_2047,N_840,In_2941);
and U2048 (N_2048,In_4169,In_4268);
or U2049 (N_2049,In_186,N_931);
or U2050 (N_2050,N_573,In_284);
and U2051 (N_2051,N_1096,N_1209);
or U2052 (N_2052,N_979,In_470);
xnor U2053 (N_2053,In_2221,N_1991);
and U2054 (N_2054,N_76,N_645);
or U2055 (N_2055,In_1459,N_1713);
and U2056 (N_2056,N_485,N_569);
nand U2057 (N_2057,N_1531,N_1749);
or U2058 (N_2058,N_1462,N_1865);
xor U2059 (N_2059,In_3824,In_239);
or U2060 (N_2060,In_187,In_2177);
nand U2061 (N_2061,In_2063,N_1730);
nor U2062 (N_2062,N_802,In_157);
xor U2063 (N_2063,N_1792,In_1240);
or U2064 (N_2064,In_4401,N_735);
xnor U2065 (N_2065,In_1932,N_749);
nand U2066 (N_2066,N_1810,N_422);
nor U2067 (N_2067,N_125,In_2484);
xor U2068 (N_2068,N_351,N_1738);
or U2069 (N_2069,N_1582,N_1308);
nor U2070 (N_2070,N_1627,In_1469);
nor U2071 (N_2071,N_693,In_3782);
nand U2072 (N_2072,N_264,N_477);
xnor U2073 (N_2073,N_1727,N_1650);
xnor U2074 (N_2074,N_854,N_499);
xnor U2075 (N_2075,N_1041,N_1860);
nor U2076 (N_2076,N_1361,In_4653);
nor U2077 (N_2077,N_389,N_1336);
xor U2078 (N_2078,In_2758,In_649);
xor U2079 (N_2079,In_4541,N_1549);
xnor U2080 (N_2080,N_917,N_464);
or U2081 (N_2081,N_1431,In_1975);
xor U2082 (N_2082,In_1018,N_397);
xor U2083 (N_2083,N_457,N_867);
nand U2084 (N_2084,In_4007,N_331);
xnor U2085 (N_2085,N_242,In_4115);
nor U2086 (N_2086,In_1589,N_28);
nor U2087 (N_2087,N_103,N_1751);
nor U2088 (N_2088,N_906,N_955);
and U2089 (N_2089,N_956,N_669);
nand U2090 (N_2090,N_1059,N_186);
nor U2091 (N_2091,N_616,N_1523);
nand U2092 (N_2092,N_210,In_846);
xnor U2093 (N_2093,In_3967,N_1270);
nor U2094 (N_2094,In_2483,N_1966);
or U2095 (N_2095,N_377,In_1124);
nor U2096 (N_2096,N_1313,N_1823);
and U2097 (N_2097,N_348,N_1995);
xor U2098 (N_2098,N_1366,N_1304);
and U2099 (N_2099,N_170,N_1229);
or U2100 (N_2100,N_1255,N_1669);
xnor U2101 (N_2101,N_1180,N_1586);
and U2102 (N_2102,N_583,N_1054);
or U2103 (N_2103,In_766,N_1965);
and U2104 (N_2104,In_2551,N_1634);
and U2105 (N_2105,N_1327,N_916);
xor U2106 (N_2106,N_1011,N_1543);
nand U2107 (N_2107,In_4299,N_74);
xnor U2108 (N_2108,N_462,In_2994);
nor U2109 (N_2109,N_740,N_1950);
or U2110 (N_2110,In_4778,N_1155);
and U2111 (N_2111,N_1430,N_1874);
xor U2112 (N_2112,N_1734,N_1970);
and U2113 (N_2113,N_1909,N_929);
nor U2114 (N_2114,N_738,N_809);
or U2115 (N_2115,In_1012,N_1680);
nand U2116 (N_2116,N_902,N_1724);
xor U2117 (N_2117,N_934,N_584);
nor U2118 (N_2118,N_1298,In_2778);
xnor U2119 (N_2119,In_2774,In_1211);
or U2120 (N_2120,N_124,N_1733);
and U2121 (N_2121,N_682,N_1329);
nor U2122 (N_2122,N_1781,N_1563);
or U2123 (N_2123,N_491,In_3190);
and U2124 (N_2124,N_1750,N_1006);
or U2125 (N_2125,In_3848,N_255);
and U2126 (N_2126,N_619,N_1773);
nor U2127 (N_2127,N_333,N_1685);
xor U2128 (N_2128,In_3273,N_527);
and U2129 (N_2129,N_1076,N_1280);
nor U2130 (N_2130,In_1418,N_1358);
xnor U2131 (N_2131,N_48,N_1375);
nand U2132 (N_2132,In_1238,N_661);
or U2133 (N_2133,N_1394,In_4045);
or U2134 (N_2134,N_79,N_32);
and U2135 (N_2135,N_742,N_252);
nor U2136 (N_2136,N_1993,N_962);
or U2137 (N_2137,N_1879,N_590);
nor U2138 (N_2138,In_717,In_3677);
nor U2139 (N_2139,In_4020,N_1900);
nor U2140 (N_2140,In_1654,N_1377);
xnor U2141 (N_2141,In_2664,N_132);
nor U2142 (N_2142,N_1964,N_1696);
nor U2143 (N_2143,In_4703,In_3017);
nor U2144 (N_2144,N_1949,N_1591);
and U2145 (N_2145,N_630,N_1776);
nand U2146 (N_2146,N_1899,N_1850);
and U2147 (N_2147,N_1580,In_452);
nor U2148 (N_2148,N_1129,N_520);
xor U2149 (N_2149,In_2377,N_1687);
nor U2150 (N_2150,In_515,N_1122);
xor U2151 (N_2151,N_1271,N_1617);
nand U2152 (N_2152,N_1633,N_224);
nor U2153 (N_2153,In_614,In_1922);
nand U2154 (N_2154,N_1887,N_1530);
and U2155 (N_2155,N_632,N_479);
and U2156 (N_2156,In_2601,N_1231);
nand U2157 (N_2157,N_678,N_1097);
and U2158 (N_2158,N_401,N_978);
and U2159 (N_2159,N_193,N_723);
or U2160 (N_2160,N_503,N_843);
or U2161 (N_2161,In_3793,N_830);
or U2162 (N_2162,In_1421,N_1843);
and U2163 (N_2163,N_273,N_1113);
and U2164 (N_2164,N_355,In_445);
xor U2165 (N_2165,N_50,In_116);
xnor U2166 (N_2166,In_4567,N_1919);
nor U2167 (N_2167,N_1483,N_49);
or U2168 (N_2168,N_1921,N_1876);
and U2169 (N_2169,N_277,In_1714);
xor U2170 (N_2170,N_155,N_539);
nor U2171 (N_2171,N_304,N_1291);
xor U2172 (N_2172,In_2230,N_1817);
and U2173 (N_2173,In_1323,N_1796);
xnor U2174 (N_2174,N_515,N_428);
xnor U2175 (N_2175,N_423,In_1849);
nand U2176 (N_2176,In_4712,In_827);
and U2177 (N_2177,In_566,N_832);
nand U2178 (N_2178,N_1584,N_176);
nand U2179 (N_2179,In_77,N_1880);
or U2180 (N_2180,N_1665,In_2593);
and U2181 (N_2181,N_1183,N_1666);
or U2182 (N_2182,N_417,N_541);
or U2183 (N_2183,N_1515,In_982);
and U2184 (N_2184,N_478,N_1756);
and U2185 (N_2185,N_703,N_629);
or U2186 (N_2186,N_612,In_3110);
or U2187 (N_2187,N_142,N_1856);
nor U2188 (N_2188,N_1249,N_1890);
nor U2189 (N_2189,In_2395,N_1267);
nand U2190 (N_2190,N_1567,N_33);
or U2191 (N_2191,N_1007,N_747);
nand U2192 (N_2192,N_1372,N_1907);
nor U2193 (N_2193,In_4596,N_1763);
nor U2194 (N_2194,N_1383,N_1095);
nor U2195 (N_2195,N_447,N_1288);
and U2196 (N_2196,N_1243,N_162);
or U2197 (N_2197,N_778,In_134);
nor U2198 (N_2198,N_725,N_870);
and U2199 (N_2199,N_1102,N_1294);
nor U2200 (N_2200,N_1925,N_1704);
nand U2201 (N_2201,N_376,N_1323);
nand U2202 (N_2202,N_392,In_121);
xor U2203 (N_2203,In_727,N_926);
and U2204 (N_2204,N_1112,N_149);
and U2205 (N_2205,N_1769,N_1926);
nor U2206 (N_2206,N_1833,In_2917);
or U2207 (N_2207,In_2210,In_1916);
and U2208 (N_2208,N_63,N_1862);
nor U2209 (N_2209,N_1962,N_1699);
nor U2210 (N_2210,N_761,N_1603);
xor U2211 (N_2211,N_1725,N_1752);
nor U2212 (N_2212,N_261,In_3792);
or U2213 (N_2213,N_1710,In_2702);
xor U2214 (N_2214,N_1740,In_294);
xnor U2215 (N_2215,N_1816,In_4801);
or U2216 (N_2216,N_1761,In_1985);
and U2217 (N_2217,In_2216,N_785);
or U2218 (N_2218,N_1565,N_1159);
nor U2219 (N_2219,In_1412,N_687);
nand U2220 (N_2220,N_1930,N_1225);
and U2221 (N_2221,N_156,In_12);
xnor U2222 (N_2222,N_945,N_101);
or U2223 (N_2223,N_1967,In_640);
xor U2224 (N_2224,N_1151,N_21);
nand U2225 (N_2225,In_1514,In_3253);
xnor U2226 (N_2226,In_1314,N_1509);
xor U2227 (N_2227,In_633,N_572);
xor U2228 (N_2228,In_336,N_1082);
and U2229 (N_2229,N_1251,N_1943);
or U2230 (N_2230,N_1958,In_2131);
or U2231 (N_2231,N_405,N_1008);
and U2232 (N_2232,N_1422,In_2289);
and U2233 (N_2233,N_896,N_954);
nand U2234 (N_2234,N_879,N_1398);
nand U2235 (N_2235,In_2290,N_1600);
xnor U2236 (N_2236,N_1148,N_1130);
or U2237 (N_2237,N_706,N_684);
nor U2238 (N_2238,N_1544,In_3485);
and U2239 (N_2239,In_4431,N_719);
xnor U2240 (N_2240,In_568,In_487);
xor U2241 (N_2241,In_3249,N_1857);
nor U2242 (N_2242,N_284,N_839);
and U2243 (N_2243,In_3294,N_560);
xnor U2244 (N_2244,In_1109,N_1069);
and U2245 (N_2245,N_1178,In_579);
nor U2246 (N_2246,In_1980,In_590);
or U2247 (N_2247,In_4886,N_568);
nor U2248 (N_2248,In_2746,N_1005);
nand U2249 (N_2249,In_3278,In_2015);
nor U2250 (N_2250,In_4859,N_108);
nand U2251 (N_2251,In_3708,N_1822);
or U2252 (N_2252,In_3426,N_1453);
and U2253 (N_2253,In_3516,N_189);
or U2254 (N_2254,N_1019,In_2006);
and U2255 (N_2255,In_4744,In_3299);
nor U2256 (N_2256,N_1078,N_1297);
or U2257 (N_2257,In_299,N_727);
nand U2258 (N_2258,N_1655,N_915);
or U2259 (N_2259,N_577,N_1149);
xor U2260 (N_2260,In_1440,N_947);
nor U2261 (N_2261,N_1293,In_2475);
nand U2262 (N_2262,N_459,In_111);
and U2263 (N_2263,In_2348,In_4670);
and U2264 (N_2264,In_3396,In_1937);
nor U2265 (N_2265,In_3604,N_1188);
and U2266 (N_2266,N_1847,In_2846);
nand U2267 (N_2267,N_800,In_2763);
nand U2268 (N_2268,N_758,N_168);
xor U2269 (N_2269,In_7,In_3134);
nor U2270 (N_2270,In_4649,In_2275);
and U2271 (N_2271,In_466,N_350);
nand U2272 (N_2272,In_4835,N_524);
and U2273 (N_2273,N_427,N_1639);
or U2274 (N_2274,N_744,N_1877);
nand U2275 (N_2275,In_4982,In_2881);
nand U2276 (N_2276,N_467,In_297);
nand U2277 (N_2277,N_1244,In_4203);
nand U2278 (N_2278,N_1640,N_1333);
nor U2279 (N_2279,N_325,In_3349);
xor U2280 (N_2280,N_886,N_433);
nor U2281 (N_2281,N_274,N_1658);
or U2282 (N_2282,N_299,N_1546);
nand U2283 (N_2283,N_1489,N_429);
or U2284 (N_2284,N_833,In_2978);
or U2285 (N_2285,N_1307,In_4976);
nand U2286 (N_2286,In_815,N_1539);
and U2287 (N_2287,N_1593,In_3277);
nand U2288 (N_2288,In_2203,N_1164);
or U2289 (N_2289,N_1806,In_682);
or U2290 (N_2290,In_943,N_1074);
xor U2291 (N_2291,N_592,N_1357);
and U2292 (N_2292,N_122,In_1448);
and U2293 (N_2293,N_59,N_949);
or U2294 (N_2294,N_77,N_498);
xnor U2295 (N_2295,In_2819,N_1741);
xor U2296 (N_2296,N_1232,N_1668);
or U2297 (N_2297,In_4734,N_455);
and U2298 (N_2298,N_1537,N_1269);
xnor U2299 (N_2299,In_4720,N_94);
or U2300 (N_2300,N_290,In_361);
xor U2301 (N_2301,N_930,N_1747);
nand U2302 (N_2302,In_3206,N_1711);
or U2303 (N_2303,N_229,N_1023);
nand U2304 (N_2304,In_4284,N_1867);
nor U2305 (N_2305,In_1334,N_212);
and U2306 (N_2306,In_3159,In_3023);
or U2307 (N_2307,N_766,N_784);
nor U2308 (N_2308,In_289,In_2648);
and U2309 (N_2309,In_4970,N_662);
xnor U2310 (N_2310,In_3238,N_1237);
nor U2311 (N_2311,N_731,N_1185);
and U2312 (N_2312,N_1980,N_1342);
or U2313 (N_2313,N_1691,N_559);
nand U2314 (N_2314,In_2362,N_58);
or U2315 (N_2315,In_4875,N_1904);
nor U2316 (N_2316,N_618,N_119);
or U2317 (N_2317,N_1983,N_548);
and U2318 (N_2318,In_25,In_1369);
and U2319 (N_2319,N_863,N_1173);
or U2320 (N_2320,N_549,N_1642);
or U2321 (N_2321,In_175,N_204);
nand U2322 (N_2322,N_1864,N_354);
or U2323 (N_2323,N_764,In_1405);
xor U2324 (N_2324,N_1230,In_1794);
nor U2325 (N_2325,N_480,N_1363);
xnor U2326 (N_2326,In_2953,N_1999);
nand U2327 (N_2327,N_891,N_52);
or U2328 (N_2328,In_4270,In_3692);
and U2329 (N_2329,N_861,N_1395);
xor U2330 (N_2330,In_3988,In_2857);
xor U2331 (N_2331,N_946,N_1310);
xnor U2332 (N_2332,In_1858,N_314);
and U2333 (N_2333,N_1093,N_932);
nor U2334 (N_2334,N_1621,In_3637);
and U2335 (N_2335,In_2646,N_1605);
nand U2336 (N_2336,In_1840,In_1398);
nor U2337 (N_2337,N_1985,N_1338);
nand U2338 (N_2338,N_1924,In_1964);
nand U2339 (N_2339,N_1292,N_1472);
nor U2340 (N_2340,In_2467,N_636);
nor U2341 (N_2341,N_413,In_1498);
nor U2342 (N_2342,In_2877,N_486);
xnor U2343 (N_2343,In_1574,In_4165);
or U2344 (N_2344,N_241,N_173);
xnor U2345 (N_2345,N_1171,In_1302);
xnor U2346 (N_2346,In_4798,N_363);
and U2347 (N_2347,N_685,In_886);
nand U2348 (N_2348,N_537,N_769);
or U2349 (N_2349,N_1091,N_871);
nor U2350 (N_2350,N_1718,N_1872);
or U2351 (N_2351,In_3241,N_1998);
and U2352 (N_2352,In_3348,In_2343);
and U2353 (N_2353,N_1670,In_1606);
nor U2354 (N_2354,N_1681,In_2339);
nand U2355 (N_2355,N_1513,In_2570);
or U2356 (N_2356,N_754,In_2239);
nor U2357 (N_2357,N_1779,In_4724);
and U2358 (N_2358,N_205,N_674);
nor U2359 (N_2359,N_1485,N_1100);
nor U2360 (N_2360,N_1503,N_175);
nor U2361 (N_2361,N_1364,N_23);
and U2362 (N_2362,N_1218,N_689);
or U2363 (N_2363,N_963,In_4615);
xor U2364 (N_2364,N_1896,In_2178);
xor U2365 (N_2365,N_1072,In_3851);
nand U2366 (N_2366,N_1719,In_2048);
or U2367 (N_2367,N_1883,N_966);
xor U2368 (N_2368,In_3400,N_1657);
and U2369 (N_2369,In_182,In_597);
or U2370 (N_2370,N_794,N_185);
nand U2371 (N_2371,N_803,N_1098);
xor U2372 (N_2372,N_1099,In_702);
nand U2373 (N_2373,In_3478,N_1316);
xor U2374 (N_2374,N_1334,N_1829);
or U2375 (N_2375,N_1858,In_2515);
xnor U2376 (N_2376,In_2324,N_1976);
nand U2377 (N_2377,In_3822,N_317);
nor U2378 (N_2378,N_1814,N_257);
nand U2379 (N_2379,N_1505,In_4493);
or U2380 (N_2380,N_436,In_2840);
xor U2381 (N_2381,N_650,N_1068);
or U2382 (N_2382,In_1313,In_2378);
and U2383 (N_2383,N_1568,N_1121);
nor U2384 (N_2384,N_1947,In_2078);
nand U2385 (N_2385,N_1077,In_3704);
nand U2386 (N_2386,N_291,N_8);
nor U2387 (N_2387,N_1257,N_375);
nor U2388 (N_2388,N_1259,N_1545);
or U2389 (N_2389,In_3949,In_2222);
nand U2390 (N_2390,In_905,N_202);
and U2391 (N_2391,N_226,N_1859);
nand U2392 (N_2392,N_1941,In_4906);
xnor U2393 (N_2393,N_40,N_1189);
and U2394 (N_2394,N_182,In_1503);
xnor U2395 (N_2395,In_4197,N_1504);
nor U2396 (N_2396,In_4354,N_659);
xor U2397 (N_2397,In_615,N_1972);
xnor U2398 (N_2398,N_704,N_159);
nor U2399 (N_2399,In_1319,In_1773);
xnor U2400 (N_2400,N_1573,N_1735);
nand U2401 (N_2401,In_3025,N_316);
xor U2402 (N_2402,In_1318,N_1433);
or U2403 (N_2403,N_1224,N_1163);
or U2404 (N_2404,N_1136,In_2317);
nor U2405 (N_2405,N_1233,N_1646);
nand U2406 (N_2406,N_1117,In_2473);
nand U2407 (N_2407,In_4501,In_1511);
nor U2408 (N_2408,N_1682,N_597);
or U2409 (N_2409,N_172,In_3029);
nand U2410 (N_2410,In_4530,In_4016);
and U2411 (N_2411,In_3923,N_1519);
or U2412 (N_2412,In_1007,N_1362);
nor U2413 (N_2413,N_91,N_20);
nor U2414 (N_2414,N_1798,N_195);
nand U2415 (N_2415,N_1533,In_2883);
and U2416 (N_2416,In_2454,N_746);
xnor U2417 (N_2417,N_1170,N_753);
nand U2418 (N_2418,N_1266,In_4163);
or U2419 (N_2419,N_968,In_559);
nand U2420 (N_2420,N_1870,N_1262);
nand U2421 (N_2421,In_2013,N_1577);
nand U2422 (N_2422,In_2864,In_277);
and U2423 (N_2423,N_174,In_352);
nand U2424 (N_2424,In_2418,In_2613);
or U2425 (N_2425,N_551,N_1106);
xor U2426 (N_2426,N_233,N_610);
nand U2427 (N_2427,In_127,N_495);
nor U2428 (N_2428,In_3976,N_795);
xnor U2429 (N_2429,N_1534,N_716);
or U2430 (N_2430,N_797,N_944);
or U2431 (N_2431,N_626,N_473);
nor U2432 (N_2432,N_1981,In_4309);
or U2433 (N_2433,In_123,N_1553);
or U2434 (N_2434,N_54,In_4085);
nand U2435 (N_2435,N_502,N_1933);
and U2436 (N_2436,In_3379,In_1728);
or U2437 (N_2437,N_1536,N_1540);
or U2438 (N_2438,N_788,N_341);
and U2439 (N_2439,N_1067,N_1278);
nand U2440 (N_2440,N_276,N_1055);
nand U2441 (N_2441,N_819,N_1683);
xor U2442 (N_2442,N_820,N_542);
xor U2443 (N_2443,In_4559,N_281);
or U2444 (N_2444,N_1335,In_2265);
nand U2445 (N_2445,N_209,In_1702);
nor U2446 (N_2446,In_4385,In_1804);
and U2447 (N_2447,In_4018,In_3868);
xor U2448 (N_2448,N_878,In_1620);
xor U2449 (N_2449,N_1835,N_900);
or U2450 (N_2450,In_3034,N_1252);
or U2451 (N_2451,N_362,In_2413);
xor U2452 (N_2452,In_1242,N_1955);
xor U2453 (N_2453,N_1982,N_1480);
xnor U2454 (N_2454,N_601,In_2718);
and U2455 (N_2455,N_1205,N_1671);
or U2456 (N_2456,N_1703,In_3714);
and U2457 (N_2457,N_849,In_2663);
nor U2458 (N_2458,N_1279,N_30);
nor U2459 (N_2459,N_1410,N_1015);
or U2460 (N_2460,In_3045,N_1187);
nand U2461 (N_2461,N_239,N_1825);
and U2462 (N_2462,N_1065,N_472);
or U2463 (N_2463,N_1245,N_1037);
or U2464 (N_2464,N_234,N_288);
or U2465 (N_2465,N_1450,In_2851);
or U2466 (N_2466,N_713,N_776);
xnor U2467 (N_2467,In_3605,N_357);
and U2468 (N_2468,N_695,In_1068);
nor U2469 (N_2469,In_3359,N_1869);
or U2470 (N_2470,In_2049,N_118);
and U2471 (N_2471,N_129,In_1960);
and U2472 (N_2472,N_231,N_1346);
and U2473 (N_2473,N_465,N_1882);
nand U2474 (N_2474,N_407,N_396);
nor U2475 (N_2475,N_1378,N_326);
and U2476 (N_2476,N_922,N_1200);
and U2477 (N_2477,N_976,N_1029);
and U2478 (N_2478,N_658,In_4432);
xnor U2479 (N_2479,N_2,N_1875);
and U2480 (N_2480,N_286,N_827);
nor U2481 (N_2481,N_837,N_338);
xnor U2482 (N_2482,N_64,N_1664);
and U2483 (N_2483,N_1135,In_2234);
or U2484 (N_2484,N_1802,In_4733);
nand U2485 (N_2485,N_975,N_821);
xor U2486 (N_2486,N_1285,N_1885);
and U2487 (N_2487,In_574,N_144);
nand U2488 (N_2488,N_1963,N_1581);
nor U2489 (N_2489,N_1114,N_793);
and U2490 (N_2490,N_14,N_1382);
or U2491 (N_2491,N_529,In_3005);
or U2492 (N_2492,In_4623,N_1246);
and U2493 (N_2493,N_576,In_2496);
or U2494 (N_2494,N_920,N_779);
or U2495 (N_2495,N_1631,N_1039);
nand U2496 (N_2496,N_1242,In_4214);
nor U2497 (N_2497,N_292,N_1490);
nor U2498 (N_2498,N_344,In_2875);
and U2499 (N_2499,N_1629,N_607);
and U2500 (N_2500,N_646,In_4426);
xor U2501 (N_2501,N_349,In_3592);
or U2502 (N_2502,In_58,In_4218);
xnor U2503 (N_2503,In_396,N_446);
nor U2504 (N_2504,In_3539,In_3419);
and U2505 (N_2505,N_578,N_665);
or U2506 (N_2506,N_1700,N_1423);
nand U2507 (N_2507,N_1922,In_3344);
xor U2508 (N_2508,In_2764,N_501);
nand U2509 (N_2509,N_734,In_4476);
xnor U2510 (N_2510,N_757,N_1208);
nor U2511 (N_2511,N_1034,In_634);
and U2512 (N_2512,N_1314,N_1004);
nand U2513 (N_2513,In_355,N_599);
xor U2514 (N_2514,N_466,In_39);
and U2515 (N_2515,N_1009,In_4230);
nand U2516 (N_2516,In_4598,N_1212);
nor U2517 (N_2517,N_1321,N_271);
and U2518 (N_2518,N_631,N_1012);
and U2519 (N_2519,N_1348,N_622);
or U2520 (N_2520,In_2437,N_1511);
xnor U2521 (N_2521,N_1649,N_648);
or U2522 (N_2522,In_4027,N_557);
xnor U2523 (N_2523,In_2487,N_550);
and U2524 (N_2524,N_1309,N_1698);
and U2525 (N_2525,N_1166,In_4981);
nor U2526 (N_2526,N_1799,In_3468);
nor U2527 (N_2527,In_4022,N_815);
nor U2528 (N_2528,In_1653,In_4371);
nor U2529 (N_2529,N_1273,In_4357);
xnor U2530 (N_2530,N_1541,In_4002);
nand U2531 (N_2531,In_2621,N_904);
or U2532 (N_2532,In_1324,N_379);
nor U2533 (N_2533,N_408,N_1559);
and U2534 (N_2534,N_567,N_845);
nor U2535 (N_2535,In_2915,N_1547);
nand U2536 (N_2536,N_1240,In_4489);
and U2537 (N_2537,N_1345,N_1311);
nand U2538 (N_2538,N_1042,N_287);
or U2539 (N_2539,In_2720,N_1254);
xnor U2540 (N_2540,In_464,In_2768);
xor U2541 (N_2541,In_881,N_591);
nor U2542 (N_2542,In_35,In_4872);
nand U2543 (N_2543,In_4468,N_594);
xor U2544 (N_2544,N_681,In_4073);
nor U2545 (N_2545,In_4239,N_1892);
or U2546 (N_2546,N_675,N_1791);
or U2547 (N_2547,In_4106,In_1939);
xnor U2548 (N_2548,N_1143,N_1051);
nand U2549 (N_2549,N_887,N_1895);
xor U2550 (N_2550,In_2408,N_836);
and U2551 (N_2551,In_3858,In_2173);
nor U2552 (N_2552,In_3509,In_3229);
or U2553 (N_2553,In_1696,In_1239);
or U2554 (N_2554,N_707,N_308);
nand U2555 (N_2555,In_4554,N_120);
nand U2556 (N_2556,N_959,N_1578);
and U2557 (N_2557,N_285,N_700);
xor U2558 (N_2558,N_200,In_4730);
and U2559 (N_2559,N_1145,N_1975);
or U2560 (N_2560,N_228,In_2219);
xnor U2561 (N_2561,In_2791,N_1848);
nand U2562 (N_2562,N_1625,N_13);
nor U2563 (N_2563,N_1268,N_42);
or U2564 (N_2564,N_1318,N_712);
nor U2565 (N_2565,N_910,N_197);
nand U2566 (N_2566,N_1610,N_360);
nand U2567 (N_2567,In_1749,In_4766);
xnor U2568 (N_2568,N_1777,N_500);
or U2569 (N_2569,In_36,In_2573);
xnor U2570 (N_2570,N_295,In_2743);
and U2571 (N_2571,In_4672,N_18);
xnor U2572 (N_2572,N_508,N_799);
and U2573 (N_2573,N_880,N_582);
or U2574 (N_2574,N_634,In_1103);
nand U2575 (N_2575,N_801,N_270);
xnor U2576 (N_2576,N_1425,In_3372);
and U2577 (N_2577,In_3157,N_1223);
xor U2578 (N_2578,In_1123,N_1554);
nand U2579 (N_2579,N_1499,N_322);
and U2580 (N_2580,In_377,N_1551);
nand U2581 (N_2581,N_106,In_3787);
xor U2582 (N_2582,N_1937,N_1745);
or U2583 (N_2583,N_494,In_3500);
or U2584 (N_2584,In_2253,In_1898);
nand U2585 (N_2585,N_1386,In_1743);
xor U2586 (N_2586,N_1815,N_1454);
and U2587 (N_2587,N_1897,N_855);
or U2588 (N_2588,N_536,N_1732);
and U2589 (N_2589,In_356,N_7);
or U2590 (N_2590,N_1,N_238);
or U2591 (N_2591,In_4938,N_490);
xnor U2592 (N_2592,N_1971,N_1021);
xnor U2593 (N_2593,N_1370,N_474);
xnor U2594 (N_2594,N_789,In_4955);
and U2595 (N_2595,N_44,N_1641);
and U2596 (N_2596,N_1127,In_2719);
nand U2597 (N_2597,In_617,In_2081);
or U2598 (N_2598,N_1566,N_1184);
or U2599 (N_2599,N_1263,N_469);
nand U2600 (N_2600,N_6,N_511);
or U2601 (N_2601,In_2032,In_1739);
or U2602 (N_2602,In_4761,N_564);
nor U2603 (N_2603,N_303,In_3120);
nand U2604 (N_2604,N_102,N_1512);
nand U2605 (N_2605,N_227,N_1821);
xor U2606 (N_2606,In_1297,N_1371);
and U2607 (N_2607,In_1176,N_722);
or U2608 (N_2608,N_1622,In_1388);
nor U2609 (N_2609,In_4586,N_382);
xor U2610 (N_2610,In_2363,N_531);
or U2611 (N_2611,N_905,In_253);
and U2612 (N_2612,N_615,N_1493);
nor U2613 (N_2613,In_1460,N_448);
nand U2614 (N_2614,N_25,In_2826);
or U2615 (N_2615,N_1306,N_1020);
or U2616 (N_2616,N_361,In_1301);
and U2617 (N_2617,In_4289,N_306);
and U2618 (N_2618,N_1968,In_5);
or U2619 (N_2619,N_368,N_1818);
or U2620 (N_2620,In_3460,In_1497);
nand U2621 (N_2621,N_269,N_272);
and U2622 (N_2622,N_398,In_4691);
xor U2623 (N_2623,In_685,In_2197);
or U2624 (N_2624,N_372,N_437);
nand U2625 (N_2625,N_1912,N_941);
and U2626 (N_2626,In_3905,N_1281);
and U2627 (N_2627,N_1574,N_1861);
nand U2628 (N_2628,N_822,N_380);
or U2629 (N_2629,N_782,In_3865);
xor U2630 (N_2630,In_4994,N_1083);
nand U2631 (N_2631,N_1144,N_1918);
and U2632 (N_2632,N_996,N_600);
or U2633 (N_2633,N_575,N_111);
nand U2634 (N_2634,N_1753,N_518);
nand U2635 (N_2635,N_1828,In_1414);
and U2636 (N_2636,In_56,N_677);
nand U2637 (N_2637,N_1596,In_811);
and U2638 (N_2638,In_3239,N_935);
nand U2639 (N_2639,N_1676,In_1322);
xor U2640 (N_2640,N_82,N_1092);
or U2641 (N_2641,N_418,N_653);
and U2642 (N_2642,In_1420,N_1914);
xnor U2643 (N_2643,N_0,In_1850);
or U2644 (N_2644,In_3573,N_481);
nor U2645 (N_2645,N_1456,N_1351);
or U2646 (N_2646,N_1615,N_705);
nand U2647 (N_2647,N_1831,N_1488);
xnor U2648 (N_2648,In_4004,In_4395);
xnor U2649 (N_2649,In_4160,In_4306);
nor U2650 (N_2650,In_4294,N_532);
or U2651 (N_2651,N_1716,N_1558);
nor U2652 (N_2652,In_2211,In_4409);
xor U2653 (N_2653,N_1186,N_571);
xnor U2654 (N_2654,N_1635,N_835);
xor U2655 (N_2655,In_4751,In_4423);
nand U2656 (N_2656,N_136,In_454);
or U2657 (N_2657,N_1873,N_1414);
nor U2658 (N_2658,N_321,N_824);
nor U2659 (N_2659,In_801,N_1328);
and U2660 (N_2660,N_513,In_27);
xor U2661 (N_2661,N_933,N_275);
nand U2662 (N_2662,N_783,N_604);
nor U2663 (N_2663,N_412,N_365);
nor U2664 (N_2664,In_3117,In_3656);
xnor U2665 (N_2665,In_810,N_461);
xor U2666 (N_2666,In_3096,In_2185);
and U2667 (N_2667,N_540,N_371);
and U2668 (N_2668,N_633,In_1228);
nand U2669 (N_2669,N_80,N_1402);
nand U2670 (N_2670,N_1134,In_572);
or U2671 (N_2671,In_4634,N_1352);
nor U2672 (N_2672,N_1973,In_2565);
and U2673 (N_2673,In_4136,N_1632);
or U2674 (N_2674,N_1013,N_928);
nand U2675 (N_2675,N_115,N_851);
and U2676 (N_2676,In_1566,N_107);
nor U2677 (N_2677,N_1905,N_846);
xnor U2678 (N_2678,N_856,In_1784);
or U2679 (N_2679,N_165,N_1415);
and U2680 (N_2680,N_517,N_1778);
or U2681 (N_2681,In_3726,N_997);
nand U2682 (N_2682,In_4888,N_127);
and U2683 (N_2683,N_923,In_2451);
nand U2684 (N_2684,In_250,N_1468);
and U2685 (N_2685,N_1626,N_1614);
and U2686 (N_2686,In_3230,In_152);
nor U2687 (N_2687,N_251,N_1057);
xor U2688 (N_2688,In_2372,In_849);
or U2689 (N_2689,N_244,In_3155);
and U2690 (N_2690,In_1927,In_4496);
nand U2691 (N_2691,N_1583,In_4086);
and U2692 (N_2692,In_651,N_1343);
nand U2693 (N_2693,In_3862,In_494);
nand U2694 (N_2694,N_1893,In_1249);
xor U2695 (N_2695,N_1886,N_279);
nor U2696 (N_2696,N_985,In_4637);
or U2697 (N_2697,N_236,In_3987);
xor U2698 (N_2698,N_1216,N_435);
nand U2699 (N_2699,N_430,N_89);
nor U2700 (N_2700,In_4572,In_3562);
and U2701 (N_2701,In_1733,In_3702);
xor U2702 (N_2702,N_1062,N_1662);
and U2703 (N_2703,N_1458,N_1595);
xor U2704 (N_2704,N_1409,N_1768);
and U2705 (N_2705,In_1080,N_253);
or U2706 (N_2706,N_1789,N_1411);
and U2707 (N_2707,N_1994,N_649);
or U2708 (N_2708,N_528,In_1041);
xnor U2709 (N_2709,N_1406,N_1760);
nor U2710 (N_2710,N_1385,N_1510);
nand U2711 (N_2711,N_1588,N_1830);
nor U2712 (N_2712,In_3077,N_1264);
and U2713 (N_2713,N_386,N_109);
xnor U2714 (N_2714,In_2293,N_449);
and U2715 (N_2715,N_1528,In_3384);
and U2716 (N_2716,N_624,N_1368);
or U2717 (N_2717,N_724,In_343);
or U2718 (N_2718,N_909,In_1888);
and U2719 (N_2719,N_1656,N_921);
nand U2720 (N_2720,N_1754,N_1868);
and U2721 (N_2721,In_1838,N_1108);
and U2722 (N_2722,N_611,N_977);
or U2723 (N_2723,N_150,In_1480);
or U2724 (N_2724,N_1174,N_1031);
and U2725 (N_2725,In_2182,In_29);
nand U2726 (N_2726,N_390,N_1672);
nor U2727 (N_2727,N_912,In_1757);
or U2728 (N_2728,In_13,In_2754);
or U2729 (N_2729,N_936,In_3448);
and U2730 (N_2730,N_538,N_1936);
and U2731 (N_2731,In_0,N_1491);
xnor U2732 (N_2732,N_1032,In_3730);
nor U2733 (N_2733,N_745,N_1535);
and U2734 (N_2734,N_621,N_399);
nand U2735 (N_2735,N_26,N_225);
or U2736 (N_2736,In_582,N_424);
nor U2737 (N_2737,N_826,In_170);
or U2738 (N_2738,N_639,N_1944);
nand U2739 (N_2739,In_436,N_78);
or U2740 (N_2740,In_2104,N_29);
xnor U2741 (N_2741,N_1461,In_2932);
nand U2742 (N_2742,N_672,N_15);
or U2743 (N_2743,In_4522,N_1451);
nor U2744 (N_2744,In_2549,In_2350);
nand U2745 (N_2745,N_1628,N_817);
and U2746 (N_2746,N_11,In_1092);
and U2747 (N_2747,N_1624,In_3183);
nor U2748 (N_2748,N_340,N_580);
and U2749 (N_2749,N_240,N_1772);
and U2750 (N_2750,N_1884,N_1359);
nand U2751 (N_2751,N_888,N_1770);
and U2752 (N_2752,N_72,N_1428);
or U2753 (N_2753,In_1826,N_998);
nor U2754 (N_2754,N_302,N_1277);
and U2755 (N_2755,In_2535,N_47);
nor U2756 (N_2756,N_143,In_3620);
xor U2757 (N_2757,In_759,In_1100);
or U2758 (N_2758,N_1623,N_603);
or U2759 (N_2759,N_750,N_777);
nand U2760 (N_2760,In_1008,N_1903);
nor U2761 (N_2761,N_90,N_452);
nand U2762 (N_2762,In_3602,N_914);
and U2763 (N_2763,N_419,N_516);
nor U2764 (N_2764,N_1988,N_337);
xor U2765 (N_2765,N_1604,In_924);
and U2766 (N_2766,N_489,N_534);
nor U2767 (N_2767,In_2352,N_1033);
and U2768 (N_2768,In_3606,N_1439);
and U2769 (N_2769,In_3715,N_439);
xor U2770 (N_2770,N_1959,In_3529);
or U2771 (N_2771,N_543,N_1190);
and U2772 (N_2772,N_1241,N_388);
xor U2773 (N_2773,N_1838,N_201);
or U2774 (N_2774,N_1840,N_589);
or U2775 (N_2775,In_80,In_2563);
and U2776 (N_2776,N_663,N_460);
or U2777 (N_2777,N_1762,N_1236);
and U2778 (N_2778,In_1387,N_1290);
and U2779 (N_2779,In_403,N_918);
or U2780 (N_2780,N_1373,In_478);
nor U2781 (N_2781,N_951,N_88);
or U2782 (N_2782,In_4600,N_117);
nor U2783 (N_2783,In_4973,N_1317);
nor U2784 (N_2784,In_2406,In_1005);
and U2785 (N_2785,N_206,N_545);
xor U2786 (N_2786,In_2469,In_302);
and U2787 (N_2787,N_890,N_248);
xnor U2788 (N_2788,In_3162,N_1403);
xnor U2789 (N_2789,In_2686,N_1355);
nand U2790 (N_2790,In_4963,In_2307);
nand U2791 (N_2791,N_289,N_640);
nand U2792 (N_2792,N_1038,N_1475);
xor U2793 (N_2793,In_4108,N_420);
nor U2794 (N_2794,In_2038,N_1132);
nand U2795 (N_2795,N_774,In_1148);
nand U2796 (N_2796,N_1284,N_1677);
or U2797 (N_2797,N_75,N_960);
and U2798 (N_2798,N_1590,N_894);
nor U2799 (N_2799,N_553,N_370);
nor U2800 (N_2800,In_1072,N_183);
and U2801 (N_2801,N_1452,In_4474);
and U2802 (N_2802,N_1369,N_1555);
or U2803 (N_2803,N_1661,N_1330);
or U2804 (N_2804,N_1550,In_2155);
or U2805 (N_2805,N_1542,N_364);
and U2806 (N_2806,In_4965,N_892);
nor U2807 (N_2807,N_1514,N_1449);
xor U2808 (N_2808,N_179,In_3269);
nand U2809 (N_2809,N_1939,N_1517);
nand U2810 (N_2810,In_688,In_4772);
and U2811 (N_2811,In_2449,N_1552);
nor U2812 (N_2812,N_1607,N_1191);
or U2813 (N_2813,In_4817,In_1926);
nand U2814 (N_2814,N_1045,In_305);
xor U2815 (N_2815,In_2012,N_1081);
and U2816 (N_2816,N_1018,In_1062);
nor U2817 (N_2817,N_697,N_1444);
and U2818 (N_2818,N_1697,N_1282);
nor U2819 (N_2819,In_1499,N_1347);
nand U2820 (N_2820,N_1800,N_1978);
nor U2821 (N_2821,N_237,In_1644);
nor U2822 (N_2822,N_1714,N_579);
nand U2823 (N_2823,N_266,In_756);
and U2824 (N_2824,N_1495,In_653);
nor U2825 (N_2825,N_1767,N_1050);
or U2826 (N_2826,N_765,In_4549);
nand U2827 (N_2827,N_898,In_4390);
nor U2828 (N_2828,N_1289,N_166);
xnor U2829 (N_2829,N_1408,In_1340);
or U2830 (N_2830,N_1638,N_373);
xnor U2831 (N_2831,N_250,N_1150);
nand U2832 (N_2832,In_4305,N_969);
xor U2833 (N_2833,N_883,N_218);
or U2834 (N_2834,N_1427,N_526);
xnor U2835 (N_2835,N_1179,N_67);
nand U2836 (N_2836,N_729,N_953);
nand U2837 (N_2837,N_721,N_1445);
and U2838 (N_2838,In_3195,N_114);
nor U2839 (N_2839,N_1780,N_307);
and U2840 (N_2840,N_1709,In_3404);
nand U2841 (N_2841,In_2531,In_1458);
xnor U2842 (N_2842,N_1047,In_271);
nand U2843 (N_2843,N_1048,In_1430);
nor U2844 (N_2844,N_808,N_406);
and U2845 (N_2845,N_1805,In_678);
and U2846 (N_2846,In_783,In_2409);
and U2847 (N_2847,N_367,N_1611);
nor U2848 (N_2848,N_563,N_1679);
and U2849 (N_2849,N_46,N_1948);
nor U2850 (N_2850,N_188,In_1576);
xor U2851 (N_2851,N_1265,N_441);
nand U2852 (N_2852,N_1125,N_1466);
or U2853 (N_2853,N_1736,N_153);
or U2854 (N_2854,In_1604,N_1470);
and U2855 (N_2855,N_148,In_3072);
nand U2856 (N_2856,In_4380,In_1877);
nand U2857 (N_2857,N_347,N_1757);
and U2858 (N_2858,N_547,N_925);
nor U2859 (N_2859,N_701,N_772);
and U2860 (N_2860,N_999,N_730);
xor U2861 (N_2861,N_1217,N_1396);
and U2862 (N_2862,In_4866,N_3);
xor U2863 (N_2863,N_558,N_1548);
or U2864 (N_2864,N_190,N_595);
nor U2865 (N_2865,In_3193,In_527);
or U2866 (N_2866,In_3038,In_3480);
and U2867 (N_2867,N_343,N_986);
or U2868 (N_2868,In_306,N_865);
or U2869 (N_2869,In_201,N_1597);
xor U2870 (N_2870,N_813,In_1380);
nor U2871 (N_2871,N_1954,In_2384);
or U2872 (N_2872,N_552,In_282);
nor U2873 (N_2873,N_507,N_1902);
nor U2874 (N_2874,N_958,N_402);
and U2875 (N_2875,N_92,N_964);
nand U2876 (N_2876,N_1300,In_3995);
nand U2877 (N_2877,N_178,In_4901);
and U2878 (N_2878,In_3530,N_1527);
xnor U2879 (N_2879,In_4066,N_1820);
nand U2880 (N_2880,N_605,N_1374);
nor U2881 (N_2881,N_1766,In_52);
nand U2882 (N_2882,N_1286,N_544);
or U2883 (N_2883,In_3557,N_699);
xor U2884 (N_2884,N_1651,In_2100);
and U2885 (N_2885,In_3089,N_1167);
nor U2886 (N_2886,N_810,In_1540);
or U2887 (N_2887,N_163,In_2273);
or U2888 (N_2888,N_456,N_1275);
xor U2889 (N_2889,N_1339,In_1350);
nand U2890 (N_2890,N_22,N_135);
or U2891 (N_2891,N_938,N_1399);
and U2892 (N_2892,In_570,N_842);
and U2893 (N_2893,N_1387,In_3222);
or U2894 (N_2894,N_1654,N_1852);
xnor U2895 (N_2895,N_1837,In_2823);
or U2896 (N_2896,N_1025,N_36);
and U2897 (N_2897,N_1807,N_458);
or U2898 (N_2898,N_161,N_1443);
nor U2899 (N_2899,N_43,N_336);
and U2900 (N_2900,In_3098,N_1219);
and U2901 (N_2901,In_2073,N_421);
nand U2902 (N_2902,In_1465,N_298);
nand U2903 (N_2903,N_1570,N_1228);
nor U2904 (N_2904,N_1846,N_294);
and U2905 (N_2905,N_841,N_1616);
nand U2906 (N_2906,In_3842,N_1643);
or U2907 (N_2907,N_714,N_1424);
xnor U2908 (N_2908,In_159,In_2288);
or U2909 (N_2909,In_1280,N_834);
nor U2910 (N_2910,N_1569,In_4233);
xor U2911 (N_2911,N_1990,N_943);
or U2912 (N_2912,In_3036,In_421);
or U2913 (N_2913,N_164,In_2740);
nor U2914 (N_2914,N_1128,N_1497);
and U2915 (N_2915,N_628,In_4351);
or U2916 (N_2916,N_1927,In_1082);
nand U2917 (N_2917,In_3673,N_762);
nand U2918 (N_2918,N_1226,N_798);
or U2919 (N_2919,In_3405,N_1878);
nor U2920 (N_2920,N_741,N_1942);
or U2921 (N_2921,In_354,N_198);
nor U2922 (N_2922,In_4527,N_1261);
xor U2923 (N_2923,N_751,N_1996);
and U2924 (N_2924,N_99,N_323);
and U2925 (N_2925,N_702,N_773);
nor U2926 (N_2926,N_1133,In_3744);
or U2927 (N_2927,In_2338,In_4317);
and U2928 (N_2928,In_4021,N_1138);
nor U2929 (N_2929,N_739,In_4410);
and U2930 (N_2930,In_2134,In_4851);
and U2931 (N_2931,N_191,N_874);
nor U2932 (N_2932,N_1989,In_3497);
nand U2933 (N_2933,N_1412,N_1248);
nand U2934 (N_2934,N_1759,N_983);
and U2935 (N_2935,In_3759,In_3119);
and U2936 (N_2936,In_3679,N_1440);
nor U2937 (N_2937,N_1391,N_1075);
or U2938 (N_2938,N_708,N_1107);
nand U2939 (N_2939,In_4184,N_391);
or U2940 (N_2940,N_1478,In_1381);
or U2941 (N_2941,N_823,N_1945);
nand U2942 (N_2942,In_3933,N_1758);
and U2943 (N_2943,N_1723,N_1238);
or U2944 (N_2944,N_1819,N_1089);
xor U2945 (N_2945,N_374,N_1526);
xnor U2946 (N_2946,In_1830,N_972);
nand U2947 (N_2947,N_434,In_1619);
nand U2948 (N_2948,N_96,In_4825);
nor U2949 (N_2949,In_427,In_1990);
xnor U2950 (N_2950,N_1589,N_211);
nand U2951 (N_2951,N_980,In_794);
or U2952 (N_2952,N_1405,N_215);
nand U2953 (N_2953,N_1487,N_1742);
nor U2954 (N_2954,N_1350,N_1484);
or U2955 (N_2955,In_2695,N_113);
xor U2956 (N_2956,In_4897,N_57);
nand U2957 (N_2957,In_2309,N_258);
nand U2958 (N_2958,N_280,In_2724);
or U2959 (N_2959,N_818,N_1101);
nand U2960 (N_2960,In_2627,In_3670);
or U2961 (N_2961,N_825,N_1931);
xnor U2962 (N_2962,N_487,N_56);
and U2963 (N_2963,In_3171,N_1156);
and U2964 (N_2964,N_1957,N_278);
xor U2965 (N_2965,N_1717,N_1421);
or U2966 (N_2966,In_880,In_4312);
or U2967 (N_2967,N_245,N_868);
or U2968 (N_2968,N_1898,N_1842);
and U2969 (N_2969,N_1003,In_4256);
or U2970 (N_2970,N_807,In_938);
and U2971 (N_2971,N_493,N_39);
and U2972 (N_2972,N_312,N_987);
nand U2973 (N_2973,In_737,N_1201);
nand U2974 (N_2974,N_167,N_606);
nand U2975 (N_2975,N_1660,N_614);
or U2976 (N_2976,N_1561,N_254);
nand U2977 (N_2977,In_4171,N_1783);
xor U2978 (N_2978,N_911,N_885);
nand U2979 (N_2979,In_2783,N_339);
or U2980 (N_2980,In_3755,N_1376);
xor U2981 (N_2981,In_1256,In_4232);
or U2982 (N_2982,In_3202,N_756);
xnor U2983 (N_2983,N_664,N_1058);
and U2984 (N_2984,In_1876,N_1705);
xnor U2985 (N_2985,In_1539,N_1612);
xnor U2986 (N_2986,In_3410,N_70);
and U2987 (N_2987,N_160,N_1997);
and U2988 (N_2988,N_324,N_1575);
nor U2989 (N_2989,In_1741,In_2215);
nand U2990 (N_2990,In_4391,N_828);
xnor U2991 (N_2991,N_1094,N_617);
or U2992 (N_2992,N_1088,N_510);
nand U2993 (N_2993,In_4762,In_4438);
xnor U2994 (N_2994,N_1426,In_3742);
nand U2995 (N_2995,N_223,N_268);
nand U2996 (N_2996,N_1502,N_1977);
and U2997 (N_2997,N_1784,N_991);
and U2998 (N_2998,N_152,In_505);
or U2999 (N_2999,In_2788,N_1465);
nand U3000 (N_3000,In_1378,N_1002);
nand U3001 (N_3001,In_4673,N_440);
nor U3002 (N_3002,N_876,N_246);
or U3003 (N_3003,In_663,N_881);
nor U3004 (N_3004,In_3378,N_10);
or U3005 (N_3005,In_3345,N_642);
nor U3006 (N_3006,N_1826,N_1115);
and U3007 (N_3007,N_1841,N_1026);
xnor U3008 (N_3008,N_194,N_763);
nor U3009 (N_3009,In_1941,N_1917);
nor U3010 (N_3010,N_1894,N_1692);
and U3011 (N_3011,N_643,N_1301);
nand U3012 (N_3012,N_319,N_1090);
nand U3013 (N_3013,N_83,In_3390);
xor U3014 (N_3014,N_1152,N_967);
or U3015 (N_3015,N_151,N_1274);
nand U3016 (N_3016,In_3463,N_562);
xor U3017 (N_3017,In_4060,N_647);
or U3018 (N_3018,In_4314,N_1221);
and U3019 (N_3019,N_387,In_2603);
and U3020 (N_3020,In_89,In_4182);
xor U3021 (N_3021,N_134,N_1960);
and U3022 (N_3022,N_1721,N_1442);
nand U3023 (N_3023,In_3927,In_203);
nand U3024 (N_3024,N_1839,In_1425);
or U3025 (N_3025,In_2704,N_775);
and U3026 (N_3026,N_1932,N_393);
nor U3027 (N_3027,N_328,N_829);
or U3028 (N_3028,In_2760,In_3099);
xor U3029 (N_3029,In_1752,In_1332);
nor U3030 (N_3030,N_1929,N_971);
xor U3031 (N_3031,N_217,In_1999);
and U3032 (N_3032,N_62,N_792);
or U3033 (N_3033,N_1956,N_812);
xor U3034 (N_3034,N_358,N_635);
nand U3035 (N_3035,N_199,N_668);
xnor U3036 (N_3036,N_445,In_2322);
xor U3037 (N_3037,N_1302,N_496);
nor U3038 (N_3038,In_2993,N_743);
nand U3039 (N_3039,N_1182,In_1624);
nor U3040 (N_3040,In_279,N_609);
nand U3041 (N_3041,N_1739,N_87);
nor U3042 (N_3042,In_4533,N_1774);
nand U3043 (N_3043,In_2507,In_60);
and U3044 (N_3044,N_1836,In_3594);
nand U3045 (N_3045,N_1529,In_1760);
nor U3046 (N_3046,N_596,In_779);
and U3047 (N_3047,N_366,In_2893);
nor U3048 (N_3048,N_69,N_1110);
nand U3049 (N_3049,N_1579,N_952);
nor U3050 (N_3050,In_4773,N_1295);
and U3051 (N_3051,In_3342,In_891);
nand U3052 (N_3052,In_780,In_460);
or U3053 (N_3053,In_3535,In_2938);
nor U3054 (N_3054,In_4082,N_908);
xnor U3055 (N_3055,In_4846,N_104);
xor U3056 (N_3056,N_736,N_1379);
and U3057 (N_3057,N_24,N_1863);
nor U3058 (N_3058,N_1177,N_901);
and U3059 (N_3059,N_282,N_1953);
xnor U3060 (N_3060,In_621,N_1419);
nor U3061 (N_3061,In_4254,In_2485);
nor U3062 (N_3062,N_19,In_1233);
xnor U3063 (N_3063,N_1176,N_1928);
nor U3064 (N_3064,In_1841,N_1694);
xnor U3065 (N_3065,In_287,N_1674);
nor U3066 (N_3066,N_146,In_2759);
or U3067 (N_3067,N_1645,In_523);
nand U3068 (N_3068,In_2987,N_1084);
and U3069 (N_3069,N_395,N_1793);
nor U3070 (N_3070,N_733,In_2848);
nand U3071 (N_3071,N_85,N_1508);
or U3072 (N_3072,N_995,In_4625);
nand U3073 (N_3073,N_1303,N_1952);
and U3074 (N_3074,N_1198,In_4510);
and U3075 (N_3075,In_2789,In_764);
or U3076 (N_3076,N_1063,N_857);
or U3077 (N_3077,N_1436,N_1030);
and U3078 (N_3078,In_1681,N_313);
xor U3079 (N_3079,N_1326,In_730);
nand U3080 (N_3080,N_409,N_1482);
or U3081 (N_3081,N_16,In_878);
nor U3082 (N_3082,N_1690,In_2560);
or U3083 (N_3083,N_243,In_3496);
nand U3084 (N_3084,N_1969,N_444);
or U3085 (N_3085,In_560,N_1222);
nor U3086 (N_3086,In_2079,N_158);
or U3087 (N_3087,In_1682,N_1214);
and U3088 (N_3088,In_2374,N_755);
and U3089 (N_3089,In_133,N_267);
nor U3090 (N_3090,N_352,N_138);
xnor U3091 (N_3091,In_4221,N_696);
and U3092 (N_3092,N_831,N_1181);
and U3093 (N_3093,N_760,N_1813);
nor U3094 (N_3094,N_1071,N_1908);
nor U3095 (N_3095,N_66,In_2884);
and U3096 (N_3096,N_1400,N_1693);
nor U3097 (N_3097,In_474,N_1203);
and U3098 (N_3098,In_2571,In_3694);
nor U3099 (N_3099,N_1227,In_4105);
nand U3100 (N_3100,N_680,In_553);
xor U3101 (N_3101,N_1923,In_785);
nor U3102 (N_3102,In_631,N_400);
or U3103 (N_3103,N_1477,In_1426);
and U3104 (N_3104,N_1283,N_1429);
xnor U3105 (N_3105,In_3055,N_471);
nand U3106 (N_3106,N_787,N_100);
nand U3107 (N_3107,N_463,N_1220);
and U3108 (N_3108,N_981,N_1141);
xnor U3109 (N_3109,N_414,N_990);
nand U3110 (N_3110,In_2373,N_1532);
or U3111 (N_3111,N_882,In_269);
or U3112 (N_3112,N_1587,In_1296);
or U3113 (N_3113,N_1834,In_1483);
nor U3114 (N_3114,In_4155,N_973);
and U3115 (N_3115,N_1432,N_432);
and U3116 (N_3116,In_4324,N_1619);
or U3117 (N_3117,N_1085,N_994);
and U3118 (N_3118,N_1079,N_1332);
nand U3119 (N_3119,In_1219,N_1853);
xor U3120 (N_3120,In_3006,N_1663);
and U3121 (N_3121,N_859,N_1979);
and U3122 (N_3122,In_1970,In_3494);
xnor U3123 (N_3123,N_786,N_126);
nand U3124 (N_3124,N_673,N_1146);
nor U3125 (N_3125,N_1647,N_1322);
and U3126 (N_3126,N_884,N_1247);
nor U3127 (N_3127,N_327,In_1933);
and U3128 (N_3128,N_965,N_1070);
nand U3129 (N_3129,In_1454,N_1299);
and U3130 (N_3130,N_1418,N_1459);
or U3131 (N_3131,N_679,N_588);
nor U3132 (N_3132,N_1471,N_1986);
or U3133 (N_3133,In_286,In_3966);
xor U3134 (N_3134,N_844,In_1647);
and U3135 (N_3135,In_3559,N_625);
xnor U3136 (N_3136,N_318,N_1434);
nor U3137 (N_3137,N_1934,N_717);
xor U3138 (N_3138,In_1577,In_893);
and U3139 (N_3139,N_249,In_3913);
nand U3140 (N_3140,N_301,N_492);
or U3141 (N_3141,N_394,In_1507);
nor U3142 (N_3142,In_2614,N_426);
xnor U3143 (N_3143,N_850,N_1105);
xor U3144 (N_3144,N_1712,N_1022);
xor U3145 (N_3145,N_546,N_623);
xor U3146 (N_3146,N_385,N_112);
or U3147 (N_3147,N_187,In_4723);
xor U3148 (N_3148,N_1729,N_1785);
or U3149 (N_3149,N_1204,N_416);
nand U3150 (N_3150,In_2824,N_644);
nor U3151 (N_3151,In_3601,N_1028);
or U3152 (N_3152,N_1755,N_660);
or U3153 (N_3153,In_4593,In_4292);
xnor U3154 (N_3154,N_1353,N_1492);
or U3155 (N_3155,N_1496,N_505);
and U3156 (N_3156,N_907,In_4547);
nor U3157 (N_3157,In_4531,In_543);
nand U3158 (N_3158,N_1844,In_1217);
nand U3159 (N_3159,N_411,In_1803);
xor U3160 (N_3160,In_2843,N_1522);
or U3161 (N_3161,N_752,N_81);
nand U3162 (N_3162,N_232,In_939);
or U3163 (N_3163,N_262,In_1039);
nand U3164 (N_3164,In_171,N_1786);
and U3165 (N_3165,N_442,N_1961);
nor U3166 (N_3166,N_1764,N_1520);
or U3167 (N_3167,N_864,N_438);
or U3168 (N_3168,N_453,N_1001);
or U3169 (N_3169,In_3609,In_2907);
nand U3170 (N_3170,N_1525,In_4838);
xnor U3171 (N_3171,In_2947,N_710);
nor U3172 (N_3172,N_1250,N_847);
or U3173 (N_3173,N_140,N_425);
nand U3174 (N_3174,N_767,In_2853);
nand U3175 (N_3175,In_2506,N_1667);
xnor U3176 (N_3176,In_4124,N_1889);
xor U3177 (N_3177,N_1594,In_1330);
nor U3178 (N_3178,N_1448,N_858);
and U3179 (N_3179,N_356,In_1291);
xnor U3180 (N_3180,N_638,N_1324);
and U3181 (N_3181,In_930,N_1276);
nand U3182 (N_3182,In_337,In_541);
xor U3183 (N_3183,N_221,N_1116);
nand U3184 (N_3184,In_3722,N_1601);
nor U3185 (N_3185,N_1109,N_65);
xnor U3186 (N_3186,N_1653,N_1731);
or U3187 (N_3187,N_141,In_2587);
nand U3188 (N_3188,N_1154,In_4855);
and U3189 (N_3189,In_314,N_1142);
nand U3190 (N_3190,N_585,In_1230);
or U3191 (N_3191,N_670,In_4948);
xnor U3192 (N_3192,N_728,N_1211);
nor U3193 (N_3193,N_791,In_3429);
nand U3194 (N_3194,N_869,N_1618);
and U3195 (N_3195,N_37,N_899);
xnor U3196 (N_3196,In_3777,In_3841);
and U3197 (N_3197,N_403,In_760);
nand U3198 (N_3198,N_220,In_4176);
or U3199 (N_3199,N_1920,N_514);
nand U3200 (N_3200,In_1844,In_3327);
nand U3201 (N_3201,N_768,N_1035);
or U3202 (N_3202,N_1812,N_875);
nand U3203 (N_3203,N_1689,In_2585);
xnor U3204 (N_3204,N_345,N_31);
or U3205 (N_3205,N_512,N_310);
xnor U3206 (N_3206,In_184,N_1344);
nand U3207 (N_3207,In_1795,N_1804);
nand U3208 (N_3208,In_2196,N_1518);
xor U3209 (N_3209,N_1516,In_3947);
xor U3210 (N_3210,In_3214,In_503);
xnor U3211 (N_3211,N_332,In_2632);
or U3212 (N_3212,N_1728,N_1500);
and U3213 (N_3213,N_1726,N_1808);
nand U3214 (N_3214,In_580,N_1169);
nand U3215 (N_3215,In_3122,N_1613);
or U3216 (N_3216,N_586,N_1404);
nand U3217 (N_3217,N_1413,N_927);
nand U3218 (N_3218,N_41,N_893);
or U3219 (N_3219,N_110,In_3475);
nor U3220 (N_3220,In_1712,N_1695);
nor U3221 (N_3221,N_71,N_1940);
or U3222 (N_3222,In_3809,In_4487);
or U3223 (N_3223,N_1938,In_4337);
nor U3224 (N_3224,N_1341,N_1407);
and U3225 (N_3225,N_718,In_3207);
or U3226 (N_3226,N_620,In_3779);
nor U3227 (N_3227,N_504,N_1193);
or U3228 (N_3228,In_937,N_919);
nor U3229 (N_3229,N_342,N_1599);
xor U3230 (N_3230,In_1111,In_4630);
or U3231 (N_3231,N_488,In_2872);
and U3232 (N_3232,N_711,N_1438);
xor U3233 (N_3233,In_679,In_2296);
xnor U3234 (N_3234,N_652,In_4803);
nand U3235 (N_3235,In_3286,In_47);
and U3236 (N_3236,N_1080,In_72);
nand U3237 (N_3237,In_3211,In_3177);
xnor U3238 (N_3238,N_781,N_475);
nor U3239 (N_3239,In_3736,N_482);
xor U3240 (N_3240,N_989,N_410);
and U3241 (N_3241,N_1319,N_1911);
and U3242 (N_3242,N_1648,N_1210);
nand U3243 (N_3243,N_1397,N_1795);
nand U3244 (N_3244,N_1194,N_1192);
or U3245 (N_3245,In_1590,N_811);
nand U3246 (N_3246,N_180,N_1161);
nor U3247 (N_3247,N_666,In_2043);
nand U3248 (N_3248,N_1637,In_1675);
nor U3249 (N_3249,In_745,In_4396);
or U3250 (N_3250,In_4128,N_1673);
nand U3251 (N_3251,In_4805,N_1707);
xnor U3252 (N_3252,In_258,N_1417);
or U3253 (N_3253,N_1305,N_1287);
and U3254 (N_3254,In_4116,N_1435);
and U3255 (N_3255,N_1437,In_2657);
or U3256 (N_3256,N_12,N_145);
or U3257 (N_3257,In_2192,N_1380);
and U3258 (N_3258,N_1609,In_272);
nor U3259 (N_3259,N_1620,N_1866);
nand U3260 (N_3260,N_1365,In_2421);
nand U3261 (N_3261,N_1602,N_554);
xnor U3262 (N_3262,In_940,In_1010);
and U3263 (N_3263,In_2341,In_2625);
nand U3264 (N_3264,In_1282,N_1086);
nand U3265 (N_3265,N_1476,N_897);
xnor U3266 (N_3266,N_1340,N_1715);
or U3267 (N_3267,In_3184,N_1014);
and U3268 (N_3268,In_661,N_330);
or U3269 (N_3269,N_561,N_381);
and U3270 (N_3270,N_1748,In_2580);
nand U3271 (N_3271,In_2501,N_1684);
or U3272 (N_3272,N_1481,N_214);
nand U3273 (N_3273,In_2419,In_4149);
or U3274 (N_3274,N_1043,In_148);
xor U3275 (N_3275,In_4152,N_1881);
xnor U3276 (N_3276,N_235,N_1782);
nor U3277 (N_3277,N_1331,N_1312);
and U3278 (N_3278,N_1066,N_852);
xor U3279 (N_3279,In_2069,N_671);
nand U3280 (N_3280,N_98,In_2813);
nor U3281 (N_3281,N_1598,N_1000);
xnor U3282 (N_3282,N_1446,N_169);
or U3283 (N_3283,N_602,N_889);
and U3284 (N_3284,N_1498,In_2874);
and U3285 (N_3285,In_1532,N_311);
xor U3286 (N_3286,N_38,N_593);
and U3287 (N_3287,In_428,N_521);
or U3288 (N_3288,In_3317,In_3674);
or U3289 (N_3289,In_3151,In_2717);
nand U3290 (N_3290,N_1790,N_315);
xnor U3291 (N_3291,N_216,In_2058);
and U3292 (N_3292,N_1474,N_1390);
xor U3293 (N_3293,In_995,N_263);
nand U3294 (N_3294,N_1199,N_1053);
nor U3295 (N_3295,In_2434,N_208);
nand U3296 (N_3296,In_1467,N_181);
nand U3297 (N_3297,N_657,N_1381);
nor U3298 (N_3298,In_1150,In_1471);
nand U3299 (N_3299,In_2204,N_948);
xor U3300 (N_3300,N_982,N_519);
nor U3301 (N_3301,In_2577,N_654);
nand U3302 (N_3302,N_1420,N_329);
nor U3303 (N_3303,In_4736,In_648);
xor U3304 (N_3304,In_3486,N_1765);
xor U3305 (N_3305,N_1630,In_3584);
nor U3306 (N_3306,N_1213,In_2635);
or U3307 (N_3307,N_814,N_431);
xnor U3308 (N_3308,N_556,In_1536);
or U3309 (N_3309,In_2345,N_1320);
nand U3310 (N_3310,N_1585,N_296);
nor U3311 (N_3311,In_4424,In_3725);
xnor U3312 (N_3312,In_622,N_913);
nand U3313 (N_3313,In_2979,N_1356);
or U3314 (N_3314,N_133,N_860);
and U3315 (N_3315,In_4080,In_4707);
and U3316 (N_3316,In_3669,In_139);
and U3317 (N_3317,N_1441,N_1708);
and U3318 (N_3318,N_937,In_2450);
and U3319 (N_3319,N_335,N_1606);
xor U3320 (N_3320,N_1479,N_247);
or U3321 (N_3321,In_4621,In_981);
and U3322 (N_3322,In_241,N_300);
xnor U3323 (N_3323,N_1473,N_988);
xor U3324 (N_3324,N_1447,N_506);
or U3325 (N_3325,In_2521,N_691);
nand U3326 (N_3326,N_207,In_4816);
xor U3327 (N_3327,N_848,N_1974);
xor U3328 (N_3328,N_1260,N_838);
or U3329 (N_3329,In_2474,N_939);
nor U3330 (N_3330,N_1197,In_2906);
xnor U3331 (N_3331,N_1467,N_219);
nor U3332 (N_3332,N_770,In_595);
nor U3333 (N_3333,In_4930,N_1557);
or U3334 (N_3334,N_476,In_2828);
and U3335 (N_3335,In_1272,N_130);
and U3336 (N_3336,N_68,N_877);
nand U3337 (N_3337,N_468,N_260);
xnor U3338 (N_3338,N_1675,N_1916);
and U3339 (N_3339,N_1854,N_131);
nand U3340 (N_3340,N_1809,N_940);
or U3341 (N_3341,N_1315,In_3625);
nor U3342 (N_3342,N_1775,In_2997);
nor U3343 (N_3343,N_1158,N_1195);
or U3344 (N_3344,In_4297,In_1362);
or U3345 (N_3345,N_1562,N_369);
nor U3346 (N_3346,N_1706,In_2457);
nor U3347 (N_3347,N_873,N_655);
nand U3348 (N_3348,N_1036,N_470);
or U3349 (N_3349,N_587,N_177);
and U3350 (N_3350,N_641,N_384);
nand U3351 (N_3351,In_4513,In_935);
or U3352 (N_3352,In_1778,In_1470);
nor U3353 (N_3353,N_1855,N_535);
nor U3354 (N_3354,N_692,N_759);
nand U3355 (N_3355,In_1166,N_1652);
xor U3356 (N_3356,In_81,N_1801);
nand U3357 (N_3357,N_121,In_2093);
and U3358 (N_3358,N_35,In_3388);
and U3359 (N_3359,N_1103,N_1337);
nand U3360 (N_3360,N_1360,N_1052);
and U3361 (N_3361,N_1024,N_533);
nor U3362 (N_3362,N_525,In_1674);
xor U3363 (N_3363,N_454,N_1367);
nor U3364 (N_3364,N_1175,N_872);
nor U3365 (N_3365,N_1016,N_522);
and U3366 (N_3366,N_297,N_1168);
and U3367 (N_3367,N_1131,N_1486);
xor U3368 (N_3368,In_3041,N_1571);
nand U3369 (N_3369,N_283,In_1255);
nor U3370 (N_3370,In_3108,N_1701);
nand U3371 (N_3371,N_95,N_17);
nand U3372 (N_3372,N_51,N_1524);
nand U3373 (N_3373,N_1811,In_395);
nand U3374 (N_3374,N_1722,N_1234);
nand U3375 (N_3375,In_3563,N_555);
nand U3376 (N_3376,N_1592,N_1017);
and U3377 (N_3377,In_1265,N_862);
xnor U3378 (N_3378,N_651,In_2972);
nand U3379 (N_3379,N_1702,In_1036);
xor U3380 (N_3380,N_574,In_1953);
and U3381 (N_3381,N_497,N_1992);
xnor U3382 (N_3382,In_40,In_2225);
nor U3383 (N_3383,N_1737,N_1073);
or U3384 (N_3384,In_3713,In_3626);
and U3385 (N_3385,N_1206,N_1087);
nand U3386 (N_3386,In_4565,In_927);
nand U3387 (N_3387,N_1794,In_3864);
or U3388 (N_3388,N_443,N_957);
nor U3389 (N_3389,N_1139,N_1771);
nand U3390 (N_3390,In_1713,In_1502);
nand U3391 (N_3391,In_3955,N_359);
nor U3392 (N_3392,In_1218,N_1040);
nor U3393 (N_3393,In_4704,N_1202);
nor U3394 (N_3394,N_683,In_1401);
and U3395 (N_3395,In_2903,N_1126);
nand U3396 (N_3396,N_1137,N_86);
nor U3397 (N_3397,N_1215,In_4627);
and U3398 (N_3398,In_3975,N_1744);
nand U3399 (N_3399,N_1906,In_2606);
nor U3400 (N_3400,In_4235,N_1196);
nand U3401 (N_3401,N_690,N_1636);
nand U3402 (N_3402,In_3254,N_698);
and U3403 (N_3403,N_1888,N_1457);
or U3404 (N_3404,In_3892,N_1891);
nand U3405 (N_3405,In_100,N_676);
nand U3406 (N_3406,N_147,N_903);
nand U3407 (N_3407,N_1659,In_3455);
nand U3408 (N_3408,N_866,N_1049);
xnor U3409 (N_3409,In_2332,In_2331);
and U3410 (N_3410,In_3623,N_1678);
xor U3411 (N_3411,N_1824,N_1401);
nor U3412 (N_3412,N_55,In_3219);
nand U3413 (N_3413,In_1289,N_265);
xor U3414 (N_3414,N_157,N_196);
or U3415 (N_3415,In_3258,N_415);
nand U3416 (N_3416,In_524,N_1384);
or U3417 (N_3417,In_68,N_1984);
and U3418 (N_3418,N_1521,N_1147);
and U3419 (N_3419,N_483,N_73);
and U3420 (N_3420,N_346,N_895);
nand U3421 (N_3421,N_715,N_1560);
nor U3422 (N_3422,N_1140,In_899);
and U3423 (N_3423,N_451,N_1915);
nand U3424 (N_3424,N_1455,In_2615);
nor U3425 (N_3425,N_1910,N_1118);
nor U3426 (N_3426,N_1564,N_116);
and U3427 (N_3427,N_1111,N_523);
and U3428 (N_3428,N_305,In_872);
nand U3429 (N_3429,N_1851,N_334);
nor U3430 (N_3430,In_174,N_1788);
xnor U3431 (N_3431,N_694,In_4013);
nor U3432 (N_3432,N_1123,N_566);
xnor U3433 (N_3433,In_4433,In_3681);
and U3434 (N_3434,N_688,N_1388);
nor U3435 (N_3435,N_222,In_490);
nor U3436 (N_3436,In_2970,In_1428);
nand U3437 (N_3437,N_1056,N_627);
and U3438 (N_3438,N_1946,In_486);
xnor U3439 (N_3439,N_686,N_1153);
nand U3440 (N_3440,In_4205,N_1987);
nand U3441 (N_3441,N_105,N_570);
nand U3442 (N_3442,In_1054,In_2443);
nor U3443 (N_3443,N_950,N_1349);
nand U3444 (N_3444,In_3639,In_1236);
xor U3445 (N_3445,N_1506,N_1494);
or U3446 (N_3446,N_709,In_3727);
nor U3447 (N_3447,N_1239,In_4322);
nand U3448 (N_3448,N_61,N_1060);
or U3449 (N_3449,N_137,N_450);
nor U3450 (N_3450,N_1296,N_154);
nand U3451 (N_3451,N_5,N_530);
and U3452 (N_3452,In_268,N_1120);
nor U3453 (N_3453,In_1303,N_1871);
and U3454 (N_3454,N_1253,In_1466);
or U3455 (N_3455,N_637,N_667);
or U3456 (N_3456,In_3895,In_4488);
xor U3457 (N_3457,N_1935,N_1157);
nor U3458 (N_3458,N_656,In_179);
nand U3459 (N_3459,In_4113,In_4852);
or U3460 (N_3460,N_816,N_1416);
nand U3461 (N_3461,N_1064,In_4795);
nand U3462 (N_3462,N_1845,N_259);
nand U3463 (N_3463,In_2552,N_732);
nor U3464 (N_3464,N_992,N_1572);
nor U3465 (N_3465,N_806,N_1688);
nor U3466 (N_3466,N_1162,N_53);
or U3467 (N_3467,N_34,N_961);
or U3468 (N_3468,In_4990,N_1507);
or U3469 (N_3469,N_203,In_818);
nor U3470 (N_3470,In_3772,N_1501);
xor U3471 (N_3471,N_737,In_4767);
and U3472 (N_3472,N_1124,In_2722);
nor U3473 (N_3473,N_9,In_1337);
and U3474 (N_3474,N_320,In_4936);
nand U3475 (N_3475,N_1644,N_1256);
nor U3476 (N_3476,N_1797,In_431);
or U3477 (N_3477,In_350,In_4349);
nor U3478 (N_3478,N_1460,N_230);
and U3479 (N_3479,In_4191,N_293);
nor U3480 (N_3480,N_184,N_984);
xnor U3481 (N_3481,In_4015,N_805);
nor U3482 (N_3482,N_1901,In_3789);
nand U3483 (N_3483,In_3482,In_2685);
or U3484 (N_3484,N_256,N_1207);
nand U3485 (N_3485,In_2103,In_4238);
xnor U3486 (N_3486,N_1354,In_2581);
nand U3487 (N_3487,N_726,N_974);
nand U3488 (N_3488,In_4793,N_1576);
nor U3489 (N_3489,In_606,N_853);
and U3490 (N_3490,N_1463,N_1743);
or U3491 (N_3491,In_3937,N_1469);
nor U3492 (N_3492,N_139,N_93);
nand U3493 (N_3493,N_1827,N_780);
nand U3494 (N_3494,N_1044,N_1258);
and U3495 (N_3495,N_484,In_3640);
or U3496 (N_3496,N_1849,N_1787);
nor U3497 (N_3497,N_1746,N_1832);
xnor U3498 (N_3498,In_2,N_4);
and U3499 (N_3499,N_383,In_4140);
nand U3500 (N_3500,N_545,N_1818);
xor U3501 (N_3501,In_3497,N_1238);
xnor U3502 (N_3502,N_491,N_239);
nand U3503 (N_3503,In_1238,In_3858);
xnor U3504 (N_3504,In_4720,In_1080);
and U3505 (N_3505,In_617,N_579);
or U3506 (N_3506,In_3674,N_585);
or U3507 (N_3507,N_550,N_583);
and U3508 (N_3508,N_1081,N_123);
nor U3509 (N_3509,N_792,N_1245);
nand U3510 (N_3510,N_1523,In_4349);
nor U3511 (N_3511,In_2875,In_702);
or U3512 (N_3512,N_1200,N_771);
and U3513 (N_3513,N_640,In_1743);
and U3514 (N_3514,N_1965,N_1346);
nand U3515 (N_3515,In_27,In_1539);
or U3516 (N_3516,N_1075,N_1223);
xor U3517 (N_3517,In_3349,In_4254);
xnor U3518 (N_3518,In_2104,N_1336);
nand U3519 (N_3519,N_1296,In_4730);
or U3520 (N_3520,N_69,In_1236);
xnor U3521 (N_3521,In_1503,N_217);
or U3522 (N_3522,N_0,In_2906);
nand U3523 (N_3523,N_411,In_2324);
and U3524 (N_3524,N_1763,In_139);
nand U3525 (N_3525,N_1059,N_54);
or U3526 (N_3526,N_433,In_4149);
nand U3527 (N_3527,N_1191,N_1692);
and U3528 (N_3528,N_645,N_1024);
xor U3529 (N_3529,N_31,In_3273);
nand U3530 (N_3530,In_377,N_785);
xnor U3531 (N_3531,N_674,N_940);
nand U3532 (N_3532,N_64,N_701);
nand U3533 (N_3533,N_1797,N_246);
xnor U3534 (N_3534,N_1683,In_2580);
or U3535 (N_3535,In_3034,N_1291);
xnor U3536 (N_3536,N_294,N_969);
and U3537 (N_3537,N_477,In_4385);
nor U3538 (N_3538,N_309,N_1070);
nand U3539 (N_3539,In_3480,N_1376);
or U3540 (N_3540,N_86,N_446);
nand U3541 (N_3541,N_450,N_1014);
nand U3542 (N_3542,N_711,N_632);
and U3543 (N_3543,N_1584,N_1452);
xnor U3544 (N_3544,In_3851,In_4106);
or U3545 (N_3545,N_1268,In_2953);
nor U3546 (N_3546,N_17,In_1148);
nand U3547 (N_3547,In_2063,N_1585);
xor U3548 (N_3548,N_707,In_1566);
or U3549 (N_3549,In_3413,N_1322);
or U3550 (N_3550,In_3626,In_1458);
xnor U3551 (N_3551,N_1349,N_782);
and U3552 (N_3552,N_155,N_103);
nand U3553 (N_3553,N_1538,In_294);
and U3554 (N_3554,N_252,N_1706);
nand U3555 (N_3555,In_1421,N_1868);
or U3556 (N_3556,N_995,In_4433);
nand U3557 (N_3557,In_2225,N_1824);
nor U3558 (N_3558,N_1355,N_1922);
or U3559 (N_3559,N_59,N_743);
nor U3560 (N_3560,N_716,N_64);
or U3561 (N_3561,N_1458,N_1963);
or U3562 (N_3562,N_105,N_1022);
nor U3563 (N_3563,N_1523,N_704);
or U3564 (N_3564,N_1559,In_1265);
nor U3565 (N_3565,N_1042,N_1225);
and U3566 (N_3566,In_2469,N_1170);
nand U3567 (N_3567,N_1984,N_23);
xnor U3568 (N_3568,In_3184,N_1691);
nor U3569 (N_3569,N_819,N_718);
and U3570 (N_3570,N_1501,N_274);
and U3571 (N_3571,In_3413,In_4798);
nor U3572 (N_3572,In_3626,N_861);
nand U3573 (N_3573,N_597,N_1866);
nand U3574 (N_3574,N_1250,N_1602);
or U3575 (N_3575,In_4086,N_450);
nand U3576 (N_3576,N_1694,N_711);
or U3577 (N_3577,N_550,N_123);
nor U3578 (N_3578,N_1413,N_1175);
nor U3579 (N_3579,N_499,N_461);
or U3580 (N_3580,In_2204,N_301);
xor U3581 (N_3581,In_649,N_1020);
and U3582 (N_3582,N_52,N_422);
nor U3583 (N_3583,N_243,In_2560);
and U3584 (N_3584,In_2454,N_712);
xor U3585 (N_3585,N_1284,In_4163);
nand U3586 (N_3586,In_3373,N_831);
nand U3587 (N_3587,N_960,In_3207);
and U3588 (N_3588,N_1803,N_1467);
nor U3589 (N_3589,In_3429,N_687);
nor U3590 (N_3590,N_1786,N_1118);
nor U3591 (N_3591,In_4772,N_379);
nand U3592 (N_3592,N_773,N_1845);
nand U3593 (N_3593,N_330,N_729);
xnor U3594 (N_3594,In_4767,In_3987);
nand U3595 (N_3595,N_469,N_1418);
and U3596 (N_3596,N_1084,N_326);
nand U3597 (N_3597,N_1756,N_634);
or U3598 (N_3598,N_989,N_1425);
or U3599 (N_3599,N_1549,In_1532);
nor U3600 (N_3600,In_1318,N_1334);
nand U3601 (N_3601,N_1566,N_1215);
and U3602 (N_3602,N_1196,N_895);
nor U3603 (N_3603,In_2239,In_2864);
nand U3604 (N_3604,N_525,N_914);
nand U3605 (N_3605,N_257,N_1123);
nor U3606 (N_3606,N_1924,N_462);
nor U3607 (N_3607,In_36,N_363);
nor U3608 (N_3608,N_1743,In_4155);
or U3609 (N_3609,N_1849,N_1698);
nand U3610 (N_3610,In_2273,N_853);
nor U3611 (N_3611,N_258,N_827);
nand U3612 (N_3612,In_1256,In_1953);
nand U3613 (N_3613,In_4549,N_822);
nor U3614 (N_3614,In_4672,N_835);
and U3615 (N_3615,N_520,N_1922);
nor U3616 (N_3616,N_166,N_1498);
or U3617 (N_3617,N_442,N_1542);
nor U3618 (N_3618,In_352,N_377);
and U3619 (N_3619,N_1091,N_919);
nand U3620 (N_3620,N_1277,N_196);
or U3621 (N_3621,N_1375,N_1277);
xnor U3622 (N_3622,N_360,In_80);
and U3623 (N_3623,N_116,N_582);
nor U3624 (N_3624,In_239,N_573);
nand U3625 (N_3625,N_1325,N_1020);
xor U3626 (N_3626,N_1555,In_483);
xnor U3627 (N_3627,N_1287,N_1602);
and U3628 (N_3628,In_633,N_91);
nand U3629 (N_3629,N_1639,In_1540);
and U3630 (N_3630,In_4875,N_168);
and U3631 (N_3631,N_1598,In_3193);
or U3632 (N_3632,N_800,In_1041);
xor U3633 (N_3633,N_120,N_390);
and U3634 (N_3634,N_707,N_119);
xor U3635 (N_3635,N_849,N_1808);
or U3636 (N_3636,N_1298,N_479);
nand U3637 (N_3637,N_1509,N_1779);
and U3638 (N_3638,N_1683,N_702);
nand U3639 (N_3639,In_1499,In_286);
or U3640 (N_3640,N_977,N_807);
xnor U3641 (N_3641,In_4888,In_1681);
nor U3642 (N_3642,N_635,In_4930);
and U3643 (N_3643,N_1415,N_1842);
nor U3644 (N_3644,In_2210,N_457);
nor U3645 (N_3645,N_1829,In_4897);
xor U3646 (N_3646,N_1130,In_4600);
xor U3647 (N_3647,N_330,In_239);
nor U3648 (N_3648,N_213,In_1334);
and U3649 (N_3649,N_532,In_4625);
xor U3650 (N_3650,N_1227,In_4066);
or U3651 (N_3651,N_569,N_563);
nand U3652 (N_3652,In_3702,N_1306);
xor U3653 (N_3653,N_1480,In_3429);
nor U3654 (N_3654,In_1322,N_1585);
xnor U3655 (N_3655,N_1068,In_2049);
xor U3656 (N_3656,In_2768,N_1517);
and U3657 (N_3657,In_4182,N_1326);
and U3658 (N_3658,N_367,N_212);
xnor U3659 (N_3659,In_3976,N_219);
nand U3660 (N_3660,In_3345,In_4312);
or U3661 (N_3661,N_157,N_976);
nor U3662 (N_3662,In_4712,N_486);
nor U3663 (N_3663,N_994,N_1422);
nor U3664 (N_3664,N_1934,N_592);
nor U3665 (N_3665,In_4981,N_618);
or U3666 (N_3666,N_1737,In_2664);
or U3667 (N_3667,N_230,N_734);
or U3668 (N_3668,In_1256,In_4965);
or U3669 (N_3669,N_601,N_1618);
nand U3670 (N_3670,In_880,N_1985);
or U3671 (N_3671,N_1300,N_912);
nand U3672 (N_3672,In_3620,N_1378);
xnor U3673 (N_3673,N_1678,N_116);
nand U3674 (N_3674,N_200,N_26);
xnor U3675 (N_3675,N_1959,In_4256);
xnor U3676 (N_3676,N_1405,N_413);
or U3677 (N_3677,N_1033,In_3345);
or U3678 (N_3678,In_4720,N_1069);
nor U3679 (N_3679,In_1330,In_1297);
nand U3680 (N_3680,N_1868,N_1597);
nand U3681 (N_3681,In_148,N_1796);
or U3682 (N_3682,N_1250,N_688);
and U3683 (N_3683,N_926,N_470);
nor U3684 (N_3684,N_482,N_581);
nor U3685 (N_3685,N_1827,N_152);
or U3686 (N_3686,In_1743,N_1664);
nand U3687 (N_3687,In_1324,In_570);
xor U3688 (N_3688,In_4852,N_1920);
xor U3689 (N_3689,N_913,N_695);
and U3690 (N_3690,N_1398,In_431);
nand U3691 (N_3691,In_1675,N_1353);
or U3692 (N_3692,In_1008,N_490);
or U3693 (N_3693,In_2947,N_1648);
nand U3694 (N_3694,In_930,In_187);
nor U3695 (N_3695,In_4349,In_3211);
nor U3696 (N_3696,N_621,N_339);
nor U3697 (N_3697,N_51,N_210);
xnor U3698 (N_3698,N_622,N_1240);
xor U3699 (N_3699,N_1064,N_940);
or U3700 (N_3700,N_1036,In_1323);
nand U3701 (N_3701,N_1212,N_348);
xnor U3702 (N_3702,N_707,In_4292);
or U3703 (N_3703,N_1228,N_325);
nand U3704 (N_3704,N_1671,N_293);
and U3705 (N_3705,N_841,N_881);
and U3706 (N_3706,N_248,N_844);
nor U3707 (N_3707,In_1985,N_1254);
xor U3708 (N_3708,In_3789,In_651);
nor U3709 (N_3709,N_1572,N_840);
or U3710 (N_3710,N_949,In_2104);
xor U3711 (N_3711,In_1454,In_1100);
xor U3712 (N_3712,N_1366,In_940);
xnor U3713 (N_3713,In_3640,N_774);
nor U3714 (N_3714,In_174,N_1901);
nand U3715 (N_3715,In_685,N_733);
nand U3716 (N_3716,N_790,In_2322);
nand U3717 (N_3717,N_41,In_4113);
or U3718 (N_3718,In_4235,In_2560);
and U3719 (N_3719,N_1667,In_3359);
or U3720 (N_3720,In_3609,N_1887);
nand U3721 (N_3721,N_402,In_3681);
nand U3722 (N_3722,In_36,N_1424);
nor U3723 (N_3723,N_1497,N_701);
or U3724 (N_3724,N_19,N_1756);
nor U3725 (N_3725,N_1685,In_4846);
xor U3726 (N_3726,N_1587,N_1117);
nand U3727 (N_3727,N_439,N_1406);
nor U3728 (N_3728,N_539,N_1076);
or U3729 (N_3729,N_1731,N_1574);
nand U3730 (N_3730,N_456,N_124);
xor U3731 (N_3731,N_262,N_1157);
nand U3732 (N_3732,N_1142,N_129);
nand U3733 (N_3733,In_3299,In_1470);
nand U3734 (N_3734,N_649,N_132);
nand U3735 (N_3735,In_1480,N_1424);
nand U3736 (N_3736,N_1201,N_410);
nand U3737 (N_3737,In_3842,N_1866);
and U3738 (N_3738,In_2474,In_649);
nand U3739 (N_3739,In_2632,N_1219);
nor U3740 (N_3740,In_4337,N_281);
xnor U3741 (N_3741,N_1567,N_1993);
or U3742 (N_3742,N_1409,In_4981);
xnor U3743 (N_3743,N_1536,In_4795);
xnor U3744 (N_3744,In_4965,In_4872);
or U3745 (N_3745,N_885,N_1164);
and U3746 (N_3746,N_1693,In_3851);
and U3747 (N_3747,N_1260,N_1206);
xor U3748 (N_3748,N_1962,N_259);
nor U3749 (N_3749,N_511,N_98);
nor U3750 (N_3750,N_650,N_523);
nand U3751 (N_3751,N_1511,N_1004);
xnor U3752 (N_3752,N_1312,N_469);
nor U3753 (N_3753,N_1074,N_1856);
xor U3754 (N_3754,In_1080,N_1303);
xor U3755 (N_3755,N_742,In_427);
nor U3756 (N_3756,N_1129,In_3485);
xor U3757 (N_3757,In_4817,In_2774);
nand U3758 (N_3758,N_1437,N_359);
nor U3759 (N_3759,N_358,N_1073);
and U3760 (N_3760,In_4306,N_1139);
xor U3761 (N_3761,N_679,In_1990);
and U3762 (N_3762,In_4294,In_4160);
nand U3763 (N_3763,In_3404,N_1620);
or U3764 (N_3764,N_612,N_829);
nand U3765 (N_3765,N_918,N_1284);
and U3766 (N_3766,N_277,N_1267);
nor U3767 (N_3767,N_1204,In_4431);
nor U3768 (N_3768,N_1251,N_1804);
nor U3769 (N_3769,In_649,N_1930);
or U3770 (N_3770,N_1240,N_1090);
or U3771 (N_3771,In_3379,N_1964);
and U3772 (N_3772,In_3674,N_857);
nand U3773 (N_3773,N_1411,N_831);
nand U3774 (N_3774,N_365,In_3241);
xnor U3775 (N_3775,In_3905,N_169);
nor U3776 (N_3776,N_915,N_1807);
or U3777 (N_3777,In_4793,N_1270);
or U3778 (N_3778,N_808,N_690);
xnor U3779 (N_3779,In_4322,N_32);
nand U3780 (N_3780,N_1965,In_3759);
or U3781 (N_3781,In_4230,In_3895);
or U3782 (N_3782,N_314,N_326);
nor U3783 (N_3783,N_1331,N_1846);
or U3784 (N_3784,N_1682,In_4306);
and U3785 (N_3785,In_282,N_841);
nor U3786 (N_3786,N_1558,N_984);
and U3787 (N_3787,N_1393,N_722);
nor U3788 (N_3788,In_3592,In_186);
and U3789 (N_3789,N_373,N_324);
or U3790 (N_3790,N_491,N_1676);
or U3791 (N_3791,N_1897,In_3677);
or U3792 (N_3792,N_50,N_1750);
nor U3793 (N_3793,N_749,In_760);
xor U3794 (N_3794,N_1390,N_625);
xor U3795 (N_3795,In_2774,N_147);
and U3796 (N_3796,N_233,In_846);
nand U3797 (N_3797,N_970,N_345);
xnor U3798 (N_3798,N_230,N_1765);
and U3799 (N_3799,In_2580,N_1185);
xnor U3800 (N_3800,N_495,N_654);
or U3801 (N_3801,N_641,N_1776);
nor U3802 (N_3802,N_1808,N_1470);
xor U3803 (N_3803,In_3494,N_1941);
and U3804 (N_3804,N_1696,N_937);
xor U3805 (N_3805,In_3400,N_750);
nand U3806 (N_3806,In_1577,In_1752);
xnor U3807 (N_3807,N_1072,N_1592);
xnor U3808 (N_3808,In_1072,In_3639);
nand U3809 (N_3809,N_680,N_660);
or U3810 (N_3810,In_1784,In_1953);
nor U3811 (N_3811,In_2615,In_3219);
xnor U3812 (N_3812,In_12,N_1233);
xor U3813 (N_3813,N_881,In_2570);
and U3814 (N_3814,In_1208,In_1148);
xor U3815 (N_3815,N_1952,In_4317);
and U3816 (N_3816,N_543,N_896);
nor U3817 (N_3817,N_1755,N_1018);
and U3818 (N_3818,N_1545,N_1844);
nand U3819 (N_3819,N_71,In_4510);
nor U3820 (N_3820,In_2997,N_1867);
and U3821 (N_3821,N_114,N_1190);
nor U3822 (N_3822,In_678,N_1152);
nand U3823 (N_3823,N_1747,N_1021);
or U3824 (N_3824,N_786,In_1280);
xnor U3825 (N_3825,N_295,N_1865);
or U3826 (N_3826,In_2338,In_3089);
nand U3827 (N_3827,N_1614,N_581);
or U3828 (N_3828,N_566,N_1635);
or U3829 (N_3829,In_2363,N_173);
and U3830 (N_3830,N_1665,In_745);
or U3831 (N_3831,In_1350,N_1967);
or U3832 (N_3832,N_1250,In_4431);
or U3833 (N_3833,N_1284,N_376);
or U3834 (N_3834,N_879,N_1761);
nor U3835 (N_3835,N_1428,N_521);
nor U3836 (N_3836,N_296,N_1647);
nand U3837 (N_3837,N_471,N_1159);
nand U3838 (N_3838,N_646,N_1043);
nand U3839 (N_3839,In_2551,N_981);
or U3840 (N_3840,N_880,N_76);
or U3841 (N_3841,N_1555,N_209);
nand U3842 (N_3842,N_382,N_683);
or U3843 (N_3843,In_2704,In_4955);
nor U3844 (N_3844,In_2348,N_316);
nor U3845 (N_3845,N_927,In_2565);
and U3846 (N_3846,N_840,In_396);
xnor U3847 (N_3847,N_1535,N_1683);
and U3848 (N_3848,N_921,N_672);
and U3849 (N_3849,N_373,In_1471);
nor U3850 (N_3850,In_3238,N_129);
and U3851 (N_3851,In_2916,In_3339);
and U3852 (N_3852,N_36,In_2038);
or U3853 (N_3853,In_3410,N_257);
or U3854 (N_3854,N_625,N_1956);
xnor U3855 (N_3855,N_1669,In_1054);
or U3856 (N_3856,In_175,In_1624);
nor U3857 (N_3857,In_3535,N_1824);
xor U3858 (N_3858,In_2993,N_1554);
nand U3859 (N_3859,N_1331,In_1383);
nor U3860 (N_3860,In_1301,In_3211);
or U3861 (N_3861,N_294,In_2531);
and U3862 (N_3862,N_249,N_1762);
or U3863 (N_3863,N_384,N_564);
nand U3864 (N_3864,N_270,N_1648);
xor U3865 (N_3865,N_1881,N_951);
nor U3866 (N_3866,In_2826,N_635);
nand U3867 (N_3867,N_978,N_1548);
nor U3868 (N_3868,In_170,N_1651);
and U3869 (N_3869,N_1328,N_1075);
and U3870 (N_3870,N_1965,In_2182);
or U3871 (N_3871,N_676,N_978);
nor U3872 (N_3872,N_666,N_1559);
nor U3873 (N_3873,In_1036,N_295);
and U3874 (N_3874,N_674,N_1294);
nor U3875 (N_3875,In_152,In_4349);
xnor U3876 (N_3876,N_1260,N_1083);
or U3877 (N_3877,N_527,N_1893);
xnor U3878 (N_3878,N_1901,N_1251);
nand U3879 (N_3879,N_325,In_590);
nand U3880 (N_3880,N_479,N_814);
or U3881 (N_3881,In_886,In_3273);
nor U3882 (N_3882,In_68,In_3535);
xor U3883 (N_3883,N_1579,In_3496);
or U3884 (N_3884,In_4317,N_1093);
and U3885 (N_3885,In_543,N_726);
nand U3886 (N_3886,In_1109,N_821);
or U3887 (N_3887,In_490,In_1497);
nand U3888 (N_3888,In_1498,N_1834);
nor U3889 (N_3889,In_2932,In_553);
or U3890 (N_3890,N_1795,N_1950);
or U3891 (N_3891,In_4938,N_234);
nor U3892 (N_3892,N_405,N_1978);
nand U3893 (N_3893,N_1873,N_1337);
xor U3894 (N_3894,N_1716,N_1928);
nand U3895 (N_3895,N_280,N_1928);
nor U3896 (N_3896,N_1764,N_1886);
xnor U3897 (N_3897,N_1320,In_2695);
and U3898 (N_3898,N_895,N_405);
and U3899 (N_3899,In_4163,N_1702);
nand U3900 (N_3900,N_42,In_4396);
or U3901 (N_3901,In_816,N_495);
nand U3902 (N_3902,N_1202,In_2506);
xor U3903 (N_3903,N_419,N_850);
nand U3904 (N_3904,N_1302,In_633);
nor U3905 (N_3905,N_412,In_1401);
and U3906 (N_3906,N_586,N_295);
nor U3907 (N_3907,In_995,N_1220);
or U3908 (N_3908,In_1876,In_2722);
nand U3909 (N_3909,N_1380,N_232);
nor U3910 (N_3910,N_1031,In_4468);
and U3911 (N_3911,In_4020,N_1633);
and U3912 (N_3912,N_1198,N_1653);
xnor U3913 (N_3913,In_3036,N_24);
and U3914 (N_3914,N_279,In_4214);
nand U3915 (N_3915,N_37,N_387);
nor U3916 (N_3916,N_377,N_1928);
or U3917 (N_3917,In_1933,In_3704);
xnor U3918 (N_3918,N_753,N_139);
and U3919 (N_3919,N_229,In_452);
or U3920 (N_3920,N_241,N_931);
xor U3921 (N_3921,In_3779,N_1152);
xnor U3922 (N_3922,N_191,In_3344);
and U3923 (N_3923,N_202,N_1254);
xnor U3924 (N_3924,In_2717,N_1823);
or U3925 (N_3925,N_360,N_1536);
or U3926 (N_3926,N_1474,N_1044);
nor U3927 (N_3927,In_1713,N_498);
nor U3928 (N_3928,In_4825,N_1559);
xnor U3929 (N_3929,N_1337,N_1572);
and U3930 (N_3930,In_1111,N_582);
or U3931 (N_3931,N_1521,N_401);
nor U3932 (N_3932,N_1068,N_638);
nor U3933 (N_3933,In_1953,N_1815);
xnor U3934 (N_3934,In_930,In_3626);
and U3935 (N_3935,N_1900,N_495);
nor U3936 (N_3936,N_438,N_1959);
nand U3937 (N_3937,In_1282,In_1467);
nor U3938 (N_3938,N_1990,In_352);
nor U3939 (N_3939,N_1146,In_3865);
and U3940 (N_3940,In_1230,In_2585);
nand U3941 (N_3941,N_76,In_3384);
and U3942 (N_3942,N_338,N_19);
or U3943 (N_3943,N_457,N_4);
xnor U3944 (N_3944,N_866,In_1337);
and U3945 (N_3945,In_780,N_153);
nor U3946 (N_3946,N_570,In_4403);
xor U3947 (N_3947,N_298,In_3211);
or U3948 (N_3948,N_1291,In_4433);
and U3949 (N_3949,In_4720,N_251);
or U3950 (N_3950,N_1724,N_950);
and U3951 (N_3951,N_458,In_745);
nor U3952 (N_3952,N_904,N_1745);
nor U3953 (N_3953,N_664,N_1122);
nand U3954 (N_3954,N_1990,N_802);
or U3955 (N_3955,N_419,In_6);
and U3956 (N_3956,N_671,N_1447);
and U3957 (N_3957,In_4445,N_795);
xor U3958 (N_3958,In_651,N_313);
or U3959 (N_3959,In_597,N_1325);
or U3960 (N_3960,N_1527,N_910);
xnor U3961 (N_3961,N_1071,In_2078);
and U3962 (N_3962,N_794,N_689);
xnor U3963 (N_3963,N_867,N_231);
or U3964 (N_3964,N_731,In_3562);
xor U3965 (N_3965,N_378,In_2506);
and U3966 (N_3966,N_829,In_2073);
and U3967 (N_3967,N_508,In_2788);
and U3968 (N_3968,In_4930,N_560);
xnor U3969 (N_3969,N_865,N_1318);
nand U3970 (N_3970,N_1682,N_1961);
or U3971 (N_3971,N_618,N_1615);
and U3972 (N_3972,N_754,N_965);
or U3973 (N_3973,N_329,In_395);
nand U3974 (N_3974,N_44,In_287);
and U3975 (N_3975,In_1314,In_3851);
xnor U3976 (N_3976,N_1576,N_1610);
or U3977 (N_3977,N_88,In_2718);
or U3978 (N_3978,N_1533,N_1182);
nand U3979 (N_3979,In_2058,N_1219);
xor U3980 (N_3980,N_1469,N_390);
nor U3981 (N_3981,N_525,N_877);
nand U3982 (N_3982,N_1223,N_1060);
nor U3983 (N_3983,In_2743,N_80);
nand U3984 (N_3984,N_111,N_1901);
and U3985 (N_3985,In_4385,N_1038);
xor U3986 (N_3986,In_3475,N_1475);
and U3987 (N_3987,N_1534,In_490);
nand U3988 (N_3988,N_613,N_1322);
nor U3989 (N_3989,N_71,N_1508);
or U3990 (N_3990,N_16,In_3714);
nand U3991 (N_3991,In_116,N_15);
nand U3992 (N_3992,N_267,N_291);
or U3993 (N_3993,N_1593,N_1886);
nor U3994 (N_3994,In_4572,N_1155);
and U3995 (N_3995,N_1359,In_2469);
or U3996 (N_3996,N_1392,In_878);
and U3997 (N_3997,In_1387,In_3702);
and U3998 (N_3998,N_1310,N_1089);
nand U3999 (N_3999,N_1534,N_413);
or U4000 (N_4000,N_2491,N_2796);
nand U4001 (N_4001,N_2339,N_2196);
nand U4002 (N_4002,N_2300,N_3023);
xnor U4003 (N_4003,N_3722,N_2839);
nor U4004 (N_4004,N_2228,N_2954);
and U4005 (N_4005,N_3470,N_3820);
xor U4006 (N_4006,N_3448,N_2390);
and U4007 (N_4007,N_2331,N_2577);
nand U4008 (N_4008,N_3889,N_3130);
nor U4009 (N_4009,N_2533,N_2226);
nor U4010 (N_4010,N_2790,N_3561);
nand U4011 (N_4011,N_3222,N_3085);
nand U4012 (N_4012,N_2972,N_2127);
nor U4013 (N_4013,N_3071,N_2673);
xnor U4014 (N_4014,N_3810,N_2111);
xor U4015 (N_4015,N_2478,N_2327);
or U4016 (N_4016,N_2132,N_3236);
nand U4017 (N_4017,N_3855,N_2671);
and U4018 (N_4018,N_3693,N_2801);
or U4019 (N_4019,N_2550,N_2675);
or U4020 (N_4020,N_3166,N_3549);
xnor U4021 (N_4021,N_2823,N_2194);
xor U4022 (N_4022,N_2290,N_2701);
nand U4023 (N_4023,N_3076,N_3501);
or U4024 (N_4024,N_3272,N_2508);
xnor U4025 (N_4025,N_3514,N_3526);
nor U4026 (N_4026,N_3370,N_2587);
nand U4027 (N_4027,N_2286,N_2988);
nor U4028 (N_4028,N_2903,N_3001);
and U4029 (N_4029,N_3535,N_3374);
nor U4030 (N_4030,N_3203,N_2465);
nand U4031 (N_4031,N_2664,N_2383);
xnor U4032 (N_4032,N_2798,N_2430);
nor U4033 (N_4033,N_2287,N_2573);
nand U4034 (N_4034,N_2686,N_3168);
nor U4035 (N_4035,N_3155,N_3079);
xnor U4036 (N_4036,N_3275,N_2984);
nor U4037 (N_4037,N_2642,N_3726);
or U4038 (N_4038,N_3433,N_3224);
nor U4039 (N_4039,N_3848,N_2107);
and U4040 (N_4040,N_2474,N_3537);
or U4041 (N_4041,N_2377,N_3532);
nand U4042 (N_4042,N_2112,N_2313);
or U4043 (N_4043,N_2546,N_3972);
xor U4044 (N_4044,N_3608,N_2494);
or U4045 (N_4045,N_3299,N_2707);
xor U4046 (N_4046,N_3120,N_2514);
nor U4047 (N_4047,N_2650,N_3131);
nor U4048 (N_4048,N_2018,N_3312);
nand U4049 (N_4049,N_3218,N_2855);
and U4050 (N_4050,N_2318,N_2856);
nor U4051 (N_4051,N_2614,N_2044);
xnor U4052 (N_4052,N_2667,N_2901);
nor U4053 (N_4053,N_3636,N_2880);
or U4054 (N_4054,N_3478,N_3183);
nand U4055 (N_4055,N_3248,N_3386);
nand U4056 (N_4056,N_2720,N_3200);
and U4057 (N_4057,N_2053,N_3933);
or U4058 (N_4058,N_2515,N_2610);
and U4059 (N_4059,N_2462,N_2799);
and U4060 (N_4060,N_3682,N_3825);
nand U4061 (N_4061,N_2469,N_3572);
nand U4062 (N_4062,N_2665,N_2236);
xnor U4063 (N_4063,N_3089,N_3714);
or U4064 (N_4064,N_3141,N_3346);
or U4065 (N_4065,N_2539,N_3372);
nor U4066 (N_4066,N_3839,N_2930);
or U4067 (N_4067,N_2402,N_3775);
xnor U4068 (N_4068,N_3685,N_3264);
xor U4069 (N_4069,N_2365,N_2633);
nor U4070 (N_4070,N_2865,N_3813);
and U4071 (N_4071,N_3475,N_2682);
nor U4072 (N_4072,N_2177,N_3927);
and U4073 (N_4073,N_2618,N_2354);
nand U4074 (N_4074,N_3195,N_3690);
and U4075 (N_4075,N_3362,N_2916);
or U4076 (N_4076,N_3755,N_3129);
and U4077 (N_4077,N_2987,N_3186);
nor U4078 (N_4078,N_3842,N_3024);
or U4079 (N_4079,N_3145,N_3122);
and U4080 (N_4080,N_3782,N_2522);
and U4081 (N_4081,N_2595,N_3093);
nor U4082 (N_4082,N_2946,N_3245);
xor U4083 (N_4083,N_3391,N_3663);
nor U4084 (N_4084,N_3880,N_2303);
xnor U4085 (N_4085,N_2911,N_3647);
nor U4086 (N_4086,N_3361,N_2311);
xor U4087 (N_4087,N_2291,N_3033);
and U4088 (N_4088,N_2548,N_2378);
or U4089 (N_4089,N_3159,N_2983);
nand U4090 (N_4090,N_3253,N_3907);
xnor U4091 (N_4091,N_2951,N_2051);
and U4092 (N_4092,N_2990,N_2712);
nand U4093 (N_4093,N_3548,N_3597);
nor U4094 (N_4094,N_2456,N_3136);
and U4095 (N_4095,N_2922,N_3844);
or U4096 (N_4096,N_3288,N_3291);
nor U4097 (N_4097,N_2971,N_3623);
and U4098 (N_4098,N_3861,N_2649);
nor U4099 (N_4099,N_3396,N_2769);
xnor U4100 (N_4100,N_2192,N_2031);
xnor U4101 (N_4101,N_2221,N_2679);
or U4102 (N_4102,N_3858,N_2117);
or U4103 (N_4103,N_3923,N_3679);
or U4104 (N_4104,N_2909,N_2738);
and U4105 (N_4105,N_2863,N_3883);
or U4106 (N_4106,N_3963,N_3571);
xor U4107 (N_4107,N_3014,N_3527);
nand U4108 (N_4108,N_2298,N_3828);
and U4109 (N_4109,N_3773,N_2939);
nor U4110 (N_4110,N_2635,N_3010);
nand U4111 (N_4111,N_3891,N_3857);
and U4112 (N_4112,N_3701,N_3601);
or U4113 (N_4113,N_2688,N_2078);
xor U4114 (N_4114,N_2316,N_3211);
xnor U4115 (N_4115,N_2200,N_3022);
xnor U4116 (N_4116,N_2892,N_2778);
nor U4117 (N_4117,N_2022,N_3710);
and U4118 (N_4118,N_2234,N_2332);
nand U4119 (N_4119,N_2202,N_2597);
and U4120 (N_4120,N_2160,N_3332);
or U4121 (N_4121,N_3622,N_3890);
nor U4122 (N_4122,N_3283,N_3951);
and U4123 (N_4123,N_3078,N_2070);
xnor U4124 (N_4124,N_2807,N_2048);
and U4125 (N_4125,N_3105,N_3335);
and U4126 (N_4126,N_2077,N_3431);
nor U4127 (N_4127,N_3325,N_3399);
or U4128 (N_4128,N_3720,N_2400);
and U4129 (N_4129,N_3653,N_2047);
or U4130 (N_4130,N_3438,N_2168);
xnor U4131 (N_4131,N_3670,N_3735);
and U4132 (N_4132,N_3007,N_2690);
nor U4133 (N_4133,N_3512,N_3991);
nor U4134 (N_4134,N_2235,N_3134);
xnor U4135 (N_4135,N_2536,N_2069);
and U4136 (N_4136,N_2758,N_3037);
and U4137 (N_4137,N_2967,N_3903);
nand U4138 (N_4138,N_3468,N_2143);
nor U4139 (N_4139,N_3942,N_3323);
nand U4140 (N_4140,N_2569,N_3841);
and U4141 (N_4141,N_2065,N_3429);
nor U4142 (N_4142,N_3821,N_3551);
nand U4143 (N_4143,N_2579,N_2193);
and U4144 (N_4144,N_2980,N_3713);
nor U4145 (N_4145,N_2099,N_2704);
nand U4146 (N_4146,N_2645,N_3614);
or U4147 (N_4147,N_3260,N_2979);
xor U4148 (N_4148,N_3924,N_3428);
nand U4149 (N_4149,N_3906,N_2443);
and U4150 (N_4150,N_3884,N_2153);
nand U4151 (N_4151,N_3294,N_3455);
and U4152 (N_4152,N_2628,N_2680);
nor U4153 (N_4153,N_2986,N_2534);
nor U4154 (N_4154,N_2350,N_3485);
and U4155 (N_4155,N_2155,N_3314);
xnor U4156 (N_4156,N_2437,N_2853);
and U4157 (N_4157,N_2557,N_3724);
nor U4158 (N_4158,N_3000,N_3021);
nor U4159 (N_4159,N_2060,N_3158);
and U4160 (N_4160,N_2761,N_3520);
or U4161 (N_4161,N_2231,N_2876);
or U4162 (N_4162,N_3055,N_3987);
and U4163 (N_4163,N_3958,N_3792);
and U4164 (N_4164,N_2483,N_2413);
or U4165 (N_4165,N_2562,N_2934);
and U4166 (N_4166,N_3280,N_2423);
and U4167 (N_4167,N_2419,N_2493);
and U4168 (N_4168,N_2725,N_3197);
nand U4169 (N_4169,N_3832,N_3424);
nor U4170 (N_4170,N_3181,N_2399);
nor U4171 (N_4171,N_2741,N_3081);
nor U4172 (N_4172,N_3586,N_2576);
nand U4173 (N_4173,N_2189,N_2715);
or U4174 (N_4174,N_2841,N_2962);
nor U4175 (N_4175,N_3780,N_3519);
xnor U4176 (N_4176,N_3761,N_2232);
xor U4177 (N_4177,N_2084,N_3384);
or U4178 (N_4178,N_2292,N_2808);
and U4179 (N_4179,N_3799,N_3975);
and U4180 (N_4180,N_2792,N_3917);
nand U4181 (N_4181,N_3699,N_2085);
nand U4182 (N_4182,N_2861,N_2130);
nand U4183 (N_4183,N_3811,N_3725);
nor U4184 (N_4184,N_2583,N_3979);
nand U4185 (N_4185,N_2834,N_3496);
nand U4186 (N_4186,N_2388,N_2382);
xor U4187 (N_4187,N_3938,N_2280);
nand U4188 (N_4188,N_3460,N_2184);
xor U4189 (N_4189,N_3697,N_2752);
nand U4190 (N_4190,N_2237,N_3498);
xor U4191 (N_4191,N_2724,N_2634);
nor U4192 (N_4192,N_3711,N_3913);
or U4193 (N_4193,N_3030,N_2197);
xor U4194 (N_4194,N_3749,N_3149);
or U4195 (N_4195,N_2185,N_2561);
xnor U4196 (N_4196,N_2136,N_3759);
and U4197 (N_4197,N_2073,N_2497);
xnor U4198 (N_4198,N_3590,N_2697);
or U4199 (N_4199,N_3150,N_2054);
nor U4200 (N_4200,N_2385,N_2351);
and U4201 (N_4201,N_2789,N_2281);
nand U4202 (N_4202,N_3268,N_3694);
xnor U4203 (N_4203,N_3124,N_3015);
nand U4204 (N_4204,N_3087,N_2468);
nand U4205 (N_4205,N_2767,N_2267);
nor U4206 (N_4206,N_2708,N_2369);
xor U4207 (N_4207,N_3503,N_2006);
nand U4208 (N_4208,N_3178,N_3067);
nand U4209 (N_4209,N_2874,N_2294);
nand U4210 (N_4210,N_2190,N_2486);
xnor U4211 (N_4211,N_2981,N_3566);
xnor U4212 (N_4212,N_3579,N_3354);
nor U4213 (N_4213,N_2081,N_2306);
xnor U4214 (N_4214,N_3407,N_2580);
nand U4215 (N_4215,N_3558,N_3649);
or U4216 (N_4216,N_2948,N_2623);
xnor U4217 (N_4217,N_2241,N_3040);
and U4218 (N_4218,N_3457,N_3472);
nor U4219 (N_4219,N_3625,N_3494);
xnor U4220 (N_4220,N_2955,N_2887);
nand U4221 (N_4221,N_3032,N_2146);
or U4222 (N_4222,N_2427,N_3121);
xnor U4223 (N_4223,N_2588,N_3247);
xor U4224 (N_4224,N_3507,N_2334);
xor U4225 (N_4225,N_2276,N_3106);
or U4226 (N_4226,N_3464,N_2510);
and U4227 (N_4227,N_3479,N_3188);
or U4228 (N_4228,N_2342,N_2651);
xor U4229 (N_4229,N_2250,N_2709);
xnor U4230 (N_4230,N_3244,N_3591);
xnor U4231 (N_4231,N_3595,N_3053);
or U4232 (N_4232,N_2366,N_2348);
and U4233 (N_4233,N_3117,N_2940);
nand U4234 (N_4234,N_3737,N_3176);
nor U4235 (N_4235,N_3426,N_3538);
nor U4236 (N_4236,N_3905,N_3356);
xor U4237 (N_4237,N_2520,N_3669);
or U4238 (N_4238,N_3400,N_3871);
nand U4239 (N_4239,N_3994,N_2964);
nor U4240 (N_4240,N_3285,N_3046);
nand U4241 (N_4241,N_3812,N_2428);
nor U4242 (N_4242,N_2759,N_2252);
nor U4243 (N_4243,N_3147,N_3047);
nor U4244 (N_4244,N_2459,N_3539);
and U4245 (N_4245,N_2182,N_3565);
xor U4246 (N_4246,N_2397,N_3350);
nand U4247 (N_4247,N_2321,N_2319);
and U4248 (N_4248,N_2858,N_2043);
nor U4249 (N_4249,N_3066,N_3297);
xnor U4250 (N_4250,N_2017,N_3419);
and U4251 (N_4251,N_2379,N_3859);
and U4252 (N_4252,N_3199,N_3395);
nand U4253 (N_4253,N_2411,N_2114);
or U4254 (N_4254,N_2552,N_3352);
and U4255 (N_4255,N_3179,N_3008);
xnor U4256 (N_4256,N_2162,N_3368);
nor U4257 (N_4257,N_3529,N_2918);
or U4258 (N_4258,N_2502,N_3326);
nand U4259 (N_4259,N_2582,N_2737);
nor U4260 (N_4260,N_3205,N_3988);
xnor U4261 (N_4261,N_3144,N_3768);
xnor U4262 (N_4262,N_3808,N_3961);
xnor U4263 (N_4263,N_3300,N_3570);
and U4264 (N_4264,N_2100,N_2326);
nor U4265 (N_4265,N_2304,N_3341);
and U4266 (N_4266,N_3292,N_3483);
or U4267 (N_4267,N_3355,N_3269);
nand U4268 (N_4268,N_2061,N_3417);
and U4269 (N_4269,N_2056,N_2008);
and U4270 (N_4270,N_2821,N_2819);
or U4271 (N_4271,N_2612,N_2352);
and U4272 (N_4272,N_3238,N_2249);
or U4273 (N_4273,N_2760,N_2615);
xor U4274 (N_4274,N_3692,N_3152);
or U4275 (N_4275,N_2782,N_2521);
nor U4276 (N_4276,N_2938,N_2825);
and U4277 (N_4277,N_3282,N_2270);
or U4278 (N_4278,N_2009,N_2970);
nand U4279 (N_4279,N_2818,N_2275);
nor U4280 (N_4280,N_3042,N_2072);
or U4281 (N_4281,N_3641,N_2963);
xor U4282 (N_4282,N_2862,N_3660);
nand U4283 (N_4283,N_2133,N_2450);
or U4284 (N_4284,N_3101,N_3786);
nor U4285 (N_4285,N_3086,N_2581);
or U4286 (N_4286,N_3926,N_3174);
nand U4287 (N_4287,N_2007,N_2713);
nand U4288 (N_4288,N_3655,N_3580);
nand U4289 (N_4289,N_2937,N_2343);
and U4290 (N_4290,N_2297,N_2148);
or U4291 (N_4291,N_2183,N_3754);
nor U4292 (N_4292,N_2999,N_3657);
nand U4293 (N_4293,N_3788,N_3111);
and U4294 (N_4294,N_2105,N_3599);
and U4295 (N_4295,N_2362,N_2519);
nand U4296 (N_4296,N_2974,N_2392);
nor U4297 (N_4297,N_3928,N_3600);
nor U4298 (N_4298,N_3207,N_2822);
nand U4299 (N_4299,N_2433,N_2259);
or U4300 (N_4300,N_3638,N_3517);
xor U4301 (N_4301,N_2142,N_2703);
xor U4302 (N_4302,N_2295,N_3072);
nor U4303 (N_4303,N_3977,N_3540);
nand U4304 (N_4304,N_2487,N_3865);
nand U4305 (N_4305,N_2416,N_3045);
or U4306 (N_4306,N_3895,N_3187);
or U4307 (N_4307,N_3161,N_3826);
and U4308 (N_4308,N_2625,N_3080);
nor U4309 (N_4309,N_3829,N_3474);
nor U4310 (N_4310,N_3437,N_2010);
nand U4311 (N_4311,N_3304,N_3967);
nand U4312 (N_4312,N_2565,N_3133);
xor U4313 (N_4313,N_2154,N_3613);
nor U4314 (N_4314,N_3665,N_2138);
and U4315 (N_4315,N_2076,N_3879);
nand U4316 (N_4316,N_3730,N_3393);
xor U4317 (N_4317,N_3367,N_3289);
and U4318 (N_4318,N_2609,N_3688);
xor U4319 (N_4319,N_2532,N_3843);
xnor U4320 (N_4320,N_2716,N_2932);
or U4321 (N_4321,N_3633,N_3956);
or U4322 (N_4322,N_3899,N_3965);
nand U4323 (N_4323,N_2421,N_2898);
or U4324 (N_4324,N_3313,N_2784);
nor U4325 (N_4325,N_2384,N_2444);
and U4326 (N_4326,N_2263,N_3493);
or U4327 (N_4327,N_2541,N_2832);
nor U4328 (N_4328,N_3056,N_2216);
xnor U4329 (N_4329,N_3266,N_3999);
nand U4330 (N_4330,N_2118,N_2302);
nand U4331 (N_4331,N_2406,N_2936);
nand U4332 (N_4332,N_2360,N_2198);
xnor U4333 (N_4333,N_2770,N_2886);
and U4334 (N_4334,N_2410,N_2809);
xor U4335 (N_4335,N_3962,N_3034);
nand U4336 (N_4336,N_2944,N_3769);
nand U4337 (N_4337,N_3993,N_3547);
nand U4338 (N_4338,N_2544,N_2900);
or U4339 (N_4339,N_2700,N_3126);
or U4340 (N_4340,N_3827,N_3220);
or U4341 (N_4341,N_3968,N_3976);
xor U4342 (N_4342,N_2030,N_3921);
and U4343 (N_4343,N_2191,N_2501);
and U4344 (N_4344,N_3552,N_3434);
or U4345 (N_4345,N_2890,N_3744);
xor U4346 (N_4346,N_2338,N_2897);
xor U4347 (N_4347,N_2919,N_3427);
nor U4348 (N_4348,N_3886,N_2079);
nand U4349 (N_4349,N_2641,N_2035);
nand U4350 (N_4350,N_3302,N_2921);
or U4351 (N_4351,N_2847,N_3898);
and U4352 (N_4352,N_3398,N_3381);
nand U4353 (N_4353,N_2367,N_2206);
nand U4354 (N_4354,N_3217,N_3945);
or U4355 (N_4355,N_2696,N_3482);
nand U4356 (N_4356,N_3846,N_2694);
nand U4357 (N_4357,N_3059,N_2066);
nor U4358 (N_4358,N_2572,N_3646);
or U4359 (N_4359,N_3077,N_3379);
nand U4360 (N_4360,N_2850,N_2989);
and U4361 (N_4361,N_2775,N_2749);
nor U4362 (N_4362,N_3619,N_2857);
or U4363 (N_4363,N_3748,N_3643);
xnor U4364 (N_4364,N_2405,N_3049);
nor U4365 (N_4365,N_3318,N_2435);
and U4366 (N_4366,N_2740,N_3787);
xor U4367 (N_4367,N_3981,N_3708);
nand U4368 (N_4368,N_2219,N_2188);
nor U4369 (N_4369,N_3480,N_2414);
xor U4370 (N_4370,N_3011,N_2055);
and U4371 (N_4371,N_2015,N_2826);
or U4372 (N_4372,N_2128,N_3851);
xor U4373 (N_4373,N_2309,N_2663);
xor U4374 (N_4374,N_2558,N_2274);
or U4375 (N_4375,N_2045,N_2417);
or U4376 (N_4376,N_2976,N_3644);
or U4377 (N_4377,N_3955,N_3637);
xnor U4378 (N_4378,N_3454,N_2912);
nand U4379 (N_4379,N_2538,N_3877);
and U4380 (N_4380,N_3330,N_3934);
or U4381 (N_4381,N_3795,N_3013);
xor U4382 (N_4382,N_3860,N_3652);
nand U4383 (N_4383,N_3113,N_3937);
and U4384 (N_4384,N_2179,N_3686);
nor U4385 (N_4385,N_3102,N_3491);
or U4386 (N_4386,N_3233,N_2455);
and U4387 (N_4387,N_3574,N_3170);
and U4388 (N_4388,N_2346,N_3522);
xnor U4389 (N_4389,N_2285,N_3068);
and U4390 (N_4390,N_3192,N_2959);
nand U4391 (N_4391,N_3242,N_3835);
and U4392 (N_4392,N_2600,N_2658);
or U4393 (N_4393,N_2093,N_3505);
and U4394 (N_4394,N_2668,N_3684);
and U4395 (N_4395,N_3734,N_2159);
nor U4396 (N_4396,N_2124,N_2968);
nand U4397 (N_4397,N_2779,N_3700);
xor U4398 (N_4398,N_2748,N_3495);
xnor U4399 (N_4399,N_2842,N_3589);
nand U4400 (N_4400,N_3626,N_3901);
nand U4401 (N_4401,N_2906,N_2699);
xor U4402 (N_4402,N_3277,N_2120);
nor U4403 (N_4403,N_3621,N_2261);
or U4404 (N_4404,N_2464,N_3984);
xor U4405 (N_4405,N_3971,N_2123);
nand U4406 (N_4406,N_2203,N_2996);
nand U4407 (N_4407,N_3337,N_2262);
and U4408 (N_4408,N_2394,N_3836);
or U4409 (N_4409,N_2205,N_2215);
and U4410 (N_4410,N_3404,N_2644);
nor U4411 (N_4411,N_3567,N_2429);
nor U4412 (N_4412,N_3257,N_2571);
or U4413 (N_4413,N_2355,N_2781);
or U4414 (N_4414,N_2794,N_2335);
nand U4415 (N_4415,N_3593,N_3488);
and U4416 (N_4416,N_2454,N_3462);
or U4417 (N_4417,N_2167,N_3333);
and U4418 (N_4418,N_2806,N_2268);
xnor U4419 (N_4419,N_2064,N_3568);
nand U4420 (N_4420,N_2966,N_3263);
nand U4421 (N_4421,N_3324,N_2604);
and U4422 (N_4422,N_3388,N_3534);
xnor U4423 (N_4423,N_2214,N_2670);
nand U4424 (N_4424,N_3058,N_3027);
or U4425 (N_4425,N_2095,N_3656);
xor U4426 (N_4426,N_2509,N_2695);
and U4427 (N_4427,N_2305,N_3894);
or U4428 (N_4428,N_2042,N_3029);
or U4429 (N_4429,N_3414,N_3351);
and U4430 (N_4430,N_3736,N_3246);
or U4431 (N_4431,N_3947,N_3801);
or U4432 (N_4432,N_2499,N_3838);
nand U4433 (N_4433,N_3774,N_3609);
or U4434 (N_4434,N_2540,N_3112);
nand U4435 (N_4435,N_2917,N_3718);
or U4436 (N_4436,N_2638,N_3756);
nor U4437 (N_4437,N_3006,N_2098);
and U4438 (N_4438,N_3138,N_2253);
xnor U4439 (N_4439,N_3467,N_3132);
nand U4440 (N_4440,N_3818,N_2101);
and U4441 (N_4441,N_2889,N_3017);
nor U4442 (N_4442,N_2905,N_2786);
nor U4443 (N_4443,N_3405,N_3051);
or U4444 (N_4444,N_2907,N_2387);
nand U4445 (N_4445,N_3658,N_3212);
and U4446 (N_4446,N_3980,N_2734);
nand U4447 (N_4447,N_3530,N_2357);
nand U4448 (N_4448,N_2706,N_2655);
and U4449 (N_4449,N_2637,N_3882);
and U4450 (N_4450,N_3342,N_2949);
nor U4451 (N_4451,N_2910,N_3797);
or U4452 (N_4452,N_2036,N_3559);
or U4453 (N_4453,N_3941,N_3107);
or U4454 (N_4454,N_3510,N_3721);
and U4455 (N_4455,N_3198,N_2091);
or U4456 (N_4456,N_2029,N_2181);
xnor U4457 (N_4457,N_2283,N_3262);
nor U4458 (N_4458,N_3650,N_3611);
or U4459 (N_4459,N_2915,N_2516);
nand U4460 (N_4460,N_3435,N_2676);
nor U4461 (N_4461,N_3261,N_2144);
nor U4462 (N_4462,N_3343,N_3819);
or U4463 (N_4463,N_3410,N_2445);
or U4464 (N_4464,N_2122,N_3369);
and U4465 (N_4465,N_3594,N_2718);
nor U4466 (N_4466,N_3583,N_3182);
nor U4467 (N_4467,N_2258,N_3635);
and U4468 (N_4468,N_2721,N_3240);
nand U4469 (N_4469,N_2381,N_2756);
nand U4470 (N_4470,N_3847,N_3002);
and U4471 (N_4471,N_3164,N_2157);
nor U4472 (N_4472,N_3208,N_2563);
and U4473 (N_4473,N_3624,N_3698);
or U4474 (N_4474,N_3406,N_2187);
and U4475 (N_4475,N_2458,N_2325);
or U4476 (N_4476,N_3303,N_2424);
nor U4477 (N_4477,N_3536,N_3091);
or U4478 (N_4478,N_3251,N_3604);
nand U4479 (N_4479,N_3508,N_3944);
or U4480 (N_4480,N_2074,N_2380);
nand U4481 (N_4481,N_3885,N_3789);
or U4482 (N_4482,N_3440,N_3691);
xor U4483 (N_4483,N_3123,N_3556);
nand U4484 (N_4484,N_2165,N_2732);
xor U4485 (N_4485,N_2598,N_2204);
or U4486 (N_4486,N_2602,N_2083);
xnor U4487 (N_4487,N_2209,N_3528);
or U4488 (N_4488,N_2643,N_2344);
xnor U4489 (N_4489,N_3321,N_3732);
or U4490 (N_4490,N_3486,N_3290);
or U4491 (N_4491,N_3378,N_2089);
and U4492 (N_4492,N_3151,N_3831);
nor U4493 (N_4493,N_2836,N_2517);
or U4494 (N_4494,N_3546,N_3767);
nor U4495 (N_4495,N_2924,N_3463);
nor U4496 (N_4496,N_3327,N_3778);
xnor U4497 (N_4497,N_3620,N_3616);
nor U4498 (N_4498,N_2866,N_2255);
nand U4499 (N_4499,N_3328,N_3403);
or U4500 (N_4500,N_2058,N_3167);
or U4501 (N_4501,N_2293,N_3715);
nand U4502 (N_4502,N_3824,N_2401);
and U4503 (N_4503,N_3659,N_2004);
xnor U4504 (N_4504,N_3544,N_2882);
nand U4505 (N_4505,N_2141,N_3349);
xor U4506 (N_4506,N_2068,N_2026);
nand U4507 (N_4507,N_2145,N_2172);
nor U4508 (N_4508,N_2272,N_3587);
nor U4509 (N_4509,N_3902,N_3723);
and U4510 (N_4510,N_2403,N_2322);
xnor U4511 (N_4511,N_2929,N_3278);
or U4512 (N_4512,N_2161,N_2931);
or U4513 (N_4513,N_3997,N_3970);
nor U4514 (N_4514,N_2125,N_2434);
nor U4515 (N_4515,N_3003,N_3794);
xor U4516 (N_4516,N_3630,N_2463);
and U4517 (N_4517,N_3109,N_2524);
nand U4518 (N_4518,N_2470,N_3163);
or U4519 (N_4519,N_2186,N_2223);
and U4520 (N_4520,N_3910,N_2363);
nor U4521 (N_4521,N_3243,N_2621);
or U4522 (N_4522,N_2791,N_2933);
xor U4523 (N_4523,N_3250,N_3276);
or U4524 (N_4524,N_2389,N_3385);
or U4525 (N_4525,N_3005,N_3939);
xor U4526 (N_4526,N_2391,N_3557);
xnor U4527 (N_4527,N_3230,N_3293);
or U4528 (N_4528,N_2845,N_2545);
nor U4529 (N_4529,N_3209,N_2827);
and U4530 (N_4530,N_3709,N_3026);
or U4531 (N_4531,N_3617,N_3985);
xor U4532 (N_4532,N_3770,N_2991);
and U4533 (N_4533,N_3518,N_2032);
or U4534 (N_4534,N_3745,N_2368);
xnor U4535 (N_4535,N_2109,N_2174);
nor U4536 (N_4536,N_2594,N_3603);
nor U4537 (N_4537,N_3430,N_2956);
and U4538 (N_4538,N_3450,N_3201);
xor U4539 (N_4539,N_2687,N_3870);
nor U4540 (N_4540,N_2337,N_2977);
or U4541 (N_4541,N_3389,N_3990);
nor U4542 (N_4542,N_3872,N_2549);
nor U4543 (N_4543,N_3607,N_3009);
xor U4544 (N_4544,N_3099,N_2038);
and U4545 (N_4545,N_2207,N_2952);
and U4546 (N_4546,N_2998,N_2049);
nor U4547 (N_4547,N_3190,N_2817);
nand U4548 (N_4548,N_3733,N_2605);
xnor U4549 (N_4549,N_3418,N_2766);
or U4550 (N_4550,N_3998,N_3764);
xnor U4551 (N_4551,N_3950,N_2590);
xor U4552 (N_4552,N_2958,N_2438);
nor U4553 (N_4553,N_2374,N_2927);
nand U4554 (N_4554,N_3800,N_2554);
or U4555 (N_4555,N_2506,N_3531);
or U4556 (N_4556,N_2376,N_2624);
and U4557 (N_4557,N_2978,N_2877);
nand U4558 (N_4558,N_3717,N_3281);
xor U4559 (N_4559,N_3887,N_3545);
nand U4560 (N_4560,N_2875,N_2531);
and U4561 (N_4561,N_2620,N_2152);
or U4562 (N_4562,N_2714,N_3206);
xnor U4563 (N_4563,N_3995,N_2677);
nand U4564 (N_4564,N_3864,N_2489);
and U4565 (N_4565,N_3409,N_3516);
nor U4566 (N_4566,N_3863,N_3287);
or U4567 (N_4567,N_3402,N_2619);
and U4568 (N_4568,N_2717,N_2868);
xnor U4569 (N_4569,N_3996,N_2243);
nand U4570 (N_4570,N_2247,N_2211);
and U4571 (N_4571,N_3319,N_2659);
nand U4572 (N_4572,N_3500,N_3322);
nor U4573 (N_4573,N_3922,N_3931);
or U4574 (N_4574,N_2525,N_2733);
and U4575 (N_4575,N_3173,N_2224);
xnor U4576 (N_4576,N_2359,N_2500);
and U4577 (N_4577,N_3598,N_2830);
nand U4578 (N_4578,N_2025,N_3443);
xnor U4579 (N_4579,N_3873,N_3779);
nand U4580 (N_4580,N_2097,N_2340);
xnor U4581 (N_4581,N_2129,N_3477);
nor U4582 (N_4582,N_3569,N_3874);
nor U4583 (N_4583,N_2094,N_3554);
nand U4584 (N_4584,N_2816,N_3807);
or U4585 (N_4585,N_2831,N_3627);
and U4586 (N_4586,N_3237,N_3274);
or U4587 (N_4587,N_3681,N_2764);
nor U4588 (N_4588,N_3359,N_2728);
nand U4589 (N_4589,N_3949,N_3677);
nor U4590 (N_4590,N_3436,N_2710);
nand U4591 (N_4591,N_3515,N_2961);
nand U4592 (N_4592,N_3075,N_3357);
or U4593 (N_4593,N_3581,N_2037);
or U4594 (N_4594,N_3084,N_3364);
and U4595 (N_4595,N_3191,N_2632);
nand U4596 (N_4596,N_3284,N_3142);
nand U4597 (N_4597,N_3948,N_2902);
and U4598 (N_4598,N_2126,N_2601);
and U4599 (N_4599,N_3560,N_3696);
nand U4600 (N_4600,N_2745,N_3766);
xor U4601 (N_4601,N_3823,N_2119);
nor U4602 (N_4602,N_2904,N_3451);
or U4603 (N_4603,N_2333,N_2838);
xnor U4604 (N_4604,N_2373,N_3849);
nor U4605 (N_4605,N_3576,N_2033);
nand U4606 (N_4606,N_2592,N_3671);
nand U4607 (N_4607,N_2505,N_3762);
xor U4608 (N_4608,N_3753,N_2953);
or U4609 (N_4609,N_3110,N_2894);
and U4610 (N_4610,N_3573,N_3490);
xor U4611 (N_4611,N_2852,N_3978);
and U4612 (N_4612,N_2451,N_3249);
and U4613 (N_4613,N_3973,N_2086);
and U4614 (N_4614,N_2498,N_2150);
and U4615 (N_4615,N_2507,N_2776);
xor U4616 (N_4616,N_3954,N_2567);
or U4617 (N_4617,N_3893,N_2242);
or U4618 (N_4618,N_2908,N_2518);
xnor U4619 (N_4619,N_2636,N_2484);
or U4620 (N_4620,N_3004,N_3504);
and U4621 (N_4621,N_3259,N_2442);
or U4622 (N_4622,N_2575,N_2349);
nand U4623 (N_4623,N_2608,N_2482);
nand U4624 (N_4624,N_2011,N_2260);
nand U4625 (N_4625,N_3983,N_2492);
or U4626 (N_4626,N_3061,N_3177);
or U4627 (N_4627,N_3674,N_2846);
or U4628 (N_4628,N_2001,N_2364);
nor U4629 (N_4629,N_3331,N_2729);
xor U4630 (N_4630,N_3137,N_3336);
nand U4631 (N_4631,N_3888,N_2864);
nand U4632 (N_4632,N_2899,N_3064);
nand U4633 (N_4633,N_2308,N_2739);
nand U4634 (N_4634,N_3592,N_2755);
nand U4635 (N_4635,N_3964,N_3096);
and U4636 (N_4636,N_3830,N_3969);
nor U4637 (N_4637,N_3408,N_2137);
nand U4638 (N_4638,N_3392,N_3308);
nand U4639 (N_4639,N_3146,N_2108);
and U4640 (N_4640,N_3306,N_2418);
xor U4641 (N_4641,N_2477,N_2914);
nand U4642 (N_4642,N_2736,N_3940);
and U4643 (N_4643,N_3044,N_3194);
and U4644 (N_4644,N_2656,N_3310);
or U4645 (N_4645,N_3311,N_3533);
nor U4646 (N_4646,N_3175,N_3481);
nor U4647 (N_4647,N_2166,N_3654);
nor U4648 (N_4648,N_3116,N_2568);
nor U4649 (N_4649,N_3960,N_3673);
nor U4650 (N_4650,N_2772,N_3866);
and U4651 (N_4651,N_3239,N_2751);
nand U4652 (N_4652,N_2969,N_3666);
nor U4653 (N_4653,N_2448,N_3878);
and U4654 (N_4654,N_3702,N_2254);
nand U4655 (N_4655,N_3449,N_3966);
and U4656 (N_4656,N_2844,N_3041);
xnor U4657 (N_4657,N_2092,N_2475);
nor U4658 (N_4658,N_2812,N_2747);
nand U4659 (N_4659,N_3425,N_3153);
or U4660 (N_4660,N_3348,N_2062);
xnor U4661 (N_4661,N_2467,N_2870);
or U4662 (N_4662,N_3751,N_2626);
and U4663 (N_4663,N_2820,N_3252);
nor U4664 (N_4664,N_2674,N_3642);
nor U4665 (N_4665,N_3513,N_3063);
and U4666 (N_4666,N_3171,N_3588);
and U4667 (N_4667,N_2630,N_3585);
or U4668 (N_4668,N_3582,N_3852);
and U4669 (N_4669,N_2684,N_2372);
nor U4670 (N_4670,N_2071,N_3128);
nor U4671 (N_4671,N_2420,N_3634);
nand U4672 (N_4672,N_3676,N_2040);
nand U4673 (N_4673,N_2441,N_2815);
nor U4674 (N_4674,N_2471,N_2324);
xnor U4675 (N_4675,N_2757,N_3876);
nor U4676 (N_4676,N_3667,N_3420);
or U4677 (N_4677,N_3881,N_3459);
and U4678 (N_4678,N_3664,N_2257);
nand U4679 (N_4679,N_2396,N_3421);
xnor U4680 (N_4680,N_2398,N_2472);
and U4681 (N_4681,N_3255,N_2301);
xnor U4682 (N_4682,N_2681,N_3380);
or U4683 (N_4683,N_2878,N_2829);
xnor U4684 (N_4684,N_2345,N_3296);
and U4685 (N_4685,N_3550,N_2965);
nand U4686 (N_4686,N_2103,N_2941);
nor U4687 (N_4687,N_3946,N_2982);
nand U4688 (N_4688,N_2669,N_2885);
nor U4689 (N_4689,N_3705,N_3837);
xor U4690 (N_4690,N_2329,N_2251);
nor U4691 (N_4691,N_2457,N_2763);
nor U4692 (N_4692,N_3932,N_3584);
or U4693 (N_4693,N_2800,N_3048);
nor U4694 (N_4694,N_2530,N_3982);
xnor U4695 (N_4695,N_2238,N_2408);
nor U4696 (N_4696,N_2135,N_3444);
xor U4697 (N_4697,N_3542,N_3305);
or U4698 (N_4698,N_2473,N_3119);
xor U4699 (N_4699,N_3760,N_3668);
nand U4700 (N_4700,N_2404,N_2893);
or U4701 (N_4701,N_2947,N_2840);
xor U4702 (N_4702,N_3069,N_3817);
nor U4703 (N_4703,N_2328,N_3555);
and U4704 (N_4704,N_2210,N_2320);
nand U4705 (N_4705,N_2466,N_2754);
nand U4706 (N_4706,N_2178,N_3763);
nand U4707 (N_4707,N_3750,N_3118);
and U4708 (N_4708,N_3757,N_3258);
xor U4709 (N_4709,N_2426,N_3360);
nor U4710 (N_4710,N_2797,N_3062);
and U4711 (N_4711,N_2529,N_2994);
and U4712 (N_4712,N_3390,N_3856);
nor U4713 (N_4713,N_3340,N_2310);
xor U4714 (N_4714,N_3095,N_3606);
nand U4715 (N_4715,N_3031,N_3316);
and U4716 (N_4716,N_2024,N_2526);
xor U4717 (N_4717,N_2692,N_3651);
xor U4718 (N_4718,N_2593,N_2678);
xnor U4719 (N_4719,N_3154,N_3804);
nor U4720 (N_4720,N_3675,N_2742);
nor U4721 (N_4721,N_2851,N_2431);
nand U4722 (N_4722,N_3957,N_2553);
and U4723 (N_4723,N_3541,N_2660);
and U4724 (N_4724,N_3054,N_2768);
or U4725 (N_4725,N_3104,N_2727);
or U4726 (N_4726,N_3256,N_2985);
and U4727 (N_4727,N_3752,N_2005);
nor U4728 (N_4728,N_2386,N_2395);
and U4729 (N_4729,N_2648,N_3456);
nand U4730 (N_4730,N_3043,N_2244);
and U4731 (N_4731,N_2719,N_3036);
nor U4732 (N_4732,N_3267,N_2314);
nor U4733 (N_4733,N_3092,N_2859);
or U4734 (N_4734,N_3487,N_2928);
nand U4735 (N_4735,N_3785,N_3073);
or U4736 (N_4736,N_2960,N_3344);
nor U4737 (N_4737,N_2811,N_3740);
xnor U4738 (N_4738,N_3432,N_2229);
nand U4739 (N_4739,N_2217,N_3458);
xnor U4740 (N_4740,N_3140,N_2361);
nor U4741 (N_4741,N_3221,N_3814);
or U4742 (N_4742,N_3387,N_3394);
or U4743 (N_4743,N_2810,N_3094);
xnor U4744 (N_4744,N_3125,N_2412);
and U4745 (N_4745,N_3439,N_2485);
xor U4746 (N_4746,N_2131,N_3279);
and U4747 (N_4747,N_2722,N_3645);
and U4748 (N_4748,N_2683,N_3226);
and U4749 (N_4749,N_2233,N_2942);
or U4750 (N_4750,N_2312,N_2096);
nor U4751 (N_4751,N_3184,N_3229);
and U4752 (N_4752,N_3959,N_3577);
nor U4753 (N_4753,N_3484,N_2867);
and U4754 (N_4754,N_2879,N_3553);
and U4755 (N_4755,N_3850,N_2041);
or U4756 (N_4756,N_2195,N_2913);
nand U4757 (N_4757,N_2271,N_2264);
nand U4758 (N_4758,N_2535,N_3050);
nor U4759 (N_4759,N_3900,N_3329);
xor U4760 (N_4760,N_2121,N_3371);
and U4761 (N_4761,N_3445,N_3413);
and U4762 (N_4762,N_3286,N_3758);
xnor U4763 (N_4763,N_2783,N_3989);
nor U4764 (N_4764,N_3992,N_3680);
or U4765 (N_4765,N_2611,N_2672);
or U4766 (N_4766,N_3743,N_2881);
nand U4767 (N_4767,N_3640,N_3090);
nor U4768 (N_4768,N_3366,N_2016);
and U4769 (N_4769,N_3039,N_2787);
xor U4770 (N_4770,N_2299,N_2653);
or U4771 (N_4771,N_2307,N_2613);
nand U4772 (N_4772,N_2503,N_3497);
or U4773 (N_4773,N_2777,N_2814);
nor U4774 (N_4774,N_2460,N_3729);
nand U4775 (N_4775,N_3270,N_3383);
nand U4776 (N_4776,N_2110,N_3727);
nand U4777 (N_4777,N_3943,N_2705);
xnor U4778 (N_4778,N_3315,N_2883);
nand U4779 (N_4779,N_2869,N_2795);
nand U4780 (N_4780,N_3214,N_2992);
xnor U4781 (N_4781,N_2284,N_3025);
xor U4782 (N_4782,N_2622,N_2585);
or U4783 (N_4783,N_3204,N_3716);
xnor U4784 (N_4784,N_3473,N_3605);
nor U4785 (N_4785,N_2584,N_2023);
or U4786 (N_4786,N_2212,N_2631);
nand U4787 (N_4787,N_2425,N_3083);
and U4788 (N_4788,N_3618,N_3628);
xnor U4789 (N_4789,N_3338,N_2277);
xor U4790 (N_4790,N_3575,N_2240);
or U4791 (N_4791,N_3441,N_3213);
and U4792 (N_4792,N_3169,N_2527);
nor U4793 (N_4793,N_2646,N_3307);
or U4794 (N_4794,N_3363,N_2835);
nand U4795 (N_4795,N_3180,N_3615);
and U4796 (N_4796,N_2014,N_2559);
or U4797 (N_4797,N_3422,N_3446);
and U4798 (N_4798,N_3365,N_3953);
nand U4799 (N_4799,N_2773,N_2158);
xnor U4800 (N_4800,N_3678,N_3452);
xnor U4801 (N_4801,N_3100,N_3358);
xnor U4802 (N_4802,N_3115,N_3228);
nor U4803 (N_4803,N_2945,N_2358);
nand U4804 (N_4804,N_2654,N_2218);
or U4805 (N_4805,N_3712,N_2726);
or U4806 (N_4806,N_3929,N_2480);
nand U4807 (N_4807,N_3317,N_3543);
or U4808 (N_4808,N_3020,N_3672);
nor U4809 (N_4809,N_3662,N_3461);
nor U4810 (N_4810,N_2606,N_2266);
nand U4811 (N_4811,N_3816,N_3793);
and U4812 (N_4812,N_2175,N_3074);
nor U4813 (N_4813,N_2731,N_3466);
and U4814 (N_4814,N_3703,N_2698);
or U4815 (N_4815,N_2201,N_3806);
nand U4816 (N_4816,N_2446,N_2488);
nand U4817 (N_4817,N_2828,N_3060);
nor U4818 (N_4818,N_3904,N_3869);
nor U4819 (N_4819,N_2513,N_2082);
and U4820 (N_4820,N_2793,N_2849);
xnor U4821 (N_4821,N_3974,N_2837);
nand U4822 (N_4822,N_2629,N_3235);
xor U4823 (N_4823,N_3098,N_2481);
nor U4824 (N_4824,N_3471,N_2063);
nand U4825 (N_4825,N_3082,N_2341);
nor U4826 (N_4826,N_3273,N_3783);
and U4827 (N_4827,N_3738,N_3661);
and U4828 (N_4828,N_2973,N_2225);
or U4829 (N_4829,N_2273,N_3632);
nor U4830 (N_4830,N_2666,N_2888);
nand U4831 (N_4831,N_2282,N_3704);
or U4832 (N_4832,N_2415,N_3165);
or U4833 (N_4833,N_3822,N_2269);
nand U4834 (N_4834,N_2156,N_2723);
nor U4835 (N_4835,N_3216,N_2000);
nor U4836 (N_4836,N_3796,N_2923);
nor U4837 (N_4837,N_2353,N_3562);
xor U4838 (N_4838,N_2657,N_2511);
and U4839 (N_4839,N_3815,N_2943);
xor U4840 (N_4840,N_2139,N_3227);
or U4841 (N_4841,N_3223,N_2019);
nor U4842 (N_4842,N_2452,N_2265);
nand U4843 (N_4843,N_3376,N_2278);
or U4844 (N_4844,N_2169,N_3231);
and U4845 (N_4845,N_3401,N_3765);
or U4846 (N_4846,N_3524,N_2432);
or U4847 (N_4847,N_2246,N_3345);
xnor U4848 (N_4848,N_2027,N_3952);
or U4849 (N_4849,N_2896,N_2547);
nor U4850 (N_4850,N_2617,N_3375);
or U4851 (N_4851,N_3492,N_2106);
xor U4852 (N_4852,N_3777,N_2685);
and U4853 (N_4853,N_3469,N_3834);
or U4854 (N_4854,N_2453,N_3382);
or U4855 (N_4855,N_2950,N_2616);
and U4856 (N_4856,N_2639,N_3802);
nor U4857 (N_4857,N_3833,N_3706);
or U4858 (N_4858,N_3805,N_2087);
nand U4859 (N_4859,N_2279,N_2804);
and U4860 (N_4860,N_3347,N_2002);
nor U4861 (N_4861,N_3127,N_3511);
nor U4862 (N_4862,N_2208,N_2034);
and U4863 (N_4863,N_2871,N_2461);
and U4864 (N_4864,N_2872,N_3339);
xnor U4865 (N_4865,N_3108,N_3476);
and U4866 (N_4866,N_3232,N_2926);
nor U4867 (N_4867,N_2336,N_2173);
nand U4868 (N_4868,N_3088,N_2599);
nor U4869 (N_4869,N_2711,N_2496);
nand U4870 (N_4870,N_2556,N_2691);
or U4871 (N_4871,N_2935,N_2689);
and U4872 (N_4872,N_3225,N_2028);
xor U4873 (N_4873,N_3747,N_2925);
nor U4874 (N_4874,N_2860,N_2447);
xnor U4875 (N_4875,N_2997,N_2115);
and U4876 (N_4876,N_2230,N_3521);
or U4877 (N_4877,N_3791,N_3234);
nor U4878 (N_4878,N_2164,N_3695);
xnor U4879 (N_4879,N_2735,N_3918);
or U4880 (N_4880,N_3103,N_3509);
or U4881 (N_4881,N_3160,N_3172);
nor U4882 (N_4882,N_3683,N_3502);
and U4883 (N_4883,N_3853,N_2296);
nand U4884 (N_4884,N_2227,N_2080);
xor U4885 (N_4885,N_3930,N_2762);
and U4886 (N_4886,N_3772,N_2957);
xnor U4887 (N_4887,N_3156,N_2134);
nor U4888 (N_4888,N_3602,N_3162);
and U4889 (N_4889,N_3185,N_2199);
and U4890 (N_4890,N_2116,N_3875);
xnor U4891 (N_4891,N_3447,N_3016);
and U4892 (N_4892,N_2113,N_2289);
and U4893 (N_4893,N_3157,N_2090);
or U4894 (N_4894,N_3648,N_2873);
or U4895 (N_4895,N_2422,N_3867);
or U4896 (N_4896,N_3892,N_3728);
and U4897 (N_4897,N_2574,N_3453);
or U4898 (N_4898,N_3739,N_3916);
xor U4899 (N_4899,N_2046,N_2409);
nor U4900 (N_4900,N_2693,N_2407);
xor U4901 (N_4901,N_3596,N_2564);
or U4902 (N_4902,N_3784,N_2170);
xor U4903 (N_4903,N_2640,N_2315);
nor U4904 (N_4904,N_3936,N_2371);
nand U4905 (N_4905,N_3809,N_2542);
or U4906 (N_4906,N_2570,N_3320);
nor U4907 (N_4907,N_2020,N_3019);
or U4908 (N_4908,N_2586,N_2780);
and U4909 (N_4909,N_2596,N_2504);
nor U4910 (N_4910,N_3412,N_3397);
nand U4911 (N_4911,N_2566,N_3803);
nor U4912 (N_4912,N_2220,N_2436);
or U4913 (N_4913,N_3038,N_2021);
or U4914 (N_4914,N_3193,N_3241);
xnor U4915 (N_4915,N_3896,N_2843);
and U4916 (N_4916,N_3525,N_2560);
xnor U4917 (N_4917,N_3489,N_2662);
nand U4918 (N_4918,N_2824,N_2356);
nor U4919 (N_4919,N_2746,N_2591);
or U4920 (N_4920,N_3897,N_2180);
xor U4921 (N_4921,N_2555,N_3919);
xor U4922 (N_4922,N_2449,N_2140);
nor U4923 (N_4923,N_3353,N_3499);
nor U4924 (N_4924,N_2088,N_2805);
and U4925 (N_4925,N_3912,N_3719);
nand U4926 (N_4926,N_3854,N_3416);
and U4927 (N_4927,N_2891,N_3629);
nor U4928 (N_4928,N_3202,N_2013);
and U4929 (N_4929,N_2884,N_3035);
and U4930 (N_4930,N_2578,N_3746);
and U4931 (N_4931,N_3707,N_2248);
and U4932 (N_4932,N_3523,N_2059);
nor U4933 (N_4933,N_2607,N_2330);
and U4934 (N_4934,N_3415,N_3210);
nand U4935 (N_4935,N_2039,N_3506);
nor U4936 (N_4936,N_2785,N_2788);
nor U4937 (N_4937,N_3298,N_3689);
xor U4938 (N_4938,N_2323,N_2476);
and U4939 (N_4939,N_2854,N_3411);
nand U4940 (N_4940,N_3271,N_2512);
xnor U4941 (N_4941,N_3143,N_2176);
or U4942 (N_4942,N_3114,N_2213);
or U4943 (N_4943,N_2317,N_3052);
or U4944 (N_4944,N_3776,N_2730);
nand U4945 (N_4945,N_3377,N_3915);
xnor U4946 (N_4946,N_3612,N_2347);
and U4947 (N_4947,N_2744,N_2551);
or U4948 (N_4948,N_2057,N_2147);
nor U4949 (N_4949,N_2848,N_3911);
and U4950 (N_4950,N_3442,N_2102);
xnor U4951 (N_4951,N_3868,N_2003);
xnor U4952 (N_4952,N_2528,N_3610);
and U4953 (N_4953,N_3309,N_2920);
and U4954 (N_4954,N_2490,N_2256);
nand U4955 (N_4955,N_3254,N_2495);
xnor U4956 (N_4956,N_3741,N_2802);
nor U4957 (N_4957,N_2239,N_2995);
nand U4958 (N_4958,N_3935,N_3423);
or U4959 (N_4959,N_3986,N_2895);
or U4960 (N_4960,N_3012,N_2627);
or U4961 (N_4961,N_2765,N_2288);
xnor U4962 (N_4962,N_2743,N_2661);
and U4963 (N_4963,N_2012,N_2479);
and U4964 (N_4964,N_3845,N_3925);
or U4965 (N_4965,N_2537,N_2702);
or U4966 (N_4966,N_2439,N_2803);
xor U4967 (N_4967,N_3215,N_2774);
or U4968 (N_4968,N_3028,N_2370);
or U4969 (N_4969,N_3097,N_3373);
xor U4970 (N_4970,N_3070,N_3909);
nand U4971 (N_4971,N_3135,N_2753);
or U4972 (N_4972,N_3920,N_3914);
and U4973 (N_4973,N_3631,N_2813);
or U4974 (N_4974,N_3798,N_2652);
and U4975 (N_4975,N_3139,N_2067);
or U4976 (N_4976,N_2993,N_3781);
and U4977 (N_4977,N_2523,N_3687);
xor U4978 (N_4978,N_3771,N_2833);
nor U4979 (N_4979,N_2149,N_2375);
xor U4980 (N_4980,N_3578,N_3057);
nand U4981 (N_4981,N_2647,N_2750);
and U4982 (N_4982,N_3840,N_2543);
nand U4983 (N_4983,N_3148,N_3301);
nand U4984 (N_4984,N_3265,N_2104);
nand U4985 (N_4985,N_3465,N_3189);
nand U4986 (N_4986,N_2075,N_3334);
nand U4987 (N_4987,N_2440,N_3065);
or U4988 (N_4988,N_2393,N_3790);
nand U4989 (N_4989,N_3731,N_2603);
nand U4990 (N_4990,N_2050,N_2052);
or U4991 (N_4991,N_3018,N_2975);
xor U4992 (N_4992,N_3196,N_2163);
xor U4993 (N_4993,N_3219,N_3295);
and U4994 (N_4994,N_2245,N_2222);
nand U4995 (N_4995,N_3862,N_2151);
nand U4996 (N_4996,N_3639,N_3563);
nand U4997 (N_4997,N_3742,N_2771);
and U4998 (N_4998,N_2171,N_2589);
nor U4999 (N_4999,N_3908,N_3564);
nand U5000 (N_5000,N_2713,N_3662);
nand U5001 (N_5001,N_3775,N_2726);
or U5002 (N_5002,N_3614,N_3640);
nand U5003 (N_5003,N_2016,N_3669);
nor U5004 (N_5004,N_3219,N_3667);
or U5005 (N_5005,N_2679,N_2582);
nand U5006 (N_5006,N_3714,N_3583);
nand U5007 (N_5007,N_3057,N_2144);
or U5008 (N_5008,N_2437,N_2102);
xnor U5009 (N_5009,N_2380,N_3307);
nand U5010 (N_5010,N_3262,N_3104);
and U5011 (N_5011,N_2920,N_3697);
nor U5012 (N_5012,N_3027,N_3421);
or U5013 (N_5013,N_3808,N_3193);
and U5014 (N_5014,N_2467,N_2972);
nor U5015 (N_5015,N_2519,N_3601);
or U5016 (N_5016,N_2693,N_2191);
and U5017 (N_5017,N_2969,N_3978);
or U5018 (N_5018,N_2348,N_2812);
xor U5019 (N_5019,N_3896,N_3692);
nor U5020 (N_5020,N_3441,N_3606);
and U5021 (N_5021,N_2809,N_3196);
xor U5022 (N_5022,N_3461,N_2513);
xnor U5023 (N_5023,N_3573,N_2167);
or U5024 (N_5024,N_2878,N_2298);
and U5025 (N_5025,N_2715,N_2895);
nand U5026 (N_5026,N_2563,N_2681);
xor U5027 (N_5027,N_3004,N_3946);
or U5028 (N_5028,N_2622,N_2496);
xor U5029 (N_5029,N_3904,N_2355);
xor U5030 (N_5030,N_3383,N_2709);
nand U5031 (N_5031,N_2900,N_2386);
or U5032 (N_5032,N_3802,N_3715);
nor U5033 (N_5033,N_2798,N_3082);
or U5034 (N_5034,N_2127,N_3031);
nor U5035 (N_5035,N_3364,N_2247);
and U5036 (N_5036,N_3914,N_3813);
nand U5037 (N_5037,N_3876,N_3451);
and U5038 (N_5038,N_2387,N_3997);
nand U5039 (N_5039,N_3109,N_3627);
and U5040 (N_5040,N_3751,N_2985);
nor U5041 (N_5041,N_2027,N_2232);
and U5042 (N_5042,N_3431,N_2172);
xor U5043 (N_5043,N_3558,N_2505);
xnor U5044 (N_5044,N_3060,N_3338);
and U5045 (N_5045,N_2750,N_2926);
and U5046 (N_5046,N_2523,N_3326);
and U5047 (N_5047,N_2036,N_2388);
nand U5048 (N_5048,N_2008,N_2608);
nor U5049 (N_5049,N_3992,N_3068);
nor U5050 (N_5050,N_3580,N_2605);
or U5051 (N_5051,N_2387,N_2025);
or U5052 (N_5052,N_3810,N_2621);
or U5053 (N_5053,N_2674,N_3427);
nand U5054 (N_5054,N_3384,N_2702);
or U5055 (N_5055,N_3007,N_3989);
xor U5056 (N_5056,N_2531,N_3665);
or U5057 (N_5057,N_2431,N_2142);
xor U5058 (N_5058,N_2358,N_3354);
xnor U5059 (N_5059,N_3913,N_3416);
and U5060 (N_5060,N_2095,N_2836);
xor U5061 (N_5061,N_3818,N_2018);
or U5062 (N_5062,N_3685,N_2701);
nor U5063 (N_5063,N_3649,N_3949);
nand U5064 (N_5064,N_2135,N_2469);
nand U5065 (N_5065,N_3355,N_3914);
or U5066 (N_5066,N_3861,N_3083);
xor U5067 (N_5067,N_2377,N_3457);
nand U5068 (N_5068,N_3839,N_3421);
or U5069 (N_5069,N_3305,N_2278);
or U5070 (N_5070,N_3079,N_3262);
or U5071 (N_5071,N_3384,N_2072);
or U5072 (N_5072,N_2329,N_2091);
xor U5073 (N_5073,N_2534,N_2505);
xnor U5074 (N_5074,N_2514,N_3636);
xor U5075 (N_5075,N_2480,N_3485);
nand U5076 (N_5076,N_3990,N_2022);
or U5077 (N_5077,N_2113,N_2299);
and U5078 (N_5078,N_3893,N_3991);
or U5079 (N_5079,N_2376,N_2836);
nand U5080 (N_5080,N_2378,N_3720);
nor U5081 (N_5081,N_2810,N_3923);
xnor U5082 (N_5082,N_3429,N_3166);
and U5083 (N_5083,N_2679,N_2154);
or U5084 (N_5084,N_3368,N_3271);
nand U5085 (N_5085,N_3115,N_3064);
or U5086 (N_5086,N_3455,N_3630);
nor U5087 (N_5087,N_3115,N_3629);
xor U5088 (N_5088,N_3100,N_3890);
xnor U5089 (N_5089,N_2839,N_2267);
nand U5090 (N_5090,N_3523,N_3451);
and U5091 (N_5091,N_2257,N_2055);
nand U5092 (N_5092,N_2657,N_2282);
xor U5093 (N_5093,N_2658,N_3361);
xnor U5094 (N_5094,N_3084,N_3481);
nor U5095 (N_5095,N_3322,N_2655);
xnor U5096 (N_5096,N_3583,N_3260);
and U5097 (N_5097,N_2473,N_2402);
or U5098 (N_5098,N_2593,N_2124);
xor U5099 (N_5099,N_3810,N_2416);
and U5100 (N_5100,N_3018,N_2334);
and U5101 (N_5101,N_2325,N_2586);
and U5102 (N_5102,N_3064,N_2260);
or U5103 (N_5103,N_2859,N_3798);
nor U5104 (N_5104,N_2800,N_3444);
or U5105 (N_5105,N_2530,N_2898);
nor U5106 (N_5106,N_3563,N_3379);
xor U5107 (N_5107,N_2926,N_3465);
or U5108 (N_5108,N_2321,N_3944);
nor U5109 (N_5109,N_2205,N_2858);
nand U5110 (N_5110,N_2620,N_3183);
nand U5111 (N_5111,N_3413,N_2766);
nand U5112 (N_5112,N_3612,N_2289);
nand U5113 (N_5113,N_2574,N_2382);
or U5114 (N_5114,N_2371,N_2380);
and U5115 (N_5115,N_2394,N_3411);
or U5116 (N_5116,N_3449,N_3598);
and U5117 (N_5117,N_2300,N_3593);
or U5118 (N_5118,N_2753,N_2367);
or U5119 (N_5119,N_3350,N_3028);
nand U5120 (N_5120,N_3034,N_3162);
or U5121 (N_5121,N_3991,N_3268);
nor U5122 (N_5122,N_2181,N_3191);
or U5123 (N_5123,N_3854,N_2084);
and U5124 (N_5124,N_3567,N_3886);
xnor U5125 (N_5125,N_3986,N_3944);
nand U5126 (N_5126,N_2259,N_3280);
xnor U5127 (N_5127,N_3393,N_2468);
nor U5128 (N_5128,N_3555,N_2279);
xnor U5129 (N_5129,N_3005,N_3040);
nor U5130 (N_5130,N_2594,N_2376);
or U5131 (N_5131,N_2842,N_2135);
or U5132 (N_5132,N_3834,N_2130);
or U5133 (N_5133,N_3473,N_2698);
nand U5134 (N_5134,N_2349,N_3793);
nor U5135 (N_5135,N_2188,N_3284);
nand U5136 (N_5136,N_3379,N_3303);
nor U5137 (N_5137,N_3809,N_2311);
and U5138 (N_5138,N_3889,N_3623);
and U5139 (N_5139,N_2213,N_3185);
nand U5140 (N_5140,N_2812,N_2845);
nand U5141 (N_5141,N_2830,N_3227);
nand U5142 (N_5142,N_3292,N_2569);
nor U5143 (N_5143,N_2270,N_3442);
nor U5144 (N_5144,N_3844,N_3265);
nand U5145 (N_5145,N_2789,N_3021);
xor U5146 (N_5146,N_3642,N_3831);
nand U5147 (N_5147,N_3300,N_2476);
xnor U5148 (N_5148,N_2627,N_3864);
or U5149 (N_5149,N_3091,N_2855);
or U5150 (N_5150,N_2443,N_2877);
nor U5151 (N_5151,N_3944,N_2464);
xnor U5152 (N_5152,N_3597,N_3327);
xor U5153 (N_5153,N_3886,N_2607);
nand U5154 (N_5154,N_2876,N_3411);
and U5155 (N_5155,N_2089,N_2445);
nor U5156 (N_5156,N_3098,N_2027);
nor U5157 (N_5157,N_2906,N_2770);
nand U5158 (N_5158,N_2467,N_2077);
xnor U5159 (N_5159,N_2680,N_3722);
nand U5160 (N_5160,N_3851,N_2907);
or U5161 (N_5161,N_2947,N_3034);
xor U5162 (N_5162,N_3981,N_3143);
xor U5163 (N_5163,N_3714,N_3197);
xor U5164 (N_5164,N_2332,N_2096);
and U5165 (N_5165,N_2620,N_3626);
or U5166 (N_5166,N_2539,N_2671);
or U5167 (N_5167,N_2124,N_3259);
xnor U5168 (N_5168,N_3671,N_2212);
and U5169 (N_5169,N_2654,N_2932);
xor U5170 (N_5170,N_3879,N_3330);
nand U5171 (N_5171,N_3872,N_3147);
nor U5172 (N_5172,N_3205,N_2334);
or U5173 (N_5173,N_2958,N_2303);
xnor U5174 (N_5174,N_3817,N_2550);
or U5175 (N_5175,N_3190,N_3570);
and U5176 (N_5176,N_3242,N_3627);
xnor U5177 (N_5177,N_3471,N_3677);
and U5178 (N_5178,N_2821,N_2060);
nand U5179 (N_5179,N_2646,N_2719);
nor U5180 (N_5180,N_2132,N_2143);
or U5181 (N_5181,N_3389,N_2989);
or U5182 (N_5182,N_2587,N_2375);
nor U5183 (N_5183,N_3521,N_2689);
xnor U5184 (N_5184,N_2967,N_2529);
nand U5185 (N_5185,N_2895,N_2150);
xor U5186 (N_5186,N_2667,N_3996);
or U5187 (N_5187,N_2318,N_2678);
nand U5188 (N_5188,N_3654,N_2451);
nor U5189 (N_5189,N_2220,N_3152);
and U5190 (N_5190,N_3302,N_2723);
nor U5191 (N_5191,N_2548,N_2727);
nand U5192 (N_5192,N_2729,N_2368);
nor U5193 (N_5193,N_3438,N_2192);
and U5194 (N_5194,N_2115,N_2075);
or U5195 (N_5195,N_3843,N_3141);
xnor U5196 (N_5196,N_2543,N_2148);
and U5197 (N_5197,N_3377,N_2584);
or U5198 (N_5198,N_2022,N_2766);
and U5199 (N_5199,N_2654,N_3252);
and U5200 (N_5200,N_3934,N_2312);
xor U5201 (N_5201,N_2096,N_3899);
nand U5202 (N_5202,N_3605,N_3457);
nand U5203 (N_5203,N_3512,N_2564);
xnor U5204 (N_5204,N_3388,N_3700);
nand U5205 (N_5205,N_3873,N_3850);
and U5206 (N_5206,N_2062,N_2552);
nand U5207 (N_5207,N_3091,N_3747);
or U5208 (N_5208,N_2015,N_2470);
nor U5209 (N_5209,N_3739,N_3798);
xor U5210 (N_5210,N_2001,N_2047);
xor U5211 (N_5211,N_2114,N_2762);
xnor U5212 (N_5212,N_2499,N_3139);
xnor U5213 (N_5213,N_3395,N_2742);
and U5214 (N_5214,N_3396,N_3491);
and U5215 (N_5215,N_3211,N_3318);
xor U5216 (N_5216,N_2642,N_2880);
nor U5217 (N_5217,N_3435,N_2124);
nor U5218 (N_5218,N_3795,N_2267);
or U5219 (N_5219,N_2213,N_3126);
nor U5220 (N_5220,N_3412,N_3692);
nand U5221 (N_5221,N_3957,N_2292);
or U5222 (N_5222,N_2082,N_3136);
xor U5223 (N_5223,N_3214,N_2697);
nand U5224 (N_5224,N_3578,N_3899);
nand U5225 (N_5225,N_2185,N_3445);
or U5226 (N_5226,N_2107,N_2258);
xnor U5227 (N_5227,N_3380,N_3920);
nor U5228 (N_5228,N_2866,N_3417);
nand U5229 (N_5229,N_2111,N_3018);
and U5230 (N_5230,N_2323,N_2130);
nand U5231 (N_5231,N_2295,N_2150);
nand U5232 (N_5232,N_3175,N_2735);
and U5233 (N_5233,N_2035,N_2878);
nand U5234 (N_5234,N_3741,N_3015);
nand U5235 (N_5235,N_2439,N_3608);
nand U5236 (N_5236,N_2744,N_3841);
and U5237 (N_5237,N_2016,N_2646);
nand U5238 (N_5238,N_2356,N_3424);
xor U5239 (N_5239,N_2059,N_3851);
xnor U5240 (N_5240,N_3826,N_2912);
nand U5241 (N_5241,N_3711,N_2811);
nor U5242 (N_5242,N_2989,N_2167);
nand U5243 (N_5243,N_2875,N_2337);
or U5244 (N_5244,N_2885,N_2348);
nand U5245 (N_5245,N_3603,N_2263);
nand U5246 (N_5246,N_3151,N_2067);
nor U5247 (N_5247,N_2942,N_2174);
nand U5248 (N_5248,N_2520,N_2085);
or U5249 (N_5249,N_3553,N_2817);
nand U5250 (N_5250,N_2319,N_3947);
or U5251 (N_5251,N_3893,N_2770);
and U5252 (N_5252,N_2246,N_3884);
nand U5253 (N_5253,N_3815,N_3999);
xor U5254 (N_5254,N_3585,N_2606);
and U5255 (N_5255,N_2682,N_2651);
xnor U5256 (N_5256,N_2412,N_3135);
and U5257 (N_5257,N_2422,N_3360);
xor U5258 (N_5258,N_3622,N_2064);
nor U5259 (N_5259,N_2839,N_2050);
nand U5260 (N_5260,N_3605,N_2724);
nor U5261 (N_5261,N_3812,N_2300);
and U5262 (N_5262,N_2830,N_3744);
nor U5263 (N_5263,N_3516,N_2734);
nand U5264 (N_5264,N_2475,N_3659);
or U5265 (N_5265,N_2989,N_3577);
and U5266 (N_5266,N_2223,N_3582);
and U5267 (N_5267,N_3606,N_3108);
and U5268 (N_5268,N_2692,N_2836);
nor U5269 (N_5269,N_3682,N_2977);
nor U5270 (N_5270,N_3711,N_2936);
xnor U5271 (N_5271,N_3648,N_3932);
and U5272 (N_5272,N_3053,N_3155);
nor U5273 (N_5273,N_3022,N_3087);
nor U5274 (N_5274,N_2033,N_2494);
nor U5275 (N_5275,N_2816,N_3559);
and U5276 (N_5276,N_2132,N_2269);
nand U5277 (N_5277,N_2237,N_2602);
and U5278 (N_5278,N_2118,N_2482);
nor U5279 (N_5279,N_3924,N_2814);
or U5280 (N_5280,N_3584,N_3153);
xor U5281 (N_5281,N_2301,N_2908);
or U5282 (N_5282,N_2724,N_3130);
and U5283 (N_5283,N_3667,N_2035);
nor U5284 (N_5284,N_2765,N_3055);
xnor U5285 (N_5285,N_2538,N_2979);
xor U5286 (N_5286,N_3681,N_3778);
or U5287 (N_5287,N_3188,N_3793);
xnor U5288 (N_5288,N_3528,N_3660);
nor U5289 (N_5289,N_2066,N_3156);
nand U5290 (N_5290,N_3819,N_2284);
nor U5291 (N_5291,N_2671,N_3400);
nand U5292 (N_5292,N_2853,N_2619);
and U5293 (N_5293,N_3615,N_2315);
nor U5294 (N_5294,N_2045,N_3353);
nand U5295 (N_5295,N_2328,N_2791);
and U5296 (N_5296,N_2672,N_2673);
xor U5297 (N_5297,N_2897,N_2780);
nor U5298 (N_5298,N_3008,N_3946);
and U5299 (N_5299,N_2461,N_2852);
or U5300 (N_5300,N_3661,N_3658);
and U5301 (N_5301,N_2074,N_2381);
nand U5302 (N_5302,N_3297,N_3458);
nand U5303 (N_5303,N_2958,N_3292);
or U5304 (N_5304,N_2654,N_3311);
nor U5305 (N_5305,N_3885,N_2679);
nand U5306 (N_5306,N_3308,N_2006);
xnor U5307 (N_5307,N_3826,N_3226);
nand U5308 (N_5308,N_2669,N_2793);
nor U5309 (N_5309,N_2459,N_3188);
xnor U5310 (N_5310,N_2381,N_2000);
or U5311 (N_5311,N_2071,N_2103);
xor U5312 (N_5312,N_3920,N_3404);
nand U5313 (N_5313,N_3212,N_2916);
or U5314 (N_5314,N_3429,N_3675);
nand U5315 (N_5315,N_2318,N_2238);
nand U5316 (N_5316,N_3757,N_2169);
nand U5317 (N_5317,N_2300,N_2718);
nand U5318 (N_5318,N_2667,N_3760);
xor U5319 (N_5319,N_3090,N_2082);
xnor U5320 (N_5320,N_3577,N_3334);
nand U5321 (N_5321,N_3868,N_3851);
nand U5322 (N_5322,N_2780,N_3183);
xnor U5323 (N_5323,N_3317,N_3861);
and U5324 (N_5324,N_2875,N_3236);
nor U5325 (N_5325,N_3899,N_2471);
or U5326 (N_5326,N_3452,N_3210);
nand U5327 (N_5327,N_3968,N_3532);
and U5328 (N_5328,N_3422,N_3754);
and U5329 (N_5329,N_2841,N_2396);
nand U5330 (N_5330,N_3925,N_2312);
or U5331 (N_5331,N_3018,N_3525);
nand U5332 (N_5332,N_3908,N_2243);
xor U5333 (N_5333,N_3644,N_2106);
xor U5334 (N_5334,N_3104,N_3647);
and U5335 (N_5335,N_3456,N_3597);
nand U5336 (N_5336,N_2584,N_3865);
or U5337 (N_5337,N_2219,N_3617);
or U5338 (N_5338,N_3986,N_2114);
or U5339 (N_5339,N_3469,N_3474);
xnor U5340 (N_5340,N_3605,N_2543);
nand U5341 (N_5341,N_3436,N_2778);
xor U5342 (N_5342,N_3352,N_3464);
xor U5343 (N_5343,N_3316,N_2500);
xor U5344 (N_5344,N_3429,N_3505);
nand U5345 (N_5345,N_3234,N_2580);
nor U5346 (N_5346,N_2246,N_3929);
and U5347 (N_5347,N_3850,N_2629);
nor U5348 (N_5348,N_3384,N_3495);
and U5349 (N_5349,N_3785,N_2136);
nor U5350 (N_5350,N_3587,N_2107);
nand U5351 (N_5351,N_3629,N_3931);
nor U5352 (N_5352,N_2229,N_2314);
nor U5353 (N_5353,N_2961,N_3378);
nand U5354 (N_5354,N_2301,N_3115);
or U5355 (N_5355,N_2173,N_3741);
and U5356 (N_5356,N_2653,N_2048);
xnor U5357 (N_5357,N_3671,N_2051);
nand U5358 (N_5358,N_2746,N_3113);
or U5359 (N_5359,N_2429,N_3731);
xor U5360 (N_5360,N_3252,N_3517);
nor U5361 (N_5361,N_3198,N_3200);
xor U5362 (N_5362,N_2301,N_2150);
or U5363 (N_5363,N_2698,N_2819);
and U5364 (N_5364,N_3025,N_2479);
and U5365 (N_5365,N_3339,N_3978);
nor U5366 (N_5366,N_3697,N_3934);
or U5367 (N_5367,N_2073,N_2595);
and U5368 (N_5368,N_3414,N_2726);
and U5369 (N_5369,N_3905,N_2981);
and U5370 (N_5370,N_3196,N_2101);
xnor U5371 (N_5371,N_2797,N_2423);
and U5372 (N_5372,N_2978,N_2660);
nand U5373 (N_5373,N_2039,N_2441);
nand U5374 (N_5374,N_2978,N_3430);
nand U5375 (N_5375,N_3129,N_2585);
nand U5376 (N_5376,N_2833,N_3898);
nor U5377 (N_5377,N_2267,N_3733);
nand U5378 (N_5378,N_2494,N_2565);
nand U5379 (N_5379,N_3294,N_3543);
nand U5380 (N_5380,N_3627,N_3417);
or U5381 (N_5381,N_2751,N_3506);
nand U5382 (N_5382,N_2721,N_3589);
nor U5383 (N_5383,N_2563,N_2510);
nand U5384 (N_5384,N_3943,N_3304);
xor U5385 (N_5385,N_2041,N_2126);
or U5386 (N_5386,N_3397,N_2699);
nand U5387 (N_5387,N_2424,N_2003);
and U5388 (N_5388,N_2580,N_3696);
nand U5389 (N_5389,N_2359,N_2005);
nor U5390 (N_5390,N_3809,N_2477);
and U5391 (N_5391,N_2851,N_2025);
nor U5392 (N_5392,N_2933,N_2924);
or U5393 (N_5393,N_2933,N_3001);
nor U5394 (N_5394,N_3507,N_2913);
and U5395 (N_5395,N_2806,N_3598);
xor U5396 (N_5396,N_2403,N_2472);
nor U5397 (N_5397,N_2024,N_3433);
xor U5398 (N_5398,N_2294,N_3100);
or U5399 (N_5399,N_2320,N_3796);
nand U5400 (N_5400,N_2955,N_3973);
and U5401 (N_5401,N_3955,N_2445);
or U5402 (N_5402,N_3219,N_2184);
nor U5403 (N_5403,N_2887,N_2285);
and U5404 (N_5404,N_2928,N_2253);
or U5405 (N_5405,N_3247,N_3325);
xnor U5406 (N_5406,N_2087,N_2016);
and U5407 (N_5407,N_3683,N_3720);
and U5408 (N_5408,N_2963,N_2971);
and U5409 (N_5409,N_2991,N_3152);
nand U5410 (N_5410,N_3513,N_2338);
xor U5411 (N_5411,N_2461,N_2880);
or U5412 (N_5412,N_3715,N_3353);
nor U5413 (N_5413,N_2263,N_3733);
nor U5414 (N_5414,N_2047,N_2077);
or U5415 (N_5415,N_2061,N_2532);
nand U5416 (N_5416,N_3997,N_2671);
nor U5417 (N_5417,N_2137,N_3030);
and U5418 (N_5418,N_3769,N_2090);
nand U5419 (N_5419,N_2225,N_3078);
nand U5420 (N_5420,N_3412,N_2967);
nand U5421 (N_5421,N_2154,N_2702);
nand U5422 (N_5422,N_2143,N_3191);
or U5423 (N_5423,N_2559,N_2713);
and U5424 (N_5424,N_3776,N_2265);
nor U5425 (N_5425,N_3070,N_3081);
and U5426 (N_5426,N_3819,N_3113);
nor U5427 (N_5427,N_3374,N_2250);
xor U5428 (N_5428,N_3153,N_2441);
xor U5429 (N_5429,N_2318,N_2803);
or U5430 (N_5430,N_2570,N_3803);
and U5431 (N_5431,N_2179,N_2555);
nor U5432 (N_5432,N_2351,N_3772);
xor U5433 (N_5433,N_3715,N_2222);
nand U5434 (N_5434,N_2944,N_3862);
nor U5435 (N_5435,N_3333,N_2818);
xnor U5436 (N_5436,N_2837,N_2042);
nor U5437 (N_5437,N_3430,N_2433);
or U5438 (N_5438,N_3439,N_2640);
and U5439 (N_5439,N_3486,N_3931);
nand U5440 (N_5440,N_3536,N_2836);
and U5441 (N_5441,N_2067,N_3575);
xor U5442 (N_5442,N_2758,N_3787);
nand U5443 (N_5443,N_2297,N_2688);
or U5444 (N_5444,N_3771,N_3359);
and U5445 (N_5445,N_2443,N_3076);
xor U5446 (N_5446,N_2474,N_3773);
nand U5447 (N_5447,N_2796,N_3252);
nand U5448 (N_5448,N_3359,N_2375);
xor U5449 (N_5449,N_2857,N_3254);
or U5450 (N_5450,N_3996,N_3672);
xor U5451 (N_5451,N_3950,N_2880);
and U5452 (N_5452,N_2262,N_2960);
nor U5453 (N_5453,N_2966,N_3264);
and U5454 (N_5454,N_2285,N_2358);
or U5455 (N_5455,N_3283,N_3938);
xnor U5456 (N_5456,N_2041,N_3416);
nand U5457 (N_5457,N_3179,N_3672);
nor U5458 (N_5458,N_2114,N_3555);
and U5459 (N_5459,N_2162,N_3917);
or U5460 (N_5460,N_2990,N_3006);
nor U5461 (N_5461,N_2059,N_2022);
xor U5462 (N_5462,N_2325,N_3603);
or U5463 (N_5463,N_2027,N_2441);
nor U5464 (N_5464,N_2258,N_3734);
and U5465 (N_5465,N_2009,N_3367);
nand U5466 (N_5466,N_2441,N_2164);
xor U5467 (N_5467,N_2637,N_2229);
and U5468 (N_5468,N_3190,N_2126);
and U5469 (N_5469,N_3804,N_2859);
and U5470 (N_5470,N_2930,N_2928);
nor U5471 (N_5471,N_3886,N_3961);
xor U5472 (N_5472,N_3320,N_2196);
or U5473 (N_5473,N_3365,N_3670);
and U5474 (N_5474,N_3705,N_3185);
nand U5475 (N_5475,N_2559,N_2102);
xnor U5476 (N_5476,N_3732,N_3459);
and U5477 (N_5477,N_2854,N_3360);
nor U5478 (N_5478,N_3656,N_3228);
nand U5479 (N_5479,N_3600,N_3049);
or U5480 (N_5480,N_2320,N_3005);
and U5481 (N_5481,N_3046,N_2553);
xnor U5482 (N_5482,N_2182,N_2229);
nor U5483 (N_5483,N_3165,N_2350);
nand U5484 (N_5484,N_2642,N_3698);
or U5485 (N_5485,N_3238,N_2778);
and U5486 (N_5486,N_2302,N_3317);
or U5487 (N_5487,N_2505,N_2965);
nand U5488 (N_5488,N_3509,N_3422);
and U5489 (N_5489,N_3281,N_2762);
and U5490 (N_5490,N_3575,N_3109);
nor U5491 (N_5491,N_2443,N_2983);
nand U5492 (N_5492,N_3596,N_2781);
or U5493 (N_5493,N_2317,N_2716);
or U5494 (N_5494,N_2778,N_2307);
xor U5495 (N_5495,N_2904,N_3472);
xor U5496 (N_5496,N_2858,N_2046);
or U5497 (N_5497,N_2097,N_3254);
xor U5498 (N_5498,N_2978,N_2416);
nand U5499 (N_5499,N_3104,N_2800);
or U5500 (N_5500,N_2782,N_2668);
nand U5501 (N_5501,N_2591,N_2460);
or U5502 (N_5502,N_3338,N_3531);
and U5503 (N_5503,N_2307,N_3955);
nor U5504 (N_5504,N_3147,N_2647);
nand U5505 (N_5505,N_3605,N_2455);
nor U5506 (N_5506,N_2411,N_3449);
nor U5507 (N_5507,N_2348,N_3338);
xor U5508 (N_5508,N_3975,N_3211);
or U5509 (N_5509,N_3406,N_3157);
nand U5510 (N_5510,N_2232,N_3565);
nand U5511 (N_5511,N_3793,N_2135);
and U5512 (N_5512,N_2394,N_3265);
nor U5513 (N_5513,N_2836,N_3604);
nand U5514 (N_5514,N_3374,N_3451);
or U5515 (N_5515,N_3473,N_3204);
or U5516 (N_5516,N_3767,N_2791);
nor U5517 (N_5517,N_3665,N_2242);
nor U5518 (N_5518,N_2509,N_3266);
or U5519 (N_5519,N_3164,N_3573);
and U5520 (N_5520,N_3729,N_2905);
xor U5521 (N_5521,N_2496,N_3348);
or U5522 (N_5522,N_3393,N_3921);
and U5523 (N_5523,N_2872,N_3266);
nor U5524 (N_5524,N_2512,N_2537);
xnor U5525 (N_5525,N_2706,N_2401);
nand U5526 (N_5526,N_2166,N_2946);
or U5527 (N_5527,N_3706,N_2750);
and U5528 (N_5528,N_3781,N_2633);
nand U5529 (N_5529,N_2075,N_3926);
nand U5530 (N_5530,N_2260,N_2826);
nand U5531 (N_5531,N_3924,N_2747);
or U5532 (N_5532,N_2346,N_3445);
xnor U5533 (N_5533,N_2510,N_3726);
or U5534 (N_5534,N_3146,N_2225);
xor U5535 (N_5535,N_2698,N_3177);
xor U5536 (N_5536,N_2180,N_3168);
or U5537 (N_5537,N_2698,N_2028);
xnor U5538 (N_5538,N_3212,N_3898);
xor U5539 (N_5539,N_3658,N_3964);
nor U5540 (N_5540,N_2243,N_3966);
xnor U5541 (N_5541,N_3624,N_2725);
and U5542 (N_5542,N_3419,N_3474);
or U5543 (N_5543,N_3013,N_3058);
xor U5544 (N_5544,N_3500,N_2509);
nand U5545 (N_5545,N_3509,N_2593);
or U5546 (N_5546,N_3854,N_3921);
and U5547 (N_5547,N_2433,N_3209);
or U5548 (N_5548,N_3049,N_2741);
nand U5549 (N_5549,N_2211,N_3308);
xor U5550 (N_5550,N_3919,N_3228);
xor U5551 (N_5551,N_2789,N_2166);
and U5552 (N_5552,N_3599,N_2462);
nor U5553 (N_5553,N_2982,N_3005);
nor U5554 (N_5554,N_3383,N_3649);
and U5555 (N_5555,N_3755,N_2721);
xor U5556 (N_5556,N_2540,N_2750);
nor U5557 (N_5557,N_2623,N_3212);
nor U5558 (N_5558,N_3196,N_2808);
and U5559 (N_5559,N_3984,N_3789);
or U5560 (N_5560,N_3117,N_2382);
xor U5561 (N_5561,N_3692,N_2466);
and U5562 (N_5562,N_2086,N_2883);
and U5563 (N_5563,N_3297,N_2553);
and U5564 (N_5564,N_3575,N_3876);
nor U5565 (N_5565,N_3924,N_3546);
nand U5566 (N_5566,N_3546,N_3177);
and U5567 (N_5567,N_2493,N_3560);
xnor U5568 (N_5568,N_2312,N_2494);
and U5569 (N_5569,N_3558,N_3722);
and U5570 (N_5570,N_2449,N_2507);
nand U5571 (N_5571,N_2597,N_2366);
and U5572 (N_5572,N_3496,N_3156);
xor U5573 (N_5573,N_2003,N_3075);
nor U5574 (N_5574,N_3702,N_2537);
xor U5575 (N_5575,N_3360,N_3016);
nor U5576 (N_5576,N_3681,N_2948);
and U5577 (N_5577,N_3269,N_3818);
and U5578 (N_5578,N_2465,N_2997);
nor U5579 (N_5579,N_2099,N_2922);
xnor U5580 (N_5580,N_2882,N_2612);
nor U5581 (N_5581,N_2391,N_3275);
nor U5582 (N_5582,N_3135,N_2641);
nor U5583 (N_5583,N_2591,N_2043);
or U5584 (N_5584,N_2812,N_2911);
and U5585 (N_5585,N_2699,N_3538);
and U5586 (N_5586,N_2840,N_2162);
and U5587 (N_5587,N_3054,N_3931);
or U5588 (N_5588,N_3685,N_2179);
xor U5589 (N_5589,N_2247,N_2612);
nor U5590 (N_5590,N_2490,N_2900);
nor U5591 (N_5591,N_2314,N_3735);
or U5592 (N_5592,N_3124,N_3073);
nor U5593 (N_5593,N_2058,N_2369);
nand U5594 (N_5594,N_2527,N_3990);
xor U5595 (N_5595,N_2562,N_2915);
nand U5596 (N_5596,N_3764,N_2523);
xnor U5597 (N_5597,N_2627,N_2908);
xnor U5598 (N_5598,N_2890,N_3526);
and U5599 (N_5599,N_3495,N_2869);
nand U5600 (N_5600,N_2112,N_2404);
or U5601 (N_5601,N_3293,N_2209);
and U5602 (N_5602,N_2635,N_2453);
xnor U5603 (N_5603,N_3255,N_3888);
and U5604 (N_5604,N_2588,N_3065);
and U5605 (N_5605,N_3562,N_3728);
xnor U5606 (N_5606,N_2340,N_2959);
nor U5607 (N_5607,N_3974,N_2282);
nand U5608 (N_5608,N_2381,N_2517);
and U5609 (N_5609,N_2084,N_2472);
xnor U5610 (N_5610,N_2068,N_3744);
and U5611 (N_5611,N_3636,N_2371);
and U5612 (N_5612,N_3148,N_3025);
nor U5613 (N_5613,N_2698,N_3926);
nand U5614 (N_5614,N_3862,N_3322);
xor U5615 (N_5615,N_3186,N_3773);
nand U5616 (N_5616,N_3558,N_3970);
nor U5617 (N_5617,N_2038,N_2405);
nand U5618 (N_5618,N_3983,N_2225);
and U5619 (N_5619,N_2258,N_2311);
or U5620 (N_5620,N_3754,N_3472);
nand U5621 (N_5621,N_2473,N_3701);
xor U5622 (N_5622,N_2319,N_3345);
nor U5623 (N_5623,N_2175,N_3097);
xnor U5624 (N_5624,N_3964,N_2386);
and U5625 (N_5625,N_2661,N_2756);
nand U5626 (N_5626,N_2889,N_3899);
or U5627 (N_5627,N_3832,N_2291);
nor U5628 (N_5628,N_2842,N_3062);
xnor U5629 (N_5629,N_3243,N_3828);
and U5630 (N_5630,N_2452,N_2977);
or U5631 (N_5631,N_2225,N_2432);
nor U5632 (N_5632,N_2764,N_2518);
nand U5633 (N_5633,N_3179,N_2696);
and U5634 (N_5634,N_3162,N_3007);
or U5635 (N_5635,N_2603,N_3022);
or U5636 (N_5636,N_2564,N_2193);
or U5637 (N_5637,N_2740,N_3490);
nor U5638 (N_5638,N_2916,N_3589);
or U5639 (N_5639,N_2126,N_3387);
nand U5640 (N_5640,N_3554,N_3207);
and U5641 (N_5641,N_2699,N_3664);
nand U5642 (N_5642,N_2383,N_3286);
nor U5643 (N_5643,N_2517,N_2597);
nor U5644 (N_5644,N_3011,N_3376);
xnor U5645 (N_5645,N_3076,N_2118);
xor U5646 (N_5646,N_3029,N_3722);
nor U5647 (N_5647,N_2040,N_2863);
nand U5648 (N_5648,N_2731,N_3445);
or U5649 (N_5649,N_3007,N_2605);
nor U5650 (N_5650,N_3300,N_3903);
or U5651 (N_5651,N_2047,N_2985);
xor U5652 (N_5652,N_2972,N_2702);
or U5653 (N_5653,N_2024,N_3249);
nor U5654 (N_5654,N_3420,N_3345);
and U5655 (N_5655,N_2103,N_2036);
or U5656 (N_5656,N_3335,N_2255);
nor U5657 (N_5657,N_3670,N_2835);
xnor U5658 (N_5658,N_2510,N_3544);
nor U5659 (N_5659,N_3767,N_2951);
and U5660 (N_5660,N_2072,N_2468);
nor U5661 (N_5661,N_3032,N_2905);
nor U5662 (N_5662,N_3842,N_2630);
and U5663 (N_5663,N_3145,N_2925);
xnor U5664 (N_5664,N_3046,N_2456);
nand U5665 (N_5665,N_3068,N_3939);
or U5666 (N_5666,N_3943,N_2329);
nand U5667 (N_5667,N_2261,N_3209);
nor U5668 (N_5668,N_2204,N_2525);
xnor U5669 (N_5669,N_3241,N_3109);
and U5670 (N_5670,N_2390,N_3147);
xor U5671 (N_5671,N_2057,N_3693);
nor U5672 (N_5672,N_2042,N_3062);
nand U5673 (N_5673,N_3041,N_3096);
and U5674 (N_5674,N_2091,N_2539);
or U5675 (N_5675,N_3772,N_2947);
nor U5676 (N_5676,N_3271,N_3961);
nand U5677 (N_5677,N_2190,N_2701);
or U5678 (N_5678,N_2944,N_3271);
nor U5679 (N_5679,N_3121,N_2902);
nand U5680 (N_5680,N_3998,N_2548);
and U5681 (N_5681,N_3388,N_3923);
xor U5682 (N_5682,N_3798,N_2473);
xor U5683 (N_5683,N_3735,N_2712);
nand U5684 (N_5684,N_3360,N_2596);
nand U5685 (N_5685,N_3096,N_2868);
and U5686 (N_5686,N_2634,N_3389);
and U5687 (N_5687,N_2510,N_2947);
xor U5688 (N_5688,N_3431,N_3109);
and U5689 (N_5689,N_2195,N_3220);
nor U5690 (N_5690,N_2142,N_2250);
nor U5691 (N_5691,N_2806,N_2903);
nand U5692 (N_5692,N_3692,N_3968);
xor U5693 (N_5693,N_3914,N_3700);
nand U5694 (N_5694,N_3181,N_2423);
nand U5695 (N_5695,N_2267,N_2168);
xor U5696 (N_5696,N_2513,N_3826);
xor U5697 (N_5697,N_3421,N_3587);
or U5698 (N_5698,N_3433,N_2842);
and U5699 (N_5699,N_3190,N_2294);
or U5700 (N_5700,N_2578,N_3600);
nand U5701 (N_5701,N_2107,N_3446);
nor U5702 (N_5702,N_3205,N_3358);
nor U5703 (N_5703,N_2562,N_3192);
or U5704 (N_5704,N_2373,N_2670);
xnor U5705 (N_5705,N_2649,N_2377);
xor U5706 (N_5706,N_3707,N_3953);
and U5707 (N_5707,N_3489,N_3405);
nand U5708 (N_5708,N_3823,N_3822);
nand U5709 (N_5709,N_2459,N_3763);
xor U5710 (N_5710,N_2651,N_3882);
nand U5711 (N_5711,N_3552,N_3120);
nor U5712 (N_5712,N_2474,N_2008);
nor U5713 (N_5713,N_2877,N_3731);
xor U5714 (N_5714,N_3951,N_3826);
and U5715 (N_5715,N_2458,N_3381);
or U5716 (N_5716,N_3241,N_3776);
xnor U5717 (N_5717,N_2970,N_3060);
nor U5718 (N_5718,N_2467,N_3083);
xnor U5719 (N_5719,N_2836,N_3357);
nand U5720 (N_5720,N_3534,N_3055);
nand U5721 (N_5721,N_3371,N_3961);
or U5722 (N_5722,N_3995,N_3087);
nand U5723 (N_5723,N_2009,N_3398);
or U5724 (N_5724,N_2256,N_3876);
nand U5725 (N_5725,N_3144,N_2091);
nand U5726 (N_5726,N_2020,N_2355);
nand U5727 (N_5727,N_3297,N_3702);
nor U5728 (N_5728,N_2715,N_3143);
nand U5729 (N_5729,N_2497,N_2603);
and U5730 (N_5730,N_2004,N_2736);
or U5731 (N_5731,N_3869,N_3665);
nand U5732 (N_5732,N_3088,N_2206);
xnor U5733 (N_5733,N_2559,N_2354);
nand U5734 (N_5734,N_3948,N_2090);
nand U5735 (N_5735,N_2728,N_2542);
or U5736 (N_5736,N_2273,N_2716);
nor U5737 (N_5737,N_2405,N_2981);
nor U5738 (N_5738,N_3085,N_2563);
xor U5739 (N_5739,N_2238,N_2608);
and U5740 (N_5740,N_2083,N_2946);
nand U5741 (N_5741,N_2778,N_2049);
xor U5742 (N_5742,N_3277,N_2703);
xor U5743 (N_5743,N_3570,N_2996);
or U5744 (N_5744,N_3413,N_2757);
xnor U5745 (N_5745,N_3440,N_2548);
xnor U5746 (N_5746,N_3038,N_2843);
nor U5747 (N_5747,N_3294,N_2910);
nand U5748 (N_5748,N_2531,N_3871);
and U5749 (N_5749,N_3931,N_3167);
and U5750 (N_5750,N_3127,N_3695);
or U5751 (N_5751,N_2927,N_3733);
xnor U5752 (N_5752,N_2307,N_3431);
and U5753 (N_5753,N_3932,N_3653);
nor U5754 (N_5754,N_2634,N_3457);
or U5755 (N_5755,N_3442,N_3551);
xnor U5756 (N_5756,N_3983,N_3464);
and U5757 (N_5757,N_2851,N_2621);
nand U5758 (N_5758,N_3458,N_2147);
nand U5759 (N_5759,N_2340,N_3274);
and U5760 (N_5760,N_2635,N_2508);
and U5761 (N_5761,N_2554,N_2434);
xnor U5762 (N_5762,N_3033,N_2653);
nand U5763 (N_5763,N_3834,N_3301);
or U5764 (N_5764,N_3928,N_2919);
or U5765 (N_5765,N_3442,N_2727);
nand U5766 (N_5766,N_3964,N_2393);
nor U5767 (N_5767,N_3442,N_2005);
and U5768 (N_5768,N_3580,N_3432);
nor U5769 (N_5769,N_3594,N_2871);
xor U5770 (N_5770,N_3075,N_2329);
nand U5771 (N_5771,N_2827,N_2363);
xnor U5772 (N_5772,N_3284,N_2368);
or U5773 (N_5773,N_2841,N_3918);
xnor U5774 (N_5774,N_3025,N_3838);
or U5775 (N_5775,N_3651,N_3890);
nor U5776 (N_5776,N_2783,N_2035);
nand U5777 (N_5777,N_3455,N_2771);
xnor U5778 (N_5778,N_2070,N_2534);
and U5779 (N_5779,N_3676,N_3159);
nor U5780 (N_5780,N_3185,N_3488);
nor U5781 (N_5781,N_2825,N_2264);
and U5782 (N_5782,N_2781,N_2391);
nor U5783 (N_5783,N_3497,N_3270);
or U5784 (N_5784,N_2367,N_3585);
nand U5785 (N_5785,N_2980,N_2326);
nand U5786 (N_5786,N_2725,N_3500);
or U5787 (N_5787,N_3037,N_2577);
and U5788 (N_5788,N_2833,N_3722);
nand U5789 (N_5789,N_2448,N_3788);
xor U5790 (N_5790,N_3164,N_3443);
and U5791 (N_5791,N_3068,N_3656);
or U5792 (N_5792,N_2240,N_3737);
nor U5793 (N_5793,N_3658,N_3023);
or U5794 (N_5794,N_3083,N_3932);
nand U5795 (N_5795,N_3296,N_3641);
or U5796 (N_5796,N_3841,N_3117);
and U5797 (N_5797,N_3107,N_2082);
or U5798 (N_5798,N_3951,N_2211);
nor U5799 (N_5799,N_3169,N_2893);
xor U5800 (N_5800,N_3553,N_2689);
xor U5801 (N_5801,N_3076,N_3083);
or U5802 (N_5802,N_2803,N_3555);
and U5803 (N_5803,N_3472,N_3047);
or U5804 (N_5804,N_3416,N_2236);
xnor U5805 (N_5805,N_2421,N_3527);
xor U5806 (N_5806,N_3979,N_3419);
and U5807 (N_5807,N_2779,N_2894);
or U5808 (N_5808,N_3788,N_2217);
and U5809 (N_5809,N_2427,N_3689);
nand U5810 (N_5810,N_3847,N_2353);
nor U5811 (N_5811,N_2487,N_2870);
nor U5812 (N_5812,N_2728,N_3561);
xor U5813 (N_5813,N_2959,N_3490);
nor U5814 (N_5814,N_3989,N_3021);
and U5815 (N_5815,N_3317,N_3040);
and U5816 (N_5816,N_3164,N_2172);
nor U5817 (N_5817,N_3315,N_2224);
xnor U5818 (N_5818,N_2882,N_2293);
or U5819 (N_5819,N_2450,N_3319);
xnor U5820 (N_5820,N_2181,N_3349);
xor U5821 (N_5821,N_2586,N_3678);
or U5822 (N_5822,N_3394,N_3259);
nand U5823 (N_5823,N_2792,N_2255);
and U5824 (N_5824,N_3214,N_2814);
nor U5825 (N_5825,N_2343,N_3331);
nand U5826 (N_5826,N_2399,N_2868);
nor U5827 (N_5827,N_2438,N_3123);
xnor U5828 (N_5828,N_2619,N_2248);
or U5829 (N_5829,N_3454,N_2857);
and U5830 (N_5830,N_3238,N_2142);
nand U5831 (N_5831,N_3494,N_3255);
and U5832 (N_5832,N_3211,N_2432);
nand U5833 (N_5833,N_2424,N_3397);
nor U5834 (N_5834,N_3895,N_2780);
or U5835 (N_5835,N_2205,N_3993);
or U5836 (N_5836,N_3174,N_2434);
or U5837 (N_5837,N_3514,N_2403);
and U5838 (N_5838,N_3211,N_2236);
xnor U5839 (N_5839,N_3320,N_3821);
xor U5840 (N_5840,N_2786,N_2200);
xnor U5841 (N_5841,N_3126,N_2234);
and U5842 (N_5842,N_2052,N_3063);
xnor U5843 (N_5843,N_2391,N_3874);
or U5844 (N_5844,N_3017,N_3954);
or U5845 (N_5845,N_3684,N_2638);
nor U5846 (N_5846,N_2592,N_3492);
nand U5847 (N_5847,N_3765,N_3915);
nor U5848 (N_5848,N_3946,N_3948);
and U5849 (N_5849,N_2174,N_3164);
nand U5850 (N_5850,N_2560,N_2535);
or U5851 (N_5851,N_2316,N_3031);
and U5852 (N_5852,N_2738,N_3316);
or U5853 (N_5853,N_2402,N_3363);
nor U5854 (N_5854,N_3184,N_2840);
nor U5855 (N_5855,N_3688,N_2174);
nor U5856 (N_5856,N_3263,N_3727);
xnor U5857 (N_5857,N_3136,N_2545);
nand U5858 (N_5858,N_3033,N_2899);
nand U5859 (N_5859,N_3443,N_3304);
xor U5860 (N_5860,N_2048,N_3692);
and U5861 (N_5861,N_3031,N_3912);
and U5862 (N_5862,N_3409,N_3185);
xnor U5863 (N_5863,N_2322,N_3752);
nand U5864 (N_5864,N_2963,N_3312);
and U5865 (N_5865,N_3826,N_3517);
nand U5866 (N_5866,N_2142,N_3473);
and U5867 (N_5867,N_2192,N_2798);
nor U5868 (N_5868,N_2690,N_2669);
and U5869 (N_5869,N_2305,N_3497);
or U5870 (N_5870,N_2627,N_3831);
and U5871 (N_5871,N_2277,N_2049);
xor U5872 (N_5872,N_3131,N_3402);
or U5873 (N_5873,N_2446,N_2054);
nor U5874 (N_5874,N_3452,N_2402);
and U5875 (N_5875,N_3143,N_2776);
and U5876 (N_5876,N_2131,N_2872);
or U5877 (N_5877,N_2064,N_2007);
and U5878 (N_5878,N_3053,N_2069);
nand U5879 (N_5879,N_3424,N_3419);
nor U5880 (N_5880,N_2135,N_2856);
xor U5881 (N_5881,N_3492,N_2714);
nand U5882 (N_5882,N_3683,N_2220);
nand U5883 (N_5883,N_3995,N_3229);
xor U5884 (N_5884,N_3965,N_3790);
nand U5885 (N_5885,N_3714,N_2282);
nand U5886 (N_5886,N_2132,N_3879);
nor U5887 (N_5887,N_3713,N_3277);
nor U5888 (N_5888,N_3718,N_3682);
nor U5889 (N_5889,N_2270,N_2885);
nand U5890 (N_5890,N_2522,N_3045);
nand U5891 (N_5891,N_2060,N_2196);
or U5892 (N_5892,N_3670,N_2162);
or U5893 (N_5893,N_3942,N_3313);
nand U5894 (N_5894,N_3049,N_2000);
xnor U5895 (N_5895,N_2884,N_2575);
and U5896 (N_5896,N_3149,N_3303);
nor U5897 (N_5897,N_2798,N_2028);
or U5898 (N_5898,N_3592,N_2714);
xor U5899 (N_5899,N_2290,N_2124);
xor U5900 (N_5900,N_2449,N_3869);
nor U5901 (N_5901,N_3872,N_3954);
nor U5902 (N_5902,N_3750,N_2860);
and U5903 (N_5903,N_2421,N_2533);
xor U5904 (N_5904,N_2442,N_3403);
xnor U5905 (N_5905,N_2805,N_3748);
nor U5906 (N_5906,N_2828,N_3456);
or U5907 (N_5907,N_3237,N_3765);
or U5908 (N_5908,N_2102,N_2302);
nand U5909 (N_5909,N_3498,N_3672);
nand U5910 (N_5910,N_2154,N_2426);
nand U5911 (N_5911,N_3620,N_3089);
or U5912 (N_5912,N_3196,N_3374);
and U5913 (N_5913,N_2304,N_3913);
nor U5914 (N_5914,N_2414,N_3414);
or U5915 (N_5915,N_2742,N_3393);
xnor U5916 (N_5916,N_2942,N_2810);
or U5917 (N_5917,N_2388,N_3805);
or U5918 (N_5918,N_2235,N_2120);
nand U5919 (N_5919,N_2285,N_3445);
nor U5920 (N_5920,N_3941,N_3705);
nor U5921 (N_5921,N_3705,N_3951);
or U5922 (N_5922,N_3432,N_2560);
nand U5923 (N_5923,N_3214,N_3004);
and U5924 (N_5924,N_3250,N_3682);
and U5925 (N_5925,N_2584,N_3745);
and U5926 (N_5926,N_3545,N_2010);
and U5927 (N_5927,N_2721,N_3800);
nor U5928 (N_5928,N_2612,N_3128);
nor U5929 (N_5929,N_3060,N_3878);
xnor U5930 (N_5930,N_2389,N_2231);
nor U5931 (N_5931,N_3096,N_3530);
or U5932 (N_5932,N_3484,N_3702);
and U5933 (N_5933,N_2097,N_2613);
xnor U5934 (N_5934,N_2532,N_2245);
and U5935 (N_5935,N_3673,N_2688);
or U5936 (N_5936,N_3904,N_3702);
nand U5937 (N_5937,N_3737,N_2942);
or U5938 (N_5938,N_2537,N_2700);
nor U5939 (N_5939,N_3473,N_3407);
xor U5940 (N_5940,N_2801,N_3967);
nand U5941 (N_5941,N_3410,N_2862);
and U5942 (N_5942,N_2934,N_2542);
nor U5943 (N_5943,N_2944,N_3072);
or U5944 (N_5944,N_2395,N_2382);
and U5945 (N_5945,N_3807,N_2475);
nor U5946 (N_5946,N_2195,N_2961);
xor U5947 (N_5947,N_2768,N_2822);
nand U5948 (N_5948,N_3939,N_3553);
nor U5949 (N_5949,N_2413,N_3727);
nor U5950 (N_5950,N_3361,N_2270);
and U5951 (N_5951,N_2865,N_2874);
and U5952 (N_5952,N_2423,N_3997);
and U5953 (N_5953,N_2913,N_2416);
nor U5954 (N_5954,N_2719,N_2105);
or U5955 (N_5955,N_3287,N_3310);
nand U5956 (N_5956,N_3597,N_2880);
nand U5957 (N_5957,N_3920,N_2756);
nand U5958 (N_5958,N_3283,N_2138);
nor U5959 (N_5959,N_2913,N_3219);
nand U5960 (N_5960,N_2531,N_3055);
nor U5961 (N_5961,N_3341,N_2104);
nor U5962 (N_5962,N_2742,N_2130);
or U5963 (N_5963,N_3211,N_3202);
nor U5964 (N_5964,N_2832,N_3339);
xor U5965 (N_5965,N_2246,N_3282);
and U5966 (N_5966,N_2725,N_3169);
or U5967 (N_5967,N_2576,N_3521);
and U5968 (N_5968,N_3904,N_3734);
xnor U5969 (N_5969,N_3971,N_2226);
nand U5970 (N_5970,N_3719,N_2201);
or U5971 (N_5971,N_3046,N_3932);
nor U5972 (N_5972,N_3352,N_3909);
nand U5973 (N_5973,N_2602,N_2730);
or U5974 (N_5974,N_3893,N_3279);
nor U5975 (N_5975,N_3089,N_2887);
xnor U5976 (N_5976,N_2035,N_2410);
nor U5977 (N_5977,N_2109,N_2908);
or U5978 (N_5978,N_2790,N_3111);
nand U5979 (N_5979,N_2165,N_2341);
and U5980 (N_5980,N_2139,N_3031);
or U5981 (N_5981,N_3748,N_2976);
and U5982 (N_5982,N_3374,N_3731);
or U5983 (N_5983,N_2037,N_2248);
xor U5984 (N_5984,N_2083,N_2823);
nor U5985 (N_5985,N_2230,N_2026);
nor U5986 (N_5986,N_2747,N_3498);
nand U5987 (N_5987,N_3660,N_2590);
and U5988 (N_5988,N_2632,N_3301);
nor U5989 (N_5989,N_2864,N_3190);
nand U5990 (N_5990,N_3261,N_3307);
xnor U5991 (N_5991,N_3578,N_2309);
nor U5992 (N_5992,N_2779,N_2155);
xnor U5993 (N_5993,N_3410,N_2254);
or U5994 (N_5994,N_2864,N_2583);
and U5995 (N_5995,N_2290,N_2224);
nor U5996 (N_5996,N_3372,N_3815);
nor U5997 (N_5997,N_2102,N_3692);
and U5998 (N_5998,N_3290,N_2825);
and U5999 (N_5999,N_2258,N_2613);
nor U6000 (N_6000,N_4241,N_5428);
xor U6001 (N_6001,N_5038,N_5738);
or U6002 (N_6002,N_4219,N_5133);
xnor U6003 (N_6003,N_5235,N_4511);
nor U6004 (N_6004,N_5983,N_4745);
nand U6005 (N_6005,N_4589,N_4918);
and U6006 (N_6006,N_4524,N_5850);
and U6007 (N_6007,N_5661,N_5331);
nand U6008 (N_6008,N_5993,N_5915);
xnor U6009 (N_6009,N_4698,N_5654);
nor U6010 (N_6010,N_4781,N_5572);
or U6011 (N_6011,N_5517,N_4240);
and U6012 (N_6012,N_5615,N_4766);
and U6013 (N_6013,N_5766,N_5744);
nor U6014 (N_6014,N_4016,N_5342);
nor U6015 (N_6015,N_4760,N_4383);
nor U6016 (N_6016,N_5505,N_4547);
xor U6017 (N_6017,N_5583,N_5734);
and U6018 (N_6018,N_5364,N_5971);
and U6019 (N_6019,N_4556,N_4818);
xor U6020 (N_6020,N_5590,N_4667);
nand U6021 (N_6021,N_5730,N_4031);
nand U6022 (N_6022,N_4289,N_4902);
nor U6023 (N_6023,N_4995,N_4183);
nor U6024 (N_6024,N_5226,N_4738);
and U6025 (N_6025,N_4139,N_4780);
xor U6026 (N_6026,N_5911,N_5834);
nor U6027 (N_6027,N_4883,N_5885);
and U6028 (N_6028,N_5122,N_4207);
nand U6029 (N_6029,N_4049,N_4854);
nand U6030 (N_6030,N_5644,N_5014);
xnor U6031 (N_6031,N_5456,N_5113);
nand U6032 (N_6032,N_5527,N_4328);
nand U6033 (N_6033,N_5145,N_5294);
xor U6034 (N_6034,N_5794,N_4969);
nand U6035 (N_6035,N_5731,N_5825);
nor U6036 (N_6036,N_5622,N_5204);
and U6037 (N_6037,N_4179,N_5628);
xor U6038 (N_6038,N_4200,N_4076);
nor U6039 (N_6039,N_5819,N_4649);
or U6040 (N_6040,N_5416,N_4164);
or U6041 (N_6041,N_5809,N_5727);
nand U6042 (N_6042,N_4157,N_4844);
or U6043 (N_6043,N_5714,N_5399);
or U6044 (N_6044,N_5659,N_4807);
xor U6045 (N_6045,N_4099,N_4478);
nor U6046 (N_6046,N_5676,N_4979);
and U6047 (N_6047,N_4506,N_5537);
nor U6048 (N_6048,N_4222,N_5435);
and U6049 (N_6049,N_5426,N_5212);
nor U6050 (N_6050,N_5323,N_4591);
xor U6051 (N_6051,N_5507,N_5540);
or U6052 (N_6052,N_5791,N_4269);
or U6053 (N_6053,N_5655,N_5251);
or U6054 (N_6054,N_5677,N_4334);
or U6055 (N_6055,N_5474,N_5196);
or U6056 (N_6056,N_5747,N_4897);
and U6057 (N_6057,N_4682,N_5601);
and U6058 (N_6058,N_4720,N_5824);
and U6059 (N_6059,N_4496,N_5402);
nor U6060 (N_6060,N_4586,N_4823);
and U6061 (N_6061,N_4508,N_5266);
nor U6062 (N_6062,N_4799,N_4683);
nand U6063 (N_6063,N_5568,N_5752);
and U6064 (N_6064,N_4041,N_5082);
nor U6065 (N_6065,N_5863,N_5599);
nor U6066 (N_6066,N_4210,N_4371);
xor U6067 (N_6067,N_5864,N_5951);
nor U6068 (N_6068,N_4488,N_5703);
or U6069 (N_6069,N_5961,N_4346);
or U6070 (N_6070,N_4726,N_4029);
and U6071 (N_6071,N_5783,N_4708);
and U6072 (N_6072,N_4609,N_4084);
or U6073 (N_6073,N_4652,N_5109);
and U6074 (N_6074,N_4864,N_5120);
and U6075 (N_6075,N_4093,N_5771);
xnor U6076 (N_6076,N_5292,N_4282);
and U6077 (N_6077,N_4774,N_4263);
or U6078 (N_6078,N_4359,N_4000);
nor U6079 (N_6079,N_4692,N_4115);
xnor U6080 (N_6080,N_4987,N_5062);
nand U6081 (N_6081,N_5952,N_5447);
and U6082 (N_6082,N_4209,N_5041);
and U6083 (N_6083,N_4929,N_5175);
nand U6084 (N_6084,N_4010,N_5262);
nor U6085 (N_6085,N_4418,N_5211);
or U6086 (N_6086,N_4160,N_4958);
nand U6087 (N_6087,N_4477,N_5822);
nand U6088 (N_6088,N_4162,N_4857);
nor U6089 (N_6089,N_4402,N_5312);
nand U6090 (N_6090,N_4023,N_4944);
nor U6091 (N_6091,N_5980,N_5999);
or U6092 (N_6092,N_4087,N_5471);
or U6093 (N_6093,N_5037,N_4009);
and U6094 (N_6094,N_5931,N_4483);
or U6095 (N_6095,N_4654,N_4975);
nand U6096 (N_6096,N_4391,N_5751);
and U6097 (N_6097,N_4980,N_4133);
or U6098 (N_6098,N_4364,N_5076);
xnor U6099 (N_6099,N_5238,N_4149);
xnor U6100 (N_6100,N_5541,N_4841);
nor U6101 (N_6101,N_5743,N_5179);
nand U6102 (N_6102,N_4990,N_5502);
nand U6103 (N_6103,N_4577,N_5278);
xor U6104 (N_6104,N_4830,N_4134);
xor U6105 (N_6105,N_5019,N_5116);
xnor U6106 (N_6106,N_4666,N_4624);
xnor U6107 (N_6107,N_4361,N_5310);
xor U6108 (N_6108,N_5207,N_5051);
and U6109 (N_6109,N_5995,N_5012);
nor U6110 (N_6110,N_4890,N_4660);
nand U6111 (N_6111,N_4629,N_4323);
or U6112 (N_6112,N_5722,N_5536);
nand U6113 (N_6113,N_5682,N_5988);
or U6114 (N_6114,N_4188,N_4317);
nor U6115 (N_6115,N_4723,N_4761);
xnor U6116 (N_6116,N_5754,N_4332);
nor U6117 (N_6117,N_5023,N_5647);
nand U6118 (N_6118,N_4439,N_5313);
nor U6119 (N_6119,N_5699,N_4779);
nor U6120 (N_6120,N_4366,N_4693);
nand U6121 (N_6121,N_5296,N_5847);
xor U6122 (N_6122,N_5845,N_4204);
nor U6123 (N_6123,N_5687,N_5081);
xor U6124 (N_6124,N_5329,N_5318);
xnor U6125 (N_6125,N_5146,N_5886);
or U6126 (N_6126,N_5693,N_4850);
and U6127 (N_6127,N_4080,N_5337);
or U6128 (N_6128,N_5220,N_4678);
or U6129 (N_6129,N_5286,N_4218);
nor U6130 (N_6130,N_5534,N_5612);
and U6131 (N_6131,N_4449,N_4287);
nor U6132 (N_6132,N_5042,N_5842);
or U6133 (N_6133,N_4753,N_5793);
nand U6134 (N_6134,N_4038,N_4325);
nand U6135 (N_6135,N_5261,N_5908);
or U6136 (N_6136,N_5945,N_5759);
nor U6137 (N_6137,N_4107,N_4297);
nand U6138 (N_6138,N_4631,N_5923);
or U6139 (N_6139,N_5798,N_5149);
xor U6140 (N_6140,N_4464,N_4942);
and U6141 (N_6141,N_4090,N_5244);
and U6142 (N_6142,N_4504,N_4071);
or U6143 (N_6143,N_5757,N_4007);
nand U6144 (N_6144,N_4814,N_5992);
xnor U6145 (N_6145,N_4394,N_5881);
nand U6146 (N_6146,N_4569,N_5136);
xor U6147 (N_6147,N_5241,N_4934);
xor U6148 (N_6148,N_4996,N_4281);
nor U6149 (N_6149,N_5413,N_4623);
or U6150 (N_6150,N_5347,N_5073);
nand U6151 (N_6151,N_5121,N_4131);
nor U6152 (N_6152,N_5603,N_4432);
or U6153 (N_6153,N_5546,N_5742);
or U6154 (N_6154,N_4896,N_5205);
nand U6155 (N_6155,N_4455,N_4369);
and U6156 (N_6156,N_4916,N_4614);
or U6157 (N_6157,N_4143,N_5267);
or U6158 (N_6158,N_4710,N_5691);
and U6159 (N_6159,N_4647,N_4978);
xor U6160 (N_6160,N_5022,N_5948);
xor U6161 (N_6161,N_4104,N_4553);
or U6162 (N_6162,N_4737,N_5724);
nor U6163 (N_6163,N_4035,N_5201);
nor U6164 (N_6164,N_4396,N_4757);
and U6165 (N_6165,N_4565,N_4214);
and U6166 (N_6166,N_5018,N_4468);
nand U6167 (N_6167,N_5796,N_5151);
and U6168 (N_6168,N_4306,N_4759);
or U6169 (N_6169,N_4842,N_4291);
nor U6170 (N_6170,N_4881,N_4911);
nor U6171 (N_6171,N_5837,N_4834);
nor U6172 (N_6172,N_4384,N_5739);
or U6173 (N_6173,N_5057,N_4509);
or U6174 (N_6174,N_4409,N_4442);
xor U6175 (N_6175,N_4051,N_5483);
xnor U6176 (N_6176,N_4410,N_5521);
or U6177 (N_6177,N_5177,N_5816);
xor U6178 (N_6178,N_4546,N_4229);
and U6179 (N_6179,N_4863,N_5446);
and U6180 (N_6180,N_4169,N_4215);
and U6181 (N_6181,N_4868,N_5884);
and U6182 (N_6182,N_5529,N_5011);
or U6183 (N_6183,N_5914,N_5533);
xor U6184 (N_6184,N_4572,N_5450);
nor U6185 (N_6185,N_5728,N_5028);
and U6186 (N_6186,N_4522,N_5518);
nor U6187 (N_6187,N_5363,N_4054);
or U6188 (N_6188,N_5336,N_4755);
nor U6189 (N_6189,N_4463,N_4785);
or U6190 (N_6190,N_5032,N_4575);
xnor U6191 (N_6191,N_4433,N_5690);
nor U6192 (N_6192,N_4889,N_5637);
or U6193 (N_6193,N_5288,N_5907);
xnor U6194 (N_6194,N_4172,N_5718);
and U6195 (N_6195,N_4327,N_5501);
or U6196 (N_6196,N_5478,N_4492);
xnor U6197 (N_6197,N_4791,N_5280);
or U6198 (N_6198,N_5110,N_5913);
nor U6199 (N_6199,N_5176,N_4680);
nor U6200 (N_6200,N_5463,N_5775);
nand U6201 (N_6201,N_5526,N_4405);
and U6202 (N_6202,N_5708,N_4004);
nand U6203 (N_6203,N_4789,N_4363);
xnor U6204 (N_6204,N_4998,N_5577);
nor U6205 (N_6205,N_5129,N_5756);
xor U6206 (N_6206,N_4940,N_4118);
nor U6207 (N_6207,N_4393,N_5372);
xnor U6208 (N_6208,N_4949,N_5575);
or U6209 (N_6209,N_4700,N_4238);
and U6210 (N_6210,N_4285,N_5341);
and U6211 (N_6211,N_5476,N_4894);
and U6212 (N_6212,N_4793,N_4947);
or U6213 (N_6213,N_4627,N_4952);
and U6214 (N_6214,N_5882,N_4158);
and U6215 (N_6215,N_5953,N_4805);
and U6216 (N_6216,N_5324,N_5264);
xor U6217 (N_6217,N_4716,N_5894);
xor U6218 (N_6218,N_4308,N_5194);
xnor U6219 (N_6219,N_4348,N_4109);
xor U6220 (N_6220,N_4168,N_5920);
nor U6221 (N_6221,N_5570,N_4273);
or U6222 (N_6222,N_5542,N_4244);
nor U6223 (N_6223,N_5573,N_4230);
and U6224 (N_6224,N_4877,N_5782);
nor U6225 (N_6225,N_4101,N_4893);
nand U6226 (N_6226,N_4420,N_5424);
nand U6227 (N_6227,N_5459,N_4267);
nand U6228 (N_6228,N_4856,N_5184);
or U6229 (N_6229,N_5202,N_5584);
nor U6230 (N_6230,N_5167,N_4258);
xor U6231 (N_6231,N_5969,N_4827);
nor U6232 (N_6232,N_4826,N_5338);
or U6233 (N_6233,N_5351,N_5680);
nand U6234 (N_6234,N_4484,N_4519);
nor U6235 (N_6235,N_5187,N_4152);
and U6236 (N_6236,N_4733,N_5436);
and U6237 (N_6237,N_5678,N_4711);
xor U6238 (N_6238,N_5094,N_4845);
xor U6239 (N_6239,N_5265,N_4573);
xnor U6240 (N_6240,N_4021,N_4879);
nor U6241 (N_6241,N_4626,N_4005);
or U6242 (N_6242,N_4968,N_5232);
and U6243 (N_6243,N_4276,N_4862);
nor U6244 (N_6244,N_5326,N_4648);
nand U6245 (N_6245,N_5069,N_4794);
nand U6246 (N_6246,N_5937,N_4239);
or U6247 (N_6247,N_4165,N_5222);
nor U6248 (N_6248,N_5611,N_4910);
or U6249 (N_6249,N_5159,N_5621);
and U6250 (N_6250,N_4319,N_4435);
xor U6251 (N_6251,N_4212,N_4389);
xor U6252 (N_6252,N_5827,N_5448);
and U6253 (N_6253,N_5270,N_5433);
or U6254 (N_6254,N_4748,N_4288);
nor U6255 (N_6255,N_4401,N_4963);
nand U6256 (N_6256,N_5500,N_5043);
xor U6257 (N_6257,N_4205,N_5972);
nand U6258 (N_6258,N_4870,N_5963);
xnor U6259 (N_6259,N_5853,N_5942);
nand U6260 (N_6260,N_5044,N_4489);
nor U6261 (N_6261,N_5561,N_5359);
and U6262 (N_6262,N_4503,N_5503);
nor U6263 (N_6263,N_4724,N_5466);
and U6264 (N_6264,N_5799,N_5921);
nor U6265 (N_6265,N_5789,N_5315);
or U6266 (N_6266,N_5150,N_4413);
or U6267 (N_6267,N_4965,N_5762);
nand U6268 (N_6268,N_5829,N_5547);
nand U6269 (N_6269,N_5906,N_5163);
and U6270 (N_6270,N_5308,N_4381);
and U6271 (N_6271,N_4182,N_4458);
nand U6272 (N_6272,N_4309,N_5048);
or U6273 (N_6273,N_5717,N_4491);
nor U6274 (N_6274,N_4596,N_4174);
or U6275 (N_6275,N_4217,N_4370);
nor U6276 (N_6276,N_5246,N_5875);
xnor U6277 (N_6277,N_4951,N_5689);
nand U6278 (N_6278,N_5200,N_4112);
nand U6279 (N_6279,N_4762,N_5373);
or U6280 (N_6280,N_4037,N_4017);
xor U6281 (N_6281,N_4154,N_4429);
and U6282 (N_6282,N_4810,N_5260);
nor U6283 (N_6283,N_4156,N_5970);
and U6284 (N_6284,N_4977,N_5625);
or U6285 (N_6285,N_4971,N_4529);
and U6286 (N_6286,N_4732,N_4772);
and U6287 (N_6287,N_4177,N_4566);
nand U6288 (N_6288,N_5454,N_4294);
xor U6289 (N_6289,N_4180,N_4608);
or U6290 (N_6290,N_4190,N_5880);
or U6291 (N_6291,N_4441,N_5815);
nor U6292 (N_6292,N_4039,N_4729);
nand U6293 (N_6293,N_5139,N_4597);
and U6294 (N_6294,N_4453,N_4690);
nor U6295 (N_6295,N_5033,N_5806);
xnor U6296 (N_6296,N_4590,N_5902);
and U6297 (N_6297,N_4661,N_4831);
or U6298 (N_6298,N_5218,N_4480);
or U6299 (N_6299,N_4262,N_5078);
xor U6300 (N_6300,N_5925,N_4034);
or U6301 (N_6301,N_5538,N_5455);
nand U6302 (N_6302,N_4593,N_5166);
and U6303 (N_6303,N_4457,N_4632);
or U6304 (N_6304,N_5753,N_5061);
xnor U6305 (N_6305,N_4820,N_5740);
nand U6306 (N_6306,N_4027,N_5157);
or U6307 (N_6307,N_5883,N_5545);
nor U6308 (N_6308,N_5685,N_4502);
and U6309 (N_6309,N_4891,N_4697);
nor U6310 (N_6310,N_4725,N_4137);
and U6311 (N_6311,N_4259,N_4053);
nor U6312 (N_6312,N_5160,N_4905);
nand U6313 (N_6313,N_4941,N_4567);
and U6314 (N_6314,N_4914,N_5732);
or U6315 (N_6315,N_5564,N_5233);
and U6316 (N_6316,N_4026,N_4835);
and U6317 (N_6317,N_5844,N_4561);
nand U6318 (N_6318,N_5903,N_5909);
nand U6319 (N_6319,N_4917,N_4178);
xor U6320 (N_6320,N_5745,N_5223);
and U6321 (N_6321,N_5831,N_5860);
or U6322 (N_6322,N_5170,N_4923);
xnor U6323 (N_6323,N_4081,N_4847);
and U6324 (N_6324,N_4639,N_4600);
or U6325 (N_6325,N_5549,N_5015);
nand U6326 (N_6326,N_5539,N_4451);
and U6327 (N_6327,N_4610,N_5105);
nor U6328 (N_6328,N_5965,N_5608);
nor U6329 (N_6329,N_5104,N_4098);
or U6330 (N_6330,N_5224,N_5375);
and U6331 (N_6331,N_5769,N_4970);
nor U6332 (N_6332,N_4321,N_4078);
and U6333 (N_6333,N_4837,N_4734);
nor U6334 (N_6334,N_5169,N_5311);
and U6335 (N_6335,N_4620,N_5898);
or U6336 (N_6336,N_4097,N_5841);
nor U6337 (N_6337,N_4520,N_5935);
or U6338 (N_6338,N_4301,N_5997);
xor U6339 (N_6339,N_4674,N_5026);
nor U6340 (N_6340,N_4022,N_4320);
or U6341 (N_6341,N_5493,N_5553);
nand U6342 (N_6342,N_4578,N_4749);
nand U6343 (N_6343,N_5996,N_4829);
nor U6344 (N_6344,N_5786,N_5522);
xnor U6345 (N_6345,N_5768,N_4279);
xor U6346 (N_6346,N_5357,N_4549);
and U6347 (N_6347,N_4904,N_5868);
xor U6348 (N_6348,N_4851,N_4006);
and U6349 (N_6349,N_4201,N_5152);
or U6350 (N_6350,N_5671,N_4465);
xor U6351 (N_6351,N_5305,N_4994);
xor U6352 (N_6352,N_5511,N_5249);
nand U6353 (N_6353,N_5662,N_5554);
or U6354 (N_6354,N_5300,N_5301);
and U6355 (N_6355,N_5623,N_5393);
and U6356 (N_6356,N_4434,N_4510);
and U6357 (N_6357,N_5939,N_4117);
xnor U6358 (N_6358,N_4299,N_4114);
or U6359 (N_6359,N_4920,N_5289);
xnor U6360 (N_6360,N_5808,N_4960);
nor U6361 (N_6361,N_5781,N_5686);
nor U6362 (N_6362,N_4602,N_4014);
nand U6363 (N_6363,N_5597,N_5297);
and U6364 (N_6364,N_4474,N_5192);
and U6365 (N_6365,N_5414,N_4028);
nand U6366 (N_6366,N_5140,N_4984);
xor U6367 (N_6367,N_4607,N_5833);
and U6368 (N_6368,N_4992,N_4326);
nor U6369 (N_6369,N_4024,N_5481);
and U6370 (N_6370,N_4040,N_4548);
nor U6371 (N_6371,N_5675,N_5928);
nor U6372 (N_6372,N_4551,N_4495);
and U6373 (N_6373,N_4494,N_5967);
nand U6374 (N_6374,N_5314,N_5968);
and U6375 (N_6375,N_4485,N_5715);
nand U6376 (N_6376,N_5635,N_5103);
xor U6377 (N_6377,N_4425,N_5592);
nand U6378 (N_6378,N_5470,N_4946);
nor U6379 (N_6379,N_4828,N_5096);
nor U6380 (N_6380,N_4900,N_5838);
nand U6381 (N_6381,N_4450,N_4903);
xor U6382 (N_6382,N_5591,N_5867);
xor U6383 (N_6383,N_4208,N_4932);
nor U6384 (N_6384,N_5544,N_5425);
nor U6385 (N_6385,N_4899,N_4873);
nand U6386 (N_6386,N_5574,N_4226);
xnor U6387 (N_6387,N_5610,N_4606);
nor U6388 (N_6388,N_4642,N_4776);
nand U6389 (N_6389,N_5700,N_5566);
or U6390 (N_6390,N_5080,N_4640);
nand U6391 (N_6391,N_4382,N_5460);
nand U6392 (N_6392,N_4331,N_4121);
xor U6393 (N_6393,N_4368,N_4421);
xor U6394 (N_6394,N_5090,N_4380);
and U6395 (N_6395,N_5343,N_4576);
or U6396 (N_6396,N_4630,N_5025);
nor U6397 (N_6397,N_4507,N_5688);
nand U6398 (N_6398,N_5231,N_5633);
nor U6399 (N_6399,N_4138,N_5763);
or U6400 (N_6400,N_4803,N_5989);
or U6401 (N_6401,N_4671,N_4280);
nand U6402 (N_6402,N_4362,N_5355);
nand U6403 (N_6403,N_5127,N_5214);
and U6404 (N_6404,N_4194,N_5029);
nor U6405 (N_6405,N_5156,N_5741);
or U6406 (N_6406,N_4096,N_5516);
nor U6407 (N_6407,N_4715,N_5692);
nand U6408 (N_6408,N_4541,N_5407);
or U6409 (N_6409,N_5190,N_5896);
or U6410 (N_6410,N_4261,N_4644);
xnor U6411 (N_6411,N_5496,N_4612);
or U6412 (N_6412,N_5852,N_4783);
xor U6413 (N_6413,N_4047,N_4094);
or U6414 (N_6414,N_4599,N_5079);
xnor U6415 (N_6415,N_5112,N_5643);
xnor U6416 (N_6416,N_5388,N_5706);
nand U6417 (N_6417,N_4908,N_4539);
or U6418 (N_6418,N_4412,N_4676);
nand U6419 (N_6419,N_5528,N_5344);
or U6420 (N_6420,N_5579,N_5394);
or U6421 (N_6421,N_4136,N_4476);
and U6422 (N_6422,N_4203,N_5982);
nor U6423 (N_6423,N_5998,N_4189);
or U6424 (N_6424,N_4592,N_4290);
nand U6425 (N_6425,N_5962,N_5475);
and U6426 (N_6426,N_5649,N_5787);
nand U6427 (N_6427,N_4153,N_5255);
nand U6428 (N_6428,N_5569,N_5091);
nand U6429 (N_6429,N_4843,N_4085);
and U6430 (N_6430,N_5940,N_4068);
and U6431 (N_6431,N_5543,N_4527);
nand U6432 (N_6432,N_4611,N_4937);
nand U6433 (N_6433,N_4782,N_5451);
nor U6434 (N_6434,N_4665,N_4801);
xor U6435 (N_6435,N_4166,N_4270);
and U6436 (N_6436,N_4679,N_5924);
nand U6437 (N_6437,N_5247,N_4838);
and U6438 (N_6438,N_4105,N_5135);
xnor U6439 (N_6439,N_5823,N_4651);
or U6440 (N_6440,N_5901,N_4479);
and U6441 (N_6441,N_5857,N_4033);
and U6442 (N_6442,N_5422,N_4415);
nor U6443 (N_6443,N_5307,N_5813);
nor U6444 (N_6444,N_4340,N_4307);
or U6445 (N_6445,N_4585,N_4388);
nand U6446 (N_6446,N_4337,N_5598);
or U6447 (N_6447,N_4354,N_5339);
xnor U6448 (N_6448,N_4408,N_5877);
nor U6449 (N_6449,N_5790,N_4641);
xnor U6450 (N_6450,N_4601,N_4045);
or U6451 (N_6451,N_5378,N_5679);
xnor U6452 (N_6452,N_5240,N_4113);
or U6453 (N_6453,N_5087,N_4141);
and U6454 (N_6454,N_4617,N_5814);
and U6455 (N_6455,N_5705,N_4574);
nor U6456 (N_6456,N_5005,N_4933);
or U6457 (N_6457,N_4176,N_4397);
nand U6458 (N_6458,N_5158,N_5368);
nand U6459 (N_6459,N_4358,N_4557);
and U6460 (N_6460,N_4251,N_5406);
nor U6461 (N_6461,N_5178,N_4123);
xnor U6462 (N_6462,N_4221,N_5108);
nand U6463 (N_6463,N_5001,N_5974);
and U6464 (N_6464,N_5683,N_5472);
nand U6465 (N_6465,N_5666,N_4231);
and U6466 (N_6466,N_5586,N_4906);
or U6467 (N_6467,N_5376,N_4315);
and U6468 (N_6468,N_4764,N_4061);
or U6469 (N_6469,N_5230,N_4437);
nand U6470 (N_6470,N_4197,N_4619);
nand U6471 (N_6471,N_4852,N_4042);
nor U6472 (N_6472,N_5327,N_5273);
and U6473 (N_6473,N_5234,N_4645);
or U6474 (N_6474,N_5431,N_5593);
or U6475 (N_6475,N_5774,N_4379);
nor U6476 (N_6476,N_5401,N_4653);
or U6477 (N_6477,N_4858,N_4670);
or U6478 (N_6478,N_5086,N_4582);
or U6479 (N_6479,N_5071,N_4846);
nor U6480 (N_6480,N_4588,N_4874);
xnor U6481 (N_6481,N_5316,N_4875);
nor U6482 (N_6482,N_4677,N_4469);
xor U6483 (N_6483,N_4770,N_4699);
nor U6484 (N_6484,N_5024,N_4773);
nand U6485 (N_6485,N_4472,N_4543);
and U6486 (N_6486,N_4861,N_5760);
or U6487 (N_6487,N_4571,N_5352);
nor U6488 (N_6488,N_5412,N_5469);
xnor U6489 (N_6489,N_4356,N_4777);
and U6490 (N_6490,N_4853,N_5007);
nor U6491 (N_6491,N_5107,N_5932);
and U6492 (N_6492,N_4691,N_4213);
nor U6493 (N_6493,N_4961,N_5933);
and U6494 (N_6494,N_5293,N_4295);
and U6495 (N_6495,N_5514,N_4806);
or U6496 (N_6496,N_4817,N_4145);
and U6497 (N_6497,N_4743,N_5302);
nor U6498 (N_6498,N_4672,N_4701);
and U6499 (N_6499,N_4075,N_5985);
xor U6500 (N_6500,N_5936,N_5990);
xnor U6501 (N_6501,N_4020,N_4568);
nor U6502 (N_6502,N_4350,N_4142);
xnor U6503 (N_6503,N_4272,N_5788);
and U6504 (N_6504,N_4092,N_5531);
nor U6505 (N_6505,N_4058,N_4884);
or U6506 (N_6506,N_4505,N_5477);
xnor U6507 (N_6507,N_4663,N_4811);
or U6508 (N_6508,N_4120,N_5148);
or U6509 (N_6509,N_4242,N_5832);
and U6510 (N_6510,N_4373,N_5869);
nor U6511 (N_6511,N_4921,N_5132);
nand U6512 (N_6512,N_4225,N_5216);
nand U6513 (N_6513,N_5171,N_5758);
and U6514 (N_6514,N_5027,N_5807);
xor U6515 (N_6515,N_4305,N_4860);
xor U6516 (N_6516,N_4129,N_4057);
nand U6517 (N_6517,N_5092,N_5978);
xnor U6518 (N_6518,N_5053,N_4030);
and U6519 (N_6519,N_4329,N_4456);
and U6520 (N_6520,N_5710,N_4709);
nand U6521 (N_6521,N_4001,N_4443);
nor U6522 (N_6522,N_4377,N_4493);
and U6523 (N_6523,N_4634,N_4278);
nand U6524 (N_6524,N_5862,N_5124);
nand U6525 (N_6525,N_4013,N_4533);
and U6526 (N_6526,N_5003,N_4615);
or U6527 (N_6527,N_5512,N_5130);
xnor U6528 (N_6528,N_4560,N_5065);
and U6529 (N_6529,N_4292,N_5185);
nor U6530 (N_6530,N_5164,N_5468);
xnor U6531 (N_6531,N_5382,N_5137);
or U6532 (N_6532,N_5445,N_5958);
or U6533 (N_6533,N_5115,N_5279);
nor U6534 (N_6534,N_4559,N_4973);
nor U6535 (N_6535,N_4750,N_4635);
nand U6536 (N_6536,N_4019,N_4945);
xnor U6537 (N_6537,N_4146,N_5749);
xnor U6538 (N_6538,N_4512,N_5750);
nand U6539 (N_6539,N_4895,N_5523);
xnor U6540 (N_6540,N_5922,N_4754);
nand U6541 (N_6541,N_4335,N_4452);
xor U6542 (N_6542,N_4416,N_5888);
xor U6543 (N_6543,N_4360,N_5846);
or U6544 (N_6544,N_5820,N_4304);
nor U6545 (N_6545,N_4719,N_4912);
or U6546 (N_6546,N_4500,N_4778);
or U6547 (N_6547,N_4414,N_4840);
or U6548 (N_6548,N_5627,N_5981);
or U6549 (N_6549,N_5055,N_5228);
or U6550 (N_6550,N_4275,N_4515);
xnor U6551 (N_6551,N_5186,N_5755);
xor U6552 (N_6552,N_5058,N_4707);
nor U6553 (N_6553,N_5034,N_5804);
xnor U6554 (N_6554,N_5144,N_5817);
and U6555 (N_6555,N_4025,N_5095);
nand U6556 (N_6556,N_4387,N_5792);
and U6557 (N_6557,N_5119,N_5905);
xor U6558 (N_6558,N_5810,N_5839);
or U6559 (N_6559,N_5640,N_5917);
nor U6560 (N_6560,N_4915,N_5046);
or U6561 (N_6561,N_4473,N_4530);
xor U6562 (N_6562,N_4398,N_5384);
nand U6563 (N_6563,N_5606,N_4077);
xor U6564 (N_6564,N_5559,N_4151);
and U6565 (N_6565,N_4739,N_4140);
or U6566 (N_6566,N_4471,N_5652);
nand U6567 (N_6567,N_4741,N_5189);
nor U6568 (N_6568,N_5117,N_4646);
nor U6569 (N_6569,N_5485,N_5765);
and U6570 (N_6570,N_5172,N_5221);
nor U6571 (N_6571,N_5208,N_5097);
nor U6572 (N_6572,N_5325,N_4181);
xnor U6573 (N_6573,N_5614,N_5440);
nand U6574 (N_6574,N_4486,N_4312);
or U6575 (N_6575,N_5889,N_4193);
and U6576 (N_6576,N_5673,N_4580);
xor U6577 (N_6577,N_4302,N_5707);
nand U6578 (N_6578,N_4531,N_4736);
or U6579 (N_6579,N_5949,N_5072);
nand U6580 (N_6580,N_4046,N_4545);
nand U6581 (N_6581,N_4943,N_5243);
nand U6582 (N_6582,N_5489,N_5966);
and U6583 (N_6583,N_5084,N_4579);
and U6584 (N_6584,N_4986,N_5154);
xor U6585 (N_6585,N_4002,N_5764);
and U6586 (N_6586,N_5947,N_4079);
nor U6587 (N_6587,N_5056,N_4704);
xor U6588 (N_6588,N_5410,N_4490);
xor U6589 (N_6589,N_4695,N_5605);
nand U6590 (N_6590,N_4342,N_4909);
and U6591 (N_6591,N_5870,N_4403);
nand U6592 (N_6592,N_5443,N_4132);
nand U6593 (N_6593,N_5126,N_4108);
and U6594 (N_6594,N_5013,N_5142);
nand U6595 (N_6595,N_5858,N_4015);
and U6596 (N_6596,N_5335,N_5462);
xor U6597 (N_6597,N_5345,N_4686);
nand U6598 (N_6598,N_5555,N_5282);
xnor U6599 (N_6599,N_5694,N_4767);
nor U6600 (N_6600,N_4746,N_4171);
or U6601 (N_6601,N_5118,N_5143);
nor U6602 (N_6602,N_5650,N_4538);
nand U6603 (N_6603,N_4769,N_5195);
xor U6604 (N_6604,N_4352,N_5106);
nor U6605 (N_6605,N_4664,N_5629);
nand U6606 (N_6606,N_4523,N_4161);
nor U6607 (N_6607,N_5367,N_5669);
or U6608 (N_6608,N_5733,N_4747);
nand U6609 (N_6609,N_5977,N_4357);
or U6610 (N_6610,N_4252,N_5320);
nand U6611 (N_6611,N_5713,N_5467);
nor U6612 (N_6612,N_4298,N_4804);
nand U6613 (N_6613,N_5257,N_4913);
nand U6614 (N_6614,N_5491,N_4106);
and U6615 (N_6615,N_5465,N_4950);
or U6616 (N_6616,N_4284,N_5276);
and U6617 (N_6617,N_4637,N_5979);
nand U6618 (N_6618,N_5390,N_5362);
nand U6619 (N_6619,N_4459,N_5391);
nand U6620 (N_6620,N_4438,N_5009);
or U6621 (N_6621,N_5490,N_5797);
xnor U6622 (N_6622,N_5719,N_5100);
nand U6623 (N_6623,N_5077,N_4236);
nand U6624 (N_6624,N_5658,N_5198);
nand U6625 (N_6625,N_5229,N_4423);
and U6626 (N_6626,N_5830,N_4470);
nor U6627 (N_6627,N_5131,N_4497);
and U6628 (N_6628,N_5580,N_5021);
nand U6629 (N_6629,N_4516,N_4657);
nor U6630 (N_6630,N_5147,N_4655);
xnor U6631 (N_6631,N_4924,N_5317);
or U6632 (N_6632,N_5895,N_5892);
nor U6633 (N_6633,N_5873,N_5298);
nor U6634 (N_6634,N_5581,N_4535);
and U6635 (N_6635,N_5562,N_4372);
xnor U6636 (N_6636,N_5291,N_5197);
xnor U6637 (N_6637,N_4659,N_4584);
nor U6638 (N_6638,N_5155,N_4246);
and U6639 (N_6639,N_4447,N_4296);
xnor U6640 (N_6640,N_4927,N_5736);
xnor U6641 (N_6641,N_4404,N_5054);
xor U6642 (N_6642,N_4056,N_5596);
nor U6643 (N_6643,N_5174,N_5479);
and U6644 (N_6644,N_5698,N_4798);
or U6645 (N_6645,N_5607,N_5994);
xnor U6646 (N_6646,N_5415,N_4839);
xor U6647 (N_6647,N_5778,N_4907);
xnor U6648 (N_6648,N_5943,N_5039);
xor U6649 (N_6649,N_4224,N_5319);
and U6650 (N_6650,N_4314,N_5099);
or U6651 (N_6651,N_5125,N_4865);
and U6652 (N_6652,N_5380,N_4999);
or U6653 (N_6653,N_4892,N_5403);
or U6654 (N_6654,N_5225,N_4250);
nor U6655 (N_6655,N_5284,N_5421);
or U6656 (N_6656,N_5210,N_4454);
nor U6657 (N_6657,N_4544,N_4540);
and U6658 (N_6658,N_5441,N_5427);
or U6659 (N_6659,N_5711,N_5887);
nor U6660 (N_6660,N_5085,N_4199);
nor U6661 (N_6661,N_5510,N_4714);
xnor U6662 (N_6662,N_4583,N_5497);
nor U6663 (N_6663,N_4253,N_5017);
nand U6664 (N_6664,N_5773,N_4175);
nor U6665 (N_6665,N_5191,N_5504);
or U6666 (N_6666,N_4407,N_4111);
xor U6667 (N_6667,N_4256,N_5213);
and U6668 (N_6668,N_4855,N_5821);
nor U6669 (N_6669,N_5386,N_4790);
xnor U6670 (N_6670,N_4248,N_5632);
nor U6671 (N_6671,N_5524,N_5729);
nor U6672 (N_6672,N_4956,N_4095);
and U6673 (N_6673,N_5464,N_5181);
or U6674 (N_6674,N_5812,N_4330);
and U6675 (N_6675,N_5173,N_4082);
or U6676 (N_6676,N_5256,N_4603);
or U6677 (N_6677,N_5239,N_4185);
or U6678 (N_6678,N_4885,N_4564);
nand U6679 (N_6679,N_5392,N_4126);
and U6680 (N_6680,N_4066,N_4048);
nor U6681 (N_6681,N_4378,N_5950);
nor U6682 (N_6682,N_4618,N_5430);
nand U6683 (N_6683,N_4266,N_4888);
nand U6684 (N_6684,N_5861,N_4625);
and U6685 (N_6685,N_5452,N_5432);
nand U6686 (N_6686,N_5532,N_4930);
or U6687 (N_6687,N_5735,N_5890);
or U6688 (N_6688,N_5854,N_4311);
nand U6689 (N_6689,N_4365,N_4953);
nand U6690 (N_6690,N_4072,N_5576);
nor U6691 (N_6691,N_4765,N_5168);
and U6692 (N_6692,N_5646,N_5803);
nor U6693 (N_6693,N_4487,N_5530);
nor U6694 (N_6694,N_4124,N_4070);
nor U6695 (N_6695,N_4255,N_4735);
xnor U6696 (N_6696,N_5976,N_4705);
and U6697 (N_6697,N_5938,N_4744);
xor U6698 (N_6698,N_4962,N_4044);
nor U6699 (N_6699,N_5826,N_5613);
and U6700 (N_6700,N_4740,N_4922);
xor U6701 (N_6701,N_4993,N_5585);
nor U6702 (N_6702,N_4675,N_5871);
nor U6703 (N_6703,N_4324,N_4498);
and U6704 (N_6704,N_5552,N_4198);
xor U6705 (N_6705,N_5134,N_5916);
nand U6706 (N_6706,N_5203,N_4802);
and U6707 (N_6707,N_4184,N_5681);
or U6708 (N_6708,N_5619,N_4460);
or U6709 (N_6709,N_4050,N_4819);
or U6710 (N_6710,N_4424,N_4245);
nor U6711 (N_6711,N_5930,N_4730);
nand U6712 (N_6712,N_5383,N_5405);
nor U6713 (N_6713,N_5776,N_4257);
and U6714 (N_6714,N_4417,N_4406);
and U6715 (N_6715,N_4669,N_5045);
or U6716 (N_6716,N_4938,N_4110);
and U6717 (N_6717,N_5609,N_4233);
xor U6718 (N_6718,N_4247,N_5849);
nand U6719 (N_6719,N_4065,N_4849);
xnor U6720 (N_6720,N_4192,N_5638);
nor U6721 (N_6721,N_5381,N_4062);
or U6722 (N_6722,N_5052,N_4202);
and U6723 (N_6723,N_4333,N_5704);
or U6724 (N_6724,N_4436,N_5944);
xnor U6725 (N_6725,N_4427,N_5340);
and U6726 (N_6726,N_4195,N_4100);
nor U6727 (N_6727,N_5458,N_4763);
nand U6728 (N_6728,N_5602,N_4681);
xnor U6729 (N_6729,N_4563,N_4440);
xnor U6730 (N_6730,N_5417,N_4867);
nor U6731 (N_6731,N_4886,N_5290);
nand U6732 (N_6732,N_5836,N_4122);
or U6733 (N_6733,N_5418,N_4605);
or U6734 (N_6734,N_5934,N_5899);
or U6735 (N_6735,N_5556,N_5138);
nand U6736 (N_6736,N_5927,N_4235);
nand U6737 (N_6737,N_4428,N_4374);
or U6738 (N_6738,N_5141,N_5515);
or U6739 (N_6739,N_4345,N_5665);
xnor U6740 (N_6740,N_5473,N_4728);
nor U6741 (N_6741,N_5350,N_4800);
nor U6742 (N_6742,N_4967,N_5957);
xnor U6743 (N_6743,N_5332,N_5361);
and U6744 (N_6744,N_5560,N_4063);
nor U6745 (N_6745,N_5802,N_5050);
or U6746 (N_6746,N_5349,N_5851);
nand U6747 (N_6747,N_4223,N_5333);
and U6748 (N_6748,N_5663,N_4206);
nor U6749 (N_6749,N_5457,N_5670);
and U6750 (N_6750,N_5964,N_5444);
and U6751 (N_6751,N_5604,N_5281);
nor U6752 (N_6752,N_4310,N_4446);
xor U6753 (N_6753,N_4191,N_4073);
nand U6754 (N_6754,N_4866,N_5217);
nand U6755 (N_6755,N_5959,N_5269);
xnor U6756 (N_6756,N_4008,N_5712);
nand U6757 (N_6757,N_4988,N_4570);
xor U6758 (N_6758,N_5321,N_4170);
and U6759 (N_6759,N_4032,N_5991);
nor U6760 (N_6760,N_5060,N_4717);
nand U6761 (N_6761,N_4825,N_5506);
or U6762 (N_6762,N_5482,N_4622);
nand U6763 (N_6763,N_5000,N_5520);
xnor U6764 (N_6764,N_5897,N_5020);
or U6765 (N_6765,N_4628,N_5617);
xnor U6766 (N_6766,N_5674,N_4127);
and U6767 (N_6767,N_4196,N_5063);
nor U6768 (N_6768,N_4931,N_5587);
nand U6769 (N_6769,N_5840,N_4972);
xor U6770 (N_6770,N_4784,N_5805);
nor U6771 (N_6771,N_4689,N_5956);
and U6772 (N_6772,N_5439,N_4018);
xnor U6773 (N_6773,N_5395,N_4525);
nand U6774 (N_6774,N_5161,N_5508);
and U6775 (N_6775,N_5165,N_5088);
and U6776 (N_6776,N_4696,N_5004);
nor U6777 (N_6777,N_5660,N_4562);
or U6778 (N_6778,N_5513,N_5709);
nor U6779 (N_6779,N_4976,N_5277);
nor U6780 (N_6780,N_4254,N_5616);
xor U6781 (N_6781,N_4859,N_5387);
nor U6782 (N_6782,N_5365,N_4928);
xor U6783 (N_6783,N_4232,N_4514);
and U6784 (N_6784,N_4621,N_4237);
nand U6785 (N_6785,N_5594,N_5429);
nor U6786 (N_6786,N_5064,N_5494);
and U6787 (N_6787,N_4959,N_5236);
xnor U6788 (N_6788,N_5835,N_5114);
nor U6789 (N_6789,N_4426,N_5565);
xnor U6790 (N_6790,N_5695,N_5283);
xor U6791 (N_6791,N_4925,N_4808);
or U6792 (N_6792,N_5245,N_5411);
and U6793 (N_6793,N_4445,N_5461);
nand U6794 (N_6794,N_4702,N_4974);
and U6795 (N_6795,N_4816,N_4086);
or U6796 (N_6796,N_4128,N_5589);
xnor U6797 (N_6797,N_5258,N_5180);
nor U6798 (N_6798,N_4303,N_5354);
xor U6799 (N_6799,N_4718,N_5737);
nand U6800 (N_6800,N_5309,N_4462);
xnor U6801 (N_6801,N_5828,N_4935);
nand U6802 (N_6802,N_5328,N_5006);
xnor U6803 (N_6803,N_4809,N_4587);
nor U6804 (N_6804,N_4534,N_4983);
or U6805 (N_6805,N_4103,N_4052);
nand U6806 (N_6806,N_5480,N_4316);
or U6807 (N_6807,N_5253,N_5111);
or U6808 (N_6808,N_4518,N_4948);
nor U6809 (N_6809,N_4982,N_4528);
nor U6810 (N_6810,N_4419,N_5519);
or U6811 (N_6811,N_5639,N_4722);
xor U6812 (N_6812,N_4880,N_4824);
or U6813 (N_6813,N_5672,N_5879);
and U6814 (N_6814,N_5334,N_5578);
nand U6815 (N_6815,N_5271,N_5397);
nor U6816 (N_6816,N_5259,N_4293);
nand U6817 (N_6817,N_5684,N_5525);
or U6818 (N_6818,N_5779,N_5811);
xnor U6819 (N_6819,N_4064,N_4668);
nor U6820 (N_6820,N_5929,N_4300);
or U6821 (N_6821,N_4227,N_5772);
xor U6822 (N_6822,N_4069,N_4521);
nand U6823 (N_6823,N_5036,N_5047);
or U6824 (N_6824,N_5716,N_5299);
xnor U6825 (N_6825,N_5696,N_5720);
nor U6826 (N_6826,N_5550,N_4771);
nor U6827 (N_6827,N_4322,N_4249);
xnor U6828 (N_6828,N_4989,N_4344);
and U6829 (N_6829,N_4243,N_4395);
nand U6830 (N_6830,N_5385,N_4919);
and U6831 (N_6831,N_5389,N_4643);
and U6832 (N_6832,N_4144,N_4964);
and U6833 (N_6833,N_4336,N_5878);
nand U6834 (N_6834,N_4731,N_5551);
nor U6835 (N_6835,N_4011,N_5449);
xnor U6836 (N_6836,N_4636,N_5182);
and U6837 (N_6837,N_4786,N_4633);
or U6838 (N_6838,N_5275,N_4475);
xnor U6839 (N_6839,N_4003,N_5859);
nand U6840 (N_6840,N_5358,N_4836);
nand U6841 (N_6841,N_5651,N_5636);
nor U6842 (N_6842,N_5254,N_4821);
and U6843 (N_6843,N_5630,N_5263);
nor U6844 (N_6844,N_5030,N_5049);
and U6845 (N_6845,N_4758,N_5668);
nand U6846 (N_6846,N_5571,N_5010);
nor U6847 (N_6847,N_5941,N_4083);
or U6848 (N_6848,N_5398,N_5960);
nand U6849 (N_6849,N_5008,N_5701);
nor U6850 (N_6850,N_5919,N_5785);
or U6851 (N_6851,N_5848,N_4173);
nand U6852 (N_6852,N_4526,N_5093);
xor U6853 (N_6853,N_5866,N_4815);
nand U6854 (N_6854,N_5618,N_4461);
xnor U6855 (N_6855,N_5548,N_4768);
xor U6856 (N_6856,N_4339,N_4694);
xor U6857 (N_6857,N_4163,N_5558);
xor U6858 (N_6858,N_4102,N_4055);
nor U6859 (N_6859,N_4887,N_5874);
and U6860 (N_6860,N_4074,N_4532);
or U6861 (N_6861,N_4658,N_5101);
and U6862 (N_6862,N_4985,N_5600);
and U6863 (N_6863,N_5242,N_4706);
or U6864 (N_6864,N_5074,N_5206);
xor U6865 (N_6865,N_4712,N_4752);
or U6866 (N_6866,N_4501,N_4130);
nor U6867 (N_6867,N_4125,N_5975);
nand U6868 (N_6868,N_4876,N_5484);
or U6869 (N_6869,N_4422,N_5487);
nor U6870 (N_6870,N_4787,N_4159);
and U6871 (N_6871,N_5645,N_5723);
nor U6872 (N_6872,N_5818,N_5656);
and U6873 (N_6873,N_4444,N_5067);
or U6874 (N_6874,N_5567,N_4673);
xnor U6875 (N_6875,N_5535,N_5396);
xor U6876 (N_6876,N_4467,N_4286);
and U6877 (N_6877,N_4349,N_4687);
xor U6878 (N_6878,N_5215,N_5453);
and U6879 (N_6879,N_5910,N_5648);
nor U6880 (N_6880,N_5035,N_5330);
nand U6881 (N_6881,N_5252,N_5404);
nand U6882 (N_6882,N_4751,N_5800);
and U6883 (N_6883,N_4313,N_5075);
nor U6884 (N_6884,N_5777,N_5702);
or U6885 (N_6885,N_4499,N_4656);
xnor U6886 (N_6886,N_5488,N_5379);
xnor U6887 (N_6887,N_4581,N_4882);
or U6888 (N_6888,N_4742,N_4283);
xor U6889 (N_6889,N_5183,N_5408);
nor U6890 (N_6890,N_5904,N_4872);
and U6891 (N_6891,N_5492,N_4390);
or U6892 (N_6892,N_4594,N_5423);
nor U6893 (N_6893,N_5973,N_5419);
nand U6894 (N_6894,N_5098,N_5926);
and U6895 (N_6895,N_5272,N_4595);
nand U6896 (N_6896,N_5102,N_5237);
nand U6897 (N_6897,N_5193,N_4150);
nor U6898 (N_6898,N_5287,N_5285);
nand U6899 (N_6899,N_4271,N_4347);
nand U6900 (N_6900,N_4060,N_5780);
or U6901 (N_6901,N_5588,N_5209);
or U6902 (N_6902,N_5040,N_4482);
nor U6903 (N_6903,N_5641,N_4954);
nand U6904 (N_6904,N_4991,N_4448);
nand U6905 (N_6905,N_5360,N_5876);
or U6906 (N_6906,N_5420,N_5128);
and U6907 (N_6907,N_5843,N_4430);
nor U6908 (N_6908,N_4059,N_5954);
nor U6909 (N_6909,N_5801,N_5918);
nor U6910 (N_6910,N_5748,N_4878);
and U6911 (N_6911,N_4537,N_4318);
or U6912 (N_6912,N_4832,N_5955);
nor U6913 (N_6913,N_5219,N_5059);
and U6914 (N_6914,N_4385,N_4431);
and U6915 (N_6915,N_5653,N_4957);
xor U6916 (N_6916,N_5893,N_4513);
or U6917 (N_6917,N_4517,N_5356);
or U6918 (N_6918,N_4936,N_5900);
or U6919 (N_6919,N_5031,N_5746);
nor U6920 (N_6920,N_5068,N_4036);
nand U6921 (N_6921,N_4598,N_5016);
xnor U6922 (N_6922,N_4264,N_5624);
xnor U6923 (N_6923,N_4089,N_5984);
and U6924 (N_6924,N_5582,N_5912);
or U6925 (N_6925,N_4341,N_5664);
xnor U6926 (N_6926,N_5442,N_4901);
nor U6927 (N_6927,N_5767,N_4155);
or U6928 (N_6928,N_4797,N_5725);
and U6929 (N_6929,N_5089,N_4135);
nor U6930 (N_6930,N_5070,N_5274);
nor U6931 (N_6931,N_5374,N_4616);
or U6932 (N_6932,N_5495,N_4955);
nand U6933 (N_6933,N_4399,N_4939);
or U6934 (N_6934,N_5434,N_5946);
and U6935 (N_6935,N_5377,N_5370);
nand U6936 (N_6936,N_5346,N_4554);
xnor U6937 (N_6937,N_5761,N_4650);
and U6938 (N_6938,N_4792,N_4116);
and U6939 (N_6939,N_5162,N_4604);
nand U6940 (N_6940,N_5784,N_5371);
xor U6941 (N_6941,N_5322,N_4812);
nor U6942 (N_6942,N_4638,N_5595);
and U6943 (N_6943,N_4662,N_4997);
nand U6944 (N_6944,N_4088,N_5369);
nor U6945 (N_6945,N_4788,N_5856);
xnor U6946 (N_6946,N_5557,N_4481);
and U6947 (N_6947,N_4833,N_4228);
nand U6948 (N_6948,N_5855,N_4187);
nand U6949 (N_6949,N_4376,N_5438);
nor U6950 (N_6950,N_5620,N_4091);
and U6951 (N_6951,N_4355,N_4220);
xnor U6952 (N_6952,N_4542,N_5153);
nand U6953 (N_6953,N_5227,N_5657);
and U6954 (N_6954,N_5986,N_4713);
nor U6955 (N_6955,N_4277,N_5199);
and U6956 (N_6956,N_4268,N_5499);
or U6957 (N_6957,N_4375,N_4211);
and U6958 (N_6958,N_5865,N_4147);
or U6959 (N_6959,N_4216,N_4966);
nand U6960 (N_6960,N_4703,N_4684);
and U6961 (N_6961,N_5726,N_5642);
and U6962 (N_6962,N_4536,N_4555);
and U6963 (N_6963,N_5295,N_4795);
and U6964 (N_6964,N_4351,N_4822);
or U6965 (N_6965,N_5721,N_4813);
and U6966 (N_6966,N_4012,N_4981);
nand U6967 (N_6967,N_5987,N_4353);
or U6968 (N_6968,N_4869,N_4274);
nor U6969 (N_6969,N_5348,N_5498);
nor U6970 (N_6970,N_5066,N_4386);
xor U6971 (N_6971,N_4926,N_5563);
and U6972 (N_6972,N_5437,N_5123);
nand U6973 (N_6973,N_5891,N_4721);
and U6974 (N_6974,N_4265,N_4067);
nand U6975 (N_6975,N_4367,N_4148);
nor U6976 (N_6976,N_5353,N_4552);
xor U6977 (N_6977,N_5795,N_4796);
nor U6978 (N_6978,N_5366,N_4343);
nand U6979 (N_6979,N_5667,N_4043);
xnor U6980 (N_6980,N_4848,N_4756);
or U6981 (N_6981,N_5306,N_4392);
or U6982 (N_6982,N_4871,N_5250);
or U6983 (N_6983,N_4234,N_5770);
nand U6984 (N_6984,N_4685,N_5509);
nor U6985 (N_6985,N_4260,N_4186);
or U6986 (N_6986,N_5626,N_5002);
nand U6987 (N_6987,N_4400,N_4550);
or U6988 (N_6988,N_4688,N_5304);
xnor U6989 (N_6989,N_4338,N_5634);
nor U6990 (N_6990,N_4167,N_5486);
and U6991 (N_6991,N_4411,N_4558);
or U6992 (N_6992,N_4119,N_5303);
xor U6993 (N_6993,N_4613,N_5268);
and U6994 (N_6994,N_5083,N_5872);
nor U6995 (N_6995,N_4466,N_5188);
and U6996 (N_6996,N_4727,N_5631);
nand U6997 (N_6997,N_4898,N_5409);
or U6998 (N_6998,N_5697,N_5400);
xor U6999 (N_6999,N_4775,N_5248);
and U7000 (N_7000,N_5235,N_5437);
nor U7001 (N_7001,N_5361,N_5088);
nor U7002 (N_7002,N_4881,N_4946);
or U7003 (N_7003,N_4057,N_4231);
nand U7004 (N_7004,N_5241,N_4709);
nand U7005 (N_7005,N_5437,N_5762);
and U7006 (N_7006,N_4636,N_4700);
nand U7007 (N_7007,N_4510,N_5357);
or U7008 (N_7008,N_5950,N_4619);
and U7009 (N_7009,N_5303,N_5795);
or U7010 (N_7010,N_4845,N_4186);
or U7011 (N_7011,N_5497,N_5839);
and U7012 (N_7012,N_5544,N_5158);
nor U7013 (N_7013,N_5864,N_4947);
or U7014 (N_7014,N_4374,N_5985);
nor U7015 (N_7015,N_4368,N_5066);
xor U7016 (N_7016,N_5375,N_5594);
nor U7017 (N_7017,N_5720,N_4964);
xor U7018 (N_7018,N_4082,N_5647);
nand U7019 (N_7019,N_5077,N_4332);
or U7020 (N_7020,N_5048,N_4584);
xor U7021 (N_7021,N_4918,N_4781);
nand U7022 (N_7022,N_5034,N_5338);
nand U7023 (N_7023,N_5203,N_5775);
and U7024 (N_7024,N_5004,N_5380);
or U7025 (N_7025,N_5132,N_4957);
or U7026 (N_7026,N_5760,N_5635);
and U7027 (N_7027,N_5332,N_5660);
xnor U7028 (N_7028,N_5190,N_5935);
nand U7029 (N_7029,N_5299,N_4116);
nor U7030 (N_7030,N_5496,N_4843);
and U7031 (N_7031,N_4388,N_4894);
and U7032 (N_7032,N_4367,N_5157);
nand U7033 (N_7033,N_5877,N_4595);
and U7034 (N_7034,N_4430,N_5631);
or U7035 (N_7035,N_4377,N_5650);
and U7036 (N_7036,N_4812,N_5625);
xnor U7037 (N_7037,N_4836,N_4422);
and U7038 (N_7038,N_4667,N_5498);
nand U7039 (N_7039,N_5189,N_5411);
nand U7040 (N_7040,N_4616,N_4012);
xnor U7041 (N_7041,N_5344,N_4937);
or U7042 (N_7042,N_4061,N_5455);
xor U7043 (N_7043,N_4145,N_5641);
nor U7044 (N_7044,N_5047,N_4946);
or U7045 (N_7045,N_5704,N_4876);
nand U7046 (N_7046,N_4718,N_4400);
nand U7047 (N_7047,N_5906,N_5013);
nand U7048 (N_7048,N_4429,N_5671);
and U7049 (N_7049,N_4950,N_5434);
and U7050 (N_7050,N_5211,N_5622);
or U7051 (N_7051,N_5596,N_4578);
or U7052 (N_7052,N_5841,N_4472);
xor U7053 (N_7053,N_5726,N_5930);
nor U7054 (N_7054,N_4134,N_4984);
or U7055 (N_7055,N_5277,N_4931);
xor U7056 (N_7056,N_5738,N_4172);
nor U7057 (N_7057,N_4496,N_5812);
nor U7058 (N_7058,N_5096,N_4233);
and U7059 (N_7059,N_5025,N_5512);
nand U7060 (N_7060,N_5439,N_4683);
nand U7061 (N_7061,N_4192,N_5388);
nand U7062 (N_7062,N_5464,N_5355);
or U7063 (N_7063,N_4630,N_5274);
xnor U7064 (N_7064,N_4144,N_4794);
xnor U7065 (N_7065,N_5179,N_4465);
and U7066 (N_7066,N_5504,N_5716);
xor U7067 (N_7067,N_4334,N_4513);
or U7068 (N_7068,N_5950,N_4732);
and U7069 (N_7069,N_4198,N_5959);
nor U7070 (N_7070,N_4990,N_5028);
nand U7071 (N_7071,N_4262,N_5496);
and U7072 (N_7072,N_5388,N_5622);
or U7073 (N_7073,N_4198,N_4843);
or U7074 (N_7074,N_5015,N_4428);
and U7075 (N_7075,N_4666,N_5452);
and U7076 (N_7076,N_5765,N_5350);
or U7077 (N_7077,N_5192,N_5439);
or U7078 (N_7078,N_5495,N_4608);
or U7079 (N_7079,N_5022,N_4771);
nor U7080 (N_7080,N_4424,N_4325);
or U7081 (N_7081,N_5089,N_5603);
nor U7082 (N_7082,N_4050,N_5551);
nor U7083 (N_7083,N_4403,N_4191);
xor U7084 (N_7084,N_5083,N_4943);
nor U7085 (N_7085,N_5830,N_5920);
xor U7086 (N_7086,N_4469,N_5766);
and U7087 (N_7087,N_5997,N_5336);
nor U7088 (N_7088,N_5230,N_4197);
nand U7089 (N_7089,N_4139,N_4440);
xnor U7090 (N_7090,N_5542,N_4513);
and U7091 (N_7091,N_4474,N_5355);
nand U7092 (N_7092,N_4481,N_5476);
and U7093 (N_7093,N_5453,N_5455);
xnor U7094 (N_7094,N_5263,N_4329);
and U7095 (N_7095,N_4924,N_5122);
nand U7096 (N_7096,N_5246,N_4432);
or U7097 (N_7097,N_4144,N_5525);
xor U7098 (N_7098,N_4901,N_4386);
xor U7099 (N_7099,N_4288,N_4313);
xor U7100 (N_7100,N_5750,N_5261);
xnor U7101 (N_7101,N_5714,N_5250);
xnor U7102 (N_7102,N_5931,N_5959);
or U7103 (N_7103,N_5111,N_4240);
nor U7104 (N_7104,N_4807,N_4126);
nand U7105 (N_7105,N_5468,N_4938);
or U7106 (N_7106,N_4960,N_5986);
nor U7107 (N_7107,N_5769,N_4201);
or U7108 (N_7108,N_4404,N_5017);
and U7109 (N_7109,N_5561,N_4112);
xor U7110 (N_7110,N_5788,N_5709);
nand U7111 (N_7111,N_4257,N_4450);
or U7112 (N_7112,N_5948,N_5757);
nand U7113 (N_7113,N_4225,N_5364);
nor U7114 (N_7114,N_4424,N_5895);
nand U7115 (N_7115,N_4243,N_5539);
xor U7116 (N_7116,N_4588,N_4758);
nor U7117 (N_7117,N_5993,N_4636);
nor U7118 (N_7118,N_5475,N_5878);
nor U7119 (N_7119,N_5636,N_5482);
nand U7120 (N_7120,N_5161,N_4050);
and U7121 (N_7121,N_4195,N_4793);
or U7122 (N_7122,N_5649,N_5852);
nand U7123 (N_7123,N_4839,N_5710);
xor U7124 (N_7124,N_5547,N_5156);
or U7125 (N_7125,N_4582,N_4882);
and U7126 (N_7126,N_5209,N_4806);
or U7127 (N_7127,N_5254,N_4050);
and U7128 (N_7128,N_5131,N_5915);
nand U7129 (N_7129,N_5993,N_4379);
and U7130 (N_7130,N_5297,N_5020);
xor U7131 (N_7131,N_4689,N_5933);
nor U7132 (N_7132,N_4947,N_4517);
nand U7133 (N_7133,N_4716,N_5171);
or U7134 (N_7134,N_5749,N_5935);
and U7135 (N_7135,N_5951,N_5054);
nor U7136 (N_7136,N_4639,N_5232);
or U7137 (N_7137,N_5744,N_5516);
or U7138 (N_7138,N_4314,N_4236);
and U7139 (N_7139,N_4812,N_5723);
nand U7140 (N_7140,N_5084,N_5143);
xor U7141 (N_7141,N_5253,N_4656);
or U7142 (N_7142,N_5597,N_5458);
nand U7143 (N_7143,N_4929,N_5981);
nand U7144 (N_7144,N_4589,N_5035);
xnor U7145 (N_7145,N_4245,N_4063);
xnor U7146 (N_7146,N_5088,N_5238);
nor U7147 (N_7147,N_4703,N_4957);
nor U7148 (N_7148,N_5513,N_5207);
nor U7149 (N_7149,N_4808,N_5191);
and U7150 (N_7150,N_4335,N_4243);
and U7151 (N_7151,N_5381,N_5860);
nor U7152 (N_7152,N_4482,N_4952);
nor U7153 (N_7153,N_4003,N_4539);
nor U7154 (N_7154,N_4848,N_4684);
nor U7155 (N_7155,N_4646,N_4109);
xnor U7156 (N_7156,N_4010,N_5446);
nand U7157 (N_7157,N_5042,N_5453);
and U7158 (N_7158,N_4408,N_4326);
xor U7159 (N_7159,N_5349,N_5302);
nor U7160 (N_7160,N_5069,N_5110);
xnor U7161 (N_7161,N_5457,N_4867);
or U7162 (N_7162,N_4617,N_5625);
xnor U7163 (N_7163,N_4595,N_4543);
nor U7164 (N_7164,N_4090,N_4858);
nand U7165 (N_7165,N_4310,N_4277);
and U7166 (N_7166,N_5617,N_4900);
or U7167 (N_7167,N_5711,N_4918);
xnor U7168 (N_7168,N_5699,N_4808);
nand U7169 (N_7169,N_5493,N_4606);
nor U7170 (N_7170,N_5633,N_4455);
xnor U7171 (N_7171,N_4175,N_4879);
xor U7172 (N_7172,N_5157,N_4741);
and U7173 (N_7173,N_5027,N_5159);
xor U7174 (N_7174,N_5034,N_4384);
nand U7175 (N_7175,N_5654,N_5543);
xor U7176 (N_7176,N_4513,N_5286);
or U7177 (N_7177,N_4004,N_5753);
or U7178 (N_7178,N_4174,N_5622);
xor U7179 (N_7179,N_4942,N_5387);
or U7180 (N_7180,N_4696,N_5682);
xnor U7181 (N_7181,N_5288,N_5882);
nor U7182 (N_7182,N_4336,N_5632);
nor U7183 (N_7183,N_4203,N_5603);
and U7184 (N_7184,N_5984,N_4300);
xnor U7185 (N_7185,N_4693,N_5321);
nor U7186 (N_7186,N_4753,N_5476);
nor U7187 (N_7187,N_5576,N_5694);
nand U7188 (N_7188,N_5360,N_5409);
nand U7189 (N_7189,N_4752,N_4722);
and U7190 (N_7190,N_5059,N_4550);
or U7191 (N_7191,N_4549,N_5544);
xor U7192 (N_7192,N_5082,N_5722);
xnor U7193 (N_7193,N_4425,N_5485);
nor U7194 (N_7194,N_4117,N_4436);
nor U7195 (N_7195,N_5777,N_4258);
nand U7196 (N_7196,N_5402,N_4333);
nor U7197 (N_7197,N_4891,N_5078);
nand U7198 (N_7198,N_4748,N_5348);
or U7199 (N_7199,N_5112,N_5576);
and U7200 (N_7200,N_5508,N_4744);
and U7201 (N_7201,N_4709,N_5548);
and U7202 (N_7202,N_4507,N_4171);
xor U7203 (N_7203,N_4548,N_4817);
or U7204 (N_7204,N_5709,N_4322);
xor U7205 (N_7205,N_4713,N_5835);
nor U7206 (N_7206,N_4829,N_5652);
xnor U7207 (N_7207,N_4300,N_4411);
nand U7208 (N_7208,N_4045,N_5079);
or U7209 (N_7209,N_4152,N_4261);
nor U7210 (N_7210,N_4215,N_4000);
nor U7211 (N_7211,N_4576,N_4852);
nand U7212 (N_7212,N_4553,N_5918);
nor U7213 (N_7213,N_5707,N_4394);
nand U7214 (N_7214,N_5032,N_5547);
nor U7215 (N_7215,N_5749,N_4525);
xor U7216 (N_7216,N_4115,N_4260);
nand U7217 (N_7217,N_4033,N_4394);
and U7218 (N_7218,N_5265,N_4150);
and U7219 (N_7219,N_4004,N_5108);
or U7220 (N_7220,N_5483,N_5883);
nor U7221 (N_7221,N_4704,N_5883);
nand U7222 (N_7222,N_4835,N_5908);
and U7223 (N_7223,N_5887,N_4491);
xor U7224 (N_7224,N_4689,N_5570);
and U7225 (N_7225,N_5809,N_5405);
nand U7226 (N_7226,N_4125,N_4515);
or U7227 (N_7227,N_5859,N_4041);
or U7228 (N_7228,N_5123,N_4510);
nor U7229 (N_7229,N_5000,N_5535);
or U7230 (N_7230,N_5355,N_4385);
or U7231 (N_7231,N_5026,N_4060);
and U7232 (N_7232,N_5276,N_5127);
nor U7233 (N_7233,N_4563,N_5707);
xnor U7234 (N_7234,N_4366,N_5986);
and U7235 (N_7235,N_4164,N_4783);
and U7236 (N_7236,N_5732,N_5136);
nand U7237 (N_7237,N_4158,N_4992);
and U7238 (N_7238,N_5780,N_4106);
and U7239 (N_7239,N_5917,N_5862);
or U7240 (N_7240,N_4956,N_4046);
or U7241 (N_7241,N_5504,N_5488);
and U7242 (N_7242,N_5225,N_5946);
xnor U7243 (N_7243,N_5816,N_5752);
nand U7244 (N_7244,N_4096,N_4155);
xor U7245 (N_7245,N_5301,N_5848);
nand U7246 (N_7246,N_4045,N_5340);
or U7247 (N_7247,N_4515,N_4143);
nor U7248 (N_7248,N_5688,N_4199);
nand U7249 (N_7249,N_5420,N_5031);
and U7250 (N_7250,N_5198,N_4520);
or U7251 (N_7251,N_4289,N_5125);
xor U7252 (N_7252,N_4242,N_4385);
or U7253 (N_7253,N_4210,N_4868);
xor U7254 (N_7254,N_4621,N_4421);
and U7255 (N_7255,N_4328,N_5959);
nand U7256 (N_7256,N_5819,N_5640);
or U7257 (N_7257,N_4679,N_5600);
nand U7258 (N_7258,N_4212,N_5608);
nor U7259 (N_7259,N_4365,N_4749);
nor U7260 (N_7260,N_5293,N_4296);
and U7261 (N_7261,N_5615,N_4447);
nand U7262 (N_7262,N_4532,N_4318);
nand U7263 (N_7263,N_5727,N_5436);
xor U7264 (N_7264,N_4981,N_4880);
nand U7265 (N_7265,N_5949,N_5576);
and U7266 (N_7266,N_4139,N_5920);
nand U7267 (N_7267,N_4062,N_4928);
xnor U7268 (N_7268,N_4068,N_4318);
xnor U7269 (N_7269,N_4303,N_5964);
or U7270 (N_7270,N_5532,N_5149);
and U7271 (N_7271,N_4938,N_5096);
and U7272 (N_7272,N_4936,N_5133);
nor U7273 (N_7273,N_4075,N_4901);
and U7274 (N_7274,N_5784,N_4151);
nand U7275 (N_7275,N_5856,N_5176);
nand U7276 (N_7276,N_4255,N_4098);
or U7277 (N_7277,N_5772,N_4535);
or U7278 (N_7278,N_4150,N_5842);
and U7279 (N_7279,N_4580,N_5624);
nor U7280 (N_7280,N_5675,N_4682);
nand U7281 (N_7281,N_5835,N_5673);
nand U7282 (N_7282,N_4091,N_4566);
xnor U7283 (N_7283,N_4986,N_4057);
nor U7284 (N_7284,N_5199,N_5715);
and U7285 (N_7285,N_5716,N_5510);
or U7286 (N_7286,N_4577,N_4010);
and U7287 (N_7287,N_4396,N_5251);
or U7288 (N_7288,N_5481,N_4029);
nor U7289 (N_7289,N_5894,N_4831);
nand U7290 (N_7290,N_4570,N_5056);
and U7291 (N_7291,N_5462,N_4458);
and U7292 (N_7292,N_5522,N_5458);
and U7293 (N_7293,N_5950,N_5998);
and U7294 (N_7294,N_4127,N_5706);
and U7295 (N_7295,N_4872,N_5714);
nor U7296 (N_7296,N_5371,N_4160);
and U7297 (N_7297,N_5465,N_5688);
xnor U7298 (N_7298,N_4781,N_4476);
nand U7299 (N_7299,N_4886,N_5097);
nor U7300 (N_7300,N_4374,N_4674);
nand U7301 (N_7301,N_5521,N_5183);
nand U7302 (N_7302,N_4419,N_5069);
nand U7303 (N_7303,N_4528,N_4202);
nor U7304 (N_7304,N_4185,N_4920);
and U7305 (N_7305,N_4604,N_5104);
nor U7306 (N_7306,N_4114,N_4169);
and U7307 (N_7307,N_5627,N_5056);
nor U7308 (N_7308,N_5742,N_4421);
nand U7309 (N_7309,N_5650,N_4730);
nor U7310 (N_7310,N_4756,N_4813);
or U7311 (N_7311,N_4493,N_4953);
xor U7312 (N_7312,N_4854,N_5892);
and U7313 (N_7313,N_5073,N_5510);
nand U7314 (N_7314,N_4941,N_4774);
nor U7315 (N_7315,N_5286,N_5004);
xnor U7316 (N_7316,N_4849,N_5730);
xnor U7317 (N_7317,N_5558,N_4532);
and U7318 (N_7318,N_5807,N_4453);
nand U7319 (N_7319,N_5745,N_5642);
nor U7320 (N_7320,N_4688,N_4400);
nor U7321 (N_7321,N_4340,N_5610);
and U7322 (N_7322,N_4318,N_5313);
xor U7323 (N_7323,N_5014,N_4901);
or U7324 (N_7324,N_5913,N_4206);
nand U7325 (N_7325,N_5020,N_5468);
or U7326 (N_7326,N_5792,N_4182);
xnor U7327 (N_7327,N_4572,N_5226);
nand U7328 (N_7328,N_5500,N_5396);
or U7329 (N_7329,N_4867,N_5221);
or U7330 (N_7330,N_5283,N_5176);
nor U7331 (N_7331,N_5084,N_5597);
or U7332 (N_7332,N_4160,N_5847);
nand U7333 (N_7333,N_4328,N_4405);
nor U7334 (N_7334,N_4591,N_5436);
and U7335 (N_7335,N_4819,N_4379);
nor U7336 (N_7336,N_4711,N_4486);
or U7337 (N_7337,N_5666,N_5495);
and U7338 (N_7338,N_5163,N_4556);
nand U7339 (N_7339,N_4274,N_5006);
nand U7340 (N_7340,N_5294,N_5703);
nor U7341 (N_7341,N_4013,N_4329);
or U7342 (N_7342,N_4226,N_4954);
or U7343 (N_7343,N_4749,N_5060);
or U7344 (N_7344,N_5512,N_4179);
xor U7345 (N_7345,N_4416,N_5283);
nor U7346 (N_7346,N_5544,N_4325);
nor U7347 (N_7347,N_4658,N_5772);
or U7348 (N_7348,N_5890,N_5392);
or U7349 (N_7349,N_4417,N_5056);
xnor U7350 (N_7350,N_5966,N_4726);
or U7351 (N_7351,N_4308,N_4963);
and U7352 (N_7352,N_5696,N_5112);
nor U7353 (N_7353,N_4870,N_5962);
xnor U7354 (N_7354,N_4078,N_4772);
or U7355 (N_7355,N_5178,N_4135);
and U7356 (N_7356,N_5794,N_4389);
or U7357 (N_7357,N_5959,N_5684);
and U7358 (N_7358,N_5644,N_4125);
xnor U7359 (N_7359,N_4727,N_4469);
nor U7360 (N_7360,N_4999,N_4460);
or U7361 (N_7361,N_5252,N_5333);
or U7362 (N_7362,N_4750,N_5952);
and U7363 (N_7363,N_4568,N_5433);
xnor U7364 (N_7364,N_5556,N_4308);
or U7365 (N_7365,N_5804,N_4124);
nor U7366 (N_7366,N_5213,N_5937);
xor U7367 (N_7367,N_5657,N_4352);
xor U7368 (N_7368,N_5926,N_4166);
xnor U7369 (N_7369,N_5954,N_4693);
or U7370 (N_7370,N_5055,N_5296);
nand U7371 (N_7371,N_4437,N_5029);
and U7372 (N_7372,N_4450,N_5827);
or U7373 (N_7373,N_5514,N_5630);
xor U7374 (N_7374,N_5293,N_5250);
and U7375 (N_7375,N_5503,N_4275);
xnor U7376 (N_7376,N_4655,N_4387);
or U7377 (N_7377,N_5620,N_4867);
xor U7378 (N_7378,N_5331,N_5487);
nand U7379 (N_7379,N_5963,N_5011);
nor U7380 (N_7380,N_5095,N_5366);
nor U7381 (N_7381,N_5822,N_4667);
or U7382 (N_7382,N_5731,N_5283);
nor U7383 (N_7383,N_4234,N_5546);
xnor U7384 (N_7384,N_4649,N_5606);
xor U7385 (N_7385,N_4513,N_5505);
nor U7386 (N_7386,N_5717,N_4750);
or U7387 (N_7387,N_4197,N_4683);
and U7388 (N_7388,N_5634,N_5541);
nor U7389 (N_7389,N_4247,N_5172);
or U7390 (N_7390,N_5084,N_5135);
xor U7391 (N_7391,N_4728,N_5380);
xor U7392 (N_7392,N_5193,N_5471);
nor U7393 (N_7393,N_5915,N_4085);
nand U7394 (N_7394,N_5490,N_5866);
and U7395 (N_7395,N_5398,N_4733);
nor U7396 (N_7396,N_4759,N_4143);
nor U7397 (N_7397,N_5127,N_4447);
xor U7398 (N_7398,N_4972,N_5325);
and U7399 (N_7399,N_5472,N_4997);
xor U7400 (N_7400,N_5706,N_5713);
xor U7401 (N_7401,N_5468,N_4029);
or U7402 (N_7402,N_5377,N_5654);
nand U7403 (N_7403,N_5610,N_5912);
nand U7404 (N_7404,N_4073,N_5949);
xor U7405 (N_7405,N_4420,N_4409);
and U7406 (N_7406,N_5173,N_5971);
nor U7407 (N_7407,N_4375,N_5441);
nand U7408 (N_7408,N_4481,N_5804);
and U7409 (N_7409,N_5013,N_5860);
nor U7410 (N_7410,N_5439,N_5523);
or U7411 (N_7411,N_4774,N_4218);
and U7412 (N_7412,N_4864,N_5069);
nand U7413 (N_7413,N_5691,N_4248);
or U7414 (N_7414,N_4802,N_5007);
or U7415 (N_7415,N_4458,N_4580);
nand U7416 (N_7416,N_4678,N_4398);
or U7417 (N_7417,N_4045,N_5322);
xnor U7418 (N_7418,N_5135,N_5960);
nand U7419 (N_7419,N_4309,N_4596);
nand U7420 (N_7420,N_4000,N_4605);
or U7421 (N_7421,N_5136,N_5626);
and U7422 (N_7422,N_4044,N_4924);
nand U7423 (N_7423,N_4141,N_5456);
or U7424 (N_7424,N_4306,N_4193);
nor U7425 (N_7425,N_4857,N_4493);
and U7426 (N_7426,N_5698,N_4004);
or U7427 (N_7427,N_4483,N_5243);
nor U7428 (N_7428,N_4104,N_4044);
nand U7429 (N_7429,N_5884,N_4225);
xor U7430 (N_7430,N_4720,N_5084);
nor U7431 (N_7431,N_5627,N_4533);
nand U7432 (N_7432,N_5742,N_4128);
xnor U7433 (N_7433,N_5818,N_5333);
or U7434 (N_7434,N_4262,N_4832);
xor U7435 (N_7435,N_5510,N_5580);
and U7436 (N_7436,N_5834,N_4731);
nor U7437 (N_7437,N_5446,N_4229);
or U7438 (N_7438,N_4205,N_5927);
nor U7439 (N_7439,N_4063,N_4733);
nor U7440 (N_7440,N_4144,N_4007);
or U7441 (N_7441,N_4323,N_5447);
and U7442 (N_7442,N_5942,N_5601);
and U7443 (N_7443,N_4270,N_4019);
xor U7444 (N_7444,N_5101,N_4482);
nand U7445 (N_7445,N_4518,N_5314);
or U7446 (N_7446,N_5404,N_5382);
xor U7447 (N_7447,N_4584,N_5898);
nand U7448 (N_7448,N_5226,N_5054);
or U7449 (N_7449,N_5539,N_4165);
xor U7450 (N_7450,N_4088,N_5326);
nor U7451 (N_7451,N_4057,N_4228);
nand U7452 (N_7452,N_4349,N_4683);
and U7453 (N_7453,N_4039,N_5504);
or U7454 (N_7454,N_4613,N_5421);
nor U7455 (N_7455,N_5135,N_5047);
nand U7456 (N_7456,N_4260,N_5465);
nand U7457 (N_7457,N_4030,N_5813);
xnor U7458 (N_7458,N_5031,N_5530);
and U7459 (N_7459,N_4513,N_4564);
and U7460 (N_7460,N_5512,N_4009);
or U7461 (N_7461,N_4196,N_4763);
xor U7462 (N_7462,N_5776,N_5346);
nand U7463 (N_7463,N_4941,N_5137);
and U7464 (N_7464,N_5702,N_5044);
or U7465 (N_7465,N_5046,N_4287);
xnor U7466 (N_7466,N_4217,N_5319);
nor U7467 (N_7467,N_4782,N_4674);
or U7468 (N_7468,N_4838,N_5568);
nand U7469 (N_7469,N_5966,N_5759);
xnor U7470 (N_7470,N_5826,N_4415);
or U7471 (N_7471,N_4396,N_5289);
or U7472 (N_7472,N_4174,N_5577);
nor U7473 (N_7473,N_5417,N_5646);
nand U7474 (N_7474,N_5512,N_4677);
nor U7475 (N_7475,N_4885,N_4008);
nand U7476 (N_7476,N_4395,N_4068);
xnor U7477 (N_7477,N_4164,N_4455);
nand U7478 (N_7478,N_4167,N_4170);
nor U7479 (N_7479,N_5919,N_5410);
nand U7480 (N_7480,N_4295,N_4824);
nor U7481 (N_7481,N_4964,N_5080);
or U7482 (N_7482,N_4023,N_4717);
xnor U7483 (N_7483,N_5825,N_5500);
or U7484 (N_7484,N_4276,N_4916);
xnor U7485 (N_7485,N_4056,N_5479);
nand U7486 (N_7486,N_4906,N_5138);
nor U7487 (N_7487,N_4647,N_4942);
or U7488 (N_7488,N_4645,N_4559);
and U7489 (N_7489,N_4983,N_4536);
nand U7490 (N_7490,N_5143,N_4663);
nand U7491 (N_7491,N_4356,N_5917);
nor U7492 (N_7492,N_4523,N_5960);
xnor U7493 (N_7493,N_5575,N_4557);
and U7494 (N_7494,N_4857,N_5962);
nand U7495 (N_7495,N_5872,N_4053);
and U7496 (N_7496,N_5719,N_4579);
and U7497 (N_7497,N_4023,N_4726);
xnor U7498 (N_7498,N_5099,N_4073);
xor U7499 (N_7499,N_4436,N_5195);
nor U7500 (N_7500,N_4273,N_4743);
and U7501 (N_7501,N_4006,N_4108);
xnor U7502 (N_7502,N_4444,N_5295);
or U7503 (N_7503,N_5401,N_5146);
xor U7504 (N_7504,N_5682,N_5992);
or U7505 (N_7505,N_5062,N_4983);
xor U7506 (N_7506,N_5908,N_5676);
nor U7507 (N_7507,N_5951,N_4903);
or U7508 (N_7508,N_5332,N_4458);
and U7509 (N_7509,N_5350,N_4250);
nand U7510 (N_7510,N_5966,N_4801);
nand U7511 (N_7511,N_4939,N_5991);
or U7512 (N_7512,N_4101,N_5760);
nand U7513 (N_7513,N_4598,N_5102);
nor U7514 (N_7514,N_4998,N_5894);
and U7515 (N_7515,N_5049,N_5773);
nand U7516 (N_7516,N_5843,N_5111);
and U7517 (N_7517,N_4468,N_5075);
nand U7518 (N_7518,N_4535,N_4534);
or U7519 (N_7519,N_4005,N_4179);
xnor U7520 (N_7520,N_5033,N_4205);
nand U7521 (N_7521,N_5489,N_5756);
xor U7522 (N_7522,N_5657,N_5221);
nor U7523 (N_7523,N_5637,N_5972);
nor U7524 (N_7524,N_5542,N_4359);
and U7525 (N_7525,N_4009,N_4753);
or U7526 (N_7526,N_4922,N_5565);
nor U7527 (N_7527,N_5830,N_5024);
nor U7528 (N_7528,N_4871,N_4177);
xnor U7529 (N_7529,N_4635,N_4367);
or U7530 (N_7530,N_5074,N_5678);
or U7531 (N_7531,N_5606,N_4224);
xnor U7532 (N_7532,N_5859,N_4869);
xor U7533 (N_7533,N_4784,N_5892);
nand U7534 (N_7534,N_5860,N_4054);
xor U7535 (N_7535,N_5304,N_5041);
and U7536 (N_7536,N_4071,N_5990);
nor U7537 (N_7537,N_5304,N_4740);
nor U7538 (N_7538,N_5902,N_4669);
xor U7539 (N_7539,N_5474,N_5329);
nor U7540 (N_7540,N_5598,N_4101);
nor U7541 (N_7541,N_5946,N_4015);
nand U7542 (N_7542,N_5843,N_5707);
or U7543 (N_7543,N_5674,N_5809);
or U7544 (N_7544,N_5933,N_4328);
and U7545 (N_7545,N_5558,N_4935);
xor U7546 (N_7546,N_4199,N_5993);
nor U7547 (N_7547,N_4724,N_4637);
nand U7548 (N_7548,N_5025,N_5528);
nand U7549 (N_7549,N_5566,N_4412);
or U7550 (N_7550,N_5415,N_4454);
or U7551 (N_7551,N_5467,N_4728);
nor U7552 (N_7552,N_5376,N_5735);
and U7553 (N_7553,N_4389,N_5334);
or U7554 (N_7554,N_5956,N_5871);
nor U7555 (N_7555,N_4682,N_5526);
and U7556 (N_7556,N_5184,N_4175);
xnor U7557 (N_7557,N_5707,N_5940);
xnor U7558 (N_7558,N_4727,N_4857);
nand U7559 (N_7559,N_4394,N_4498);
or U7560 (N_7560,N_5699,N_5506);
and U7561 (N_7561,N_4927,N_4218);
nor U7562 (N_7562,N_5244,N_5190);
nor U7563 (N_7563,N_4649,N_5437);
xnor U7564 (N_7564,N_4525,N_5988);
xor U7565 (N_7565,N_4507,N_5998);
nand U7566 (N_7566,N_4281,N_4108);
nor U7567 (N_7567,N_4775,N_4884);
nand U7568 (N_7568,N_4373,N_4771);
or U7569 (N_7569,N_4677,N_4788);
and U7570 (N_7570,N_4709,N_5615);
or U7571 (N_7571,N_4433,N_5569);
or U7572 (N_7572,N_4637,N_5535);
nor U7573 (N_7573,N_5185,N_5611);
or U7574 (N_7574,N_5597,N_5738);
xnor U7575 (N_7575,N_4576,N_5526);
xor U7576 (N_7576,N_5988,N_4660);
xor U7577 (N_7577,N_4406,N_5441);
xor U7578 (N_7578,N_4510,N_5184);
nand U7579 (N_7579,N_4774,N_4805);
or U7580 (N_7580,N_4500,N_4907);
nor U7581 (N_7581,N_5487,N_4800);
xor U7582 (N_7582,N_4694,N_4461);
xor U7583 (N_7583,N_4551,N_4158);
xor U7584 (N_7584,N_4197,N_5581);
xnor U7585 (N_7585,N_5240,N_4416);
or U7586 (N_7586,N_5203,N_5880);
or U7587 (N_7587,N_4633,N_5457);
nor U7588 (N_7588,N_4342,N_5451);
nor U7589 (N_7589,N_5979,N_4553);
and U7590 (N_7590,N_4386,N_5568);
and U7591 (N_7591,N_5771,N_5343);
nor U7592 (N_7592,N_4405,N_5042);
and U7593 (N_7593,N_5923,N_5603);
or U7594 (N_7594,N_5539,N_5970);
nor U7595 (N_7595,N_4904,N_5533);
nor U7596 (N_7596,N_4658,N_5166);
and U7597 (N_7597,N_5321,N_4294);
nor U7598 (N_7598,N_4933,N_5828);
nor U7599 (N_7599,N_4510,N_5616);
nor U7600 (N_7600,N_4383,N_4115);
and U7601 (N_7601,N_5344,N_4550);
xnor U7602 (N_7602,N_5601,N_5616);
and U7603 (N_7603,N_5144,N_5247);
xnor U7604 (N_7604,N_4903,N_5867);
xor U7605 (N_7605,N_5680,N_4687);
xnor U7606 (N_7606,N_4364,N_5102);
xnor U7607 (N_7607,N_4845,N_4863);
and U7608 (N_7608,N_4696,N_5217);
nor U7609 (N_7609,N_4684,N_5553);
and U7610 (N_7610,N_5353,N_5524);
and U7611 (N_7611,N_4879,N_5296);
xor U7612 (N_7612,N_5812,N_5682);
nand U7613 (N_7613,N_5583,N_4564);
and U7614 (N_7614,N_5720,N_5053);
nor U7615 (N_7615,N_4437,N_5997);
and U7616 (N_7616,N_5109,N_5603);
nor U7617 (N_7617,N_5499,N_4565);
nor U7618 (N_7618,N_4528,N_4070);
xor U7619 (N_7619,N_4781,N_5899);
nand U7620 (N_7620,N_4095,N_4739);
and U7621 (N_7621,N_4127,N_4025);
xor U7622 (N_7622,N_4215,N_4471);
nand U7623 (N_7623,N_4417,N_4507);
nand U7624 (N_7624,N_5824,N_4007);
or U7625 (N_7625,N_4241,N_4125);
nand U7626 (N_7626,N_4591,N_5831);
nand U7627 (N_7627,N_4535,N_5333);
nand U7628 (N_7628,N_4193,N_5119);
nand U7629 (N_7629,N_5268,N_5417);
or U7630 (N_7630,N_4451,N_5782);
xor U7631 (N_7631,N_4846,N_4706);
xor U7632 (N_7632,N_5830,N_5345);
xor U7633 (N_7633,N_5344,N_4222);
xor U7634 (N_7634,N_4408,N_4509);
nand U7635 (N_7635,N_5968,N_4145);
or U7636 (N_7636,N_4894,N_4301);
and U7637 (N_7637,N_5822,N_5420);
and U7638 (N_7638,N_5001,N_4769);
nand U7639 (N_7639,N_4269,N_5773);
or U7640 (N_7640,N_4030,N_5737);
nand U7641 (N_7641,N_5299,N_5694);
or U7642 (N_7642,N_4791,N_5285);
and U7643 (N_7643,N_5343,N_4096);
nor U7644 (N_7644,N_4873,N_4882);
or U7645 (N_7645,N_5735,N_4294);
and U7646 (N_7646,N_5069,N_4936);
xor U7647 (N_7647,N_4455,N_4413);
or U7648 (N_7648,N_5059,N_4684);
or U7649 (N_7649,N_5817,N_4301);
and U7650 (N_7650,N_5409,N_4811);
nand U7651 (N_7651,N_4778,N_5152);
or U7652 (N_7652,N_5294,N_5545);
nand U7653 (N_7653,N_4250,N_5934);
xor U7654 (N_7654,N_4996,N_5912);
and U7655 (N_7655,N_5016,N_4216);
nand U7656 (N_7656,N_4736,N_5348);
and U7657 (N_7657,N_4790,N_4536);
or U7658 (N_7658,N_4802,N_5735);
or U7659 (N_7659,N_5307,N_4230);
nor U7660 (N_7660,N_4210,N_4261);
and U7661 (N_7661,N_5196,N_4082);
nor U7662 (N_7662,N_4974,N_4251);
nor U7663 (N_7663,N_4704,N_4608);
and U7664 (N_7664,N_5106,N_4053);
nor U7665 (N_7665,N_4868,N_5467);
or U7666 (N_7666,N_4645,N_5376);
nor U7667 (N_7667,N_4046,N_5856);
or U7668 (N_7668,N_5995,N_4700);
nor U7669 (N_7669,N_4905,N_4593);
xor U7670 (N_7670,N_5680,N_4298);
nand U7671 (N_7671,N_5682,N_5371);
and U7672 (N_7672,N_4693,N_4657);
nor U7673 (N_7673,N_5271,N_5640);
nand U7674 (N_7674,N_4225,N_5055);
or U7675 (N_7675,N_4257,N_4017);
nand U7676 (N_7676,N_5151,N_5429);
nor U7677 (N_7677,N_4413,N_5592);
and U7678 (N_7678,N_4836,N_4105);
xor U7679 (N_7679,N_4007,N_5159);
or U7680 (N_7680,N_5061,N_4422);
xnor U7681 (N_7681,N_5188,N_4503);
and U7682 (N_7682,N_4313,N_4612);
nor U7683 (N_7683,N_4573,N_5499);
nand U7684 (N_7684,N_5391,N_4872);
nor U7685 (N_7685,N_4867,N_4774);
and U7686 (N_7686,N_5415,N_5533);
or U7687 (N_7687,N_4521,N_5980);
nor U7688 (N_7688,N_4832,N_5934);
xor U7689 (N_7689,N_4241,N_4840);
and U7690 (N_7690,N_5939,N_5670);
or U7691 (N_7691,N_5648,N_5093);
nand U7692 (N_7692,N_5687,N_4361);
nand U7693 (N_7693,N_5131,N_5314);
nor U7694 (N_7694,N_4633,N_4868);
nor U7695 (N_7695,N_4127,N_5917);
and U7696 (N_7696,N_4380,N_4179);
nand U7697 (N_7697,N_4619,N_5184);
nor U7698 (N_7698,N_4169,N_5149);
and U7699 (N_7699,N_5603,N_4086);
xor U7700 (N_7700,N_4416,N_5364);
or U7701 (N_7701,N_5941,N_4196);
xor U7702 (N_7702,N_4705,N_4300);
and U7703 (N_7703,N_4577,N_4325);
nand U7704 (N_7704,N_5346,N_4734);
nand U7705 (N_7705,N_5658,N_4017);
and U7706 (N_7706,N_4041,N_5148);
xor U7707 (N_7707,N_5078,N_4545);
and U7708 (N_7708,N_4880,N_5589);
and U7709 (N_7709,N_5126,N_4055);
or U7710 (N_7710,N_5610,N_5840);
xnor U7711 (N_7711,N_5493,N_4500);
nor U7712 (N_7712,N_5771,N_5839);
and U7713 (N_7713,N_4623,N_4899);
nor U7714 (N_7714,N_5440,N_4501);
and U7715 (N_7715,N_4314,N_5832);
and U7716 (N_7716,N_5974,N_5783);
nand U7717 (N_7717,N_5882,N_5941);
nor U7718 (N_7718,N_5568,N_4102);
and U7719 (N_7719,N_5761,N_4529);
nand U7720 (N_7720,N_5307,N_5982);
and U7721 (N_7721,N_4040,N_4919);
nand U7722 (N_7722,N_5309,N_4284);
nand U7723 (N_7723,N_4796,N_4242);
and U7724 (N_7724,N_4975,N_5974);
nor U7725 (N_7725,N_4845,N_4987);
nand U7726 (N_7726,N_5632,N_5577);
xnor U7727 (N_7727,N_4910,N_4856);
nand U7728 (N_7728,N_4045,N_4246);
and U7729 (N_7729,N_4304,N_5678);
nor U7730 (N_7730,N_4935,N_4238);
and U7731 (N_7731,N_5514,N_5153);
nor U7732 (N_7732,N_4560,N_5578);
and U7733 (N_7733,N_5652,N_4554);
xnor U7734 (N_7734,N_5443,N_5821);
and U7735 (N_7735,N_4663,N_4213);
or U7736 (N_7736,N_4708,N_4590);
xnor U7737 (N_7737,N_5960,N_5620);
nand U7738 (N_7738,N_5187,N_4035);
nor U7739 (N_7739,N_4764,N_4193);
xnor U7740 (N_7740,N_4406,N_4014);
xor U7741 (N_7741,N_4528,N_4608);
xnor U7742 (N_7742,N_5297,N_5921);
and U7743 (N_7743,N_4660,N_5851);
nand U7744 (N_7744,N_5407,N_4113);
or U7745 (N_7745,N_4661,N_4691);
xnor U7746 (N_7746,N_4267,N_5170);
xor U7747 (N_7747,N_5187,N_5203);
nand U7748 (N_7748,N_4310,N_5622);
xnor U7749 (N_7749,N_4472,N_4932);
and U7750 (N_7750,N_5652,N_5935);
and U7751 (N_7751,N_5405,N_4198);
xor U7752 (N_7752,N_4837,N_4604);
nand U7753 (N_7753,N_5012,N_5022);
and U7754 (N_7754,N_4725,N_4830);
nand U7755 (N_7755,N_5406,N_5954);
nand U7756 (N_7756,N_5550,N_4229);
nand U7757 (N_7757,N_5469,N_4630);
and U7758 (N_7758,N_5165,N_4699);
nor U7759 (N_7759,N_5890,N_4931);
xnor U7760 (N_7760,N_4958,N_4752);
or U7761 (N_7761,N_4356,N_4355);
nor U7762 (N_7762,N_5312,N_4910);
xor U7763 (N_7763,N_4416,N_4389);
nand U7764 (N_7764,N_4400,N_4456);
nand U7765 (N_7765,N_5745,N_5809);
nor U7766 (N_7766,N_4956,N_5129);
or U7767 (N_7767,N_4342,N_5348);
and U7768 (N_7768,N_4772,N_5762);
or U7769 (N_7769,N_5971,N_4973);
nand U7770 (N_7770,N_5177,N_5950);
nand U7771 (N_7771,N_5969,N_5528);
or U7772 (N_7772,N_5099,N_5682);
and U7773 (N_7773,N_4611,N_5682);
nor U7774 (N_7774,N_4038,N_4564);
and U7775 (N_7775,N_4149,N_4767);
and U7776 (N_7776,N_5337,N_4032);
or U7777 (N_7777,N_4466,N_5294);
and U7778 (N_7778,N_5511,N_5592);
nand U7779 (N_7779,N_4953,N_4289);
nor U7780 (N_7780,N_5462,N_4486);
nor U7781 (N_7781,N_4311,N_5432);
xnor U7782 (N_7782,N_5959,N_5511);
or U7783 (N_7783,N_5236,N_5888);
nor U7784 (N_7784,N_4215,N_4596);
xor U7785 (N_7785,N_5602,N_5364);
nor U7786 (N_7786,N_5128,N_4168);
and U7787 (N_7787,N_5114,N_4604);
xor U7788 (N_7788,N_5976,N_4501);
xnor U7789 (N_7789,N_5375,N_5875);
xnor U7790 (N_7790,N_4515,N_5960);
nand U7791 (N_7791,N_4516,N_5569);
nand U7792 (N_7792,N_4614,N_4947);
or U7793 (N_7793,N_4907,N_5272);
or U7794 (N_7794,N_5734,N_4049);
and U7795 (N_7795,N_5377,N_4914);
and U7796 (N_7796,N_5759,N_5168);
xnor U7797 (N_7797,N_4935,N_5738);
or U7798 (N_7798,N_5131,N_5536);
nand U7799 (N_7799,N_4712,N_5850);
xnor U7800 (N_7800,N_5967,N_4512);
xnor U7801 (N_7801,N_4928,N_4938);
nor U7802 (N_7802,N_5852,N_4449);
or U7803 (N_7803,N_5332,N_4984);
xor U7804 (N_7804,N_5750,N_5529);
and U7805 (N_7805,N_4593,N_5884);
nand U7806 (N_7806,N_5566,N_4688);
and U7807 (N_7807,N_5740,N_5447);
nand U7808 (N_7808,N_4989,N_5707);
or U7809 (N_7809,N_4234,N_5399);
nand U7810 (N_7810,N_4934,N_5435);
or U7811 (N_7811,N_5644,N_4839);
nor U7812 (N_7812,N_5321,N_5593);
nand U7813 (N_7813,N_4673,N_5337);
nand U7814 (N_7814,N_4799,N_4717);
or U7815 (N_7815,N_5729,N_4256);
and U7816 (N_7816,N_4596,N_5408);
nor U7817 (N_7817,N_5315,N_5856);
nand U7818 (N_7818,N_4592,N_4410);
and U7819 (N_7819,N_4602,N_4408);
or U7820 (N_7820,N_4340,N_5163);
or U7821 (N_7821,N_5057,N_4616);
or U7822 (N_7822,N_5134,N_4057);
xnor U7823 (N_7823,N_4521,N_5731);
or U7824 (N_7824,N_5650,N_4841);
nor U7825 (N_7825,N_5377,N_5303);
nor U7826 (N_7826,N_4977,N_4860);
xnor U7827 (N_7827,N_4270,N_5881);
and U7828 (N_7828,N_5644,N_4315);
and U7829 (N_7829,N_4190,N_5293);
and U7830 (N_7830,N_5892,N_5270);
xnor U7831 (N_7831,N_5589,N_4954);
xnor U7832 (N_7832,N_5569,N_5007);
nor U7833 (N_7833,N_5067,N_4882);
nor U7834 (N_7834,N_4697,N_4262);
xnor U7835 (N_7835,N_4134,N_4372);
and U7836 (N_7836,N_4130,N_5462);
nand U7837 (N_7837,N_5400,N_4360);
and U7838 (N_7838,N_4334,N_5503);
nor U7839 (N_7839,N_5156,N_5002);
nor U7840 (N_7840,N_5413,N_5415);
xnor U7841 (N_7841,N_5665,N_5922);
and U7842 (N_7842,N_5662,N_5876);
or U7843 (N_7843,N_4115,N_5350);
xnor U7844 (N_7844,N_5625,N_4040);
or U7845 (N_7845,N_4685,N_5363);
or U7846 (N_7846,N_4854,N_5962);
xnor U7847 (N_7847,N_4217,N_4598);
or U7848 (N_7848,N_4336,N_4122);
nand U7849 (N_7849,N_4410,N_4300);
and U7850 (N_7850,N_4641,N_4695);
nand U7851 (N_7851,N_5329,N_5523);
xnor U7852 (N_7852,N_4894,N_5024);
nor U7853 (N_7853,N_4641,N_5999);
or U7854 (N_7854,N_5203,N_5961);
nand U7855 (N_7855,N_5266,N_4652);
nor U7856 (N_7856,N_5100,N_5141);
and U7857 (N_7857,N_4732,N_5860);
or U7858 (N_7858,N_4425,N_5005);
xnor U7859 (N_7859,N_5238,N_5361);
and U7860 (N_7860,N_5317,N_4565);
nor U7861 (N_7861,N_4168,N_5213);
nor U7862 (N_7862,N_5352,N_5358);
and U7863 (N_7863,N_4984,N_4160);
nor U7864 (N_7864,N_4341,N_5381);
xor U7865 (N_7865,N_4058,N_4531);
and U7866 (N_7866,N_4274,N_4079);
nand U7867 (N_7867,N_4114,N_4979);
or U7868 (N_7868,N_5787,N_5564);
nor U7869 (N_7869,N_4173,N_4817);
or U7870 (N_7870,N_4387,N_4019);
and U7871 (N_7871,N_4306,N_5446);
or U7872 (N_7872,N_4473,N_5626);
or U7873 (N_7873,N_4252,N_4060);
or U7874 (N_7874,N_4850,N_5077);
nor U7875 (N_7875,N_5694,N_4700);
and U7876 (N_7876,N_5809,N_4084);
nor U7877 (N_7877,N_4043,N_5730);
nor U7878 (N_7878,N_5351,N_4064);
and U7879 (N_7879,N_4242,N_5519);
nor U7880 (N_7880,N_4646,N_5822);
and U7881 (N_7881,N_5325,N_5207);
or U7882 (N_7882,N_5319,N_4728);
nor U7883 (N_7883,N_5749,N_4390);
nand U7884 (N_7884,N_4079,N_5085);
or U7885 (N_7885,N_5914,N_5009);
and U7886 (N_7886,N_5941,N_5282);
nor U7887 (N_7887,N_5175,N_5718);
and U7888 (N_7888,N_4262,N_4541);
nor U7889 (N_7889,N_4098,N_4838);
or U7890 (N_7890,N_4023,N_5985);
and U7891 (N_7891,N_4330,N_5020);
and U7892 (N_7892,N_5255,N_4947);
nor U7893 (N_7893,N_4343,N_5497);
or U7894 (N_7894,N_4948,N_4949);
nor U7895 (N_7895,N_5532,N_4456);
xnor U7896 (N_7896,N_4154,N_4138);
or U7897 (N_7897,N_4558,N_4640);
or U7898 (N_7898,N_5557,N_4452);
nand U7899 (N_7899,N_5229,N_5432);
xor U7900 (N_7900,N_4988,N_4859);
nand U7901 (N_7901,N_4274,N_5061);
and U7902 (N_7902,N_5279,N_5613);
and U7903 (N_7903,N_5034,N_5331);
xor U7904 (N_7904,N_4735,N_4875);
or U7905 (N_7905,N_4790,N_4178);
and U7906 (N_7906,N_4780,N_5924);
nor U7907 (N_7907,N_4273,N_4114);
or U7908 (N_7908,N_5548,N_4703);
xor U7909 (N_7909,N_5640,N_4493);
or U7910 (N_7910,N_4393,N_4503);
or U7911 (N_7911,N_4432,N_5317);
or U7912 (N_7912,N_5756,N_5326);
nor U7913 (N_7913,N_5639,N_5643);
and U7914 (N_7914,N_5362,N_4099);
or U7915 (N_7915,N_5120,N_5587);
xnor U7916 (N_7916,N_5037,N_4399);
nand U7917 (N_7917,N_4816,N_5900);
and U7918 (N_7918,N_4170,N_5845);
nor U7919 (N_7919,N_4105,N_4111);
and U7920 (N_7920,N_4725,N_4167);
nand U7921 (N_7921,N_5387,N_5614);
or U7922 (N_7922,N_4682,N_5811);
nand U7923 (N_7923,N_4598,N_4894);
nand U7924 (N_7924,N_5742,N_5388);
nand U7925 (N_7925,N_4918,N_4150);
nor U7926 (N_7926,N_4682,N_5276);
xnor U7927 (N_7927,N_5557,N_4953);
or U7928 (N_7928,N_5274,N_4919);
or U7929 (N_7929,N_5855,N_4912);
nand U7930 (N_7930,N_5285,N_4376);
nand U7931 (N_7931,N_4258,N_5166);
nand U7932 (N_7932,N_4282,N_4507);
and U7933 (N_7933,N_5244,N_4964);
nand U7934 (N_7934,N_5124,N_4446);
and U7935 (N_7935,N_5526,N_5143);
and U7936 (N_7936,N_4964,N_4001);
xnor U7937 (N_7937,N_4863,N_4766);
nor U7938 (N_7938,N_5281,N_5549);
nor U7939 (N_7939,N_4411,N_5406);
and U7940 (N_7940,N_5850,N_5938);
nand U7941 (N_7941,N_5786,N_5652);
nand U7942 (N_7942,N_5892,N_5101);
and U7943 (N_7943,N_5497,N_5960);
and U7944 (N_7944,N_5491,N_5156);
xor U7945 (N_7945,N_4668,N_4955);
xor U7946 (N_7946,N_5806,N_4043);
nor U7947 (N_7947,N_5119,N_5718);
nor U7948 (N_7948,N_4325,N_5985);
and U7949 (N_7949,N_5766,N_4968);
xnor U7950 (N_7950,N_5345,N_5698);
nor U7951 (N_7951,N_5113,N_5263);
or U7952 (N_7952,N_5697,N_4636);
and U7953 (N_7953,N_4148,N_4534);
or U7954 (N_7954,N_5165,N_4714);
nor U7955 (N_7955,N_4065,N_4861);
and U7956 (N_7956,N_5235,N_4680);
nand U7957 (N_7957,N_4461,N_4035);
nand U7958 (N_7958,N_5127,N_4340);
nand U7959 (N_7959,N_4461,N_4576);
nor U7960 (N_7960,N_4558,N_5876);
and U7961 (N_7961,N_5340,N_4877);
nand U7962 (N_7962,N_5021,N_4370);
xnor U7963 (N_7963,N_4236,N_4605);
or U7964 (N_7964,N_5995,N_4910);
xor U7965 (N_7965,N_4595,N_5840);
nor U7966 (N_7966,N_5174,N_5175);
and U7967 (N_7967,N_5434,N_4695);
xor U7968 (N_7968,N_4948,N_5785);
nand U7969 (N_7969,N_5479,N_5777);
nand U7970 (N_7970,N_5731,N_4910);
nor U7971 (N_7971,N_5629,N_5612);
and U7972 (N_7972,N_5095,N_5176);
nand U7973 (N_7973,N_4322,N_4520);
nand U7974 (N_7974,N_4180,N_4829);
xor U7975 (N_7975,N_5725,N_4062);
and U7976 (N_7976,N_4437,N_5692);
nor U7977 (N_7977,N_4124,N_5246);
and U7978 (N_7978,N_5768,N_5745);
nor U7979 (N_7979,N_5527,N_5971);
nand U7980 (N_7980,N_4864,N_5466);
xnor U7981 (N_7981,N_5690,N_5361);
and U7982 (N_7982,N_5716,N_5808);
and U7983 (N_7983,N_4509,N_4293);
nand U7984 (N_7984,N_5260,N_4009);
nor U7985 (N_7985,N_4754,N_5796);
or U7986 (N_7986,N_5407,N_5111);
or U7987 (N_7987,N_4126,N_4325);
or U7988 (N_7988,N_4634,N_5343);
and U7989 (N_7989,N_4339,N_5402);
nor U7990 (N_7990,N_4807,N_4909);
or U7991 (N_7991,N_5086,N_4611);
xnor U7992 (N_7992,N_4625,N_5998);
and U7993 (N_7993,N_5358,N_4277);
nor U7994 (N_7994,N_4263,N_4589);
and U7995 (N_7995,N_5834,N_4111);
and U7996 (N_7996,N_4601,N_4786);
nand U7997 (N_7997,N_5834,N_4267);
nor U7998 (N_7998,N_5521,N_5882);
nand U7999 (N_7999,N_5566,N_4039);
and U8000 (N_8000,N_7427,N_6589);
nand U8001 (N_8001,N_6241,N_7714);
nor U8002 (N_8002,N_6822,N_6855);
or U8003 (N_8003,N_6335,N_7007);
nor U8004 (N_8004,N_7382,N_6323);
and U8005 (N_8005,N_6264,N_7064);
nand U8006 (N_8006,N_7393,N_7275);
nor U8007 (N_8007,N_6370,N_7837);
or U8008 (N_8008,N_7149,N_6240);
nor U8009 (N_8009,N_6140,N_7969);
nand U8010 (N_8010,N_7437,N_6563);
nor U8011 (N_8011,N_6372,N_7178);
nand U8012 (N_8012,N_7310,N_6986);
and U8013 (N_8013,N_7904,N_7550);
nand U8014 (N_8014,N_6384,N_7465);
nand U8015 (N_8015,N_6745,N_6162);
and U8016 (N_8016,N_7892,N_6319);
or U8017 (N_8017,N_7679,N_7506);
nor U8018 (N_8018,N_6266,N_7908);
and U8019 (N_8019,N_7971,N_7603);
nand U8020 (N_8020,N_6223,N_7419);
or U8021 (N_8021,N_6750,N_6772);
nand U8022 (N_8022,N_7758,N_7907);
nand U8023 (N_8023,N_7355,N_6925);
and U8024 (N_8024,N_7811,N_6255);
and U8025 (N_8025,N_7773,N_6485);
or U8026 (N_8026,N_7775,N_6183);
xnor U8027 (N_8027,N_7937,N_7162);
nand U8028 (N_8028,N_6990,N_6306);
nor U8029 (N_8029,N_6678,N_6890);
nor U8030 (N_8030,N_7566,N_6824);
nand U8031 (N_8031,N_7186,N_6254);
and U8032 (N_8032,N_7111,N_7745);
or U8033 (N_8033,N_6314,N_7863);
xor U8034 (N_8034,N_7120,N_7739);
or U8035 (N_8035,N_6521,N_7501);
or U8036 (N_8036,N_7831,N_7502);
nand U8037 (N_8037,N_6818,N_6560);
nor U8038 (N_8038,N_7420,N_6035);
and U8039 (N_8039,N_6505,N_7759);
nor U8040 (N_8040,N_6917,N_6624);
nand U8041 (N_8041,N_7700,N_7658);
nand U8042 (N_8042,N_6561,N_7598);
or U8043 (N_8043,N_6086,N_7050);
xor U8044 (N_8044,N_6136,N_6126);
or U8045 (N_8045,N_6340,N_6756);
nand U8046 (N_8046,N_6702,N_6186);
or U8047 (N_8047,N_6765,N_7191);
nand U8048 (N_8048,N_6840,N_6937);
or U8049 (N_8049,N_7099,N_6064);
or U8050 (N_8050,N_7877,N_6615);
and U8051 (N_8051,N_6111,N_7792);
nor U8052 (N_8052,N_6337,N_7042);
and U8053 (N_8053,N_7023,N_6009);
nand U8054 (N_8054,N_7358,N_6435);
nand U8055 (N_8055,N_7504,N_6565);
and U8056 (N_8056,N_6175,N_7970);
or U8057 (N_8057,N_6315,N_7839);
or U8058 (N_8058,N_6070,N_7314);
xnor U8059 (N_8059,N_7737,N_7810);
xnor U8060 (N_8060,N_6671,N_7469);
and U8061 (N_8061,N_6737,N_6530);
or U8062 (N_8062,N_7172,N_6815);
xor U8063 (N_8063,N_7161,N_7114);
nand U8064 (N_8064,N_6098,N_7479);
and U8065 (N_8065,N_6614,N_6396);
or U8066 (N_8066,N_6284,N_7905);
nor U8067 (N_8067,N_7915,N_7798);
nand U8068 (N_8068,N_6960,N_6873);
nand U8069 (N_8069,N_6891,N_7097);
nor U8070 (N_8070,N_6930,N_6845);
nor U8071 (N_8071,N_7194,N_6146);
xor U8072 (N_8072,N_6177,N_7637);
or U8073 (N_8073,N_7112,N_7140);
and U8074 (N_8074,N_6655,N_6522);
xnor U8075 (N_8075,N_6653,N_6871);
and U8076 (N_8076,N_7360,N_7132);
nor U8077 (N_8077,N_6688,N_7075);
xor U8078 (N_8078,N_7574,N_7176);
xor U8079 (N_8079,N_6101,N_7978);
or U8080 (N_8080,N_7865,N_7734);
or U8081 (N_8081,N_6041,N_7919);
xnor U8082 (N_8082,N_7183,N_7345);
xor U8083 (N_8083,N_7922,N_7941);
or U8084 (N_8084,N_7975,N_6328);
or U8085 (N_8085,N_6885,N_7681);
and U8086 (N_8086,N_7832,N_6191);
xnor U8087 (N_8087,N_6692,N_7932);
xor U8088 (N_8088,N_7680,N_7306);
xnor U8089 (N_8089,N_6385,N_6099);
nand U8090 (N_8090,N_7422,N_6279);
nor U8091 (N_8091,N_6131,N_6116);
and U8092 (N_8092,N_6346,N_6812);
xor U8093 (N_8093,N_6420,N_6034);
xor U8094 (N_8094,N_6302,N_6163);
nor U8095 (N_8095,N_6414,N_7282);
and U8096 (N_8096,N_6967,N_6612);
xor U8097 (N_8097,N_6458,N_6120);
nor U8098 (N_8098,N_6575,N_7763);
nor U8099 (N_8099,N_7193,N_6091);
nand U8100 (N_8100,N_6499,N_7782);
nor U8101 (N_8101,N_7640,N_7109);
xor U8102 (N_8102,N_7032,N_7418);
nor U8103 (N_8103,N_7646,N_6348);
or U8104 (N_8104,N_6501,N_7685);
and U8105 (N_8105,N_6578,N_7035);
nor U8106 (N_8106,N_7890,N_6043);
and U8107 (N_8107,N_7648,N_6428);
nor U8108 (N_8108,N_7968,N_6044);
xor U8109 (N_8109,N_7561,N_7215);
nor U8110 (N_8110,N_6569,N_6767);
or U8111 (N_8111,N_7198,N_7499);
xnor U8112 (N_8112,N_6675,N_6180);
nor U8113 (N_8113,N_7476,N_7600);
xnor U8114 (N_8114,N_7579,N_7138);
xnor U8115 (N_8115,N_6906,N_7014);
and U8116 (N_8116,N_6640,N_6293);
nor U8117 (N_8117,N_7088,N_7096);
nor U8118 (N_8118,N_6536,N_6790);
nand U8119 (N_8119,N_7587,N_6493);
and U8120 (N_8120,N_7742,N_6978);
nor U8121 (N_8121,N_6392,N_6069);
and U8122 (N_8122,N_6416,N_7185);
xor U8123 (N_8123,N_6461,N_7069);
nor U8124 (N_8124,N_6877,N_6651);
and U8125 (N_8125,N_6998,N_7724);
xnor U8126 (N_8126,N_7405,N_7697);
nand U8127 (N_8127,N_6915,N_6491);
xnor U8128 (N_8128,N_6940,N_6540);
and U8129 (N_8129,N_7616,N_7033);
xnor U8130 (N_8130,N_7066,N_7662);
nand U8131 (N_8131,N_7743,N_7268);
xor U8132 (N_8132,N_7725,N_7979);
xor U8133 (N_8133,N_7187,N_6492);
nand U8134 (N_8134,N_6637,N_7934);
nor U8135 (N_8135,N_7399,N_7993);
xor U8136 (N_8136,N_6247,N_6141);
nor U8137 (N_8137,N_7342,N_6579);
or U8138 (N_8138,N_7354,N_7816);
and U8139 (N_8139,N_6122,N_7131);
or U8140 (N_8140,N_7959,N_7361);
or U8141 (N_8141,N_6053,N_6789);
xnor U8142 (N_8142,N_7087,N_6061);
or U8143 (N_8143,N_7486,N_6841);
nand U8144 (N_8144,N_6332,N_7982);
and U8145 (N_8145,N_7580,N_6572);
and U8146 (N_8146,N_7693,N_6992);
xnor U8147 (N_8147,N_7206,N_6063);
xor U8148 (N_8148,N_7166,N_6574);
nor U8149 (N_8149,N_7404,N_7348);
or U8150 (N_8150,N_6798,N_6271);
or U8151 (N_8151,N_7551,N_6333);
and U8152 (N_8152,N_7108,N_6219);
nor U8153 (N_8153,N_7226,N_7933);
nand U8154 (N_8154,N_6145,N_6934);
or U8155 (N_8155,N_6135,N_6151);
nor U8156 (N_8156,N_7411,N_6365);
nand U8157 (N_8157,N_6759,N_7954);
nor U8158 (N_8158,N_6261,N_7458);
xor U8159 (N_8159,N_6113,N_6794);
xnor U8160 (N_8160,N_6797,N_7398);
or U8161 (N_8161,N_6339,N_6460);
nor U8162 (N_8162,N_6788,N_6431);
or U8163 (N_8163,N_6218,N_6698);
and U8164 (N_8164,N_7895,N_7562);
or U8165 (N_8165,N_7433,N_6415);
nor U8166 (N_8166,N_7536,N_6801);
and U8167 (N_8167,N_7860,N_7813);
nor U8168 (N_8168,N_6029,N_6948);
and U8169 (N_8169,N_6022,N_7723);
nor U8170 (N_8170,N_7535,N_7462);
and U8171 (N_8171,N_6094,N_6996);
and U8172 (N_8172,N_6581,N_7727);
xnor U8173 (N_8173,N_7844,N_6610);
xor U8174 (N_8174,N_7689,N_7105);
xor U8175 (N_8175,N_6665,N_6443);
nand U8176 (N_8176,N_7871,N_7488);
nor U8177 (N_8177,N_6733,N_6526);
and U8178 (N_8178,N_6107,N_6826);
and U8179 (N_8179,N_6344,N_6926);
nor U8180 (N_8180,N_6246,N_6080);
and U8181 (N_8181,N_7833,N_7443);
nor U8182 (N_8182,N_6310,N_7869);
xor U8183 (N_8183,N_6213,N_7841);
or U8184 (N_8184,N_6452,N_6825);
nor U8185 (N_8185,N_6831,N_7036);
nor U8186 (N_8186,N_6961,N_7164);
nor U8187 (N_8187,N_6495,N_7068);
nand U8188 (N_8188,N_6426,N_7079);
xor U8189 (N_8189,N_7948,N_7591);
or U8190 (N_8190,N_6320,N_7736);
xor U8191 (N_8191,N_6618,N_7421);
xor U8192 (N_8192,N_7874,N_6123);
xor U8193 (N_8193,N_7690,N_6763);
xor U8194 (N_8194,N_7704,N_7258);
or U8195 (N_8195,N_6016,N_7264);
and U8196 (N_8196,N_6676,N_7675);
xor U8197 (N_8197,N_6504,N_6931);
nand U8198 (N_8198,N_7912,N_7677);
and U8199 (N_8199,N_6580,N_6033);
xnor U8200 (N_8200,N_6601,N_7717);
nand U8201 (N_8201,N_7425,N_7756);
or U8202 (N_8202,N_7546,N_6820);
or U8203 (N_8203,N_7402,N_7651);
and U8204 (N_8204,N_7063,N_7925);
xor U8205 (N_8205,N_6245,N_6976);
or U8206 (N_8206,N_7791,N_6429);
xor U8207 (N_8207,N_6073,N_7503);
nor U8208 (N_8208,N_6525,N_7243);
and U8209 (N_8209,N_7262,N_7189);
nand U8210 (N_8210,N_7468,N_6630);
nand U8211 (N_8211,N_7156,N_7179);
or U8212 (N_8212,N_7249,N_6259);
xor U8213 (N_8213,N_7080,N_7853);
and U8214 (N_8214,N_7913,N_7668);
nand U8215 (N_8215,N_7999,N_7389);
or U8216 (N_8216,N_7167,N_7093);
nor U8217 (N_8217,N_6628,N_6250);
nand U8218 (N_8218,N_6235,N_7926);
nand U8219 (N_8219,N_6500,N_7357);
xor U8220 (N_8220,N_7766,N_7632);
and U8221 (N_8221,N_6634,N_7103);
xor U8222 (N_8222,N_6403,N_7362);
nor U8223 (N_8223,N_7726,N_6714);
and U8224 (N_8224,N_6078,N_7686);
xor U8225 (N_8225,N_7224,N_7441);
nand U8226 (N_8226,N_6411,N_7514);
xnor U8227 (N_8227,N_6418,N_6483);
and U8228 (N_8228,N_6467,N_7082);
nand U8229 (N_8229,N_7820,N_6887);
nor U8230 (N_8230,N_7383,N_7128);
xor U8231 (N_8231,N_6353,N_6555);
nand U8232 (N_8232,N_7928,N_7130);
or U8233 (N_8233,N_7430,N_6673);
or U8234 (N_8234,N_6090,N_7721);
xnor U8235 (N_8235,N_6853,N_7211);
or U8236 (N_8236,N_6055,N_7842);
nor U8237 (N_8237,N_7116,N_6524);
nand U8238 (N_8238,N_6898,N_6938);
nand U8239 (N_8239,N_6739,N_7478);
or U8240 (N_8240,N_7586,N_6636);
or U8241 (N_8241,N_6728,N_7322);
xor U8242 (N_8242,N_7802,N_7576);
nor U8243 (N_8243,N_7942,N_7494);
or U8244 (N_8244,N_6780,N_6660);
nor U8245 (N_8245,N_7448,N_6918);
nor U8246 (N_8246,N_7021,N_6686);
or U8247 (N_8247,N_6771,N_6298);
and U8248 (N_8248,N_6980,N_6030);
or U8249 (N_8249,N_6256,N_6024);
nand U8250 (N_8250,N_7822,N_7622);
nor U8251 (N_8251,N_6103,N_7744);
or U8252 (N_8252,N_7328,N_6129);
and U8253 (N_8253,N_7988,N_6587);
xnor U8254 (N_8254,N_6953,N_6008);
nor U8255 (N_8255,N_6550,N_7049);
nand U8256 (N_8256,N_6512,N_6260);
and U8257 (N_8257,N_7228,N_6814);
nand U8258 (N_8258,N_6547,N_6457);
or U8259 (N_8259,N_6642,N_6562);
or U8260 (N_8260,N_6791,N_6139);
or U8261 (N_8261,N_7929,N_6907);
nor U8262 (N_8262,N_7715,N_7254);
nand U8263 (N_8263,N_6047,N_7955);
or U8264 (N_8264,N_6272,N_6672);
and U8265 (N_8265,N_7412,N_7558);
nand U8266 (N_8266,N_7594,N_7327);
or U8267 (N_8267,N_6023,N_7118);
or U8268 (N_8268,N_6697,N_7720);
and U8269 (N_8269,N_7024,N_7223);
or U8270 (N_8270,N_7920,N_6622);
or U8271 (N_8271,N_6632,N_6280);
and U8272 (N_8272,N_6347,N_7438);
or U8273 (N_8273,N_6004,N_7770);
or U8274 (N_8274,N_6590,N_6072);
nand U8275 (N_8275,N_6856,N_7298);
nor U8276 (N_8276,N_6768,N_7573);
or U8277 (N_8277,N_6345,N_7692);
or U8278 (N_8278,N_7879,N_7409);
xnor U8279 (N_8279,N_6313,N_6923);
nand U8280 (N_8280,N_6723,N_7170);
nand U8281 (N_8281,N_7529,N_7150);
nand U8282 (N_8282,N_7481,N_6699);
nand U8283 (N_8283,N_7391,N_6317);
or U8284 (N_8284,N_6423,N_7017);
xor U8285 (N_8285,N_7455,N_7626);
nand U8286 (N_8286,N_6515,N_6189);
and U8287 (N_8287,N_7589,N_7649);
and U8288 (N_8288,N_6577,N_6503);
and U8289 (N_8289,N_6117,N_6731);
nor U8290 (N_8290,N_6706,N_7144);
xor U8291 (N_8291,N_6666,N_6963);
nand U8292 (N_8292,N_6785,N_7366);
nor U8293 (N_8293,N_7921,N_7305);
or U8294 (N_8294,N_6405,N_6970);
and U8295 (N_8295,N_7559,N_6496);
and U8296 (N_8296,N_6427,N_7076);
or U8297 (N_8297,N_7463,N_6851);
and U8298 (N_8298,N_7799,N_6067);
and U8299 (N_8299,N_7034,N_7682);
and U8300 (N_8300,N_6463,N_7266);
xor U8301 (N_8301,N_6708,N_7983);
and U8302 (N_8302,N_7623,N_6764);
or U8303 (N_8303,N_6582,N_6710);
nor U8304 (N_8304,N_6902,N_6670);
and U8305 (N_8305,N_6330,N_7577);
nor U8306 (N_8306,N_6208,N_6480);
or U8307 (N_8307,N_7741,N_6397);
xnor U8308 (N_8308,N_6349,N_6751);
nand U8309 (N_8309,N_6879,N_7147);
and U8310 (N_8310,N_7006,N_6296);
or U8311 (N_8311,N_6805,N_7270);
xor U8312 (N_8312,N_7136,N_7171);
nor U8313 (N_8313,N_6045,N_6051);
nor U8314 (N_8314,N_7701,N_6903);
nor U8315 (N_8315,N_6231,N_6417);
xor U8316 (N_8316,N_6506,N_7683);
and U8317 (N_8317,N_7825,N_7512);
nand U8318 (N_8318,N_6559,N_6015);
nor U8319 (N_8319,N_6534,N_7091);
nand U8320 (N_8320,N_7301,N_6529);
and U8321 (N_8321,N_7663,N_7731);
or U8322 (N_8322,N_6031,N_7849);
xor U8323 (N_8323,N_6509,N_6944);
or U8324 (N_8324,N_6881,N_7208);
and U8325 (N_8325,N_6644,N_7625);
nor U8326 (N_8326,N_7073,N_6957);
or U8327 (N_8327,N_7062,N_7380);
and U8328 (N_8328,N_7180,N_6594);
nor U8329 (N_8329,N_6721,N_6884);
nor U8330 (N_8330,N_7331,N_6849);
nand U8331 (N_8331,N_7340,N_7245);
or U8332 (N_8332,N_6584,N_7319);
or U8333 (N_8333,N_7875,N_6050);
nor U8334 (N_8334,N_6278,N_7552);
or U8335 (N_8335,N_7259,N_7516);
and U8336 (N_8336,N_6558,N_7220);
xnor U8337 (N_8337,N_6071,N_7896);
xnor U8338 (N_8338,N_7403,N_7547);
or U8339 (N_8339,N_6276,N_6571);
and U8340 (N_8340,N_6437,N_6715);
nand U8341 (N_8341,N_7210,N_6199);
and U8342 (N_8342,N_6746,N_7492);
nand U8343 (N_8343,N_7583,N_7753);
nor U8344 (N_8344,N_6952,N_6874);
or U8345 (N_8345,N_6696,N_6650);
and U8346 (N_8346,N_6413,N_7751);
nand U8347 (N_8347,N_6479,N_6987);
or U8348 (N_8348,N_7316,N_7273);
nand U8349 (N_8349,N_6220,N_7370);
nand U8350 (N_8350,N_7521,N_7363);
nor U8351 (N_8351,N_7263,N_6221);
nor U8352 (N_8352,N_7369,N_6065);
and U8353 (N_8353,N_6484,N_6950);
or U8354 (N_8354,N_7219,N_6544);
or U8355 (N_8355,N_7752,N_7661);
nand U8356 (N_8356,N_6664,N_6677);
nand U8357 (N_8357,N_6886,N_7851);
nand U8358 (N_8358,N_6943,N_7192);
and U8359 (N_8359,N_7949,N_6020);
nand U8360 (N_8360,N_6857,N_6685);
nor U8361 (N_8361,N_6170,N_7058);
and U8362 (N_8362,N_6424,N_6324);
xnor U8363 (N_8363,N_7055,N_6597);
and U8364 (N_8364,N_7564,N_6846);
or U8365 (N_8365,N_7522,N_6389);
and U8366 (N_8366,N_6309,N_7154);
nor U8367 (N_8367,N_7817,N_6681);
and U8368 (N_8368,N_6629,N_6487);
nor U8369 (N_8369,N_6916,N_6649);
xor U8370 (N_8370,N_7859,N_6011);
nor U8371 (N_8371,N_7713,N_6032);
nand U8372 (N_8372,N_7368,N_6108);
nor U8373 (N_8373,N_7688,N_6425);
xnor U8374 (N_8374,N_6573,N_7010);
xor U8375 (N_8375,N_7397,N_6088);
xnor U8376 (N_8376,N_7025,N_7801);
xnor U8377 (N_8377,N_6876,N_7257);
xnor U8378 (N_8378,N_7894,N_7635);
nor U8379 (N_8379,N_6956,N_7840);
xor U8380 (N_8380,N_7196,N_7045);
nand U8381 (N_8381,N_7041,N_6109);
and U8382 (N_8382,N_6007,N_6158);
or U8383 (N_8383,N_6894,N_6982);
and U8384 (N_8384,N_7325,N_6726);
nor U8385 (N_8385,N_6369,N_6985);
nand U8386 (N_8386,N_7239,N_6154);
nor U8387 (N_8387,N_7292,N_7803);
and U8388 (N_8388,N_7394,N_7652);
xor U8389 (N_8389,N_6367,N_7181);
or U8390 (N_8390,N_6176,N_7671);
nor U8391 (N_8391,N_7960,N_7065);
or U8392 (N_8392,N_6795,N_7195);
and U8393 (N_8393,N_7237,N_7485);
or U8394 (N_8394,N_7980,N_7207);
xnor U8395 (N_8395,N_6167,N_6134);
or U8396 (N_8396,N_7523,N_6687);
nand U8397 (N_8397,N_6478,N_7538);
nor U8398 (N_8398,N_7755,N_7706);
xnor U8399 (N_8399,N_7267,N_7784);
or U8400 (N_8400,N_6038,N_6476);
nand U8401 (N_8401,N_6603,N_7789);
or U8402 (N_8402,N_7235,N_7809);
nor U8403 (N_8403,N_6784,N_7990);
xnor U8404 (N_8404,N_7104,N_7555);
xor U8405 (N_8405,N_7148,N_7344);
xor U8406 (N_8406,N_7054,N_6647);
xor U8407 (N_8407,N_7406,N_6893);
nand U8408 (N_8408,N_7870,N_7324);
xnor U8409 (N_8409,N_6212,N_6769);
or U8410 (N_8410,N_7864,N_6527);
nand U8411 (N_8411,N_7563,N_6519);
xnor U8412 (N_8412,N_6188,N_6087);
or U8413 (N_8413,N_6124,N_6277);
or U8414 (N_8414,N_6355,N_7709);
nor U8415 (N_8415,N_7650,N_6740);
nor U8416 (N_8416,N_6823,N_6786);
nand U8417 (N_8417,N_6294,N_7029);
or U8418 (N_8418,N_6583,N_6837);
nand U8419 (N_8419,N_6844,N_7381);
xor U8420 (N_8420,N_7991,N_6779);
nor U8421 (N_8421,N_6502,N_6935);
xnor U8422 (N_8422,N_7606,N_6174);
and U8423 (N_8423,N_6516,N_6184);
or U8424 (N_8424,N_6734,N_6148);
nor U8425 (N_8425,N_6102,N_6236);
nor U8426 (N_8426,N_6471,N_6439);
and U8427 (N_8427,N_7276,N_7457);
and U8428 (N_8428,N_7155,N_6548);
nor U8429 (N_8429,N_7647,N_7216);
nor U8430 (N_8430,N_6566,N_7255);
or U8431 (N_8431,N_6546,N_6198);
or U8432 (N_8432,N_7777,N_7557);
nor U8433 (N_8433,N_7746,N_6895);
nand U8434 (N_8434,N_7044,N_6026);
xnor U8435 (N_8435,N_7101,N_6171);
or U8436 (N_8436,N_6747,N_7326);
xor U8437 (N_8437,N_7269,N_7423);
nand U8438 (N_8438,N_7053,N_6018);
xor U8439 (N_8439,N_6762,N_6766);
nand U8440 (N_8440,N_6468,N_7214);
or U8441 (N_8441,N_7442,N_7694);
and U8442 (N_8442,N_6444,N_6079);
nand U8443 (N_8443,N_6889,N_6659);
or U8444 (N_8444,N_7277,N_6984);
nor U8445 (N_8445,N_6991,N_7039);
nor U8446 (N_8446,N_6507,N_7473);
nor U8447 (N_8447,N_7795,N_7893);
xor U8448 (N_8448,N_6375,N_7601);
nor U8449 (N_8449,N_6568,N_7133);
nand U8450 (N_8450,N_6811,N_7401);
nor U8451 (N_8451,N_7785,N_7530);
and U8452 (N_8452,N_7918,N_6625);
or U8453 (N_8453,N_7554,N_6159);
nor U8454 (N_8454,N_7629,N_7260);
or U8455 (N_8455,N_6211,N_6738);
nor U8456 (N_8456,N_6588,N_7365);
xor U8457 (N_8457,N_7936,N_6989);
nand U8458 (N_8458,N_7227,N_6924);
or U8459 (N_8459,N_6060,N_6497);
nor U8460 (N_8460,N_6862,N_7923);
nand U8461 (N_8461,N_6813,N_6719);
nand U8462 (N_8462,N_7371,N_6858);
or U8463 (N_8463,N_6210,N_7061);
and U8464 (N_8464,N_7994,N_6914);
or U8465 (N_8465,N_7735,N_7716);
or U8466 (N_8466,N_7655,N_7317);
nand U8467 (N_8467,N_6274,N_6334);
nor U8468 (N_8468,N_7379,N_6808);
xor U8469 (N_8469,N_6513,N_6994);
or U8470 (N_8470,N_6226,N_6336);
or U8471 (N_8471,N_6363,N_7500);
or U8472 (N_8472,N_6402,N_7542);
xnor U8473 (N_8473,N_7318,N_6358);
nand U8474 (N_8474,N_7639,N_7122);
nor U8475 (N_8475,N_7445,N_7575);
nand U8476 (N_8476,N_7060,N_7461);
nor U8477 (N_8477,N_6596,N_6722);
nand U8478 (N_8478,N_6251,N_7549);
and U8479 (N_8479,N_6755,N_7519);
and U8480 (N_8480,N_7609,N_7084);
or U8481 (N_8481,N_6127,N_7410);
and U8482 (N_8482,N_7160,N_7838);
or U8483 (N_8483,N_6354,N_7852);
or U8484 (N_8484,N_7608,N_6446);
or U8485 (N_8485,N_7786,N_6248);
nand U8486 (N_8486,N_7856,N_7480);
or U8487 (N_8487,N_7703,N_7762);
nand U8488 (N_8488,N_7250,N_7687);
or U8489 (N_8489,N_7177,N_7669);
nor U8490 (N_8490,N_6633,N_6643);
nand U8491 (N_8491,N_7887,N_7158);
nand U8492 (N_8492,N_7888,N_7508);
and U8493 (N_8493,N_6850,N_6627);
and U8494 (N_8494,N_6743,N_6754);
xor U8495 (N_8495,N_6690,N_7855);
xor U8496 (N_8496,N_7184,N_7779);
xnor U8497 (N_8497,N_7299,N_6979);
or U8498 (N_8498,N_7578,N_7607);
or U8499 (N_8499,N_7987,N_7986);
or U8500 (N_8500,N_6433,N_7854);
nand U8501 (N_8501,N_7311,N_7173);
xor U8502 (N_8502,N_6028,N_7627);
nand U8503 (N_8503,N_7885,N_6908);
or U8504 (N_8504,N_6966,N_6783);
xor U8505 (N_8505,N_7051,N_7951);
and U8506 (N_8506,N_7056,N_7595);
and U8507 (N_8507,N_6693,N_7436);
xnor U8508 (N_8508,N_6475,N_7621);
nand U8509 (N_8509,N_6974,N_7152);
or U8510 (N_8510,N_7287,N_7916);
or U8511 (N_8511,N_7452,N_7336);
or U8512 (N_8512,N_7279,N_7944);
xnor U8513 (N_8513,N_6449,N_7572);
nor U8514 (N_8514,N_6451,N_6341);
nand U8515 (N_8515,N_7560,N_7303);
nor U8516 (N_8516,N_7238,N_6883);
or U8517 (N_8517,N_6804,N_7083);
or U8518 (N_8518,N_7891,N_7234);
nand U8519 (N_8519,N_7761,N_7013);
or U8520 (N_8520,N_6166,N_6753);
or U8521 (N_8521,N_6912,N_7902);
or U8522 (N_8522,N_6608,N_7028);
nand U8523 (N_8523,N_7927,N_7300);
nand U8524 (N_8524,N_6459,N_7372);
and U8525 (N_8525,N_7684,N_7212);
nand U8526 (N_8526,N_7898,N_7197);
xnor U8527 (N_8527,N_6379,N_6816);
nor U8528 (N_8528,N_6181,N_6904);
or U8529 (N_8529,N_6230,N_6517);
nand U8530 (N_8530,N_7593,N_7272);
xnor U8531 (N_8531,N_7347,N_6172);
nand U8532 (N_8532,N_6381,N_6056);
nor U8533 (N_8533,N_7037,N_7643);
nor U8534 (N_8534,N_6639,N_7280);
or U8535 (N_8535,N_6932,N_6421);
nor U8536 (N_8536,N_6455,N_6861);
nor U8537 (N_8537,N_7539,N_7989);
or U8538 (N_8538,N_6679,N_7966);
and U8539 (N_8539,N_7884,N_7910);
nor U8540 (N_8540,N_7571,N_6453);
nand U8541 (N_8541,N_7533,N_6286);
nor U8542 (N_8542,N_7806,N_7783);
nand U8543 (N_8543,N_7001,N_7861);
and U8544 (N_8544,N_7163,N_7828);
or U8545 (N_8545,N_7829,N_7387);
xor U8546 (N_8546,N_7540,N_7435);
or U8547 (N_8547,N_7175,N_6292);
or U8548 (N_8548,N_7581,N_6273);
nand U8549 (N_8549,N_6287,N_7092);
nand U8550 (N_8550,N_6169,N_6173);
nor U8551 (N_8551,N_6981,N_6720);
or U8552 (N_8552,N_7511,N_7780);
or U8553 (N_8553,N_6125,N_6267);
xor U8554 (N_8554,N_7498,N_6867);
or U8555 (N_8555,N_6378,N_7534);
or U8556 (N_8556,N_6371,N_6342);
or U8557 (N_8557,N_7788,N_6312);
and U8558 (N_8558,N_7698,N_6598);
xnor U8559 (N_8559,N_6775,N_7107);
nand U8560 (N_8560,N_6983,N_6133);
nand U8561 (N_8561,N_6322,N_6288);
xor U8562 (N_8562,N_7222,N_6204);
nor U8563 (N_8563,N_7330,N_7641);
and U8564 (N_8564,N_7346,N_6835);
or U8565 (N_8565,N_7961,N_6465);
or U8566 (N_8566,N_7545,N_7602);
nor U8567 (N_8567,N_6012,N_7353);
and U8568 (N_8568,N_6195,N_7477);
and U8569 (N_8569,N_7938,N_6239);
xnor U8570 (N_8570,N_6374,N_6541);
and U8571 (N_8571,N_6607,N_7283);
and U8572 (N_8572,N_6075,N_6570);
or U8573 (N_8573,N_6318,N_6165);
xnor U8574 (N_8574,N_6532,N_6695);
nand U8575 (N_8575,N_6238,N_6661);
xor U8576 (N_8576,N_7444,N_6326);
or U8577 (N_8577,N_7011,N_6006);
nor U8578 (N_8578,N_7190,N_6445);
nand U8579 (N_8579,N_6593,N_6782);
nand U8580 (N_8580,N_7836,N_6839);
nor U8581 (N_8581,N_7141,N_6712);
nand U8582 (N_8582,N_6511,N_6498);
and U8583 (N_8583,N_7781,N_7146);
xor U8584 (N_8584,N_6711,N_7981);
xnor U8585 (N_8585,N_7794,N_6860);
nor U8586 (N_8586,N_6683,N_6488);
nand U8587 (N_8587,N_7230,N_6110);
and U8588 (N_8588,N_7957,N_6652);
nor U8589 (N_8589,N_6399,N_7413);
and U8590 (N_8590,N_7707,N_6951);
or U8591 (N_8591,N_6000,N_6949);
nor U8592 (N_8592,N_7225,N_6658);
nand U8593 (N_8593,N_7945,N_7159);
nand U8594 (N_8594,N_7285,N_7467);
nand U8595 (N_8595,N_7483,N_7857);
xnor U8596 (N_8596,N_7899,N_6486);
xor U8597 (N_8597,N_6535,N_6263);
xnor U8598 (N_8598,N_6234,N_6977);
or U8599 (N_8599,N_6833,N_7553);
xnor U8600 (N_8600,N_7732,N_6096);
nor U8601 (N_8601,N_7914,N_6473);
nor U8602 (N_8602,N_7673,N_7872);
xnor U8603 (N_8603,N_6209,N_7135);
and U8604 (N_8604,N_7124,N_7205);
xor U8605 (N_8605,N_6197,N_7390);
xor U8606 (N_8606,N_7143,N_6836);
and U8607 (N_8607,N_7610,N_6729);
xnor U8608 (N_8608,N_7656,N_6168);
nand U8609 (N_8609,N_6185,N_7434);
nor U8610 (N_8610,N_6806,N_7653);
and U8611 (N_8611,N_6549,N_6899);
and U8612 (N_8612,N_7524,N_6252);
nand U8613 (N_8613,N_7209,N_6817);
and U8614 (N_8614,N_6407,N_6537);
and U8615 (N_8615,N_6508,N_7375);
nand U8616 (N_8616,N_6888,N_6275);
xor U8617 (N_8617,N_6422,N_6842);
and U8618 (N_8618,N_7556,N_7525);
nor U8619 (N_8619,N_7518,N_7078);
or U8620 (N_8620,N_6228,N_7286);
or U8621 (N_8621,N_6338,N_6291);
and U8622 (N_8622,N_7295,N_6510);
xor U8623 (N_8623,N_7567,N_6115);
nand U8624 (N_8624,N_7787,N_6447);
nor U8625 (N_8625,N_6440,N_6048);
nand U8626 (N_8626,N_6377,N_7098);
nand U8627 (N_8627,N_7520,N_6289);
nor U8628 (N_8628,N_6864,N_6972);
nor U8629 (N_8629,N_7240,N_7510);
xor U8630 (N_8630,N_7985,N_6905);
nor U8631 (N_8631,N_7634,N_6058);
and U8632 (N_8632,N_6357,N_6704);
nand U8633 (N_8633,N_6939,N_7826);
and U8634 (N_8634,N_7901,N_6434);
and U8635 (N_8635,N_6626,N_6591);
xnor U8636 (N_8636,N_6155,N_7672);
nor U8637 (N_8637,N_7474,N_6376);
xnor U8638 (N_8638,N_6013,N_6114);
nor U8639 (N_8639,N_6222,N_7747);
or U8640 (N_8640,N_6436,N_6466);
nand U8641 (N_8641,N_6062,N_6217);
nand U8642 (N_8642,N_7491,N_7281);
or U8643 (N_8643,N_7233,N_6616);
xnor U8644 (N_8644,N_7376,N_7095);
or U8645 (N_8645,N_6147,N_6327);
xnor U8646 (N_8646,N_7699,N_6773);
xnor U8647 (N_8647,N_6838,N_6684);
xor U8648 (N_8648,N_7384,N_7200);
or U8649 (N_8649,N_7617,N_6599);
xor U8650 (N_8650,N_7417,N_6928);
or U8651 (N_8651,N_6393,N_6490);
nand U8652 (N_8652,N_7440,N_7392);
nor U8653 (N_8653,N_7995,N_7008);
nand U8654 (N_8654,N_6001,N_6933);
or U8655 (N_8655,N_7660,N_6859);
and U8656 (N_8656,N_7998,N_6395);
nand U8657 (N_8657,N_7090,N_6303);
or U8658 (N_8658,N_6809,N_6359);
and U8659 (N_8659,N_7174,N_6406);
or U8660 (N_8660,N_7248,N_6454);
nor U8661 (N_8661,N_6225,N_6143);
or U8662 (N_8662,N_7909,N_7772);
or U8663 (N_8663,N_7628,N_7696);
and U8664 (N_8664,N_6605,N_7102);
nor U8665 (N_8665,N_6648,N_6988);
nand U8666 (N_8666,N_7415,N_7456);
xor U8667 (N_8667,N_6366,N_6361);
and U8668 (N_8668,N_7016,N_6713);
nand U8669 (N_8669,N_7339,N_6297);
nand U8670 (N_8670,N_6538,N_6299);
nand U8671 (N_8671,N_6304,N_7796);
and U8672 (N_8672,N_6863,N_6606);
xnor U8673 (N_8673,N_6682,N_7447);
nor U8674 (N_8674,N_6964,N_7862);
and U8675 (N_8675,N_6142,N_7352);
xnor U8676 (N_8676,N_7315,N_6157);
nor U8677 (N_8677,N_7897,N_7288);
or U8678 (N_8678,N_6866,N_7867);
and U8679 (N_8679,N_7965,N_6761);
or U8680 (N_8680,N_7962,N_7620);
or U8681 (N_8681,N_6997,N_6481);
xnor U8682 (N_8682,N_6777,N_7261);
or U8683 (N_8683,N_7244,N_6257);
nand U8684 (N_8684,N_6046,N_6796);
xnor U8685 (N_8685,N_6200,N_7738);
xor U8686 (N_8686,N_6042,N_6609);
nor U8687 (N_8687,N_7086,N_6554);
or U8688 (N_8688,N_6082,N_6380);
nand U8689 (N_8689,N_7373,N_6130);
nand U8690 (N_8690,N_7242,N_6694);
nand U8691 (N_8691,N_7819,N_7931);
xor U8692 (N_8692,N_7880,N_7309);
or U8693 (N_8693,N_7843,N_7251);
xor U8694 (N_8694,N_6190,N_7515);
xnor U8695 (N_8695,N_7431,N_6160);
or U8696 (N_8696,N_6656,N_6442);
or U8697 (N_8697,N_6450,N_7719);
or U8698 (N_8698,N_6520,N_6669);
nand U8699 (N_8699,N_6623,N_6999);
nor U8700 (N_8700,N_7030,N_7695);
or U8701 (N_8701,N_7236,N_7129);
nor U8702 (N_8702,N_7125,N_6432);
and U8703 (N_8703,N_6464,N_6388);
nand U8704 (N_8704,N_6270,N_6595);
nand U8705 (N_8705,N_6909,N_7807);
and U8706 (N_8706,N_7253,N_7484);
nor U8707 (N_8707,N_7590,N_7284);
nand U8708 (N_8708,N_6821,N_7271);
nor U8709 (N_8709,N_6282,N_7454);
nand U8710 (N_8710,N_7302,N_6631);
nand U8711 (N_8711,N_7830,N_7824);
xnor U8712 (N_8712,N_6128,N_6205);
nor U8713 (N_8713,N_7568,N_6958);
and U8714 (N_8714,N_7472,N_7338);
xor U8715 (N_8715,N_7702,N_7790);
nor U8716 (N_8716,N_6368,N_6586);
or U8717 (N_8717,N_6705,N_7847);
nor U8718 (N_8718,N_6819,N_7489);
and U8719 (N_8719,N_6039,N_6531);
nand U8720 (N_8720,N_6242,N_7085);
nand U8721 (N_8721,N_7946,N_6576);
and U8722 (N_8722,N_7115,N_7071);
xnor U8723 (N_8723,N_7749,N_7505);
and U8724 (N_8724,N_7113,N_7048);
nor U8725 (N_8725,N_7597,N_7611);
nand U8726 (N_8726,N_7015,N_7881);
or U8727 (N_8727,N_7077,N_6408);
and U8728 (N_8728,N_6946,N_7351);
or U8729 (N_8729,N_7570,N_7614);
xor U8730 (N_8730,N_6178,N_6691);
nand U8731 (N_8731,N_6489,N_6021);
xor U8732 (N_8732,N_7517,N_7997);
xor U8733 (N_8733,N_6965,N_6438);
and U8734 (N_8734,N_6741,N_6744);
and U8735 (N_8735,N_6118,N_6456);
nand U8736 (N_8736,N_7182,N_6774);
xnor U8737 (N_8737,N_7636,N_6716);
nand U8738 (N_8738,N_7953,N_6232);
xor U8739 (N_8739,N_7121,N_6703);
xor U8740 (N_8740,N_6258,N_7110);
nor U8741 (N_8741,N_7889,N_7100);
nand U8742 (N_8742,N_7585,N_6077);
nand U8743 (N_8743,N_7711,N_6927);
xnor U8744 (N_8744,N_6364,N_6237);
and U8745 (N_8745,N_7026,N_7312);
nor U8746 (N_8746,N_7203,N_7057);
nand U8747 (N_8747,N_6718,N_7134);
and U8748 (N_8748,N_6727,N_7619);
xnor U8749 (N_8749,N_6193,N_6757);
and U8750 (N_8750,N_7604,N_7332);
xor U8751 (N_8751,N_6089,N_6621);
or U8752 (N_8752,N_6105,N_7814);
nand U8753 (N_8753,N_7691,N_6095);
xor U8754 (N_8754,N_6880,N_7012);
nor U8755 (N_8755,N_6373,N_7883);
nor U8756 (N_8756,N_7667,N_6828);
or U8757 (N_8757,N_7665,N_6973);
and U8758 (N_8758,N_6229,N_7333);
and U8759 (N_8759,N_6083,N_7018);
xnor U8760 (N_8760,N_6602,N_6352);
nor U8761 (N_8761,N_6093,N_6410);
or U8762 (N_8762,N_6325,N_7967);
xor U8763 (N_8763,N_7126,N_7526);
or U8764 (N_8764,N_6638,N_7106);
xor U8765 (N_8765,N_7396,N_7544);
xor U8766 (N_8766,N_7157,N_7657);
xnor U8767 (N_8767,N_6224,N_6002);
nor U8768 (N_8768,N_7072,N_6494);
xor U8769 (N_8769,N_7776,N_6268);
nor U8770 (N_8770,N_7052,N_7878);
xor U8771 (N_8771,N_6202,N_7769);
nand U8772 (N_8772,N_6617,N_7343);
nand U8773 (N_8773,N_7548,N_7618);
nor U8774 (N_8774,N_7977,N_7202);
and U8775 (N_8775,N_6567,N_6350);
xnor U8776 (N_8776,N_7644,N_6390);
nand U8777 (N_8777,N_6900,N_6802);
nand U8778 (N_8778,N_7605,N_7385);
nand U8779 (N_8779,N_7232,N_6611);
and U8780 (N_8780,N_7323,N_7674);
xor U8781 (N_8781,N_7426,N_6085);
and U8782 (N_8782,N_6482,N_6604);
nor U8783 (N_8783,N_6799,N_7470);
xnor U8784 (N_8784,N_7710,N_6138);
and U8785 (N_8785,N_7497,N_6144);
nor U8786 (N_8786,N_7337,N_7019);
and U8787 (N_8787,N_7424,N_7475);
nand U8788 (N_8788,N_6843,N_7308);
xnor U8789 (N_8789,N_6793,N_7708);
or U8790 (N_8790,N_6156,N_6149);
nor U8791 (N_8791,N_7757,N_7670);
or U8792 (N_8792,N_7527,N_6019);
and U8793 (N_8793,N_6872,N_6736);
and U8794 (N_8794,N_7868,N_7296);
nor U8795 (N_8795,N_7117,N_6954);
nor U8796 (N_8796,N_7313,N_6412);
and U8797 (N_8797,N_7451,N_6321);
nand U8798 (N_8798,N_7845,N_6360);
xor U8799 (N_8799,N_6187,N_6929);
xnor U8800 (N_8800,N_6331,N_7217);
or U8801 (N_8801,N_6878,N_6585);
nand U8802 (N_8802,N_6539,N_7320);
nor U8803 (N_8803,N_7040,N_6285);
nor U8804 (N_8804,N_6945,N_6832);
and U8805 (N_8805,N_7229,N_7973);
nand U8806 (N_8806,N_7613,N_6092);
nand U8807 (N_8807,N_6005,N_6057);
xor U8808 (N_8808,N_6758,N_7615);
nand U8809 (N_8809,N_7005,N_6781);
or U8810 (N_8810,N_7070,N_6295);
and U8811 (N_8811,N_7213,N_7654);
xor U8812 (N_8812,N_7569,N_6641);
and U8813 (N_8813,N_7750,N_7231);
nor U8814 (N_8814,N_6387,N_7031);
and U8815 (N_8815,N_6201,N_7046);
or U8816 (N_8816,N_7407,N_7906);
nand U8817 (N_8817,N_7432,N_7378);
and U8818 (N_8818,N_7341,N_6474);
and U8819 (N_8819,N_7730,N_7256);
nor U8820 (N_8820,N_7374,N_7291);
or U8821 (N_8821,N_7356,N_6362);
and U8822 (N_8822,N_6619,N_6897);
or U8823 (N_8823,N_7367,N_6316);
and U8824 (N_8824,N_6654,N_6896);
xor U8825 (N_8825,N_6132,N_6441);
or U8826 (N_8826,N_6830,N_6730);
and U8827 (N_8827,N_7464,N_7359);
or U8828 (N_8828,N_6523,N_7119);
nor U8829 (N_8829,N_6760,N_6081);
or U8830 (N_8830,N_7638,N_7002);
xor U8831 (N_8831,N_7764,N_7835);
nor U8832 (N_8832,N_6735,N_7588);
and U8833 (N_8833,N_6847,N_7247);
nand U8834 (N_8834,N_6305,N_6192);
nor U8835 (N_8835,N_7297,N_7976);
or U8836 (N_8836,N_6552,N_7000);
nor U8837 (N_8837,N_6419,N_6680);
nand U8838 (N_8838,N_7507,N_7047);
and U8839 (N_8839,N_6792,N_6551);
or U8840 (N_8840,N_6329,N_6137);
or U8841 (N_8841,N_7349,N_6301);
nand U8842 (N_8842,N_6382,N_6036);
or U8843 (N_8843,N_6343,N_7754);
nand U8844 (N_8844,N_7850,N_6153);
and U8845 (N_8845,N_7678,N_6564);
xnor U8846 (N_8846,N_6283,N_7950);
or U8847 (N_8847,N_7705,N_6076);
nand U8848 (N_8848,N_6748,N_6469);
or U8849 (N_8849,N_6752,N_6968);
nor U8850 (N_8850,N_7165,N_7142);
nor U8851 (N_8851,N_6100,N_6613);
nor U8852 (N_8852,N_7460,N_6725);
nand U8853 (N_8853,N_6959,N_6203);
and U8854 (N_8854,N_7329,N_7428);
xor U8855 (N_8855,N_6807,N_6645);
or U8856 (N_8856,N_7408,N_6962);
xor U8857 (N_8857,N_7350,N_7924);
xnor U8858 (N_8858,N_7565,N_7972);
and U8859 (N_8859,N_7659,N_7963);
or U8860 (N_8860,N_7123,N_6401);
nand U8861 (N_8861,N_7771,N_7496);
and U8862 (N_8862,N_6514,N_7471);
nand U8863 (N_8863,N_7917,N_6383);
nand U8864 (N_8864,N_6206,N_6955);
nand U8865 (N_8865,N_7531,N_6179);
xor U8866 (N_8866,N_7139,N_6911);
nand U8867 (N_8867,N_7509,N_7094);
or U8868 (N_8868,N_6971,N_7939);
nand U8869 (N_8869,N_6920,N_6037);
xor U8870 (N_8870,N_7774,N_7416);
xnor U8871 (N_8871,N_6253,N_7958);
or U8872 (N_8872,N_7151,N_7612);
or U8873 (N_8873,N_7582,N_7022);
xnor U8874 (N_8874,N_7137,N_7386);
nor U8875 (N_8875,N_7274,N_7265);
nor U8876 (N_8876,N_7541,N_7278);
and U8877 (N_8877,N_6827,N_6112);
xnor U8878 (N_8878,N_6533,N_7188);
nor U8879 (N_8879,N_7974,N_6732);
nor U8880 (N_8880,N_6054,N_7020);
or U8881 (N_8881,N_6281,N_6216);
nor U8882 (N_8882,N_6667,N_6942);
and U8883 (N_8883,N_7513,N_6707);
xnor U8884 (N_8884,N_7866,N_6701);
or U8885 (N_8885,N_6668,N_7168);
or U8886 (N_8886,N_6635,N_7089);
nand U8887 (N_8887,N_7388,N_6084);
xnor U8888 (N_8888,N_7027,N_6936);
or U8889 (N_8889,N_7493,N_7903);
and U8890 (N_8890,N_7992,N_6662);
nand U8891 (N_8891,N_6243,N_6300);
nor U8892 (N_8892,N_6472,N_7943);
nand U8893 (N_8893,N_6674,N_6848);
or U8894 (N_8894,N_6040,N_7289);
nand U8895 (N_8895,N_7778,N_7848);
or U8896 (N_8896,N_6409,N_7858);
xnor U8897 (N_8897,N_6869,N_7081);
or U8898 (N_8898,N_6249,N_6307);
and U8899 (N_8899,N_7827,N_6742);
and U8900 (N_8900,N_7768,N_6803);
and U8901 (N_8901,N_7074,N_7952);
and U8902 (N_8902,N_6700,N_6106);
or U8903 (N_8903,N_6657,N_6121);
xor U8904 (N_8904,N_7009,N_6356);
and U8905 (N_8905,N_6620,N_6901);
xor U8906 (N_8906,N_6400,N_7722);
nor U8907 (N_8907,N_7728,N_7414);
or U8908 (N_8908,N_7935,N_6066);
nand U8909 (N_8909,N_6969,N_6150);
nor U8910 (N_8910,N_6027,N_7400);
xor U8911 (N_8911,N_6404,N_6553);
xnor U8912 (N_8912,N_7145,N_7334);
nor U8913 (N_8913,N_7767,N_6975);
and U8914 (N_8914,N_6941,N_6059);
nand U8915 (N_8915,N_6182,N_7153);
or U8916 (N_8916,N_6269,N_6462);
or U8917 (N_8917,N_6290,N_7818);
nand U8918 (N_8918,N_6068,N_7290);
nand U8919 (N_8919,N_6800,N_6870);
and U8920 (N_8920,N_6910,N_7718);
or U8921 (N_8921,N_7450,N_7712);
xor U8922 (N_8922,N_6545,N_6543);
nor U8923 (N_8923,N_7429,N_7446);
nand U8924 (N_8924,N_6207,N_6074);
or U8925 (N_8925,N_7733,N_7930);
and U8926 (N_8926,N_7624,N_7873);
nand U8927 (N_8927,N_7676,N_7439);
or U8928 (N_8928,N_6689,N_7364);
and U8929 (N_8929,N_6875,N_7466);
and U8930 (N_8930,N_7241,N_7252);
xor U8931 (N_8931,N_7940,N_6477);
nand U8932 (N_8932,N_7482,N_6164);
nand U8933 (N_8933,N_7876,N_6049);
and U8934 (N_8934,N_6161,N_7537);
and U8935 (N_8935,N_6556,N_7630);
xnor U8936 (N_8936,N_6663,N_7201);
nor U8937 (N_8937,N_6311,N_7911);
or U8938 (N_8938,N_6119,N_7834);
xnor U8939 (N_8939,N_7808,N_6194);
nor U8940 (N_8940,N_6600,N_6386);
nand U8941 (N_8941,N_7631,N_7584);
and U8942 (N_8942,N_6351,N_6227);
or U8943 (N_8943,N_7760,N_6717);
or U8944 (N_8944,N_7218,N_7294);
or U8945 (N_8945,N_6868,N_7821);
and U8946 (N_8946,N_6854,N_6196);
xnor U8947 (N_8947,N_6947,N_6017);
nor U8948 (N_8948,N_6391,N_7490);
and U8949 (N_8949,N_6003,N_7127);
or U8950 (N_8950,N_6244,N_7199);
and U8951 (N_8951,N_7812,N_7846);
and U8952 (N_8952,N_6995,N_7307);
nand U8953 (N_8953,N_7642,N_6052);
xnor U8954 (N_8954,N_7321,N_6215);
nand U8955 (N_8955,N_7645,N_6865);
and U8956 (N_8956,N_7495,N_7996);
and U8957 (N_8957,N_6724,N_7043);
or U8958 (N_8958,N_7815,N_7003);
nor U8959 (N_8959,N_6528,N_7453);
nor U8960 (N_8960,N_6265,N_7797);
nand U8961 (N_8961,N_7765,N_7459);
or U8962 (N_8962,N_6922,N_7882);
or U8963 (N_8963,N_6770,N_7293);
or U8964 (N_8964,N_6892,N_7804);
and U8965 (N_8965,N_6262,N_7395);
nor U8966 (N_8966,N_7204,N_7246);
and U8967 (N_8967,N_7633,N_6749);
xnor U8968 (N_8968,N_7740,N_6913);
nor U8969 (N_8969,N_6829,N_7900);
nand U8970 (N_8970,N_6152,N_7793);
nand U8971 (N_8971,N_6919,N_6776);
and U8972 (N_8972,N_6810,N_6394);
or U8973 (N_8973,N_6010,N_6709);
or U8974 (N_8974,N_6592,N_6542);
or U8975 (N_8975,N_7599,N_7964);
or U8976 (N_8976,N_7377,N_7532);
nand U8977 (N_8977,N_7664,N_7805);
and U8978 (N_8978,N_7956,N_7004);
xnor U8979 (N_8979,N_6233,N_7487);
and U8980 (N_8980,N_6308,N_7169);
or U8981 (N_8981,N_6014,N_6834);
or U8982 (N_8982,N_6882,N_7543);
or U8983 (N_8983,N_6025,N_6646);
nor U8984 (N_8984,N_7304,N_6518);
nand U8985 (N_8985,N_7335,N_6778);
and U8986 (N_8986,N_7059,N_7038);
and U8987 (N_8987,N_7984,N_6921);
or U8988 (N_8988,N_7596,N_7886);
and U8989 (N_8989,N_6448,N_6557);
nor U8990 (N_8990,N_7592,N_7666);
xor U8991 (N_8991,N_6993,N_7449);
and U8992 (N_8992,N_6430,N_6214);
xor U8993 (N_8993,N_7067,N_7823);
nor U8994 (N_8994,N_7947,N_7800);
and U8995 (N_8995,N_6470,N_7528);
and U8996 (N_8996,N_6398,N_6097);
nor U8997 (N_8997,N_6104,N_6787);
nand U8998 (N_8998,N_6852,N_7729);
and U8999 (N_8999,N_7748,N_7221);
xnor U9000 (N_9000,N_6204,N_6740);
nand U9001 (N_9001,N_7886,N_6092);
or U9002 (N_9002,N_7214,N_6144);
and U9003 (N_9003,N_7647,N_7230);
and U9004 (N_9004,N_7940,N_7656);
nand U9005 (N_9005,N_6835,N_6347);
or U9006 (N_9006,N_7989,N_6642);
and U9007 (N_9007,N_7965,N_6723);
or U9008 (N_9008,N_6844,N_6766);
nor U9009 (N_9009,N_7000,N_6581);
or U9010 (N_9010,N_7293,N_7485);
or U9011 (N_9011,N_7876,N_6248);
and U9012 (N_9012,N_6803,N_7086);
and U9013 (N_9013,N_6039,N_7677);
nand U9014 (N_9014,N_6580,N_6657);
or U9015 (N_9015,N_7591,N_7890);
or U9016 (N_9016,N_6788,N_6712);
and U9017 (N_9017,N_6477,N_7469);
xnor U9018 (N_9018,N_6845,N_6941);
nand U9019 (N_9019,N_6310,N_6880);
nand U9020 (N_9020,N_6041,N_7285);
nand U9021 (N_9021,N_6317,N_6580);
xnor U9022 (N_9022,N_6368,N_7926);
nand U9023 (N_9023,N_7322,N_6966);
nand U9024 (N_9024,N_7651,N_7035);
nand U9025 (N_9025,N_7053,N_6108);
and U9026 (N_9026,N_6410,N_6735);
or U9027 (N_9027,N_7666,N_6825);
nand U9028 (N_9028,N_7207,N_7015);
xor U9029 (N_9029,N_7965,N_6549);
nand U9030 (N_9030,N_7469,N_7794);
xor U9031 (N_9031,N_7169,N_7164);
nand U9032 (N_9032,N_6737,N_6571);
nor U9033 (N_9033,N_7602,N_6334);
nor U9034 (N_9034,N_7058,N_6507);
and U9035 (N_9035,N_6480,N_6721);
nand U9036 (N_9036,N_7257,N_7289);
nand U9037 (N_9037,N_7355,N_6631);
xor U9038 (N_9038,N_7053,N_7543);
nand U9039 (N_9039,N_7602,N_7990);
nand U9040 (N_9040,N_6316,N_7858);
xnor U9041 (N_9041,N_7126,N_6676);
nand U9042 (N_9042,N_6279,N_7624);
xor U9043 (N_9043,N_7572,N_6775);
and U9044 (N_9044,N_6581,N_7522);
nor U9045 (N_9045,N_7696,N_7727);
xnor U9046 (N_9046,N_6891,N_7898);
and U9047 (N_9047,N_6113,N_7649);
xnor U9048 (N_9048,N_6658,N_7583);
or U9049 (N_9049,N_7316,N_6139);
nor U9050 (N_9050,N_6669,N_7628);
xnor U9051 (N_9051,N_6910,N_7224);
and U9052 (N_9052,N_7347,N_7174);
and U9053 (N_9053,N_7205,N_7220);
xor U9054 (N_9054,N_6436,N_7472);
xor U9055 (N_9055,N_6042,N_7122);
nor U9056 (N_9056,N_7116,N_7321);
and U9057 (N_9057,N_7865,N_6854);
nand U9058 (N_9058,N_6354,N_6808);
xor U9059 (N_9059,N_7700,N_7112);
or U9060 (N_9060,N_7978,N_7036);
and U9061 (N_9061,N_7532,N_7084);
nor U9062 (N_9062,N_6424,N_7930);
nand U9063 (N_9063,N_6233,N_6270);
or U9064 (N_9064,N_6121,N_7145);
xor U9065 (N_9065,N_6397,N_6291);
and U9066 (N_9066,N_6538,N_6739);
or U9067 (N_9067,N_7991,N_6706);
nand U9068 (N_9068,N_7533,N_7247);
and U9069 (N_9069,N_6303,N_6172);
and U9070 (N_9070,N_6937,N_6331);
or U9071 (N_9071,N_7824,N_6454);
xor U9072 (N_9072,N_7887,N_6853);
or U9073 (N_9073,N_7758,N_6029);
nand U9074 (N_9074,N_7851,N_6315);
or U9075 (N_9075,N_6009,N_7638);
and U9076 (N_9076,N_7417,N_7139);
or U9077 (N_9077,N_7962,N_6492);
nor U9078 (N_9078,N_6614,N_6229);
and U9079 (N_9079,N_7464,N_6658);
or U9080 (N_9080,N_7047,N_6151);
or U9081 (N_9081,N_7232,N_6793);
or U9082 (N_9082,N_6121,N_7570);
and U9083 (N_9083,N_6424,N_6399);
nand U9084 (N_9084,N_7949,N_7590);
xor U9085 (N_9085,N_7365,N_6554);
and U9086 (N_9086,N_7038,N_7826);
nor U9087 (N_9087,N_7015,N_7089);
and U9088 (N_9088,N_7473,N_6559);
or U9089 (N_9089,N_7289,N_7652);
nand U9090 (N_9090,N_7259,N_6741);
nand U9091 (N_9091,N_6904,N_7985);
xnor U9092 (N_9092,N_6553,N_7806);
xnor U9093 (N_9093,N_7155,N_6646);
nor U9094 (N_9094,N_7431,N_6472);
nor U9095 (N_9095,N_7819,N_6748);
and U9096 (N_9096,N_7403,N_7222);
and U9097 (N_9097,N_6864,N_6835);
nor U9098 (N_9098,N_6735,N_7606);
xnor U9099 (N_9099,N_6341,N_6603);
xnor U9100 (N_9100,N_6681,N_6901);
xor U9101 (N_9101,N_7643,N_7095);
nor U9102 (N_9102,N_6620,N_6009);
nor U9103 (N_9103,N_6187,N_7484);
xor U9104 (N_9104,N_6160,N_7321);
nand U9105 (N_9105,N_7489,N_6450);
nor U9106 (N_9106,N_6542,N_7956);
nor U9107 (N_9107,N_6713,N_7644);
xor U9108 (N_9108,N_7620,N_7796);
and U9109 (N_9109,N_7916,N_7242);
or U9110 (N_9110,N_6452,N_7083);
xnor U9111 (N_9111,N_6624,N_6172);
or U9112 (N_9112,N_7499,N_7609);
or U9113 (N_9113,N_6598,N_6863);
nor U9114 (N_9114,N_6044,N_7619);
and U9115 (N_9115,N_7854,N_7809);
xor U9116 (N_9116,N_6783,N_6473);
or U9117 (N_9117,N_7015,N_7379);
nand U9118 (N_9118,N_6175,N_7459);
nor U9119 (N_9119,N_6202,N_6870);
nand U9120 (N_9120,N_6186,N_7853);
xnor U9121 (N_9121,N_6078,N_7875);
nand U9122 (N_9122,N_6947,N_7189);
nor U9123 (N_9123,N_7909,N_6924);
or U9124 (N_9124,N_7890,N_7066);
nand U9125 (N_9125,N_6654,N_6537);
nor U9126 (N_9126,N_7332,N_7822);
or U9127 (N_9127,N_7991,N_7487);
nand U9128 (N_9128,N_7424,N_6666);
nand U9129 (N_9129,N_7075,N_6534);
xnor U9130 (N_9130,N_6743,N_6018);
and U9131 (N_9131,N_7223,N_6486);
and U9132 (N_9132,N_7614,N_7125);
and U9133 (N_9133,N_7777,N_7125);
xor U9134 (N_9134,N_7168,N_7924);
and U9135 (N_9135,N_7671,N_6881);
or U9136 (N_9136,N_7388,N_6720);
xor U9137 (N_9137,N_7098,N_7647);
xnor U9138 (N_9138,N_6391,N_6467);
or U9139 (N_9139,N_7768,N_7138);
xnor U9140 (N_9140,N_7142,N_6058);
nand U9141 (N_9141,N_6864,N_7950);
nor U9142 (N_9142,N_7142,N_6389);
and U9143 (N_9143,N_6023,N_7058);
nand U9144 (N_9144,N_6269,N_7737);
nand U9145 (N_9145,N_7597,N_7150);
nand U9146 (N_9146,N_6049,N_7664);
and U9147 (N_9147,N_6332,N_7909);
nand U9148 (N_9148,N_6425,N_7021);
and U9149 (N_9149,N_6773,N_6699);
nor U9150 (N_9150,N_7006,N_7730);
xor U9151 (N_9151,N_6369,N_6326);
or U9152 (N_9152,N_7134,N_6847);
or U9153 (N_9153,N_7062,N_7914);
nand U9154 (N_9154,N_7982,N_6650);
or U9155 (N_9155,N_7872,N_6841);
nand U9156 (N_9156,N_6728,N_7770);
nand U9157 (N_9157,N_6304,N_6557);
and U9158 (N_9158,N_6442,N_7978);
nor U9159 (N_9159,N_6330,N_7770);
nor U9160 (N_9160,N_7614,N_7479);
nor U9161 (N_9161,N_6106,N_7872);
nand U9162 (N_9162,N_6337,N_6376);
nand U9163 (N_9163,N_6844,N_6231);
xor U9164 (N_9164,N_7482,N_7352);
nand U9165 (N_9165,N_7581,N_7633);
nand U9166 (N_9166,N_7191,N_6516);
and U9167 (N_9167,N_6334,N_7222);
or U9168 (N_9168,N_7857,N_7144);
xor U9169 (N_9169,N_7030,N_7023);
xor U9170 (N_9170,N_7770,N_6261);
and U9171 (N_9171,N_6218,N_7168);
or U9172 (N_9172,N_6514,N_6635);
xnor U9173 (N_9173,N_6120,N_6958);
and U9174 (N_9174,N_7768,N_6185);
nand U9175 (N_9175,N_7694,N_7409);
nand U9176 (N_9176,N_6952,N_7653);
xor U9177 (N_9177,N_6332,N_7043);
or U9178 (N_9178,N_7563,N_7270);
nand U9179 (N_9179,N_6138,N_6649);
and U9180 (N_9180,N_7750,N_6032);
nor U9181 (N_9181,N_6652,N_6005);
nand U9182 (N_9182,N_6890,N_7181);
nand U9183 (N_9183,N_7755,N_6299);
nand U9184 (N_9184,N_7768,N_7822);
xnor U9185 (N_9185,N_6991,N_7350);
xor U9186 (N_9186,N_7926,N_6510);
and U9187 (N_9187,N_7031,N_6767);
xnor U9188 (N_9188,N_6309,N_6293);
and U9189 (N_9189,N_7145,N_7758);
xnor U9190 (N_9190,N_6843,N_6756);
xnor U9191 (N_9191,N_7284,N_6602);
or U9192 (N_9192,N_7565,N_7501);
nand U9193 (N_9193,N_7310,N_7408);
and U9194 (N_9194,N_7799,N_7695);
xnor U9195 (N_9195,N_7578,N_6626);
or U9196 (N_9196,N_6442,N_6135);
nor U9197 (N_9197,N_7145,N_7680);
and U9198 (N_9198,N_7116,N_6437);
xnor U9199 (N_9199,N_7723,N_7752);
or U9200 (N_9200,N_6914,N_7936);
xnor U9201 (N_9201,N_7055,N_7069);
and U9202 (N_9202,N_7831,N_6280);
nand U9203 (N_9203,N_6201,N_7969);
nand U9204 (N_9204,N_6580,N_6562);
nor U9205 (N_9205,N_6701,N_6034);
nor U9206 (N_9206,N_6746,N_6446);
or U9207 (N_9207,N_6263,N_7973);
nor U9208 (N_9208,N_7816,N_6941);
or U9209 (N_9209,N_6538,N_6699);
and U9210 (N_9210,N_6513,N_7094);
nand U9211 (N_9211,N_7283,N_7932);
nand U9212 (N_9212,N_6640,N_6093);
nand U9213 (N_9213,N_7332,N_7725);
xnor U9214 (N_9214,N_7448,N_7261);
nand U9215 (N_9215,N_6450,N_7314);
or U9216 (N_9216,N_7059,N_6260);
and U9217 (N_9217,N_6909,N_7794);
xnor U9218 (N_9218,N_6969,N_7702);
xnor U9219 (N_9219,N_6545,N_6442);
nor U9220 (N_9220,N_7958,N_7709);
nor U9221 (N_9221,N_6244,N_7415);
and U9222 (N_9222,N_6510,N_7963);
nand U9223 (N_9223,N_6518,N_7458);
and U9224 (N_9224,N_7140,N_7221);
or U9225 (N_9225,N_6106,N_7352);
or U9226 (N_9226,N_6184,N_7086);
and U9227 (N_9227,N_7761,N_7527);
or U9228 (N_9228,N_6372,N_6206);
xor U9229 (N_9229,N_6354,N_6226);
or U9230 (N_9230,N_7878,N_6544);
nand U9231 (N_9231,N_6005,N_7392);
xor U9232 (N_9232,N_7741,N_7867);
nand U9233 (N_9233,N_7266,N_7333);
nand U9234 (N_9234,N_6523,N_7893);
nor U9235 (N_9235,N_7725,N_7637);
or U9236 (N_9236,N_7586,N_7224);
nor U9237 (N_9237,N_6701,N_7252);
nand U9238 (N_9238,N_7022,N_6221);
xnor U9239 (N_9239,N_6601,N_6524);
and U9240 (N_9240,N_6126,N_6373);
and U9241 (N_9241,N_7544,N_7701);
and U9242 (N_9242,N_6376,N_7156);
or U9243 (N_9243,N_6449,N_6353);
or U9244 (N_9244,N_7561,N_6791);
nand U9245 (N_9245,N_7991,N_6696);
nor U9246 (N_9246,N_7516,N_7405);
and U9247 (N_9247,N_7516,N_6977);
nor U9248 (N_9248,N_7747,N_7833);
xor U9249 (N_9249,N_6248,N_7051);
xnor U9250 (N_9250,N_7384,N_7235);
nor U9251 (N_9251,N_6194,N_6063);
or U9252 (N_9252,N_7442,N_6819);
and U9253 (N_9253,N_7077,N_7631);
and U9254 (N_9254,N_6867,N_7786);
xor U9255 (N_9255,N_7678,N_7693);
and U9256 (N_9256,N_7724,N_6504);
nor U9257 (N_9257,N_7909,N_7340);
nand U9258 (N_9258,N_7505,N_7594);
or U9259 (N_9259,N_6242,N_6523);
xor U9260 (N_9260,N_7965,N_6279);
nand U9261 (N_9261,N_7492,N_6264);
nor U9262 (N_9262,N_6794,N_6131);
nand U9263 (N_9263,N_6336,N_7969);
nand U9264 (N_9264,N_7755,N_6641);
and U9265 (N_9265,N_7761,N_6829);
and U9266 (N_9266,N_7970,N_7067);
or U9267 (N_9267,N_6946,N_6993);
nor U9268 (N_9268,N_6187,N_7606);
nor U9269 (N_9269,N_6621,N_6296);
or U9270 (N_9270,N_6028,N_7231);
or U9271 (N_9271,N_7795,N_7640);
and U9272 (N_9272,N_6548,N_7719);
and U9273 (N_9273,N_7451,N_6974);
nor U9274 (N_9274,N_7427,N_7415);
nor U9275 (N_9275,N_7303,N_7608);
nor U9276 (N_9276,N_6912,N_7691);
and U9277 (N_9277,N_7001,N_7671);
nand U9278 (N_9278,N_7698,N_6090);
and U9279 (N_9279,N_6650,N_6584);
nor U9280 (N_9280,N_7757,N_7589);
and U9281 (N_9281,N_6681,N_6611);
nor U9282 (N_9282,N_6142,N_7543);
and U9283 (N_9283,N_7198,N_7315);
nor U9284 (N_9284,N_6972,N_7975);
nand U9285 (N_9285,N_7771,N_6085);
nor U9286 (N_9286,N_6586,N_6163);
nor U9287 (N_9287,N_7554,N_6654);
or U9288 (N_9288,N_6249,N_6766);
xor U9289 (N_9289,N_6191,N_7535);
xor U9290 (N_9290,N_6020,N_7124);
and U9291 (N_9291,N_7651,N_6630);
and U9292 (N_9292,N_6836,N_6879);
and U9293 (N_9293,N_6269,N_6360);
and U9294 (N_9294,N_7700,N_6630);
nor U9295 (N_9295,N_7374,N_6913);
and U9296 (N_9296,N_6488,N_7030);
xor U9297 (N_9297,N_6942,N_7490);
or U9298 (N_9298,N_7795,N_7165);
or U9299 (N_9299,N_6129,N_7746);
nand U9300 (N_9300,N_6858,N_6872);
xnor U9301 (N_9301,N_7761,N_7445);
and U9302 (N_9302,N_6571,N_7142);
xnor U9303 (N_9303,N_7404,N_7770);
and U9304 (N_9304,N_6077,N_6268);
nor U9305 (N_9305,N_6812,N_7260);
nor U9306 (N_9306,N_6621,N_7056);
or U9307 (N_9307,N_6836,N_7210);
nor U9308 (N_9308,N_6249,N_7691);
or U9309 (N_9309,N_6598,N_7271);
nor U9310 (N_9310,N_7343,N_7404);
xor U9311 (N_9311,N_7469,N_6867);
xor U9312 (N_9312,N_6397,N_7996);
or U9313 (N_9313,N_6386,N_7019);
and U9314 (N_9314,N_7380,N_7783);
nor U9315 (N_9315,N_6949,N_6224);
xnor U9316 (N_9316,N_6253,N_6845);
nor U9317 (N_9317,N_6160,N_6639);
and U9318 (N_9318,N_7537,N_6508);
nor U9319 (N_9319,N_7750,N_7021);
nor U9320 (N_9320,N_6018,N_7773);
or U9321 (N_9321,N_7080,N_6576);
nor U9322 (N_9322,N_6836,N_6705);
or U9323 (N_9323,N_7547,N_6295);
nand U9324 (N_9324,N_6240,N_6420);
nand U9325 (N_9325,N_6044,N_7147);
or U9326 (N_9326,N_7297,N_7585);
nor U9327 (N_9327,N_6219,N_7244);
nor U9328 (N_9328,N_7681,N_6628);
xnor U9329 (N_9329,N_7592,N_7381);
or U9330 (N_9330,N_7041,N_7721);
nand U9331 (N_9331,N_7101,N_7439);
nor U9332 (N_9332,N_7123,N_7397);
and U9333 (N_9333,N_6552,N_6065);
nor U9334 (N_9334,N_6503,N_7118);
and U9335 (N_9335,N_7976,N_7229);
or U9336 (N_9336,N_7925,N_7533);
nand U9337 (N_9337,N_7601,N_7171);
nand U9338 (N_9338,N_6854,N_7846);
xor U9339 (N_9339,N_6643,N_7456);
or U9340 (N_9340,N_6470,N_7392);
and U9341 (N_9341,N_6403,N_7299);
or U9342 (N_9342,N_6456,N_6153);
nand U9343 (N_9343,N_7450,N_7346);
xor U9344 (N_9344,N_7410,N_7196);
nand U9345 (N_9345,N_7709,N_7112);
and U9346 (N_9346,N_6340,N_6702);
nor U9347 (N_9347,N_7758,N_6766);
or U9348 (N_9348,N_6209,N_6491);
and U9349 (N_9349,N_6440,N_6922);
nand U9350 (N_9350,N_6960,N_7434);
nor U9351 (N_9351,N_6007,N_7323);
nor U9352 (N_9352,N_6796,N_7239);
xor U9353 (N_9353,N_7224,N_6996);
and U9354 (N_9354,N_7606,N_6088);
or U9355 (N_9355,N_7100,N_7178);
nand U9356 (N_9356,N_6369,N_6436);
xnor U9357 (N_9357,N_7872,N_7584);
and U9358 (N_9358,N_6177,N_6302);
xor U9359 (N_9359,N_6955,N_6379);
xor U9360 (N_9360,N_6869,N_7344);
xnor U9361 (N_9361,N_6737,N_7231);
xnor U9362 (N_9362,N_7135,N_6837);
and U9363 (N_9363,N_6002,N_7664);
or U9364 (N_9364,N_7354,N_6581);
and U9365 (N_9365,N_6070,N_7350);
or U9366 (N_9366,N_6247,N_7946);
nand U9367 (N_9367,N_7986,N_7230);
xnor U9368 (N_9368,N_6707,N_7423);
xnor U9369 (N_9369,N_6097,N_6317);
nor U9370 (N_9370,N_7852,N_6858);
and U9371 (N_9371,N_6290,N_6242);
and U9372 (N_9372,N_7278,N_6217);
xnor U9373 (N_9373,N_6328,N_7074);
nor U9374 (N_9374,N_6061,N_7128);
or U9375 (N_9375,N_7283,N_6509);
and U9376 (N_9376,N_7105,N_7647);
xnor U9377 (N_9377,N_7111,N_7353);
xnor U9378 (N_9378,N_7549,N_6191);
or U9379 (N_9379,N_6234,N_7718);
or U9380 (N_9380,N_7991,N_7152);
nor U9381 (N_9381,N_6141,N_7286);
nor U9382 (N_9382,N_7001,N_6220);
xor U9383 (N_9383,N_7468,N_7177);
xor U9384 (N_9384,N_6129,N_6133);
or U9385 (N_9385,N_7607,N_6390);
xnor U9386 (N_9386,N_6424,N_6368);
or U9387 (N_9387,N_6878,N_7502);
nand U9388 (N_9388,N_7730,N_7559);
or U9389 (N_9389,N_7024,N_7290);
xnor U9390 (N_9390,N_6811,N_6138);
and U9391 (N_9391,N_7310,N_6913);
or U9392 (N_9392,N_7335,N_7495);
nand U9393 (N_9393,N_7822,N_7403);
xnor U9394 (N_9394,N_7698,N_6772);
nor U9395 (N_9395,N_7411,N_6840);
nor U9396 (N_9396,N_7758,N_7856);
nand U9397 (N_9397,N_6312,N_7474);
and U9398 (N_9398,N_6165,N_7282);
and U9399 (N_9399,N_7893,N_7508);
nand U9400 (N_9400,N_6828,N_7397);
xor U9401 (N_9401,N_7108,N_6392);
nand U9402 (N_9402,N_6286,N_7168);
nor U9403 (N_9403,N_6899,N_7255);
nand U9404 (N_9404,N_7150,N_7823);
and U9405 (N_9405,N_6369,N_7360);
nor U9406 (N_9406,N_7810,N_6608);
nand U9407 (N_9407,N_6314,N_6152);
nand U9408 (N_9408,N_6267,N_6386);
xnor U9409 (N_9409,N_7432,N_6678);
and U9410 (N_9410,N_6177,N_7654);
nand U9411 (N_9411,N_6964,N_6838);
nor U9412 (N_9412,N_7250,N_6276);
xnor U9413 (N_9413,N_6044,N_7723);
nor U9414 (N_9414,N_7015,N_7570);
or U9415 (N_9415,N_7644,N_6446);
and U9416 (N_9416,N_6824,N_6801);
xor U9417 (N_9417,N_6918,N_6206);
nor U9418 (N_9418,N_7782,N_6482);
xor U9419 (N_9419,N_7140,N_6126);
or U9420 (N_9420,N_7607,N_6407);
or U9421 (N_9421,N_6001,N_6268);
nor U9422 (N_9422,N_7422,N_6088);
xor U9423 (N_9423,N_7966,N_6551);
or U9424 (N_9424,N_7456,N_6339);
and U9425 (N_9425,N_7939,N_6331);
nand U9426 (N_9426,N_7571,N_7889);
and U9427 (N_9427,N_7403,N_6715);
or U9428 (N_9428,N_7870,N_7448);
or U9429 (N_9429,N_6159,N_7637);
or U9430 (N_9430,N_6699,N_7868);
and U9431 (N_9431,N_7078,N_7424);
nor U9432 (N_9432,N_7447,N_6558);
or U9433 (N_9433,N_6599,N_7260);
and U9434 (N_9434,N_6797,N_6383);
and U9435 (N_9435,N_7191,N_7111);
nand U9436 (N_9436,N_7563,N_6390);
and U9437 (N_9437,N_6518,N_6080);
nor U9438 (N_9438,N_6149,N_6784);
or U9439 (N_9439,N_7854,N_7551);
nand U9440 (N_9440,N_6344,N_6416);
nand U9441 (N_9441,N_7694,N_7878);
xor U9442 (N_9442,N_6608,N_7609);
nand U9443 (N_9443,N_7224,N_6058);
or U9444 (N_9444,N_7218,N_6994);
nand U9445 (N_9445,N_7953,N_7309);
and U9446 (N_9446,N_6733,N_6774);
nand U9447 (N_9447,N_7808,N_6364);
and U9448 (N_9448,N_7104,N_6260);
nand U9449 (N_9449,N_7242,N_6025);
nand U9450 (N_9450,N_6112,N_6386);
xnor U9451 (N_9451,N_6102,N_6243);
nand U9452 (N_9452,N_6010,N_6445);
or U9453 (N_9453,N_6497,N_6582);
and U9454 (N_9454,N_7507,N_6312);
nand U9455 (N_9455,N_6533,N_7564);
and U9456 (N_9456,N_7973,N_6373);
nor U9457 (N_9457,N_6420,N_7195);
and U9458 (N_9458,N_6308,N_6386);
nand U9459 (N_9459,N_7061,N_6758);
xnor U9460 (N_9460,N_6385,N_6352);
or U9461 (N_9461,N_6588,N_7570);
xnor U9462 (N_9462,N_7955,N_7891);
nand U9463 (N_9463,N_6583,N_7695);
xor U9464 (N_9464,N_6215,N_7334);
nor U9465 (N_9465,N_6891,N_7106);
nor U9466 (N_9466,N_7853,N_6397);
nand U9467 (N_9467,N_7612,N_6942);
or U9468 (N_9468,N_6070,N_6140);
nand U9469 (N_9469,N_7679,N_6035);
nor U9470 (N_9470,N_7297,N_6106);
xor U9471 (N_9471,N_7663,N_6738);
nor U9472 (N_9472,N_7046,N_6355);
nor U9473 (N_9473,N_7171,N_6227);
nor U9474 (N_9474,N_7811,N_7621);
xor U9475 (N_9475,N_7993,N_7885);
or U9476 (N_9476,N_6183,N_7598);
or U9477 (N_9477,N_6224,N_6779);
nor U9478 (N_9478,N_6216,N_7938);
and U9479 (N_9479,N_7201,N_7797);
nand U9480 (N_9480,N_6844,N_7241);
nand U9481 (N_9481,N_6600,N_6671);
or U9482 (N_9482,N_7499,N_7148);
nand U9483 (N_9483,N_7029,N_7558);
nand U9484 (N_9484,N_7562,N_7022);
and U9485 (N_9485,N_6578,N_6448);
or U9486 (N_9486,N_7143,N_7540);
or U9487 (N_9487,N_6417,N_6433);
or U9488 (N_9488,N_7497,N_7610);
nor U9489 (N_9489,N_7982,N_6995);
and U9490 (N_9490,N_6475,N_7469);
xor U9491 (N_9491,N_7251,N_7654);
nand U9492 (N_9492,N_7978,N_6085);
or U9493 (N_9493,N_6095,N_6782);
nor U9494 (N_9494,N_7801,N_7078);
nor U9495 (N_9495,N_6295,N_7762);
or U9496 (N_9496,N_6070,N_6230);
or U9497 (N_9497,N_7009,N_7423);
or U9498 (N_9498,N_6653,N_7433);
and U9499 (N_9499,N_7438,N_7719);
or U9500 (N_9500,N_7316,N_7783);
nand U9501 (N_9501,N_6630,N_7582);
or U9502 (N_9502,N_6566,N_6364);
nor U9503 (N_9503,N_7438,N_6756);
and U9504 (N_9504,N_6926,N_6067);
or U9505 (N_9505,N_7408,N_7347);
nand U9506 (N_9506,N_7285,N_6647);
nand U9507 (N_9507,N_6100,N_6799);
nand U9508 (N_9508,N_6062,N_6842);
or U9509 (N_9509,N_6660,N_6649);
nand U9510 (N_9510,N_6308,N_7139);
and U9511 (N_9511,N_6635,N_7479);
nand U9512 (N_9512,N_6355,N_6904);
nor U9513 (N_9513,N_7228,N_6104);
and U9514 (N_9514,N_7501,N_7273);
nor U9515 (N_9515,N_6872,N_6335);
or U9516 (N_9516,N_7468,N_6015);
nor U9517 (N_9517,N_7661,N_6693);
nand U9518 (N_9518,N_7752,N_6714);
xnor U9519 (N_9519,N_6586,N_6032);
nor U9520 (N_9520,N_6986,N_7271);
or U9521 (N_9521,N_7319,N_7496);
xor U9522 (N_9522,N_7205,N_7753);
xor U9523 (N_9523,N_6309,N_6175);
xor U9524 (N_9524,N_7555,N_6532);
xor U9525 (N_9525,N_7037,N_6945);
xor U9526 (N_9526,N_6043,N_7904);
nand U9527 (N_9527,N_6704,N_7002);
nor U9528 (N_9528,N_7116,N_7331);
nand U9529 (N_9529,N_6663,N_6159);
nor U9530 (N_9530,N_7562,N_6466);
and U9531 (N_9531,N_6850,N_7606);
nand U9532 (N_9532,N_7480,N_6986);
or U9533 (N_9533,N_7051,N_6061);
and U9534 (N_9534,N_7758,N_7700);
nand U9535 (N_9535,N_6535,N_7547);
and U9536 (N_9536,N_6881,N_6097);
or U9537 (N_9537,N_7792,N_7600);
and U9538 (N_9538,N_6115,N_6924);
or U9539 (N_9539,N_7240,N_7768);
or U9540 (N_9540,N_7769,N_7639);
xnor U9541 (N_9541,N_6738,N_7515);
and U9542 (N_9542,N_7924,N_7167);
and U9543 (N_9543,N_6860,N_6712);
nor U9544 (N_9544,N_6383,N_6863);
nor U9545 (N_9545,N_7328,N_7126);
nor U9546 (N_9546,N_6717,N_7022);
and U9547 (N_9547,N_6306,N_6375);
nand U9548 (N_9548,N_6835,N_7219);
nor U9549 (N_9549,N_6016,N_6303);
or U9550 (N_9550,N_7689,N_7808);
nand U9551 (N_9551,N_6641,N_7597);
nand U9552 (N_9552,N_7019,N_6571);
xor U9553 (N_9553,N_6130,N_6239);
nor U9554 (N_9554,N_7128,N_7108);
xor U9555 (N_9555,N_6054,N_7613);
and U9556 (N_9556,N_6794,N_7863);
and U9557 (N_9557,N_6390,N_7940);
or U9558 (N_9558,N_6418,N_7679);
nand U9559 (N_9559,N_7238,N_7629);
and U9560 (N_9560,N_6433,N_6121);
nor U9561 (N_9561,N_7731,N_6143);
xor U9562 (N_9562,N_6180,N_7219);
nor U9563 (N_9563,N_7116,N_7580);
nor U9564 (N_9564,N_6059,N_7291);
and U9565 (N_9565,N_6795,N_7600);
nand U9566 (N_9566,N_6772,N_6680);
and U9567 (N_9567,N_6259,N_7853);
or U9568 (N_9568,N_7318,N_6293);
xnor U9569 (N_9569,N_7477,N_6849);
xnor U9570 (N_9570,N_6073,N_6253);
nor U9571 (N_9571,N_6057,N_6294);
and U9572 (N_9572,N_7707,N_6295);
and U9573 (N_9573,N_7053,N_6863);
nor U9574 (N_9574,N_7184,N_7646);
nand U9575 (N_9575,N_6267,N_6321);
or U9576 (N_9576,N_6578,N_7176);
xnor U9577 (N_9577,N_7570,N_7830);
and U9578 (N_9578,N_7455,N_7331);
and U9579 (N_9579,N_6609,N_7238);
nor U9580 (N_9580,N_6268,N_7057);
or U9581 (N_9581,N_6564,N_6526);
or U9582 (N_9582,N_6987,N_7855);
or U9583 (N_9583,N_7913,N_7616);
or U9584 (N_9584,N_6163,N_7471);
or U9585 (N_9585,N_7726,N_7472);
xor U9586 (N_9586,N_6478,N_6379);
nand U9587 (N_9587,N_7666,N_7202);
and U9588 (N_9588,N_7871,N_6153);
and U9589 (N_9589,N_6200,N_7950);
nand U9590 (N_9590,N_6919,N_6430);
nand U9591 (N_9591,N_7420,N_7227);
xnor U9592 (N_9592,N_7635,N_6102);
or U9593 (N_9593,N_7386,N_6670);
nand U9594 (N_9594,N_6374,N_6543);
nand U9595 (N_9595,N_7667,N_7344);
nand U9596 (N_9596,N_7577,N_6013);
or U9597 (N_9597,N_6997,N_6866);
nand U9598 (N_9598,N_6523,N_6931);
xnor U9599 (N_9599,N_6980,N_6758);
nand U9600 (N_9600,N_6573,N_7059);
nor U9601 (N_9601,N_7087,N_6786);
xnor U9602 (N_9602,N_7563,N_6352);
nor U9603 (N_9603,N_7491,N_6249);
nor U9604 (N_9604,N_6493,N_7268);
nand U9605 (N_9605,N_6963,N_7934);
xor U9606 (N_9606,N_7557,N_6442);
nand U9607 (N_9607,N_6180,N_7144);
and U9608 (N_9608,N_7926,N_6271);
or U9609 (N_9609,N_7632,N_6253);
and U9610 (N_9610,N_6834,N_6606);
and U9611 (N_9611,N_7541,N_7753);
or U9612 (N_9612,N_7986,N_6598);
nor U9613 (N_9613,N_6256,N_6150);
nand U9614 (N_9614,N_7344,N_6650);
xnor U9615 (N_9615,N_7158,N_7508);
and U9616 (N_9616,N_7363,N_7343);
nor U9617 (N_9617,N_6945,N_6102);
nor U9618 (N_9618,N_6505,N_6028);
and U9619 (N_9619,N_7119,N_7147);
or U9620 (N_9620,N_7555,N_7323);
or U9621 (N_9621,N_7746,N_6419);
and U9622 (N_9622,N_6128,N_7701);
and U9623 (N_9623,N_7498,N_6981);
or U9624 (N_9624,N_6161,N_7988);
or U9625 (N_9625,N_6185,N_7920);
nor U9626 (N_9626,N_7166,N_6351);
nand U9627 (N_9627,N_6518,N_7138);
nand U9628 (N_9628,N_6760,N_7064);
xor U9629 (N_9629,N_6535,N_6262);
and U9630 (N_9630,N_7687,N_7810);
nor U9631 (N_9631,N_7644,N_6879);
nor U9632 (N_9632,N_7429,N_7033);
xnor U9633 (N_9633,N_6615,N_6337);
and U9634 (N_9634,N_6276,N_7652);
xor U9635 (N_9635,N_6837,N_7131);
xor U9636 (N_9636,N_7502,N_7387);
and U9637 (N_9637,N_7832,N_6981);
nor U9638 (N_9638,N_7597,N_6756);
nor U9639 (N_9639,N_6856,N_6839);
and U9640 (N_9640,N_6112,N_7317);
or U9641 (N_9641,N_6812,N_6481);
or U9642 (N_9642,N_6460,N_7548);
nor U9643 (N_9643,N_6474,N_7613);
nand U9644 (N_9644,N_6684,N_7762);
and U9645 (N_9645,N_7435,N_6904);
xor U9646 (N_9646,N_7956,N_7479);
or U9647 (N_9647,N_7396,N_6160);
nor U9648 (N_9648,N_7377,N_6431);
or U9649 (N_9649,N_7183,N_7402);
nand U9650 (N_9650,N_7642,N_6513);
nand U9651 (N_9651,N_7597,N_7190);
nand U9652 (N_9652,N_6827,N_6058);
and U9653 (N_9653,N_7833,N_7892);
xor U9654 (N_9654,N_7985,N_6358);
nor U9655 (N_9655,N_7692,N_6145);
nand U9656 (N_9656,N_7735,N_7081);
nor U9657 (N_9657,N_6989,N_7411);
nand U9658 (N_9658,N_7212,N_7795);
xnor U9659 (N_9659,N_6678,N_6895);
or U9660 (N_9660,N_6421,N_6879);
xnor U9661 (N_9661,N_6791,N_6585);
nand U9662 (N_9662,N_7796,N_7326);
xor U9663 (N_9663,N_6640,N_6804);
nor U9664 (N_9664,N_6170,N_7030);
nand U9665 (N_9665,N_7860,N_6075);
and U9666 (N_9666,N_6514,N_6769);
or U9667 (N_9667,N_6962,N_6220);
xnor U9668 (N_9668,N_7708,N_7000);
or U9669 (N_9669,N_6074,N_6447);
nand U9670 (N_9670,N_6273,N_7984);
or U9671 (N_9671,N_7103,N_6332);
nor U9672 (N_9672,N_6572,N_6235);
nor U9673 (N_9673,N_6880,N_7154);
nor U9674 (N_9674,N_7369,N_7651);
or U9675 (N_9675,N_6170,N_6083);
nor U9676 (N_9676,N_7738,N_6171);
nand U9677 (N_9677,N_6346,N_7657);
and U9678 (N_9678,N_7302,N_7398);
or U9679 (N_9679,N_7846,N_7325);
nor U9680 (N_9680,N_7569,N_6177);
xnor U9681 (N_9681,N_6031,N_7184);
or U9682 (N_9682,N_6048,N_6487);
or U9683 (N_9683,N_7684,N_7086);
and U9684 (N_9684,N_6222,N_7183);
nand U9685 (N_9685,N_6013,N_6471);
xor U9686 (N_9686,N_6498,N_7356);
nor U9687 (N_9687,N_7134,N_6459);
nor U9688 (N_9688,N_6259,N_6240);
nor U9689 (N_9689,N_7911,N_6397);
and U9690 (N_9690,N_7852,N_7303);
nand U9691 (N_9691,N_7985,N_6760);
and U9692 (N_9692,N_7200,N_6889);
nand U9693 (N_9693,N_7780,N_7323);
or U9694 (N_9694,N_7634,N_6865);
and U9695 (N_9695,N_7876,N_7232);
xnor U9696 (N_9696,N_6131,N_6388);
and U9697 (N_9697,N_6237,N_6659);
or U9698 (N_9698,N_7828,N_6261);
or U9699 (N_9699,N_6784,N_6911);
and U9700 (N_9700,N_7272,N_7098);
or U9701 (N_9701,N_6265,N_7218);
and U9702 (N_9702,N_6917,N_6709);
or U9703 (N_9703,N_6471,N_7439);
and U9704 (N_9704,N_6684,N_6727);
or U9705 (N_9705,N_7254,N_7982);
and U9706 (N_9706,N_7930,N_6893);
nand U9707 (N_9707,N_6082,N_7557);
nand U9708 (N_9708,N_6621,N_6261);
or U9709 (N_9709,N_6146,N_7042);
or U9710 (N_9710,N_7443,N_7063);
nand U9711 (N_9711,N_6774,N_7576);
xor U9712 (N_9712,N_6388,N_7567);
nand U9713 (N_9713,N_6584,N_6124);
xnor U9714 (N_9714,N_6801,N_7270);
xor U9715 (N_9715,N_7173,N_7685);
nor U9716 (N_9716,N_7879,N_6657);
nand U9717 (N_9717,N_6255,N_6694);
xor U9718 (N_9718,N_7732,N_6867);
nor U9719 (N_9719,N_6478,N_7535);
or U9720 (N_9720,N_7935,N_7642);
xnor U9721 (N_9721,N_7590,N_7264);
and U9722 (N_9722,N_7219,N_6044);
xor U9723 (N_9723,N_6628,N_7287);
or U9724 (N_9724,N_7071,N_6969);
nor U9725 (N_9725,N_7374,N_6053);
nor U9726 (N_9726,N_6464,N_6181);
and U9727 (N_9727,N_6149,N_6494);
or U9728 (N_9728,N_6224,N_7537);
and U9729 (N_9729,N_6288,N_6975);
nand U9730 (N_9730,N_7121,N_6519);
and U9731 (N_9731,N_6371,N_7779);
xor U9732 (N_9732,N_7723,N_7709);
nand U9733 (N_9733,N_7140,N_7767);
nor U9734 (N_9734,N_7952,N_6531);
or U9735 (N_9735,N_7391,N_7422);
nor U9736 (N_9736,N_7108,N_7373);
or U9737 (N_9737,N_6000,N_6291);
nor U9738 (N_9738,N_6067,N_6925);
and U9739 (N_9739,N_6148,N_6773);
xnor U9740 (N_9740,N_6233,N_7723);
nand U9741 (N_9741,N_7959,N_7409);
nor U9742 (N_9742,N_7308,N_7176);
xnor U9743 (N_9743,N_7772,N_7504);
or U9744 (N_9744,N_7785,N_7744);
nor U9745 (N_9745,N_6682,N_6458);
and U9746 (N_9746,N_7667,N_7910);
xor U9747 (N_9747,N_7061,N_7420);
nand U9748 (N_9748,N_6728,N_6878);
xor U9749 (N_9749,N_6574,N_7045);
xor U9750 (N_9750,N_7339,N_6164);
nor U9751 (N_9751,N_6779,N_6300);
xnor U9752 (N_9752,N_7447,N_6443);
nand U9753 (N_9753,N_6668,N_6119);
xnor U9754 (N_9754,N_6000,N_6369);
nor U9755 (N_9755,N_7559,N_7997);
and U9756 (N_9756,N_7268,N_7474);
xor U9757 (N_9757,N_7865,N_6260);
or U9758 (N_9758,N_6059,N_6362);
nor U9759 (N_9759,N_7489,N_6053);
and U9760 (N_9760,N_6399,N_7572);
nand U9761 (N_9761,N_6633,N_7864);
and U9762 (N_9762,N_7270,N_7669);
nor U9763 (N_9763,N_7446,N_7549);
nor U9764 (N_9764,N_7619,N_7770);
nand U9765 (N_9765,N_7380,N_6244);
and U9766 (N_9766,N_7949,N_6875);
nand U9767 (N_9767,N_7939,N_7185);
and U9768 (N_9768,N_7846,N_6511);
and U9769 (N_9769,N_7786,N_6537);
nor U9770 (N_9770,N_6636,N_7803);
nor U9771 (N_9771,N_7100,N_6524);
nand U9772 (N_9772,N_7993,N_6917);
or U9773 (N_9773,N_7474,N_7806);
xor U9774 (N_9774,N_7836,N_7753);
nand U9775 (N_9775,N_6483,N_7979);
nand U9776 (N_9776,N_6412,N_6930);
and U9777 (N_9777,N_7104,N_6914);
nand U9778 (N_9778,N_6159,N_6232);
nor U9779 (N_9779,N_7024,N_6184);
and U9780 (N_9780,N_7140,N_7937);
nand U9781 (N_9781,N_6248,N_6274);
and U9782 (N_9782,N_6324,N_7828);
and U9783 (N_9783,N_7490,N_7364);
xor U9784 (N_9784,N_7753,N_6201);
nand U9785 (N_9785,N_6575,N_6086);
and U9786 (N_9786,N_6948,N_7536);
xor U9787 (N_9787,N_7443,N_7077);
or U9788 (N_9788,N_6260,N_7274);
or U9789 (N_9789,N_7170,N_6714);
xnor U9790 (N_9790,N_6355,N_7183);
xor U9791 (N_9791,N_6009,N_6726);
and U9792 (N_9792,N_6019,N_7953);
or U9793 (N_9793,N_7440,N_6018);
nand U9794 (N_9794,N_6754,N_7656);
nand U9795 (N_9795,N_7451,N_7452);
or U9796 (N_9796,N_7527,N_7467);
nor U9797 (N_9797,N_7847,N_7495);
nor U9798 (N_9798,N_6026,N_6199);
nand U9799 (N_9799,N_7493,N_7735);
xor U9800 (N_9800,N_7738,N_7777);
and U9801 (N_9801,N_6234,N_6547);
or U9802 (N_9802,N_7148,N_6876);
nor U9803 (N_9803,N_6915,N_6309);
nand U9804 (N_9804,N_7169,N_6071);
nand U9805 (N_9805,N_7262,N_6253);
or U9806 (N_9806,N_7519,N_6867);
xnor U9807 (N_9807,N_7966,N_7036);
nor U9808 (N_9808,N_6027,N_7873);
nor U9809 (N_9809,N_7099,N_7660);
and U9810 (N_9810,N_7088,N_6771);
nand U9811 (N_9811,N_7034,N_6738);
xor U9812 (N_9812,N_7656,N_6159);
nand U9813 (N_9813,N_7870,N_6366);
nor U9814 (N_9814,N_6814,N_6111);
xnor U9815 (N_9815,N_7823,N_7841);
xnor U9816 (N_9816,N_6452,N_7246);
or U9817 (N_9817,N_6243,N_6065);
xor U9818 (N_9818,N_7134,N_6269);
and U9819 (N_9819,N_6154,N_7730);
or U9820 (N_9820,N_7494,N_7285);
xnor U9821 (N_9821,N_7744,N_6790);
nor U9822 (N_9822,N_6030,N_7146);
xor U9823 (N_9823,N_6164,N_6203);
and U9824 (N_9824,N_7081,N_7434);
or U9825 (N_9825,N_6864,N_7782);
nand U9826 (N_9826,N_6822,N_6939);
nor U9827 (N_9827,N_7006,N_6845);
or U9828 (N_9828,N_7075,N_7462);
nor U9829 (N_9829,N_7705,N_7124);
and U9830 (N_9830,N_6704,N_7596);
or U9831 (N_9831,N_7804,N_6626);
and U9832 (N_9832,N_6370,N_6543);
nand U9833 (N_9833,N_6385,N_7642);
or U9834 (N_9834,N_6705,N_7679);
xnor U9835 (N_9835,N_6474,N_6288);
or U9836 (N_9836,N_6962,N_7594);
and U9837 (N_9837,N_7765,N_6531);
and U9838 (N_9838,N_7890,N_7062);
nand U9839 (N_9839,N_7247,N_7133);
xor U9840 (N_9840,N_6863,N_6378);
nand U9841 (N_9841,N_7770,N_6393);
nor U9842 (N_9842,N_6920,N_7391);
nand U9843 (N_9843,N_7442,N_7793);
and U9844 (N_9844,N_6536,N_6663);
xor U9845 (N_9845,N_7710,N_7938);
nand U9846 (N_9846,N_7783,N_7612);
or U9847 (N_9847,N_6681,N_7559);
xor U9848 (N_9848,N_7046,N_6896);
nor U9849 (N_9849,N_7514,N_7168);
nor U9850 (N_9850,N_7559,N_6727);
or U9851 (N_9851,N_6815,N_6151);
nor U9852 (N_9852,N_7234,N_6883);
and U9853 (N_9853,N_6755,N_7757);
and U9854 (N_9854,N_6001,N_7157);
or U9855 (N_9855,N_7321,N_6203);
nor U9856 (N_9856,N_7612,N_7823);
nand U9857 (N_9857,N_6680,N_7147);
nand U9858 (N_9858,N_6686,N_7894);
nor U9859 (N_9859,N_7104,N_7033);
nor U9860 (N_9860,N_6929,N_7344);
xor U9861 (N_9861,N_7364,N_7223);
nand U9862 (N_9862,N_6463,N_7365);
and U9863 (N_9863,N_6759,N_7726);
nand U9864 (N_9864,N_7246,N_6991);
nand U9865 (N_9865,N_7907,N_6820);
nand U9866 (N_9866,N_7301,N_6906);
nor U9867 (N_9867,N_7125,N_6560);
nor U9868 (N_9868,N_7962,N_6520);
xnor U9869 (N_9869,N_6582,N_6303);
and U9870 (N_9870,N_6501,N_6436);
and U9871 (N_9871,N_7239,N_7574);
or U9872 (N_9872,N_7522,N_6763);
xnor U9873 (N_9873,N_6526,N_6441);
or U9874 (N_9874,N_6256,N_6113);
xor U9875 (N_9875,N_7195,N_7526);
xor U9876 (N_9876,N_7871,N_7751);
nor U9877 (N_9877,N_6495,N_7049);
nor U9878 (N_9878,N_7941,N_7243);
nand U9879 (N_9879,N_7035,N_6418);
nand U9880 (N_9880,N_6122,N_6118);
and U9881 (N_9881,N_7741,N_6151);
or U9882 (N_9882,N_7580,N_6570);
nor U9883 (N_9883,N_6268,N_7773);
and U9884 (N_9884,N_7056,N_6995);
or U9885 (N_9885,N_6752,N_7032);
xnor U9886 (N_9886,N_7432,N_6440);
and U9887 (N_9887,N_6152,N_6312);
or U9888 (N_9888,N_7425,N_7809);
and U9889 (N_9889,N_7603,N_6007);
xnor U9890 (N_9890,N_6325,N_7593);
nand U9891 (N_9891,N_7107,N_6491);
and U9892 (N_9892,N_6813,N_7944);
or U9893 (N_9893,N_6159,N_6119);
nor U9894 (N_9894,N_7379,N_6739);
nand U9895 (N_9895,N_6084,N_6175);
nand U9896 (N_9896,N_6696,N_6093);
nor U9897 (N_9897,N_7174,N_7684);
nand U9898 (N_9898,N_6217,N_7198);
nand U9899 (N_9899,N_7131,N_6558);
nor U9900 (N_9900,N_6391,N_7000);
and U9901 (N_9901,N_7453,N_6060);
nor U9902 (N_9902,N_7892,N_6734);
and U9903 (N_9903,N_7056,N_7996);
nand U9904 (N_9904,N_7291,N_7930);
nor U9905 (N_9905,N_6397,N_7405);
xnor U9906 (N_9906,N_7905,N_7095);
xnor U9907 (N_9907,N_6446,N_6692);
xor U9908 (N_9908,N_7765,N_6796);
nor U9909 (N_9909,N_6571,N_6973);
xnor U9910 (N_9910,N_7793,N_7802);
or U9911 (N_9911,N_7583,N_6366);
nand U9912 (N_9912,N_6078,N_7524);
xor U9913 (N_9913,N_6197,N_6890);
and U9914 (N_9914,N_7379,N_7778);
nor U9915 (N_9915,N_6081,N_6459);
and U9916 (N_9916,N_7240,N_7012);
and U9917 (N_9917,N_6185,N_6394);
nand U9918 (N_9918,N_7350,N_6085);
xnor U9919 (N_9919,N_7873,N_7224);
xnor U9920 (N_9920,N_7254,N_6234);
nand U9921 (N_9921,N_7608,N_7449);
nor U9922 (N_9922,N_6426,N_6955);
xnor U9923 (N_9923,N_6816,N_6690);
xnor U9924 (N_9924,N_7316,N_6577);
and U9925 (N_9925,N_7571,N_7044);
nor U9926 (N_9926,N_7459,N_6177);
xnor U9927 (N_9927,N_6923,N_7367);
nand U9928 (N_9928,N_7793,N_7287);
xor U9929 (N_9929,N_7200,N_6209);
nand U9930 (N_9930,N_6912,N_6873);
nor U9931 (N_9931,N_6483,N_6252);
xnor U9932 (N_9932,N_7685,N_7902);
and U9933 (N_9933,N_6504,N_7338);
or U9934 (N_9934,N_6380,N_7577);
xnor U9935 (N_9935,N_7327,N_7877);
or U9936 (N_9936,N_7110,N_6114);
nor U9937 (N_9937,N_7070,N_6037);
and U9938 (N_9938,N_6621,N_6186);
nand U9939 (N_9939,N_7612,N_7698);
xnor U9940 (N_9940,N_6475,N_6759);
and U9941 (N_9941,N_6831,N_7592);
and U9942 (N_9942,N_7593,N_6532);
nor U9943 (N_9943,N_7129,N_7959);
and U9944 (N_9944,N_7541,N_7253);
or U9945 (N_9945,N_7517,N_6952);
nand U9946 (N_9946,N_6719,N_7883);
nor U9947 (N_9947,N_7880,N_7050);
and U9948 (N_9948,N_7498,N_6598);
xor U9949 (N_9949,N_7318,N_6738);
xor U9950 (N_9950,N_7292,N_7442);
and U9951 (N_9951,N_6264,N_7294);
xnor U9952 (N_9952,N_7020,N_7391);
nor U9953 (N_9953,N_7474,N_7237);
xor U9954 (N_9954,N_6124,N_6173);
and U9955 (N_9955,N_7933,N_7620);
and U9956 (N_9956,N_6287,N_7300);
and U9957 (N_9957,N_6267,N_7812);
and U9958 (N_9958,N_7282,N_7680);
xor U9959 (N_9959,N_6689,N_6216);
nand U9960 (N_9960,N_6278,N_7968);
nor U9961 (N_9961,N_6020,N_7019);
xor U9962 (N_9962,N_7474,N_7330);
nand U9963 (N_9963,N_6057,N_7139);
xor U9964 (N_9964,N_7861,N_6710);
xnor U9965 (N_9965,N_7978,N_7845);
nand U9966 (N_9966,N_6895,N_7130);
nand U9967 (N_9967,N_6922,N_6039);
nand U9968 (N_9968,N_6783,N_6313);
nor U9969 (N_9969,N_7144,N_6146);
or U9970 (N_9970,N_6453,N_6320);
and U9971 (N_9971,N_6740,N_6610);
nor U9972 (N_9972,N_6214,N_6879);
xnor U9973 (N_9973,N_7435,N_7039);
and U9974 (N_9974,N_6413,N_7766);
or U9975 (N_9975,N_6993,N_7263);
xnor U9976 (N_9976,N_6031,N_7078);
and U9977 (N_9977,N_6132,N_6740);
xnor U9978 (N_9978,N_7441,N_6236);
nor U9979 (N_9979,N_7293,N_7994);
xnor U9980 (N_9980,N_7344,N_7135);
and U9981 (N_9981,N_7298,N_6137);
nand U9982 (N_9982,N_7846,N_7725);
and U9983 (N_9983,N_6551,N_6918);
xor U9984 (N_9984,N_7429,N_7541);
xnor U9985 (N_9985,N_6321,N_6125);
and U9986 (N_9986,N_6982,N_6006);
nor U9987 (N_9987,N_6838,N_6747);
xnor U9988 (N_9988,N_6181,N_7992);
xnor U9989 (N_9989,N_6630,N_6855);
nor U9990 (N_9990,N_7825,N_6771);
or U9991 (N_9991,N_7180,N_7351);
or U9992 (N_9992,N_6826,N_6509);
and U9993 (N_9993,N_6836,N_7410);
nor U9994 (N_9994,N_6717,N_6422);
xnor U9995 (N_9995,N_6633,N_7033);
xor U9996 (N_9996,N_6428,N_7145);
xnor U9997 (N_9997,N_6049,N_6694);
nand U9998 (N_9998,N_7214,N_7751);
xnor U9999 (N_9999,N_6268,N_6430);
nor U10000 (N_10000,N_9299,N_9282);
nand U10001 (N_10001,N_9012,N_8612);
or U10002 (N_10002,N_8012,N_8502);
xor U10003 (N_10003,N_8275,N_8062);
nand U10004 (N_10004,N_9937,N_9710);
nand U10005 (N_10005,N_9560,N_9641);
nor U10006 (N_10006,N_8183,N_9973);
nor U10007 (N_10007,N_9956,N_9201);
or U10008 (N_10008,N_9343,N_8703);
xor U10009 (N_10009,N_8604,N_8425);
and U10010 (N_10010,N_9346,N_9608);
and U10011 (N_10011,N_9593,N_9393);
or U10012 (N_10012,N_8319,N_9635);
nand U10013 (N_10013,N_9403,N_9506);
and U10014 (N_10014,N_8130,N_8462);
and U10015 (N_10015,N_9578,N_8761);
or U10016 (N_10016,N_8261,N_8938);
or U10017 (N_10017,N_8980,N_9002);
nand U10018 (N_10018,N_9888,N_8246);
and U10019 (N_10019,N_9048,N_8005);
or U10020 (N_10020,N_8890,N_8335);
xnor U10021 (N_10021,N_8811,N_9075);
xnor U10022 (N_10022,N_8599,N_8777);
nor U10023 (N_10023,N_9337,N_9032);
and U10024 (N_10024,N_9358,N_8251);
or U10025 (N_10025,N_8635,N_9064);
nand U10026 (N_10026,N_8067,N_8881);
xnor U10027 (N_10027,N_9893,N_9111);
nand U10028 (N_10028,N_8239,N_9312);
xor U10029 (N_10029,N_9263,N_9985);
or U10030 (N_10030,N_8792,N_9689);
nand U10031 (N_10031,N_9160,N_9394);
or U10032 (N_10032,N_8467,N_9638);
xor U10033 (N_10033,N_8954,N_8033);
nor U10034 (N_10034,N_9601,N_9600);
and U10035 (N_10035,N_8059,N_8390);
or U10036 (N_10036,N_8464,N_9882);
and U10037 (N_10037,N_9826,N_8798);
and U10038 (N_10038,N_8397,N_8747);
nor U10039 (N_10039,N_8073,N_8273);
and U10040 (N_10040,N_8822,N_9382);
nand U10041 (N_10041,N_9930,N_8258);
xnor U10042 (N_10042,N_8541,N_9784);
nand U10043 (N_10043,N_8169,N_9490);
xnor U10044 (N_10044,N_9069,N_8816);
nand U10045 (N_10045,N_9190,N_9361);
nor U10046 (N_10046,N_9768,N_8308);
nand U10047 (N_10047,N_8937,N_9468);
and U10048 (N_10048,N_8374,N_9141);
nand U10049 (N_10049,N_9325,N_9106);
or U10050 (N_10050,N_9955,N_8297);
and U10051 (N_10051,N_8671,N_8241);
and U10052 (N_10052,N_9505,N_9721);
xor U10053 (N_10053,N_9860,N_8440);
nor U10054 (N_10054,N_8368,N_9744);
or U10055 (N_10055,N_9268,N_8101);
nor U10056 (N_10056,N_9835,N_8447);
or U10057 (N_10057,N_8933,N_9166);
nand U10058 (N_10058,N_9034,N_9712);
xor U10059 (N_10059,N_9293,N_8334);
nand U10060 (N_10060,N_9483,N_8842);
nand U10061 (N_10061,N_9953,N_8354);
nor U10062 (N_10062,N_8892,N_8564);
or U10063 (N_10063,N_8164,N_8090);
xor U10064 (N_10064,N_8898,N_8883);
or U10065 (N_10065,N_9199,N_8548);
nand U10066 (N_10066,N_9253,N_8158);
nor U10067 (N_10067,N_8787,N_9179);
and U10068 (N_10068,N_9339,N_8204);
xor U10069 (N_10069,N_9651,N_8605);
and U10070 (N_10070,N_8365,N_9197);
xnor U10071 (N_10071,N_9234,N_9997);
xor U10072 (N_10072,N_8807,N_8106);
xor U10073 (N_10073,N_8518,N_9847);
and U10074 (N_10074,N_9340,N_8831);
and U10075 (N_10075,N_8270,N_9598);
nand U10076 (N_10076,N_9760,N_9836);
and U10077 (N_10077,N_8461,N_9164);
nand U10078 (N_10078,N_9728,N_9516);
or U10079 (N_10079,N_9866,N_8056);
nand U10080 (N_10080,N_8810,N_9103);
nor U10081 (N_10081,N_8233,N_9925);
nor U10082 (N_10082,N_8125,N_8473);
and U10083 (N_10083,N_8602,N_8855);
nand U10084 (N_10084,N_8439,N_8424);
xnor U10085 (N_10085,N_8338,N_9515);
and U10086 (N_10086,N_8290,N_8885);
nor U10087 (N_10087,N_8804,N_8770);
and U10088 (N_10088,N_9513,N_8267);
nor U10089 (N_10089,N_8459,N_9162);
and U10090 (N_10090,N_9135,N_9238);
xor U10091 (N_10091,N_8003,N_8438);
xnor U10092 (N_10092,N_8510,N_8597);
xor U10093 (N_10093,N_8946,N_9846);
nand U10094 (N_10094,N_9306,N_9862);
or U10095 (N_10095,N_9999,N_8663);
xor U10096 (N_10096,N_9390,N_9143);
or U10097 (N_10097,N_9399,N_8555);
nor U10098 (N_10098,N_8725,N_8401);
and U10099 (N_10099,N_9745,N_8880);
nand U10100 (N_10100,N_8114,N_8790);
xor U10101 (N_10101,N_9616,N_9709);
or U10102 (N_10102,N_9964,N_8958);
and U10103 (N_10103,N_9184,N_8395);
nand U10104 (N_10104,N_8480,N_9633);
nand U10105 (N_10105,N_8847,N_9706);
nand U10106 (N_10106,N_9518,N_9020);
and U10107 (N_10107,N_8908,N_9491);
and U10108 (N_10108,N_8330,N_9961);
and U10109 (N_10109,N_8601,N_8455);
and U10110 (N_10110,N_8017,N_8861);
nor U10111 (N_10111,N_8607,N_9574);
and U10112 (N_10112,N_8317,N_8479);
nor U10113 (N_10113,N_8384,N_8626);
xnor U10114 (N_10114,N_8252,N_8208);
nor U10115 (N_10115,N_9829,N_9137);
nand U10116 (N_10116,N_9503,N_8926);
xor U10117 (N_10117,N_9752,N_8497);
xnor U10118 (N_10118,N_8882,N_9100);
or U10119 (N_10119,N_9940,N_9704);
or U10120 (N_10120,N_8491,N_8965);
nand U10121 (N_10121,N_8736,N_9645);
nand U10122 (N_10122,N_8347,N_9440);
nand U10123 (N_10123,N_8194,N_9548);
and U10124 (N_10124,N_9045,N_9051);
xnor U10125 (N_10125,N_9039,N_9705);
or U10126 (N_10126,N_9279,N_8760);
nand U10127 (N_10127,N_8919,N_9521);
or U10128 (N_10128,N_8232,N_8595);
or U10129 (N_10129,N_9605,N_8474);
and U10130 (N_10130,N_8535,N_8503);
xnor U10131 (N_10131,N_8051,N_9001);
nand U10132 (N_10132,N_9031,N_8360);
or U10133 (N_10133,N_9566,N_9392);
nand U10134 (N_10134,N_9102,N_9428);
or U10135 (N_10135,N_9384,N_9804);
nand U10136 (N_10136,N_8746,N_8293);
nand U10137 (N_10137,N_8469,N_9292);
xnor U10138 (N_10138,N_9624,N_9758);
nor U10139 (N_10139,N_8292,N_8490);
xnor U10140 (N_10140,N_9195,N_9870);
nor U10141 (N_10141,N_9854,N_8206);
xor U10142 (N_10142,N_8123,N_9932);
or U10143 (N_10143,N_8930,N_9599);
nand U10144 (N_10144,N_9063,N_9678);
nand U10145 (N_10145,N_8442,N_8572);
xor U10146 (N_10146,N_9708,N_8435);
xnor U10147 (N_10147,N_9900,N_9910);
xnor U10148 (N_10148,N_9404,N_8098);
xnor U10149 (N_10149,N_9167,N_9542);
or U10150 (N_10150,N_8421,N_8304);
nand U10151 (N_10151,N_8887,N_8496);
or U10152 (N_10152,N_9747,N_8013);
and U10153 (N_10153,N_8551,N_9919);
xnor U10154 (N_10154,N_8333,N_9058);
and U10155 (N_10155,N_8507,N_8078);
nand U10156 (N_10156,N_8515,N_9298);
or U10157 (N_10157,N_9014,N_8296);
nand U10158 (N_10158,N_8225,N_9591);
nand U10159 (N_10159,N_9099,N_9732);
or U10160 (N_10160,N_8398,N_9280);
xor U10161 (N_10161,N_9356,N_9650);
xnor U10162 (N_10162,N_9785,N_8534);
nand U10163 (N_10163,N_8314,N_9996);
and U10164 (N_10164,N_8007,N_8137);
nor U10165 (N_10165,N_8744,N_8618);
nand U10166 (N_10166,N_8077,N_8035);
xor U10167 (N_10167,N_9916,N_8878);
nand U10168 (N_10168,N_9969,N_9381);
and U10169 (N_10169,N_8756,N_9363);
or U10170 (N_10170,N_8237,N_9774);
nor U10171 (N_10171,N_9266,N_9439);
or U10172 (N_10172,N_8951,N_9296);
nand U10173 (N_10173,N_8886,N_8594);
or U10174 (N_10174,N_9791,N_9350);
and U10175 (N_10175,N_9487,N_9083);
nand U10176 (N_10176,N_9848,N_9669);
nand U10177 (N_10177,N_8672,N_8524);
xor U10178 (N_10178,N_8531,N_9530);
nand U10179 (N_10179,N_9289,N_9587);
and U10180 (N_10180,N_9070,N_8924);
xor U10181 (N_10181,N_9278,N_9686);
nand U10182 (N_10182,N_8606,N_9733);
and U10183 (N_10183,N_8287,N_8231);
xnor U10184 (N_10184,N_9093,N_9006);
xnor U10185 (N_10185,N_9005,N_8034);
nor U10186 (N_10186,N_8321,N_8363);
xor U10187 (N_10187,N_8656,N_9746);
or U10188 (N_10188,N_8916,N_8876);
and U10189 (N_10189,N_8378,N_8889);
nor U10190 (N_10190,N_8274,N_8103);
xnor U10191 (N_10191,N_8543,N_8433);
or U10192 (N_10192,N_8493,N_9713);
xnor U10193 (N_10193,N_8817,N_9833);
nor U10194 (N_10194,N_9907,N_8848);
nor U10195 (N_10195,N_9693,N_9665);
and U10196 (N_10196,N_9484,N_8661);
and U10197 (N_10197,N_8339,N_8533);
xor U10198 (N_10198,N_9896,N_9016);
or U10199 (N_10199,N_9975,N_9823);
or U10200 (N_10200,N_8131,N_9522);
and U10201 (N_10201,N_9569,N_8973);
or U10202 (N_10202,N_9396,N_9986);
and U10203 (N_10203,N_9189,N_9938);
xnor U10204 (N_10204,N_8836,N_9323);
or U10205 (N_10205,N_8687,N_8808);
nand U10206 (N_10206,N_8598,N_8659);
nor U10207 (N_10207,N_8870,N_9239);
or U10208 (N_10208,N_8961,N_9628);
nand U10209 (N_10209,N_9287,N_9853);
nand U10210 (N_10210,N_9105,N_8990);
and U10211 (N_10211,N_9313,N_8040);
nor U10212 (N_10212,N_9764,N_8662);
xor U10213 (N_10213,N_9783,N_9376);
xor U10214 (N_10214,N_9407,N_9088);
or U10215 (N_10215,N_8085,N_8104);
or U10216 (N_10216,N_8228,N_9030);
or U10217 (N_10217,N_9004,N_8568);
or U10218 (N_10218,N_8868,N_8453);
or U10219 (N_10219,N_9442,N_9364);
nor U10220 (N_10220,N_9885,N_8132);
nand U10221 (N_10221,N_9305,N_9327);
xor U10222 (N_10222,N_9463,N_9801);
and U10223 (N_10223,N_8146,N_9556);
or U10224 (N_10224,N_9772,N_8858);
xor U10225 (N_10225,N_8843,N_9884);
xor U10226 (N_10226,N_9723,N_9603);
or U10227 (N_10227,N_9540,N_9345);
and U10228 (N_10228,N_8043,N_9320);
xor U10229 (N_10229,N_8942,N_9731);
nor U10230 (N_10230,N_8920,N_8818);
and U10231 (N_10231,N_9617,N_8238);
nand U10232 (N_10232,N_8782,N_8501);
nor U10233 (N_10233,N_9497,N_8837);
or U10234 (N_10234,N_9615,N_9037);
nor U10235 (N_10235,N_9149,N_9450);
xnor U10236 (N_10236,N_9228,N_9445);
or U10237 (N_10237,N_9262,N_9013);
and U10238 (N_10238,N_8295,N_8018);
and U10239 (N_10239,N_9061,N_8648);
nand U10240 (N_10240,N_8989,N_9080);
nand U10241 (N_10241,N_8445,N_8224);
xor U10242 (N_10242,N_9691,N_9104);
xnor U10243 (N_10243,N_9684,N_8888);
or U10244 (N_10244,N_8751,N_8812);
xor U10245 (N_10245,N_9073,N_8563);
xor U10246 (N_10246,N_9794,N_9694);
or U10247 (N_10247,N_9604,N_9679);
xor U10248 (N_10248,N_9511,N_8617);
or U10249 (N_10249,N_9010,N_9789);
xor U10250 (N_10250,N_8894,N_9269);
and U10251 (N_10251,N_8097,N_8190);
and U10252 (N_10252,N_8879,N_8021);
nor U10253 (N_10253,N_9057,N_8336);
or U10254 (N_10254,N_9215,N_8576);
nand U10255 (N_10255,N_9056,N_9673);
or U10256 (N_10256,N_9495,N_9003);
or U10257 (N_10257,N_8715,N_8799);
xnor U10258 (N_10258,N_9781,N_8466);
nor U10259 (N_10259,N_9811,N_8081);
nor U10260 (N_10260,N_8695,N_9580);
and U10261 (N_10261,N_9901,N_9116);
xnor U10262 (N_10262,N_9478,N_8630);
nand U10263 (N_10263,N_8209,N_9682);
xor U10264 (N_10264,N_8849,N_9295);
or U10265 (N_10265,N_8144,N_9276);
nor U10266 (N_10266,N_9748,N_9216);
and U10267 (N_10267,N_9523,N_8823);
nor U10268 (N_10268,N_8762,N_9182);
nand U10269 (N_10269,N_9720,N_9391);
or U10270 (N_10270,N_9769,N_9437);
nand U10271 (N_10271,N_8446,N_9231);
nor U10272 (N_10272,N_8558,N_9881);
and U10273 (N_10273,N_9777,N_8122);
or U10274 (N_10274,N_8596,N_9904);
and U10275 (N_10275,N_9634,N_8159);
nor U10276 (N_10276,N_8119,N_9147);
and U10277 (N_10277,N_8934,N_8872);
xnor U10278 (N_10278,N_8147,N_8982);
nand U10279 (N_10279,N_8484,N_9368);
nand U10280 (N_10280,N_8839,N_9512);
or U10281 (N_10281,N_9419,N_9606);
or U10282 (N_10282,N_8245,N_9692);
or U10283 (N_10283,N_8136,N_9802);
xnor U10284 (N_10284,N_8773,N_8824);
and U10285 (N_10285,N_9328,N_8352);
nor U10286 (N_10286,N_9741,N_9547);
xnor U10287 (N_10287,N_9819,N_8904);
or U10288 (N_10288,N_8504,N_8896);
nand U10289 (N_10289,N_8302,N_8305);
nor U10290 (N_10290,N_8320,N_8544);
or U10291 (N_10291,N_9755,N_8629);
nor U10292 (N_10292,N_9475,N_8083);
or U10293 (N_10293,N_8996,N_8701);
nor U10294 (N_10294,N_9157,N_9387);
and U10295 (N_10295,N_8436,N_8652);
or U10296 (N_10296,N_9563,N_8577);
or U10297 (N_10297,N_9869,N_9214);
and U10298 (N_10298,N_9089,N_8181);
xnor U10299 (N_10299,N_9433,N_9132);
nor U10300 (N_10300,N_8884,N_9845);
or U10301 (N_10301,N_9824,N_8070);
or U10302 (N_10302,N_8223,N_8102);
and U10303 (N_10303,N_9400,N_9409);
nor U10304 (N_10304,N_8399,N_8774);
nor U10305 (N_10305,N_8328,N_8082);
and U10306 (N_10306,N_9595,N_8430);
xnor U10307 (N_10307,N_8364,N_8023);
nand U10308 (N_10308,N_9378,N_9696);
nand U10309 (N_10309,N_9960,N_9229);
nor U10310 (N_10310,N_9859,N_8180);
and U10311 (N_10311,N_8367,N_8264);
or U10312 (N_10312,N_8278,N_8707);
or U10313 (N_10313,N_8192,N_9922);
nand U10314 (N_10314,N_8277,N_9575);
xor U10315 (N_10315,N_9294,N_9796);
xor U10316 (N_10316,N_8111,N_8240);
or U10317 (N_10317,N_9174,N_8341);
xor U10318 (N_10318,N_9561,N_8443);
nand U10319 (N_10319,N_8387,N_8720);
xor U10320 (N_10320,N_8113,N_9555);
nor U10321 (N_10321,N_9637,N_8488);
or U10322 (N_10322,N_9485,N_8814);
and U10323 (N_10323,N_8813,N_8706);
and U10324 (N_10324,N_9441,N_9492);
nor U10325 (N_10325,N_9719,N_9386);
or U10326 (N_10326,N_8199,N_9993);
xnor U10327 (N_10327,N_8451,N_8570);
or U10328 (N_10328,N_9762,N_8344);
or U10329 (N_10329,N_9590,N_8897);
nand U10330 (N_10330,N_8500,N_8668);
nand U10331 (N_10331,N_8684,N_8422);
nand U10332 (N_10332,N_8120,N_8259);
nand U10333 (N_10333,N_8366,N_8348);
or U10334 (N_10334,N_8895,N_8355);
xor U10335 (N_10335,N_8255,N_8554);
nor U10336 (N_10336,N_9357,N_9979);
or U10337 (N_10337,N_8681,N_9281);
or U10338 (N_10338,N_8521,N_9607);
xnor U10339 (N_10339,N_8693,N_8699);
or U10340 (N_10340,N_8143,N_8586);
and U10341 (N_10341,N_8875,N_8080);
and U10342 (N_10342,N_9610,N_8910);
or U10343 (N_10343,N_9009,N_8647);
nand U10344 (N_10344,N_8903,N_8389);
and U10345 (N_10345,N_8786,N_9086);
nor U10346 (N_10346,N_9864,N_9308);
or U10347 (N_10347,N_9488,N_8195);
and U10348 (N_10348,N_9314,N_8441);
nand U10349 (N_10349,N_9486,N_8528);
xor U10350 (N_10350,N_9942,N_9571);
nor U10351 (N_10351,N_9277,N_8189);
nor U10352 (N_10352,N_9177,N_8417);
nand U10353 (N_10353,N_9476,N_9092);
nor U10354 (N_10354,N_9798,N_9360);
nor U10355 (N_10355,N_8306,N_8685);
nand U10356 (N_10356,N_8283,N_9886);
and U10357 (N_10357,N_8394,N_8514);
nor U10358 (N_10358,N_9291,N_9788);
nand U10359 (N_10359,N_8712,N_8509);
or U10360 (N_10360,N_8832,N_9676);
xor U10361 (N_10361,N_8863,N_8205);
nand U10362 (N_10362,N_8489,N_9987);
or U10363 (N_10363,N_9941,N_9221);
or U10364 (N_10364,N_8001,N_8625);
nor U10365 (N_10365,N_8105,N_9931);
and U10366 (N_10366,N_8675,N_9108);
nand U10367 (N_10367,N_8212,N_9156);
nor U10368 (N_10368,N_8037,N_8669);
nand U10369 (N_10369,N_8505,N_9427);
nand U10370 (N_10370,N_9423,N_8976);
and U10371 (N_10371,N_9420,N_8769);
nor U10372 (N_10372,N_9481,N_9098);
or U10373 (N_10373,N_8767,N_9572);
and U10374 (N_10374,N_8830,N_8950);
nand U10375 (N_10375,N_9243,N_8312);
xnor U10376 (N_10376,N_8128,N_9027);
nand U10377 (N_10377,N_9145,N_9648);
nand U10378 (N_10378,N_9352,N_8207);
or U10379 (N_10379,N_9218,N_9892);
xor U10380 (N_10380,N_9366,N_9480);
and U10381 (N_10381,N_8643,N_9677);
or U10382 (N_10382,N_8028,N_9401);
xor U10383 (N_10383,N_8250,N_8187);
and U10384 (N_10384,N_9568,N_9303);
nand U10385 (N_10385,N_8135,N_8853);
nor U10386 (N_10386,N_9347,N_9991);
or U10387 (N_10387,N_9341,N_8115);
xor U10388 (N_10388,N_9954,N_8527);
xor U10389 (N_10389,N_8310,N_9756);
nor U10390 (N_10390,N_8415,N_9059);
or U10391 (N_10391,N_8867,N_8030);
nor U10392 (N_10392,N_9438,N_9096);
nor U10393 (N_10393,N_9271,N_9510);
nand U10394 (N_10394,N_8550,N_9091);
xor U10395 (N_10395,N_9715,N_9256);
or U10396 (N_10396,N_8449,N_8616);
or U10397 (N_10397,N_9933,N_8846);
or U10398 (N_10398,N_9545,N_9496);
nor U10399 (N_10399,N_8957,N_9178);
or U10400 (N_10400,N_8175,N_8027);
or U10401 (N_10401,N_9793,N_8765);
nor U10402 (N_10402,N_8286,N_8713);
and U10403 (N_10403,N_9119,N_9342);
xnor U10404 (N_10404,N_8385,N_8351);
or U10405 (N_10405,N_9071,N_9799);
or U10406 (N_10406,N_9222,N_8188);
nor U10407 (N_10407,N_8088,N_8949);
nor U10408 (N_10408,N_8191,N_8121);
and U10409 (N_10409,N_9735,N_8087);
xor U10410 (N_10410,N_9553,N_8580);
nor U10411 (N_10411,N_8414,N_9375);
xnor U10412 (N_10412,N_9716,N_8815);
nor U10413 (N_10413,N_9994,N_9385);
nor U10414 (N_10414,N_9434,N_9537);
nand U10415 (N_10415,N_8176,N_9332);
xnor U10416 (N_10416,N_9115,N_8517);
and U10417 (N_10417,N_8561,N_9127);
xnor U10418 (N_10418,N_8029,N_9326);
and U10419 (N_10419,N_9773,N_9584);
or U10420 (N_10420,N_8112,N_9274);
or U10421 (N_10421,N_8731,N_8047);
and U10422 (N_10422,N_8906,N_9915);
xor U10423 (N_10423,N_8962,N_8089);
xor U10424 (N_10424,N_9597,N_9176);
xor U10425 (N_10425,N_8069,N_8827);
nand U10426 (N_10426,N_9068,N_8741);
nand U10427 (N_10427,N_8257,N_9072);
or U10428 (N_10428,N_9626,N_9751);
and U10429 (N_10429,N_8150,N_9579);
nor U10430 (N_10430,N_8780,N_9133);
xor U10431 (N_10431,N_9588,N_9398);
or U10432 (N_10432,N_8755,N_9675);
nor U10433 (N_10433,N_8107,N_9778);
or U10434 (N_10434,N_8649,N_9525);
and U10435 (N_10435,N_8752,N_8862);
nor U10436 (N_10436,N_8281,N_8981);
xnor U10437 (N_10437,N_8271,N_8032);
or U10438 (N_10438,N_8757,N_8410);
xor U10439 (N_10439,N_9672,N_8009);
nor U10440 (N_10440,N_9021,N_8710);
and U10441 (N_10441,N_8022,N_8392);
xor U10442 (N_10442,N_9895,N_8728);
or U10443 (N_10443,N_8722,N_8019);
nand U10444 (N_10444,N_9657,N_8763);
and U10445 (N_10445,N_8569,N_9464);
nor U10446 (N_10446,N_9336,N_8809);
nand U10447 (N_10447,N_8840,N_8860);
nand U10448 (N_10448,N_9015,N_9454);
nor U10449 (N_10449,N_9078,N_9539);
and U10450 (N_10450,N_9887,N_8641);
or U10451 (N_10451,N_8260,N_9165);
or U10452 (N_10452,N_9204,N_9154);
and U10453 (N_10453,N_9408,N_9087);
xor U10454 (N_10454,N_9144,N_8519);
nor U10455 (N_10455,N_9319,N_9499);
nand U10456 (N_10456,N_9532,N_8127);
and U10457 (N_10457,N_8468,N_8494);
or U10458 (N_10458,N_8382,N_9620);
or U10459 (N_10459,N_8579,N_8075);
or U10460 (N_10460,N_9076,N_8393);
nor U10461 (N_10461,N_8476,N_8915);
nor U10462 (N_10462,N_9335,N_8778);
or U10463 (N_10463,N_8953,N_8611);
nand U10464 (N_10464,N_9036,N_8615);
nand U10465 (N_10465,N_9890,N_9223);
nor U10466 (N_10466,N_8593,N_9302);
nand U10467 (N_10467,N_8049,N_8913);
nor U10468 (N_10468,N_9644,N_8613);
and U10469 (N_10469,N_8284,N_9443);
or U10470 (N_10470,N_8483,N_9035);
and U10471 (N_10471,N_9192,N_8186);
and U10472 (N_10472,N_9081,N_9458);
nor U10473 (N_10473,N_8999,N_8738);
nand U10474 (N_10474,N_9576,N_8637);
nand U10475 (N_10475,N_9007,N_9924);
xnor U10476 (N_10476,N_8993,N_9429);
or U10477 (N_10477,N_8071,N_8301);
xnor U10478 (N_10478,N_9008,N_8664);
xnor U10479 (N_10479,N_8588,N_8654);
nand U10480 (N_10480,N_9285,N_8218);
xnor U10481 (N_10481,N_8138,N_9988);
and U10482 (N_10482,N_8557,N_9564);
nand U10483 (N_10483,N_9730,N_8581);
or U10484 (N_10484,N_9260,N_9315);
and U10485 (N_10485,N_8061,N_8053);
nand U10486 (N_10486,N_9871,N_9631);
and U10487 (N_10487,N_9508,N_9703);
nor U10488 (N_10488,N_8794,N_9541);
or U10489 (N_10489,N_8216,N_8427);
xnor U10490 (N_10490,N_8977,N_9185);
or U10491 (N_10491,N_9202,N_8529);
and U10492 (N_10492,N_9200,N_9805);
or U10493 (N_10493,N_8487,N_9984);
nand U10494 (N_10494,N_8869,N_8987);
xnor U10495 (N_10495,N_9196,N_8679);
nand U10496 (N_10496,N_9911,N_9943);
xor U10497 (N_10497,N_8724,N_8513);
nor U10498 (N_10498,N_9354,N_8673);
or U10499 (N_10499,N_9642,N_9544);
and U10500 (N_10500,N_9857,N_8733);
and U10501 (N_10501,N_9462,N_9849);
or U10502 (N_10502,N_9533,N_9951);
nor U10503 (N_10503,N_9270,N_9169);
or U10504 (N_10504,N_9383,N_9586);
nand U10505 (N_10505,N_9711,N_9850);
or U10506 (N_10506,N_9140,N_8093);
and U10507 (N_10507,N_9338,N_8655);
or U10508 (N_10508,N_8300,N_8789);
nand U10509 (N_10509,N_8506,N_8621);
or U10510 (N_10510,N_9412,N_8676);
nand U10511 (N_10511,N_8431,N_8791);
nor U10512 (N_10512,N_8921,N_8620);
nand U10513 (N_10513,N_8745,N_9577);
and U10514 (N_10514,N_9444,N_8622);
and U10515 (N_10515,N_8316,N_8134);
and U10516 (N_10516,N_9632,N_8266);
xor U10517 (N_10517,N_9466,N_9998);
nor U10518 (N_10518,N_9583,N_8540);
or U10519 (N_10519,N_8975,N_8873);
and U10520 (N_10520,N_8754,N_9797);
xor U10521 (N_10521,N_8289,N_8429);
xor U10522 (N_10522,N_8696,N_9821);
nand U10523 (N_10523,N_8750,N_9334);
nand U10524 (N_10524,N_8388,N_9992);
nand U10525 (N_10525,N_8508,N_8269);
or U10526 (N_10526,N_8165,N_8140);
nor U10527 (N_10527,N_9842,N_9225);
and U10528 (N_10528,N_9172,N_9244);
nand U10529 (N_10529,N_9552,N_9117);
nor U10530 (N_10530,N_8179,N_8243);
xnor U10531 (N_10531,N_8567,N_8096);
and U10532 (N_10532,N_8511,N_8381);
or U10533 (N_10533,N_8325,N_9257);
nand U10534 (N_10534,N_9971,N_9683);
nand U10535 (N_10535,N_9416,N_9858);
nand U10536 (N_10536,N_9473,N_9477);
or U10537 (N_10537,N_8646,N_8939);
or U10538 (N_10538,N_9908,N_9406);
xor U10539 (N_10539,N_8149,N_9671);
and U10540 (N_10540,N_9699,N_9000);
nor U10541 (N_10541,N_8856,N_9921);
nand U10542 (N_10542,N_8917,N_8587);
nand U10543 (N_10543,N_9025,N_9687);
nand U10544 (N_10544,N_9841,N_8833);
and U10545 (N_10545,N_8219,N_9324);
and U10546 (N_10546,N_9529,N_9242);
nor U10547 (N_10547,N_8171,N_9422);
or U10548 (N_10548,N_9163,N_9602);
nand U10549 (N_10549,N_8779,N_9681);
or U10550 (N_10550,N_9148,N_9920);
xor U10551 (N_10551,N_9249,N_9779);
or U10552 (N_10552,N_8262,N_8156);
nand U10553 (N_10553,N_8226,N_8324);
nand U10554 (N_10554,N_9814,N_8979);
and U10555 (N_10555,N_9235,N_8160);
nor U10556 (N_10556,N_9877,N_9531);
nor U10557 (N_10557,N_8691,N_9952);
nand U10558 (N_10558,N_8729,N_8714);
and U10559 (N_10559,N_8955,N_9557);
nand U10560 (N_10560,N_9151,N_9471);
or U10561 (N_10561,N_9660,N_8553);
and U10562 (N_10562,N_9333,N_9424);
and U10563 (N_10563,N_8922,N_9055);
or U10564 (N_10564,N_8859,N_8829);
and U10565 (N_10565,N_8994,N_9374);
nor U10566 (N_10566,N_9489,N_8079);
and U10567 (N_10567,N_9161,N_9198);
or U10568 (N_10568,N_9934,N_9203);
or U10569 (N_10569,N_8845,N_9300);
and U10570 (N_10570,N_9504,N_9136);
nor U10571 (N_10571,N_9067,N_9873);
nand U10572 (N_10572,N_8772,N_8369);
and U10573 (N_10573,N_9968,N_8370);
xor U10574 (N_10574,N_8350,N_8076);
xor U10575 (N_10575,N_8705,N_9655);
nand U10576 (N_10576,N_8457,N_8844);
and U10577 (N_10577,N_9248,N_9912);
nor U10578 (N_10578,N_9872,N_8197);
nor U10579 (N_10579,N_8349,N_9348);
xor U10580 (N_10580,N_8698,N_9230);
or U10581 (N_10581,N_8161,N_8038);
xnor U10582 (N_10582,N_9207,N_9656);
and U10583 (N_10583,N_9317,N_9958);
or U10584 (N_10584,N_9421,N_8371);
or U10585 (N_10585,N_9046,N_9507);
or U10586 (N_10586,N_8986,N_9630);
nand U10587 (N_10587,N_8766,N_9159);
or U10588 (N_10588,N_9213,N_9664);
or U10589 (N_10589,N_8063,N_8585);
nor U10590 (N_10590,N_9962,N_8072);
xor U10591 (N_10591,N_9134,N_8638);
nor U10592 (N_10592,N_9582,N_8124);
or U10593 (N_10593,N_9558,N_9241);
and U10594 (N_10594,N_8562,N_8559);
and U10595 (N_10595,N_8329,N_9524);
or U10596 (N_10596,N_9452,N_8658);
xnor U10597 (N_10597,N_9265,N_8182);
xnor U10598 (N_10598,N_8475,N_8935);
or U10599 (N_10599,N_9629,N_9876);
xor U10600 (N_10600,N_8413,N_9379);
xnor U10601 (N_10601,N_8653,N_9123);
nor U10602 (N_10602,N_9372,N_9766);
nor U10603 (N_10603,N_9698,N_9989);
and U10604 (N_10604,N_8645,N_8279);
nand U10605 (N_10605,N_8759,N_9188);
xor U10606 (N_10606,N_9043,N_9124);
nor U10607 (N_10607,N_8552,N_8864);
or U10608 (N_10608,N_8905,N_8574);
nand U10609 (N_10609,N_9726,N_8141);
nor U10610 (N_10610,N_9868,N_9074);
nand U10611 (N_10611,N_9549,N_9446);
xor U10612 (N_10612,N_8865,N_9410);
xnor U10613 (N_10613,N_9844,N_8717);
xnor U10614 (N_10614,N_9502,N_9702);
nand U10615 (N_10615,N_8697,N_9661);
nor U10616 (N_10616,N_8634,N_8084);
or U10617 (N_10617,N_9874,N_9573);
xor U10618 (N_10618,N_8343,N_9026);
nor U10619 (N_10619,N_9436,N_8781);
nor U10620 (N_10620,N_9377,N_9084);
nor U10621 (N_10621,N_8583,N_9066);
or U10622 (N_10622,N_8603,N_9131);
nand U10623 (N_10623,N_8014,N_8784);
nand U10624 (N_10624,N_8155,N_8450);
or U10625 (N_10625,N_8590,N_9535);
nor U10626 (N_10626,N_8866,N_8456);
xor U10627 (N_10627,N_8825,N_8402);
and U10628 (N_10628,N_9240,N_9659);
or U10629 (N_10629,N_8008,N_9967);
xor U10630 (N_10630,N_9205,N_9152);
nand U10631 (N_10631,N_8704,N_9749);
nor U10632 (N_10632,N_9236,N_8086);
nand U10633 (N_10633,N_9120,N_9771);
and U10634 (N_10634,N_9310,N_9767);
xor U10635 (N_10635,N_9170,N_9114);
or U10636 (N_10636,N_9095,N_8795);
nor U10637 (N_10637,N_9359,N_9139);
and U10638 (N_10638,N_8793,N_8948);
or U10639 (N_10639,N_8565,N_8584);
xor U10640 (N_10640,N_9861,N_9722);
and U10641 (N_10641,N_9570,N_9742);
nand U10642 (N_10642,N_9594,N_8797);
or U10643 (N_10643,N_9193,N_8709);
nand U10644 (N_10644,N_8608,N_8229);
and U10645 (N_10645,N_8525,N_9898);
nor U10646 (N_10646,N_9674,N_9211);
nand U10647 (N_10647,N_9776,N_8900);
xor U10648 (N_10648,N_9286,N_9432);
or U10649 (N_10649,N_8444,N_9554);
and U10650 (N_10650,N_9697,N_9737);
xnor U10651 (N_10651,N_9267,N_9247);
nor U10652 (N_10652,N_9094,N_9902);
or U10653 (N_10653,N_8142,N_9331);
nand U10654 (N_10654,N_9304,N_9183);
nor U10655 (N_10655,N_9990,N_9917);
or U10656 (N_10656,N_8834,N_9171);
nand U10657 (N_10657,N_9329,N_8230);
xnor U10658 (N_10658,N_9321,N_8313);
or U10659 (N_10659,N_9498,N_8992);
or U10660 (N_10660,N_8404,N_9581);
nand U10661 (N_10661,N_8060,N_8841);
or U10662 (N_10662,N_8893,N_8177);
and U10663 (N_10663,N_8386,N_8902);
and U10664 (N_10664,N_8362,N_8054);
xnor U10665 (N_10665,N_9695,N_8337);
or U10666 (N_10666,N_9186,N_9453);
xnor U10667 (N_10667,N_8636,N_8057);
xor U10668 (N_10668,N_8185,N_8995);
or U10669 (N_10669,N_8523,N_8650);
xor U10670 (N_10670,N_8126,N_9950);
xor U10671 (N_10671,N_8326,N_9318);
and U10672 (N_10672,N_9810,N_9033);
nand U10673 (N_10673,N_9623,N_9138);
nor U10674 (N_10674,N_8925,N_8734);
nand U10675 (N_10675,N_9717,N_9362);
and U10676 (N_10676,N_9472,N_9828);
xor U10677 (N_10677,N_9936,N_9976);
xor U10678 (N_10678,N_8211,N_9817);
and U10679 (N_10679,N_8633,N_8148);
or U10680 (N_10680,N_9840,N_8091);
and U10681 (N_10681,N_9206,N_8345);
and U10682 (N_10682,N_8221,N_8819);
and U10683 (N_10683,N_9224,N_9113);
xor U10684 (N_10684,N_8299,N_8575);
and U10685 (N_10685,N_8678,N_8416);
xor U10686 (N_10686,N_9519,N_8151);
nand U10687 (N_10687,N_9322,N_8952);
or U10688 (N_10688,N_9663,N_8055);
nor U10689 (N_10689,N_8743,N_8247);
nor U10690 (N_10690,N_9038,N_9612);
xor U10691 (N_10691,N_8623,N_9928);
xor U10692 (N_10692,N_9809,N_9923);
xnor U10693 (N_10693,N_8796,N_9380);
nor U10694 (N_10694,N_9112,N_9040);
nand U10695 (N_10695,N_8667,N_9237);
nand U10696 (N_10696,N_8536,N_8971);
nor U10697 (N_10697,N_9044,N_9725);
and U10698 (N_10698,N_9469,N_9782);
and U10699 (N_10699,N_9959,N_9977);
and U10700 (N_10700,N_9272,N_9806);
or U10701 (N_10701,N_8478,N_9736);
and U10702 (N_10702,N_8168,N_9418);
nand U10703 (N_10703,N_9351,N_9640);
xnor U10704 (N_10704,N_9546,N_9914);
xor U10705 (N_10705,N_8294,N_8802);
nor U10706 (N_10706,N_9812,N_8758);
and U10707 (N_10707,N_9685,N_9050);
or U10708 (N_10708,N_8960,N_8108);
nand U10709 (N_10709,N_9365,N_8482);
nor U10710 (N_10710,N_8391,N_8539);
nor U10711 (N_10711,N_8983,N_8800);
xor U10712 (N_10712,N_8944,N_8852);
nand U10713 (N_10713,N_9662,N_8152);
nor U10714 (N_10714,N_9750,N_9101);
nor U10715 (N_10715,N_9625,N_8788);
nor U10716 (N_10716,N_8006,N_9926);
xnor U10717 (N_10717,N_9413,N_9150);
xnor U10718 (N_10718,N_9621,N_9929);
xor U10719 (N_10719,N_9972,N_9851);
or U10720 (N_10720,N_8265,N_9456);
or U10721 (N_10721,N_8640,N_8050);
nand U10722 (N_10722,N_8046,N_8025);
nand U10723 (N_10723,N_9718,N_9765);
nand U10724 (N_10724,N_9209,N_8931);
nor U10725 (N_10725,N_8520,N_9252);
nand U10726 (N_10726,N_8448,N_9808);
nor U10727 (N_10727,N_8923,N_9897);
nand U10728 (N_10728,N_9187,N_9125);
nor U10729 (N_10729,N_9827,N_8307);
nand U10730 (N_10730,N_9023,N_8614);
nor U10731 (N_10731,N_9018,N_8560);
xor U10732 (N_10732,N_9909,N_8748);
nand U10733 (N_10733,N_9028,N_9775);
nand U10734 (N_10734,N_8470,N_8065);
nand U10735 (N_10735,N_8322,N_9639);
nand U10736 (N_10736,N_9284,N_9110);
or U10737 (N_10737,N_8826,N_8624);
nor U10738 (N_10738,N_9011,N_8174);
nand U10739 (N_10739,N_9543,N_9077);
xnor U10740 (N_10740,N_8170,N_8407);
xor U10741 (N_10741,N_8682,N_9613);
nor U10742 (N_10742,N_9652,N_8632);
or U10743 (N_10743,N_8139,N_8803);
xor U10744 (N_10744,N_8463,N_8718);
nor U10745 (N_10745,N_9017,N_8465);
xnor U10746 (N_10746,N_8651,N_9838);
and U10747 (N_10747,N_9493,N_8997);
and U10748 (N_10748,N_8011,N_9754);
nand U10749 (N_10749,N_9173,N_9889);
or U10750 (N_10750,N_9180,N_8372);
xor U10751 (N_10751,N_8838,N_9122);
or U10752 (N_10752,N_8735,N_9405);
and U10753 (N_10753,N_8066,N_8964);
nor U10754 (N_10754,N_8485,N_9527);
nand U10755 (N_10755,N_9815,N_8700);
nand U10756 (N_10756,N_9734,N_8998);
and U10757 (N_10757,N_8291,N_9474);
or U10758 (N_10758,N_8272,N_9795);
xor U10759 (N_10759,N_9668,N_9417);
and U10760 (N_10760,N_8566,N_8331);
nor U10761 (N_10761,N_8254,N_8162);
xor U10762 (N_10762,N_8891,N_9370);
xnor U10763 (N_10763,N_8686,N_9153);
nand U10764 (N_10764,N_8437,N_9618);
nand U10765 (N_10765,N_9459,N_9983);
nand U10766 (N_10766,N_8178,N_9479);
nand U10767 (N_10767,N_8377,N_9807);
and U10768 (N_10768,N_8173,N_9666);
nor U10769 (N_10769,N_8031,N_9551);
and U10770 (N_10770,N_9275,N_9927);
nor U10771 (N_10771,N_8771,N_9863);
or U10772 (N_10772,N_9259,N_9753);
xnor U10773 (N_10773,N_9054,N_9622);
and U10774 (N_10774,N_8592,N_8692);
nand U10775 (N_10775,N_8409,N_9949);
nand U10776 (N_10776,N_8721,N_8298);
nor U10777 (N_10777,N_9875,N_9389);
or U10778 (N_10778,N_8244,N_9449);
nor U10779 (N_10779,N_8538,N_8821);
or U10780 (N_10780,N_9792,N_9643);
or U10781 (N_10781,N_9550,N_9097);
and U10782 (N_10782,N_9818,N_8418);
xor U10783 (N_10783,N_8984,N_9448);
xor U10784 (N_10784,N_9780,N_8163);
or U10785 (N_10785,N_8909,N_9461);
nor U10786 (N_10786,N_8911,N_9283);
nor U10787 (N_10787,N_8522,N_9042);
xor U10788 (N_10788,N_8309,N_8600);
nor U10789 (N_10789,N_9109,N_9611);
or U10790 (N_10790,N_9041,N_8133);
or U10791 (N_10791,N_8991,N_8753);
xor U10792 (N_10792,N_9494,N_9970);
and U10793 (N_10793,N_8966,N_9946);
or U10794 (N_10794,N_8198,N_9232);
nor U10795 (N_10795,N_8406,N_8730);
and U10796 (N_10796,N_8665,N_9724);
nand U10797 (N_10797,N_9395,N_8217);
and U10798 (N_10798,N_9273,N_8723);
nor U10799 (N_10799,N_9536,N_9688);
or U10800 (N_10800,N_8315,N_8153);
nor U10801 (N_10801,N_8432,N_8201);
or U10802 (N_10802,N_8549,N_8545);
nand U10803 (N_10803,N_9903,N_8235);
nand U10804 (N_10804,N_8234,N_8184);
or U10805 (N_10805,N_9619,N_9146);
nand U10806 (N_10806,N_9800,N_9614);
and U10807 (N_10807,N_8420,N_9210);
nand U10808 (N_10808,N_9261,N_9520);
nor U10809 (N_10809,N_9843,N_9654);
or U10810 (N_10810,N_8256,N_8094);
nor U10811 (N_10811,N_9670,N_8985);
and U10812 (N_10812,N_8901,N_8002);
nor U10813 (N_10813,N_8742,N_9264);
nand U10814 (N_10814,N_9307,N_9899);
or U10815 (N_10815,N_8379,N_8740);
nand U10816 (N_10816,N_9738,N_8222);
nor U10817 (N_10817,N_9680,N_9130);
and U10818 (N_10818,N_9451,N_8945);
or U10819 (N_10819,N_8412,N_8353);
or U10820 (N_10820,N_9879,N_8775);
nor U10821 (N_10821,N_9447,N_9837);
and U10822 (N_10822,N_9770,N_9085);
xor U10823 (N_10823,N_8591,N_8694);
nand U10824 (N_10824,N_9052,N_9355);
nand U10825 (N_10825,N_9935,N_9065);
or U10826 (N_10826,N_9254,N_8196);
nor U10827 (N_10827,N_9609,N_9049);
and U10828 (N_10828,N_8214,N_8332);
nand U10829 (N_10829,N_9024,N_8428);
xnor U10830 (N_10830,N_9980,N_9107);
xnor U10831 (N_10831,N_8276,N_8627);
and U10832 (N_10832,N_8854,N_8783);
nor U10833 (N_10833,N_8213,N_8110);
nand U10834 (N_10834,N_9019,N_9787);
nand U10835 (N_10835,N_8268,N_8118);
xor U10836 (N_10836,N_8737,N_8578);
xnor U10837 (N_10837,N_8280,N_8874);
or U10838 (N_10838,N_9330,N_8666);
xnor U10839 (N_10839,N_8010,N_9430);
xnor U10840 (N_10840,N_9415,N_8210);
or U10841 (N_10841,N_9729,N_9053);
nand U10842 (N_10842,N_9528,N_9966);
and U10843 (N_10843,N_8941,N_9029);
xor U10844 (N_10844,N_9965,N_9714);
or U10845 (N_10845,N_8249,N_9743);
or U10846 (N_10846,N_9559,N_9208);
nand U10847 (N_10847,N_9646,N_9367);
nand U10848 (N_10848,N_9288,N_9825);
nand U10849 (N_10849,N_8683,N_8914);
or U10850 (N_10850,N_8288,N_9126);
xnor U10851 (N_10851,N_8020,N_8039);
and U10852 (N_10852,N_8099,N_8024);
nand U10853 (N_10853,N_8499,N_9701);
or U10854 (N_10854,N_9482,N_8458);
nand U10855 (N_10855,N_8318,N_8628);
nor U10856 (N_10856,N_9128,N_8726);
and U10857 (N_10857,N_9411,N_9831);
nand U10858 (N_10858,N_9534,N_8145);
xnor U10859 (N_10859,N_8373,N_8340);
nor U10860 (N_10860,N_9290,N_9500);
and U10861 (N_10861,N_8036,N_9425);
nand U10862 (N_10862,N_8719,N_9759);
xnor U10863 (N_10863,N_9457,N_9974);
xor U10864 (N_10864,N_8356,N_9832);
nor U10865 (N_10865,N_9431,N_8912);
or U10866 (N_10866,N_8573,N_9667);
and U10867 (N_10867,N_8498,N_9636);
nand U10868 (N_10868,N_8166,N_9562);
or U10869 (N_10869,N_8045,N_8471);
or U10870 (N_10870,N_8172,N_8486);
or U10871 (N_10871,N_9414,N_9727);
nor U10872 (N_10872,N_8967,N_8492);
and U10873 (N_10873,N_9690,N_8947);
xnor U10874 (N_10874,N_8068,N_8936);
nor U10875 (N_10875,N_9121,N_8582);
nor U10876 (N_10876,N_8850,N_8380);
nor U10877 (N_10877,N_8711,N_9344);
xor U10878 (N_10878,N_9349,N_8154);
or U10879 (N_10879,N_9526,N_8674);
and U10880 (N_10880,N_8969,N_9647);
nor U10881 (N_10881,N_9834,N_9118);
or U10882 (N_10882,N_8358,N_8959);
xor U10883 (N_10883,N_8532,N_8015);
or U10884 (N_10884,N_8639,N_8253);
xnor U10885 (N_10885,N_9316,N_9227);
and U10886 (N_10886,N_8857,N_8716);
and U10887 (N_10887,N_8689,N_9251);
nand U10888 (N_10888,N_8516,N_8026);
nor U10889 (N_10889,N_9947,N_8323);
nor U10890 (N_10890,N_8801,N_9906);
nand U10891 (N_10891,N_9649,N_9191);
or U10892 (N_10892,N_9509,N_9233);
and U10893 (N_10893,N_8248,N_9939);
nor U10894 (N_10894,N_8242,N_8956);
xor U10895 (N_10895,N_9878,N_9891);
nor U10896 (N_10896,N_9309,N_8477);
xnor U10897 (N_10897,N_9060,N_8928);
nor U10898 (N_10898,N_8571,N_8042);
and U10899 (N_10899,N_9470,N_9082);
or U10900 (N_10900,N_9803,N_8215);
nand U10901 (N_10901,N_8657,N_8327);
xnor U10902 (N_10902,N_9246,N_9369);
and U10903 (N_10903,N_9371,N_8547);
nand U10904 (N_10904,N_9158,N_9852);
nand U10905 (N_10905,N_9816,N_9839);
nand U10906 (N_10906,N_9565,N_9627);
or U10907 (N_10907,N_8806,N_8342);
or U10908 (N_10908,N_9658,N_8100);
nand U10909 (N_10909,N_8481,N_8460);
nand U10910 (N_10910,N_8263,N_8851);
nor U10911 (N_10911,N_8375,N_8546);
xnor U10912 (N_10912,N_8988,N_9589);
xor U10913 (N_10913,N_8785,N_8589);
xor U10914 (N_10914,N_8052,N_8927);
nand U10915 (N_10915,N_9194,N_9181);
nand U10916 (N_10916,N_9963,N_8702);
nand U10917 (N_10917,N_9301,N_9467);
and U10918 (N_10918,N_9514,N_8157);
nand U10919 (N_10919,N_8642,N_9592);
and U10920 (N_10920,N_8203,N_8899);
nand U10921 (N_10921,N_8495,N_9913);
nand U10922 (N_10922,N_9353,N_9948);
nor U10923 (N_10923,N_8285,N_9981);
nor U10924 (N_10924,N_8346,N_9813);
nor U10925 (N_10925,N_9944,N_9957);
xor U10926 (N_10926,N_9700,N_9250);
nand U10927 (N_10927,N_9757,N_9880);
and U10928 (N_10928,N_8454,N_8220);
or U10929 (N_10929,N_9761,N_9918);
nand U10930 (N_10930,N_8680,N_9707);
or U10931 (N_10931,N_9397,N_9129);
nor U10932 (N_10932,N_9219,N_8619);
or U10933 (N_10933,N_9175,N_8690);
xor U10934 (N_10934,N_9786,N_9426);
or U10935 (N_10935,N_9142,N_8805);
nor U10936 (N_10936,N_9855,N_9047);
or U10937 (N_10937,N_9388,N_8426);
nor U10938 (N_10938,N_9820,N_8472);
xnor U10939 (N_10939,N_9435,N_8727);
xnor U10940 (N_10940,N_8968,N_8871);
and U10941 (N_10941,N_9168,N_8776);
or U10942 (N_10942,N_9311,N_8542);
xnor U10943 (N_10943,N_8907,N_9739);
nand U10944 (N_10944,N_8396,N_8405);
nor U10945 (N_10945,N_9373,N_9517);
nand U10946 (N_10946,N_8820,N_8688);
nand U10947 (N_10947,N_9945,N_8357);
nor U10948 (N_10948,N_8452,N_8311);
nor U10949 (N_10949,N_8116,N_9258);
and U10950 (N_10950,N_8383,N_8940);
xnor U10951 (N_10951,N_8092,N_8828);
nand U10952 (N_10952,N_8193,N_8932);
nor U10953 (N_10953,N_9982,N_8708);
and U10954 (N_10954,N_9567,N_8000);
and U10955 (N_10955,N_9995,N_8303);
xnor U10956 (N_10956,N_9245,N_8918);
nand U10957 (N_10957,N_9883,N_8530);
or U10958 (N_10958,N_8419,N_9212);
nand U10959 (N_10959,N_8408,N_8403);
and U10960 (N_10960,N_8376,N_8670);
nor U10961 (N_10961,N_8972,N_8109);
nor U10962 (N_10962,N_8044,N_8411);
xor U10963 (N_10963,N_9538,N_8129);
nand U10964 (N_10964,N_8167,N_9455);
or U10965 (N_10965,N_8739,N_8117);
and U10966 (N_10966,N_9978,N_8048);
nor U10967 (N_10967,N_8631,N_8974);
and U10968 (N_10968,N_8764,N_8526);
xor U10969 (N_10969,N_9653,N_8660);
or U10970 (N_10970,N_9585,N_8202);
nor U10971 (N_10971,N_8609,N_9022);
nand U10972 (N_10972,N_8359,N_9596);
nor U10973 (N_10973,N_8095,N_8877);
and U10974 (N_10974,N_8644,N_8556);
nor U10975 (N_10975,N_9822,N_8929);
xnor U10976 (N_10976,N_8512,N_9402);
or U10977 (N_10977,N_8282,N_9905);
nand U10978 (N_10978,N_9465,N_9220);
nor U10979 (N_10979,N_8016,N_9090);
xor U10980 (N_10980,N_9740,N_9867);
nand U10981 (N_10981,N_8677,N_9501);
nand U10982 (N_10982,N_8400,N_8227);
nand U10983 (N_10983,N_8200,N_8978);
and U10984 (N_10984,N_9830,N_8537);
nand U10985 (N_10985,N_8732,N_8361);
nor U10986 (N_10986,N_9865,N_8236);
or U10987 (N_10987,N_8768,N_8041);
and U10988 (N_10988,N_8970,N_8610);
or U10989 (N_10989,N_8004,N_9894);
nand U10990 (N_10990,N_9255,N_8943);
and U10991 (N_10991,N_9062,N_8434);
nor U10992 (N_10992,N_8064,N_9790);
or U10993 (N_10993,N_8963,N_9079);
xor U10994 (N_10994,N_9763,N_9856);
or U10995 (N_10995,N_8423,N_9460);
nand U10996 (N_10996,N_8835,N_8058);
or U10997 (N_10997,N_9217,N_8749);
and U10998 (N_10998,N_8074,N_9297);
xnor U10999 (N_10999,N_9155,N_9226);
xor U11000 (N_11000,N_8001,N_9269);
nor U11001 (N_11001,N_8580,N_8875);
nand U11002 (N_11002,N_8046,N_8117);
xor U11003 (N_11003,N_9019,N_9568);
and U11004 (N_11004,N_9055,N_9201);
or U11005 (N_11005,N_8192,N_9402);
nand U11006 (N_11006,N_9080,N_8395);
xor U11007 (N_11007,N_8920,N_9995);
or U11008 (N_11008,N_8598,N_9776);
nand U11009 (N_11009,N_9608,N_8759);
or U11010 (N_11010,N_9643,N_9109);
xnor U11011 (N_11011,N_9036,N_8563);
nor U11012 (N_11012,N_9530,N_8590);
nand U11013 (N_11013,N_9829,N_8228);
xnor U11014 (N_11014,N_8427,N_8087);
nor U11015 (N_11015,N_9267,N_8408);
and U11016 (N_11016,N_9625,N_9826);
or U11017 (N_11017,N_9204,N_8731);
nor U11018 (N_11018,N_9308,N_8714);
or U11019 (N_11019,N_8606,N_8313);
nand U11020 (N_11020,N_9640,N_9468);
nand U11021 (N_11021,N_8172,N_8643);
and U11022 (N_11022,N_9671,N_8528);
nor U11023 (N_11023,N_8753,N_9329);
nor U11024 (N_11024,N_8541,N_8876);
xnor U11025 (N_11025,N_9983,N_8564);
nor U11026 (N_11026,N_9897,N_9154);
xor U11027 (N_11027,N_9257,N_9784);
xor U11028 (N_11028,N_9302,N_9994);
nor U11029 (N_11029,N_9225,N_8611);
xnor U11030 (N_11030,N_9670,N_9723);
or U11031 (N_11031,N_8968,N_8567);
xnor U11032 (N_11032,N_9011,N_8704);
and U11033 (N_11033,N_9210,N_9766);
and U11034 (N_11034,N_9014,N_8040);
xnor U11035 (N_11035,N_8913,N_9976);
and U11036 (N_11036,N_9295,N_9767);
xor U11037 (N_11037,N_9465,N_8713);
xor U11038 (N_11038,N_9377,N_9489);
xor U11039 (N_11039,N_8604,N_8817);
and U11040 (N_11040,N_9547,N_9250);
or U11041 (N_11041,N_8580,N_9459);
nor U11042 (N_11042,N_9875,N_9524);
or U11043 (N_11043,N_9231,N_8717);
and U11044 (N_11044,N_8818,N_9623);
nand U11045 (N_11045,N_8572,N_8707);
nor U11046 (N_11046,N_9022,N_8857);
nand U11047 (N_11047,N_9381,N_9156);
or U11048 (N_11048,N_9395,N_8890);
nor U11049 (N_11049,N_9406,N_8621);
nor U11050 (N_11050,N_9251,N_8799);
or U11051 (N_11051,N_8420,N_9129);
or U11052 (N_11052,N_8159,N_8857);
nand U11053 (N_11053,N_9070,N_9144);
nand U11054 (N_11054,N_9749,N_9456);
nand U11055 (N_11055,N_9038,N_9857);
or U11056 (N_11056,N_9610,N_9985);
and U11057 (N_11057,N_8212,N_9928);
and U11058 (N_11058,N_9035,N_8390);
or U11059 (N_11059,N_9095,N_8603);
nand U11060 (N_11060,N_9161,N_8232);
nor U11061 (N_11061,N_9292,N_9114);
xnor U11062 (N_11062,N_8402,N_9619);
and U11063 (N_11063,N_9689,N_9478);
xnor U11064 (N_11064,N_9643,N_8686);
xor U11065 (N_11065,N_9269,N_9659);
nor U11066 (N_11066,N_8341,N_9705);
nor U11067 (N_11067,N_8842,N_8820);
and U11068 (N_11068,N_8585,N_9428);
and U11069 (N_11069,N_8115,N_8434);
and U11070 (N_11070,N_8970,N_8743);
and U11071 (N_11071,N_8628,N_9067);
nor U11072 (N_11072,N_9300,N_9639);
xor U11073 (N_11073,N_8566,N_8391);
nand U11074 (N_11074,N_9831,N_9531);
xor U11075 (N_11075,N_9697,N_9878);
xnor U11076 (N_11076,N_8047,N_8895);
nand U11077 (N_11077,N_9582,N_8296);
xor U11078 (N_11078,N_8394,N_9363);
nand U11079 (N_11079,N_9003,N_9139);
nand U11080 (N_11080,N_8159,N_8008);
xnor U11081 (N_11081,N_9853,N_9645);
xnor U11082 (N_11082,N_9286,N_8825);
and U11083 (N_11083,N_8936,N_9605);
xnor U11084 (N_11084,N_8642,N_9841);
xnor U11085 (N_11085,N_9521,N_9867);
and U11086 (N_11086,N_9035,N_8645);
or U11087 (N_11087,N_8989,N_9624);
nor U11088 (N_11088,N_8938,N_9892);
and U11089 (N_11089,N_8568,N_8979);
and U11090 (N_11090,N_9895,N_8393);
and U11091 (N_11091,N_9514,N_8376);
xor U11092 (N_11092,N_8060,N_8979);
or U11093 (N_11093,N_9561,N_8205);
nor U11094 (N_11094,N_8485,N_9900);
or U11095 (N_11095,N_8989,N_8233);
xnor U11096 (N_11096,N_9927,N_8666);
nand U11097 (N_11097,N_8935,N_8172);
nor U11098 (N_11098,N_8617,N_8493);
nor U11099 (N_11099,N_9768,N_8762);
xnor U11100 (N_11100,N_8916,N_8850);
nor U11101 (N_11101,N_9415,N_8120);
nor U11102 (N_11102,N_8300,N_9204);
and U11103 (N_11103,N_9211,N_9920);
or U11104 (N_11104,N_8343,N_9335);
nor U11105 (N_11105,N_8535,N_9631);
xor U11106 (N_11106,N_9890,N_9821);
xnor U11107 (N_11107,N_9786,N_9067);
and U11108 (N_11108,N_8565,N_9740);
and U11109 (N_11109,N_9234,N_8648);
or U11110 (N_11110,N_8184,N_8946);
nor U11111 (N_11111,N_8372,N_9408);
and U11112 (N_11112,N_8897,N_9199);
xor U11113 (N_11113,N_8101,N_9842);
nor U11114 (N_11114,N_9828,N_8579);
xnor U11115 (N_11115,N_8200,N_8638);
or U11116 (N_11116,N_8703,N_9628);
and U11117 (N_11117,N_9507,N_9883);
or U11118 (N_11118,N_8062,N_9656);
nand U11119 (N_11119,N_9574,N_8636);
nand U11120 (N_11120,N_8328,N_9535);
nand U11121 (N_11121,N_9343,N_9676);
or U11122 (N_11122,N_8799,N_9111);
or U11123 (N_11123,N_9072,N_8601);
and U11124 (N_11124,N_9111,N_9696);
and U11125 (N_11125,N_8048,N_9934);
nor U11126 (N_11126,N_8884,N_9937);
nand U11127 (N_11127,N_9004,N_9293);
or U11128 (N_11128,N_8531,N_9320);
and U11129 (N_11129,N_8270,N_9983);
nor U11130 (N_11130,N_8116,N_8283);
xnor U11131 (N_11131,N_9925,N_8980);
xor U11132 (N_11132,N_9837,N_9695);
and U11133 (N_11133,N_9114,N_9077);
nand U11134 (N_11134,N_8040,N_8713);
and U11135 (N_11135,N_8358,N_8566);
xnor U11136 (N_11136,N_8862,N_8515);
and U11137 (N_11137,N_9928,N_9230);
and U11138 (N_11138,N_9628,N_9821);
or U11139 (N_11139,N_9344,N_8410);
nand U11140 (N_11140,N_9501,N_8918);
or U11141 (N_11141,N_8626,N_9343);
or U11142 (N_11142,N_8541,N_8717);
or U11143 (N_11143,N_9435,N_9525);
xor U11144 (N_11144,N_8438,N_8983);
nand U11145 (N_11145,N_9817,N_8051);
and U11146 (N_11146,N_8638,N_9547);
nand U11147 (N_11147,N_8294,N_9046);
or U11148 (N_11148,N_8332,N_9146);
xnor U11149 (N_11149,N_9512,N_9204);
nor U11150 (N_11150,N_8014,N_8274);
nor U11151 (N_11151,N_9305,N_9384);
nand U11152 (N_11152,N_8998,N_9554);
xnor U11153 (N_11153,N_9169,N_9327);
nor U11154 (N_11154,N_9565,N_8035);
xnor U11155 (N_11155,N_9892,N_8535);
and U11156 (N_11156,N_8763,N_9662);
xor U11157 (N_11157,N_9990,N_8173);
nor U11158 (N_11158,N_8350,N_8554);
nand U11159 (N_11159,N_9941,N_9841);
xnor U11160 (N_11160,N_9267,N_8201);
and U11161 (N_11161,N_9629,N_8079);
or U11162 (N_11162,N_9805,N_8140);
xor U11163 (N_11163,N_9262,N_8253);
nor U11164 (N_11164,N_8651,N_8048);
or U11165 (N_11165,N_8426,N_8066);
nand U11166 (N_11166,N_9400,N_8158);
and U11167 (N_11167,N_9661,N_8407);
or U11168 (N_11168,N_8268,N_9550);
nor U11169 (N_11169,N_8931,N_9993);
nor U11170 (N_11170,N_9041,N_8740);
or U11171 (N_11171,N_8432,N_8946);
nor U11172 (N_11172,N_8470,N_9645);
xnor U11173 (N_11173,N_9253,N_9719);
nand U11174 (N_11174,N_9291,N_8122);
nor U11175 (N_11175,N_9675,N_8071);
and U11176 (N_11176,N_9453,N_9361);
or U11177 (N_11177,N_9342,N_8419);
xnor U11178 (N_11178,N_9059,N_8460);
xnor U11179 (N_11179,N_9704,N_8926);
xor U11180 (N_11180,N_9598,N_9778);
nor U11181 (N_11181,N_8574,N_8827);
or U11182 (N_11182,N_9426,N_9751);
and U11183 (N_11183,N_8021,N_9157);
xnor U11184 (N_11184,N_8123,N_9251);
and U11185 (N_11185,N_8470,N_8108);
xnor U11186 (N_11186,N_9946,N_8810);
nor U11187 (N_11187,N_9921,N_8882);
xnor U11188 (N_11188,N_9049,N_9438);
nand U11189 (N_11189,N_9304,N_8347);
or U11190 (N_11190,N_9462,N_9487);
xnor U11191 (N_11191,N_8320,N_9877);
or U11192 (N_11192,N_8546,N_8207);
and U11193 (N_11193,N_8245,N_8050);
or U11194 (N_11194,N_8373,N_9991);
nand U11195 (N_11195,N_8652,N_8987);
and U11196 (N_11196,N_9456,N_8675);
and U11197 (N_11197,N_9464,N_8053);
xnor U11198 (N_11198,N_8605,N_9435);
or U11199 (N_11199,N_9985,N_9529);
and U11200 (N_11200,N_8282,N_8846);
nand U11201 (N_11201,N_9690,N_9315);
nand U11202 (N_11202,N_9037,N_8220);
and U11203 (N_11203,N_8583,N_8911);
nor U11204 (N_11204,N_9450,N_9820);
or U11205 (N_11205,N_9534,N_8731);
xor U11206 (N_11206,N_9055,N_8867);
or U11207 (N_11207,N_9560,N_9557);
or U11208 (N_11208,N_8960,N_8770);
xor U11209 (N_11209,N_8681,N_8614);
nor U11210 (N_11210,N_9180,N_8334);
and U11211 (N_11211,N_9886,N_8805);
and U11212 (N_11212,N_9243,N_9582);
xnor U11213 (N_11213,N_9621,N_9167);
nor U11214 (N_11214,N_9502,N_9761);
or U11215 (N_11215,N_8111,N_8456);
and U11216 (N_11216,N_8274,N_8787);
nor U11217 (N_11217,N_9081,N_8767);
nand U11218 (N_11218,N_8836,N_8774);
nand U11219 (N_11219,N_9984,N_9106);
or U11220 (N_11220,N_8344,N_9612);
or U11221 (N_11221,N_8501,N_8251);
and U11222 (N_11222,N_8207,N_9447);
or U11223 (N_11223,N_8726,N_9620);
and U11224 (N_11224,N_8220,N_9425);
and U11225 (N_11225,N_8516,N_8933);
nand U11226 (N_11226,N_8899,N_9311);
or U11227 (N_11227,N_8654,N_8310);
nor U11228 (N_11228,N_9368,N_9711);
and U11229 (N_11229,N_8782,N_9547);
or U11230 (N_11230,N_9181,N_9495);
nor U11231 (N_11231,N_9793,N_9339);
nor U11232 (N_11232,N_8355,N_8776);
xnor U11233 (N_11233,N_8064,N_9034);
and U11234 (N_11234,N_8439,N_8451);
nand U11235 (N_11235,N_9875,N_9269);
nand U11236 (N_11236,N_8428,N_9161);
nand U11237 (N_11237,N_9040,N_8356);
and U11238 (N_11238,N_8943,N_9195);
and U11239 (N_11239,N_8759,N_9905);
or U11240 (N_11240,N_8899,N_8690);
nand U11241 (N_11241,N_9086,N_8050);
nor U11242 (N_11242,N_8096,N_9877);
nor U11243 (N_11243,N_8999,N_9579);
and U11244 (N_11244,N_9044,N_8910);
or U11245 (N_11245,N_9209,N_9249);
or U11246 (N_11246,N_8450,N_8644);
and U11247 (N_11247,N_8869,N_9871);
or U11248 (N_11248,N_9583,N_9265);
or U11249 (N_11249,N_9045,N_8162);
nor U11250 (N_11250,N_9729,N_9673);
xnor U11251 (N_11251,N_9635,N_8992);
or U11252 (N_11252,N_8413,N_8722);
and U11253 (N_11253,N_9076,N_8385);
nor U11254 (N_11254,N_8389,N_9962);
nor U11255 (N_11255,N_9251,N_9874);
nor U11256 (N_11256,N_9829,N_8502);
and U11257 (N_11257,N_8148,N_9291);
xnor U11258 (N_11258,N_9034,N_8263);
or U11259 (N_11259,N_9998,N_9656);
nor U11260 (N_11260,N_8266,N_9493);
xor U11261 (N_11261,N_8764,N_9289);
xor U11262 (N_11262,N_9056,N_9573);
xnor U11263 (N_11263,N_9597,N_9776);
and U11264 (N_11264,N_8451,N_8624);
and U11265 (N_11265,N_9927,N_9568);
and U11266 (N_11266,N_8618,N_9985);
xnor U11267 (N_11267,N_8392,N_8848);
xnor U11268 (N_11268,N_9299,N_8301);
xor U11269 (N_11269,N_8308,N_9930);
nor U11270 (N_11270,N_8294,N_9289);
or U11271 (N_11271,N_8249,N_8933);
nor U11272 (N_11272,N_9547,N_9464);
or U11273 (N_11273,N_9717,N_8182);
nand U11274 (N_11274,N_9123,N_8391);
nand U11275 (N_11275,N_8786,N_8293);
and U11276 (N_11276,N_8732,N_8022);
nand U11277 (N_11277,N_8857,N_9797);
and U11278 (N_11278,N_8091,N_9108);
and U11279 (N_11279,N_9213,N_8181);
nand U11280 (N_11280,N_8709,N_8256);
nand U11281 (N_11281,N_9714,N_9865);
nand U11282 (N_11282,N_9900,N_8624);
nor U11283 (N_11283,N_8179,N_8139);
nand U11284 (N_11284,N_8681,N_9899);
nor U11285 (N_11285,N_9619,N_8554);
or U11286 (N_11286,N_9865,N_9531);
nand U11287 (N_11287,N_8647,N_9080);
or U11288 (N_11288,N_8309,N_8850);
or U11289 (N_11289,N_8319,N_8859);
nor U11290 (N_11290,N_9344,N_9223);
or U11291 (N_11291,N_8711,N_8161);
or U11292 (N_11292,N_8124,N_9395);
nand U11293 (N_11293,N_9020,N_9177);
nand U11294 (N_11294,N_8189,N_9837);
xnor U11295 (N_11295,N_9408,N_9688);
xnor U11296 (N_11296,N_8268,N_8414);
nor U11297 (N_11297,N_8859,N_9272);
xnor U11298 (N_11298,N_8990,N_9813);
or U11299 (N_11299,N_8141,N_8273);
or U11300 (N_11300,N_8567,N_9664);
nand U11301 (N_11301,N_8259,N_8702);
and U11302 (N_11302,N_9575,N_9399);
nor U11303 (N_11303,N_8033,N_9174);
and U11304 (N_11304,N_8543,N_8668);
or U11305 (N_11305,N_8286,N_8691);
nand U11306 (N_11306,N_9600,N_8230);
nand U11307 (N_11307,N_9822,N_9318);
or U11308 (N_11308,N_8426,N_9283);
nor U11309 (N_11309,N_9861,N_9798);
or U11310 (N_11310,N_9587,N_9905);
xor U11311 (N_11311,N_8210,N_8700);
and U11312 (N_11312,N_9455,N_9549);
and U11313 (N_11313,N_8551,N_8633);
nor U11314 (N_11314,N_8775,N_9597);
nor U11315 (N_11315,N_8521,N_8415);
nor U11316 (N_11316,N_9009,N_8486);
nand U11317 (N_11317,N_8389,N_8001);
nand U11318 (N_11318,N_8467,N_9597);
or U11319 (N_11319,N_9229,N_9626);
xnor U11320 (N_11320,N_8115,N_8329);
and U11321 (N_11321,N_9752,N_8302);
nor U11322 (N_11322,N_8713,N_8380);
or U11323 (N_11323,N_9311,N_9126);
or U11324 (N_11324,N_8995,N_9779);
or U11325 (N_11325,N_8156,N_8241);
and U11326 (N_11326,N_8822,N_9770);
nand U11327 (N_11327,N_8951,N_9674);
nor U11328 (N_11328,N_8812,N_8043);
nor U11329 (N_11329,N_9124,N_9338);
nand U11330 (N_11330,N_8492,N_8097);
or U11331 (N_11331,N_9697,N_9722);
nand U11332 (N_11332,N_9123,N_8555);
nor U11333 (N_11333,N_8040,N_9401);
or U11334 (N_11334,N_9618,N_8658);
xnor U11335 (N_11335,N_8109,N_9275);
or U11336 (N_11336,N_8762,N_9479);
nand U11337 (N_11337,N_8066,N_9240);
and U11338 (N_11338,N_8155,N_9469);
and U11339 (N_11339,N_9768,N_9844);
nand U11340 (N_11340,N_8727,N_9523);
nand U11341 (N_11341,N_9774,N_8864);
or U11342 (N_11342,N_9979,N_9939);
nor U11343 (N_11343,N_8041,N_9302);
or U11344 (N_11344,N_8233,N_9976);
or U11345 (N_11345,N_9335,N_9712);
or U11346 (N_11346,N_9046,N_8271);
nand U11347 (N_11347,N_8860,N_8997);
nor U11348 (N_11348,N_9968,N_9815);
and U11349 (N_11349,N_9286,N_8419);
nor U11350 (N_11350,N_8279,N_9975);
nand U11351 (N_11351,N_9917,N_9552);
and U11352 (N_11352,N_9317,N_8835);
or U11353 (N_11353,N_8736,N_8111);
xor U11354 (N_11354,N_8508,N_8530);
xor U11355 (N_11355,N_8427,N_8553);
xnor U11356 (N_11356,N_9985,N_8686);
nand U11357 (N_11357,N_8636,N_9941);
nand U11358 (N_11358,N_8781,N_9788);
xnor U11359 (N_11359,N_8680,N_8967);
nor U11360 (N_11360,N_9486,N_8313);
or U11361 (N_11361,N_8170,N_9476);
xnor U11362 (N_11362,N_8838,N_9971);
nand U11363 (N_11363,N_8491,N_8105);
or U11364 (N_11364,N_8236,N_8088);
and U11365 (N_11365,N_8978,N_9615);
xnor U11366 (N_11366,N_8229,N_9496);
and U11367 (N_11367,N_8376,N_8302);
or U11368 (N_11368,N_9139,N_8058);
xnor U11369 (N_11369,N_9680,N_9067);
xor U11370 (N_11370,N_9362,N_8325);
nand U11371 (N_11371,N_8308,N_8716);
or U11372 (N_11372,N_9830,N_8356);
nor U11373 (N_11373,N_9297,N_8734);
nand U11374 (N_11374,N_8939,N_8547);
or U11375 (N_11375,N_8436,N_9067);
xor U11376 (N_11376,N_9785,N_9395);
nor U11377 (N_11377,N_8034,N_9725);
nor U11378 (N_11378,N_9442,N_9001);
xnor U11379 (N_11379,N_8819,N_8700);
and U11380 (N_11380,N_9857,N_8260);
or U11381 (N_11381,N_8813,N_9493);
nand U11382 (N_11382,N_9070,N_8316);
nand U11383 (N_11383,N_9579,N_8173);
xor U11384 (N_11384,N_8365,N_9683);
and U11385 (N_11385,N_8678,N_9766);
or U11386 (N_11386,N_8540,N_9750);
xor U11387 (N_11387,N_8762,N_9316);
xor U11388 (N_11388,N_9693,N_8152);
xnor U11389 (N_11389,N_9530,N_9824);
nand U11390 (N_11390,N_8900,N_8528);
nor U11391 (N_11391,N_9506,N_8115);
or U11392 (N_11392,N_8579,N_9235);
xnor U11393 (N_11393,N_9397,N_9196);
nor U11394 (N_11394,N_9119,N_8239);
xnor U11395 (N_11395,N_9122,N_9507);
and U11396 (N_11396,N_9099,N_9702);
and U11397 (N_11397,N_8968,N_9149);
nand U11398 (N_11398,N_8167,N_9781);
nand U11399 (N_11399,N_9460,N_9070);
nor U11400 (N_11400,N_9012,N_8209);
and U11401 (N_11401,N_8398,N_8160);
and U11402 (N_11402,N_9187,N_8176);
nand U11403 (N_11403,N_8545,N_8364);
xnor U11404 (N_11404,N_8733,N_9577);
and U11405 (N_11405,N_9547,N_9627);
or U11406 (N_11406,N_8158,N_8131);
or U11407 (N_11407,N_9851,N_9167);
xor U11408 (N_11408,N_9370,N_8517);
nand U11409 (N_11409,N_9445,N_9325);
nor U11410 (N_11410,N_8642,N_8163);
nor U11411 (N_11411,N_9819,N_9863);
nand U11412 (N_11412,N_9035,N_9823);
xnor U11413 (N_11413,N_8341,N_8248);
nor U11414 (N_11414,N_9507,N_8793);
or U11415 (N_11415,N_9999,N_8330);
nand U11416 (N_11416,N_9239,N_8887);
nor U11417 (N_11417,N_8490,N_8324);
xor U11418 (N_11418,N_8371,N_9455);
nor U11419 (N_11419,N_8556,N_8726);
xnor U11420 (N_11420,N_8805,N_8540);
and U11421 (N_11421,N_9575,N_8049);
nand U11422 (N_11422,N_9970,N_8578);
and U11423 (N_11423,N_8813,N_8318);
nor U11424 (N_11424,N_8314,N_8710);
xnor U11425 (N_11425,N_8020,N_8250);
xnor U11426 (N_11426,N_8509,N_9201);
nand U11427 (N_11427,N_9312,N_8289);
nand U11428 (N_11428,N_9006,N_9650);
and U11429 (N_11429,N_9839,N_8215);
and U11430 (N_11430,N_8042,N_8933);
or U11431 (N_11431,N_8787,N_8300);
nand U11432 (N_11432,N_9602,N_9042);
xnor U11433 (N_11433,N_8373,N_9287);
or U11434 (N_11434,N_8981,N_9498);
xnor U11435 (N_11435,N_8960,N_8454);
nand U11436 (N_11436,N_8479,N_9864);
and U11437 (N_11437,N_9074,N_8516);
and U11438 (N_11438,N_9491,N_9981);
and U11439 (N_11439,N_8172,N_9098);
xor U11440 (N_11440,N_9449,N_9266);
and U11441 (N_11441,N_8825,N_9788);
or U11442 (N_11442,N_8088,N_9062);
and U11443 (N_11443,N_8864,N_8059);
and U11444 (N_11444,N_8009,N_9683);
or U11445 (N_11445,N_8559,N_9630);
xnor U11446 (N_11446,N_8906,N_8466);
or U11447 (N_11447,N_9646,N_8929);
nor U11448 (N_11448,N_9348,N_8893);
nor U11449 (N_11449,N_9893,N_9842);
or U11450 (N_11450,N_8579,N_8713);
and U11451 (N_11451,N_9024,N_8983);
and U11452 (N_11452,N_9569,N_9216);
and U11453 (N_11453,N_9479,N_9481);
or U11454 (N_11454,N_8443,N_8990);
xnor U11455 (N_11455,N_8159,N_9753);
xnor U11456 (N_11456,N_8828,N_8756);
nand U11457 (N_11457,N_8851,N_9789);
and U11458 (N_11458,N_9515,N_8250);
nand U11459 (N_11459,N_9217,N_9623);
or U11460 (N_11460,N_8494,N_9054);
xnor U11461 (N_11461,N_9198,N_8182);
xor U11462 (N_11462,N_9802,N_9191);
xor U11463 (N_11463,N_8722,N_8595);
nor U11464 (N_11464,N_8392,N_8584);
and U11465 (N_11465,N_9417,N_9731);
nor U11466 (N_11466,N_8480,N_9500);
nor U11467 (N_11467,N_8149,N_8612);
or U11468 (N_11468,N_8728,N_8948);
and U11469 (N_11469,N_8574,N_9590);
xor U11470 (N_11470,N_9273,N_9184);
and U11471 (N_11471,N_9617,N_8028);
xnor U11472 (N_11472,N_9774,N_9079);
and U11473 (N_11473,N_8149,N_9148);
and U11474 (N_11474,N_8462,N_9920);
nand U11475 (N_11475,N_8651,N_8471);
xor U11476 (N_11476,N_8031,N_9211);
or U11477 (N_11477,N_8638,N_9102);
nor U11478 (N_11478,N_8262,N_9384);
nand U11479 (N_11479,N_8260,N_9747);
or U11480 (N_11480,N_8614,N_8717);
nand U11481 (N_11481,N_9053,N_8866);
xnor U11482 (N_11482,N_9683,N_8737);
and U11483 (N_11483,N_8537,N_8696);
and U11484 (N_11484,N_9015,N_8852);
nor U11485 (N_11485,N_8391,N_9036);
or U11486 (N_11486,N_9301,N_9051);
nor U11487 (N_11487,N_9611,N_8031);
nand U11488 (N_11488,N_8141,N_8048);
xor U11489 (N_11489,N_8292,N_8818);
xnor U11490 (N_11490,N_8109,N_8132);
or U11491 (N_11491,N_8136,N_8638);
or U11492 (N_11492,N_8207,N_9488);
and U11493 (N_11493,N_8036,N_8139);
nor U11494 (N_11494,N_9771,N_9045);
nor U11495 (N_11495,N_8526,N_8814);
nand U11496 (N_11496,N_8630,N_8875);
nor U11497 (N_11497,N_8369,N_8117);
and U11498 (N_11498,N_9292,N_8072);
and U11499 (N_11499,N_8267,N_8506);
nand U11500 (N_11500,N_9002,N_8425);
and U11501 (N_11501,N_8399,N_9674);
nor U11502 (N_11502,N_9480,N_8094);
and U11503 (N_11503,N_9104,N_8586);
nor U11504 (N_11504,N_8236,N_8902);
or U11505 (N_11505,N_8359,N_8271);
xor U11506 (N_11506,N_9163,N_8630);
nand U11507 (N_11507,N_9022,N_8788);
and U11508 (N_11508,N_8723,N_8127);
xnor U11509 (N_11509,N_9378,N_8924);
nor U11510 (N_11510,N_9591,N_9336);
xnor U11511 (N_11511,N_9972,N_8982);
xnor U11512 (N_11512,N_8890,N_9920);
nor U11513 (N_11513,N_8540,N_8738);
nor U11514 (N_11514,N_8674,N_8554);
or U11515 (N_11515,N_8142,N_9612);
xor U11516 (N_11516,N_8194,N_9594);
nand U11517 (N_11517,N_8496,N_9054);
and U11518 (N_11518,N_8868,N_9586);
or U11519 (N_11519,N_9440,N_8904);
or U11520 (N_11520,N_9580,N_8266);
xor U11521 (N_11521,N_9413,N_8203);
xor U11522 (N_11522,N_8452,N_8433);
and U11523 (N_11523,N_9027,N_8551);
or U11524 (N_11524,N_8815,N_9889);
or U11525 (N_11525,N_9684,N_9524);
and U11526 (N_11526,N_8267,N_9414);
nand U11527 (N_11527,N_9010,N_9739);
and U11528 (N_11528,N_9249,N_8927);
and U11529 (N_11529,N_9776,N_8488);
xnor U11530 (N_11530,N_9959,N_9370);
or U11531 (N_11531,N_9723,N_9041);
or U11532 (N_11532,N_9004,N_9686);
nor U11533 (N_11533,N_9285,N_8932);
or U11534 (N_11534,N_8036,N_9984);
nand U11535 (N_11535,N_8439,N_8987);
xnor U11536 (N_11536,N_8204,N_9515);
or U11537 (N_11537,N_9351,N_9850);
nand U11538 (N_11538,N_8522,N_8035);
or U11539 (N_11539,N_8004,N_9669);
and U11540 (N_11540,N_8471,N_9169);
nand U11541 (N_11541,N_8308,N_9645);
xor U11542 (N_11542,N_8368,N_9465);
nor U11543 (N_11543,N_9446,N_9056);
nand U11544 (N_11544,N_9895,N_9719);
nand U11545 (N_11545,N_9465,N_9795);
nand U11546 (N_11546,N_8014,N_9143);
nand U11547 (N_11547,N_9476,N_8363);
or U11548 (N_11548,N_8428,N_9246);
xnor U11549 (N_11549,N_9394,N_9405);
nand U11550 (N_11550,N_9967,N_8938);
xor U11551 (N_11551,N_9375,N_8977);
xnor U11552 (N_11552,N_8947,N_9646);
xor U11553 (N_11553,N_9814,N_8195);
or U11554 (N_11554,N_9195,N_8331);
xnor U11555 (N_11555,N_8658,N_9555);
nor U11556 (N_11556,N_8808,N_8492);
or U11557 (N_11557,N_8491,N_9544);
and U11558 (N_11558,N_8178,N_8645);
nand U11559 (N_11559,N_9988,N_8020);
nor U11560 (N_11560,N_8341,N_9805);
and U11561 (N_11561,N_8852,N_8748);
nor U11562 (N_11562,N_9053,N_9065);
or U11563 (N_11563,N_9363,N_9638);
xnor U11564 (N_11564,N_9050,N_9981);
and U11565 (N_11565,N_8732,N_8235);
or U11566 (N_11566,N_8749,N_9498);
and U11567 (N_11567,N_9980,N_8914);
nand U11568 (N_11568,N_9524,N_9013);
nand U11569 (N_11569,N_9994,N_8856);
or U11570 (N_11570,N_8205,N_8044);
nand U11571 (N_11571,N_9206,N_9448);
or U11572 (N_11572,N_8103,N_9905);
nor U11573 (N_11573,N_9859,N_9213);
xor U11574 (N_11574,N_9318,N_9883);
and U11575 (N_11575,N_8006,N_9644);
nand U11576 (N_11576,N_8518,N_9064);
or U11577 (N_11577,N_8351,N_8270);
or U11578 (N_11578,N_9292,N_8392);
nand U11579 (N_11579,N_9203,N_9441);
xor U11580 (N_11580,N_8991,N_9532);
and U11581 (N_11581,N_9845,N_9507);
and U11582 (N_11582,N_9912,N_9324);
xnor U11583 (N_11583,N_8635,N_8933);
or U11584 (N_11584,N_9816,N_8100);
nor U11585 (N_11585,N_9700,N_8543);
xor U11586 (N_11586,N_9375,N_9739);
and U11587 (N_11587,N_8292,N_9118);
and U11588 (N_11588,N_8808,N_8839);
nand U11589 (N_11589,N_8891,N_9056);
nor U11590 (N_11590,N_9521,N_9681);
nor U11591 (N_11591,N_9142,N_9436);
and U11592 (N_11592,N_8417,N_9158);
or U11593 (N_11593,N_9178,N_8212);
xor U11594 (N_11594,N_9710,N_8203);
xor U11595 (N_11595,N_8277,N_8789);
nand U11596 (N_11596,N_9476,N_9217);
nor U11597 (N_11597,N_9890,N_9697);
and U11598 (N_11598,N_8166,N_8233);
or U11599 (N_11599,N_9351,N_8495);
nand U11600 (N_11600,N_8462,N_8688);
nand U11601 (N_11601,N_9474,N_8316);
or U11602 (N_11602,N_9907,N_9695);
and U11603 (N_11603,N_8913,N_8419);
nand U11604 (N_11604,N_8043,N_8229);
xnor U11605 (N_11605,N_8168,N_9006);
and U11606 (N_11606,N_8646,N_9151);
and U11607 (N_11607,N_9569,N_9748);
xnor U11608 (N_11608,N_8093,N_9778);
xnor U11609 (N_11609,N_9176,N_8051);
or U11610 (N_11610,N_8088,N_9826);
nor U11611 (N_11611,N_9824,N_9334);
and U11612 (N_11612,N_9429,N_8162);
and U11613 (N_11613,N_8412,N_9357);
nor U11614 (N_11614,N_8252,N_9578);
xnor U11615 (N_11615,N_9918,N_9890);
nor U11616 (N_11616,N_9086,N_8202);
nor U11617 (N_11617,N_8508,N_8314);
nor U11618 (N_11618,N_8682,N_8621);
or U11619 (N_11619,N_9138,N_9964);
xor U11620 (N_11620,N_8115,N_9342);
and U11621 (N_11621,N_9298,N_9576);
nor U11622 (N_11622,N_8658,N_9641);
or U11623 (N_11623,N_8879,N_9925);
and U11624 (N_11624,N_9343,N_8398);
nor U11625 (N_11625,N_8845,N_8519);
nand U11626 (N_11626,N_8899,N_9760);
nor U11627 (N_11627,N_8217,N_8066);
xnor U11628 (N_11628,N_9941,N_8600);
or U11629 (N_11629,N_8222,N_9301);
and U11630 (N_11630,N_9855,N_8171);
and U11631 (N_11631,N_9602,N_9120);
xor U11632 (N_11632,N_8448,N_9434);
xor U11633 (N_11633,N_9458,N_9046);
nand U11634 (N_11634,N_8424,N_9658);
xor U11635 (N_11635,N_9708,N_8533);
or U11636 (N_11636,N_9174,N_9542);
nand U11637 (N_11637,N_9244,N_8889);
nand U11638 (N_11638,N_9582,N_8826);
and U11639 (N_11639,N_9018,N_9758);
or U11640 (N_11640,N_9964,N_8389);
or U11641 (N_11641,N_9901,N_9106);
or U11642 (N_11642,N_8473,N_8670);
nand U11643 (N_11643,N_8867,N_8438);
nor U11644 (N_11644,N_9442,N_9116);
nand U11645 (N_11645,N_8891,N_8150);
nand U11646 (N_11646,N_8053,N_8688);
nor U11647 (N_11647,N_9650,N_9941);
nand U11648 (N_11648,N_9217,N_9655);
and U11649 (N_11649,N_9454,N_9815);
nand U11650 (N_11650,N_9098,N_9418);
nor U11651 (N_11651,N_8685,N_8452);
nor U11652 (N_11652,N_8144,N_9282);
nor U11653 (N_11653,N_8853,N_9622);
or U11654 (N_11654,N_8542,N_8350);
and U11655 (N_11655,N_9666,N_8547);
or U11656 (N_11656,N_8162,N_9299);
and U11657 (N_11657,N_8242,N_9934);
and U11658 (N_11658,N_8278,N_8806);
or U11659 (N_11659,N_9298,N_8006);
or U11660 (N_11660,N_9329,N_8712);
or U11661 (N_11661,N_9240,N_9446);
and U11662 (N_11662,N_8653,N_9728);
and U11663 (N_11663,N_8285,N_9659);
and U11664 (N_11664,N_9738,N_9392);
xor U11665 (N_11665,N_8245,N_8372);
xor U11666 (N_11666,N_9783,N_8711);
xor U11667 (N_11667,N_8660,N_8733);
xor U11668 (N_11668,N_9990,N_8640);
xnor U11669 (N_11669,N_8968,N_9505);
nand U11670 (N_11670,N_9025,N_9822);
or U11671 (N_11671,N_8636,N_8703);
or U11672 (N_11672,N_8041,N_9989);
and U11673 (N_11673,N_9513,N_9539);
nor U11674 (N_11674,N_9388,N_9089);
and U11675 (N_11675,N_8530,N_9568);
or U11676 (N_11676,N_9485,N_8123);
nand U11677 (N_11677,N_8430,N_8881);
nand U11678 (N_11678,N_9938,N_8716);
xnor U11679 (N_11679,N_8409,N_8616);
nand U11680 (N_11680,N_8759,N_9498);
nand U11681 (N_11681,N_8410,N_8000);
nand U11682 (N_11682,N_8868,N_9458);
nand U11683 (N_11683,N_8918,N_9984);
xnor U11684 (N_11684,N_8320,N_8039);
or U11685 (N_11685,N_9379,N_8763);
xor U11686 (N_11686,N_8050,N_9449);
nand U11687 (N_11687,N_9689,N_8436);
nor U11688 (N_11688,N_8360,N_8743);
and U11689 (N_11689,N_9992,N_8412);
and U11690 (N_11690,N_9611,N_9321);
nand U11691 (N_11691,N_9825,N_9617);
nor U11692 (N_11692,N_9746,N_9738);
and U11693 (N_11693,N_9015,N_8287);
or U11694 (N_11694,N_9163,N_8583);
xnor U11695 (N_11695,N_8081,N_8911);
and U11696 (N_11696,N_8997,N_9896);
nor U11697 (N_11697,N_8433,N_8775);
or U11698 (N_11698,N_9235,N_8710);
nand U11699 (N_11699,N_9641,N_9358);
and U11700 (N_11700,N_9524,N_9825);
or U11701 (N_11701,N_9555,N_9567);
xor U11702 (N_11702,N_8789,N_9191);
xor U11703 (N_11703,N_9767,N_9936);
xnor U11704 (N_11704,N_8364,N_8916);
and U11705 (N_11705,N_8466,N_9347);
or U11706 (N_11706,N_8790,N_9423);
or U11707 (N_11707,N_9796,N_8531);
or U11708 (N_11708,N_8556,N_8981);
or U11709 (N_11709,N_9762,N_8744);
or U11710 (N_11710,N_9408,N_8986);
nand U11711 (N_11711,N_8057,N_8519);
nor U11712 (N_11712,N_8315,N_8942);
xnor U11713 (N_11713,N_9314,N_9219);
xor U11714 (N_11714,N_9752,N_9239);
or U11715 (N_11715,N_8148,N_9447);
or U11716 (N_11716,N_9593,N_9340);
nor U11717 (N_11717,N_8327,N_8185);
nor U11718 (N_11718,N_9339,N_8667);
xnor U11719 (N_11719,N_9249,N_9837);
nand U11720 (N_11720,N_9862,N_9105);
nor U11721 (N_11721,N_8918,N_8516);
nand U11722 (N_11722,N_9960,N_8024);
or U11723 (N_11723,N_9273,N_9161);
nor U11724 (N_11724,N_9998,N_9579);
nor U11725 (N_11725,N_8163,N_8190);
nor U11726 (N_11726,N_9138,N_9366);
and U11727 (N_11727,N_9536,N_8783);
and U11728 (N_11728,N_8770,N_8363);
or U11729 (N_11729,N_9081,N_9787);
and U11730 (N_11730,N_8808,N_8813);
nor U11731 (N_11731,N_9897,N_8026);
nor U11732 (N_11732,N_8298,N_8514);
xnor U11733 (N_11733,N_8001,N_9686);
and U11734 (N_11734,N_8836,N_9850);
or U11735 (N_11735,N_9628,N_8696);
and U11736 (N_11736,N_8885,N_8056);
nor U11737 (N_11737,N_9126,N_9001);
or U11738 (N_11738,N_8441,N_8069);
xor U11739 (N_11739,N_8260,N_9670);
nand U11740 (N_11740,N_8385,N_9310);
nand U11741 (N_11741,N_8496,N_9749);
nand U11742 (N_11742,N_8963,N_9017);
nand U11743 (N_11743,N_9634,N_9789);
nand U11744 (N_11744,N_8361,N_8226);
nand U11745 (N_11745,N_9004,N_8815);
nor U11746 (N_11746,N_9983,N_9219);
xnor U11747 (N_11747,N_8794,N_9046);
and U11748 (N_11748,N_9368,N_8193);
xor U11749 (N_11749,N_8707,N_9603);
xnor U11750 (N_11750,N_9401,N_8819);
nand U11751 (N_11751,N_8638,N_8123);
or U11752 (N_11752,N_8925,N_9681);
nor U11753 (N_11753,N_8731,N_9831);
nand U11754 (N_11754,N_9995,N_8722);
and U11755 (N_11755,N_9416,N_8751);
and U11756 (N_11756,N_8445,N_9131);
xnor U11757 (N_11757,N_8039,N_9402);
nor U11758 (N_11758,N_8544,N_9771);
and U11759 (N_11759,N_8100,N_8951);
or U11760 (N_11760,N_9841,N_9892);
nand U11761 (N_11761,N_9343,N_8173);
or U11762 (N_11762,N_8198,N_9274);
nand U11763 (N_11763,N_8117,N_8953);
nor U11764 (N_11764,N_9177,N_8036);
or U11765 (N_11765,N_9990,N_8912);
or U11766 (N_11766,N_9695,N_9514);
and U11767 (N_11767,N_8803,N_9882);
and U11768 (N_11768,N_8713,N_9426);
and U11769 (N_11769,N_8582,N_8272);
xnor U11770 (N_11770,N_9196,N_8098);
nor U11771 (N_11771,N_8739,N_9225);
nor U11772 (N_11772,N_9682,N_9085);
or U11773 (N_11773,N_8258,N_8246);
or U11774 (N_11774,N_8630,N_9088);
nand U11775 (N_11775,N_8585,N_8757);
xnor U11776 (N_11776,N_8871,N_8506);
and U11777 (N_11777,N_8124,N_8143);
and U11778 (N_11778,N_8163,N_9170);
nand U11779 (N_11779,N_9162,N_9927);
and U11780 (N_11780,N_9824,N_8383);
nor U11781 (N_11781,N_9375,N_9026);
nor U11782 (N_11782,N_8588,N_8194);
or U11783 (N_11783,N_9549,N_9469);
nand U11784 (N_11784,N_9889,N_8141);
and U11785 (N_11785,N_8382,N_8134);
nand U11786 (N_11786,N_9071,N_9360);
and U11787 (N_11787,N_9988,N_8744);
nand U11788 (N_11788,N_9512,N_9339);
and U11789 (N_11789,N_8358,N_9630);
nor U11790 (N_11790,N_9757,N_8746);
nor U11791 (N_11791,N_9544,N_8348);
or U11792 (N_11792,N_8617,N_9193);
or U11793 (N_11793,N_9402,N_9094);
or U11794 (N_11794,N_8039,N_9771);
or U11795 (N_11795,N_9404,N_8595);
xnor U11796 (N_11796,N_8653,N_9360);
nand U11797 (N_11797,N_8683,N_9960);
nand U11798 (N_11798,N_8943,N_8913);
nor U11799 (N_11799,N_8150,N_9601);
and U11800 (N_11800,N_9665,N_9982);
nor U11801 (N_11801,N_9954,N_8066);
or U11802 (N_11802,N_8179,N_9787);
nand U11803 (N_11803,N_9208,N_8098);
nor U11804 (N_11804,N_9974,N_9641);
or U11805 (N_11805,N_9688,N_9967);
nor U11806 (N_11806,N_9008,N_8549);
nand U11807 (N_11807,N_9593,N_9890);
and U11808 (N_11808,N_8084,N_9261);
xor U11809 (N_11809,N_8320,N_8684);
nand U11810 (N_11810,N_8692,N_9563);
xnor U11811 (N_11811,N_9783,N_8043);
and U11812 (N_11812,N_8043,N_8699);
nor U11813 (N_11813,N_9123,N_9030);
nand U11814 (N_11814,N_8281,N_8406);
xnor U11815 (N_11815,N_9918,N_9708);
xnor U11816 (N_11816,N_8296,N_8112);
xor U11817 (N_11817,N_8130,N_8083);
xor U11818 (N_11818,N_9350,N_8286);
xor U11819 (N_11819,N_8802,N_9720);
or U11820 (N_11820,N_8451,N_8544);
nor U11821 (N_11821,N_8727,N_8962);
xnor U11822 (N_11822,N_9207,N_8012);
and U11823 (N_11823,N_9747,N_8802);
and U11824 (N_11824,N_9192,N_8053);
nor U11825 (N_11825,N_9807,N_9055);
nor U11826 (N_11826,N_8928,N_8737);
nand U11827 (N_11827,N_8295,N_9947);
xor U11828 (N_11828,N_9436,N_9734);
or U11829 (N_11829,N_9581,N_9496);
nand U11830 (N_11830,N_9712,N_9893);
and U11831 (N_11831,N_8529,N_8913);
and U11832 (N_11832,N_9837,N_8434);
or U11833 (N_11833,N_9746,N_9799);
or U11834 (N_11834,N_8671,N_9270);
nor U11835 (N_11835,N_8038,N_8448);
and U11836 (N_11836,N_9794,N_8718);
and U11837 (N_11837,N_8438,N_8663);
or U11838 (N_11838,N_8823,N_8700);
xnor U11839 (N_11839,N_8582,N_8471);
xor U11840 (N_11840,N_9045,N_8967);
xnor U11841 (N_11841,N_8526,N_8293);
xor U11842 (N_11842,N_8572,N_8640);
or U11843 (N_11843,N_8331,N_8448);
xor U11844 (N_11844,N_8115,N_9980);
or U11845 (N_11845,N_9321,N_8101);
and U11846 (N_11846,N_9847,N_9861);
nand U11847 (N_11847,N_8398,N_8607);
and U11848 (N_11848,N_9986,N_9607);
nand U11849 (N_11849,N_9946,N_9980);
nand U11850 (N_11850,N_8410,N_8902);
nor U11851 (N_11851,N_9588,N_8071);
nand U11852 (N_11852,N_9730,N_8333);
and U11853 (N_11853,N_8191,N_8435);
nor U11854 (N_11854,N_8528,N_8087);
xor U11855 (N_11855,N_9104,N_8035);
nand U11856 (N_11856,N_8254,N_8761);
nor U11857 (N_11857,N_9218,N_8544);
and U11858 (N_11858,N_9361,N_8735);
or U11859 (N_11859,N_8014,N_9219);
xor U11860 (N_11860,N_9538,N_8629);
and U11861 (N_11861,N_9515,N_8096);
and U11862 (N_11862,N_8069,N_8170);
or U11863 (N_11863,N_8678,N_8648);
xor U11864 (N_11864,N_9148,N_9944);
or U11865 (N_11865,N_8777,N_9751);
nand U11866 (N_11866,N_8847,N_8665);
xor U11867 (N_11867,N_8679,N_8013);
nand U11868 (N_11868,N_8668,N_9728);
and U11869 (N_11869,N_8309,N_9359);
nand U11870 (N_11870,N_8724,N_9804);
and U11871 (N_11871,N_8651,N_8546);
and U11872 (N_11872,N_8987,N_8240);
nor U11873 (N_11873,N_9508,N_8829);
and U11874 (N_11874,N_9013,N_8923);
xnor U11875 (N_11875,N_8784,N_9703);
nand U11876 (N_11876,N_9642,N_8472);
nor U11877 (N_11877,N_8714,N_9731);
or U11878 (N_11878,N_8391,N_9565);
xnor U11879 (N_11879,N_8351,N_8300);
or U11880 (N_11880,N_9522,N_9971);
and U11881 (N_11881,N_9286,N_8924);
or U11882 (N_11882,N_9778,N_9684);
or U11883 (N_11883,N_9841,N_8576);
xnor U11884 (N_11884,N_8181,N_8339);
xor U11885 (N_11885,N_8115,N_8603);
nor U11886 (N_11886,N_8267,N_8900);
and U11887 (N_11887,N_9645,N_8300);
nand U11888 (N_11888,N_9722,N_9603);
nand U11889 (N_11889,N_9576,N_9119);
and U11890 (N_11890,N_9659,N_9543);
nor U11891 (N_11891,N_9233,N_9166);
and U11892 (N_11892,N_8599,N_9607);
or U11893 (N_11893,N_8496,N_9811);
nor U11894 (N_11894,N_9658,N_9201);
nand U11895 (N_11895,N_8330,N_8770);
or U11896 (N_11896,N_9439,N_8741);
nor U11897 (N_11897,N_9253,N_9027);
xnor U11898 (N_11898,N_9010,N_9602);
nor U11899 (N_11899,N_8501,N_9358);
nand U11900 (N_11900,N_9895,N_8198);
or U11901 (N_11901,N_8908,N_8749);
or U11902 (N_11902,N_8765,N_8393);
nand U11903 (N_11903,N_9616,N_9130);
or U11904 (N_11904,N_8462,N_9437);
nand U11905 (N_11905,N_8103,N_9803);
and U11906 (N_11906,N_9600,N_8640);
nor U11907 (N_11907,N_8635,N_8349);
and U11908 (N_11908,N_8106,N_8491);
nor U11909 (N_11909,N_8837,N_8956);
or U11910 (N_11910,N_8796,N_8790);
xor U11911 (N_11911,N_9429,N_9209);
nor U11912 (N_11912,N_9373,N_8158);
xnor U11913 (N_11913,N_9790,N_9513);
xnor U11914 (N_11914,N_8553,N_8927);
nand U11915 (N_11915,N_8836,N_9834);
nand U11916 (N_11916,N_9745,N_8548);
and U11917 (N_11917,N_8404,N_8018);
nor U11918 (N_11918,N_9887,N_9997);
nand U11919 (N_11919,N_8136,N_8900);
nor U11920 (N_11920,N_8657,N_9367);
xnor U11921 (N_11921,N_8428,N_8296);
or U11922 (N_11922,N_9832,N_8188);
nand U11923 (N_11923,N_9693,N_9333);
xor U11924 (N_11924,N_8184,N_9212);
and U11925 (N_11925,N_9663,N_8589);
nand U11926 (N_11926,N_8578,N_9723);
and U11927 (N_11927,N_9225,N_8408);
nor U11928 (N_11928,N_9710,N_8541);
nor U11929 (N_11929,N_9360,N_8626);
xnor U11930 (N_11930,N_8162,N_9761);
or U11931 (N_11931,N_8399,N_8212);
or U11932 (N_11932,N_9881,N_8981);
or U11933 (N_11933,N_8293,N_8780);
and U11934 (N_11934,N_8175,N_8909);
and U11935 (N_11935,N_9616,N_8710);
nor U11936 (N_11936,N_9732,N_8430);
xnor U11937 (N_11937,N_8201,N_9415);
or U11938 (N_11938,N_9167,N_8149);
or U11939 (N_11939,N_8332,N_8936);
nand U11940 (N_11940,N_8663,N_9665);
nor U11941 (N_11941,N_9270,N_9804);
nor U11942 (N_11942,N_9918,N_9488);
nand U11943 (N_11943,N_8703,N_9910);
or U11944 (N_11944,N_8741,N_9847);
xnor U11945 (N_11945,N_9338,N_9712);
or U11946 (N_11946,N_8473,N_8262);
and U11947 (N_11947,N_9936,N_9938);
xor U11948 (N_11948,N_8913,N_9127);
and U11949 (N_11949,N_9101,N_8279);
or U11950 (N_11950,N_9883,N_8483);
and U11951 (N_11951,N_9326,N_8645);
nor U11952 (N_11952,N_8925,N_8955);
nor U11953 (N_11953,N_9464,N_8106);
and U11954 (N_11954,N_9093,N_8023);
nand U11955 (N_11955,N_8094,N_9960);
nor U11956 (N_11956,N_9687,N_8107);
or U11957 (N_11957,N_9489,N_8451);
nand U11958 (N_11958,N_9696,N_9898);
or U11959 (N_11959,N_9352,N_8150);
or U11960 (N_11960,N_8298,N_9229);
xnor U11961 (N_11961,N_8332,N_9567);
or U11962 (N_11962,N_8238,N_8349);
nor U11963 (N_11963,N_8065,N_8512);
nor U11964 (N_11964,N_8492,N_9208);
or U11965 (N_11965,N_9287,N_9462);
xnor U11966 (N_11966,N_8881,N_9320);
and U11967 (N_11967,N_9401,N_8342);
xnor U11968 (N_11968,N_8930,N_8773);
and U11969 (N_11969,N_8084,N_8823);
and U11970 (N_11970,N_9775,N_8992);
or U11971 (N_11971,N_9696,N_9821);
and U11972 (N_11972,N_9951,N_9824);
nor U11973 (N_11973,N_8961,N_9674);
xor U11974 (N_11974,N_8890,N_8610);
xor U11975 (N_11975,N_9427,N_9407);
nor U11976 (N_11976,N_9238,N_9825);
or U11977 (N_11977,N_8422,N_9514);
xnor U11978 (N_11978,N_9285,N_9966);
nand U11979 (N_11979,N_9578,N_9641);
xnor U11980 (N_11980,N_9721,N_9219);
and U11981 (N_11981,N_9202,N_9499);
nor U11982 (N_11982,N_8210,N_9103);
nand U11983 (N_11983,N_8293,N_9374);
nor U11984 (N_11984,N_8037,N_8938);
and U11985 (N_11985,N_8466,N_9911);
or U11986 (N_11986,N_8804,N_8641);
nor U11987 (N_11987,N_9144,N_8616);
or U11988 (N_11988,N_9528,N_8422);
and U11989 (N_11989,N_9144,N_8805);
xnor U11990 (N_11990,N_9053,N_9051);
and U11991 (N_11991,N_8032,N_9356);
xnor U11992 (N_11992,N_8656,N_9053);
nor U11993 (N_11993,N_9929,N_8526);
nor U11994 (N_11994,N_8406,N_8748);
xor U11995 (N_11995,N_9546,N_8293);
nand U11996 (N_11996,N_9902,N_9206);
or U11997 (N_11997,N_9542,N_9927);
xnor U11998 (N_11998,N_8117,N_8778);
nand U11999 (N_11999,N_9405,N_9529);
xnor U12000 (N_12000,N_11526,N_10921);
or U12001 (N_12001,N_10623,N_10713);
nor U12002 (N_12002,N_11758,N_10379);
xor U12003 (N_12003,N_10664,N_11942);
and U12004 (N_12004,N_11671,N_10828);
and U12005 (N_12005,N_11280,N_11733);
and U12006 (N_12006,N_11795,N_11098);
xor U12007 (N_12007,N_11558,N_10047);
nor U12008 (N_12008,N_10423,N_11804);
nand U12009 (N_12009,N_10791,N_10621);
nor U12010 (N_12010,N_10200,N_11231);
or U12011 (N_12011,N_10308,N_10861);
xnor U12012 (N_12012,N_10909,N_10689);
and U12013 (N_12013,N_10708,N_11361);
nor U12014 (N_12014,N_11463,N_10278);
xor U12015 (N_12015,N_10454,N_11063);
nand U12016 (N_12016,N_11118,N_10866);
nor U12017 (N_12017,N_10803,N_11834);
and U12018 (N_12018,N_10416,N_10818);
or U12019 (N_12019,N_11051,N_10127);
nand U12020 (N_12020,N_11845,N_10449);
and U12021 (N_12021,N_10907,N_11213);
and U12022 (N_12022,N_10187,N_10966);
nor U12023 (N_12023,N_10654,N_11170);
xnor U12024 (N_12024,N_11099,N_10191);
or U12025 (N_12025,N_11689,N_11979);
and U12026 (N_12026,N_11315,N_10383);
or U12027 (N_12027,N_11174,N_10168);
or U12028 (N_12028,N_10555,N_10351);
or U12029 (N_12029,N_11175,N_11000);
or U12030 (N_12030,N_10928,N_10843);
xnor U12031 (N_12031,N_11256,N_10270);
nor U12032 (N_12032,N_11387,N_11821);
or U12033 (N_12033,N_11591,N_11250);
nor U12034 (N_12034,N_10381,N_10853);
nand U12035 (N_12035,N_10114,N_11489);
nand U12036 (N_12036,N_11934,N_11987);
nor U12037 (N_12037,N_10437,N_11546);
and U12038 (N_12038,N_11582,N_11117);
xor U12039 (N_12039,N_11478,N_11624);
nor U12040 (N_12040,N_11841,N_10789);
nor U12041 (N_12041,N_11792,N_11798);
nand U12042 (N_12042,N_10135,N_11364);
xnor U12043 (N_12043,N_11220,N_10296);
xnor U12044 (N_12044,N_11293,N_11755);
and U12045 (N_12045,N_11778,N_11880);
xor U12046 (N_12046,N_10656,N_10371);
and U12047 (N_12047,N_10960,N_11669);
xnor U12048 (N_12048,N_10865,N_10939);
xnor U12049 (N_12049,N_10076,N_10011);
and U12050 (N_12050,N_10409,N_10983);
nor U12051 (N_12051,N_10574,N_11286);
or U12052 (N_12052,N_10505,N_10233);
or U12053 (N_12053,N_11948,N_11857);
nand U12054 (N_12054,N_11791,N_10164);
nor U12055 (N_12055,N_11865,N_11663);
nand U12056 (N_12056,N_10304,N_10862);
nand U12057 (N_12057,N_10985,N_11074);
xor U12058 (N_12058,N_10489,N_10754);
xnor U12059 (N_12059,N_11352,N_10847);
and U12060 (N_12060,N_11242,N_10156);
nor U12061 (N_12061,N_11868,N_11877);
or U12062 (N_12062,N_11405,N_10659);
xor U12063 (N_12063,N_11818,N_11105);
nand U12064 (N_12064,N_10801,N_10638);
xor U12065 (N_12065,N_10998,N_11221);
and U12066 (N_12066,N_11159,N_11422);
and U12067 (N_12067,N_11125,N_11548);
or U12068 (N_12068,N_11785,N_10008);
nor U12069 (N_12069,N_10685,N_10086);
or U12070 (N_12070,N_10007,N_11045);
xnor U12071 (N_12071,N_10232,N_11907);
nor U12072 (N_12072,N_11727,N_11980);
nand U12073 (N_12073,N_10071,N_11020);
xnor U12074 (N_12074,N_11057,N_11744);
and U12075 (N_12075,N_11413,N_11533);
nand U12076 (N_12076,N_10279,N_10498);
nand U12077 (N_12077,N_11529,N_11557);
or U12078 (N_12078,N_11813,N_11985);
and U12079 (N_12079,N_10082,N_11436);
nor U12080 (N_12080,N_11323,N_11540);
nand U12081 (N_12081,N_10312,N_11205);
nand U12082 (N_12082,N_11937,N_10065);
xor U12083 (N_12083,N_11282,N_10397);
nor U12084 (N_12084,N_10870,N_11404);
or U12085 (N_12085,N_10272,N_11815);
or U12086 (N_12086,N_11986,N_11332);
nand U12087 (N_12087,N_11883,N_11399);
and U12088 (N_12088,N_11717,N_10003);
nor U12089 (N_12089,N_10223,N_10267);
nor U12090 (N_12090,N_11534,N_11563);
xnor U12091 (N_12091,N_11092,N_10752);
xnor U12092 (N_12092,N_11324,N_10937);
and U12093 (N_12093,N_10745,N_10771);
and U12094 (N_12094,N_11803,N_11326);
xor U12095 (N_12095,N_11124,N_11475);
nor U12096 (N_12096,N_10063,N_10766);
xor U12097 (N_12097,N_11071,N_10502);
nand U12098 (N_12098,N_10821,N_10069);
xnor U12099 (N_12099,N_10367,N_10260);
nand U12100 (N_12100,N_11029,N_11470);
xor U12101 (N_12101,N_10629,N_10221);
xnor U12102 (N_12102,N_11501,N_11660);
nand U12103 (N_12103,N_11701,N_11925);
and U12104 (N_12104,N_11973,N_10427);
nor U12105 (N_12105,N_11162,N_11599);
nand U12106 (N_12106,N_10612,N_10341);
and U12107 (N_12107,N_11629,N_11579);
nor U12108 (N_12108,N_11334,N_10228);
nand U12109 (N_12109,N_10350,N_10347);
or U12110 (N_12110,N_11716,N_10276);
and U12111 (N_12111,N_11156,N_11278);
and U12112 (N_12112,N_10701,N_10052);
xor U12113 (N_12113,N_10642,N_11357);
or U12114 (N_12114,N_11208,N_10424);
and U12115 (N_12115,N_10070,N_10706);
xor U12116 (N_12116,N_11692,N_11197);
nor U12117 (N_12117,N_10806,N_11659);
and U12118 (N_12118,N_10478,N_10465);
nand U12119 (N_12119,N_11911,N_10229);
xor U12120 (N_12120,N_10788,N_10984);
nor U12121 (N_12121,N_10744,N_10564);
or U12122 (N_12122,N_10036,N_11210);
nor U12123 (N_12123,N_11995,N_10401);
nand U12124 (N_12124,N_10503,N_10429);
and U12125 (N_12125,N_11955,N_10722);
or U12126 (N_12126,N_10293,N_11161);
and U12127 (N_12127,N_10339,N_10869);
nor U12128 (N_12128,N_11759,N_10412);
nand U12129 (N_12129,N_11371,N_11137);
nand U12130 (N_12130,N_10531,N_10469);
and U12131 (N_12131,N_10194,N_11694);
nand U12132 (N_12132,N_10980,N_11447);
nand U12133 (N_12133,N_10849,N_10370);
nor U12134 (N_12134,N_10743,N_11956);
nor U12135 (N_12135,N_10206,N_11508);
and U12136 (N_12136,N_11183,N_11492);
or U12137 (N_12137,N_10475,N_10760);
nand U12138 (N_12138,N_10002,N_11592);
nor U12139 (N_12139,N_10729,N_11377);
or U12140 (N_12140,N_10222,N_11917);
xnor U12141 (N_12141,N_10961,N_11554);
nand U12142 (N_12142,N_11732,N_11584);
and U12143 (N_12143,N_10438,N_10787);
or U12144 (N_12144,N_10518,N_11662);
nand U12145 (N_12145,N_11199,N_11498);
xor U12146 (N_12146,N_11780,N_10411);
nand U12147 (N_12147,N_10731,N_10521);
or U12148 (N_12148,N_11258,N_11106);
or U12149 (N_12149,N_10702,N_10216);
xor U12150 (N_12150,N_10636,N_10259);
and U12151 (N_12151,N_10652,N_11914);
and U12152 (N_12152,N_11648,N_11551);
xnor U12153 (N_12153,N_11835,N_11353);
xnor U12154 (N_12154,N_11887,N_10833);
nand U12155 (N_12155,N_11076,N_10275);
and U12156 (N_12156,N_10524,N_10378);
nor U12157 (N_12157,N_10212,N_10068);
nor U12158 (N_12158,N_10889,N_11151);
nor U12159 (N_12159,N_11449,N_10770);
and U12160 (N_12160,N_11643,N_11451);
xor U12161 (N_12161,N_10802,N_11038);
nor U12162 (N_12162,N_10895,N_11951);
xor U12163 (N_12163,N_11861,N_10320);
or U12164 (N_12164,N_10558,N_11120);
xor U12165 (N_12165,N_10679,N_11247);
nor U12166 (N_12166,N_10736,N_10274);
and U12167 (N_12167,N_10313,N_11612);
and U12168 (N_12168,N_11539,N_10657);
and U12169 (N_12169,N_10448,N_10101);
or U12170 (N_12170,N_11516,N_11430);
nor U12171 (N_12171,N_11163,N_10342);
nand U12172 (N_12172,N_10039,N_10358);
and U12173 (N_12173,N_10737,N_10408);
or U12174 (N_12174,N_10607,N_11035);
and U12175 (N_12175,N_10352,N_10917);
and U12176 (N_12176,N_11375,N_11686);
and U12177 (N_12177,N_11356,N_10115);
nand U12178 (N_12178,N_11276,N_11906);
nand U12179 (N_12179,N_10203,N_10360);
nand U12180 (N_12180,N_10123,N_11677);
nand U12181 (N_12181,N_10871,N_11201);
nor U12182 (N_12182,N_10768,N_11916);
nand U12183 (N_12183,N_11314,N_10667);
xor U12184 (N_12184,N_10482,N_10125);
nand U12185 (N_12185,N_10635,N_10319);
or U12186 (N_12186,N_11645,N_11506);
nand U12187 (N_12187,N_10170,N_10160);
and U12188 (N_12188,N_11752,N_11424);
and U12189 (N_12189,N_11412,N_11748);
and U12190 (N_12190,N_11972,N_10954);
and U12191 (N_12191,N_10023,N_10285);
and U12192 (N_12192,N_10244,N_10345);
and U12193 (N_12193,N_10709,N_10525);
nand U12194 (N_12194,N_11093,N_11679);
and U12195 (N_12195,N_11851,N_10747);
nand U12196 (N_12196,N_11479,N_10051);
nand U12197 (N_12197,N_11445,N_10691);
nand U12198 (N_12198,N_10060,N_11010);
xor U12199 (N_12199,N_10318,N_11053);
nor U12200 (N_12200,N_11497,N_11634);
xor U12201 (N_12201,N_11613,N_10800);
xnor U12202 (N_12202,N_11774,N_11427);
xnor U12203 (N_12203,N_11022,N_10050);
nand U12204 (N_12204,N_10450,N_11823);
or U12205 (N_12205,N_10458,N_11116);
or U12206 (N_12206,N_11127,N_11376);
nor U12207 (N_12207,N_11503,N_10585);
and U12208 (N_12208,N_10824,N_10120);
or U12209 (N_12209,N_10220,N_11739);
and U12210 (N_12210,N_10337,N_11039);
nand U12211 (N_12211,N_11989,N_10660);
xnor U12212 (N_12212,N_11146,N_11908);
xor U12213 (N_12213,N_11500,N_10653);
nor U12214 (N_12214,N_10924,N_10882);
and U12215 (N_12215,N_11085,N_11933);
nor U12216 (N_12216,N_10377,N_11188);
nor U12217 (N_12217,N_10354,N_11396);
xnor U12218 (N_12218,N_11829,N_10035);
or U12219 (N_12219,N_10850,N_10490);
nand U12220 (N_12220,N_10488,N_11615);
and U12221 (N_12221,N_10305,N_10034);
and U12222 (N_12222,N_10933,N_10395);
or U12223 (N_12223,N_11650,N_10440);
nand U12224 (N_12224,N_11299,N_11670);
and U12225 (N_12225,N_11912,N_11607);
and U12226 (N_12226,N_10561,N_11087);
or U12227 (N_12227,N_11913,N_10193);
or U12228 (N_12228,N_10947,N_11729);
or U12229 (N_12229,N_11448,N_10471);
and U12230 (N_12230,N_11415,N_11464);
nand U12231 (N_12231,N_11982,N_11594);
xnor U12232 (N_12232,N_10362,N_10732);
nor U12233 (N_12233,N_10710,N_10179);
xor U12234 (N_12234,N_10523,N_10648);
nor U12235 (N_12235,N_11443,N_11229);
nand U12236 (N_12236,N_11084,N_11454);
or U12237 (N_12237,N_11617,N_11915);
nor U12238 (N_12238,N_11067,N_11460);
nor U12239 (N_12239,N_11423,N_10663);
nor U12240 (N_12240,N_10603,N_11062);
and U12241 (N_12241,N_10852,N_11721);
nand U12242 (N_12242,N_11627,N_11606);
or U12243 (N_12243,N_10447,N_11378);
or U12244 (N_12244,N_10565,N_10217);
or U12245 (N_12245,N_11013,N_11630);
nand U12246 (N_12246,N_11355,N_10303);
or U12247 (N_12247,N_11570,N_11941);
or U12248 (N_12248,N_10616,N_11988);
nand U12249 (N_12249,N_10528,N_10451);
xor U12250 (N_12250,N_10887,N_10992);
xor U12251 (N_12251,N_11015,N_10751);
and U12252 (N_12252,N_10672,N_11573);
xnor U12253 (N_12253,N_10631,N_10999);
nand U12254 (N_12254,N_11469,N_11674);
nor U12255 (N_12255,N_11603,N_10057);
xor U12256 (N_12256,N_11090,N_10157);
and U12257 (N_12257,N_10746,N_11262);
and U12258 (N_12258,N_11317,N_10322);
or U12259 (N_12259,N_10460,N_11321);
and U12260 (N_12260,N_10972,N_10455);
nor U12261 (N_12261,N_10935,N_11490);
and U12262 (N_12262,N_11653,N_11292);
nand U12263 (N_12263,N_11924,N_10340);
nand U12264 (N_12264,N_10749,N_11585);
nor U12265 (N_12265,N_10507,N_11943);
or U12266 (N_12266,N_10131,N_10236);
or U12267 (N_12267,N_10552,N_10380);
nand U12268 (N_12268,N_10155,N_11958);
and U12269 (N_12269,N_10913,N_10669);
xor U12270 (N_12270,N_11854,N_10598);
nor U12271 (N_12271,N_11388,N_10282);
xnor U12272 (N_12272,N_11224,N_11896);
and U12273 (N_12273,N_10899,N_11919);
xor U12274 (N_12274,N_11947,N_10798);
or U12275 (N_12275,N_10541,N_10868);
or U12276 (N_12276,N_10431,N_10624);
nand U12277 (N_12277,N_10263,N_11799);
xor U12278 (N_12278,N_11938,N_10095);
or U12279 (N_12279,N_10444,N_10159);
or U12280 (N_12280,N_10517,N_11935);
nor U12281 (N_12281,N_10986,N_10767);
or U12282 (N_12282,N_10464,N_11164);
nor U12283 (N_12283,N_11187,N_10715);
nand U12284 (N_12284,N_11893,N_10905);
xor U12285 (N_12285,N_11034,N_10625);
or U12286 (N_12286,N_11771,N_11006);
nor U12287 (N_12287,N_11754,N_10392);
nor U12288 (N_12288,N_11143,N_11059);
or U12289 (N_12289,N_11527,N_10826);
or U12290 (N_12290,N_10599,N_10297);
and U12291 (N_12291,N_11306,N_11347);
nor U12292 (N_12292,N_10396,N_11888);
xnor U12293 (N_12293,N_11745,N_10329);
nand U12294 (N_12294,N_11235,N_11564);
and U12295 (N_12295,N_10261,N_10480);
xor U12296 (N_12296,N_10099,N_11403);
nor U12297 (N_12297,N_11216,N_11976);
nand U12298 (N_12298,N_10094,N_11605);
or U12299 (N_12299,N_10851,N_11891);
xor U12300 (N_12300,N_10662,N_11994);
nand U12301 (N_12301,N_10765,N_10860);
or U12302 (N_12302,N_11273,N_10201);
or U12303 (N_12303,N_11962,N_11138);
and U12304 (N_12304,N_11052,N_11265);
xor U12305 (N_12305,N_11940,N_10514);
xor U12306 (N_12306,N_11636,N_11419);
xnor U12307 (N_12307,N_10911,N_10334);
and U12308 (N_12308,N_10647,N_11008);
nor U12309 (N_12309,N_10483,N_11900);
nor U12310 (N_12310,N_10012,N_10443);
xor U12311 (N_12311,N_11275,N_11708);
xor U12312 (N_12312,N_11075,N_10775);
and U12313 (N_12313,N_11036,N_10863);
or U12314 (N_12314,N_11066,N_10759);
nand U12315 (N_12315,N_10515,N_10891);
nor U12316 (N_12316,N_11810,N_10545);
xnor U12317 (N_12317,N_11168,N_11268);
xnor U12318 (N_12318,N_11576,N_10205);
xor U12319 (N_12319,N_10922,N_10727);
or U12320 (N_12320,N_11244,N_11549);
xor U12321 (N_12321,N_10129,N_10512);
and U12322 (N_12322,N_10250,N_11738);
xnor U12323 (N_12323,N_10557,N_10024);
nand U12324 (N_12324,N_11391,N_10147);
or U12325 (N_12325,N_11971,N_11190);
nor U12326 (N_12326,N_11722,N_11824);
nor U12327 (N_12327,N_10753,N_10888);
or U12328 (N_12328,N_11048,N_10038);
and U12329 (N_12329,N_11113,N_10323);
nor U12330 (N_12330,N_10477,N_10173);
or U12331 (N_12331,N_11144,N_11171);
nand U12332 (N_12332,N_11202,N_10916);
xor U12333 (N_12333,N_10466,N_10509);
and U12334 (N_12334,N_10608,N_11885);
and U12335 (N_12335,N_11567,N_11510);
or U12336 (N_12336,N_10110,N_11044);
xor U12337 (N_12337,N_10277,N_11227);
and U12338 (N_12338,N_10777,N_11393);
nand U12339 (N_12339,N_10835,N_11316);
nor U12340 (N_12340,N_10720,N_10428);
or U12341 (N_12341,N_10133,N_11860);
or U12342 (N_12342,N_11593,N_10687);
xor U12343 (N_12343,N_11237,N_10809);
nor U12344 (N_12344,N_10848,N_11750);
and U12345 (N_12345,N_10959,N_10467);
xor U12346 (N_12346,N_11909,N_10901);
or U12347 (N_12347,N_10769,N_11248);
xnor U12348 (N_12348,N_11525,N_10814);
nor U12349 (N_12349,N_11148,N_11609);
nand U12350 (N_12350,N_11610,N_10717);
nand U12351 (N_12351,N_10606,N_11776);
nand U12352 (N_12352,N_10617,N_10453);
or U12353 (N_12353,N_11646,N_11474);
xnor U12354 (N_12354,N_11274,N_10426);
and U12355 (N_12355,N_11728,N_11209);
or U12356 (N_12356,N_10433,N_11439);
nor U12357 (N_12357,N_10779,N_10317);
nor U12358 (N_12358,N_11358,N_11441);
nor U12359 (N_12359,N_10725,N_10927);
nand U12360 (N_12360,N_10761,N_11743);
xor U12361 (N_12361,N_10167,N_11485);
nor U12362 (N_12362,N_11203,N_10000);
nor U12363 (N_12363,N_11822,N_11442);
nor U12364 (N_12364,N_10877,N_10721);
or U12365 (N_12365,N_10019,N_10841);
nor U12366 (N_12366,N_11484,N_10846);
nand U12367 (N_12367,N_11886,N_10988);
nor U12368 (N_12368,N_11327,N_10590);
nor U12369 (N_12369,N_11132,N_10748);
or U12370 (N_12370,N_10876,N_11191);
nor U12371 (N_12371,N_11329,N_11179);
xor U12372 (N_12372,N_11236,N_11046);
or U12373 (N_12373,N_10910,N_11488);
and U12374 (N_12374,N_10945,N_10857);
and U12375 (N_12375,N_10387,N_11031);
and U12376 (N_12376,N_10361,N_11450);
nand U12377 (N_12377,N_10398,N_11807);
or U12378 (N_12378,N_11668,N_11505);
and U12379 (N_12379,N_11899,N_11769);
xnor U12380 (N_12380,N_11507,N_11984);
nor U12381 (N_12381,N_11263,N_10655);
nand U12382 (N_12382,N_10001,N_10182);
or U12383 (N_12383,N_10122,N_11267);
nor U12384 (N_12384,N_10252,N_11751);
xnor U12385 (N_12385,N_11999,N_11608);
or U12386 (N_12386,N_11339,N_10837);
nand U12387 (N_12387,N_10511,N_11724);
xnor U12388 (N_12388,N_11328,N_10836);
xor U12389 (N_12389,N_10080,N_11392);
and U12390 (N_12390,N_11407,N_10690);
and U12391 (N_12391,N_11359,N_11058);
and U12392 (N_12392,N_10124,N_10364);
or U12393 (N_12393,N_10724,N_11047);
nor U12394 (N_12394,N_11016,N_10703);
nor U12395 (N_12395,N_10680,N_11012);
nand U12396 (N_12396,N_10773,N_10365);
nor U12397 (N_12397,N_10487,N_11736);
and U12398 (N_12398,N_10534,N_11672);
xor U12399 (N_12399,N_10587,N_10243);
or U12400 (N_12400,N_11255,N_10950);
and U12401 (N_12401,N_11310,N_10560);
nand U12402 (N_12402,N_11963,N_11700);
and U12403 (N_12403,N_11307,N_10461);
xor U12404 (N_12404,N_11904,N_11600);
and U12405 (N_12405,N_11461,N_10884);
nand U12406 (N_12406,N_10042,N_10031);
nand U12407 (N_12407,N_10235,N_10299);
and U12408 (N_12408,N_11495,N_10704);
and U12409 (N_12409,N_11903,N_10879);
nand U12410 (N_12410,N_11444,N_10577);
nand U12411 (N_12411,N_11869,N_10148);
nor U12412 (N_12412,N_10643,N_11079);
xor U12413 (N_12413,N_10302,N_10912);
xor U12414 (N_12414,N_11487,N_11402);
and U12415 (N_12415,N_10384,N_10499);
xor U12416 (N_12416,N_11383,N_10309);
nor U12417 (N_12417,N_11720,N_10356);
and U12418 (N_12418,N_11465,N_10357);
and U12419 (N_12419,N_10786,N_11409);
xnor U12420 (N_12420,N_10314,N_10626);
nand U12421 (N_12421,N_10256,N_11481);
xor U12422 (N_12422,N_10674,N_11102);
nand U12423 (N_12423,N_11457,N_11097);
or U12424 (N_12424,N_11195,N_10258);
and U12425 (N_12425,N_10963,N_10609);
or U12426 (N_12426,N_11298,N_10178);
nand U12427 (N_12427,N_10926,N_10018);
nand U12428 (N_12428,N_11491,N_10716);
or U12429 (N_12429,N_10808,N_10832);
xor U12430 (N_12430,N_11875,N_10237);
nand U12431 (N_12431,N_10794,N_11167);
xnor U12432 (N_12432,N_10439,N_11054);
and U12433 (N_12433,N_10472,N_10015);
or U12434 (N_12434,N_11206,N_10538);
or U12435 (N_12435,N_11335,N_10897);
or U12436 (N_12436,N_10991,N_10714);
and U12437 (N_12437,N_11840,N_11477);
or U12438 (N_12438,N_10310,N_11513);
nand U12439 (N_12439,N_11568,N_11726);
or U12440 (N_12440,N_11846,N_10742);
or U12441 (N_12441,N_11142,N_11462);
nor U12442 (N_12442,N_11333,N_11867);
or U12443 (N_12443,N_10807,N_11486);
xor U12444 (N_12444,N_11243,N_11003);
or U12445 (N_12445,N_11658,N_11043);
xor U12446 (N_12446,N_11217,N_11100);
nor U12447 (N_12447,N_10158,N_10064);
and U12448 (N_12448,N_11344,N_10359);
nor U12449 (N_12449,N_11096,N_10301);
or U12450 (N_12450,N_11476,N_10563);
xnor U12451 (N_12451,N_11115,N_10254);
nand U12452 (N_12452,N_11808,N_11433);
or U12453 (N_12453,N_11432,N_11435);
xnor U12454 (N_12454,N_10496,N_11260);
and U12455 (N_12455,N_10586,N_10349);
or U12456 (N_12456,N_10782,N_10854);
or U12457 (N_12457,N_11801,N_10022);
and U12458 (N_12458,N_10500,N_11800);
nor U12459 (N_12459,N_10711,N_11850);
nor U12460 (N_12460,N_11204,N_10805);
nor U12461 (N_12461,N_11775,N_10955);
nand U12462 (N_12462,N_10953,N_10739);
nand U12463 (N_12463,N_10688,N_10695);
or U12464 (N_12464,N_11400,N_10958);
and U12465 (N_12465,N_11014,N_11587);
or U12466 (N_12466,N_11186,N_10874);
xor U12467 (N_12467,N_10738,N_10032);
and U12468 (N_12468,N_11473,N_11779);
xor U12469 (N_12469,N_10468,N_10632);
or U12470 (N_12470,N_11680,N_11398);
nor U12471 (N_12471,N_10078,N_11251);
nand U12472 (N_12472,N_10493,N_10949);
or U12473 (N_12473,N_11882,N_11996);
nand U12474 (N_12474,N_11723,N_11426);
nand U12475 (N_12475,N_11429,N_10343);
nor U12476 (N_12476,N_11635,N_10198);
xnor U12477 (N_12477,N_10962,N_11556);
nand U12478 (N_12478,N_10315,N_11588);
or U12479 (N_12479,N_11181,N_10062);
and U12480 (N_12480,N_11437,N_10929);
xnor U12481 (N_12481,N_11968,N_11543);
or U12482 (N_12482,N_10251,N_10088);
nor U12483 (N_12483,N_10644,N_11196);
xnor U12484 (N_12484,N_11531,N_11777);
xor U12485 (N_12485,N_11812,N_10734);
or U12486 (N_12486,N_11081,N_10407);
or U12487 (N_12487,N_10758,N_11380);
nor U12488 (N_12488,N_11932,N_11301);
or U12489 (N_12489,N_10693,N_11862);
xor U12490 (N_12490,N_11420,N_11033);
and U12491 (N_12491,N_11898,N_11655);
xor U12492 (N_12492,N_10675,N_10594);
nand U12493 (N_12493,N_11336,N_10941);
or U12494 (N_12494,N_10096,N_10676);
nor U12495 (N_12495,N_10089,N_11849);
nand U12496 (N_12496,N_10591,N_11421);
or U12497 (N_12497,N_11688,N_10614);
nand U12498 (N_12498,N_10634,N_10306);
and U12499 (N_12499,N_11965,N_11974);
nor U12500 (N_12500,N_11050,N_10210);
or U12501 (N_12501,N_11590,N_11628);
xnor U12502 (N_12502,N_10369,N_11586);
or U12503 (N_12503,N_11337,N_10896);
or U12504 (N_12504,N_11158,N_11788);
nor U12505 (N_12505,N_11559,N_10185);
nand U12506 (N_12506,N_10162,N_11103);
and U12507 (N_12507,N_11682,N_11784);
nor U12508 (N_12508,N_10875,N_10171);
nand U12509 (N_12509,N_10046,N_10973);
or U12510 (N_12510,N_10700,N_11730);
and U12511 (N_12511,N_10822,N_11219);
nand U12512 (N_12512,N_11345,N_10938);
nand U12513 (N_12513,N_11561,N_10829);
or U12514 (N_12514,N_10119,N_10640);
or U12515 (N_12515,N_11390,N_11705);
or U12516 (N_12516,N_10283,N_11453);
xor U12517 (N_12517,N_10213,N_11319);
xnor U12518 (N_12518,N_11767,N_10040);
nand U12519 (N_12519,N_11657,N_10280);
xor U12520 (N_12520,N_11320,N_10268);
and U12521 (N_12521,N_11418,N_11305);
or U12522 (N_12522,N_11604,N_11770);
xnor U12523 (N_12523,N_11456,N_10957);
or U12524 (N_12524,N_10161,N_10390);
xor U12525 (N_12525,N_11483,N_11532);
and U12526 (N_12526,N_11026,N_11766);
nor U12527 (N_12527,N_10627,N_11362);
xor U12528 (N_12528,N_10964,N_11581);
nor U12529 (N_12529,N_10696,N_10967);
or U12530 (N_12530,N_10537,N_10348);
and U12531 (N_12531,N_10755,N_10442);
and U12532 (N_12532,N_10338,N_10793);
or U12533 (N_12533,N_10421,N_11990);
and U12534 (N_12534,N_10940,N_11389);
or U12535 (N_12535,N_11575,N_10994);
xnor U12536 (N_12536,N_11311,N_11953);
nor U12537 (N_12537,N_11166,N_11112);
nor U12538 (N_12538,N_10831,N_10055);
nand U12539 (N_12539,N_11707,N_11123);
nand U12540 (N_12540,N_10976,N_10571);
nor U12541 (N_12541,N_10300,N_11240);
or U12542 (N_12542,N_11842,N_10479);
xor U12543 (N_12543,N_11828,N_10376);
xnor U12544 (N_12544,N_11690,N_10615);
nor U12545 (N_12545,N_10651,N_11787);
and U12546 (N_12546,N_10569,N_10637);
and U12547 (N_12547,N_10249,N_11272);
xnor U12548 (N_12548,N_11446,N_10014);
xor U12549 (N_12549,N_11773,N_10473);
and U12550 (N_12550,N_11340,N_10838);
nor U12551 (N_12551,N_11459,N_10112);
xnor U12552 (N_12552,N_11825,N_11772);
nor U12553 (N_12553,N_10353,N_11654);
and U12554 (N_12554,N_11366,N_11249);
nand U12555 (N_12555,N_10195,N_10136);
and U12556 (N_12556,N_11330,N_11710);
xnor U12557 (N_12557,N_10346,N_11408);
and U12558 (N_12558,N_10692,N_11839);
and U12559 (N_12559,N_10415,N_11083);
nor U12560 (N_12560,N_11009,N_11864);
nor U12561 (N_12561,N_11515,N_11637);
or U12562 (N_12562,N_10436,N_10430);
or U12563 (N_12563,N_11578,N_11107);
and U12564 (N_12564,N_11141,N_11626);
nor U12565 (N_12565,N_10165,N_10948);
xor U12566 (N_12566,N_11295,N_11431);
nor U12567 (N_12567,N_10106,N_10255);
nand U12568 (N_12568,N_11341,N_10906);
and U12569 (N_12569,N_10718,N_11541);
or U12570 (N_12570,N_10199,N_10501);
nor U12571 (N_12571,N_11597,N_10242);
nor U12572 (N_12572,N_11215,N_10219);
xnor U12573 (N_12573,N_10997,N_10741);
xor U12574 (N_12574,N_10234,N_10815);
nand U12575 (N_12575,N_11737,N_11121);
nand U12576 (N_12576,N_11011,N_10247);
nand U12577 (N_12577,N_11198,N_11833);
xor U12578 (N_12578,N_11351,N_11762);
xor U12579 (N_12579,N_10904,N_10081);
or U12580 (N_12580,N_11194,N_10970);
xnor U12581 (N_12581,N_10978,N_10344);
or U12582 (N_12582,N_10017,N_11698);
and U12583 (N_12583,N_11831,N_11147);
or U12584 (N_12584,N_11023,N_11502);
nor U12585 (N_12585,N_11343,N_10045);
or U12586 (N_12586,N_10211,N_10522);
and U12587 (N_12587,N_10611,N_11379);
nor U12588 (N_12588,N_10075,N_10620);
or U12589 (N_12589,N_11897,N_10589);
nand U12590 (N_12590,N_11111,N_11673);
xnor U12591 (N_12591,N_10400,N_11847);
nand U12592 (N_12592,N_10004,N_11565);
nand U12593 (N_12593,N_11040,N_10134);
and U12594 (N_12594,N_10665,N_11583);
xor U12595 (N_12595,N_10979,N_11931);
nand U12596 (N_12596,N_11768,N_10130);
nand U12597 (N_12597,N_10446,N_10292);
xor U12598 (N_12598,N_10605,N_11765);
nand U12599 (N_12599,N_10102,N_11683);
or U12600 (N_12600,N_11856,N_11625);
nor U12601 (N_12601,N_10061,N_11920);
or U12602 (N_12602,N_11753,N_11859);
or U12603 (N_12603,N_11269,N_11218);
nand U12604 (N_12604,N_11930,N_10990);
xor U12605 (N_12605,N_10154,N_11675);
or U12606 (N_12606,N_10033,N_10079);
and U12607 (N_12607,N_10286,N_11239);
nor U12608 (N_12608,N_10619,N_10149);
nand U12609 (N_12609,N_11297,N_10712);
or U12610 (N_12610,N_11018,N_11266);
or U12611 (N_12611,N_11382,N_10542);
nand U12612 (N_12612,N_10269,N_10529);
xnor U12613 (N_12613,N_11261,N_11863);
xnor U12614 (N_12614,N_11618,N_10981);
nand U12615 (N_12615,N_10476,N_10048);
and U12616 (N_12616,N_10764,N_11782);
and U12617 (N_12617,N_10326,N_11661);
or U12618 (N_12618,N_11397,N_10037);
nand U12619 (N_12619,N_10010,N_11620);
nand U12620 (N_12620,N_11304,N_11331);
xor U12621 (N_12621,N_11878,N_10190);
nor U12622 (N_12622,N_11135,N_11535);
nor U12623 (N_12623,N_11950,N_10118);
or U12624 (N_12624,N_11145,N_10239);
nand U12625 (N_12625,N_11718,N_10823);
and U12626 (N_12626,N_11601,N_10686);
nor U12627 (N_12627,N_10628,N_11440);
nor U12628 (N_12628,N_11522,N_11078);
nand U12629 (N_12629,N_11291,N_10117);
xor U12630 (N_12630,N_10989,N_10915);
and U12631 (N_12631,N_10658,N_10332);
and U12632 (N_12632,N_10355,N_11060);
or U12633 (N_12633,N_11927,N_10996);
and U12634 (N_12634,N_10241,N_11172);
xnor U12635 (N_12635,N_10995,N_10462);
nand U12636 (N_12636,N_10900,N_10215);
or U12637 (N_12637,N_11428,N_10097);
and U12638 (N_12638,N_10230,N_10054);
nand U12639 (N_12639,N_10084,N_11279);
nand U12640 (N_12640,N_10385,N_11827);
nor U12641 (N_12641,N_10287,N_11954);
and U12642 (N_12642,N_10580,N_10740);
nor U12643 (N_12643,N_10183,N_10819);
xor U12644 (N_12644,N_10020,N_10330);
or U12645 (N_12645,N_11623,N_11296);
nor U12646 (N_12646,N_10867,N_11232);
nand U12647 (N_12647,N_10386,N_10266);
nand U12648 (N_12648,N_11553,N_10494);
xor U12649 (N_12649,N_10683,N_10914);
nor U12650 (N_12650,N_10181,N_10872);
xor U12651 (N_12651,N_11064,N_11017);
xnor U12652 (N_12652,N_10568,N_10925);
or U12653 (N_12653,N_11702,N_11374);
or U12654 (N_12654,N_10366,N_10952);
xnor U12655 (N_12655,N_11154,N_11611);
or U12656 (N_12656,N_11641,N_11318);
nor U12657 (N_12657,N_10481,N_11806);
or U12658 (N_12658,N_11691,N_11109);
and U12659 (N_12659,N_11245,N_11129);
nor U12660 (N_12660,N_10418,N_11095);
nor U12661 (N_12661,N_10785,N_11030);
and U12662 (N_12662,N_10214,N_11873);
xor U12663 (N_12663,N_10600,N_10093);
nor U12664 (N_12664,N_10049,N_11056);
or U12665 (N_12665,N_10971,N_11406);
and U12666 (N_12666,N_11055,N_11385);
nand U12667 (N_12667,N_11523,N_11836);
nand U12668 (N_12668,N_10641,N_11281);
nor U12669 (N_12669,N_10067,N_10295);
xnor U12670 (N_12670,N_10026,N_10009);
nor U12671 (N_12671,N_10810,N_11119);
or U12672 (N_12672,N_10799,N_10452);
nor U12673 (N_12673,N_10597,N_11193);
nor U12674 (N_12674,N_11458,N_10812);
nor U12675 (N_12675,N_10845,N_11520);
xnor U12676 (N_12676,N_10333,N_10410);
or U12677 (N_12677,N_11499,N_11844);
nand U12678 (N_12678,N_10543,N_10016);
nor U12679 (N_12679,N_10484,N_11967);
or U12680 (N_12680,N_11959,N_10327);
nor U12681 (N_12681,N_11619,N_11816);
or U12682 (N_12682,N_10248,N_11892);
nor U12683 (N_12683,N_10546,N_11425);
xnor U12684 (N_12684,N_10678,N_11482);
xor U12685 (N_12685,N_10965,N_10495);
and U12686 (N_12686,N_10240,N_11134);
or U12687 (N_12687,N_11667,N_11509);
xor U12688 (N_12688,N_11354,N_11157);
nor U12689 (N_12689,N_11566,N_11870);
nand U12690 (N_12690,N_10169,N_10108);
nand U12691 (N_12691,N_10830,N_10774);
and U12692 (N_12692,N_10140,N_11802);
xnor U12693 (N_12693,N_10394,N_11858);
nand U12694 (N_12694,N_11969,N_11416);
nand U12695 (N_12695,N_11952,N_11019);
and U12696 (N_12696,N_10728,N_11589);
nor U12697 (N_12697,N_10265,N_10582);
nor U12698 (N_12698,N_10820,N_11936);
and U12699 (N_12699,N_10920,N_10284);
nand U12700 (N_12700,N_10459,N_11290);
or U12701 (N_12701,N_11685,N_10307);
nand U12702 (N_12702,N_10059,N_11518);
and U12703 (N_12703,N_10224,N_10677);
and U12704 (N_12704,N_11894,N_10321);
or U12705 (N_12705,N_11411,N_10289);
nor U12706 (N_12706,N_11104,N_11741);
nand U12707 (N_12707,N_10883,N_11160);
or U12708 (N_12708,N_11760,N_10698);
nor U12709 (N_12709,N_11289,N_10630);
nor U12710 (N_12710,N_11562,N_10128);
nor U12711 (N_12711,N_11150,N_10006);
and U12712 (N_12712,N_10707,N_11368);
xnor U12713 (N_12713,N_10422,N_10264);
or U12714 (N_12714,N_11504,N_11128);
and U12715 (N_12715,N_10238,N_10153);
and U12716 (N_12716,N_10028,N_10649);
and U12717 (N_12717,N_11226,N_11838);
xnor U12718 (N_12718,N_10116,N_11876);
and U12719 (N_12719,N_10109,N_10368);
nor U12720 (N_12720,N_11287,N_11921);
and U12721 (N_12721,N_10919,N_11761);
xor U12722 (N_12722,N_10549,N_10196);
nand U12723 (N_12723,N_10029,N_11853);
or U12724 (N_12724,N_11480,N_11225);
or U12725 (N_12725,N_11234,N_10595);
and U12726 (N_12726,N_11696,N_11763);
or U12727 (N_12727,N_11580,N_10934);
and U12728 (N_12728,N_11746,N_11820);
and U12729 (N_12729,N_11725,N_10813);
and U12730 (N_12730,N_11756,N_11638);
nor U12731 (N_12731,N_11905,N_11572);
or U12732 (N_12732,N_11027,N_11252);
or U12733 (N_12733,N_10510,N_11246);
or U12734 (N_12734,N_10750,N_10192);
xnor U12735 (N_12735,N_11961,N_10834);
nand U12736 (N_12736,N_10811,N_11598);
xor U12737 (N_12737,N_10144,N_10930);
nor U12738 (N_12738,N_11595,N_10497);
and U12739 (N_12739,N_11666,N_11731);
or U12740 (N_12740,N_10573,N_10723);
or U12741 (N_12741,N_11536,N_11169);
xor U12742 (N_12742,N_10592,N_11678);
nand U12743 (N_12743,N_11631,N_11001);
and U12744 (N_12744,N_10311,N_11571);
nand U12745 (N_12745,N_10946,N_10902);
or U12746 (N_12746,N_11676,N_10163);
or U12747 (N_12747,N_11438,N_11152);
nor U12748 (N_12748,N_10816,N_11560);
or U12749 (N_12749,N_10670,N_11997);
or U12750 (N_12750,N_11313,N_11182);
xor U12751 (N_12751,N_11949,N_11512);
xor U12752 (N_12752,N_10797,N_11241);
or U12753 (N_12753,N_11080,N_11699);
nor U12754 (N_12754,N_11061,N_10673);
xnor U12755 (N_12755,N_10058,N_10298);
nand U12756 (N_12756,N_10878,N_10146);
and U12757 (N_12757,N_10873,N_11094);
or U12758 (N_12758,N_11796,N_11681);
and U12759 (N_12759,N_10005,N_10208);
or U12760 (N_12760,N_11714,N_11642);
and U12761 (N_12761,N_11302,N_11656);
and U12762 (N_12762,N_11131,N_11918);
or U12763 (N_12763,N_10575,N_11467);
nor U12764 (N_12764,N_11693,N_10290);
or U12765 (N_12765,N_11277,N_10325);
nand U12766 (N_12766,N_11639,N_10257);
or U12767 (N_12767,N_11222,N_11715);
or U12768 (N_12768,N_10103,N_11089);
or U12769 (N_12769,N_10572,N_11367);
and U12770 (N_12770,N_11719,N_11149);
and U12771 (N_12771,N_11664,N_11069);
or U12772 (N_12772,N_10918,N_10083);
nor U12773 (N_12773,N_11545,N_11466);
xor U12774 (N_12774,N_11735,N_10827);
nor U12775 (N_12775,N_11826,N_10139);
nor U12776 (N_12776,N_10197,N_11401);
and U12777 (N_12777,N_10540,N_10554);
nand U12778 (N_12778,N_11238,N_11348);
xnor U12779 (N_12779,N_11855,N_11088);
and U12780 (N_12780,N_10399,N_10363);
or U12781 (N_12781,N_11879,N_11155);
nor U12782 (N_12782,N_11496,N_11712);
and U12783 (N_12783,N_10757,N_10425);
or U12784 (N_12784,N_11514,N_11257);
nand U12785 (N_12785,N_10726,N_11021);
nand U12786 (N_12786,N_11342,N_11394);
nor U12787 (N_12787,N_11212,N_11811);
nor U12788 (N_12788,N_10559,N_10374);
or U12789 (N_12789,N_10073,N_11005);
and U12790 (N_12790,N_10581,N_11068);
nor U12791 (N_12791,N_10942,N_10977);
or U12792 (N_12792,N_10646,N_11902);
nor U12793 (N_12793,N_11472,N_11285);
xor U12794 (N_12794,N_10610,N_11910);
nor U12795 (N_12795,N_11228,N_11747);
xnor U12796 (N_12796,N_11180,N_11881);
or U12797 (N_12797,N_10633,N_11537);
nand U12798 (N_12798,N_10262,N_10666);
xor U12799 (N_12799,N_11524,N_10445);
nor U12800 (N_12800,N_11647,N_11684);
nand U12801 (N_12801,N_11992,N_11709);
xnor U12802 (N_12802,N_11300,N_10535);
nor U12803 (N_12803,N_11852,N_11007);
and U12804 (N_12804,N_11395,N_11651);
xnor U12805 (N_12805,N_10982,N_11455);
or U12806 (N_12806,N_10968,N_11957);
nor U12807 (N_12807,N_10733,N_11805);
nand U12808 (N_12808,N_10856,N_10516);
and U12809 (N_12809,N_11004,N_11814);
xnor U12810 (N_12810,N_10113,N_10253);
and U12811 (N_12811,N_10417,N_11369);
xnor U12812 (N_12812,N_10388,N_10470);
nand U12813 (N_12813,N_10336,N_10100);
and U12814 (N_12814,N_11874,N_11706);
nand U12815 (N_12815,N_10375,N_10578);
xor U12816 (N_12816,N_10886,N_10566);
or U12817 (N_12817,N_11640,N_11200);
or U12818 (N_12818,N_11960,N_11632);
nor U12819 (N_12819,N_11596,N_10404);
nor U12820 (N_12820,N_10457,N_11176);
xor U12821 (N_12821,N_10288,N_10583);
and U12822 (N_12822,N_10756,N_11945);
or U12823 (N_12823,N_10576,N_10596);
or U12824 (N_12824,N_11086,N_10402);
nand U12825 (N_12825,N_11384,N_10138);
or U12826 (N_12826,N_11264,N_10530);
and U12827 (N_12827,N_11621,N_10188);
nand U12828 (N_12828,N_11072,N_11797);
or U12829 (N_12829,N_10231,N_10441);
or U12830 (N_12830,N_10639,N_10435);
and U12831 (N_12831,N_11189,N_10143);
nor U12832 (N_12832,N_10226,N_11926);
xnor U12833 (N_12833,N_11065,N_10783);
xor U12834 (N_12834,N_10533,N_10372);
nor U12835 (N_12835,N_10890,N_10645);
xnor U12836 (N_12836,N_11713,N_10795);
and U12837 (N_12837,N_11283,N_10104);
nor U12838 (N_12838,N_11002,N_10705);
xor U12839 (N_12839,N_10694,N_11230);
or U12840 (N_12840,N_11309,N_10414);
and U12841 (N_12841,N_10072,N_10778);
nor U12842 (N_12842,N_11024,N_11288);
nor U12843 (N_12843,N_11819,N_10172);
or U12844 (N_12844,N_11122,N_10570);
and U12845 (N_12845,N_10281,N_10174);
nand U12846 (N_12846,N_10855,N_11519);
xnor U12847 (N_12847,N_10413,N_10719);
and U12848 (N_12848,N_11928,N_10520);
and U12849 (N_12849,N_10532,N_10987);
or U12850 (N_12850,N_10601,N_11665);
xnor U12851 (N_12851,N_11697,N_10207);
and U12852 (N_12852,N_11783,N_10246);
xnor U12853 (N_12853,N_10550,N_10092);
nor U12854 (N_12854,N_11223,N_11872);
and U12855 (N_12855,N_10844,N_11964);
and U12856 (N_12856,N_10772,N_10682);
nor U12857 (N_12857,N_11126,N_10613);
nand U12858 (N_12858,N_10804,N_11809);
and U12859 (N_12859,N_10463,N_10186);
and U12860 (N_12860,N_11192,N_10974);
or U12861 (N_12861,N_11794,N_10842);
or U12862 (N_12862,N_11978,N_11901);
xor U12863 (N_12863,N_11410,N_10790);
nand U12864 (N_12864,N_10839,N_10077);
nand U12865 (N_12865,N_10137,N_11975);
nor U12866 (N_12866,N_10735,N_11173);
or U12867 (N_12867,N_10021,N_10858);
nand U12868 (N_12868,N_10776,N_10943);
or U12869 (N_12869,N_10556,N_11550);
nor U12870 (N_12870,N_11644,N_11544);
nand U12871 (N_12871,N_11703,N_10166);
xor U12872 (N_12872,N_10406,N_10030);
nand U12873 (N_12873,N_11542,N_10881);
and U12874 (N_12874,N_10013,N_10697);
or U12875 (N_12875,N_11929,N_11695);
xor U12876 (N_12876,N_11895,N_10331);
xnor U12877 (N_12877,N_11848,N_10456);
xor U12878 (N_12878,N_11025,N_10419);
nand U12879 (N_12879,N_10864,N_10335);
nor U12880 (N_12880,N_11889,N_10781);
and U12881 (N_12881,N_10373,N_10893);
nand U12882 (N_12882,N_11614,N_11789);
xor U12883 (N_12883,N_10491,N_11185);
nor U12884 (N_12884,N_11704,N_10403);
nand U12885 (N_12885,N_10142,N_10141);
nand U12886 (N_12886,N_10126,N_11294);
and U12887 (N_12887,N_10041,N_11843);
nor U12888 (N_12888,N_10661,N_11091);
xor U12889 (N_12889,N_10043,N_10107);
or U12890 (N_12890,N_11468,N_10291);
xnor U12891 (N_12891,N_11452,N_10175);
xnor U12892 (N_12892,N_10382,N_11569);
and U12893 (N_12893,N_11032,N_10324);
or U12894 (N_12894,N_11871,N_11493);
nand U12895 (N_12895,N_10763,N_10923);
or U12896 (N_12896,N_10602,N_10604);
nor U12897 (N_12897,N_10551,N_10506);
nor U12898 (N_12898,N_11077,N_11130);
or U12899 (N_12899,N_11471,N_10931);
or U12900 (N_12900,N_10588,N_10796);
or U12901 (N_12901,N_11346,N_10053);
nand U12902 (N_12902,N_10121,N_11939);
nor U12903 (N_12903,N_10681,N_10825);
and U12904 (N_12904,N_11214,N_11622);
xnor U12905 (N_12905,N_11153,N_11312);
nor U12906 (N_12906,N_10504,N_11830);
xnor U12907 (N_12907,N_11981,N_10526);
and U12908 (N_12908,N_10859,N_11757);
or U12909 (N_12909,N_10539,N_11207);
nor U12910 (N_12910,N_11049,N_11923);
or U12911 (N_12911,N_10090,N_10548);
nand U12912 (N_12912,N_10209,N_10519);
and U12913 (N_12913,N_11165,N_10245);
nor U12914 (N_12914,N_10684,N_10622);
and U12915 (N_12915,N_11254,N_11073);
nor U12916 (N_12916,N_10189,N_10150);
xnor U12917 (N_12917,N_10105,N_11370);
nand U12918 (N_12918,N_11259,N_11817);
nand U12919 (N_12919,N_10420,N_10393);
nand U12920 (N_12920,N_10544,N_10951);
nand U12921 (N_12921,N_11136,N_11308);
nand U12922 (N_12922,N_11602,N_10152);
or U12923 (N_12923,N_11946,N_10840);
nor U12924 (N_12924,N_10492,N_10730);
or U12925 (N_12925,N_10176,N_11977);
nor U12926 (N_12926,N_10547,N_10880);
nand U12927 (N_12927,N_10391,N_11577);
nor U12928 (N_12928,N_11177,N_11734);
nor U12929 (N_12929,N_11616,N_10650);
xnor U12930 (N_12930,N_11742,N_10508);
nor U12931 (N_12931,N_11786,N_11037);
nor U12932 (N_12932,N_11890,N_10027);
nor U12933 (N_12933,N_10044,N_10405);
nand U12934 (N_12934,N_10567,N_10562);
and U12935 (N_12935,N_10593,N_11284);
nand U12936 (N_12936,N_10184,N_10792);
or U12937 (N_12937,N_10817,N_10087);
and U12938 (N_12938,N_10762,N_11414);
or U12939 (N_12939,N_11082,N_11521);
nor U12940 (N_12940,N_10056,N_10066);
nand U12941 (N_12941,N_10894,N_10294);
nor U12942 (N_12942,N_11211,N_11530);
nand U12943 (N_12943,N_10151,N_10091);
xor U12944 (N_12944,N_10132,N_11338);
nand U12945 (N_12945,N_10177,N_11041);
nand U12946 (N_12946,N_11552,N_10485);
nand U12947 (N_12947,N_10074,N_11998);
or U12948 (N_12948,N_10486,N_10668);
xor U12949 (N_12949,N_11373,N_10885);
and U12950 (N_12950,N_11381,N_11253);
xor U12951 (N_12951,N_10474,N_10536);
and U12952 (N_12952,N_11372,N_11983);
or U12953 (N_12953,N_10699,N_10671);
or U12954 (N_12954,N_11781,N_11970);
xor U12955 (N_12955,N_11574,N_11790);
xor U12956 (N_12956,N_11793,N_10098);
or U12957 (N_12957,N_11386,N_11832);
nand U12958 (N_12958,N_11070,N_11350);
xnor U12959 (N_12959,N_11133,N_10145);
nand U12960 (N_12960,N_10204,N_11837);
or U12961 (N_12961,N_10218,N_11028);
xor U12962 (N_12962,N_10784,N_10993);
or U12963 (N_12963,N_11042,N_10892);
nand U12964 (N_12964,N_10434,N_10273);
xnor U12965 (N_12965,N_10513,N_10969);
or U12966 (N_12966,N_11991,N_11365);
or U12967 (N_12967,N_10944,N_10903);
and U12968 (N_12968,N_11139,N_11360);
nand U12969 (N_12969,N_11271,N_11555);
nor U12970 (N_12970,N_10328,N_11108);
nor U12971 (N_12971,N_10202,N_11178);
or U12972 (N_12972,N_11944,N_11517);
nor U12973 (N_12973,N_10898,N_10956);
nand U12974 (N_12974,N_11233,N_11538);
nor U12975 (N_12975,N_10316,N_10227);
and U12976 (N_12976,N_11922,N_10618);
nor U12977 (N_12977,N_10271,N_11687);
and U12978 (N_12978,N_10932,N_11884);
and U12979 (N_12979,N_10389,N_11110);
nor U12980 (N_12980,N_11966,N_10527);
and U12981 (N_12981,N_10085,N_11140);
xnor U12982 (N_12982,N_11511,N_11652);
or U12983 (N_12983,N_10025,N_11434);
xnor U12984 (N_12984,N_11363,N_11711);
xnor U12985 (N_12985,N_10225,N_11528);
nor U12986 (N_12986,N_10180,N_11270);
nand U12987 (N_12987,N_10780,N_11993);
nand U12988 (N_12988,N_11649,N_11101);
or U12989 (N_12989,N_11633,N_10111);
xor U12990 (N_12990,N_10553,N_11114);
xnor U12991 (N_12991,N_10579,N_11184);
and U12992 (N_12992,N_10432,N_11349);
or U12993 (N_12993,N_11749,N_10975);
and U12994 (N_12994,N_11764,N_11740);
nand U12995 (N_12995,N_11866,N_11322);
nor U12996 (N_12996,N_11494,N_11417);
and U12997 (N_12997,N_11547,N_11303);
and U12998 (N_12998,N_10908,N_11325);
xnor U12999 (N_12999,N_10936,N_10584);
nand U13000 (N_13000,N_10351,N_11400);
nand U13001 (N_13001,N_10953,N_11880);
nand U13002 (N_13002,N_10388,N_10237);
nand U13003 (N_13003,N_11190,N_10510);
nor U13004 (N_13004,N_11412,N_11503);
and U13005 (N_13005,N_11591,N_11055);
nand U13006 (N_13006,N_10568,N_11234);
nand U13007 (N_13007,N_11569,N_11414);
and U13008 (N_13008,N_11016,N_11693);
or U13009 (N_13009,N_10647,N_11010);
or U13010 (N_13010,N_11540,N_11312);
nand U13011 (N_13011,N_10701,N_10622);
or U13012 (N_13012,N_11943,N_10344);
xor U13013 (N_13013,N_10788,N_10029);
nand U13014 (N_13014,N_10218,N_10909);
and U13015 (N_13015,N_10118,N_10087);
nand U13016 (N_13016,N_10417,N_10048);
nor U13017 (N_13017,N_10387,N_11154);
and U13018 (N_13018,N_10855,N_11323);
xnor U13019 (N_13019,N_11054,N_11013);
or U13020 (N_13020,N_11765,N_11602);
or U13021 (N_13021,N_11200,N_11064);
or U13022 (N_13022,N_11657,N_10301);
or U13023 (N_13023,N_10011,N_11912);
nor U13024 (N_13024,N_10545,N_11471);
nor U13025 (N_13025,N_10798,N_10470);
nor U13026 (N_13026,N_11881,N_10338);
nand U13027 (N_13027,N_11457,N_11660);
nor U13028 (N_13028,N_10838,N_11099);
and U13029 (N_13029,N_10652,N_11710);
nand U13030 (N_13030,N_11870,N_11644);
or U13031 (N_13031,N_11811,N_10000);
or U13032 (N_13032,N_10739,N_11874);
and U13033 (N_13033,N_10903,N_11521);
xor U13034 (N_13034,N_11805,N_11099);
nor U13035 (N_13035,N_10537,N_11355);
nor U13036 (N_13036,N_11574,N_10539);
xnor U13037 (N_13037,N_11403,N_11167);
and U13038 (N_13038,N_10226,N_10578);
nor U13039 (N_13039,N_11273,N_11889);
nand U13040 (N_13040,N_11817,N_10408);
or U13041 (N_13041,N_11805,N_10234);
xor U13042 (N_13042,N_10015,N_10045);
and U13043 (N_13043,N_11916,N_11537);
nand U13044 (N_13044,N_10830,N_10992);
nor U13045 (N_13045,N_11465,N_11409);
xnor U13046 (N_13046,N_10786,N_10809);
nor U13047 (N_13047,N_10929,N_11443);
or U13048 (N_13048,N_11484,N_11935);
and U13049 (N_13049,N_11697,N_10730);
and U13050 (N_13050,N_10830,N_11504);
or U13051 (N_13051,N_10399,N_10461);
or U13052 (N_13052,N_11689,N_10895);
and U13053 (N_13053,N_11743,N_10758);
and U13054 (N_13054,N_10001,N_11824);
nand U13055 (N_13055,N_11179,N_10652);
and U13056 (N_13056,N_10340,N_10352);
nor U13057 (N_13057,N_10420,N_10198);
or U13058 (N_13058,N_11433,N_10731);
or U13059 (N_13059,N_11367,N_11321);
and U13060 (N_13060,N_10735,N_11901);
nor U13061 (N_13061,N_11466,N_11638);
xnor U13062 (N_13062,N_11620,N_10922);
nand U13063 (N_13063,N_11140,N_11560);
nand U13064 (N_13064,N_10968,N_11232);
and U13065 (N_13065,N_10752,N_10086);
nand U13066 (N_13066,N_10419,N_10542);
or U13067 (N_13067,N_10458,N_11778);
or U13068 (N_13068,N_10855,N_11701);
and U13069 (N_13069,N_11795,N_11709);
xnor U13070 (N_13070,N_10527,N_10042);
or U13071 (N_13071,N_10538,N_10044);
xor U13072 (N_13072,N_10220,N_10090);
xor U13073 (N_13073,N_11581,N_10255);
and U13074 (N_13074,N_10099,N_10272);
and U13075 (N_13075,N_10099,N_11406);
and U13076 (N_13076,N_11318,N_10471);
nand U13077 (N_13077,N_11812,N_11747);
nor U13078 (N_13078,N_10717,N_11060);
nor U13079 (N_13079,N_10452,N_10507);
xnor U13080 (N_13080,N_11079,N_10845);
nand U13081 (N_13081,N_10046,N_11411);
or U13082 (N_13082,N_10941,N_11310);
nor U13083 (N_13083,N_11065,N_11102);
xnor U13084 (N_13084,N_10869,N_11089);
and U13085 (N_13085,N_10432,N_10323);
xor U13086 (N_13086,N_10513,N_11125);
nor U13087 (N_13087,N_10918,N_11652);
or U13088 (N_13088,N_11201,N_11812);
and U13089 (N_13089,N_11658,N_10705);
and U13090 (N_13090,N_11296,N_11611);
xnor U13091 (N_13091,N_11755,N_10775);
nand U13092 (N_13092,N_11725,N_11016);
nand U13093 (N_13093,N_10371,N_11841);
nand U13094 (N_13094,N_11924,N_10629);
nand U13095 (N_13095,N_10302,N_11162);
and U13096 (N_13096,N_11159,N_10091);
and U13097 (N_13097,N_10302,N_10376);
xor U13098 (N_13098,N_11687,N_11591);
and U13099 (N_13099,N_10913,N_11614);
and U13100 (N_13100,N_10280,N_11825);
or U13101 (N_13101,N_10846,N_10839);
nand U13102 (N_13102,N_10822,N_10375);
xor U13103 (N_13103,N_10136,N_10729);
xnor U13104 (N_13104,N_10279,N_11116);
nor U13105 (N_13105,N_11894,N_10407);
xor U13106 (N_13106,N_11271,N_11630);
or U13107 (N_13107,N_11167,N_11307);
nand U13108 (N_13108,N_10165,N_10181);
nor U13109 (N_13109,N_11089,N_10546);
or U13110 (N_13110,N_10821,N_10630);
xor U13111 (N_13111,N_11483,N_10441);
and U13112 (N_13112,N_11441,N_11825);
xnor U13113 (N_13113,N_11070,N_11034);
nand U13114 (N_13114,N_11610,N_10379);
or U13115 (N_13115,N_10422,N_10839);
xor U13116 (N_13116,N_11587,N_11753);
and U13117 (N_13117,N_10092,N_10473);
nand U13118 (N_13118,N_10037,N_10711);
nand U13119 (N_13119,N_11498,N_11713);
nor U13120 (N_13120,N_10707,N_11412);
xnor U13121 (N_13121,N_10891,N_10168);
and U13122 (N_13122,N_10975,N_11435);
xor U13123 (N_13123,N_10550,N_10002);
nand U13124 (N_13124,N_11100,N_11471);
nand U13125 (N_13125,N_10384,N_11459);
nand U13126 (N_13126,N_10504,N_11761);
nand U13127 (N_13127,N_10978,N_10092);
xor U13128 (N_13128,N_10328,N_11409);
xnor U13129 (N_13129,N_11303,N_10440);
or U13130 (N_13130,N_10174,N_11843);
nand U13131 (N_13131,N_11550,N_11295);
or U13132 (N_13132,N_10037,N_11983);
and U13133 (N_13133,N_10772,N_11364);
xnor U13134 (N_13134,N_10571,N_11909);
xor U13135 (N_13135,N_10431,N_11539);
nor U13136 (N_13136,N_11109,N_10488);
or U13137 (N_13137,N_10914,N_11050);
nor U13138 (N_13138,N_10043,N_10396);
nor U13139 (N_13139,N_11963,N_11510);
nand U13140 (N_13140,N_11891,N_11890);
xnor U13141 (N_13141,N_11286,N_10360);
nand U13142 (N_13142,N_10472,N_10081);
or U13143 (N_13143,N_10110,N_10849);
xnor U13144 (N_13144,N_11505,N_11722);
xnor U13145 (N_13145,N_11795,N_10661);
and U13146 (N_13146,N_11620,N_11621);
or U13147 (N_13147,N_11086,N_11823);
or U13148 (N_13148,N_10175,N_11622);
xor U13149 (N_13149,N_11513,N_11644);
and U13150 (N_13150,N_11874,N_11886);
and U13151 (N_13151,N_10642,N_10969);
xnor U13152 (N_13152,N_10072,N_10860);
nor U13153 (N_13153,N_11712,N_11250);
nand U13154 (N_13154,N_11431,N_10743);
xnor U13155 (N_13155,N_11546,N_10351);
xnor U13156 (N_13156,N_11173,N_11322);
xor U13157 (N_13157,N_10276,N_10290);
xnor U13158 (N_13158,N_11093,N_10346);
nand U13159 (N_13159,N_10690,N_11990);
nor U13160 (N_13160,N_11940,N_10012);
nor U13161 (N_13161,N_11009,N_10267);
nand U13162 (N_13162,N_10287,N_11488);
nor U13163 (N_13163,N_10577,N_11945);
and U13164 (N_13164,N_11782,N_11083);
xor U13165 (N_13165,N_11006,N_10064);
xnor U13166 (N_13166,N_11875,N_10624);
or U13167 (N_13167,N_10078,N_10230);
nor U13168 (N_13168,N_11688,N_11223);
or U13169 (N_13169,N_10365,N_10758);
xor U13170 (N_13170,N_10070,N_11658);
nand U13171 (N_13171,N_11238,N_10005);
nor U13172 (N_13172,N_11631,N_11791);
nand U13173 (N_13173,N_11420,N_10852);
nor U13174 (N_13174,N_11476,N_10242);
xor U13175 (N_13175,N_10034,N_11747);
xnor U13176 (N_13176,N_10409,N_11701);
nor U13177 (N_13177,N_10315,N_11920);
and U13178 (N_13178,N_10171,N_10039);
and U13179 (N_13179,N_11455,N_11719);
xnor U13180 (N_13180,N_10484,N_10957);
and U13181 (N_13181,N_10338,N_10580);
xnor U13182 (N_13182,N_11193,N_11516);
nor U13183 (N_13183,N_11750,N_10259);
xnor U13184 (N_13184,N_10293,N_11527);
nand U13185 (N_13185,N_10576,N_11956);
nor U13186 (N_13186,N_10124,N_10296);
xnor U13187 (N_13187,N_11947,N_11756);
nand U13188 (N_13188,N_10751,N_10236);
or U13189 (N_13189,N_11260,N_10692);
nor U13190 (N_13190,N_10689,N_10455);
nor U13191 (N_13191,N_11622,N_10291);
nand U13192 (N_13192,N_10619,N_10305);
nand U13193 (N_13193,N_11914,N_10545);
nor U13194 (N_13194,N_10919,N_11864);
xor U13195 (N_13195,N_11612,N_10028);
xnor U13196 (N_13196,N_10232,N_11932);
and U13197 (N_13197,N_10236,N_10662);
xnor U13198 (N_13198,N_11292,N_10589);
nor U13199 (N_13199,N_10527,N_10217);
nand U13200 (N_13200,N_10085,N_11131);
nand U13201 (N_13201,N_11350,N_11532);
nand U13202 (N_13202,N_11949,N_11777);
or U13203 (N_13203,N_10737,N_10249);
and U13204 (N_13204,N_11562,N_11714);
nor U13205 (N_13205,N_11509,N_11860);
xnor U13206 (N_13206,N_11953,N_10393);
nand U13207 (N_13207,N_10740,N_10727);
and U13208 (N_13208,N_11040,N_11830);
nand U13209 (N_13209,N_10543,N_10561);
nand U13210 (N_13210,N_11338,N_11830);
or U13211 (N_13211,N_11166,N_10631);
nor U13212 (N_13212,N_11190,N_11420);
xor U13213 (N_13213,N_10441,N_11266);
or U13214 (N_13214,N_10097,N_11256);
or U13215 (N_13215,N_10163,N_11782);
or U13216 (N_13216,N_11975,N_10839);
and U13217 (N_13217,N_10259,N_10028);
and U13218 (N_13218,N_11453,N_10297);
and U13219 (N_13219,N_10634,N_11825);
and U13220 (N_13220,N_10061,N_11097);
and U13221 (N_13221,N_10796,N_10866);
nand U13222 (N_13222,N_11938,N_11770);
or U13223 (N_13223,N_10122,N_10478);
or U13224 (N_13224,N_11490,N_10694);
xnor U13225 (N_13225,N_11396,N_11492);
or U13226 (N_13226,N_10945,N_10288);
or U13227 (N_13227,N_10441,N_10132);
or U13228 (N_13228,N_10732,N_11565);
or U13229 (N_13229,N_11383,N_10459);
xnor U13230 (N_13230,N_11790,N_10412);
nor U13231 (N_13231,N_11348,N_11283);
and U13232 (N_13232,N_10334,N_11461);
or U13233 (N_13233,N_11390,N_11067);
and U13234 (N_13234,N_11541,N_10547);
or U13235 (N_13235,N_11275,N_11113);
nand U13236 (N_13236,N_11458,N_10972);
and U13237 (N_13237,N_11333,N_10638);
and U13238 (N_13238,N_11851,N_10923);
or U13239 (N_13239,N_10232,N_11751);
nor U13240 (N_13240,N_10491,N_10300);
xnor U13241 (N_13241,N_11361,N_11318);
nand U13242 (N_13242,N_10867,N_11596);
nand U13243 (N_13243,N_10798,N_11845);
nand U13244 (N_13244,N_11897,N_11564);
xnor U13245 (N_13245,N_10995,N_10006);
or U13246 (N_13246,N_10021,N_11882);
and U13247 (N_13247,N_11240,N_10963);
nor U13248 (N_13248,N_11371,N_10962);
and U13249 (N_13249,N_11022,N_11412);
nor U13250 (N_13250,N_10379,N_11284);
and U13251 (N_13251,N_11788,N_10311);
and U13252 (N_13252,N_11623,N_10623);
xor U13253 (N_13253,N_10783,N_11380);
or U13254 (N_13254,N_10390,N_11164);
or U13255 (N_13255,N_11848,N_11470);
or U13256 (N_13256,N_11985,N_10763);
and U13257 (N_13257,N_11024,N_10854);
and U13258 (N_13258,N_11419,N_11305);
or U13259 (N_13259,N_11512,N_11557);
or U13260 (N_13260,N_10287,N_10409);
nand U13261 (N_13261,N_11702,N_11535);
or U13262 (N_13262,N_10258,N_10349);
xor U13263 (N_13263,N_11570,N_10651);
nor U13264 (N_13264,N_10338,N_11017);
nor U13265 (N_13265,N_10259,N_11653);
and U13266 (N_13266,N_10401,N_11322);
or U13267 (N_13267,N_11348,N_11204);
and U13268 (N_13268,N_11495,N_11570);
or U13269 (N_13269,N_11628,N_11490);
or U13270 (N_13270,N_10594,N_11595);
and U13271 (N_13271,N_11310,N_10933);
nand U13272 (N_13272,N_11807,N_11349);
nor U13273 (N_13273,N_11745,N_10798);
or U13274 (N_13274,N_10748,N_11462);
or U13275 (N_13275,N_10569,N_10330);
nor U13276 (N_13276,N_10321,N_10285);
nor U13277 (N_13277,N_11166,N_10409);
nor U13278 (N_13278,N_11530,N_11471);
or U13279 (N_13279,N_10071,N_11110);
nor U13280 (N_13280,N_10161,N_10056);
or U13281 (N_13281,N_10940,N_11527);
nor U13282 (N_13282,N_10343,N_10417);
xor U13283 (N_13283,N_11327,N_11261);
and U13284 (N_13284,N_10405,N_10719);
nor U13285 (N_13285,N_10861,N_11982);
and U13286 (N_13286,N_11920,N_10173);
or U13287 (N_13287,N_11090,N_11704);
and U13288 (N_13288,N_11083,N_10418);
and U13289 (N_13289,N_11121,N_11458);
or U13290 (N_13290,N_11769,N_11587);
xnor U13291 (N_13291,N_11287,N_10249);
or U13292 (N_13292,N_11463,N_10840);
or U13293 (N_13293,N_11748,N_11783);
nor U13294 (N_13294,N_10049,N_10496);
or U13295 (N_13295,N_11332,N_11203);
and U13296 (N_13296,N_10796,N_11569);
nand U13297 (N_13297,N_10748,N_11355);
nor U13298 (N_13298,N_10063,N_10446);
nor U13299 (N_13299,N_11337,N_10776);
nor U13300 (N_13300,N_11990,N_11201);
nand U13301 (N_13301,N_11672,N_10322);
or U13302 (N_13302,N_10270,N_11044);
xnor U13303 (N_13303,N_10501,N_10521);
nor U13304 (N_13304,N_11550,N_11216);
and U13305 (N_13305,N_11347,N_10340);
xor U13306 (N_13306,N_10342,N_10215);
xor U13307 (N_13307,N_11011,N_11911);
xnor U13308 (N_13308,N_10418,N_11943);
xnor U13309 (N_13309,N_10078,N_11872);
and U13310 (N_13310,N_11170,N_10716);
or U13311 (N_13311,N_10417,N_10441);
and U13312 (N_13312,N_11729,N_11151);
nand U13313 (N_13313,N_10087,N_10412);
and U13314 (N_13314,N_10548,N_11512);
xnor U13315 (N_13315,N_11001,N_10593);
or U13316 (N_13316,N_10609,N_10071);
or U13317 (N_13317,N_10055,N_10609);
nor U13318 (N_13318,N_11656,N_11187);
and U13319 (N_13319,N_10966,N_10463);
nand U13320 (N_13320,N_11872,N_10265);
nor U13321 (N_13321,N_11928,N_11735);
and U13322 (N_13322,N_11924,N_11775);
xor U13323 (N_13323,N_11952,N_10266);
xor U13324 (N_13324,N_10044,N_11573);
and U13325 (N_13325,N_11284,N_10827);
and U13326 (N_13326,N_11444,N_11584);
or U13327 (N_13327,N_11458,N_11939);
xnor U13328 (N_13328,N_10985,N_10858);
nor U13329 (N_13329,N_11429,N_10370);
or U13330 (N_13330,N_10757,N_10040);
or U13331 (N_13331,N_10018,N_11308);
or U13332 (N_13332,N_11498,N_10514);
and U13333 (N_13333,N_11079,N_11633);
and U13334 (N_13334,N_10347,N_10449);
and U13335 (N_13335,N_10944,N_10291);
xnor U13336 (N_13336,N_10195,N_10377);
or U13337 (N_13337,N_11954,N_11939);
xnor U13338 (N_13338,N_10408,N_11637);
or U13339 (N_13339,N_10657,N_10875);
xor U13340 (N_13340,N_10788,N_10166);
or U13341 (N_13341,N_11694,N_11373);
and U13342 (N_13342,N_11298,N_11009);
and U13343 (N_13343,N_11085,N_11696);
nor U13344 (N_13344,N_11316,N_10972);
nor U13345 (N_13345,N_11024,N_11787);
or U13346 (N_13346,N_10226,N_10798);
or U13347 (N_13347,N_10547,N_10612);
nor U13348 (N_13348,N_10985,N_10114);
and U13349 (N_13349,N_10222,N_11454);
or U13350 (N_13350,N_11659,N_11375);
nand U13351 (N_13351,N_10926,N_10302);
nor U13352 (N_13352,N_10966,N_11626);
or U13353 (N_13353,N_10640,N_11749);
or U13354 (N_13354,N_10746,N_10416);
and U13355 (N_13355,N_10461,N_10255);
nor U13356 (N_13356,N_10678,N_11249);
nand U13357 (N_13357,N_10600,N_10790);
and U13358 (N_13358,N_11048,N_11195);
nand U13359 (N_13359,N_11302,N_10518);
and U13360 (N_13360,N_10310,N_10458);
and U13361 (N_13361,N_11762,N_10749);
or U13362 (N_13362,N_11651,N_11210);
or U13363 (N_13363,N_11347,N_11718);
and U13364 (N_13364,N_10475,N_10783);
xor U13365 (N_13365,N_11375,N_11243);
nand U13366 (N_13366,N_10484,N_10830);
xor U13367 (N_13367,N_11324,N_11792);
or U13368 (N_13368,N_10291,N_11699);
and U13369 (N_13369,N_11142,N_11459);
or U13370 (N_13370,N_10626,N_10553);
or U13371 (N_13371,N_11019,N_11004);
xor U13372 (N_13372,N_11704,N_11725);
xor U13373 (N_13373,N_10432,N_10476);
nor U13374 (N_13374,N_10873,N_11321);
or U13375 (N_13375,N_11226,N_10622);
nor U13376 (N_13376,N_10019,N_10269);
and U13377 (N_13377,N_10085,N_11329);
nor U13378 (N_13378,N_10480,N_10801);
nor U13379 (N_13379,N_11065,N_10692);
nor U13380 (N_13380,N_11498,N_10931);
nand U13381 (N_13381,N_11232,N_11172);
nand U13382 (N_13382,N_10873,N_11222);
or U13383 (N_13383,N_11760,N_11322);
nor U13384 (N_13384,N_11621,N_11177);
and U13385 (N_13385,N_11057,N_10771);
nand U13386 (N_13386,N_11580,N_10298);
xor U13387 (N_13387,N_11918,N_10499);
nor U13388 (N_13388,N_10725,N_11576);
xnor U13389 (N_13389,N_11850,N_10143);
nand U13390 (N_13390,N_10486,N_11419);
nor U13391 (N_13391,N_10838,N_10996);
nand U13392 (N_13392,N_11736,N_11529);
or U13393 (N_13393,N_10465,N_10755);
xor U13394 (N_13394,N_10808,N_11059);
xnor U13395 (N_13395,N_11648,N_11848);
or U13396 (N_13396,N_11298,N_11171);
nor U13397 (N_13397,N_10746,N_11876);
nand U13398 (N_13398,N_10310,N_10740);
nand U13399 (N_13399,N_11122,N_10122);
nand U13400 (N_13400,N_11943,N_10571);
xnor U13401 (N_13401,N_10460,N_11841);
xnor U13402 (N_13402,N_11140,N_11398);
nor U13403 (N_13403,N_10287,N_11997);
or U13404 (N_13404,N_11772,N_10686);
xor U13405 (N_13405,N_11076,N_11077);
nor U13406 (N_13406,N_10135,N_11337);
and U13407 (N_13407,N_10849,N_10163);
xor U13408 (N_13408,N_11233,N_10968);
xnor U13409 (N_13409,N_11844,N_10065);
xor U13410 (N_13410,N_11973,N_10290);
nor U13411 (N_13411,N_11679,N_10714);
nand U13412 (N_13412,N_10866,N_11145);
nand U13413 (N_13413,N_11987,N_11794);
xnor U13414 (N_13414,N_11532,N_10108);
and U13415 (N_13415,N_10988,N_10586);
or U13416 (N_13416,N_11940,N_11814);
or U13417 (N_13417,N_11300,N_10264);
nor U13418 (N_13418,N_10086,N_10726);
or U13419 (N_13419,N_11678,N_11528);
xnor U13420 (N_13420,N_11803,N_11245);
xor U13421 (N_13421,N_10525,N_10977);
and U13422 (N_13422,N_10056,N_11616);
and U13423 (N_13423,N_10784,N_11816);
xnor U13424 (N_13424,N_11581,N_10468);
xnor U13425 (N_13425,N_10587,N_10139);
xor U13426 (N_13426,N_11246,N_11955);
nor U13427 (N_13427,N_10198,N_11308);
nand U13428 (N_13428,N_11169,N_10074);
nor U13429 (N_13429,N_10053,N_10230);
xor U13430 (N_13430,N_10819,N_10933);
xor U13431 (N_13431,N_10470,N_10852);
xor U13432 (N_13432,N_10765,N_11399);
nor U13433 (N_13433,N_11387,N_11098);
and U13434 (N_13434,N_10924,N_11118);
or U13435 (N_13435,N_11730,N_10927);
and U13436 (N_13436,N_10610,N_11746);
nand U13437 (N_13437,N_11566,N_10484);
nor U13438 (N_13438,N_10989,N_10243);
xor U13439 (N_13439,N_10997,N_11705);
nor U13440 (N_13440,N_10708,N_10460);
xnor U13441 (N_13441,N_10845,N_10332);
nand U13442 (N_13442,N_11134,N_11565);
nor U13443 (N_13443,N_10750,N_10226);
and U13444 (N_13444,N_10664,N_10843);
or U13445 (N_13445,N_10680,N_10274);
nand U13446 (N_13446,N_11606,N_10281);
nor U13447 (N_13447,N_10610,N_10312);
and U13448 (N_13448,N_11126,N_10981);
nor U13449 (N_13449,N_10014,N_11357);
and U13450 (N_13450,N_10989,N_11418);
or U13451 (N_13451,N_10281,N_11330);
or U13452 (N_13452,N_10751,N_11917);
nand U13453 (N_13453,N_10962,N_10134);
nor U13454 (N_13454,N_10238,N_10233);
or U13455 (N_13455,N_11430,N_11980);
or U13456 (N_13456,N_11709,N_10506);
xor U13457 (N_13457,N_11293,N_10310);
xor U13458 (N_13458,N_10754,N_11585);
or U13459 (N_13459,N_11282,N_10254);
and U13460 (N_13460,N_11690,N_10490);
xnor U13461 (N_13461,N_10870,N_10507);
or U13462 (N_13462,N_11961,N_11555);
nand U13463 (N_13463,N_10003,N_11777);
and U13464 (N_13464,N_11659,N_10410);
or U13465 (N_13465,N_11453,N_11846);
or U13466 (N_13466,N_10019,N_11188);
xor U13467 (N_13467,N_10297,N_11967);
nand U13468 (N_13468,N_10945,N_10809);
nor U13469 (N_13469,N_11579,N_11427);
xnor U13470 (N_13470,N_10561,N_10885);
or U13471 (N_13471,N_10008,N_10900);
xor U13472 (N_13472,N_10683,N_10118);
and U13473 (N_13473,N_10530,N_11290);
nand U13474 (N_13474,N_10320,N_11975);
xor U13475 (N_13475,N_11800,N_11120);
nor U13476 (N_13476,N_11669,N_10208);
nand U13477 (N_13477,N_11540,N_10658);
nand U13478 (N_13478,N_10591,N_10975);
nand U13479 (N_13479,N_11616,N_10154);
or U13480 (N_13480,N_11315,N_11559);
xnor U13481 (N_13481,N_11504,N_10607);
and U13482 (N_13482,N_10622,N_10324);
nand U13483 (N_13483,N_10200,N_10156);
or U13484 (N_13484,N_11691,N_10744);
xor U13485 (N_13485,N_10027,N_11806);
nor U13486 (N_13486,N_10582,N_11243);
nand U13487 (N_13487,N_11007,N_11475);
or U13488 (N_13488,N_11020,N_11723);
xnor U13489 (N_13489,N_11718,N_10994);
xor U13490 (N_13490,N_11127,N_11274);
and U13491 (N_13491,N_11234,N_11491);
or U13492 (N_13492,N_10080,N_11263);
nor U13493 (N_13493,N_11229,N_11730);
nor U13494 (N_13494,N_10846,N_11987);
xor U13495 (N_13495,N_11219,N_10307);
nor U13496 (N_13496,N_11514,N_11978);
or U13497 (N_13497,N_10460,N_11520);
nand U13498 (N_13498,N_11344,N_10562);
nand U13499 (N_13499,N_10378,N_11995);
xor U13500 (N_13500,N_11810,N_10171);
and U13501 (N_13501,N_11835,N_11148);
xor U13502 (N_13502,N_10476,N_10037);
nand U13503 (N_13503,N_10003,N_10019);
nand U13504 (N_13504,N_11945,N_10213);
and U13505 (N_13505,N_10662,N_10637);
nand U13506 (N_13506,N_10656,N_10018);
or U13507 (N_13507,N_10897,N_10733);
nand U13508 (N_13508,N_11437,N_11594);
or U13509 (N_13509,N_10130,N_11682);
and U13510 (N_13510,N_11983,N_11334);
nor U13511 (N_13511,N_10862,N_10176);
nor U13512 (N_13512,N_11371,N_10817);
nand U13513 (N_13513,N_11571,N_10328);
nor U13514 (N_13514,N_11594,N_11775);
xnor U13515 (N_13515,N_11480,N_10503);
xor U13516 (N_13516,N_11786,N_11920);
xnor U13517 (N_13517,N_10677,N_10541);
xnor U13518 (N_13518,N_11973,N_11926);
nor U13519 (N_13519,N_11298,N_10912);
and U13520 (N_13520,N_11287,N_10667);
xnor U13521 (N_13521,N_11036,N_10784);
and U13522 (N_13522,N_11519,N_11975);
and U13523 (N_13523,N_10292,N_11818);
nand U13524 (N_13524,N_10647,N_11303);
nor U13525 (N_13525,N_11329,N_11183);
and U13526 (N_13526,N_11814,N_11646);
nor U13527 (N_13527,N_11662,N_11784);
and U13528 (N_13528,N_11917,N_10917);
nand U13529 (N_13529,N_10548,N_10202);
nor U13530 (N_13530,N_10311,N_11895);
or U13531 (N_13531,N_10297,N_10321);
nor U13532 (N_13532,N_10741,N_10507);
nand U13533 (N_13533,N_11043,N_11689);
and U13534 (N_13534,N_10590,N_10002);
nand U13535 (N_13535,N_10090,N_10820);
and U13536 (N_13536,N_10923,N_11859);
xor U13537 (N_13537,N_10722,N_11772);
nor U13538 (N_13538,N_11637,N_10832);
xnor U13539 (N_13539,N_10860,N_10378);
xor U13540 (N_13540,N_11460,N_10819);
xnor U13541 (N_13541,N_10015,N_11583);
xor U13542 (N_13542,N_11808,N_10775);
nand U13543 (N_13543,N_11515,N_11516);
xor U13544 (N_13544,N_11272,N_10831);
nand U13545 (N_13545,N_10958,N_11438);
or U13546 (N_13546,N_11266,N_10674);
nand U13547 (N_13547,N_10673,N_10026);
xor U13548 (N_13548,N_10906,N_11818);
and U13549 (N_13549,N_10365,N_10770);
nor U13550 (N_13550,N_10629,N_11639);
and U13551 (N_13551,N_11538,N_11507);
nand U13552 (N_13552,N_11743,N_11793);
and U13553 (N_13553,N_11042,N_11959);
nand U13554 (N_13554,N_10472,N_11775);
or U13555 (N_13555,N_10885,N_11675);
and U13556 (N_13556,N_11891,N_11323);
nand U13557 (N_13557,N_10170,N_10790);
nor U13558 (N_13558,N_10762,N_11675);
nor U13559 (N_13559,N_11444,N_11730);
and U13560 (N_13560,N_11317,N_11768);
and U13561 (N_13561,N_11207,N_11777);
nand U13562 (N_13562,N_10232,N_11217);
nand U13563 (N_13563,N_10115,N_10008);
or U13564 (N_13564,N_10053,N_10429);
and U13565 (N_13565,N_11026,N_11504);
nor U13566 (N_13566,N_10590,N_11016);
nand U13567 (N_13567,N_11606,N_10940);
xnor U13568 (N_13568,N_11940,N_11427);
xnor U13569 (N_13569,N_11483,N_10623);
nand U13570 (N_13570,N_10614,N_11402);
xnor U13571 (N_13571,N_10254,N_10941);
and U13572 (N_13572,N_10370,N_10248);
or U13573 (N_13573,N_11670,N_10207);
nor U13574 (N_13574,N_10112,N_11248);
xor U13575 (N_13575,N_11568,N_11630);
nand U13576 (N_13576,N_11424,N_10869);
nand U13577 (N_13577,N_11441,N_10369);
nor U13578 (N_13578,N_10896,N_11542);
nand U13579 (N_13579,N_11257,N_10629);
and U13580 (N_13580,N_10273,N_11755);
and U13581 (N_13581,N_10140,N_11871);
xor U13582 (N_13582,N_10570,N_10514);
xnor U13583 (N_13583,N_10322,N_10813);
nor U13584 (N_13584,N_10370,N_11056);
nand U13585 (N_13585,N_10166,N_11709);
nand U13586 (N_13586,N_11850,N_11633);
nor U13587 (N_13587,N_11500,N_11184);
or U13588 (N_13588,N_11568,N_11523);
nand U13589 (N_13589,N_10477,N_11440);
or U13590 (N_13590,N_10759,N_10605);
and U13591 (N_13591,N_10108,N_11950);
nand U13592 (N_13592,N_10484,N_10795);
or U13593 (N_13593,N_10022,N_11597);
nand U13594 (N_13594,N_10898,N_10746);
nand U13595 (N_13595,N_11105,N_10195);
nor U13596 (N_13596,N_11782,N_10791);
or U13597 (N_13597,N_10478,N_11488);
xor U13598 (N_13598,N_10384,N_10204);
nand U13599 (N_13599,N_10178,N_11555);
nor U13600 (N_13600,N_11813,N_10569);
nor U13601 (N_13601,N_10136,N_10091);
or U13602 (N_13602,N_10432,N_11540);
xor U13603 (N_13603,N_10161,N_10846);
nor U13604 (N_13604,N_11802,N_11864);
nor U13605 (N_13605,N_10882,N_11325);
nor U13606 (N_13606,N_11148,N_10770);
nor U13607 (N_13607,N_11312,N_11481);
nor U13608 (N_13608,N_10726,N_11562);
xor U13609 (N_13609,N_11355,N_10131);
nor U13610 (N_13610,N_10069,N_11215);
and U13611 (N_13611,N_11046,N_11641);
xor U13612 (N_13612,N_11653,N_11991);
xor U13613 (N_13613,N_11554,N_11795);
nor U13614 (N_13614,N_10207,N_10795);
nor U13615 (N_13615,N_10854,N_11718);
nor U13616 (N_13616,N_11078,N_11741);
or U13617 (N_13617,N_10963,N_11998);
nor U13618 (N_13618,N_11138,N_10049);
nand U13619 (N_13619,N_11014,N_11280);
xnor U13620 (N_13620,N_10581,N_11123);
xnor U13621 (N_13621,N_10926,N_11569);
nand U13622 (N_13622,N_11435,N_10817);
nand U13623 (N_13623,N_11217,N_11003);
or U13624 (N_13624,N_10249,N_10595);
nand U13625 (N_13625,N_10403,N_11793);
or U13626 (N_13626,N_10287,N_10738);
nand U13627 (N_13627,N_11865,N_11966);
and U13628 (N_13628,N_10163,N_10315);
nor U13629 (N_13629,N_10039,N_11171);
nand U13630 (N_13630,N_11074,N_11451);
nor U13631 (N_13631,N_10168,N_11819);
nand U13632 (N_13632,N_11764,N_10448);
or U13633 (N_13633,N_11242,N_10766);
and U13634 (N_13634,N_11759,N_10586);
nand U13635 (N_13635,N_10066,N_11800);
nor U13636 (N_13636,N_11606,N_10984);
or U13637 (N_13637,N_10437,N_11489);
or U13638 (N_13638,N_10663,N_10274);
nor U13639 (N_13639,N_10967,N_11635);
and U13640 (N_13640,N_10099,N_11715);
and U13641 (N_13641,N_10657,N_10493);
or U13642 (N_13642,N_10097,N_10533);
xor U13643 (N_13643,N_10789,N_11775);
xor U13644 (N_13644,N_10033,N_11071);
xnor U13645 (N_13645,N_11741,N_10915);
nand U13646 (N_13646,N_11862,N_11317);
xor U13647 (N_13647,N_11366,N_11004);
and U13648 (N_13648,N_10835,N_10201);
nand U13649 (N_13649,N_11414,N_10693);
xnor U13650 (N_13650,N_10475,N_11632);
and U13651 (N_13651,N_11595,N_11883);
xnor U13652 (N_13652,N_10155,N_10446);
and U13653 (N_13653,N_11848,N_10137);
nor U13654 (N_13654,N_10084,N_11276);
or U13655 (N_13655,N_10091,N_11128);
or U13656 (N_13656,N_11528,N_11507);
nor U13657 (N_13657,N_10703,N_11142);
or U13658 (N_13658,N_10528,N_11727);
and U13659 (N_13659,N_11451,N_10925);
and U13660 (N_13660,N_10517,N_11588);
xor U13661 (N_13661,N_10971,N_11250);
nand U13662 (N_13662,N_11447,N_11239);
nor U13663 (N_13663,N_11203,N_11312);
nand U13664 (N_13664,N_11678,N_11981);
xor U13665 (N_13665,N_10402,N_10221);
or U13666 (N_13666,N_10649,N_10081);
nand U13667 (N_13667,N_11308,N_10349);
and U13668 (N_13668,N_11700,N_11229);
and U13669 (N_13669,N_10528,N_11916);
nor U13670 (N_13670,N_11315,N_10724);
and U13671 (N_13671,N_11562,N_11326);
and U13672 (N_13672,N_10367,N_10637);
nor U13673 (N_13673,N_10734,N_10091);
nand U13674 (N_13674,N_10899,N_11937);
or U13675 (N_13675,N_10138,N_11091);
nor U13676 (N_13676,N_10842,N_10816);
or U13677 (N_13677,N_10908,N_10867);
and U13678 (N_13678,N_10710,N_11377);
and U13679 (N_13679,N_11314,N_10338);
and U13680 (N_13680,N_10358,N_10501);
nand U13681 (N_13681,N_11965,N_10457);
nor U13682 (N_13682,N_11976,N_11472);
nand U13683 (N_13683,N_11243,N_10623);
and U13684 (N_13684,N_10426,N_10711);
nor U13685 (N_13685,N_11375,N_10089);
or U13686 (N_13686,N_11224,N_10649);
and U13687 (N_13687,N_11680,N_10609);
nor U13688 (N_13688,N_11154,N_10128);
nand U13689 (N_13689,N_10382,N_10077);
nand U13690 (N_13690,N_11328,N_11525);
xor U13691 (N_13691,N_11964,N_10159);
and U13692 (N_13692,N_10865,N_11026);
nor U13693 (N_13693,N_10201,N_10351);
and U13694 (N_13694,N_10034,N_11068);
nand U13695 (N_13695,N_10773,N_11607);
nand U13696 (N_13696,N_11359,N_10139);
nor U13697 (N_13697,N_10459,N_10453);
or U13698 (N_13698,N_11781,N_11175);
or U13699 (N_13699,N_10956,N_10988);
xnor U13700 (N_13700,N_10915,N_11069);
nor U13701 (N_13701,N_10235,N_10945);
nand U13702 (N_13702,N_11756,N_11786);
nor U13703 (N_13703,N_11008,N_10180);
and U13704 (N_13704,N_11037,N_10968);
nand U13705 (N_13705,N_11885,N_11264);
nand U13706 (N_13706,N_10615,N_11351);
nand U13707 (N_13707,N_10301,N_11982);
xor U13708 (N_13708,N_10054,N_10503);
nand U13709 (N_13709,N_10607,N_10327);
xor U13710 (N_13710,N_11303,N_10883);
or U13711 (N_13711,N_10053,N_11154);
nand U13712 (N_13712,N_10024,N_11455);
nor U13713 (N_13713,N_10724,N_10443);
nand U13714 (N_13714,N_11433,N_10009);
or U13715 (N_13715,N_11099,N_10433);
or U13716 (N_13716,N_11952,N_10563);
xor U13717 (N_13717,N_11843,N_10513);
nand U13718 (N_13718,N_11432,N_11217);
and U13719 (N_13719,N_10543,N_11361);
or U13720 (N_13720,N_10483,N_10320);
xnor U13721 (N_13721,N_10706,N_11178);
and U13722 (N_13722,N_11964,N_11362);
nand U13723 (N_13723,N_10768,N_11752);
nor U13724 (N_13724,N_10412,N_11853);
and U13725 (N_13725,N_11531,N_10515);
or U13726 (N_13726,N_11766,N_11654);
nand U13727 (N_13727,N_11380,N_11754);
nand U13728 (N_13728,N_10518,N_11139);
nand U13729 (N_13729,N_10370,N_10143);
nor U13730 (N_13730,N_10115,N_11157);
or U13731 (N_13731,N_10860,N_10068);
nand U13732 (N_13732,N_11128,N_10070);
nor U13733 (N_13733,N_11692,N_10616);
xor U13734 (N_13734,N_11150,N_11981);
xnor U13735 (N_13735,N_10042,N_11070);
nor U13736 (N_13736,N_11324,N_10766);
or U13737 (N_13737,N_11658,N_11730);
nor U13738 (N_13738,N_10496,N_11959);
and U13739 (N_13739,N_11937,N_10269);
and U13740 (N_13740,N_11948,N_11843);
xor U13741 (N_13741,N_11277,N_10785);
nand U13742 (N_13742,N_10930,N_10468);
nor U13743 (N_13743,N_11711,N_10373);
xor U13744 (N_13744,N_10470,N_11608);
xnor U13745 (N_13745,N_10334,N_11639);
xnor U13746 (N_13746,N_11545,N_11699);
xnor U13747 (N_13747,N_11469,N_11309);
or U13748 (N_13748,N_10624,N_11894);
nor U13749 (N_13749,N_10818,N_10891);
nor U13750 (N_13750,N_10426,N_10667);
and U13751 (N_13751,N_11232,N_10188);
or U13752 (N_13752,N_10662,N_11826);
nor U13753 (N_13753,N_10648,N_11260);
xnor U13754 (N_13754,N_11520,N_10904);
or U13755 (N_13755,N_10150,N_11858);
or U13756 (N_13756,N_10932,N_11130);
or U13757 (N_13757,N_11675,N_10063);
xor U13758 (N_13758,N_10114,N_11327);
and U13759 (N_13759,N_11677,N_10442);
nor U13760 (N_13760,N_11578,N_11296);
nor U13761 (N_13761,N_10942,N_11583);
or U13762 (N_13762,N_11180,N_11117);
nand U13763 (N_13763,N_11449,N_10479);
xor U13764 (N_13764,N_10282,N_11324);
xor U13765 (N_13765,N_10759,N_10308);
and U13766 (N_13766,N_11305,N_11441);
nor U13767 (N_13767,N_11176,N_11743);
nand U13768 (N_13768,N_11827,N_11377);
and U13769 (N_13769,N_10585,N_10905);
nor U13770 (N_13770,N_11296,N_10638);
nor U13771 (N_13771,N_10261,N_11082);
nor U13772 (N_13772,N_11297,N_10325);
or U13773 (N_13773,N_11785,N_11752);
or U13774 (N_13774,N_11725,N_10326);
and U13775 (N_13775,N_11993,N_11072);
and U13776 (N_13776,N_10837,N_11927);
and U13777 (N_13777,N_10279,N_10724);
and U13778 (N_13778,N_11813,N_10534);
nor U13779 (N_13779,N_10040,N_10428);
or U13780 (N_13780,N_10569,N_10228);
and U13781 (N_13781,N_10744,N_11788);
xnor U13782 (N_13782,N_10628,N_11053);
xor U13783 (N_13783,N_10763,N_11750);
nor U13784 (N_13784,N_11532,N_10287);
nand U13785 (N_13785,N_10097,N_11072);
xor U13786 (N_13786,N_11847,N_11625);
nand U13787 (N_13787,N_10115,N_10233);
or U13788 (N_13788,N_10604,N_11928);
nand U13789 (N_13789,N_10745,N_11929);
and U13790 (N_13790,N_10588,N_11683);
and U13791 (N_13791,N_11893,N_11674);
and U13792 (N_13792,N_11282,N_10757);
nor U13793 (N_13793,N_10129,N_10468);
or U13794 (N_13794,N_10239,N_10575);
nand U13795 (N_13795,N_11281,N_11934);
nor U13796 (N_13796,N_11218,N_11585);
nor U13797 (N_13797,N_11731,N_11873);
or U13798 (N_13798,N_10747,N_10218);
and U13799 (N_13799,N_11918,N_11667);
nand U13800 (N_13800,N_11350,N_10678);
and U13801 (N_13801,N_11077,N_10468);
xnor U13802 (N_13802,N_10652,N_11484);
nor U13803 (N_13803,N_10137,N_10170);
nand U13804 (N_13804,N_11668,N_11163);
and U13805 (N_13805,N_11522,N_10757);
and U13806 (N_13806,N_11780,N_10029);
nor U13807 (N_13807,N_11846,N_10995);
xnor U13808 (N_13808,N_10042,N_11366);
or U13809 (N_13809,N_10995,N_10693);
xor U13810 (N_13810,N_11037,N_10960);
xnor U13811 (N_13811,N_10202,N_11288);
and U13812 (N_13812,N_10821,N_11744);
xnor U13813 (N_13813,N_10626,N_11252);
nand U13814 (N_13814,N_11129,N_11975);
xnor U13815 (N_13815,N_10033,N_11333);
and U13816 (N_13816,N_11677,N_11912);
xor U13817 (N_13817,N_10198,N_11980);
nor U13818 (N_13818,N_10237,N_10702);
xor U13819 (N_13819,N_10079,N_11005);
and U13820 (N_13820,N_11747,N_11446);
xor U13821 (N_13821,N_11640,N_10278);
nor U13822 (N_13822,N_11564,N_11221);
xnor U13823 (N_13823,N_11996,N_10559);
and U13824 (N_13824,N_10070,N_10090);
nor U13825 (N_13825,N_11030,N_11782);
and U13826 (N_13826,N_11323,N_10132);
nor U13827 (N_13827,N_11261,N_10697);
xnor U13828 (N_13828,N_10728,N_10542);
and U13829 (N_13829,N_10360,N_11696);
xor U13830 (N_13830,N_10814,N_11026);
nand U13831 (N_13831,N_11754,N_11081);
or U13832 (N_13832,N_11729,N_11047);
and U13833 (N_13833,N_11854,N_11537);
xnor U13834 (N_13834,N_11679,N_11783);
nor U13835 (N_13835,N_10323,N_11807);
nand U13836 (N_13836,N_10298,N_10609);
nor U13837 (N_13837,N_11472,N_11563);
nand U13838 (N_13838,N_10961,N_11327);
and U13839 (N_13839,N_10783,N_11628);
nor U13840 (N_13840,N_10548,N_11708);
and U13841 (N_13841,N_11526,N_10736);
or U13842 (N_13842,N_10980,N_10985);
or U13843 (N_13843,N_11972,N_11542);
xor U13844 (N_13844,N_11922,N_10040);
xor U13845 (N_13845,N_10161,N_11586);
or U13846 (N_13846,N_11614,N_10550);
nor U13847 (N_13847,N_11177,N_10106);
nand U13848 (N_13848,N_11657,N_11155);
nand U13849 (N_13849,N_10232,N_11875);
nor U13850 (N_13850,N_10447,N_10151);
nand U13851 (N_13851,N_10638,N_10570);
or U13852 (N_13852,N_10933,N_10382);
and U13853 (N_13853,N_11298,N_11566);
nor U13854 (N_13854,N_10208,N_10101);
xnor U13855 (N_13855,N_10533,N_10009);
xnor U13856 (N_13856,N_11390,N_11600);
or U13857 (N_13857,N_10315,N_11915);
or U13858 (N_13858,N_11539,N_11347);
and U13859 (N_13859,N_10519,N_11235);
and U13860 (N_13860,N_11347,N_10642);
xnor U13861 (N_13861,N_11435,N_10146);
or U13862 (N_13862,N_10055,N_11331);
xnor U13863 (N_13863,N_11437,N_11843);
or U13864 (N_13864,N_11144,N_10235);
or U13865 (N_13865,N_11203,N_11806);
nor U13866 (N_13866,N_10606,N_11882);
and U13867 (N_13867,N_11411,N_11798);
nand U13868 (N_13868,N_11866,N_10108);
or U13869 (N_13869,N_10785,N_10453);
and U13870 (N_13870,N_11566,N_11386);
nor U13871 (N_13871,N_10426,N_11380);
or U13872 (N_13872,N_11028,N_10810);
nor U13873 (N_13873,N_11264,N_11194);
nor U13874 (N_13874,N_10104,N_10494);
xnor U13875 (N_13875,N_11284,N_11145);
or U13876 (N_13876,N_11632,N_10894);
xor U13877 (N_13877,N_10812,N_11961);
xnor U13878 (N_13878,N_11540,N_10534);
nand U13879 (N_13879,N_10409,N_11153);
and U13880 (N_13880,N_10236,N_11997);
and U13881 (N_13881,N_11506,N_10822);
xnor U13882 (N_13882,N_11553,N_10202);
nand U13883 (N_13883,N_10489,N_10304);
nand U13884 (N_13884,N_10030,N_10719);
nand U13885 (N_13885,N_10943,N_11539);
and U13886 (N_13886,N_11801,N_10461);
and U13887 (N_13887,N_11554,N_10513);
and U13888 (N_13888,N_11728,N_11802);
nand U13889 (N_13889,N_11235,N_10295);
and U13890 (N_13890,N_10065,N_10405);
and U13891 (N_13891,N_11525,N_11533);
xnor U13892 (N_13892,N_11212,N_11102);
nand U13893 (N_13893,N_10428,N_11245);
nor U13894 (N_13894,N_11075,N_10301);
xnor U13895 (N_13895,N_11013,N_11736);
nand U13896 (N_13896,N_11946,N_11818);
xnor U13897 (N_13897,N_10681,N_10063);
nor U13898 (N_13898,N_11344,N_11479);
nand U13899 (N_13899,N_11528,N_11837);
xor U13900 (N_13900,N_10570,N_11172);
and U13901 (N_13901,N_11423,N_11225);
nor U13902 (N_13902,N_11832,N_10163);
nand U13903 (N_13903,N_11901,N_10505);
xor U13904 (N_13904,N_10814,N_10542);
nor U13905 (N_13905,N_11781,N_11182);
nand U13906 (N_13906,N_11946,N_11325);
and U13907 (N_13907,N_10794,N_11328);
or U13908 (N_13908,N_10585,N_10927);
and U13909 (N_13909,N_10750,N_10471);
xnor U13910 (N_13910,N_10221,N_10330);
or U13911 (N_13911,N_11649,N_10089);
nand U13912 (N_13912,N_10924,N_10356);
nor U13913 (N_13913,N_11252,N_10255);
or U13914 (N_13914,N_11058,N_10366);
or U13915 (N_13915,N_11955,N_11182);
and U13916 (N_13916,N_10187,N_10140);
and U13917 (N_13917,N_11894,N_10638);
xnor U13918 (N_13918,N_11704,N_11141);
nor U13919 (N_13919,N_11820,N_11971);
or U13920 (N_13920,N_11458,N_11783);
and U13921 (N_13921,N_10047,N_11753);
nand U13922 (N_13922,N_11352,N_10910);
nor U13923 (N_13923,N_11961,N_10950);
nor U13924 (N_13924,N_11070,N_10457);
nand U13925 (N_13925,N_11816,N_11248);
xnor U13926 (N_13926,N_10467,N_10527);
or U13927 (N_13927,N_11592,N_11944);
or U13928 (N_13928,N_11281,N_10307);
nor U13929 (N_13929,N_11064,N_11877);
and U13930 (N_13930,N_10439,N_10973);
and U13931 (N_13931,N_10453,N_11866);
or U13932 (N_13932,N_10760,N_10127);
or U13933 (N_13933,N_10609,N_11876);
nor U13934 (N_13934,N_10232,N_10945);
nand U13935 (N_13935,N_10124,N_11728);
and U13936 (N_13936,N_11026,N_11128);
xnor U13937 (N_13937,N_11035,N_11378);
xor U13938 (N_13938,N_11532,N_10581);
or U13939 (N_13939,N_10396,N_10648);
xor U13940 (N_13940,N_10813,N_11311);
nor U13941 (N_13941,N_10356,N_11887);
nor U13942 (N_13942,N_11816,N_11881);
xnor U13943 (N_13943,N_11783,N_11002);
or U13944 (N_13944,N_11342,N_11134);
or U13945 (N_13945,N_11678,N_11780);
xnor U13946 (N_13946,N_10739,N_10307);
xor U13947 (N_13947,N_11648,N_10765);
xor U13948 (N_13948,N_10339,N_10801);
and U13949 (N_13949,N_10412,N_10443);
nor U13950 (N_13950,N_11921,N_11924);
or U13951 (N_13951,N_10093,N_10168);
xnor U13952 (N_13952,N_11106,N_10023);
nor U13953 (N_13953,N_11695,N_11465);
or U13954 (N_13954,N_10955,N_11280);
nand U13955 (N_13955,N_10183,N_10028);
nor U13956 (N_13956,N_10945,N_11696);
and U13957 (N_13957,N_11787,N_10315);
xnor U13958 (N_13958,N_10893,N_10660);
nand U13959 (N_13959,N_11675,N_11980);
or U13960 (N_13960,N_11539,N_10588);
or U13961 (N_13961,N_10655,N_11709);
and U13962 (N_13962,N_11455,N_10583);
nor U13963 (N_13963,N_11680,N_10104);
xor U13964 (N_13964,N_11266,N_11896);
or U13965 (N_13965,N_10905,N_11345);
xnor U13966 (N_13966,N_10670,N_10622);
and U13967 (N_13967,N_11801,N_10462);
and U13968 (N_13968,N_10985,N_10479);
nand U13969 (N_13969,N_10896,N_10573);
nor U13970 (N_13970,N_10227,N_10129);
and U13971 (N_13971,N_10652,N_11500);
and U13972 (N_13972,N_10348,N_11821);
nor U13973 (N_13973,N_10478,N_11145);
xnor U13974 (N_13974,N_11937,N_11003);
nand U13975 (N_13975,N_10557,N_11966);
nor U13976 (N_13976,N_11333,N_11831);
xnor U13977 (N_13977,N_11790,N_10972);
nor U13978 (N_13978,N_10066,N_11124);
or U13979 (N_13979,N_10296,N_11915);
xnor U13980 (N_13980,N_10821,N_11531);
or U13981 (N_13981,N_11810,N_10358);
xor U13982 (N_13982,N_11095,N_11357);
or U13983 (N_13983,N_11800,N_11897);
and U13984 (N_13984,N_10671,N_10337);
and U13985 (N_13985,N_10583,N_10356);
xnor U13986 (N_13986,N_11991,N_11587);
nor U13987 (N_13987,N_10410,N_11452);
xnor U13988 (N_13988,N_11607,N_10852);
nor U13989 (N_13989,N_10425,N_10184);
or U13990 (N_13990,N_11832,N_11665);
nor U13991 (N_13991,N_10110,N_10114);
and U13992 (N_13992,N_11732,N_10414);
nor U13993 (N_13993,N_10563,N_11897);
nand U13994 (N_13994,N_11314,N_11826);
xnor U13995 (N_13995,N_11146,N_11017);
nor U13996 (N_13996,N_10681,N_11765);
nor U13997 (N_13997,N_10088,N_11643);
and U13998 (N_13998,N_11841,N_10038);
xnor U13999 (N_13999,N_10172,N_10096);
xor U14000 (N_14000,N_12621,N_13811);
nand U14001 (N_14001,N_13162,N_12034);
nand U14002 (N_14002,N_12714,N_12271);
xnor U14003 (N_14003,N_12517,N_12269);
and U14004 (N_14004,N_13922,N_12758);
xnor U14005 (N_14005,N_13023,N_12023);
or U14006 (N_14006,N_13862,N_12975);
nand U14007 (N_14007,N_13789,N_12777);
nor U14008 (N_14008,N_12501,N_12727);
xor U14009 (N_14009,N_12660,N_12837);
nand U14010 (N_14010,N_12265,N_12891);
and U14011 (N_14011,N_13988,N_12091);
and U14012 (N_14012,N_12244,N_12429);
nand U14013 (N_14013,N_13658,N_12450);
and U14014 (N_14014,N_13364,N_12619);
nand U14015 (N_14015,N_13823,N_13516);
and U14016 (N_14016,N_12054,N_12305);
nor U14017 (N_14017,N_13461,N_13555);
xor U14018 (N_14018,N_12536,N_13844);
and U14019 (N_14019,N_13170,N_12513);
nor U14020 (N_14020,N_13664,N_13424);
nand U14021 (N_14021,N_12459,N_12327);
and U14022 (N_14022,N_13764,N_12260);
nor U14023 (N_14023,N_12398,N_13877);
nor U14024 (N_14024,N_12437,N_12721);
nor U14025 (N_14025,N_13401,N_13523);
xnor U14026 (N_14026,N_12148,N_13778);
and U14027 (N_14027,N_13260,N_12942);
xnor U14028 (N_14028,N_12609,N_12208);
xor U14029 (N_14029,N_12041,N_13472);
xor U14030 (N_14030,N_12066,N_12038);
or U14031 (N_14031,N_12951,N_12635);
and U14032 (N_14032,N_13052,N_12578);
xnor U14033 (N_14033,N_13590,N_13095);
xnor U14034 (N_14034,N_12362,N_12728);
xnor U14035 (N_14035,N_12070,N_13887);
nand U14036 (N_14036,N_12137,N_13770);
nand U14037 (N_14037,N_12734,N_13258);
nand U14038 (N_14038,N_13596,N_13346);
nor U14039 (N_14039,N_13627,N_12707);
or U14040 (N_14040,N_13347,N_13528);
nand U14041 (N_14041,N_13728,N_13402);
nand U14042 (N_14042,N_12959,N_13598);
nand U14043 (N_14043,N_13883,N_12141);
xor U14044 (N_14044,N_12793,N_13431);
nand U14045 (N_14045,N_12620,N_12982);
and U14046 (N_14046,N_12639,N_13654);
xnor U14047 (N_14047,N_13915,N_12961);
nor U14048 (N_14048,N_13466,N_13135);
xnor U14049 (N_14049,N_12008,N_13827);
xor U14050 (N_14050,N_13803,N_13145);
nor U14051 (N_14051,N_12126,N_12489);
xor U14052 (N_14052,N_13699,N_13924);
xnor U14053 (N_14053,N_12644,N_12209);
nand U14054 (N_14054,N_13409,N_13666);
and U14055 (N_14055,N_13551,N_13760);
nand U14056 (N_14056,N_13386,N_12596);
and U14057 (N_14057,N_13489,N_12622);
or U14058 (N_14058,N_12523,N_12544);
or U14059 (N_14059,N_13259,N_12476);
nor U14060 (N_14060,N_12934,N_12974);
nand U14061 (N_14061,N_12992,N_13861);
nand U14062 (N_14062,N_13412,N_13394);
nand U14063 (N_14063,N_12379,N_13410);
nor U14064 (N_14064,N_12955,N_12742);
or U14065 (N_14065,N_13018,N_13396);
or U14066 (N_14066,N_13467,N_13136);
xor U14067 (N_14067,N_12252,N_13650);
and U14068 (N_14068,N_12462,N_13263);
and U14069 (N_14069,N_13281,N_12520);
xnor U14070 (N_14070,N_12706,N_13423);
or U14071 (N_14071,N_12823,N_12345);
nor U14072 (N_14072,N_13389,N_12401);
nor U14073 (N_14073,N_13985,N_13697);
nor U14074 (N_14074,N_12599,N_12096);
xor U14075 (N_14075,N_13578,N_13477);
and U14076 (N_14076,N_12083,N_13583);
and U14077 (N_14077,N_12545,N_13940);
and U14078 (N_14078,N_12205,N_13054);
nor U14079 (N_14079,N_12086,N_12568);
nand U14080 (N_14080,N_12831,N_13439);
and U14081 (N_14081,N_12119,N_13214);
and U14082 (N_14082,N_13548,N_13662);
and U14083 (N_14083,N_12580,N_13397);
nor U14084 (N_14084,N_13117,N_12525);
and U14085 (N_14085,N_13031,N_13190);
xnor U14086 (N_14086,N_13568,N_12120);
nor U14087 (N_14087,N_12024,N_13299);
nor U14088 (N_14088,N_12464,N_12369);
or U14089 (N_14089,N_12419,N_13616);
xor U14090 (N_14090,N_12819,N_13320);
nand U14091 (N_14091,N_12511,N_13206);
nand U14092 (N_14092,N_12025,N_13575);
and U14093 (N_14093,N_12512,N_12176);
and U14094 (N_14094,N_12189,N_12496);
nand U14095 (N_14095,N_12431,N_12297);
nand U14096 (N_14096,N_13788,N_13367);
nand U14097 (N_14097,N_13672,N_13769);
nor U14098 (N_14098,N_13264,N_13027);
nand U14099 (N_14099,N_12357,N_12550);
xnor U14100 (N_14100,N_12801,N_13607);
xnor U14101 (N_14101,N_13092,N_12627);
or U14102 (N_14102,N_13975,N_13909);
or U14103 (N_14103,N_12661,N_13348);
and U14104 (N_14104,N_13148,N_12076);
nor U14105 (N_14105,N_12842,N_13865);
or U14106 (N_14106,N_12902,N_13632);
xor U14107 (N_14107,N_12163,N_12057);
or U14108 (N_14108,N_13783,N_12172);
and U14109 (N_14109,N_13327,N_12486);
xor U14110 (N_14110,N_13330,N_13663);
and U14111 (N_14111,N_13942,N_13504);
xor U14112 (N_14112,N_13029,N_12637);
or U14113 (N_14113,N_12118,N_12900);
nand U14114 (N_14114,N_13073,N_13597);
or U14115 (N_14115,N_12233,N_13373);
xor U14116 (N_14116,N_12745,N_13043);
nor U14117 (N_14117,N_13237,N_12301);
or U14118 (N_14118,N_13983,N_12941);
or U14119 (N_14119,N_12918,N_13208);
nor U14120 (N_14120,N_13995,N_13161);
xor U14121 (N_14121,N_13384,N_12864);
xnor U14122 (N_14122,N_13318,N_13475);
nand U14123 (N_14123,N_12534,N_13441);
or U14124 (N_14124,N_12908,N_12111);
nor U14125 (N_14125,N_12946,N_13956);
nand U14126 (N_14126,N_13335,N_13715);
nor U14127 (N_14127,N_12863,N_12963);
xor U14128 (N_14128,N_12711,N_12216);
xnor U14129 (N_14129,N_12591,N_12457);
xor U14130 (N_14130,N_13154,N_13670);
xnor U14131 (N_14131,N_12700,N_13229);
nand U14132 (N_14132,N_12328,N_13037);
nand U14133 (N_14133,N_13338,N_12556);
and U14134 (N_14134,N_13171,N_12535);
nor U14135 (N_14135,N_13351,N_13970);
or U14136 (N_14136,N_13668,N_12870);
xnor U14137 (N_14137,N_13453,N_12257);
or U14138 (N_14138,N_12883,N_13837);
xor U14139 (N_14139,N_12505,N_13741);
and U14140 (N_14140,N_13797,N_13560);
xnor U14141 (N_14141,N_13533,N_13566);
nand U14142 (N_14142,N_13074,N_12330);
nand U14143 (N_14143,N_12887,N_13511);
nor U14144 (N_14144,N_12344,N_12844);
nor U14145 (N_14145,N_12720,N_12434);
nand U14146 (N_14146,N_13552,N_13251);
and U14147 (N_14147,N_13382,N_13687);
nand U14148 (N_14148,N_12791,N_12962);
nor U14149 (N_14149,N_13964,N_13456);
or U14150 (N_14150,N_13089,N_13957);
nand U14151 (N_14151,N_12387,N_12248);
nand U14152 (N_14152,N_13468,N_13825);
or U14153 (N_14153,N_12895,N_13896);
nor U14154 (N_14154,N_12651,N_13767);
and U14155 (N_14155,N_12697,N_12164);
or U14156 (N_14156,N_12125,N_13250);
xor U14157 (N_14157,N_12368,N_12866);
nor U14158 (N_14158,N_13619,N_12798);
or U14159 (N_14159,N_12061,N_13064);
nor U14160 (N_14160,N_12004,N_13725);
and U14161 (N_14161,N_13180,N_13897);
xor U14162 (N_14162,N_13355,N_13143);
nor U14163 (N_14163,N_13990,N_12068);
nor U14164 (N_14164,N_12717,N_13682);
or U14165 (N_14165,N_12846,N_13657);
or U14166 (N_14166,N_12084,N_12173);
xor U14167 (N_14167,N_13199,N_12736);
xnor U14168 (N_14168,N_12017,N_13804);
nand U14169 (N_14169,N_12931,N_13509);
or U14170 (N_14170,N_13480,N_12056);
and U14171 (N_14171,N_13539,N_13246);
nand U14172 (N_14172,N_13033,N_12985);
and U14173 (N_14173,N_13813,N_13950);
or U14174 (N_14174,N_13028,N_12080);
and U14175 (N_14175,N_13809,N_12543);
or U14176 (N_14176,N_13659,N_13763);
and U14177 (N_14177,N_12147,N_12191);
xnor U14178 (N_14178,N_13391,N_13230);
or U14179 (N_14179,N_12658,N_12286);
nor U14180 (N_14180,N_12333,N_12442);
and U14181 (N_14181,N_13352,N_13243);
xor U14182 (N_14182,N_12220,N_12217);
and U14183 (N_14183,N_12641,N_12200);
nand U14184 (N_14184,N_12779,N_12263);
nand U14185 (N_14185,N_13300,N_12557);
nor U14186 (N_14186,N_13071,N_12304);
nand U14187 (N_14187,N_12806,N_13164);
xor U14188 (N_14188,N_12821,N_13128);
xnor U14189 (N_14189,N_13131,N_13853);
nand U14190 (N_14190,N_13139,N_12753);
and U14191 (N_14191,N_12789,N_13458);
and U14192 (N_14192,N_13100,N_12548);
nand U14193 (N_14193,N_12022,N_13044);
xnor U14194 (N_14194,N_12324,N_13935);
nand U14195 (N_14195,N_13189,N_13637);
and U14196 (N_14196,N_13280,N_12136);
or U14197 (N_14197,N_12766,N_12944);
and U14198 (N_14198,N_12293,N_12378);
or U14199 (N_14199,N_12461,N_12843);
and U14200 (N_14200,N_12146,N_13540);
and U14201 (N_14201,N_13780,N_12029);
or U14202 (N_14202,N_13313,N_13898);
or U14203 (N_14203,N_13297,N_12987);
nor U14204 (N_14204,N_13270,N_13278);
xor U14205 (N_14205,N_13012,N_13223);
xor U14206 (N_14206,N_12785,N_13432);
or U14207 (N_14207,N_12978,N_12834);
xor U14208 (N_14208,N_13009,N_12782);
nor U14209 (N_14209,N_12225,N_12285);
nor U14210 (N_14210,N_13236,N_12813);
nand U14211 (N_14211,N_12530,N_12308);
or U14212 (N_14212,N_13217,N_13919);
nand U14213 (N_14213,N_12958,N_12047);
nor U14214 (N_14214,N_13091,N_13062);
nand U14215 (N_14215,N_13416,N_13717);
xor U14216 (N_14216,N_12059,N_13448);
nor U14217 (N_14217,N_12007,N_13706);
or U14218 (N_14218,N_13179,N_12219);
xnor U14219 (N_14219,N_13003,N_12935);
or U14220 (N_14220,N_13869,N_12010);
nor U14221 (N_14221,N_12049,N_13253);
or U14222 (N_14222,N_13872,N_13067);
and U14223 (N_14223,N_13928,N_13541);
or U14224 (N_14224,N_13363,N_13361);
xnor U14225 (N_14225,N_12889,N_13153);
or U14226 (N_14226,N_13269,N_12521);
nor U14227 (N_14227,N_13016,N_13852);
xor U14228 (N_14228,N_12073,N_12704);
nand U14229 (N_14229,N_13201,N_12236);
xor U14230 (N_14230,N_12183,N_13221);
nor U14231 (N_14231,N_13104,N_12374);
and U14232 (N_14232,N_12677,N_12207);
xnor U14233 (N_14233,N_12764,N_13951);
nand U14234 (N_14234,N_13714,N_13017);
nor U14235 (N_14235,N_13974,N_12417);
nor U14236 (N_14236,N_12816,N_12593);
nand U14237 (N_14237,N_12759,N_13188);
xnor U14238 (N_14238,N_13709,N_12203);
nor U14239 (N_14239,N_12185,N_12321);
or U14240 (N_14240,N_13061,N_12940);
or U14241 (N_14241,N_13010,N_12649);
nand U14242 (N_14242,N_13537,N_13166);
or U14243 (N_14243,N_13870,N_13362);
and U14244 (N_14244,N_12326,N_12625);
nand U14245 (N_14245,N_12581,N_12048);
xnor U14246 (N_14246,N_12776,N_13357);
nor U14247 (N_14247,N_13965,N_13090);
xor U14248 (N_14248,N_12972,N_12830);
xnor U14249 (N_14249,N_12192,N_13077);
nand U14250 (N_14250,N_13726,N_13337);
nand U14251 (N_14251,N_13864,N_13372);
or U14252 (N_14252,N_13365,N_13249);
nand U14253 (N_14253,N_12320,N_13773);
nand U14254 (N_14254,N_13748,N_12366);
and U14255 (N_14255,N_13200,N_12629);
or U14256 (N_14256,N_13058,N_13354);
or U14257 (N_14257,N_13271,N_12762);
xor U14258 (N_14258,N_12748,N_13169);
and U14259 (N_14259,N_13833,N_12569);
and U14260 (N_14260,N_13903,N_12896);
and U14261 (N_14261,N_12733,N_12970);
nor U14262 (N_14262,N_12969,N_13910);
nand U14263 (N_14263,N_13045,N_13634);
xnor U14264 (N_14264,N_13007,N_12381);
nand U14265 (N_14265,N_12538,N_12926);
xnor U14266 (N_14266,N_13737,N_12334);
nor U14267 (N_14267,N_12829,N_12309);
nor U14268 (N_14268,N_12675,N_13937);
nand U14269 (N_14269,N_13945,N_13488);
and U14270 (N_14270,N_13437,N_13425);
nor U14271 (N_14271,N_12913,N_12740);
nor U14272 (N_14272,N_13265,N_12143);
and U14273 (N_14273,N_12968,N_12838);
xor U14274 (N_14274,N_13857,N_13105);
or U14275 (N_14275,N_12037,N_13806);
nor U14276 (N_14276,N_12983,N_13195);
or U14277 (N_14277,N_13859,N_12994);
xor U14278 (N_14278,N_12355,N_13931);
xnor U14279 (N_14279,N_13233,N_13839);
and U14280 (N_14280,N_13304,N_13157);
xnor U14281 (N_14281,N_13828,N_12161);
xor U14282 (N_14282,N_13652,N_12647);
nor U14283 (N_14283,N_13899,N_12528);
or U14284 (N_14284,N_12522,N_13810);
xor U14285 (N_14285,N_13621,N_12905);
and U14286 (N_14286,N_13505,N_12425);
or U14287 (N_14287,N_12370,N_12341);
or U14288 (N_14288,N_12188,N_13359);
xor U14289 (N_14289,N_13081,N_13563);
nor U14290 (N_14290,N_12139,N_12155);
or U14291 (N_14291,N_12854,N_13691);
or U14292 (N_14292,N_12104,N_13589);
and U14293 (N_14293,N_12473,N_13805);
nor U14294 (N_14294,N_12346,N_13601);
or U14295 (N_14295,N_12919,N_12853);
xor U14296 (N_14296,N_12453,N_13522);
or U14297 (N_14297,N_13078,N_13298);
xnor U14298 (N_14298,N_12703,N_12712);
and U14299 (N_14299,N_13414,N_13655);
and U14300 (N_14300,N_13464,N_12045);
nand U14301 (N_14301,N_12768,N_13836);
nor U14302 (N_14302,N_12588,N_12395);
nand U14303 (N_14303,N_13776,N_13499);
and U14304 (N_14304,N_12805,N_13826);
and U14305 (N_14305,N_12373,N_13585);
nor U14306 (N_14306,N_12912,N_13317);
or U14307 (N_14307,N_13182,N_12995);
nor U14308 (N_14308,N_12165,N_13186);
xor U14309 (N_14309,N_13344,N_12065);
and U14310 (N_14310,N_13422,N_13377);
or U14311 (N_14311,N_13000,N_12563);
xnor U14312 (N_14312,N_12325,N_12726);
xor U14313 (N_14313,N_12744,N_12484);
and U14314 (N_14314,N_12615,N_12474);
and U14315 (N_14315,N_13876,N_12289);
xor U14316 (N_14316,N_12986,N_13938);
xor U14317 (N_14317,N_12645,N_13577);
or U14318 (N_14318,N_12212,N_12901);
and U14319 (N_14319,N_13106,N_13707);
nand U14320 (N_14320,N_13415,N_12943);
nor U14321 (N_14321,N_13724,N_13015);
nand U14322 (N_14322,N_12678,N_13411);
and U14323 (N_14323,N_12755,N_13754);
nand U14324 (N_14324,N_12053,N_13683);
xor U14325 (N_14325,N_12732,N_12775);
and U14326 (N_14326,N_12804,N_12526);
and U14327 (N_14327,N_12685,N_13759);
nand U14328 (N_14328,N_13679,N_13315);
nor U14329 (N_14329,N_13267,N_12796);
and U14330 (N_14330,N_13483,N_13216);
nand U14331 (N_14331,N_12890,N_12094);
and U14332 (N_14332,N_13930,N_13309);
nand U14333 (N_14333,N_12152,N_13019);
or U14334 (N_14334,N_12290,N_12452);
or U14335 (N_14335,N_12662,N_12067);
xor U14336 (N_14336,N_13305,N_12306);
and U14337 (N_14337,N_12549,N_12062);
nand U14338 (N_14338,N_13629,N_12154);
nor U14339 (N_14339,N_13600,N_13992);
and U14340 (N_14340,N_13656,N_12093);
nand U14341 (N_14341,N_13450,N_13534);
xor U14342 (N_14342,N_13639,N_12030);
or U14343 (N_14343,N_12198,N_12175);
and U14344 (N_14344,N_12767,N_13503);
and U14345 (N_14345,N_12696,N_13158);
or U14346 (N_14346,N_13495,N_12936);
nand U14347 (N_14347,N_12773,N_13701);
nor U14348 (N_14348,N_13614,N_13660);
nand U14349 (N_14349,N_12903,N_13481);
nand U14350 (N_14350,N_13113,N_12235);
and U14351 (N_14351,N_13508,N_12052);
nor U14352 (N_14352,N_12784,N_12638);
or U14353 (N_14353,N_13736,N_13474);
nor U14354 (N_14354,N_13526,N_12214);
and U14355 (N_14355,N_12412,N_12110);
xnor U14356 (N_14356,N_12769,N_13675);
nand U14357 (N_14357,N_13604,N_12221);
xnor U14358 (N_14358,N_12230,N_13832);
nor U14359 (N_14359,N_12018,N_12405);
and U14360 (N_14360,N_12190,N_13841);
xor U14361 (N_14361,N_12817,N_13635);
xor U14362 (N_14362,N_13623,N_13417);
xnor U14363 (N_14363,N_13349,N_13376);
or U14364 (N_14364,N_13093,N_12433);
nand U14365 (N_14365,N_13421,N_12443);
and U14366 (N_14366,N_12404,N_12710);
or U14367 (N_14367,N_13119,N_12331);
nor U14368 (N_14368,N_13677,N_13676);
nor U14369 (N_14369,N_12210,N_13399);
nand U14370 (N_14370,N_12998,N_12546);
nor U14371 (N_14371,N_12151,N_13661);
xnor U14372 (N_14372,N_12674,N_13114);
xor U14373 (N_14373,N_12015,N_12131);
nor U14374 (N_14374,N_13068,N_13066);
nand U14375 (N_14375,N_12640,N_12044);
nor U14376 (N_14376,N_13907,N_13339);
and U14377 (N_14377,N_12624,N_12652);
xnor U14378 (N_14378,N_13514,N_13690);
nor U14379 (N_14379,N_12140,N_12441);
or U14380 (N_14380,N_12403,N_12855);
xnor U14381 (N_14381,N_13969,N_12224);
and U14382 (N_14382,N_13213,N_12466);
nand U14383 (N_14383,N_12689,N_13333);
xnor U14384 (N_14384,N_12988,N_12507);
or U14385 (N_14385,N_12449,N_12444);
and U14386 (N_14386,N_13149,N_13004);
nand U14387 (N_14387,N_12105,N_13184);
or U14388 (N_14388,N_13231,N_12514);
and U14389 (N_14389,N_12106,N_12026);
nand U14390 (N_14390,N_12835,N_12349);
and U14391 (N_14391,N_12885,N_13484);
nand U14392 (N_14392,N_13746,N_13490);
xnor U14393 (N_14393,N_13025,N_13099);
or U14394 (N_14394,N_12980,N_12339);
and U14395 (N_14395,N_13144,N_13151);
xnor U14396 (N_14396,N_12012,N_13102);
nor U14397 (N_14397,N_13711,N_13856);
or U14398 (N_14398,N_13406,N_12623);
xnor U14399 (N_14399,N_13020,N_13847);
and U14400 (N_14400,N_12033,N_13288);
nand U14401 (N_14401,N_12232,N_12876);
nand U14402 (N_14402,N_12976,N_12268);
nor U14403 (N_14403,N_13550,N_12575);
and U14404 (N_14404,N_12950,N_12158);
and U14405 (N_14405,N_13486,N_12856);
xnor U14406 (N_14406,N_12351,N_13374);
nand U14407 (N_14407,N_13294,N_13591);
nor U14408 (N_14408,N_13643,N_12127);
nor U14409 (N_14409,N_13881,N_13220);
or U14410 (N_14410,N_13408,N_12089);
nand U14411 (N_14411,N_12731,N_12423);
nand U14412 (N_14412,N_12307,N_12868);
nand U14413 (N_14413,N_13047,N_12234);
xnor U14414 (N_14414,N_13603,N_13863);
xnor U14415 (N_14415,N_13479,N_12256);
nand U14416 (N_14416,N_12613,N_12541);
nor U14417 (N_14417,N_13311,N_13642);
nor U14418 (N_14418,N_13400,N_12803);
or U14419 (N_14419,N_13168,N_12187);
or U14420 (N_14420,N_12611,N_13048);
nand U14421 (N_14421,N_12006,N_13611);
nand U14422 (N_14422,N_13358,N_13625);
xnor U14423 (N_14423,N_13610,N_12240);
xnor U14424 (N_14424,N_12348,N_12312);
and U14425 (N_14425,N_13174,N_13118);
nand U14426 (N_14426,N_12284,N_13996);
xnor U14427 (N_14427,N_12427,N_12494);
xor U14428 (N_14428,N_13124,N_12953);
xnor U14429 (N_14429,N_13702,N_12595);
or U14430 (N_14430,N_13757,N_12971);
and U14431 (N_14431,N_13430,N_13569);
or U14432 (N_14432,N_12617,N_13713);
xor U14433 (N_14433,N_12894,N_12997);
nor U14434 (N_14434,N_13482,N_12359);
xnor U14435 (N_14435,N_13984,N_13096);
nand U14436 (N_14436,N_13860,N_13167);
or U14437 (N_14437,N_13226,N_13491);
and U14438 (N_14438,N_13648,N_12222);
nor U14439 (N_14439,N_12999,N_12394);
or U14440 (N_14440,N_13981,N_13120);
nand U14441 (N_14441,N_13427,N_13172);
or U14442 (N_14442,N_12150,N_13842);
nand U14443 (N_14443,N_12562,N_13319);
or U14444 (N_14444,N_13649,N_13274);
xor U14445 (N_14445,N_12532,N_13039);
xnor U14446 (N_14446,N_13973,N_13292);
or U14447 (N_14447,N_13262,N_13605);
and U14448 (N_14448,N_13185,N_12113);
or U14449 (N_14449,N_13807,N_12787);
nor U14450 (N_14450,N_12383,N_13248);
nor U14451 (N_14451,N_13532,N_13133);
and U14452 (N_14452,N_12414,N_12977);
xor U14453 (N_14453,N_12709,N_13556);
or U14454 (N_14454,N_12099,N_12589);
nor U14455 (N_14455,N_13447,N_13356);
and U14456 (N_14456,N_12238,N_12107);
xnor U14457 (N_14457,N_13465,N_13586);
or U14458 (N_14458,N_13991,N_13176);
nor U14459 (N_14459,N_12211,N_13177);
xor U14460 (N_14460,N_13094,N_12179);
nand U14461 (N_14461,N_12991,N_13761);
nor U14462 (N_14462,N_12979,N_12747);
and U14463 (N_14463,N_12166,N_13669);
or U14464 (N_14464,N_12114,N_12402);
nor U14465 (N_14465,N_13429,N_12739);
nor U14466 (N_14466,N_12656,N_13946);
and U14467 (N_14467,N_13147,N_13006);
nor U14468 (N_14468,N_12223,N_13261);
and U14469 (N_14469,N_12914,N_13943);
xnor U14470 (N_14470,N_12391,N_12646);
nor U14471 (N_14471,N_13116,N_12552);
xor U14472 (N_14472,N_12115,N_13204);
nand U14473 (N_14473,N_13041,N_12565);
xor U14474 (N_14474,N_13350,N_12392);
xor U14475 (N_14475,N_12439,N_12071);
xor U14476 (N_14476,N_12249,N_12292);
or U14477 (N_14477,N_12583,N_12456);
nor U14478 (N_14478,N_12138,N_12828);
nor U14479 (N_14479,N_13059,N_12701);
xnor U14480 (N_14480,N_12409,N_12181);
and U14481 (N_14481,N_12799,N_12833);
xnor U14482 (N_14482,N_13613,N_13911);
nor U14483 (N_14483,N_12035,N_13287);
xor U14484 (N_14484,N_13933,N_13470);
nor U14485 (N_14485,N_12072,N_12451);
nor U14486 (N_14486,N_12261,N_12653);
nor U14487 (N_14487,N_13570,N_13908);
nor U14488 (N_14488,N_13747,N_12278);
nor U14489 (N_14489,N_12797,N_12245);
nor U14490 (N_14490,N_12648,N_13443);
or U14491 (N_14491,N_13460,N_12122);
xor U14492 (N_14492,N_12276,N_13111);
nor U14493 (N_14493,N_13155,N_13684);
nor U14494 (N_14494,N_12472,N_13112);
nor U14495 (N_14495,N_13390,N_13801);
nand U14496 (N_14496,N_13520,N_13463);
nand U14497 (N_14497,N_13868,N_12664);
nand U14498 (N_14498,N_13492,N_13192);
and U14499 (N_14499,N_13507,N_12332);
nand U14500 (N_14500,N_12917,N_12280);
nor U14501 (N_14501,N_12195,N_12614);
xor U14502 (N_14502,N_13183,N_13793);
and U14503 (N_14503,N_12168,N_12407);
and U14504 (N_14504,N_13301,N_12347);
or U14505 (N_14505,N_13678,N_12531);
or U14506 (N_14506,N_12227,N_13434);
nor U14507 (N_14507,N_13609,N_12186);
xor U14508 (N_14508,N_13719,N_13873);
nor U14509 (N_14509,N_12482,N_12760);
nand U14510 (N_14510,N_12718,N_12241);
and U14511 (N_14511,N_12342,N_12947);
nor U14512 (N_14512,N_12862,N_12133);
nor U14513 (N_14513,N_12681,N_13846);
nand U14514 (N_14514,N_13593,N_12471);
nor U14515 (N_14515,N_12586,N_13976);
nor U14516 (N_14516,N_13257,N_12371);
nor U14517 (N_14517,N_13925,N_12719);
and U14518 (N_14518,N_13316,N_12898);
or U14519 (N_14519,N_12920,N_12322);
or U14520 (N_14520,N_12087,N_13703);
nor U14521 (N_14521,N_13291,N_13673);
xor U14522 (N_14522,N_12508,N_13755);
xor U14523 (N_14523,N_12515,N_12281);
and U14524 (N_14524,N_13245,N_13051);
xnor U14525 (N_14525,N_13816,N_12415);
xnor U14526 (N_14526,N_13360,N_12178);
nor U14527 (N_14527,N_13275,N_13721);
nor U14528 (N_14528,N_12650,N_13562);
xnor U14529 (N_14529,N_12364,N_12690);
nand U14530 (N_14530,N_13108,N_12966);
and U14531 (N_14531,N_13784,N_13446);
nor U14532 (N_14532,N_12295,N_13955);
or U14533 (N_14533,N_12663,N_13238);
or U14534 (N_14534,N_12852,N_12691);
nand U14535 (N_14535,N_12673,N_12723);
or U14536 (N_14536,N_12399,N_12795);
or U14537 (N_14537,N_13695,N_12516);
or U14538 (N_14538,N_12888,N_12922);
xor U14539 (N_14539,N_13917,N_12079);
or U14540 (N_14540,N_12375,N_13024);
xnor U14541 (N_14541,N_12610,N_13653);
and U14542 (N_14542,N_13038,N_12577);
and U14543 (N_14543,N_13843,N_13057);
nor U14544 (N_14544,N_13014,N_12790);
nor U14545 (N_14545,N_13921,N_12708);
and U14546 (N_14546,N_12353,N_12386);
or U14547 (N_14547,N_13215,N_13980);
or U14548 (N_14548,N_13734,N_13752);
or U14549 (N_14549,N_12272,N_12134);
nor U14550 (N_14550,N_13326,N_12050);
nand U14551 (N_14551,N_12906,N_12877);
and U14552 (N_14552,N_13314,N_13125);
or U14553 (N_14553,N_13579,N_12128);
and U14554 (N_14554,N_12820,N_12682);
nand U14555 (N_14555,N_13130,N_12825);
or U14556 (N_14556,N_12377,N_13786);
or U14557 (N_14557,N_13893,N_12448);
nand U14558 (N_14558,N_13718,N_12875);
or U14559 (N_14559,N_13849,N_13247);
nor U14560 (N_14560,N_12028,N_13543);
or U14561 (N_14561,N_12213,N_12410);
nor U14562 (N_14562,N_12822,N_12440);
nor U14563 (N_14563,N_12911,N_12561);
nand U14564 (N_14564,N_13971,N_12078);
xor U14565 (N_14565,N_12098,N_12698);
and U14566 (N_14566,N_12487,N_13395);
or U14567 (N_14567,N_12074,N_13599);
xor U14568 (N_14568,N_12800,N_12435);
or U14569 (N_14569,N_13065,N_13584);
and U14570 (N_14570,N_12116,N_13889);
and U14571 (N_14571,N_13912,N_13875);
or U14572 (N_14572,N_13498,N_13224);
nand U14573 (N_14573,N_13779,N_12882);
nor U14574 (N_14574,N_12483,N_12576);
or U14575 (N_14575,N_12046,N_12695);
xor U14576 (N_14576,N_12117,N_13011);
nand U14577 (N_14577,N_12335,N_13594);
and U14578 (N_14578,N_13733,N_13252);
nor U14579 (N_14579,N_12848,N_12454);
nand U14580 (N_14580,N_13080,N_13765);
and U14581 (N_14581,N_12291,N_12478);
and U14582 (N_14582,N_13002,N_13606);
xnor U14583 (N_14583,N_13030,N_13999);
xor U14584 (N_14584,N_13704,N_12989);
and U14585 (N_14585,N_12361,N_12849);
and U14586 (N_14586,N_13075,N_13063);
nor U14587 (N_14587,N_12606,N_13978);
nor U14588 (N_14588,N_13972,N_12380);
and U14589 (N_14589,N_13927,N_13282);
or U14590 (N_14590,N_12356,N_12812);
or U14591 (N_14591,N_12628,N_12460);
and U14592 (N_14592,N_13444,N_13542);
nand U14593 (N_14593,N_13830,N_12430);
or U14594 (N_14594,N_13729,N_12382);
or U14595 (N_14595,N_13165,N_13771);
nor U14596 (N_14596,N_13502,N_12503);
nor U14597 (N_14597,N_13471,N_13581);
xor U14598 (N_14598,N_13743,N_12097);
nand U14599 (N_14599,N_12201,N_12036);
nand U14600 (N_14600,N_12679,N_12878);
xnor U14601 (N_14601,N_13496,N_13953);
nor U14602 (N_14602,N_13564,N_12019);
or U14603 (N_14603,N_12300,N_13109);
nor U14604 (N_14604,N_12716,N_12555);
or U14605 (N_14605,N_13266,N_13561);
nand U14606 (N_14606,N_13554,N_12850);
xnor U14607 (N_14607,N_12964,N_13032);
and U14608 (N_14608,N_13325,N_12749);
nor U14609 (N_14609,N_12879,N_12884);
nand U14610 (N_14610,N_13510,N_13798);
or U14611 (N_14611,N_13273,N_12996);
nand U14612 (N_14612,N_13110,N_13982);
nor U14613 (N_14613,N_13628,N_13799);
nand U14614 (N_14614,N_12927,N_13055);
nor U14615 (N_14615,N_13815,N_13366);
xnor U14616 (N_14616,N_13934,N_13608);
nand U14617 (N_14617,N_12069,N_12671);
or U14618 (N_14618,N_12318,N_12954);
nor U14619 (N_14619,N_13196,N_12510);
or U14620 (N_14620,N_13735,N_12930);
nand U14621 (N_14621,N_12329,N_12529);
nor U14622 (N_14622,N_12929,N_12250);
and U14623 (N_14623,N_13840,N_13892);
or U14624 (N_14624,N_13920,N_12794);
nor U14625 (N_14625,N_12389,N_12488);
nand U14626 (N_14626,N_12090,N_13531);
or U14627 (N_14627,N_12527,N_12169);
or U14628 (N_14628,N_12874,N_13817);
xnor U14629 (N_14629,N_12206,N_12783);
and U14630 (N_14630,N_12693,N_13225);
xor U14631 (N_14631,N_13385,N_12860);
and U14632 (N_14632,N_13744,N_13835);
xor U14633 (N_14633,N_12949,N_13134);
xnor U14634 (N_14634,N_13152,N_12746);
xor U14635 (N_14635,N_13205,N_13671);
and U14636 (N_14636,N_13756,N_12909);
or U14637 (N_14637,N_12124,N_13254);
and U14638 (N_14638,N_12253,N_12547);
or U14639 (N_14639,N_13775,N_13285);
nand U14640 (N_14640,N_12818,N_13939);
nand U14641 (N_14641,N_12702,N_12063);
nor U14642 (N_14642,N_13521,N_12851);
xnor U14643 (N_14643,N_13538,N_13913);
xor U14644 (N_14644,N_13478,N_12493);
nor U14645 (N_14645,N_12101,N_13138);
nor U14646 (N_14646,N_12129,N_13622);
nor U14647 (N_14647,N_13159,N_13076);
xnor U14648 (N_14648,N_12824,N_12204);
and U14649 (N_14649,N_13500,N_13567);
nand U14650 (N_14650,N_13888,N_12132);
nand U14651 (N_14651,N_12730,N_12757);
nand U14652 (N_14652,N_13440,N_13203);
or U14653 (N_14653,N_12587,N_12631);
or U14654 (N_14654,N_12317,N_13885);
nor U14655 (N_14655,N_12772,N_13485);
and U14656 (N_14656,N_13963,N_12103);
nor U14657 (N_14657,N_12765,N_12315);
nand U14658 (N_14658,N_12737,N_13886);
nand U14659 (N_14659,N_13941,N_12159);
xor U14660 (N_14660,N_12495,N_13345);
nand U14661 (N_14661,N_13553,N_13302);
nand U14662 (N_14662,N_13272,N_13947);
xor U14663 (N_14663,N_13966,N_12319);
xnor U14664 (N_14664,N_12607,N_13459);
xnor U14665 (N_14665,N_12447,N_12400);
nor U14666 (N_14666,N_12060,N_13914);
xnor U14667 (N_14667,N_13722,N_13380);
nand U14668 (N_14668,N_13122,N_12490);
nor U14669 (N_14669,N_13751,N_12761);
nor U14670 (N_14670,N_12579,N_12886);
or U14671 (N_14671,N_12396,N_12756);
or U14672 (N_14672,N_12725,N_13546);
nor U14673 (N_14673,N_13086,N_13800);
or U14674 (N_14674,N_13035,N_13381);
nand U14675 (N_14675,N_12130,N_12925);
xnor U14676 (N_14676,N_13328,N_12258);
xor U14677 (N_14677,N_12215,N_13615);
or U14678 (N_14678,N_12560,N_12102);
nand U14679 (N_14679,N_12670,N_13487);
xnor U14680 (N_14680,N_12492,N_13993);
xnor U14681 (N_14681,N_13878,N_12055);
xnor U14682 (N_14682,N_13083,N_13519);
xor U14683 (N_14683,N_12600,N_13536);
or U14684 (N_14684,N_12519,N_13121);
and U14685 (N_14685,N_13565,N_13831);
xor U14686 (N_14686,N_12872,N_12633);
and U14687 (N_14687,N_12752,N_13227);
nand U14688 (N_14688,N_12873,N_13242);
or U14689 (N_14689,N_13693,N_12153);
nor U14690 (N_14690,N_13322,N_13895);
nor U14691 (N_14691,N_12310,N_13060);
and U14692 (N_14692,N_12729,N_12741);
or U14693 (N_14693,N_13187,N_12277);
xnor U14694 (N_14694,N_12585,N_12171);
nor U14695 (N_14695,N_13462,N_13084);
or U14696 (N_14696,N_12475,N_13867);
xnor U14697 (N_14697,N_12014,N_13680);
nand U14698 (N_14698,N_13334,N_12180);
nor U14699 (N_14699,N_13904,N_13962);
or U14700 (N_14700,N_13276,N_13644);
or U14701 (N_14701,N_12021,N_13329);
nor U14702 (N_14702,N_13812,N_12524);
xor U14703 (N_14703,N_13636,N_12567);
nor U14704 (N_14704,N_13774,N_12384);
nor U14705 (N_14705,N_12666,N_13087);
nor U14706 (N_14706,N_13088,N_13640);
or U14707 (N_14707,N_13383,N_12597);
or U14708 (N_14708,N_12455,N_13766);
nor U14709 (N_14709,N_12463,N_12770);
nand U14710 (N_14710,N_13126,N_12182);
or U14711 (N_14711,N_12254,N_13900);
xor U14712 (N_14712,N_12956,N_13103);
nand U14713 (N_14713,N_12612,N_13438);
or U14714 (N_14714,N_12156,N_12857);
xnor U14715 (N_14715,N_12299,N_13960);
nand U14716 (N_14716,N_12603,N_13008);
or U14717 (N_14717,N_12932,N_12665);
or U14718 (N_14718,N_12422,N_12338);
xnor U14719 (N_14719,N_13858,N_13306);
and U14720 (N_14720,N_12559,N_12807);
xor U14721 (N_14721,N_12426,N_12683);
xnor U14722 (N_14722,N_12584,N_13290);
or U14723 (N_14723,N_12509,N_12916);
nor U14724 (N_14724,N_12479,N_13712);
nand U14725 (N_14725,N_13944,N_13574);
and U14726 (N_14726,N_13056,N_13515);
nand U14727 (N_14727,N_12602,N_13716);
and U14728 (N_14728,N_13961,N_13626);
or U14729 (N_14729,N_12287,N_12467);
nand U14730 (N_14730,N_13689,N_13557);
or U14731 (N_14731,N_13193,N_13219);
nor U14732 (N_14732,N_12432,N_12288);
or U14733 (N_14733,N_12810,N_12808);
nand U14734 (N_14734,N_12273,N_13730);
xor U14735 (N_14735,N_13781,N_12899);
xnor U14736 (N_14736,N_13371,N_13049);
nand U14737 (N_14737,N_13240,N_13796);
nand U14738 (N_14738,N_12081,N_13738);
nand U14739 (N_14739,N_13977,N_12397);
or U14740 (N_14740,N_12242,N_12420);
xor U14741 (N_14741,N_13332,N_12100);
or U14742 (N_14742,N_13255,N_13244);
xnor U14743 (N_14743,N_13645,N_13884);
nand U14744 (N_14744,N_13082,N_12194);
nand U14745 (N_14745,N_13494,N_12497);
and U14746 (N_14746,N_12771,N_13323);
xor U14747 (N_14747,N_12376,N_12694);
or U14748 (N_14748,N_13241,N_13968);
and U14749 (N_14749,N_13127,N_13405);
nand U14750 (N_14750,N_12788,N_13178);
nor U14751 (N_14751,N_12485,N_12121);
and U14752 (N_14752,N_12313,N_13795);
nand U14753 (N_14753,N_12112,N_13293);
or U14754 (N_14754,N_13705,N_13512);
or U14755 (N_14755,N_13501,N_12246);
or U14756 (N_14756,N_13851,N_13378);
nor U14757 (N_14757,N_13822,N_13918);
nand U14758 (N_14758,N_13692,N_13854);
and U14759 (N_14759,N_13808,N_12571);
nand U14760 (N_14760,N_13517,N_12196);
xnor U14761 (N_14761,N_13700,N_12616);
or U14762 (N_14762,N_13994,N_13544);
and U14763 (N_14763,N_13341,N_13140);
nand U14764 (N_14764,N_12655,N_12239);
and U14765 (N_14765,N_13638,N_12643);
nand U14766 (N_14766,N_13005,N_13156);
nor U14767 (N_14767,N_12667,N_13753);
xnor U14768 (N_14768,N_12780,N_13173);
nand U14769 (N_14769,N_12945,N_13954);
xnor U14770 (N_14770,N_13630,N_13279);
nand U14771 (N_14771,N_12705,N_12303);
nor U14772 (N_14772,N_13129,N_13959);
xnor U14773 (N_14773,N_12385,N_12247);
nand U14774 (N_14774,N_12928,N_12296);
nand U14775 (N_14775,N_13549,N_13449);
nor U14776 (N_14776,N_13079,N_12157);
nor U14777 (N_14777,N_13469,N_12418);
xor U14778 (N_14778,N_13150,N_12064);
or U14779 (N_14779,N_13518,N_13454);
nor U14780 (N_14780,N_12792,N_12294);
nor U14781 (N_14781,N_12684,N_13286);
xor U14782 (N_14782,N_13790,N_12781);
nor U14783 (N_14783,N_13455,N_12880);
nand U14784 (N_14784,N_12095,N_13207);
nor U14785 (N_14785,N_13310,N_13026);
or U14786 (N_14786,N_12582,N_13633);
or U14787 (N_14787,N_12910,N_12408);
and U14788 (N_14788,N_12088,N_12270);
nand U14789 (N_14789,N_13997,N_13595);
nand U14790 (N_14790,N_13407,N_12938);
xor U14791 (N_14791,N_12274,N_13681);
xor U14792 (N_14792,N_12406,N_12003);
xnor U14793 (N_14793,N_12144,N_12573);
and U14794 (N_14794,N_12993,N_13525);
xnor U14795 (N_14795,N_12750,N_13979);
or U14796 (N_14796,N_12160,N_13894);
nor U14797 (N_14797,N_12657,N_12537);
and U14798 (N_14798,N_12424,N_13785);
xnor U14799 (N_14799,N_12499,N_13436);
nor U14800 (N_14800,N_12553,N_12262);
or U14801 (N_14801,N_13046,N_13720);
and U14802 (N_14802,N_12283,N_13620);
nor U14803 (N_14803,N_12388,N_13905);
xnor U14804 (N_14804,N_12445,N_12533);
nor U14805 (N_14805,N_13529,N_13340);
and U14806 (N_14806,N_13283,N_12847);
xnor U14807 (N_14807,N_13821,N_12869);
xnor U14808 (N_14808,N_13393,N_12699);
xor U14809 (N_14809,N_12032,N_12570);
or U14810 (N_14810,N_13493,N_12601);
nand U14811 (N_14811,N_13353,N_12354);
xnor U14812 (N_14812,N_12352,N_12881);
or U14813 (N_14813,N_12162,N_13413);
nor U14814 (N_14814,N_12921,N_13451);
nor U14815 (N_14815,N_13392,N_12841);
or U14816 (N_14816,N_12618,N_13289);
nor U14817 (N_14817,N_12506,N_12957);
nor U14818 (N_14818,N_13902,N_12815);
xnor U14819 (N_14819,N_13592,N_12811);
xnor U14820 (N_14820,N_13142,N_13824);
or U14821 (N_14821,N_12871,N_13232);
xnor U14822 (N_14822,N_12867,N_12566);
nand U14823 (N_14823,N_12011,N_13547);
and U14824 (N_14824,N_13435,N_12859);
nand U14825 (N_14825,N_12827,N_13070);
or U14826 (N_14826,N_12438,N_12594);
or U14827 (N_14827,N_12668,N_12952);
or U14828 (N_14828,N_13428,N_13222);
xnor U14829 (N_14829,N_13343,N_12915);
or U14830 (N_14830,N_13617,N_13782);
nand U14831 (N_14831,N_12170,N_13948);
nor U14832 (N_14832,N_13321,N_13141);
or U14833 (N_14833,N_12715,N_13097);
nand U14834 (N_14834,N_12365,N_12016);
and U14835 (N_14835,N_12840,N_13426);
nor U14836 (N_14836,N_12686,N_13602);
or U14837 (N_14837,N_12039,N_12724);
or U14838 (N_14838,N_12642,N_12193);
nor U14839 (N_14839,N_13228,N_13936);
and U14840 (N_14840,N_12428,N_13891);
xor U14841 (N_14841,N_13694,N_12446);
xor U14842 (N_14842,N_13558,N_13160);
nand U14843 (N_14843,N_12390,N_13476);
nor U14844 (N_14844,N_12343,N_12763);
xor U14845 (N_14845,N_12372,N_13723);
and U14846 (N_14846,N_12167,N_13021);
xnor U14847 (N_14847,N_12202,N_12832);
or U14848 (N_14848,N_12413,N_13218);
or U14849 (N_14849,N_12558,N_12363);
xnor U14850 (N_14850,N_13452,N_13442);
and U14851 (N_14851,N_12897,N_12149);
nor U14852 (N_14852,N_12275,N_13618);
nand U14853 (N_14853,N_13987,N_12923);
xor U14854 (N_14854,N_12077,N_13819);
xnor U14855 (N_14855,N_13879,N_12687);
nand U14856 (N_14856,N_13013,N_13571);
or U14857 (N_14857,N_12350,N_12311);
xnor U14858 (N_14858,N_13958,N_12123);
nor U14859 (N_14859,N_12845,N_12713);
xor U14860 (N_14860,N_12360,N_13211);
or U14861 (N_14861,N_13001,N_12778);
nor U14862 (N_14862,N_12680,N_12314);
and U14863 (N_14863,N_12416,N_12367);
and U14864 (N_14864,N_13387,N_12279);
and U14865 (N_14865,N_12142,N_12393);
nand U14866 (N_14866,N_12865,N_13175);
and U14867 (N_14867,N_13665,N_12237);
and U14868 (N_14868,N_12937,N_12814);
and U14869 (N_14869,N_12839,N_12540);
xor U14870 (N_14870,N_13587,N_12005);
nor U14871 (N_14871,N_13698,N_12470);
and U14872 (N_14872,N_13588,N_12502);
xor U14873 (N_14873,N_12564,N_12145);
xor U14874 (N_14874,N_12688,N_13573);
and U14875 (N_14875,N_13132,N_12858);
and U14876 (N_14876,N_13040,N_12554);
nand U14877 (N_14877,N_13880,N_13740);
and U14878 (N_14878,N_12001,N_13818);
and U14879 (N_14879,N_12043,N_12477);
and U14880 (N_14880,N_13838,N_13580);
nand U14881 (N_14881,N_13146,N_12491);
and U14882 (N_14882,N_13932,N_13906);
nand U14883 (N_14883,N_13686,N_12904);
xnor U14884 (N_14884,N_13181,N_13331);
and U14885 (N_14885,N_12826,N_12480);
or U14886 (N_14886,N_13949,N_13209);
nor U14887 (N_14887,N_13710,N_12743);
and U14888 (N_14888,N_12013,N_13814);
and U14889 (N_14889,N_12654,N_12722);
xor U14890 (N_14890,N_13202,N_13403);
and U14891 (N_14891,N_12135,N_13530);
and U14892 (N_14892,N_13191,N_12990);
nor U14893 (N_14893,N_13419,N_12002);
nand U14894 (N_14894,N_12634,N_13647);
and U14895 (N_14895,N_12981,N_12174);
nor U14896 (N_14896,N_13998,N_13745);
or U14897 (N_14897,N_12075,N_12539);
or U14898 (N_14898,N_13398,N_13882);
nand U14899 (N_14899,N_12973,N_13742);
xor U14900 (N_14900,N_13572,N_13256);
or U14901 (N_14901,N_13388,N_13696);
or U14902 (N_14902,N_13473,N_12659);
or U14903 (N_14903,N_12738,N_13194);
or U14904 (N_14904,N_12626,N_12598);
or U14905 (N_14905,N_13069,N_13513);
and U14906 (N_14906,N_13239,N_12960);
or U14907 (N_14907,N_12893,N_12676);
or U14908 (N_14908,N_13989,N_12218);
and U14909 (N_14909,N_12551,N_12735);
xor U14910 (N_14910,N_13708,N_12058);
nand U14911 (N_14911,N_13777,N_13829);
nand U14912 (N_14912,N_13303,N_12000);
xor U14913 (N_14913,N_13445,N_12774);
nand U14914 (N_14914,N_13667,N_12184);
nand U14915 (N_14915,N_12605,N_13022);
nand U14916 (N_14916,N_12809,N_13631);
nand U14917 (N_14917,N_13308,N_12933);
or U14918 (N_14918,N_12243,N_12266);
nand U14919 (N_14919,N_13612,N_13506);
or U14920 (N_14920,N_13050,N_13923);
nor U14921 (N_14921,N_13277,N_12948);
xor U14922 (N_14922,N_12197,N_12282);
xnor U14923 (N_14923,N_13234,N_13646);
nor U14924 (N_14924,N_13848,N_13866);
and U14925 (N_14925,N_13115,N_13820);
or U14926 (N_14926,N_12630,N_12302);
nand U14927 (N_14927,N_12042,N_13794);
nand U14928 (N_14928,N_12264,N_12754);
and U14929 (N_14929,N_12009,N_13916);
nor U14930 (N_14930,N_13792,N_13952);
and U14931 (N_14931,N_12177,N_13901);
nand U14932 (N_14932,N_12458,N_12421);
and U14933 (N_14933,N_12229,N_13379);
nand U14934 (N_14934,N_13524,N_13535);
and U14935 (N_14935,N_12108,N_13688);
or U14936 (N_14936,N_12336,N_13235);
and U14937 (N_14937,N_13674,N_12267);
or U14938 (N_14938,N_13834,N_12786);
and U14939 (N_14939,N_12604,N_12337);
and U14940 (N_14940,N_13324,N_12259);
xor U14941 (N_14941,N_13198,N_13370);
nand U14942 (N_14942,N_12836,N_12468);
and U14943 (N_14943,N_12939,N_13336);
or U14944 (N_14944,N_13197,N_12255);
or U14945 (N_14945,N_13967,N_13107);
or U14946 (N_14946,N_13929,N_13072);
nor U14947 (N_14947,N_12861,N_13036);
nand U14948 (N_14948,N_12608,N_13085);
and U14949 (N_14949,N_12082,N_13871);
nand U14950 (N_14950,N_12518,N_13685);
xor U14951 (N_14951,N_13284,N_12590);
and U14952 (N_14952,N_12092,N_13772);
or U14953 (N_14953,N_12340,N_13527);
nand U14954 (N_14954,N_12040,N_13890);
and U14955 (N_14955,N_12027,N_13053);
xnor U14956 (N_14956,N_13727,N_13101);
or U14957 (N_14957,N_12574,N_13295);
nor U14958 (N_14958,N_12228,N_12020);
or U14959 (N_14959,N_13098,N_12500);
and U14960 (N_14960,N_13457,N_12636);
xnor U14961 (N_14961,N_12031,N_13137);
and U14962 (N_14962,N_13768,N_12323);
or U14963 (N_14963,N_12924,N_13497);
nor U14964 (N_14964,N_12251,N_12316);
and U14965 (N_14965,N_13420,N_13762);
xor U14966 (N_14966,N_12109,N_13418);
nor U14967 (N_14967,N_12231,N_13268);
or U14968 (N_14968,N_13787,N_12051);
or U14969 (N_14969,N_13651,N_12465);
or U14970 (N_14970,N_13855,N_13042);
or U14971 (N_14971,N_13576,N_12892);
nor U14972 (N_14972,N_12965,N_12085);
and U14973 (N_14973,N_12411,N_13732);
or U14974 (N_14974,N_13624,N_12907);
nand U14975 (N_14975,N_12751,N_12498);
nand U14976 (N_14976,N_13369,N_13641);
xor U14977 (N_14977,N_13874,N_13845);
and U14978 (N_14978,N_13750,N_12469);
xor U14979 (N_14979,N_13433,N_13404);
xnor U14980 (N_14980,N_13739,N_12481);
or U14981 (N_14981,N_12298,N_13034);
nor U14982 (N_14982,N_13342,N_13307);
or U14983 (N_14983,N_13791,N_13296);
xnor U14984 (N_14984,N_12504,N_13545);
xnor U14985 (N_14985,N_13375,N_13163);
xnor U14986 (N_14986,N_12592,N_12967);
or U14987 (N_14987,N_12669,N_12802);
nand U14988 (N_14988,N_12226,N_13749);
or U14989 (N_14989,N_13123,N_12358);
nor U14990 (N_14990,N_12199,N_12984);
or U14991 (N_14991,N_12542,N_13312);
or U14992 (N_14992,N_13731,N_13582);
or U14993 (N_14993,N_13926,N_13758);
nand U14994 (N_14994,N_13850,N_13210);
nand U14995 (N_14995,N_13212,N_12692);
and U14996 (N_14996,N_12436,N_12672);
or U14997 (N_14997,N_13986,N_13802);
nor U14998 (N_14998,N_12632,N_13559);
and U14999 (N_14999,N_13368,N_12572);
nor U15000 (N_15000,N_13952,N_13527);
and U15001 (N_15001,N_13227,N_13124);
nor U15002 (N_15002,N_13279,N_13594);
and U15003 (N_15003,N_13038,N_12858);
nand U15004 (N_15004,N_13951,N_13661);
xor U15005 (N_15005,N_12852,N_12617);
nand U15006 (N_15006,N_12526,N_13616);
nand U15007 (N_15007,N_13036,N_12411);
nor U15008 (N_15008,N_13912,N_13114);
or U15009 (N_15009,N_13889,N_12419);
and U15010 (N_15010,N_12388,N_12112);
or U15011 (N_15011,N_13287,N_13484);
nor U15012 (N_15012,N_13249,N_12218);
and U15013 (N_15013,N_12817,N_12101);
and U15014 (N_15014,N_13087,N_13787);
or U15015 (N_15015,N_12319,N_12398);
and U15016 (N_15016,N_13726,N_13442);
nor U15017 (N_15017,N_13405,N_12138);
or U15018 (N_15018,N_13756,N_13335);
or U15019 (N_15019,N_12140,N_12423);
nor U15020 (N_15020,N_13333,N_12256);
xor U15021 (N_15021,N_12942,N_13324);
nand U15022 (N_15022,N_12249,N_12362);
and U15023 (N_15023,N_13050,N_13052);
or U15024 (N_15024,N_13042,N_13833);
nand U15025 (N_15025,N_12011,N_12485);
nor U15026 (N_15026,N_12381,N_13063);
nand U15027 (N_15027,N_12093,N_13186);
nand U15028 (N_15028,N_12993,N_12299);
or U15029 (N_15029,N_13766,N_12135);
xor U15030 (N_15030,N_12716,N_13658);
nor U15031 (N_15031,N_13556,N_13300);
and U15032 (N_15032,N_12985,N_12743);
and U15033 (N_15033,N_12547,N_12656);
xnor U15034 (N_15034,N_12884,N_12607);
nand U15035 (N_15035,N_12284,N_13926);
or U15036 (N_15036,N_13541,N_12576);
and U15037 (N_15037,N_13977,N_13401);
xor U15038 (N_15038,N_12062,N_12181);
xor U15039 (N_15039,N_12662,N_12946);
or U15040 (N_15040,N_12399,N_13349);
xor U15041 (N_15041,N_13873,N_12016);
and U15042 (N_15042,N_12164,N_12947);
or U15043 (N_15043,N_13252,N_12048);
nor U15044 (N_15044,N_13451,N_13122);
xor U15045 (N_15045,N_13147,N_13894);
nor U15046 (N_15046,N_12666,N_12926);
xor U15047 (N_15047,N_12198,N_12284);
and U15048 (N_15048,N_13944,N_13283);
nor U15049 (N_15049,N_13935,N_12648);
xnor U15050 (N_15050,N_12675,N_12660);
or U15051 (N_15051,N_13729,N_12802);
nand U15052 (N_15052,N_12832,N_12050);
or U15053 (N_15053,N_13255,N_12004);
nor U15054 (N_15054,N_13753,N_13294);
xor U15055 (N_15055,N_13226,N_13972);
or U15056 (N_15056,N_12899,N_12076);
and U15057 (N_15057,N_12534,N_12929);
and U15058 (N_15058,N_13256,N_12219);
nor U15059 (N_15059,N_12586,N_13727);
nor U15060 (N_15060,N_12848,N_13556);
or U15061 (N_15061,N_13168,N_12784);
xor U15062 (N_15062,N_13269,N_12548);
and U15063 (N_15063,N_12433,N_13619);
nor U15064 (N_15064,N_13386,N_12377);
or U15065 (N_15065,N_12709,N_13002);
and U15066 (N_15066,N_13182,N_12512);
or U15067 (N_15067,N_12857,N_12253);
nor U15068 (N_15068,N_13879,N_13486);
nor U15069 (N_15069,N_12030,N_13368);
or U15070 (N_15070,N_13970,N_12812);
and U15071 (N_15071,N_13829,N_12656);
or U15072 (N_15072,N_12073,N_13059);
and U15073 (N_15073,N_13471,N_12796);
or U15074 (N_15074,N_13890,N_12907);
and U15075 (N_15075,N_12436,N_12332);
and U15076 (N_15076,N_12436,N_13501);
nand U15077 (N_15077,N_13672,N_13788);
nor U15078 (N_15078,N_12559,N_12968);
or U15079 (N_15079,N_13914,N_13417);
nand U15080 (N_15080,N_13726,N_12400);
nand U15081 (N_15081,N_13442,N_13780);
and U15082 (N_15082,N_13399,N_12059);
and U15083 (N_15083,N_12014,N_12125);
or U15084 (N_15084,N_12015,N_12089);
nand U15085 (N_15085,N_12504,N_13453);
xor U15086 (N_15086,N_12236,N_13215);
nor U15087 (N_15087,N_13894,N_12809);
nor U15088 (N_15088,N_12233,N_12839);
or U15089 (N_15089,N_13060,N_12219);
xor U15090 (N_15090,N_13717,N_13302);
nand U15091 (N_15091,N_12713,N_12908);
xnor U15092 (N_15092,N_12610,N_13093);
nand U15093 (N_15093,N_13106,N_13338);
nand U15094 (N_15094,N_12648,N_12750);
xnor U15095 (N_15095,N_12352,N_12758);
xnor U15096 (N_15096,N_13824,N_13534);
or U15097 (N_15097,N_13458,N_12670);
and U15098 (N_15098,N_12905,N_12061);
xor U15099 (N_15099,N_12528,N_13906);
nand U15100 (N_15100,N_12991,N_13982);
and U15101 (N_15101,N_13301,N_13603);
nand U15102 (N_15102,N_12350,N_13298);
and U15103 (N_15103,N_12222,N_12743);
or U15104 (N_15104,N_13640,N_12839);
nand U15105 (N_15105,N_13814,N_12667);
xnor U15106 (N_15106,N_12906,N_13891);
nor U15107 (N_15107,N_12779,N_13287);
or U15108 (N_15108,N_12208,N_13173);
and U15109 (N_15109,N_13157,N_13560);
nand U15110 (N_15110,N_13565,N_12866);
and U15111 (N_15111,N_13802,N_13555);
or U15112 (N_15112,N_12886,N_12581);
or U15113 (N_15113,N_13389,N_12583);
or U15114 (N_15114,N_12150,N_13633);
xor U15115 (N_15115,N_12702,N_13003);
or U15116 (N_15116,N_12037,N_13187);
or U15117 (N_15117,N_12560,N_13138);
xnor U15118 (N_15118,N_13522,N_12077);
nand U15119 (N_15119,N_12678,N_13309);
or U15120 (N_15120,N_13122,N_13073);
nor U15121 (N_15121,N_13027,N_12586);
and U15122 (N_15122,N_12729,N_12399);
nand U15123 (N_15123,N_12812,N_12292);
nor U15124 (N_15124,N_13912,N_13880);
or U15125 (N_15125,N_13601,N_12030);
nor U15126 (N_15126,N_12017,N_13871);
nor U15127 (N_15127,N_12572,N_12078);
xnor U15128 (N_15128,N_12440,N_13670);
xnor U15129 (N_15129,N_13811,N_13724);
nor U15130 (N_15130,N_12196,N_12992);
or U15131 (N_15131,N_13613,N_13296);
nor U15132 (N_15132,N_12541,N_12858);
nor U15133 (N_15133,N_13007,N_12071);
nand U15134 (N_15134,N_13844,N_12528);
and U15135 (N_15135,N_12692,N_13064);
xnor U15136 (N_15136,N_13729,N_13519);
nor U15137 (N_15137,N_13962,N_12478);
nor U15138 (N_15138,N_13931,N_12719);
xor U15139 (N_15139,N_12340,N_13110);
and U15140 (N_15140,N_12772,N_12371);
xor U15141 (N_15141,N_13596,N_13974);
or U15142 (N_15142,N_13193,N_12962);
and U15143 (N_15143,N_13466,N_13557);
nand U15144 (N_15144,N_13049,N_12896);
nand U15145 (N_15145,N_13578,N_12493);
and U15146 (N_15146,N_12769,N_13501);
nor U15147 (N_15147,N_12500,N_12933);
or U15148 (N_15148,N_13320,N_13458);
and U15149 (N_15149,N_12391,N_13939);
and U15150 (N_15150,N_13292,N_12932);
nor U15151 (N_15151,N_13487,N_12077);
or U15152 (N_15152,N_13798,N_12702);
nor U15153 (N_15153,N_13621,N_13157);
or U15154 (N_15154,N_12355,N_12516);
nor U15155 (N_15155,N_12879,N_13942);
or U15156 (N_15156,N_13227,N_13995);
nor U15157 (N_15157,N_13094,N_13848);
and U15158 (N_15158,N_12186,N_12590);
and U15159 (N_15159,N_12168,N_12426);
nor U15160 (N_15160,N_12482,N_13830);
and U15161 (N_15161,N_13359,N_12403);
nor U15162 (N_15162,N_13437,N_12351);
nand U15163 (N_15163,N_12963,N_12838);
and U15164 (N_15164,N_13625,N_13107);
nand U15165 (N_15165,N_13323,N_12216);
or U15166 (N_15166,N_12563,N_12472);
and U15167 (N_15167,N_12775,N_12598);
nor U15168 (N_15168,N_12066,N_13644);
xor U15169 (N_15169,N_12855,N_12547);
or U15170 (N_15170,N_12670,N_13217);
nor U15171 (N_15171,N_13905,N_13916);
and U15172 (N_15172,N_13668,N_12478);
or U15173 (N_15173,N_12938,N_12254);
or U15174 (N_15174,N_13787,N_13567);
nand U15175 (N_15175,N_12904,N_13426);
nand U15176 (N_15176,N_13390,N_12130);
or U15177 (N_15177,N_13238,N_13917);
or U15178 (N_15178,N_12910,N_12739);
xnor U15179 (N_15179,N_12497,N_12484);
xor U15180 (N_15180,N_13296,N_12252);
and U15181 (N_15181,N_12636,N_13185);
nand U15182 (N_15182,N_12839,N_13918);
or U15183 (N_15183,N_12198,N_12139);
nand U15184 (N_15184,N_12549,N_13926);
and U15185 (N_15185,N_12633,N_12836);
nand U15186 (N_15186,N_12705,N_13269);
nor U15187 (N_15187,N_13992,N_12048);
and U15188 (N_15188,N_12609,N_12884);
and U15189 (N_15189,N_12998,N_13099);
nor U15190 (N_15190,N_13732,N_13203);
or U15191 (N_15191,N_13567,N_13721);
nand U15192 (N_15192,N_12179,N_12365);
and U15193 (N_15193,N_12625,N_13711);
nand U15194 (N_15194,N_13423,N_13363);
nor U15195 (N_15195,N_13849,N_12172);
and U15196 (N_15196,N_12367,N_13428);
nor U15197 (N_15197,N_12730,N_13083);
nand U15198 (N_15198,N_12345,N_12614);
nand U15199 (N_15199,N_13881,N_12626);
and U15200 (N_15200,N_12463,N_13601);
nor U15201 (N_15201,N_12573,N_12687);
or U15202 (N_15202,N_13121,N_12165);
and U15203 (N_15203,N_12924,N_12405);
or U15204 (N_15204,N_12234,N_13482);
and U15205 (N_15205,N_12634,N_13297);
nor U15206 (N_15206,N_12139,N_13119);
or U15207 (N_15207,N_12114,N_13038);
nor U15208 (N_15208,N_12007,N_12141);
and U15209 (N_15209,N_12590,N_12455);
or U15210 (N_15210,N_12099,N_13268);
nor U15211 (N_15211,N_12485,N_12847);
or U15212 (N_15212,N_12661,N_12847);
and U15213 (N_15213,N_12274,N_13045);
and U15214 (N_15214,N_12470,N_12598);
and U15215 (N_15215,N_13809,N_12162);
and U15216 (N_15216,N_12214,N_13979);
nand U15217 (N_15217,N_12133,N_12903);
and U15218 (N_15218,N_13470,N_12878);
xor U15219 (N_15219,N_12614,N_13583);
nand U15220 (N_15220,N_12036,N_12932);
xnor U15221 (N_15221,N_13153,N_13996);
xnor U15222 (N_15222,N_12266,N_13961);
xor U15223 (N_15223,N_12055,N_13540);
nand U15224 (N_15224,N_13530,N_12375);
or U15225 (N_15225,N_12002,N_12007);
and U15226 (N_15226,N_13348,N_12986);
or U15227 (N_15227,N_13954,N_13306);
nand U15228 (N_15228,N_12274,N_12130);
nor U15229 (N_15229,N_12792,N_13013);
nor U15230 (N_15230,N_13146,N_13378);
nand U15231 (N_15231,N_13720,N_13871);
and U15232 (N_15232,N_12576,N_13762);
or U15233 (N_15233,N_12579,N_12755);
nand U15234 (N_15234,N_13441,N_13001);
xor U15235 (N_15235,N_13491,N_12327);
and U15236 (N_15236,N_12274,N_13903);
xnor U15237 (N_15237,N_13475,N_13389);
nor U15238 (N_15238,N_12546,N_12808);
nand U15239 (N_15239,N_13019,N_13528);
and U15240 (N_15240,N_12117,N_13350);
and U15241 (N_15241,N_12284,N_12234);
or U15242 (N_15242,N_13210,N_13019);
or U15243 (N_15243,N_12475,N_13075);
and U15244 (N_15244,N_13046,N_13765);
nand U15245 (N_15245,N_13843,N_13568);
xnor U15246 (N_15246,N_13509,N_12618);
and U15247 (N_15247,N_13521,N_12867);
nand U15248 (N_15248,N_13813,N_12170);
xnor U15249 (N_15249,N_12143,N_13314);
nand U15250 (N_15250,N_12237,N_13524);
nand U15251 (N_15251,N_12616,N_12787);
nor U15252 (N_15252,N_13527,N_12985);
and U15253 (N_15253,N_12361,N_12198);
xnor U15254 (N_15254,N_12783,N_12152);
xor U15255 (N_15255,N_13296,N_13483);
xnor U15256 (N_15256,N_12870,N_13151);
and U15257 (N_15257,N_12093,N_13885);
xor U15258 (N_15258,N_13153,N_13607);
xor U15259 (N_15259,N_13536,N_13617);
and U15260 (N_15260,N_12222,N_13987);
xnor U15261 (N_15261,N_13490,N_12341);
nor U15262 (N_15262,N_12026,N_12704);
or U15263 (N_15263,N_13159,N_13686);
nand U15264 (N_15264,N_13370,N_12662);
xor U15265 (N_15265,N_13074,N_13557);
nor U15266 (N_15266,N_12392,N_13722);
nand U15267 (N_15267,N_13715,N_12515);
and U15268 (N_15268,N_13671,N_13830);
or U15269 (N_15269,N_12380,N_13765);
nand U15270 (N_15270,N_12338,N_12587);
nor U15271 (N_15271,N_13469,N_13692);
or U15272 (N_15272,N_12594,N_13509);
and U15273 (N_15273,N_12633,N_12950);
nor U15274 (N_15274,N_13148,N_12627);
nor U15275 (N_15275,N_13941,N_12025);
xor U15276 (N_15276,N_12458,N_12797);
xor U15277 (N_15277,N_12159,N_13002);
nand U15278 (N_15278,N_13325,N_13037);
nor U15279 (N_15279,N_12835,N_12936);
xnor U15280 (N_15280,N_12159,N_13942);
nor U15281 (N_15281,N_12785,N_12584);
nor U15282 (N_15282,N_12728,N_12621);
and U15283 (N_15283,N_12165,N_12791);
and U15284 (N_15284,N_12562,N_12087);
nand U15285 (N_15285,N_13153,N_12763);
nand U15286 (N_15286,N_13063,N_13231);
or U15287 (N_15287,N_12469,N_12519);
nand U15288 (N_15288,N_12757,N_12571);
nor U15289 (N_15289,N_13434,N_13570);
nor U15290 (N_15290,N_12833,N_12845);
xnor U15291 (N_15291,N_13323,N_13484);
nand U15292 (N_15292,N_12176,N_12428);
xnor U15293 (N_15293,N_12793,N_13931);
nor U15294 (N_15294,N_12683,N_12617);
nand U15295 (N_15295,N_12200,N_13773);
nor U15296 (N_15296,N_13601,N_12773);
or U15297 (N_15297,N_12593,N_13376);
nor U15298 (N_15298,N_13280,N_13129);
nand U15299 (N_15299,N_12577,N_13562);
or U15300 (N_15300,N_13675,N_12706);
and U15301 (N_15301,N_13867,N_12746);
nand U15302 (N_15302,N_13778,N_13783);
nor U15303 (N_15303,N_12357,N_13075);
or U15304 (N_15304,N_12989,N_13109);
or U15305 (N_15305,N_12201,N_13945);
and U15306 (N_15306,N_12012,N_12860);
nand U15307 (N_15307,N_13277,N_13051);
xor U15308 (N_15308,N_12973,N_12199);
xnor U15309 (N_15309,N_13623,N_13655);
nor U15310 (N_15310,N_13077,N_12184);
nand U15311 (N_15311,N_13306,N_13703);
nand U15312 (N_15312,N_13805,N_12100);
xor U15313 (N_15313,N_13295,N_12247);
or U15314 (N_15314,N_13454,N_12047);
or U15315 (N_15315,N_12606,N_13014);
nand U15316 (N_15316,N_13430,N_13904);
nand U15317 (N_15317,N_12319,N_13836);
xnor U15318 (N_15318,N_12203,N_12956);
nand U15319 (N_15319,N_12187,N_13973);
and U15320 (N_15320,N_13247,N_13682);
nand U15321 (N_15321,N_12472,N_12860);
or U15322 (N_15322,N_12688,N_13961);
and U15323 (N_15323,N_13500,N_13141);
nand U15324 (N_15324,N_12443,N_12942);
nand U15325 (N_15325,N_12488,N_13031);
or U15326 (N_15326,N_12704,N_12730);
nand U15327 (N_15327,N_12405,N_12016);
nand U15328 (N_15328,N_12903,N_13604);
nand U15329 (N_15329,N_13155,N_13538);
xor U15330 (N_15330,N_12841,N_13836);
or U15331 (N_15331,N_13015,N_12005);
or U15332 (N_15332,N_12111,N_12935);
nor U15333 (N_15333,N_12093,N_12990);
xor U15334 (N_15334,N_13325,N_13824);
nand U15335 (N_15335,N_12442,N_12014);
nand U15336 (N_15336,N_13833,N_12233);
and U15337 (N_15337,N_13195,N_13476);
and U15338 (N_15338,N_13209,N_13765);
or U15339 (N_15339,N_13682,N_12065);
or U15340 (N_15340,N_13007,N_12648);
and U15341 (N_15341,N_12589,N_13267);
or U15342 (N_15342,N_13322,N_13102);
xnor U15343 (N_15343,N_12389,N_13834);
or U15344 (N_15344,N_13794,N_13701);
or U15345 (N_15345,N_12577,N_13615);
and U15346 (N_15346,N_12805,N_13092);
nor U15347 (N_15347,N_13047,N_13210);
or U15348 (N_15348,N_13992,N_12709);
nand U15349 (N_15349,N_13744,N_12027);
and U15350 (N_15350,N_12410,N_12575);
and U15351 (N_15351,N_12245,N_13898);
and U15352 (N_15352,N_12151,N_12496);
and U15353 (N_15353,N_13559,N_13910);
and U15354 (N_15354,N_13122,N_13859);
nor U15355 (N_15355,N_12347,N_13971);
and U15356 (N_15356,N_12752,N_12872);
nand U15357 (N_15357,N_12072,N_12584);
or U15358 (N_15358,N_13937,N_12906);
nor U15359 (N_15359,N_13917,N_12709);
or U15360 (N_15360,N_13368,N_12638);
nand U15361 (N_15361,N_13214,N_13197);
nand U15362 (N_15362,N_13845,N_12792);
or U15363 (N_15363,N_12175,N_12401);
nor U15364 (N_15364,N_13200,N_13775);
or U15365 (N_15365,N_12438,N_12644);
xnor U15366 (N_15366,N_12230,N_12218);
and U15367 (N_15367,N_12906,N_12737);
xor U15368 (N_15368,N_12798,N_12212);
xnor U15369 (N_15369,N_13647,N_12022);
and U15370 (N_15370,N_13668,N_12031);
or U15371 (N_15371,N_12967,N_13453);
or U15372 (N_15372,N_12657,N_12074);
xor U15373 (N_15373,N_12356,N_12786);
xor U15374 (N_15374,N_13530,N_12559);
and U15375 (N_15375,N_12136,N_13772);
or U15376 (N_15376,N_13211,N_12362);
nor U15377 (N_15377,N_12820,N_13614);
or U15378 (N_15378,N_13366,N_12616);
or U15379 (N_15379,N_13539,N_12079);
xnor U15380 (N_15380,N_13340,N_13406);
and U15381 (N_15381,N_12108,N_12484);
nor U15382 (N_15382,N_13307,N_12834);
xnor U15383 (N_15383,N_12251,N_13569);
nor U15384 (N_15384,N_12499,N_13492);
xor U15385 (N_15385,N_13932,N_13701);
nand U15386 (N_15386,N_13563,N_13337);
and U15387 (N_15387,N_12038,N_13794);
nor U15388 (N_15388,N_13801,N_13456);
nand U15389 (N_15389,N_12081,N_12002);
xor U15390 (N_15390,N_12641,N_12079);
nor U15391 (N_15391,N_13580,N_12200);
and U15392 (N_15392,N_13968,N_13301);
nand U15393 (N_15393,N_12193,N_13710);
nand U15394 (N_15394,N_12619,N_13717);
xnor U15395 (N_15395,N_13508,N_12523);
nor U15396 (N_15396,N_12679,N_12741);
nand U15397 (N_15397,N_13137,N_12737);
xnor U15398 (N_15398,N_13536,N_13183);
and U15399 (N_15399,N_13824,N_12071);
nor U15400 (N_15400,N_13968,N_13411);
or U15401 (N_15401,N_12322,N_12362);
nand U15402 (N_15402,N_12336,N_13890);
or U15403 (N_15403,N_13457,N_13815);
nor U15404 (N_15404,N_13227,N_13940);
or U15405 (N_15405,N_13152,N_13806);
and U15406 (N_15406,N_12949,N_12236);
or U15407 (N_15407,N_13655,N_12783);
nand U15408 (N_15408,N_13302,N_13053);
nor U15409 (N_15409,N_12390,N_13918);
or U15410 (N_15410,N_12389,N_12129);
and U15411 (N_15411,N_13235,N_13412);
xor U15412 (N_15412,N_12790,N_12897);
and U15413 (N_15413,N_12371,N_12110);
or U15414 (N_15414,N_13493,N_13989);
nor U15415 (N_15415,N_13401,N_13345);
nand U15416 (N_15416,N_12968,N_12369);
nor U15417 (N_15417,N_13546,N_12503);
and U15418 (N_15418,N_12129,N_12225);
nand U15419 (N_15419,N_12448,N_13484);
nor U15420 (N_15420,N_13630,N_12015);
nand U15421 (N_15421,N_12672,N_13917);
or U15422 (N_15422,N_12836,N_13888);
xor U15423 (N_15423,N_12480,N_13165);
nor U15424 (N_15424,N_12582,N_13283);
or U15425 (N_15425,N_13999,N_12686);
nor U15426 (N_15426,N_13999,N_12526);
nand U15427 (N_15427,N_13037,N_13176);
or U15428 (N_15428,N_12621,N_13724);
or U15429 (N_15429,N_12809,N_12808);
or U15430 (N_15430,N_13326,N_13854);
nand U15431 (N_15431,N_13441,N_12064);
or U15432 (N_15432,N_12264,N_13112);
nor U15433 (N_15433,N_12215,N_12177);
or U15434 (N_15434,N_12606,N_12776);
xor U15435 (N_15435,N_13170,N_12673);
and U15436 (N_15436,N_13829,N_12716);
xor U15437 (N_15437,N_12048,N_13066);
xnor U15438 (N_15438,N_12589,N_13716);
nor U15439 (N_15439,N_13332,N_12831);
nand U15440 (N_15440,N_12085,N_13358);
nor U15441 (N_15441,N_12978,N_12747);
xnor U15442 (N_15442,N_13479,N_12057);
nand U15443 (N_15443,N_13085,N_12766);
nand U15444 (N_15444,N_12731,N_12532);
nor U15445 (N_15445,N_13320,N_13197);
nor U15446 (N_15446,N_12177,N_13280);
and U15447 (N_15447,N_13904,N_13928);
nand U15448 (N_15448,N_13127,N_12605);
nand U15449 (N_15449,N_12856,N_12156);
or U15450 (N_15450,N_12052,N_13633);
nand U15451 (N_15451,N_12964,N_12334);
or U15452 (N_15452,N_12847,N_12727);
and U15453 (N_15453,N_12679,N_13337);
and U15454 (N_15454,N_13483,N_13545);
xnor U15455 (N_15455,N_12877,N_13411);
nand U15456 (N_15456,N_13874,N_12536);
or U15457 (N_15457,N_12939,N_13750);
xor U15458 (N_15458,N_13931,N_13934);
nand U15459 (N_15459,N_13746,N_12592);
xnor U15460 (N_15460,N_13068,N_13483);
nand U15461 (N_15461,N_12478,N_12088);
nor U15462 (N_15462,N_13572,N_13647);
xor U15463 (N_15463,N_13159,N_13584);
or U15464 (N_15464,N_13251,N_12814);
nor U15465 (N_15465,N_12360,N_13122);
or U15466 (N_15466,N_12614,N_12676);
nor U15467 (N_15467,N_12411,N_13681);
and U15468 (N_15468,N_13922,N_13689);
and U15469 (N_15469,N_13515,N_13679);
or U15470 (N_15470,N_13990,N_13800);
or U15471 (N_15471,N_13471,N_13575);
and U15472 (N_15472,N_13932,N_12878);
nor U15473 (N_15473,N_13814,N_13936);
nor U15474 (N_15474,N_13397,N_13043);
xor U15475 (N_15475,N_12425,N_13886);
or U15476 (N_15476,N_12141,N_13279);
nand U15477 (N_15477,N_12227,N_13270);
and U15478 (N_15478,N_12422,N_12714);
or U15479 (N_15479,N_13583,N_12272);
and U15480 (N_15480,N_13221,N_12189);
nand U15481 (N_15481,N_12184,N_12992);
and U15482 (N_15482,N_12118,N_13809);
or U15483 (N_15483,N_13120,N_12557);
or U15484 (N_15484,N_13275,N_13308);
nor U15485 (N_15485,N_12509,N_12043);
nand U15486 (N_15486,N_12326,N_13687);
nor U15487 (N_15487,N_12167,N_12955);
or U15488 (N_15488,N_13971,N_12022);
xor U15489 (N_15489,N_13341,N_13645);
xnor U15490 (N_15490,N_13898,N_12234);
xor U15491 (N_15491,N_12250,N_13018);
xnor U15492 (N_15492,N_13901,N_12774);
xnor U15493 (N_15493,N_12325,N_12546);
xor U15494 (N_15494,N_13654,N_13420);
xor U15495 (N_15495,N_12088,N_12683);
or U15496 (N_15496,N_13845,N_13233);
xor U15497 (N_15497,N_13598,N_13058);
xnor U15498 (N_15498,N_13796,N_12207);
or U15499 (N_15499,N_12683,N_13837);
or U15500 (N_15500,N_12170,N_13602);
xnor U15501 (N_15501,N_13173,N_13188);
and U15502 (N_15502,N_12262,N_12571);
or U15503 (N_15503,N_13483,N_13753);
nand U15504 (N_15504,N_13685,N_12311);
nand U15505 (N_15505,N_12017,N_12350);
or U15506 (N_15506,N_12829,N_13254);
nor U15507 (N_15507,N_12958,N_13378);
nor U15508 (N_15508,N_13168,N_12940);
xor U15509 (N_15509,N_13954,N_12360);
xor U15510 (N_15510,N_12511,N_13070);
xor U15511 (N_15511,N_12701,N_12718);
nor U15512 (N_15512,N_13043,N_13470);
nand U15513 (N_15513,N_12862,N_13809);
or U15514 (N_15514,N_13315,N_12894);
nor U15515 (N_15515,N_12957,N_12578);
and U15516 (N_15516,N_13658,N_12162);
and U15517 (N_15517,N_13921,N_12995);
or U15518 (N_15518,N_12110,N_13707);
or U15519 (N_15519,N_12810,N_13235);
or U15520 (N_15520,N_12272,N_13350);
nand U15521 (N_15521,N_13521,N_12779);
or U15522 (N_15522,N_13821,N_13269);
or U15523 (N_15523,N_12714,N_13569);
nand U15524 (N_15524,N_13130,N_12285);
xor U15525 (N_15525,N_12218,N_13807);
nor U15526 (N_15526,N_12135,N_12056);
nor U15527 (N_15527,N_12640,N_12654);
or U15528 (N_15528,N_13604,N_13040);
nor U15529 (N_15529,N_13124,N_12466);
xnor U15530 (N_15530,N_12696,N_12538);
nand U15531 (N_15531,N_12084,N_12954);
or U15532 (N_15532,N_13858,N_12293);
and U15533 (N_15533,N_13257,N_13973);
or U15534 (N_15534,N_13594,N_13754);
and U15535 (N_15535,N_12883,N_13057);
xnor U15536 (N_15536,N_12622,N_12231);
and U15537 (N_15537,N_13043,N_13536);
nor U15538 (N_15538,N_13530,N_12962);
nor U15539 (N_15539,N_13398,N_13985);
xor U15540 (N_15540,N_12161,N_13800);
or U15541 (N_15541,N_12301,N_12163);
or U15542 (N_15542,N_12406,N_12688);
or U15543 (N_15543,N_13194,N_12741);
or U15544 (N_15544,N_13064,N_12921);
and U15545 (N_15545,N_12431,N_13788);
or U15546 (N_15546,N_12787,N_12711);
nor U15547 (N_15547,N_12789,N_13955);
nor U15548 (N_15548,N_13901,N_13913);
xor U15549 (N_15549,N_13588,N_13781);
and U15550 (N_15550,N_12346,N_12717);
or U15551 (N_15551,N_13630,N_12693);
or U15552 (N_15552,N_13337,N_13889);
xor U15553 (N_15553,N_12489,N_12400);
nor U15554 (N_15554,N_12232,N_13816);
and U15555 (N_15555,N_12603,N_13913);
and U15556 (N_15556,N_13942,N_12856);
or U15557 (N_15557,N_13988,N_13964);
or U15558 (N_15558,N_13096,N_13956);
and U15559 (N_15559,N_12556,N_12243);
and U15560 (N_15560,N_13419,N_13564);
and U15561 (N_15561,N_13838,N_12776);
nor U15562 (N_15562,N_13786,N_13369);
xnor U15563 (N_15563,N_12962,N_12927);
or U15564 (N_15564,N_12392,N_13410);
nor U15565 (N_15565,N_12881,N_12436);
and U15566 (N_15566,N_12619,N_12188);
and U15567 (N_15567,N_12733,N_13845);
nand U15568 (N_15568,N_12348,N_13493);
and U15569 (N_15569,N_12285,N_13934);
nand U15570 (N_15570,N_12468,N_12098);
nand U15571 (N_15571,N_12255,N_13255);
xor U15572 (N_15572,N_13637,N_13054);
nor U15573 (N_15573,N_13010,N_12587);
nor U15574 (N_15574,N_13057,N_13007);
or U15575 (N_15575,N_12821,N_12610);
nand U15576 (N_15576,N_12567,N_12233);
or U15577 (N_15577,N_13590,N_13183);
or U15578 (N_15578,N_13841,N_12339);
and U15579 (N_15579,N_12302,N_12268);
nand U15580 (N_15580,N_12557,N_13357);
xor U15581 (N_15581,N_12736,N_12672);
nor U15582 (N_15582,N_12709,N_13658);
and U15583 (N_15583,N_12730,N_13878);
nand U15584 (N_15584,N_13571,N_13951);
and U15585 (N_15585,N_12902,N_13537);
xor U15586 (N_15586,N_12919,N_13152);
and U15587 (N_15587,N_13655,N_12416);
or U15588 (N_15588,N_12962,N_13257);
nand U15589 (N_15589,N_12113,N_13250);
xnor U15590 (N_15590,N_12165,N_13761);
xnor U15591 (N_15591,N_13387,N_13015);
or U15592 (N_15592,N_12806,N_12725);
nand U15593 (N_15593,N_12158,N_12416);
xnor U15594 (N_15594,N_12058,N_12406);
and U15595 (N_15595,N_13221,N_13864);
and U15596 (N_15596,N_13208,N_12308);
nand U15597 (N_15597,N_13265,N_12086);
or U15598 (N_15598,N_12580,N_13285);
nor U15599 (N_15599,N_12175,N_13136);
and U15600 (N_15600,N_13759,N_13527);
xnor U15601 (N_15601,N_13031,N_13658);
xor U15602 (N_15602,N_13684,N_12381);
nor U15603 (N_15603,N_13350,N_12950);
and U15604 (N_15604,N_12990,N_12132);
xor U15605 (N_15605,N_13394,N_12200);
xor U15606 (N_15606,N_12908,N_13287);
or U15607 (N_15607,N_12201,N_12583);
or U15608 (N_15608,N_12836,N_12948);
or U15609 (N_15609,N_12056,N_13270);
xor U15610 (N_15610,N_13938,N_12871);
nor U15611 (N_15611,N_12781,N_13871);
nand U15612 (N_15612,N_12348,N_12649);
nand U15613 (N_15613,N_12924,N_13051);
or U15614 (N_15614,N_13421,N_13429);
or U15615 (N_15615,N_13902,N_13036);
or U15616 (N_15616,N_13473,N_13889);
xor U15617 (N_15617,N_13273,N_12386);
or U15618 (N_15618,N_13106,N_12934);
and U15619 (N_15619,N_12597,N_13694);
xor U15620 (N_15620,N_13075,N_13204);
nor U15621 (N_15621,N_12426,N_12106);
and U15622 (N_15622,N_13816,N_13151);
nand U15623 (N_15623,N_13575,N_13704);
and U15624 (N_15624,N_12798,N_12173);
nand U15625 (N_15625,N_12255,N_13541);
and U15626 (N_15626,N_12448,N_12565);
xor U15627 (N_15627,N_13813,N_12567);
nand U15628 (N_15628,N_12714,N_13477);
nor U15629 (N_15629,N_13647,N_12452);
xnor U15630 (N_15630,N_12203,N_12614);
nor U15631 (N_15631,N_12439,N_12820);
nand U15632 (N_15632,N_12096,N_12996);
xor U15633 (N_15633,N_12517,N_12624);
and U15634 (N_15634,N_12202,N_13993);
nand U15635 (N_15635,N_13349,N_12817);
nor U15636 (N_15636,N_13631,N_12307);
xnor U15637 (N_15637,N_12132,N_13227);
and U15638 (N_15638,N_13284,N_13184);
and U15639 (N_15639,N_13341,N_12586);
nand U15640 (N_15640,N_13440,N_13085);
nor U15641 (N_15641,N_12705,N_12508);
and U15642 (N_15642,N_13232,N_13011);
nand U15643 (N_15643,N_13069,N_12912);
or U15644 (N_15644,N_13973,N_13343);
or U15645 (N_15645,N_12298,N_12693);
nand U15646 (N_15646,N_13612,N_13431);
or U15647 (N_15647,N_12072,N_12926);
xnor U15648 (N_15648,N_13020,N_13365);
nand U15649 (N_15649,N_12082,N_12130);
and U15650 (N_15650,N_13601,N_12920);
and U15651 (N_15651,N_12840,N_13544);
xor U15652 (N_15652,N_13811,N_13873);
xor U15653 (N_15653,N_13167,N_13243);
and U15654 (N_15654,N_12910,N_12973);
or U15655 (N_15655,N_12812,N_13093);
nand U15656 (N_15656,N_13600,N_13335);
nor U15657 (N_15657,N_13217,N_12140);
and U15658 (N_15658,N_12243,N_13785);
nor U15659 (N_15659,N_12757,N_12005);
nor U15660 (N_15660,N_12286,N_12857);
nand U15661 (N_15661,N_13209,N_13387);
nand U15662 (N_15662,N_12157,N_13676);
nand U15663 (N_15663,N_12007,N_13353);
or U15664 (N_15664,N_13408,N_12664);
nand U15665 (N_15665,N_12501,N_12742);
and U15666 (N_15666,N_12100,N_13227);
and U15667 (N_15667,N_12647,N_13376);
or U15668 (N_15668,N_12722,N_12894);
or U15669 (N_15669,N_13747,N_12619);
nand U15670 (N_15670,N_12812,N_13971);
or U15671 (N_15671,N_12258,N_13511);
or U15672 (N_15672,N_12005,N_12411);
and U15673 (N_15673,N_12075,N_12506);
or U15674 (N_15674,N_12782,N_12918);
nor U15675 (N_15675,N_12675,N_13490);
nand U15676 (N_15676,N_13946,N_13994);
nor U15677 (N_15677,N_13093,N_12553);
and U15678 (N_15678,N_12411,N_12178);
nand U15679 (N_15679,N_12811,N_13985);
and U15680 (N_15680,N_13161,N_13594);
nor U15681 (N_15681,N_12629,N_13171);
nand U15682 (N_15682,N_13278,N_13281);
nor U15683 (N_15683,N_13766,N_12203);
and U15684 (N_15684,N_12676,N_12345);
nand U15685 (N_15685,N_12485,N_13888);
or U15686 (N_15686,N_12783,N_12682);
or U15687 (N_15687,N_12367,N_12779);
xnor U15688 (N_15688,N_12463,N_13703);
xor U15689 (N_15689,N_13185,N_12162);
and U15690 (N_15690,N_12860,N_12572);
and U15691 (N_15691,N_12201,N_12774);
and U15692 (N_15692,N_13987,N_13531);
nor U15693 (N_15693,N_12805,N_12116);
and U15694 (N_15694,N_13994,N_13810);
nand U15695 (N_15695,N_12499,N_13493);
and U15696 (N_15696,N_13635,N_12424);
nor U15697 (N_15697,N_12919,N_12020);
or U15698 (N_15698,N_13380,N_13128);
or U15699 (N_15699,N_12288,N_13454);
or U15700 (N_15700,N_13567,N_12662);
xnor U15701 (N_15701,N_12483,N_12249);
nor U15702 (N_15702,N_12403,N_12234);
nand U15703 (N_15703,N_12659,N_13600);
nand U15704 (N_15704,N_12062,N_13763);
nor U15705 (N_15705,N_13789,N_12123);
xnor U15706 (N_15706,N_13258,N_13760);
nor U15707 (N_15707,N_13247,N_12900);
nand U15708 (N_15708,N_13576,N_12493);
nand U15709 (N_15709,N_13273,N_12196);
nor U15710 (N_15710,N_13285,N_12034);
nand U15711 (N_15711,N_13224,N_13301);
nor U15712 (N_15712,N_12285,N_13683);
xnor U15713 (N_15713,N_13159,N_13579);
or U15714 (N_15714,N_12331,N_13738);
xnor U15715 (N_15715,N_12663,N_13656);
nor U15716 (N_15716,N_12066,N_13449);
xnor U15717 (N_15717,N_13672,N_13372);
xnor U15718 (N_15718,N_13884,N_12737);
nor U15719 (N_15719,N_12480,N_13100);
nor U15720 (N_15720,N_12958,N_13780);
nor U15721 (N_15721,N_12106,N_13892);
or U15722 (N_15722,N_13191,N_13710);
nor U15723 (N_15723,N_12650,N_12187);
nand U15724 (N_15724,N_13404,N_13088);
nand U15725 (N_15725,N_12677,N_12658);
xnor U15726 (N_15726,N_13741,N_12101);
nand U15727 (N_15727,N_13752,N_13558);
nand U15728 (N_15728,N_13308,N_12067);
nor U15729 (N_15729,N_12930,N_13719);
nor U15730 (N_15730,N_12484,N_13796);
or U15731 (N_15731,N_12946,N_13081);
xor U15732 (N_15732,N_12428,N_13310);
nand U15733 (N_15733,N_12937,N_13242);
xnor U15734 (N_15734,N_13837,N_13210);
xnor U15735 (N_15735,N_13696,N_13975);
nand U15736 (N_15736,N_12215,N_13090);
nand U15737 (N_15737,N_13587,N_13772);
xnor U15738 (N_15738,N_13952,N_13700);
and U15739 (N_15739,N_13465,N_13573);
or U15740 (N_15740,N_12236,N_13386);
xnor U15741 (N_15741,N_13719,N_13607);
nand U15742 (N_15742,N_13133,N_12867);
nor U15743 (N_15743,N_12788,N_12297);
nand U15744 (N_15744,N_13946,N_12679);
and U15745 (N_15745,N_13860,N_12187);
nand U15746 (N_15746,N_12189,N_13270);
nor U15747 (N_15747,N_13098,N_13217);
nor U15748 (N_15748,N_12797,N_13170);
nor U15749 (N_15749,N_13556,N_12297);
nor U15750 (N_15750,N_13549,N_13657);
xnor U15751 (N_15751,N_12076,N_13866);
or U15752 (N_15752,N_12248,N_13859);
nand U15753 (N_15753,N_12478,N_12094);
xnor U15754 (N_15754,N_13770,N_12833);
or U15755 (N_15755,N_13496,N_13177);
nor U15756 (N_15756,N_13390,N_12258);
nand U15757 (N_15757,N_12173,N_12754);
nand U15758 (N_15758,N_13174,N_12909);
nand U15759 (N_15759,N_12088,N_13547);
xnor U15760 (N_15760,N_12345,N_12891);
nand U15761 (N_15761,N_13741,N_13652);
xnor U15762 (N_15762,N_12273,N_12386);
or U15763 (N_15763,N_12404,N_12582);
nand U15764 (N_15764,N_13213,N_13576);
xnor U15765 (N_15765,N_12819,N_13254);
and U15766 (N_15766,N_12085,N_13219);
or U15767 (N_15767,N_12507,N_12469);
or U15768 (N_15768,N_13813,N_13820);
or U15769 (N_15769,N_12330,N_12424);
and U15770 (N_15770,N_12494,N_13876);
and U15771 (N_15771,N_12182,N_12559);
nand U15772 (N_15772,N_12456,N_12169);
or U15773 (N_15773,N_13250,N_12102);
xor U15774 (N_15774,N_12618,N_12199);
nand U15775 (N_15775,N_12346,N_12799);
xnor U15776 (N_15776,N_12990,N_12874);
nand U15777 (N_15777,N_12371,N_13225);
and U15778 (N_15778,N_12890,N_12274);
nand U15779 (N_15779,N_12440,N_13521);
xor U15780 (N_15780,N_12739,N_13125);
nor U15781 (N_15781,N_12499,N_13462);
nand U15782 (N_15782,N_12067,N_13892);
and U15783 (N_15783,N_12250,N_13147);
nand U15784 (N_15784,N_13339,N_12365);
and U15785 (N_15785,N_13320,N_13420);
and U15786 (N_15786,N_12364,N_12409);
and U15787 (N_15787,N_12623,N_13779);
or U15788 (N_15788,N_12980,N_13429);
xnor U15789 (N_15789,N_12499,N_12741);
xor U15790 (N_15790,N_13660,N_12761);
nor U15791 (N_15791,N_13400,N_12672);
nor U15792 (N_15792,N_12566,N_13206);
xor U15793 (N_15793,N_13654,N_12741);
and U15794 (N_15794,N_13733,N_13739);
or U15795 (N_15795,N_12658,N_12780);
nor U15796 (N_15796,N_13017,N_12160);
and U15797 (N_15797,N_13942,N_13165);
or U15798 (N_15798,N_12797,N_13509);
or U15799 (N_15799,N_13446,N_13549);
and U15800 (N_15800,N_13528,N_13492);
xnor U15801 (N_15801,N_12575,N_12018);
nand U15802 (N_15802,N_13241,N_12318);
xnor U15803 (N_15803,N_13142,N_12445);
nand U15804 (N_15804,N_13859,N_12283);
or U15805 (N_15805,N_13889,N_12762);
or U15806 (N_15806,N_13139,N_12969);
xnor U15807 (N_15807,N_12560,N_13805);
nand U15808 (N_15808,N_13369,N_13567);
xor U15809 (N_15809,N_13122,N_12519);
nand U15810 (N_15810,N_13641,N_13181);
xnor U15811 (N_15811,N_13157,N_12231);
nor U15812 (N_15812,N_12190,N_12109);
nor U15813 (N_15813,N_12234,N_13006);
nor U15814 (N_15814,N_12480,N_12469);
or U15815 (N_15815,N_13281,N_13219);
nor U15816 (N_15816,N_12524,N_12741);
xnor U15817 (N_15817,N_12341,N_13148);
nand U15818 (N_15818,N_12921,N_12478);
nand U15819 (N_15819,N_13544,N_12746);
nand U15820 (N_15820,N_12755,N_13552);
nor U15821 (N_15821,N_12943,N_13551);
nor U15822 (N_15822,N_12729,N_12158);
xor U15823 (N_15823,N_12658,N_13541);
nand U15824 (N_15824,N_12685,N_13104);
xnor U15825 (N_15825,N_13061,N_12404);
nor U15826 (N_15826,N_13039,N_12065);
or U15827 (N_15827,N_12120,N_12751);
or U15828 (N_15828,N_12956,N_13204);
xnor U15829 (N_15829,N_13874,N_13875);
nor U15830 (N_15830,N_12691,N_12742);
or U15831 (N_15831,N_13229,N_12213);
nand U15832 (N_15832,N_13714,N_13312);
nor U15833 (N_15833,N_13576,N_12763);
nor U15834 (N_15834,N_13321,N_12118);
nand U15835 (N_15835,N_12708,N_13774);
or U15836 (N_15836,N_13582,N_13033);
xnor U15837 (N_15837,N_13250,N_13298);
nand U15838 (N_15838,N_13888,N_13531);
nor U15839 (N_15839,N_12736,N_13177);
nand U15840 (N_15840,N_12036,N_12591);
or U15841 (N_15841,N_12509,N_12262);
and U15842 (N_15842,N_13662,N_12212);
and U15843 (N_15843,N_13293,N_13085);
xor U15844 (N_15844,N_12217,N_13991);
xor U15845 (N_15845,N_12539,N_13276);
and U15846 (N_15846,N_12619,N_12624);
xnor U15847 (N_15847,N_12762,N_12771);
nor U15848 (N_15848,N_13952,N_12047);
nor U15849 (N_15849,N_13547,N_12846);
xor U15850 (N_15850,N_13880,N_13441);
or U15851 (N_15851,N_13062,N_12658);
nor U15852 (N_15852,N_13032,N_13513);
or U15853 (N_15853,N_13658,N_12212);
nor U15854 (N_15854,N_13574,N_13272);
and U15855 (N_15855,N_12937,N_13222);
xor U15856 (N_15856,N_13504,N_12100);
nor U15857 (N_15857,N_12533,N_13416);
nor U15858 (N_15858,N_12306,N_13088);
nor U15859 (N_15859,N_12185,N_13536);
or U15860 (N_15860,N_13159,N_12548);
or U15861 (N_15861,N_13417,N_12389);
nand U15862 (N_15862,N_13291,N_12979);
nand U15863 (N_15863,N_13943,N_13881);
and U15864 (N_15864,N_13342,N_12372);
or U15865 (N_15865,N_13855,N_13308);
and U15866 (N_15866,N_13595,N_13729);
or U15867 (N_15867,N_12444,N_13601);
nor U15868 (N_15868,N_12483,N_12242);
xor U15869 (N_15869,N_13098,N_13956);
nand U15870 (N_15870,N_12883,N_13858);
nor U15871 (N_15871,N_13341,N_13728);
nor U15872 (N_15872,N_13654,N_13534);
nand U15873 (N_15873,N_13938,N_12827);
xor U15874 (N_15874,N_12210,N_13162);
or U15875 (N_15875,N_12276,N_12752);
or U15876 (N_15876,N_13802,N_12797);
or U15877 (N_15877,N_13153,N_12482);
nor U15878 (N_15878,N_12317,N_12569);
xor U15879 (N_15879,N_12530,N_12804);
nand U15880 (N_15880,N_12436,N_13451);
nand U15881 (N_15881,N_13252,N_13584);
nor U15882 (N_15882,N_13640,N_12489);
xor U15883 (N_15883,N_12748,N_12637);
and U15884 (N_15884,N_13089,N_13364);
and U15885 (N_15885,N_13242,N_12550);
nand U15886 (N_15886,N_13602,N_13253);
nand U15887 (N_15887,N_12113,N_12373);
xnor U15888 (N_15888,N_12714,N_13920);
or U15889 (N_15889,N_13855,N_12593);
nand U15890 (N_15890,N_13710,N_12307);
nand U15891 (N_15891,N_13716,N_13663);
xnor U15892 (N_15892,N_13190,N_12872);
nor U15893 (N_15893,N_13692,N_12461);
xor U15894 (N_15894,N_13485,N_12393);
nand U15895 (N_15895,N_12627,N_13350);
nor U15896 (N_15896,N_12993,N_13716);
nor U15897 (N_15897,N_12448,N_12024);
nand U15898 (N_15898,N_12346,N_13737);
nor U15899 (N_15899,N_12353,N_12791);
or U15900 (N_15900,N_13436,N_13983);
nor U15901 (N_15901,N_13681,N_12308);
nand U15902 (N_15902,N_12424,N_12339);
or U15903 (N_15903,N_12459,N_13606);
or U15904 (N_15904,N_12782,N_12240);
or U15905 (N_15905,N_13004,N_12356);
nor U15906 (N_15906,N_12120,N_12701);
or U15907 (N_15907,N_13253,N_13240);
and U15908 (N_15908,N_13572,N_12670);
or U15909 (N_15909,N_13105,N_13193);
nor U15910 (N_15910,N_12556,N_12977);
xnor U15911 (N_15911,N_13970,N_13232);
or U15912 (N_15912,N_12081,N_13145);
xor U15913 (N_15913,N_13418,N_12771);
xnor U15914 (N_15914,N_12376,N_12172);
nor U15915 (N_15915,N_13122,N_13838);
xor U15916 (N_15916,N_13456,N_12833);
and U15917 (N_15917,N_13648,N_12881);
and U15918 (N_15918,N_13695,N_13254);
xnor U15919 (N_15919,N_12260,N_13263);
or U15920 (N_15920,N_12776,N_12489);
nor U15921 (N_15921,N_12841,N_12925);
nor U15922 (N_15922,N_12890,N_12884);
nand U15923 (N_15923,N_13755,N_13466);
nor U15924 (N_15924,N_13025,N_13611);
nand U15925 (N_15925,N_12539,N_13112);
nor U15926 (N_15926,N_13056,N_12067);
or U15927 (N_15927,N_13807,N_13798);
xnor U15928 (N_15928,N_13022,N_13852);
or U15929 (N_15929,N_12989,N_12637);
nor U15930 (N_15930,N_13638,N_13448);
xor U15931 (N_15931,N_12430,N_13045);
or U15932 (N_15932,N_12740,N_12915);
xnor U15933 (N_15933,N_12459,N_13208);
nand U15934 (N_15934,N_13873,N_13804);
and U15935 (N_15935,N_12769,N_12927);
and U15936 (N_15936,N_12614,N_13452);
nor U15937 (N_15937,N_13351,N_12760);
nand U15938 (N_15938,N_13232,N_13294);
nand U15939 (N_15939,N_12184,N_13290);
nor U15940 (N_15940,N_13317,N_13702);
or U15941 (N_15941,N_13345,N_13138);
nor U15942 (N_15942,N_12162,N_12719);
and U15943 (N_15943,N_13061,N_13831);
xor U15944 (N_15944,N_13568,N_13361);
or U15945 (N_15945,N_12966,N_13433);
and U15946 (N_15946,N_12739,N_12660);
nand U15947 (N_15947,N_12463,N_13454);
or U15948 (N_15948,N_13170,N_13068);
and U15949 (N_15949,N_12926,N_12248);
nor U15950 (N_15950,N_13717,N_12400);
or U15951 (N_15951,N_12961,N_12012);
or U15952 (N_15952,N_13456,N_13509);
and U15953 (N_15953,N_12340,N_13750);
nand U15954 (N_15954,N_13328,N_12613);
and U15955 (N_15955,N_13504,N_13900);
nor U15956 (N_15956,N_12799,N_12631);
xnor U15957 (N_15957,N_13301,N_13020);
and U15958 (N_15958,N_12753,N_12148);
nor U15959 (N_15959,N_13382,N_12648);
nand U15960 (N_15960,N_13660,N_12172);
nor U15961 (N_15961,N_12267,N_12186);
nor U15962 (N_15962,N_13306,N_13638);
nand U15963 (N_15963,N_13874,N_13421);
nand U15964 (N_15964,N_12158,N_13650);
or U15965 (N_15965,N_13488,N_13358);
nand U15966 (N_15966,N_13170,N_13016);
nor U15967 (N_15967,N_12382,N_13687);
nor U15968 (N_15968,N_13160,N_13223);
and U15969 (N_15969,N_12309,N_12716);
and U15970 (N_15970,N_13669,N_12294);
xor U15971 (N_15971,N_13101,N_12312);
nor U15972 (N_15972,N_13650,N_13595);
nand U15973 (N_15973,N_12087,N_12535);
nand U15974 (N_15974,N_12100,N_13090);
xnor U15975 (N_15975,N_13241,N_12395);
nor U15976 (N_15976,N_13065,N_12560);
and U15977 (N_15977,N_13351,N_12545);
nand U15978 (N_15978,N_13373,N_13404);
or U15979 (N_15979,N_13392,N_13175);
or U15980 (N_15980,N_13771,N_12112);
or U15981 (N_15981,N_12527,N_12884);
nor U15982 (N_15982,N_13868,N_13045);
nand U15983 (N_15983,N_13981,N_12314);
and U15984 (N_15984,N_13052,N_13198);
nor U15985 (N_15985,N_12599,N_13554);
or U15986 (N_15986,N_13270,N_12681);
xor U15987 (N_15987,N_12688,N_13515);
and U15988 (N_15988,N_13450,N_12511);
xor U15989 (N_15989,N_13475,N_12597);
and U15990 (N_15990,N_13070,N_12028);
xnor U15991 (N_15991,N_13601,N_13995);
and U15992 (N_15992,N_13382,N_13844);
nand U15993 (N_15993,N_12640,N_12101);
and U15994 (N_15994,N_13302,N_13330);
or U15995 (N_15995,N_12632,N_13790);
nand U15996 (N_15996,N_13728,N_12522);
and U15997 (N_15997,N_13430,N_12241);
nor U15998 (N_15998,N_13541,N_12136);
nor U15999 (N_15999,N_13205,N_12410);
or U16000 (N_16000,N_15186,N_15752);
xnor U16001 (N_16001,N_14867,N_14405);
nor U16002 (N_16002,N_14213,N_15581);
and U16003 (N_16003,N_14234,N_14317);
nand U16004 (N_16004,N_14595,N_15905);
and U16005 (N_16005,N_14268,N_14382);
nor U16006 (N_16006,N_14763,N_15377);
or U16007 (N_16007,N_15511,N_14798);
xor U16008 (N_16008,N_14009,N_14462);
xor U16009 (N_16009,N_14486,N_14244);
nor U16010 (N_16010,N_15745,N_15322);
or U16011 (N_16011,N_15915,N_15487);
nor U16012 (N_16012,N_15221,N_14929);
nor U16013 (N_16013,N_15174,N_14037);
nand U16014 (N_16014,N_15357,N_14396);
or U16015 (N_16015,N_14573,N_14022);
nor U16016 (N_16016,N_15200,N_14576);
or U16017 (N_16017,N_15716,N_14957);
and U16018 (N_16018,N_14250,N_14696);
nand U16019 (N_16019,N_15721,N_15091);
or U16020 (N_16020,N_15197,N_14948);
xor U16021 (N_16021,N_14888,N_14899);
nand U16022 (N_16022,N_14121,N_14032);
nand U16023 (N_16023,N_15268,N_14509);
and U16024 (N_16024,N_15757,N_14316);
nor U16025 (N_16025,N_14094,N_15630);
nand U16026 (N_16026,N_14113,N_15894);
nand U16027 (N_16027,N_14143,N_15619);
nor U16028 (N_16028,N_15201,N_14707);
nand U16029 (N_16029,N_15566,N_15374);
nor U16030 (N_16030,N_15154,N_15399);
nor U16031 (N_16031,N_14089,N_14669);
nor U16032 (N_16032,N_14521,N_15868);
xor U16033 (N_16033,N_15016,N_14528);
or U16034 (N_16034,N_14066,N_14102);
nor U16035 (N_16035,N_14851,N_14108);
or U16036 (N_16036,N_15147,N_15259);
nand U16037 (N_16037,N_14178,N_15576);
nor U16038 (N_16038,N_14709,N_15832);
xnor U16039 (N_16039,N_14255,N_14839);
nand U16040 (N_16040,N_14532,N_15983);
nor U16041 (N_16041,N_14515,N_14799);
nor U16042 (N_16042,N_15215,N_14500);
and U16043 (N_16043,N_14972,N_14917);
nand U16044 (N_16044,N_15559,N_15125);
nand U16045 (N_16045,N_15499,N_14788);
xnor U16046 (N_16046,N_14270,N_15714);
nand U16047 (N_16047,N_14564,N_15993);
nor U16048 (N_16048,N_14133,N_15209);
or U16049 (N_16049,N_14923,N_15638);
and U16050 (N_16050,N_15073,N_15635);
xnor U16051 (N_16051,N_15067,N_15738);
and U16052 (N_16052,N_14645,N_15611);
nor U16053 (N_16053,N_14263,N_15519);
and U16054 (N_16054,N_14750,N_15381);
nor U16055 (N_16055,N_14451,N_15942);
nor U16056 (N_16056,N_14442,N_14075);
or U16057 (N_16057,N_15945,N_15601);
xor U16058 (N_16058,N_15937,N_15303);
xnor U16059 (N_16059,N_15903,N_15312);
nand U16060 (N_16060,N_14909,N_15204);
nor U16061 (N_16061,N_14218,N_15673);
and U16062 (N_16062,N_14099,N_15114);
nand U16063 (N_16063,N_15033,N_15177);
nand U16064 (N_16064,N_14552,N_15934);
xor U16065 (N_16065,N_14424,N_15065);
xnor U16066 (N_16066,N_15838,N_15086);
nand U16067 (N_16067,N_15090,N_14474);
or U16068 (N_16068,N_14780,N_15867);
nor U16069 (N_16069,N_14057,N_14512);
nand U16070 (N_16070,N_15830,N_15421);
nand U16071 (N_16071,N_14273,N_14119);
xor U16072 (N_16072,N_14012,N_14704);
xor U16073 (N_16073,N_14240,N_15495);
nor U16074 (N_16074,N_15040,N_15012);
and U16075 (N_16075,N_15916,N_14334);
and U16076 (N_16076,N_15483,N_14242);
nand U16077 (N_16077,N_14578,N_14694);
or U16078 (N_16078,N_14772,N_15530);
nand U16079 (N_16079,N_15320,N_15331);
or U16080 (N_16080,N_14706,N_14294);
nand U16081 (N_16081,N_14693,N_14630);
and U16082 (N_16082,N_15473,N_14196);
and U16083 (N_16083,N_14664,N_14949);
or U16084 (N_16084,N_14077,N_14737);
nand U16085 (N_16085,N_14953,N_15363);
xor U16086 (N_16086,N_15685,N_14292);
nand U16087 (N_16087,N_14103,N_14175);
and U16088 (N_16088,N_15663,N_15648);
nor U16089 (N_16089,N_15893,N_14874);
and U16090 (N_16090,N_15129,N_15340);
and U16091 (N_16091,N_14388,N_15857);
nor U16092 (N_16092,N_14990,N_14079);
xor U16093 (N_16093,N_14766,N_15346);
nor U16094 (N_16094,N_15626,N_14768);
nor U16095 (N_16095,N_14655,N_15737);
or U16096 (N_16096,N_15094,N_15475);
and U16097 (N_16097,N_15116,N_14914);
nand U16098 (N_16098,N_14942,N_15624);
and U16099 (N_16099,N_14026,N_15080);
or U16100 (N_16100,N_14078,N_14735);
and U16101 (N_16101,N_15370,N_15068);
nand U16102 (N_16102,N_14385,N_15613);
nand U16103 (N_16103,N_14201,N_15369);
xor U16104 (N_16104,N_15152,N_15183);
or U16105 (N_16105,N_14393,N_14035);
nand U16106 (N_16106,N_14025,N_14215);
or U16107 (N_16107,N_15731,N_14973);
or U16108 (N_16108,N_15072,N_15769);
xor U16109 (N_16109,N_15438,N_15647);
xor U16110 (N_16110,N_15967,N_14599);
nand U16111 (N_16111,N_15609,N_14369);
xnor U16112 (N_16112,N_14863,N_14351);
nor U16113 (N_16113,N_15866,N_14376);
xor U16114 (N_16114,N_14427,N_14116);
and U16115 (N_16115,N_14871,N_14115);
nor U16116 (N_16116,N_15289,N_14907);
or U16117 (N_16117,N_15429,N_14819);
nor U16118 (N_16118,N_15840,N_15284);
xor U16119 (N_16119,N_14995,N_15664);
and U16120 (N_16120,N_15833,N_14505);
nand U16121 (N_16121,N_15546,N_15598);
or U16122 (N_16122,N_14588,N_14643);
or U16123 (N_16123,N_14997,N_15575);
or U16124 (N_16124,N_14674,N_14232);
xor U16125 (N_16125,N_14177,N_14940);
nor U16126 (N_16126,N_14721,N_15407);
nor U16127 (N_16127,N_15235,N_14168);
or U16128 (N_16128,N_14549,N_15747);
nor U16129 (N_16129,N_14455,N_14280);
or U16130 (N_16130,N_15127,N_14120);
and U16131 (N_16131,N_15538,N_14597);
nor U16132 (N_16132,N_14181,N_14620);
nor U16133 (N_16133,N_15654,N_15311);
nand U16134 (N_16134,N_15217,N_14767);
nor U16135 (N_16135,N_15749,N_15006);
and U16136 (N_16136,N_14151,N_15310);
nor U16137 (N_16137,N_14651,N_14147);
xor U16138 (N_16138,N_14619,N_15213);
xor U16139 (N_16139,N_15496,N_14987);
and U16140 (N_16140,N_14412,N_14739);
or U16141 (N_16141,N_15314,N_15264);
or U16142 (N_16142,N_14876,N_15105);
nand U16143 (N_16143,N_15921,N_14345);
xnor U16144 (N_16144,N_15489,N_15179);
and U16145 (N_16145,N_14493,N_14904);
or U16146 (N_16146,N_15274,N_14145);
nor U16147 (N_16147,N_14033,N_14587);
xor U16148 (N_16148,N_14327,N_15972);
nand U16149 (N_16149,N_14323,N_14098);
nor U16150 (N_16150,N_15301,N_14258);
and U16151 (N_16151,N_14279,N_15912);
and U16152 (N_16152,N_15100,N_14807);
and U16153 (N_16153,N_15155,N_14671);
nand U16154 (N_16154,N_14295,N_14642);
nor U16155 (N_16155,N_15004,N_14123);
or U16156 (N_16156,N_14503,N_14966);
and U16157 (N_16157,N_14809,N_15002);
nand U16158 (N_16158,N_15076,N_15468);
nand U16159 (N_16159,N_15614,N_14269);
nor U16160 (N_16160,N_15777,N_14004);
nand U16161 (N_16161,N_14996,N_15275);
or U16162 (N_16162,N_15359,N_14383);
nor U16163 (N_16163,N_14541,N_15656);
or U16164 (N_16164,N_15389,N_15232);
nand U16165 (N_16165,N_14525,N_14600);
nor U16166 (N_16166,N_14373,N_14530);
xor U16167 (N_16167,N_15957,N_15978);
xor U16168 (N_16168,N_14374,N_15774);
or U16169 (N_16169,N_15587,N_14017);
and U16170 (N_16170,N_15266,N_15296);
and U16171 (N_16171,N_15189,N_15435);
and U16172 (N_16172,N_15782,N_14624);
nor U16173 (N_16173,N_14924,N_14325);
xor U16174 (N_16174,N_15641,N_14076);
and U16175 (N_16175,N_14372,N_14538);
xor U16176 (N_16176,N_14992,N_15940);
nand U16177 (N_16177,N_14824,N_15115);
nand U16178 (N_16178,N_14598,N_14744);
nand U16179 (N_16179,N_14591,N_15554);
nand U16180 (N_16180,N_15662,N_14061);
xnor U16181 (N_16181,N_14014,N_14933);
and U16182 (N_16182,N_14641,N_15740);
xnor U16183 (N_16183,N_15616,N_15456);
nor U16184 (N_16184,N_15474,N_15084);
or U16185 (N_16185,N_15350,N_15533);
and U16186 (N_16186,N_15805,N_14575);
and U16187 (N_16187,N_14833,N_14231);
xor U16188 (N_16188,N_14106,N_15578);
nor U16189 (N_16189,N_15427,N_15168);
nor U16190 (N_16190,N_15053,N_14358);
xnor U16191 (N_16191,N_14795,N_14746);
or U16192 (N_16192,N_15979,N_15313);
or U16193 (N_16193,N_14592,N_15172);
or U16194 (N_16194,N_15842,N_14853);
or U16195 (N_16195,N_14485,N_14324);
xor U16196 (N_16196,N_15078,N_15584);
nor U16197 (N_16197,N_15552,N_15280);
xor U16198 (N_16198,N_14332,N_14375);
and U16199 (N_16199,N_15397,N_15282);
nand U16200 (N_16200,N_15410,N_15079);
or U16201 (N_16201,N_14127,N_14105);
and U16202 (N_16202,N_15454,N_15964);
and U16203 (N_16203,N_15477,N_14790);
xor U16204 (N_16204,N_14760,N_15096);
or U16205 (N_16205,N_15674,N_14813);
nand U16206 (N_16206,N_15527,N_15884);
nand U16207 (N_16207,N_14056,N_15253);
xnor U16208 (N_16208,N_14858,N_15060);
xor U16209 (N_16209,N_14524,N_15193);
and U16210 (N_16210,N_15862,N_15831);
nor U16211 (N_16211,N_14237,N_15117);
or U16212 (N_16212,N_14705,N_14734);
nand U16213 (N_16213,N_14457,N_14381);
nor U16214 (N_16214,N_14691,N_14342);
nand U16215 (N_16215,N_14313,N_15387);
nand U16216 (N_16216,N_14986,N_15623);
and U16217 (N_16217,N_14417,N_15759);
and U16218 (N_16218,N_15678,N_15974);
or U16219 (N_16219,N_15005,N_15953);
and U16220 (N_16220,N_14310,N_15743);
xnor U16221 (N_16221,N_15844,N_15514);
or U16222 (N_16222,N_14665,N_15419);
or U16223 (N_16223,N_15826,N_15327);
xnor U16224 (N_16224,N_15988,N_15283);
nand U16225 (N_16225,N_15412,N_14781);
nor U16226 (N_16226,N_15702,N_14783);
nor U16227 (N_16227,N_15099,N_14900);
nor U16228 (N_16228,N_15706,N_15902);
nand U16229 (N_16229,N_15118,N_15599);
nand U16230 (N_16230,N_14446,N_15890);
nor U16231 (N_16231,N_15064,N_15020);
and U16232 (N_16232,N_14330,N_15741);
xor U16233 (N_16233,N_14960,N_14138);
nor U16234 (N_16234,N_15691,N_14680);
xor U16235 (N_16235,N_14341,N_15765);
nor U16236 (N_16236,N_15515,N_14171);
or U16237 (N_16237,N_14019,N_15355);
nand U16238 (N_16238,N_15285,N_15265);
nand U16239 (N_16239,N_14303,N_14366);
xor U16240 (N_16240,N_14445,N_14610);
and U16241 (N_16241,N_14319,N_14498);
and U16242 (N_16242,N_15877,N_14208);
xor U16243 (N_16243,N_15956,N_14754);
nand U16244 (N_16244,N_14956,N_15476);
nor U16245 (N_16245,N_14305,N_15700);
nand U16246 (N_16246,N_14639,N_15491);
and U16247 (N_16247,N_15243,N_15290);
or U16248 (N_16248,N_15651,N_15582);
or U16249 (N_16249,N_14540,N_15037);
or U16250 (N_16250,N_15698,N_14774);
and U16251 (N_16251,N_15169,N_15795);
or U16252 (N_16252,N_15593,N_14981);
nand U16253 (N_16253,N_15182,N_15398);
and U16254 (N_16254,N_14093,N_15430);
nor U16255 (N_16255,N_15316,N_15657);
xor U16256 (N_16256,N_15501,N_15985);
nand U16257 (N_16257,N_15439,N_14873);
or U16258 (N_16258,N_14190,N_14055);
nand U16259 (N_16259,N_14002,N_15778);
or U16260 (N_16260,N_15879,N_14632);
xor U16261 (N_16261,N_14742,N_14036);
xor U16262 (N_16262,N_15208,N_15690);
and U16263 (N_16263,N_14663,N_15408);
xor U16264 (N_16264,N_14666,N_15404);
or U16265 (N_16265,N_14561,N_14164);
or U16266 (N_16266,N_15755,N_15464);
xnor U16267 (N_16267,N_15211,N_15242);
xnor U16268 (N_16268,N_14869,N_14355);
or U16269 (N_16269,N_14413,N_14608);
nand U16270 (N_16270,N_14596,N_15718);
xnor U16271 (N_16271,N_15267,N_14761);
nor U16272 (N_16272,N_14927,N_15845);
xnor U16273 (N_16273,N_14048,N_15991);
nor U16274 (N_16274,N_15181,N_14901);
xnor U16275 (N_16275,N_14502,N_15136);
nor U16276 (N_16276,N_15085,N_15949);
nor U16277 (N_16277,N_15922,N_14193);
and U16278 (N_16278,N_14884,N_14932);
nand U16279 (N_16279,N_14826,N_14364);
nor U16280 (N_16280,N_14203,N_15770);
or U16281 (N_16281,N_14365,N_15665);
xnor U16282 (N_16282,N_15571,N_15590);
nor U16283 (N_16283,N_15110,N_14534);
nand U16284 (N_16284,N_15908,N_14647);
or U16285 (N_16285,N_15711,N_15695);
xor U16286 (N_16286,N_14830,N_14659);
xnor U16287 (N_16287,N_15637,N_14160);
nor U16288 (N_16288,N_14343,N_15071);
nand U16289 (N_16289,N_14891,N_14702);
or U16290 (N_16290,N_14452,N_15403);
nand U16291 (N_16291,N_15560,N_15803);
and U16292 (N_16292,N_15302,N_15853);
or U16293 (N_16293,N_15083,N_14444);
or U16294 (N_16294,N_15708,N_14741);
xor U16295 (N_16295,N_14660,N_15895);
nor U16296 (N_16296,N_14510,N_14640);
and U16297 (N_16297,N_14267,N_14233);
or U16298 (N_16298,N_14377,N_14321);
and U16299 (N_16299,N_14110,N_15325);
nor U16300 (N_16300,N_15141,N_15886);
or U16301 (N_16301,N_14834,N_15195);
nand U16302 (N_16302,N_15022,N_14216);
and U16303 (N_16303,N_15380,N_15286);
nand U16304 (N_16304,N_15825,N_15874);
and U16305 (N_16305,N_15423,N_14349);
nor U16306 (N_16306,N_14314,N_15863);
and U16307 (N_16307,N_14829,N_15277);
nor U16308 (N_16308,N_15750,N_15097);
nand U16309 (N_16309,N_15939,N_14423);
nand U16310 (N_16310,N_15732,N_14636);
or U16311 (N_16311,N_15612,N_15586);
and U16312 (N_16312,N_14835,N_14565);
nand U16313 (N_16313,N_15535,N_15353);
nor U16314 (N_16314,N_14410,N_14315);
or U16315 (N_16315,N_14285,N_15223);
and U16316 (N_16316,N_15692,N_15846);
and U16317 (N_16317,N_15335,N_15163);
and U16318 (N_16318,N_15332,N_15725);
and U16319 (N_16319,N_14063,N_15220);
nor U16320 (N_16320,N_14729,N_14003);
nand U16321 (N_16321,N_14703,N_14985);
xnor U16322 (N_16322,N_15192,N_15968);
or U16323 (N_16323,N_15278,N_14522);
nor U16324 (N_16324,N_14080,N_14387);
and U16325 (N_16325,N_14519,N_15245);
and U16326 (N_16326,N_15416,N_14015);
and U16327 (N_16327,N_15437,N_14714);
nor U16328 (N_16328,N_14163,N_14794);
nor U16329 (N_16329,N_14887,N_14222);
xor U16330 (N_16330,N_15442,N_15140);
and U16331 (N_16331,N_14769,N_14477);
nand U16332 (N_16332,N_14889,N_14842);
and U16333 (N_16333,N_14545,N_14980);
and U16334 (N_16334,N_14225,N_14910);
xor U16335 (N_16335,N_15362,N_15864);
xor U16336 (N_16336,N_14261,N_15185);
or U16337 (N_16337,N_14574,N_14149);
xnor U16338 (N_16338,N_15009,N_14898);
xor U16339 (N_16339,N_15579,N_15859);
and U16340 (N_16340,N_15287,N_14837);
or U16341 (N_16341,N_14939,N_14840);
nand U16342 (N_16342,N_15402,N_15384);
nor U16343 (N_16343,N_14131,N_15783);
and U16344 (N_16344,N_14846,N_15528);
and U16345 (N_16345,N_14569,N_15951);
nor U16346 (N_16346,N_15870,N_14958);
xnor U16347 (N_16347,N_15134,N_15167);
nand U16348 (N_16348,N_14125,N_14803);
and U16349 (N_16349,N_15001,N_14437);
xnor U16350 (N_16350,N_15524,N_14389);
nor U16351 (N_16351,N_14938,N_15773);
or U16352 (N_16352,N_15920,N_15622);
nor U16353 (N_16353,N_14018,N_15173);
or U16354 (N_16354,N_14649,N_15032);
xor U16355 (N_16355,N_15126,N_15919);
nand U16356 (N_16356,N_15679,N_14609);
nand U16357 (N_16357,N_14811,N_15390);
or U16358 (N_16358,N_15447,N_15038);
nand U16359 (N_16359,N_14260,N_14712);
nand U16360 (N_16360,N_14426,N_14407);
or U16361 (N_16361,N_14999,N_15300);
nor U16362 (N_16362,N_15931,N_14150);
and U16363 (N_16363,N_14453,N_14007);
or U16364 (N_16364,N_15950,N_15043);
xnor U16365 (N_16365,N_15452,N_14129);
or U16366 (N_16366,N_14013,N_15052);
or U16367 (N_16367,N_14205,N_15015);
or U16368 (N_16368,N_14802,N_15976);
xnor U16369 (N_16369,N_15165,N_14084);
or U16370 (N_16370,N_14625,N_14081);
or U16371 (N_16371,N_15415,N_14652);
and U16372 (N_16372,N_15900,N_14964);
and U16373 (N_16373,N_15361,N_14634);
nor U16374 (N_16374,N_15761,N_14085);
xor U16375 (N_16375,N_15689,N_14724);
and U16376 (N_16376,N_14613,N_15170);
nor U16377 (N_16377,N_15156,N_15502);
or U16378 (N_16378,N_14926,N_15520);
and U16379 (N_16379,N_15260,N_15561);
or U16380 (N_16380,N_14144,N_15629);
and U16381 (N_16381,N_14153,N_15132);
nand U16382 (N_16382,N_14132,N_14879);
nand U16383 (N_16383,N_15449,N_15434);
nand U16384 (N_16384,N_15379,N_15971);
or U16385 (N_16385,N_15104,N_14159);
nor U16386 (N_16386,N_14491,N_15810);
and U16387 (N_16387,N_15047,N_14539);
or U16388 (N_16388,N_15789,N_15329);
xor U16389 (N_16389,N_14611,N_15443);
nand U16390 (N_16390,N_15540,N_15161);
nand U16391 (N_16391,N_14302,N_15339);
or U16392 (N_16392,N_14362,N_14275);
and U16393 (N_16393,N_14350,N_15343);
or U16394 (N_16394,N_14134,N_14386);
or U16395 (N_16395,N_15279,N_15400);
xnor U16396 (N_16396,N_15876,N_15748);
or U16397 (N_16397,N_15639,N_15351);
xor U16398 (N_16398,N_14661,N_15544);
or U16399 (N_16399,N_15734,N_14687);
xor U16400 (N_16400,N_14265,N_14771);
nor U16401 (N_16401,N_14725,N_15724);
xnor U16402 (N_16402,N_14400,N_15425);
nand U16403 (N_16403,N_14058,N_14053);
and U16404 (N_16404,N_14135,N_15035);
nor U16405 (N_16405,N_14277,N_15391);
or U16406 (N_16406,N_14011,N_15786);
nor U16407 (N_16407,N_14301,N_14281);
and U16408 (N_16408,N_14631,N_15345);
nand U16409 (N_16409,N_14204,N_14320);
nand U16410 (N_16410,N_14097,N_15969);
nand U16411 (N_16411,N_15828,N_14379);
xor U16412 (N_16412,N_15615,N_14402);
nor U16413 (N_16413,N_14047,N_14975);
nor U16414 (N_16414,N_14299,N_15045);
xor U16415 (N_16415,N_15550,N_15467);
or U16416 (N_16416,N_14091,N_14797);
or U16417 (N_16417,N_14194,N_15553);
nor U16418 (N_16418,N_14675,N_14069);
or U16419 (N_16419,N_14656,N_15694);
nor U16420 (N_16420,N_15249,N_14928);
and U16421 (N_16421,N_15675,N_14906);
xnor U16422 (N_16422,N_15021,N_14392);
or U16423 (N_16423,N_14390,N_14584);
nand U16424 (N_16424,N_14844,N_15932);
and U16425 (N_16425,N_15779,N_15291);
or U16426 (N_16426,N_15030,N_15461);
nor U16427 (N_16427,N_14757,N_14023);
and U16428 (N_16428,N_14915,N_15224);
and U16429 (N_16429,N_15162,N_14291);
and U16430 (N_16430,N_14676,N_14180);
nor U16431 (N_16431,N_14049,N_14139);
or U16432 (N_16432,N_15070,N_14235);
xor U16433 (N_16433,N_14513,N_14447);
nand U16434 (N_16434,N_14117,N_15677);
nand U16435 (N_16435,N_15946,N_15927);
nand U16436 (N_16436,N_15471,N_14126);
xnor U16437 (N_16437,N_15089,N_15119);
xor U16438 (N_16438,N_14165,N_14715);
nor U16439 (N_16439,N_14494,N_14841);
nand U16440 (N_16440,N_15742,N_14554);
nand U16441 (N_16441,N_14662,N_15981);
nand U16442 (N_16442,N_15372,N_14287);
nor U16443 (N_16443,N_14527,N_14068);
and U16444 (N_16444,N_15225,N_14679);
nor U16445 (N_16445,N_15762,N_15356);
nand U16446 (N_16446,N_15926,N_15848);
xor U16447 (N_16447,N_14759,N_15505);
xnor U16448 (N_16448,N_15898,N_14536);
nor U16449 (N_16449,N_14738,N_14657);
nand U16450 (N_16450,N_14067,N_15796);
xnor U16451 (N_16451,N_15472,N_14852);
xnor U16452 (N_16452,N_14209,N_15653);
nor U16453 (N_16453,N_14967,N_15814);
and U16454 (N_16454,N_15563,N_14843);
nor U16455 (N_16455,N_14397,N_14850);
nand U16456 (N_16456,N_14154,N_15093);
or U16457 (N_16457,N_14248,N_15906);
xor U16458 (N_16458,N_14517,N_14367);
nand U16459 (N_16459,N_15050,N_14866);
xnor U16460 (N_16460,N_15634,N_14582);
nor U16461 (N_16461,N_14475,N_14221);
xnor U16462 (N_16462,N_15298,N_15891);
nand U16463 (N_16463,N_15426,N_14030);
nor U16464 (N_16464,N_15448,N_14770);
nand U16465 (N_16465,N_15056,N_15992);
xor U16466 (N_16466,N_14622,N_14006);
nand U16467 (N_16467,N_15872,N_15240);
and U16468 (N_16468,N_15843,N_15807);
and U16469 (N_16469,N_14988,N_14831);
nand U16470 (N_16470,N_14855,N_14492);
xnor U16471 (N_16471,N_15219,N_14736);
xnor U16472 (N_16472,N_15855,N_15348);
nand U16473 (N_16473,N_15526,N_15112);
and U16474 (N_16474,N_14618,N_14473);
or U16475 (N_16475,N_14810,N_14471);
nand U16476 (N_16476,N_15658,N_15710);
nor U16477 (N_16477,N_15250,N_15366);
and U16478 (N_16478,N_14878,N_14827);
nand U16479 (N_16479,N_15564,N_14883);
or U16480 (N_16480,N_15809,N_15234);
nand U16481 (N_16481,N_15341,N_14629);
or U16482 (N_16482,N_15354,N_14758);
xnor U16483 (N_16483,N_14989,N_15959);
nand U16484 (N_16484,N_14217,N_15124);
and U16485 (N_16485,N_14214,N_14935);
nand U16486 (N_16486,N_15414,N_15555);
nor U16487 (N_16487,N_15371,N_14581);
nor U16488 (N_16488,N_14572,N_15824);
and U16489 (N_16489,N_15108,N_15739);
or U16490 (N_16490,N_14488,N_15405);
or U16491 (N_16491,N_14380,N_15817);
or U16492 (N_16492,N_15897,N_15813);
xnor U16493 (N_16493,N_15851,N_14416);
nand U16494 (N_16494,N_14060,N_14146);
or U16495 (N_16495,N_15568,N_15460);
nand U16496 (N_16496,N_15081,N_14290);
xor U16497 (N_16497,N_14441,N_14563);
and U16498 (N_16498,N_14463,N_15498);
nand U16499 (N_16499,N_15202,N_15263);
or U16500 (N_16500,N_15881,N_15930);
or U16501 (N_16501,N_14732,N_15861);
nor U16502 (N_16502,N_15508,N_14408);
and U16503 (N_16503,N_14628,N_15948);
nand U16504 (N_16504,N_14043,N_14580);
and U16505 (N_16505,N_15055,N_15196);
nand U16506 (N_16506,N_14777,N_15486);
nor U16507 (N_16507,N_14965,N_15000);
or U16508 (N_16508,N_15693,N_14847);
and U16509 (N_16509,N_14677,N_15984);
nor U16510 (N_16510,N_14568,N_15226);
nor U16511 (N_16511,N_15929,N_14456);
nand U16512 (N_16512,N_14249,N_15763);
nand U16513 (N_16513,N_15621,N_15228);
or U16514 (N_16514,N_14224,N_15328);
nand U16515 (N_16515,N_14309,N_15645);
and U16516 (N_16516,N_15176,N_15049);
nand U16517 (N_16517,N_15395,N_14678);
nand U16518 (N_16518,N_14601,N_15482);
or U16519 (N_16519,N_14185,N_15138);
nand U16520 (N_16520,N_14422,N_14912);
xor U16521 (N_16521,N_15066,N_15148);
nor U16522 (N_16522,N_14238,N_14791);
xnor U16523 (N_16523,N_15596,N_15239);
and U16524 (N_16524,N_14637,N_15917);
or U16525 (N_16525,N_15247,N_15970);
xnor U16526 (N_16526,N_15781,N_14930);
nor U16527 (N_16527,N_14466,N_15157);
or U16528 (N_16528,N_14354,N_14559);
nand U16529 (N_16529,N_14436,N_15018);
xor U16530 (N_16530,N_14481,N_15367);
and U16531 (N_16531,N_14179,N_14348);
nand U16532 (N_16532,N_14976,N_14823);
or U16533 (N_16533,N_15820,N_15788);
nand U16534 (N_16534,N_14860,N_15669);
xor U16535 (N_16535,N_14562,N_14962);
and U16536 (N_16536,N_14586,N_15334);
and U16537 (N_16537,N_15835,N_15042);
or U16538 (N_16538,N_15484,N_14191);
xnor U16539 (N_16539,N_15941,N_15470);
and U16540 (N_16540,N_14136,N_14166);
or U16541 (N_16541,N_15713,N_15936);
nor U16542 (N_16542,N_15107,N_14667);
nand U16543 (N_16543,N_14245,N_14499);
and U16544 (N_16544,N_15241,N_14751);
nor U16545 (N_16545,N_15406,N_15744);
or U16546 (N_16546,N_15592,N_14708);
or U16547 (N_16547,N_15799,N_14590);
xnor U16548 (N_16548,N_14692,N_15980);
xnor U16549 (N_16549,N_14368,N_15998);
xor U16550 (N_16550,N_15292,N_15420);
or U16551 (N_16551,N_14278,N_15997);
or U16552 (N_16552,N_14728,N_15982);
xnor U16553 (N_16553,N_14478,N_15558);
and U16554 (N_16554,N_15146,N_15494);
nand U16555 (N_16555,N_14192,N_15446);
xnor U16556 (N_16556,N_15701,N_15466);
xor U16557 (N_16557,N_15704,N_14646);
nor U16558 (N_16558,N_15194,N_14257);
xnor U16559 (N_16559,N_14779,N_14921);
nor U16560 (N_16560,N_15212,N_15054);
nand U16561 (N_16561,N_14176,N_15276);
or U16562 (N_16562,N_14259,N_14336);
or U16563 (N_16563,N_14922,N_15028);
and U16564 (N_16564,N_14027,N_15650);
or U16565 (N_16565,N_15865,N_14710);
and U16566 (N_16566,N_14284,N_15150);
or U16567 (N_16567,N_14968,N_15756);
xor U16568 (N_16568,N_14993,N_14311);
and U16569 (N_16569,N_15604,N_14096);
and U16570 (N_16570,N_14604,N_15850);
and U16571 (N_16571,N_14585,N_15251);
nand U16572 (N_16572,N_15506,N_15503);
nand U16573 (N_16573,N_14419,N_15504);
or U16574 (N_16574,N_14434,N_14583);
xnor U16575 (N_16575,N_15368,N_14832);
and U16576 (N_16576,N_14892,N_14378);
and U16577 (N_16577,N_15059,N_15591);
nor U16578 (N_16578,N_14420,N_14148);
or U16579 (N_16579,N_14229,N_15440);
xnor U16580 (N_16580,N_14688,N_14062);
nand U16581 (N_16581,N_14363,N_15288);
or U16582 (N_16582,N_14950,N_15888);
or U16583 (N_16583,N_14885,N_15297);
xor U16584 (N_16584,N_14683,N_14415);
xnor U16585 (N_16585,N_15122,N_14083);
nor U16586 (N_16586,N_15676,N_14230);
or U16587 (N_16587,N_14100,N_14223);
xnor U16588 (N_16588,N_15871,N_14438);
nor U16589 (N_16589,N_14685,N_15547);
nor U16590 (N_16590,N_14607,N_15557);
or U16591 (N_16591,N_15914,N_15834);
or U16592 (N_16592,N_15383,N_14200);
or U16593 (N_16593,N_15510,N_14395);
nand U16594 (N_16594,N_14161,N_15620);
nor U16595 (N_16595,N_14352,N_14140);
xnor U16596 (N_16596,N_14755,N_15730);
and U16597 (N_16597,N_14040,N_15246);
xnor U16598 (N_16598,N_15913,N_14207);
nor U16599 (N_16599,N_15733,N_14394);
and U16600 (N_16600,N_14838,N_14182);
nand U16601 (N_16601,N_15901,N_14482);
nand U16602 (N_16602,N_15507,N_15827);
nor U16603 (N_16603,N_15411,N_15409);
and U16604 (N_16604,N_14088,N_14142);
xor U16605 (N_16605,N_14606,N_15203);
or U16606 (N_16606,N_15309,N_14944);
xnor U16607 (N_16607,N_15766,N_14195);
xor U16608 (N_16608,N_15342,N_15523);
and U16609 (N_16609,N_14211,N_15024);
xnor U16610 (N_16610,N_14241,N_14338);
nor U16611 (N_16611,N_15462,N_15588);
or U16612 (N_16612,N_15159,N_14753);
xnor U16613 (N_16613,N_15166,N_14716);
xor U16614 (N_16614,N_14699,N_15655);
and U16615 (N_16615,N_15019,N_15918);
xnor U16616 (N_16616,N_14745,N_14551);
xor U16617 (N_16617,N_15458,N_14785);
nor U16618 (N_16618,N_14733,N_14893);
and U16619 (N_16619,N_15802,N_15109);
or U16620 (N_16620,N_14340,N_15023);
or U16621 (N_16621,N_15352,N_14817);
or U16622 (N_16622,N_15633,N_15441);
xor U16623 (N_16623,N_15269,N_14954);
nand U16624 (N_16624,N_14199,N_15088);
nand U16625 (N_16625,N_14723,N_14210);
nand U16626 (N_16626,N_15376,N_15727);
and U16627 (N_16627,N_14862,N_14672);
and U16628 (N_16628,N_15349,N_14429);
nor U16629 (N_16629,N_14896,N_14686);
xnor U16630 (N_16630,N_14360,N_15760);
or U16631 (N_16631,N_14254,N_15534);
nand U16632 (N_16632,N_14936,N_15882);
nand U16633 (N_16633,N_15281,N_15808);
and U16634 (N_16634,N_14202,N_14256);
nor U16635 (N_16635,N_15190,N_15819);
and U16636 (N_16636,N_15670,N_15837);
and U16637 (N_16637,N_15436,N_14087);
and U16638 (N_16638,N_14065,N_14370);
nand U16639 (N_16639,N_15378,N_14947);
or U16640 (N_16640,N_14300,N_15092);
or U16641 (N_16641,N_15536,N_14322);
nor U16642 (N_16642,N_15517,N_14991);
nor U16643 (N_16643,N_14000,N_14016);
and U16644 (N_16644,N_15237,N_15726);
xnor U16645 (N_16645,N_14589,N_15562);
nand U16646 (N_16646,N_15772,N_14266);
xor U16647 (N_16647,N_14480,N_14895);
nand U16648 (N_16648,N_15617,N_15244);
or U16649 (N_16649,N_14952,N_14228);
nor U16650 (N_16650,N_15758,N_14518);
or U16651 (N_16651,N_15597,N_14749);
xnor U16652 (N_16652,N_15797,N_14024);
xnor U16653 (N_16653,N_15767,N_14546);
nand U16654 (N_16654,N_15705,N_15643);
or U16655 (N_16655,N_15537,N_14052);
nand U16656 (N_16656,N_15063,N_15516);
nor U16657 (N_16657,N_15644,N_15883);
nand U16658 (N_16658,N_15010,N_14614);
or U16659 (N_16659,N_14430,N_14567);
nand U16660 (N_16660,N_15618,N_15792);
and U16661 (N_16661,N_15149,N_15227);
nand U16662 (N_16662,N_14252,N_14740);
or U16663 (N_16663,N_15995,N_15026);
nor U16664 (N_16664,N_14700,N_15074);
nor U16665 (N_16665,N_15158,N_14848);
nand U16666 (N_16666,N_15315,N_14183);
nand U16667 (N_16667,N_14535,N_15923);
xor U16668 (N_16668,N_15175,N_15935);
nor U16669 (N_16669,N_15632,N_14875);
nand U16670 (N_16670,N_15144,N_14946);
nor U16671 (N_16671,N_15385,N_15602);
xnor U16672 (N_16672,N_14713,N_14347);
xnor U16673 (N_16673,N_14391,N_15873);
and U16674 (N_16674,N_15509,N_14526);
nand U16675 (N_16675,N_15735,N_15580);
nor U16676 (N_16676,N_14542,N_15880);
or U16677 (N_16677,N_14726,N_14668);
nand U16678 (N_16678,N_14118,N_15989);
and U16679 (N_16679,N_15424,N_15034);
and U16680 (N_16680,N_15143,N_14919);
nor U16681 (N_16681,N_15382,N_15459);
nand U16682 (N_16682,N_15233,N_14306);
xnor U16683 (N_16683,N_14198,N_15583);
or U16684 (N_16684,N_15671,N_15990);
nor U16685 (N_16685,N_14157,N_14616);
or U16686 (N_16686,N_14414,N_15999);
nor U16687 (N_16687,N_15326,N_14289);
nand U16688 (N_16688,N_15911,N_15057);
nor U16689 (N_16689,N_14130,N_15994);
or U16690 (N_16690,N_14805,N_14752);
xnor U16691 (N_16691,N_14886,N_14226);
xor U16692 (N_16692,N_15252,N_15128);
or U16693 (N_16693,N_14961,N_15954);
and U16694 (N_16694,N_14398,N_15373);
nor U16695 (N_16695,N_15860,N_15493);
and U16696 (N_16696,N_14978,N_14428);
xnor U16697 (N_16697,N_15965,N_14635);
or U16698 (N_16698,N_15787,N_14765);
nand U16699 (N_16699,N_15659,N_15330);
nor U16700 (N_16700,N_15338,N_14697);
or U16701 (N_16701,N_14064,N_14558);
nor U16702 (N_16702,N_15258,N_14339);
xor U16703 (N_16703,N_14174,N_15723);
nor U16704 (N_16704,N_14286,N_14925);
nor U16705 (N_16705,N_14570,N_14274);
or U16706 (N_16706,N_15261,N_15027);
nand U16707 (N_16707,N_14054,N_14356);
or U16708 (N_16708,N_15392,N_14484);
nand U16709 (N_16709,N_14916,N_14792);
and U16710 (N_16710,N_14095,N_15102);
nor U16711 (N_16711,N_14421,N_15642);
xnor U16712 (N_16712,N_14406,N_14894);
and U16713 (N_16713,N_14816,N_15736);
nand U16714 (N_16714,N_15565,N_14184);
nand U16715 (N_16715,N_14603,N_15801);
nor U16716 (N_16716,N_14653,N_14044);
or U16717 (N_16717,N_15542,N_14431);
nor U16718 (N_16718,N_14778,N_14727);
nand U16719 (N_16719,N_14974,N_14072);
and U16720 (N_16720,N_15753,N_14051);
xor U16721 (N_16721,N_15551,N_14654);
nor U16722 (N_16722,N_15139,N_14756);
nor U16723 (N_16723,N_14731,N_15014);
nand U16724 (N_16724,N_15444,N_15746);
or U16725 (N_16725,N_14808,N_15490);
xor U16726 (N_16726,N_15270,N_15944);
xnor U16727 (N_16727,N_14312,N_14271);
or U16728 (N_16728,N_14815,N_14308);
and U16729 (N_16729,N_15605,N_14553);
or U16730 (N_16730,N_15822,N_15318);
and U16731 (N_16731,N_14031,N_14821);
nand U16732 (N_16732,N_15776,N_15793);
nor U16733 (N_16733,N_14882,N_15512);
or U16734 (N_16734,N_15687,N_15847);
xor U16735 (N_16735,N_15171,N_15841);
nand U16736 (N_16736,N_15388,N_14468);
and U16737 (N_16737,N_15393,N_14717);
nor U16738 (N_16738,N_14152,N_14167);
xnor U16739 (N_16739,N_14508,N_14571);
nor U16740 (N_16740,N_15003,N_15728);
nor U16741 (N_16741,N_15525,N_15103);
or U16742 (N_16742,N_15130,N_14864);
and U16743 (N_16743,N_14820,N_14784);
or U16744 (N_16744,N_14418,N_14516);
nand U16745 (N_16745,N_14353,N_14796);
nand U16746 (N_16746,N_15113,N_14247);
nand U16747 (N_16747,N_15818,N_14227);
xor U16748 (N_16748,N_14461,N_15492);
or U16749 (N_16749,N_14951,N_14050);
xnor U16750 (N_16750,N_14433,N_15222);
and U16751 (N_16751,N_15358,N_14304);
or U16752 (N_16752,N_15323,N_15131);
or U16753 (N_16753,N_14711,N_15570);
and U16754 (N_16754,N_15469,N_14681);
or U16755 (N_16755,N_14162,N_15660);
nor U16756 (N_16756,N_14764,N_14557);
and U16757 (N_16757,N_15816,N_14288);
xnor U16758 (N_16758,N_14828,N_14617);
nor U16759 (N_16759,N_14937,N_15907);
or U16760 (N_16760,N_15567,N_14326);
nand U16761 (N_16761,N_15029,N_14219);
and U16762 (N_16762,N_14128,N_15943);
nor U16763 (N_16763,N_14998,N_15142);
or U16764 (N_16764,N_15973,N_14460);
xnor U16765 (N_16765,N_14501,N_14543);
nor U16766 (N_16766,N_14548,N_14695);
xnor U16767 (N_16767,N_14789,N_15058);
nor U16768 (N_16768,N_15048,N_14903);
xor U16769 (N_16769,N_15646,N_15652);
nor U16770 (N_16770,N_14359,N_15087);
and U16771 (N_16771,N_14001,N_15480);
or U16772 (N_16772,N_15960,N_14908);
nor U16773 (N_16773,N_14483,N_15722);
xor U16774 (N_16774,N_14220,N_15529);
or U16775 (N_16775,N_14296,N_14822);
nand U16776 (N_16776,N_15684,N_15145);
and U16777 (N_16777,N_14849,N_14854);
nand U16778 (N_16778,N_14690,N_14403);
nor U16779 (N_16779,N_15719,N_14111);
and U16780 (N_16780,N_15075,N_14644);
nor U16781 (N_16781,N_14682,N_15878);
nand U16782 (N_16782,N_14520,N_14467);
and U16783 (N_16783,N_14470,N_15336);
and U16784 (N_16784,N_14934,N_15854);
and U16785 (N_16785,N_15095,N_14870);
nor U16786 (N_16786,N_14856,N_15543);
nand U16787 (N_16787,N_15031,N_15887);
nand U16788 (N_16788,N_14298,N_15885);
nor U16789 (N_16789,N_15821,N_14747);
nand U16790 (N_16790,N_15497,N_14172);
and U16791 (N_16791,N_14931,N_15123);
or U16792 (N_16792,N_14719,N_15899);
xor U16793 (N_16793,N_14722,N_14448);
nor U16794 (N_16794,N_15712,N_15295);
xnor U16795 (N_16795,N_15522,N_15273);
or U16796 (N_16796,N_15852,N_14845);
and U16797 (N_16797,N_15039,N_15703);
xnor U16798 (N_16798,N_14038,N_15513);
nor U16799 (N_16799,N_15337,N_15573);
xor U16800 (N_16800,N_15764,N_15683);
nor U16801 (N_16801,N_15608,N_15306);
or U16802 (N_16802,N_14059,N_15305);
xnor U16803 (N_16803,N_15996,N_14107);
or U16804 (N_16804,N_15481,N_14877);
or U16805 (N_16805,N_15210,N_14092);
nor U16806 (N_16806,N_14042,N_14029);
or U16807 (N_16807,N_14371,N_14633);
and U16808 (N_16808,N_15610,N_14905);
nor U16809 (N_16809,N_14073,N_14490);
and U16810 (N_16810,N_14566,N_14529);
xnor U16811 (N_16811,N_14070,N_15829);
nand U16812 (N_16812,N_14156,N_15178);
or U16813 (N_16813,N_15133,N_14977);
xor U16814 (N_16814,N_14443,N_15649);
xnor U16815 (N_16815,N_14335,N_14086);
xnor U16816 (N_16816,N_14800,N_15082);
or U16817 (N_16817,N_15780,N_14439);
nand U16818 (N_16818,N_15455,N_15606);
nand U16819 (N_16819,N_14212,N_15046);
or U16820 (N_16820,N_15418,N_15680);
and U16821 (N_16821,N_15206,N_14623);
and U16822 (N_16822,N_14114,N_14773);
and U16823 (N_16823,N_14082,N_14272);
and U16824 (N_16824,N_15518,N_14806);
xor U16825 (N_16825,N_15077,N_15977);
or U16826 (N_16826,N_14169,N_15625);
nand U16827 (N_16827,N_15715,N_14333);
nand U16828 (N_16828,N_15453,N_14812);
and U16829 (N_16829,N_14602,N_15036);
and U16830 (N_16830,N_14401,N_15961);
nor U16831 (N_16831,N_15600,N_15198);
xor U16832 (N_16832,N_15257,N_15463);
nand U16833 (N_16833,N_14264,N_14955);
nand U16834 (N_16834,N_15365,N_15603);
nor U16835 (N_16835,N_14173,N_15858);
nand U16836 (N_16836,N_15307,N_15812);
or U16837 (N_16837,N_15904,N_14028);
nor U16838 (N_16838,N_15229,N_14297);
and U16839 (N_16839,N_14698,N_15214);
nand U16840 (N_16840,N_15422,N_15433);
xnor U16841 (N_16841,N_15294,N_14684);
and U16842 (N_16842,N_15800,N_14861);
or U16843 (N_16843,N_15751,N_15098);
nand U16844 (N_16844,N_15595,N_14911);
or U16845 (N_16845,N_15928,N_14718);
and U16846 (N_16846,N_14404,N_15754);
nand U16847 (N_16847,N_14979,N_15101);
xor U16848 (N_16848,N_15457,N_14034);
xor U16849 (N_16849,N_15254,N_14902);
nand U16850 (N_16850,N_14577,N_15798);
and U16851 (N_16851,N_14627,N_15696);
xor U16852 (N_16852,N_15304,N_15187);
nor U16853 (N_16853,N_14435,N_15717);
nand U16854 (N_16854,N_14186,N_15347);
xor U16855 (N_16855,N_15428,N_14090);
xnor U16856 (N_16856,N_14020,N_14648);
and U16857 (N_16857,N_14544,N_14787);
xor U16858 (N_16858,N_15933,N_15062);
and U16859 (N_16859,N_15396,N_14331);
and U16860 (N_16860,N_14246,N_14459);
or U16861 (N_16861,N_15111,N_14329);
nor U16862 (N_16862,N_15299,N_14670);
nand U16863 (N_16863,N_15248,N_15025);
xor U16864 (N_16864,N_14818,N_15216);
and U16865 (N_16865,N_14579,N_14775);
or U16866 (N_16866,N_15051,N_14786);
and U16867 (N_16867,N_15106,N_15811);
nand U16868 (N_16868,N_14399,N_15666);
and U16869 (N_16869,N_14605,N_15485);
nand U16870 (N_16870,N_15975,N_15231);
nand U16871 (N_16871,N_15849,N_15791);
xnor U16872 (N_16872,N_15790,N_15069);
xor U16873 (N_16873,N_14836,N_14638);
nor U16874 (N_16874,N_15667,N_14293);
nand U16875 (N_16875,N_15636,N_15445);
and U16876 (N_16876,N_15044,N_14141);
and U16877 (N_16877,N_15308,N_15577);
nand U16878 (N_16878,N_15806,N_15531);
nand U16879 (N_16879,N_14045,N_15771);
and U16880 (N_16880,N_15205,N_15465);
xnor U16881 (N_16881,N_14612,N_14814);
or U16882 (N_16882,N_15697,N_14658);
or U16883 (N_16883,N_14865,N_15889);
xor U16884 (N_16884,N_14283,N_15594);
nor U16885 (N_16885,N_15413,N_14472);
and U16886 (N_16886,N_15682,N_15333);
and U16887 (N_16887,N_15451,N_14189);
xor U16888 (N_16888,N_14109,N_14074);
xor U16889 (N_16889,N_14101,N_14615);
or U16890 (N_16890,N_14122,N_15386);
and U16891 (N_16891,N_14983,N_14650);
xnor U16892 (N_16892,N_14046,N_14357);
and U16893 (N_16893,N_14793,N_14010);
nand U16894 (N_16894,N_14450,N_15548);
xnor U16895 (N_16895,N_14825,N_15293);
nand U16896 (N_16896,N_14555,N_15432);
or U16897 (N_16897,N_15768,N_14920);
or U16898 (N_16898,N_14041,N_15184);
and U16899 (N_16899,N_14243,N_15262);
nor U16900 (N_16900,N_15688,N_14945);
and U16901 (N_16901,N_14112,N_14547);
nor U16902 (N_16902,N_15775,N_15836);
or U16903 (N_16903,N_14730,N_14550);
nor U16904 (N_16904,N_15585,N_14124);
xnor U16905 (N_16905,N_15823,N_14005);
xnor U16906 (N_16906,N_15317,N_15417);
nor U16907 (N_16907,N_15896,N_14188);
xnor U16908 (N_16908,N_15627,N_14943);
and U16909 (N_16909,N_15008,N_14307);
xor U16910 (N_16910,N_14872,N_15007);
or U16911 (N_16911,N_15364,N_14801);
and U16912 (N_16912,N_14689,N_14963);
nand U16913 (N_16913,N_15804,N_15135);
nand U16914 (N_16914,N_14361,N_14495);
and U16915 (N_16915,N_15574,N_14449);
nand U16916 (N_16916,N_15925,N_15924);
or U16917 (N_16917,N_15236,N_15607);
xnor U16918 (N_16918,N_14476,N_14941);
or U16919 (N_16919,N_15218,N_14626);
xor U16920 (N_16920,N_15668,N_15394);
or U16921 (N_16921,N_14701,N_15164);
or U16922 (N_16922,N_14762,N_14982);
nand U16923 (N_16923,N_14881,N_14913);
nand U16924 (N_16924,N_14868,N_14282);
and U16925 (N_16925,N_14262,N_14720);
and U16926 (N_16926,N_14984,N_15815);
xnor U16927 (N_16927,N_14489,N_14454);
or U16928 (N_16928,N_15952,N_15785);
nor U16929 (N_16929,N_14857,N_15191);
nand U16930 (N_16930,N_14504,N_15869);
nor U16931 (N_16931,N_15875,N_15401);
nor U16932 (N_16932,N_15720,N_14804);
nand U16933 (N_16933,N_14970,N_14506);
nand U16934 (N_16934,N_15856,N_14497);
xnor U16935 (N_16935,N_14346,N_14344);
or U16936 (N_16936,N_15255,N_15500);
or U16937 (N_16937,N_14158,N_14197);
nand U16938 (N_16938,N_15344,N_15180);
or U16939 (N_16939,N_15375,N_15938);
nor U16940 (N_16940,N_15631,N_15151);
or U16941 (N_16941,N_14594,N_14748);
nand U16942 (N_16942,N_14560,N_15545);
nand U16943 (N_16943,N_15319,N_15892);
nor U16944 (N_16944,N_14425,N_15199);
or U16945 (N_16945,N_15986,N_14537);
nor U16946 (N_16946,N_14440,N_15572);
nand U16947 (N_16947,N_15707,N_15532);
xnor U16948 (N_16948,N_14782,N_15230);
nand U16949 (N_16949,N_14621,N_14337);
nor U16950 (N_16950,N_15188,N_15041);
xnor U16951 (N_16951,N_14959,N_14511);
and U16952 (N_16952,N_14432,N_14523);
or U16953 (N_16953,N_15958,N_14859);
nor U16954 (N_16954,N_15238,N_14593);
xor U16955 (N_16955,N_15910,N_14239);
nor U16956 (N_16956,N_15672,N_14533);
and U16957 (N_16957,N_14897,N_14236);
xor U16958 (N_16958,N_15709,N_14465);
xor U16959 (N_16959,N_14071,N_14155);
and U16960 (N_16960,N_15947,N_14039);
and U16961 (N_16961,N_14384,N_15839);
nand U16962 (N_16962,N_15955,N_15569);
nor U16963 (N_16963,N_14251,N_15017);
xor U16964 (N_16964,N_15137,N_14170);
xnor U16965 (N_16965,N_15207,N_14971);
nand U16966 (N_16966,N_15521,N_14104);
nand U16967 (N_16967,N_15153,N_14458);
xnor U16968 (N_16968,N_15681,N_15272);
nand U16969 (N_16969,N_14469,N_14137);
nor U16970 (N_16970,N_14187,N_14479);
nand U16971 (N_16971,N_14206,N_14531);
nand U16972 (N_16972,N_15987,N_14514);
and U16973 (N_16973,N_15556,N_15966);
nor U16974 (N_16974,N_14890,N_14507);
nor U16975 (N_16975,N_15628,N_15431);
xnor U16976 (N_16976,N_15120,N_14328);
nor U16977 (N_16977,N_14673,N_14487);
nor U16978 (N_16978,N_15360,N_15013);
and U16979 (N_16979,N_14556,N_15909);
and U16980 (N_16980,N_15061,N_15160);
nand U16981 (N_16981,N_15640,N_15478);
or U16982 (N_16982,N_15729,N_14276);
nor U16983 (N_16983,N_15321,N_14021);
or U16984 (N_16984,N_14969,N_15324);
xor U16985 (N_16985,N_15539,N_15686);
and U16986 (N_16986,N_14880,N_15256);
nand U16987 (N_16987,N_15661,N_14776);
nor U16988 (N_16988,N_14496,N_15963);
or U16989 (N_16989,N_14743,N_15589);
xnor U16990 (N_16990,N_15121,N_15699);
xnor U16991 (N_16991,N_14411,N_15549);
and U16992 (N_16992,N_14464,N_14994);
nor U16993 (N_16993,N_15784,N_14318);
and U16994 (N_16994,N_15011,N_14008);
xor U16995 (N_16995,N_15541,N_15962);
or U16996 (N_16996,N_15488,N_15479);
and U16997 (N_16997,N_14918,N_14409);
nand U16998 (N_16998,N_15450,N_14253);
nand U16999 (N_16999,N_15271,N_15794);
xnor U17000 (N_17000,N_15615,N_15960);
xor U17001 (N_17001,N_14289,N_14657);
and U17002 (N_17002,N_15340,N_14615);
or U17003 (N_17003,N_14195,N_14956);
or U17004 (N_17004,N_14978,N_15870);
nor U17005 (N_17005,N_15686,N_15205);
nand U17006 (N_17006,N_14689,N_14384);
and U17007 (N_17007,N_15546,N_14303);
and U17008 (N_17008,N_15700,N_14326);
or U17009 (N_17009,N_14108,N_14043);
nor U17010 (N_17010,N_14507,N_14404);
or U17011 (N_17011,N_14283,N_14906);
nand U17012 (N_17012,N_14350,N_15553);
nand U17013 (N_17013,N_15296,N_15598);
nor U17014 (N_17014,N_15977,N_15964);
xor U17015 (N_17015,N_15949,N_14348);
xnor U17016 (N_17016,N_14501,N_15805);
and U17017 (N_17017,N_14029,N_14272);
nand U17018 (N_17018,N_15262,N_14264);
and U17019 (N_17019,N_15585,N_14632);
or U17020 (N_17020,N_15258,N_15721);
nand U17021 (N_17021,N_14587,N_15733);
or U17022 (N_17022,N_14851,N_14988);
nand U17023 (N_17023,N_14384,N_15652);
or U17024 (N_17024,N_15211,N_14107);
nor U17025 (N_17025,N_15005,N_14672);
xor U17026 (N_17026,N_15711,N_15905);
nand U17027 (N_17027,N_15866,N_15310);
nand U17028 (N_17028,N_14665,N_15687);
nor U17029 (N_17029,N_14371,N_14612);
and U17030 (N_17030,N_15237,N_14298);
nor U17031 (N_17031,N_14881,N_15851);
nor U17032 (N_17032,N_14159,N_14931);
or U17033 (N_17033,N_15919,N_14388);
xor U17034 (N_17034,N_15888,N_15221);
and U17035 (N_17035,N_14709,N_15976);
nand U17036 (N_17036,N_15216,N_15947);
xor U17037 (N_17037,N_14255,N_15458);
xnor U17038 (N_17038,N_14435,N_14385);
nor U17039 (N_17039,N_15064,N_15366);
nand U17040 (N_17040,N_14782,N_15380);
or U17041 (N_17041,N_15916,N_14635);
and U17042 (N_17042,N_14548,N_15834);
and U17043 (N_17043,N_14516,N_14114);
nor U17044 (N_17044,N_15699,N_15859);
and U17045 (N_17045,N_15005,N_14544);
nor U17046 (N_17046,N_14474,N_15505);
xnor U17047 (N_17047,N_14601,N_14416);
xnor U17048 (N_17048,N_14552,N_15211);
or U17049 (N_17049,N_15211,N_15838);
nand U17050 (N_17050,N_15364,N_14054);
nor U17051 (N_17051,N_15495,N_14739);
and U17052 (N_17052,N_14367,N_14490);
nor U17053 (N_17053,N_15311,N_15259);
and U17054 (N_17054,N_14139,N_14761);
xnor U17055 (N_17055,N_15619,N_14426);
xnor U17056 (N_17056,N_14190,N_15277);
and U17057 (N_17057,N_14638,N_14815);
nand U17058 (N_17058,N_15723,N_15315);
nand U17059 (N_17059,N_15897,N_14765);
nor U17060 (N_17060,N_14254,N_15909);
xnor U17061 (N_17061,N_15342,N_14575);
nor U17062 (N_17062,N_15251,N_15429);
or U17063 (N_17063,N_15040,N_15052);
or U17064 (N_17064,N_14806,N_15625);
nand U17065 (N_17065,N_14701,N_15199);
xor U17066 (N_17066,N_14896,N_15663);
or U17067 (N_17067,N_14748,N_14875);
nand U17068 (N_17068,N_14499,N_14702);
nor U17069 (N_17069,N_15695,N_15227);
nand U17070 (N_17070,N_15779,N_15695);
nand U17071 (N_17071,N_15960,N_15551);
nand U17072 (N_17072,N_15017,N_15856);
xnor U17073 (N_17073,N_14888,N_14423);
xnor U17074 (N_17074,N_15700,N_14803);
and U17075 (N_17075,N_15165,N_14239);
or U17076 (N_17076,N_14309,N_15711);
or U17077 (N_17077,N_14587,N_15505);
xnor U17078 (N_17078,N_14892,N_14947);
nand U17079 (N_17079,N_15274,N_15186);
nor U17080 (N_17080,N_14168,N_15661);
and U17081 (N_17081,N_14424,N_15909);
nor U17082 (N_17082,N_15717,N_14870);
nand U17083 (N_17083,N_15187,N_14065);
nor U17084 (N_17084,N_14045,N_14492);
or U17085 (N_17085,N_15934,N_14060);
or U17086 (N_17086,N_15761,N_15970);
or U17087 (N_17087,N_14528,N_15222);
nand U17088 (N_17088,N_15423,N_14964);
or U17089 (N_17089,N_14434,N_15178);
or U17090 (N_17090,N_15720,N_15291);
nor U17091 (N_17091,N_15960,N_14356);
nand U17092 (N_17092,N_14854,N_15235);
and U17093 (N_17093,N_15343,N_15246);
nor U17094 (N_17094,N_14207,N_14382);
and U17095 (N_17095,N_14291,N_15644);
xnor U17096 (N_17096,N_15675,N_14207);
nor U17097 (N_17097,N_14767,N_15144);
and U17098 (N_17098,N_15340,N_15861);
or U17099 (N_17099,N_15640,N_15180);
or U17100 (N_17100,N_15933,N_15070);
nor U17101 (N_17101,N_14891,N_15025);
nand U17102 (N_17102,N_15828,N_15113);
or U17103 (N_17103,N_15616,N_15246);
or U17104 (N_17104,N_15819,N_14081);
nand U17105 (N_17105,N_14092,N_14626);
nor U17106 (N_17106,N_14285,N_15729);
and U17107 (N_17107,N_14736,N_14202);
or U17108 (N_17108,N_15229,N_14851);
xor U17109 (N_17109,N_14704,N_14438);
and U17110 (N_17110,N_15599,N_14685);
xor U17111 (N_17111,N_14480,N_14630);
xnor U17112 (N_17112,N_15269,N_14303);
nand U17113 (N_17113,N_15424,N_15279);
nand U17114 (N_17114,N_15696,N_14638);
and U17115 (N_17115,N_14098,N_15557);
or U17116 (N_17116,N_14552,N_15571);
nand U17117 (N_17117,N_14710,N_15631);
and U17118 (N_17118,N_15558,N_14168);
and U17119 (N_17119,N_14098,N_15967);
nor U17120 (N_17120,N_15257,N_15909);
and U17121 (N_17121,N_14217,N_14763);
xor U17122 (N_17122,N_14585,N_15510);
nor U17123 (N_17123,N_15966,N_15814);
or U17124 (N_17124,N_14347,N_14036);
xnor U17125 (N_17125,N_14190,N_14796);
or U17126 (N_17126,N_15619,N_15269);
nand U17127 (N_17127,N_15858,N_15321);
nand U17128 (N_17128,N_14340,N_15973);
and U17129 (N_17129,N_15399,N_14353);
and U17130 (N_17130,N_14991,N_15555);
or U17131 (N_17131,N_14177,N_14064);
or U17132 (N_17132,N_14856,N_15538);
nand U17133 (N_17133,N_15925,N_14030);
or U17134 (N_17134,N_14014,N_14754);
or U17135 (N_17135,N_14721,N_14501);
and U17136 (N_17136,N_15123,N_15337);
and U17137 (N_17137,N_15835,N_15232);
xnor U17138 (N_17138,N_15536,N_15586);
or U17139 (N_17139,N_14927,N_15813);
nand U17140 (N_17140,N_14531,N_15008);
and U17141 (N_17141,N_14771,N_14485);
xor U17142 (N_17142,N_14861,N_14958);
or U17143 (N_17143,N_14060,N_14417);
or U17144 (N_17144,N_15209,N_15826);
or U17145 (N_17145,N_14915,N_15443);
and U17146 (N_17146,N_14577,N_15268);
nor U17147 (N_17147,N_14098,N_14630);
and U17148 (N_17148,N_15754,N_14073);
and U17149 (N_17149,N_14804,N_14450);
nand U17150 (N_17150,N_14980,N_15440);
and U17151 (N_17151,N_15330,N_14962);
and U17152 (N_17152,N_14172,N_14706);
and U17153 (N_17153,N_15908,N_15742);
and U17154 (N_17154,N_14645,N_15220);
nor U17155 (N_17155,N_15983,N_14670);
nand U17156 (N_17156,N_14801,N_14978);
or U17157 (N_17157,N_14221,N_14053);
nor U17158 (N_17158,N_14619,N_14263);
xor U17159 (N_17159,N_14753,N_14573);
nor U17160 (N_17160,N_15365,N_14952);
nand U17161 (N_17161,N_15255,N_14737);
nand U17162 (N_17162,N_15416,N_15135);
and U17163 (N_17163,N_15823,N_14980);
xor U17164 (N_17164,N_15232,N_14538);
nor U17165 (N_17165,N_15681,N_15481);
nor U17166 (N_17166,N_15014,N_14250);
nand U17167 (N_17167,N_14280,N_15275);
and U17168 (N_17168,N_14809,N_15363);
nor U17169 (N_17169,N_15863,N_14614);
nand U17170 (N_17170,N_15543,N_14613);
and U17171 (N_17171,N_14545,N_15120);
or U17172 (N_17172,N_15931,N_15434);
nand U17173 (N_17173,N_14707,N_14379);
nor U17174 (N_17174,N_14748,N_15727);
nand U17175 (N_17175,N_15202,N_14729);
nor U17176 (N_17176,N_14731,N_15467);
nor U17177 (N_17177,N_15079,N_15919);
or U17178 (N_17178,N_14177,N_14394);
or U17179 (N_17179,N_15684,N_14713);
xnor U17180 (N_17180,N_15646,N_14280);
or U17181 (N_17181,N_15039,N_15148);
xor U17182 (N_17182,N_14140,N_15952);
nor U17183 (N_17183,N_15363,N_15292);
nor U17184 (N_17184,N_14265,N_14860);
or U17185 (N_17185,N_14688,N_14919);
nor U17186 (N_17186,N_15059,N_15479);
nor U17187 (N_17187,N_15844,N_15811);
and U17188 (N_17188,N_14462,N_14686);
nor U17189 (N_17189,N_14882,N_14745);
nor U17190 (N_17190,N_15645,N_15294);
or U17191 (N_17191,N_14990,N_15018);
xnor U17192 (N_17192,N_14019,N_15426);
nor U17193 (N_17193,N_15047,N_15789);
nor U17194 (N_17194,N_15333,N_15075);
and U17195 (N_17195,N_15884,N_14861);
nand U17196 (N_17196,N_15858,N_14528);
and U17197 (N_17197,N_15224,N_14074);
or U17198 (N_17198,N_15551,N_14055);
nor U17199 (N_17199,N_14400,N_14563);
or U17200 (N_17200,N_14755,N_15258);
and U17201 (N_17201,N_15567,N_14298);
or U17202 (N_17202,N_15035,N_14329);
and U17203 (N_17203,N_14733,N_14885);
or U17204 (N_17204,N_15550,N_14828);
nor U17205 (N_17205,N_14059,N_15640);
nand U17206 (N_17206,N_15713,N_15915);
and U17207 (N_17207,N_14799,N_14141);
or U17208 (N_17208,N_14332,N_14100);
or U17209 (N_17209,N_14066,N_15312);
and U17210 (N_17210,N_14858,N_14379);
nand U17211 (N_17211,N_15548,N_14556);
xnor U17212 (N_17212,N_15834,N_14443);
and U17213 (N_17213,N_14528,N_15855);
and U17214 (N_17214,N_14124,N_14540);
nand U17215 (N_17215,N_14264,N_15429);
nand U17216 (N_17216,N_14595,N_14804);
xnor U17217 (N_17217,N_14020,N_14494);
xor U17218 (N_17218,N_14641,N_15174);
xor U17219 (N_17219,N_14044,N_15541);
xor U17220 (N_17220,N_15847,N_15551);
nor U17221 (N_17221,N_15808,N_14276);
nor U17222 (N_17222,N_14961,N_14525);
and U17223 (N_17223,N_14416,N_14459);
and U17224 (N_17224,N_15540,N_14879);
xnor U17225 (N_17225,N_15950,N_15470);
nand U17226 (N_17226,N_15137,N_15736);
nand U17227 (N_17227,N_14018,N_14825);
nor U17228 (N_17228,N_15114,N_14727);
xnor U17229 (N_17229,N_14354,N_14108);
or U17230 (N_17230,N_14467,N_14774);
xor U17231 (N_17231,N_15300,N_14454);
or U17232 (N_17232,N_14424,N_14541);
nand U17233 (N_17233,N_15393,N_15671);
or U17234 (N_17234,N_14508,N_15654);
xnor U17235 (N_17235,N_15842,N_14876);
or U17236 (N_17236,N_15541,N_15242);
nand U17237 (N_17237,N_14744,N_15239);
and U17238 (N_17238,N_15642,N_15721);
nor U17239 (N_17239,N_14610,N_14661);
nor U17240 (N_17240,N_14989,N_14881);
and U17241 (N_17241,N_15047,N_14040);
and U17242 (N_17242,N_14054,N_15279);
xnor U17243 (N_17243,N_15705,N_15404);
xor U17244 (N_17244,N_15909,N_15056);
nand U17245 (N_17245,N_14065,N_15858);
or U17246 (N_17246,N_14821,N_14015);
and U17247 (N_17247,N_15785,N_15305);
and U17248 (N_17248,N_14694,N_14891);
nor U17249 (N_17249,N_15926,N_14982);
or U17250 (N_17250,N_15617,N_15199);
or U17251 (N_17251,N_15959,N_15318);
xnor U17252 (N_17252,N_14456,N_15511);
xnor U17253 (N_17253,N_14293,N_15295);
xnor U17254 (N_17254,N_15101,N_14188);
xnor U17255 (N_17255,N_14697,N_14872);
nor U17256 (N_17256,N_14287,N_15799);
xor U17257 (N_17257,N_15035,N_14872);
and U17258 (N_17258,N_15595,N_15902);
and U17259 (N_17259,N_14629,N_14857);
or U17260 (N_17260,N_15198,N_15178);
nand U17261 (N_17261,N_14155,N_14351);
or U17262 (N_17262,N_14690,N_14427);
nor U17263 (N_17263,N_15979,N_15171);
xor U17264 (N_17264,N_14148,N_15903);
or U17265 (N_17265,N_15965,N_15605);
nor U17266 (N_17266,N_14267,N_14707);
nand U17267 (N_17267,N_15352,N_15518);
nor U17268 (N_17268,N_15917,N_14745);
nand U17269 (N_17269,N_15728,N_14899);
and U17270 (N_17270,N_15751,N_14823);
or U17271 (N_17271,N_15003,N_15517);
or U17272 (N_17272,N_14446,N_15894);
or U17273 (N_17273,N_14558,N_14575);
nand U17274 (N_17274,N_14482,N_14685);
nor U17275 (N_17275,N_14116,N_14096);
and U17276 (N_17276,N_15711,N_15683);
xor U17277 (N_17277,N_14002,N_14978);
or U17278 (N_17278,N_14920,N_14989);
and U17279 (N_17279,N_15955,N_14301);
and U17280 (N_17280,N_14274,N_15120);
nor U17281 (N_17281,N_14387,N_14028);
nor U17282 (N_17282,N_14179,N_15901);
nor U17283 (N_17283,N_15928,N_14648);
or U17284 (N_17284,N_15719,N_14045);
nand U17285 (N_17285,N_15686,N_15673);
nor U17286 (N_17286,N_15489,N_14354);
nand U17287 (N_17287,N_15570,N_15157);
and U17288 (N_17288,N_15146,N_15841);
or U17289 (N_17289,N_14887,N_15621);
xnor U17290 (N_17290,N_15727,N_14981);
or U17291 (N_17291,N_15318,N_15202);
nor U17292 (N_17292,N_14559,N_15735);
or U17293 (N_17293,N_15686,N_15325);
xor U17294 (N_17294,N_14862,N_15199);
xor U17295 (N_17295,N_15577,N_14237);
or U17296 (N_17296,N_14546,N_15974);
xnor U17297 (N_17297,N_15868,N_14107);
xor U17298 (N_17298,N_14087,N_14039);
xor U17299 (N_17299,N_14603,N_15701);
nor U17300 (N_17300,N_14797,N_15504);
or U17301 (N_17301,N_15188,N_15205);
nor U17302 (N_17302,N_14779,N_15663);
nor U17303 (N_17303,N_15464,N_14214);
nand U17304 (N_17304,N_15877,N_15204);
nor U17305 (N_17305,N_15578,N_15562);
and U17306 (N_17306,N_14162,N_14438);
or U17307 (N_17307,N_15724,N_15867);
xor U17308 (N_17308,N_15523,N_14023);
xor U17309 (N_17309,N_14492,N_14160);
nor U17310 (N_17310,N_15904,N_15309);
or U17311 (N_17311,N_14748,N_15039);
xnor U17312 (N_17312,N_14011,N_15123);
or U17313 (N_17313,N_14344,N_14982);
nand U17314 (N_17314,N_14387,N_15477);
or U17315 (N_17315,N_14047,N_15861);
nor U17316 (N_17316,N_14815,N_14506);
xor U17317 (N_17317,N_14722,N_14245);
nand U17318 (N_17318,N_15163,N_14769);
nand U17319 (N_17319,N_15141,N_14970);
or U17320 (N_17320,N_14500,N_15996);
nand U17321 (N_17321,N_14856,N_14416);
nor U17322 (N_17322,N_14418,N_14224);
xor U17323 (N_17323,N_15142,N_14963);
or U17324 (N_17324,N_15557,N_15137);
nand U17325 (N_17325,N_15007,N_15291);
nand U17326 (N_17326,N_14346,N_14451);
nor U17327 (N_17327,N_15348,N_14757);
and U17328 (N_17328,N_14563,N_14860);
xor U17329 (N_17329,N_15701,N_15932);
or U17330 (N_17330,N_15100,N_15922);
nor U17331 (N_17331,N_15195,N_15226);
nand U17332 (N_17332,N_14907,N_14961);
xor U17333 (N_17333,N_14151,N_14742);
nand U17334 (N_17334,N_15409,N_15281);
and U17335 (N_17335,N_14656,N_15799);
nand U17336 (N_17336,N_14780,N_14769);
or U17337 (N_17337,N_14713,N_15300);
xnor U17338 (N_17338,N_14276,N_14249);
or U17339 (N_17339,N_14889,N_15871);
or U17340 (N_17340,N_14333,N_14723);
and U17341 (N_17341,N_14092,N_15898);
and U17342 (N_17342,N_14902,N_14996);
nand U17343 (N_17343,N_14090,N_15101);
nand U17344 (N_17344,N_14728,N_14206);
and U17345 (N_17345,N_14664,N_15004);
nand U17346 (N_17346,N_14998,N_14546);
nand U17347 (N_17347,N_14583,N_14608);
nor U17348 (N_17348,N_15016,N_14769);
nor U17349 (N_17349,N_14456,N_14489);
or U17350 (N_17350,N_14593,N_15542);
and U17351 (N_17351,N_15747,N_15232);
or U17352 (N_17352,N_14170,N_14428);
or U17353 (N_17353,N_14661,N_15339);
nand U17354 (N_17354,N_14270,N_15428);
xnor U17355 (N_17355,N_14842,N_14873);
nand U17356 (N_17356,N_14230,N_14574);
and U17357 (N_17357,N_14035,N_14824);
nor U17358 (N_17358,N_14373,N_15341);
or U17359 (N_17359,N_14785,N_15900);
nand U17360 (N_17360,N_15510,N_14870);
and U17361 (N_17361,N_14800,N_14473);
and U17362 (N_17362,N_15236,N_14161);
nor U17363 (N_17363,N_15951,N_15343);
nand U17364 (N_17364,N_14584,N_15941);
or U17365 (N_17365,N_14594,N_15119);
nor U17366 (N_17366,N_15691,N_14038);
or U17367 (N_17367,N_14442,N_14251);
xnor U17368 (N_17368,N_14434,N_15089);
and U17369 (N_17369,N_14732,N_14511);
nand U17370 (N_17370,N_15128,N_15789);
or U17371 (N_17371,N_15181,N_15119);
nand U17372 (N_17372,N_14752,N_15305);
nand U17373 (N_17373,N_15934,N_14088);
nand U17374 (N_17374,N_15133,N_15293);
nand U17375 (N_17375,N_15135,N_15643);
and U17376 (N_17376,N_15498,N_14662);
or U17377 (N_17377,N_14914,N_15133);
xnor U17378 (N_17378,N_15369,N_14572);
nand U17379 (N_17379,N_15643,N_15334);
or U17380 (N_17380,N_14675,N_15713);
and U17381 (N_17381,N_15500,N_15136);
or U17382 (N_17382,N_15026,N_15321);
and U17383 (N_17383,N_15711,N_14994);
and U17384 (N_17384,N_15625,N_14530);
and U17385 (N_17385,N_14392,N_14865);
nand U17386 (N_17386,N_14360,N_15336);
and U17387 (N_17387,N_14785,N_15016);
xor U17388 (N_17388,N_14398,N_15237);
nand U17389 (N_17389,N_14821,N_15625);
or U17390 (N_17390,N_14721,N_14045);
nor U17391 (N_17391,N_14779,N_14818);
nand U17392 (N_17392,N_15389,N_15637);
nor U17393 (N_17393,N_14572,N_15692);
xnor U17394 (N_17394,N_14550,N_14693);
or U17395 (N_17395,N_15809,N_15583);
xnor U17396 (N_17396,N_14375,N_14252);
nand U17397 (N_17397,N_15720,N_14068);
xor U17398 (N_17398,N_15982,N_15287);
nand U17399 (N_17399,N_15460,N_15039);
xor U17400 (N_17400,N_15518,N_15845);
and U17401 (N_17401,N_14694,N_14121);
nand U17402 (N_17402,N_15055,N_14250);
or U17403 (N_17403,N_15195,N_14619);
nor U17404 (N_17404,N_14287,N_15768);
and U17405 (N_17405,N_15146,N_14729);
xor U17406 (N_17406,N_14576,N_15287);
or U17407 (N_17407,N_15301,N_15207);
or U17408 (N_17408,N_14979,N_15763);
and U17409 (N_17409,N_15551,N_15934);
and U17410 (N_17410,N_15252,N_14637);
nor U17411 (N_17411,N_15690,N_15031);
or U17412 (N_17412,N_15126,N_14012);
and U17413 (N_17413,N_15656,N_14670);
xor U17414 (N_17414,N_15931,N_14157);
nor U17415 (N_17415,N_15019,N_14084);
or U17416 (N_17416,N_15189,N_15656);
nand U17417 (N_17417,N_15239,N_14798);
or U17418 (N_17418,N_15325,N_15829);
and U17419 (N_17419,N_14294,N_15838);
xor U17420 (N_17420,N_14461,N_15193);
nor U17421 (N_17421,N_14067,N_14766);
nand U17422 (N_17422,N_14608,N_14795);
or U17423 (N_17423,N_14259,N_14197);
or U17424 (N_17424,N_14219,N_15951);
and U17425 (N_17425,N_14031,N_15975);
or U17426 (N_17426,N_14779,N_15932);
nand U17427 (N_17427,N_14026,N_14947);
or U17428 (N_17428,N_15962,N_14256);
nand U17429 (N_17429,N_14929,N_14805);
or U17430 (N_17430,N_14688,N_15932);
xnor U17431 (N_17431,N_14275,N_14133);
and U17432 (N_17432,N_14031,N_15476);
xor U17433 (N_17433,N_14690,N_15228);
or U17434 (N_17434,N_14519,N_15281);
or U17435 (N_17435,N_14158,N_14584);
nor U17436 (N_17436,N_14032,N_15141);
xor U17437 (N_17437,N_14313,N_14772);
nand U17438 (N_17438,N_14986,N_15596);
or U17439 (N_17439,N_14600,N_15024);
nor U17440 (N_17440,N_15636,N_15158);
nand U17441 (N_17441,N_15846,N_14304);
nor U17442 (N_17442,N_14546,N_14395);
or U17443 (N_17443,N_14868,N_14221);
nand U17444 (N_17444,N_15151,N_15464);
nand U17445 (N_17445,N_15402,N_14012);
nand U17446 (N_17446,N_14284,N_14574);
nor U17447 (N_17447,N_15568,N_14594);
nand U17448 (N_17448,N_14398,N_14928);
and U17449 (N_17449,N_14675,N_14002);
and U17450 (N_17450,N_14849,N_14109);
xnor U17451 (N_17451,N_14527,N_14695);
and U17452 (N_17452,N_15311,N_15691);
nand U17453 (N_17453,N_15102,N_14473);
xnor U17454 (N_17454,N_14761,N_15216);
nand U17455 (N_17455,N_15839,N_15611);
and U17456 (N_17456,N_14136,N_14528);
or U17457 (N_17457,N_14575,N_15866);
nand U17458 (N_17458,N_14452,N_15741);
and U17459 (N_17459,N_14698,N_14131);
xnor U17460 (N_17460,N_14731,N_14448);
nor U17461 (N_17461,N_14692,N_14660);
nand U17462 (N_17462,N_15353,N_14013);
xnor U17463 (N_17463,N_14311,N_14479);
nor U17464 (N_17464,N_14012,N_15090);
nand U17465 (N_17465,N_15213,N_14417);
or U17466 (N_17466,N_15995,N_15051);
nor U17467 (N_17467,N_14818,N_15638);
nor U17468 (N_17468,N_14266,N_14391);
nor U17469 (N_17469,N_15719,N_15514);
and U17470 (N_17470,N_14430,N_15500);
or U17471 (N_17471,N_15678,N_15461);
and U17472 (N_17472,N_15532,N_15086);
nand U17473 (N_17473,N_14540,N_15853);
or U17474 (N_17474,N_14411,N_14019);
nand U17475 (N_17475,N_15147,N_15944);
or U17476 (N_17476,N_15651,N_15312);
xor U17477 (N_17477,N_15475,N_15822);
nand U17478 (N_17478,N_15200,N_14139);
xnor U17479 (N_17479,N_15224,N_14202);
or U17480 (N_17480,N_15555,N_15997);
nor U17481 (N_17481,N_15027,N_14786);
and U17482 (N_17482,N_14807,N_15688);
and U17483 (N_17483,N_14131,N_14194);
nand U17484 (N_17484,N_14463,N_15278);
and U17485 (N_17485,N_15778,N_15166);
and U17486 (N_17486,N_15128,N_14561);
xor U17487 (N_17487,N_15447,N_15967);
nor U17488 (N_17488,N_15111,N_15057);
nor U17489 (N_17489,N_14162,N_15616);
or U17490 (N_17490,N_14851,N_15490);
xor U17491 (N_17491,N_15456,N_14970);
and U17492 (N_17492,N_14473,N_14954);
xnor U17493 (N_17493,N_14533,N_14878);
and U17494 (N_17494,N_14399,N_14503);
nand U17495 (N_17495,N_15366,N_14549);
nor U17496 (N_17496,N_14512,N_15035);
nor U17497 (N_17497,N_15244,N_14794);
and U17498 (N_17498,N_15693,N_15127);
xnor U17499 (N_17499,N_15679,N_14484);
xnor U17500 (N_17500,N_14037,N_15528);
xor U17501 (N_17501,N_15852,N_15323);
xor U17502 (N_17502,N_14973,N_15759);
nand U17503 (N_17503,N_15503,N_14118);
or U17504 (N_17504,N_14062,N_14662);
or U17505 (N_17505,N_14967,N_15624);
and U17506 (N_17506,N_14105,N_15291);
or U17507 (N_17507,N_15578,N_14151);
xnor U17508 (N_17508,N_15225,N_15717);
or U17509 (N_17509,N_14663,N_14541);
nand U17510 (N_17510,N_14994,N_14999);
nor U17511 (N_17511,N_14596,N_15464);
xor U17512 (N_17512,N_14834,N_15740);
or U17513 (N_17513,N_14370,N_15828);
xnor U17514 (N_17514,N_14753,N_14554);
nand U17515 (N_17515,N_14158,N_14787);
xnor U17516 (N_17516,N_14028,N_15746);
nor U17517 (N_17517,N_15852,N_14629);
nand U17518 (N_17518,N_14619,N_14233);
xnor U17519 (N_17519,N_15506,N_15116);
nor U17520 (N_17520,N_14256,N_14685);
or U17521 (N_17521,N_14907,N_14261);
nand U17522 (N_17522,N_14052,N_15150);
and U17523 (N_17523,N_14224,N_15412);
nor U17524 (N_17524,N_14137,N_15513);
xnor U17525 (N_17525,N_15555,N_15206);
or U17526 (N_17526,N_15006,N_14201);
and U17527 (N_17527,N_14116,N_15070);
nand U17528 (N_17528,N_15949,N_15675);
nor U17529 (N_17529,N_14762,N_14556);
or U17530 (N_17530,N_15679,N_15317);
nand U17531 (N_17531,N_15408,N_14670);
or U17532 (N_17532,N_15465,N_14747);
xnor U17533 (N_17533,N_15792,N_14693);
and U17534 (N_17534,N_15477,N_14607);
or U17535 (N_17535,N_14032,N_14612);
xor U17536 (N_17536,N_15052,N_14388);
and U17537 (N_17537,N_14524,N_15116);
xor U17538 (N_17538,N_15876,N_14328);
xor U17539 (N_17539,N_14374,N_14039);
and U17540 (N_17540,N_15218,N_15696);
or U17541 (N_17541,N_15655,N_15557);
and U17542 (N_17542,N_14164,N_14454);
and U17543 (N_17543,N_14992,N_14910);
xor U17544 (N_17544,N_14680,N_15020);
xnor U17545 (N_17545,N_14633,N_14104);
nand U17546 (N_17546,N_15349,N_15180);
nand U17547 (N_17547,N_15228,N_14211);
nand U17548 (N_17548,N_14340,N_14611);
xor U17549 (N_17549,N_14709,N_15474);
nand U17550 (N_17550,N_15398,N_14484);
nor U17551 (N_17551,N_15154,N_14492);
nor U17552 (N_17552,N_14716,N_15234);
xor U17553 (N_17553,N_14495,N_15435);
and U17554 (N_17554,N_14322,N_15428);
and U17555 (N_17555,N_14633,N_15545);
or U17556 (N_17556,N_15355,N_15781);
nand U17557 (N_17557,N_15405,N_15362);
nor U17558 (N_17558,N_14984,N_14566);
nor U17559 (N_17559,N_14889,N_15738);
xnor U17560 (N_17560,N_15863,N_15115);
or U17561 (N_17561,N_15011,N_14729);
xor U17562 (N_17562,N_14088,N_14732);
and U17563 (N_17563,N_15410,N_14001);
xnor U17564 (N_17564,N_14998,N_15203);
nand U17565 (N_17565,N_14805,N_15386);
nor U17566 (N_17566,N_15709,N_15035);
nor U17567 (N_17567,N_15826,N_14744);
or U17568 (N_17568,N_15638,N_15121);
nor U17569 (N_17569,N_15197,N_15283);
xor U17570 (N_17570,N_15319,N_15154);
nand U17571 (N_17571,N_14779,N_14360);
nand U17572 (N_17572,N_15650,N_14141);
xnor U17573 (N_17573,N_14620,N_15121);
and U17574 (N_17574,N_14094,N_15213);
nor U17575 (N_17575,N_15720,N_15200);
nor U17576 (N_17576,N_14404,N_15094);
xor U17577 (N_17577,N_14491,N_15896);
nor U17578 (N_17578,N_14530,N_15354);
and U17579 (N_17579,N_15183,N_15735);
xor U17580 (N_17580,N_15208,N_14157);
and U17581 (N_17581,N_15940,N_14557);
nand U17582 (N_17582,N_15083,N_15489);
or U17583 (N_17583,N_14977,N_15979);
nand U17584 (N_17584,N_14596,N_14602);
nor U17585 (N_17585,N_15088,N_14884);
nand U17586 (N_17586,N_15266,N_14770);
xnor U17587 (N_17587,N_14916,N_14622);
xnor U17588 (N_17588,N_15075,N_14477);
xnor U17589 (N_17589,N_14043,N_15675);
nand U17590 (N_17590,N_14366,N_15979);
or U17591 (N_17591,N_14930,N_14155);
or U17592 (N_17592,N_15091,N_14426);
nor U17593 (N_17593,N_14680,N_14496);
nand U17594 (N_17594,N_15121,N_15178);
and U17595 (N_17595,N_14789,N_14552);
and U17596 (N_17596,N_15037,N_15127);
and U17597 (N_17597,N_14089,N_15443);
xor U17598 (N_17598,N_15078,N_14616);
nor U17599 (N_17599,N_14665,N_14447);
xor U17600 (N_17600,N_14022,N_14665);
xnor U17601 (N_17601,N_15485,N_15697);
nor U17602 (N_17602,N_15004,N_15644);
nand U17603 (N_17603,N_15860,N_15402);
and U17604 (N_17604,N_14000,N_14503);
nor U17605 (N_17605,N_14179,N_15882);
or U17606 (N_17606,N_15310,N_14168);
xnor U17607 (N_17607,N_15602,N_14055);
and U17608 (N_17608,N_14964,N_15621);
nand U17609 (N_17609,N_15908,N_14001);
or U17610 (N_17610,N_14869,N_15067);
or U17611 (N_17611,N_14239,N_14598);
xnor U17612 (N_17612,N_15576,N_15928);
and U17613 (N_17613,N_15381,N_14269);
nor U17614 (N_17614,N_15255,N_14088);
nand U17615 (N_17615,N_14496,N_14893);
nor U17616 (N_17616,N_15462,N_14660);
nand U17617 (N_17617,N_14147,N_15461);
nor U17618 (N_17618,N_14310,N_15402);
or U17619 (N_17619,N_15130,N_14272);
and U17620 (N_17620,N_15830,N_15124);
and U17621 (N_17621,N_14712,N_14263);
nor U17622 (N_17622,N_14974,N_14061);
nor U17623 (N_17623,N_15844,N_15989);
nor U17624 (N_17624,N_15741,N_15333);
xnor U17625 (N_17625,N_14348,N_14890);
xor U17626 (N_17626,N_15786,N_14661);
or U17627 (N_17627,N_15857,N_14338);
xor U17628 (N_17628,N_15207,N_15300);
or U17629 (N_17629,N_14009,N_15320);
xnor U17630 (N_17630,N_14928,N_14816);
or U17631 (N_17631,N_15597,N_14528);
and U17632 (N_17632,N_14969,N_15918);
xor U17633 (N_17633,N_15826,N_14528);
xor U17634 (N_17634,N_14216,N_15491);
nand U17635 (N_17635,N_15109,N_14438);
nor U17636 (N_17636,N_14047,N_15615);
xor U17637 (N_17637,N_15211,N_14540);
nor U17638 (N_17638,N_14104,N_14813);
nand U17639 (N_17639,N_15485,N_14326);
nor U17640 (N_17640,N_15072,N_14423);
or U17641 (N_17641,N_15230,N_14966);
nand U17642 (N_17642,N_14142,N_15552);
nor U17643 (N_17643,N_15535,N_14759);
or U17644 (N_17644,N_14044,N_15244);
and U17645 (N_17645,N_14038,N_15289);
xnor U17646 (N_17646,N_15296,N_14535);
nor U17647 (N_17647,N_15361,N_15600);
nand U17648 (N_17648,N_15398,N_14578);
and U17649 (N_17649,N_14843,N_15038);
or U17650 (N_17650,N_14075,N_14649);
nor U17651 (N_17651,N_14219,N_15830);
and U17652 (N_17652,N_15832,N_14417);
or U17653 (N_17653,N_15146,N_15966);
xor U17654 (N_17654,N_14065,N_15424);
xnor U17655 (N_17655,N_14309,N_15008);
xor U17656 (N_17656,N_15698,N_14583);
and U17657 (N_17657,N_14689,N_15153);
or U17658 (N_17658,N_15143,N_15553);
nor U17659 (N_17659,N_14323,N_15819);
or U17660 (N_17660,N_14032,N_14195);
nor U17661 (N_17661,N_15024,N_15370);
and U17662 (N_17662,N_15476,N_15271);
or U17663 (N_17663,N_14428,N_14500);
and U17664 (N_17664,N_14663,N_15738);
and U17665 (N_17665,N_15166,N_15989);
nand U17666 (N_17666,N_14930,N_15284);
or U17667 (N_17667,N_15456,N_14031);
nor U17668 (N_17668,N_14868,N_15357);
xnor U17669 (N_17669,N_14706,N_15210);
or U17670 (N_17670,N_14971,N_14383);
xor U17671 (N_17671,N_14322,N_14876);
and U17672 (N_17672,N_14164,N_15148);
or U17673 (N_17673,N_15882,N_14299);
nor U17674 (N_17674,N_15950,N_15969);
nand U17675 (N_17675,N_14228,N_15140);
xnor U17676 (N_17676,N_15692,N_15439);
nor U17677 (N_17677,N_14706,N_15224);
and U17678 (N_17678,N_14023,N_14515);
xnor U17679 (N_17679,N_15854,N_14304);
xnor U17680 (N_17680,N_15528,N_15176);
and U17681 (N_17681,N_15222,N_15809);
xor U17682 (N_17682,N_14228,N_15003);
nand U17683 (N_17683,N_15975,N_14977);
xnor U17684 (N_17684,N_15244,N_14428);
or U17685 (N_17685,N_14461,N_14997);
xnor U17686 (N_17686,N_15088,N_15501);
nor U17687 (N_17687,N_15544,N_14494);
xor U17688 (N_17688,N_14742,N_14746);
xor U17689 (N_17689,N_14743,N_15719);
xnor U17690 (N_17690,N_15959,N_15026);
and U17691 (N_17691,N_14594,N_15431);
and U17692 (N_17692,N_15986,N_15425);
and U17693 (N_17693,N_14150,N_14326);
xnor U17694 (N_17694,N_15569,N_14320);
and U17695 (N_17695,N_15912,N_14656);
and U17696 (N_17696,N_14048,N_15685);
nand U17697 (N_17697,N_14353,N_15744);
nor U17698 (N_17698,N_15238,N_14280);
xnor U17699 (N_17699,N_15019,N_15766);
nand U17700 (N_17700,N_14887,N_15282);
nand U17701 (N_17701,N_14030,N_15499);
xor U17702 (N_17702,N_15552,N_15370);
xor U17703 (N_17703,N_14910,N_14406);
nor U17704 (N_17704,N_14352,N_14222);
xnor U17705 (N_17705,N_14207,N_14722);
and U17706 (N_17706,N_15035,N_14630);
xor U17707 (N_17707,N_15404,N_14963);
xnor U17708 (N_17708,N_14364,N_15113);
and U17709 (N_17709,N_14354,N_15006);
xor U17710 (N_17710,N_15598,N_14447);
nor U17711 (N_17711,N_14608,N_15173);
nand U17712 (N_17712,N_15259,N_14414);
xnor U17713 (N_17713,N_14654,N_15471);
or U17714 (N_17714,N_15653,N_14283);
nand U17715 (N_17715,N_15802,N_15346);
nand U17716 (N_17716,N_15338,N_15370);
nand U17717 (N_17717,N_14511,N_15792);
nand U17718 (N_17718,N_14995,N_15675);
and U17719 (N_17719,N_14859,N_15522);
xnor U17720 (N_17720,N_14511,N_15992);
xor U17721 (N_17721,N_15282,N_14963);
nand U17722 (N_17722,N_14375,N_15229);
nor U17723 (N_17723,N_15538,N_15325);
xor U17724 (N_17724,N_15545,N_14747);
and U17725 (N_17725,N_14556,N_14152);
nand U17726 (N_17726,N_14309,N_14579);
nor U17727 (N_17727,N_14682,N_15591);
or U17728 (N_17728,N_14696,N_15383);
nor U17729 (N_17729,N_14629,N_14187);
xnor U17730 (N_17730,N_14540,N_15990);
and U17731 (N_17731,N_14605,N_15296);
nor U17732 (N_17732,N_15507,N_15805);
nor U17733 (N_17733,N_14444,N_14457);
xnor U17734 (N_17734,N_14909,N_15600);
and U17735 (N_17735,N_14830,N_14693);
xor U17736 (N_17736,N_14281,N_15507);
nor U17737 (N_17737,N_15672,N_15364);
or U17738 (N_17738,N_15554,N_14483);
xor U17739 (N_17739,N_14594,N_14183);
or U17740 (N_17740,N_14194,N_14348);
xnor U17741 (N_17741,N_14775,N_14369);
nand U17742 (N_17742,N_15496,N_15337);
xor U17743 (N_17743,N_14228,N_15205);
nand U17744 (N_17744,N_15377,N_15192);
nor U17745 (N_17745,N_14561,N_14244);
xor U17746 (N_17746,N_15560,N_14588);
and U17747 (N_17747,N_15306,N_14080);
and U17748 (N_17748,N_14443,N_14106);
or U17749 (N_17749,N_15627,N_15273);
and U17750 (N_17750,N_15415,N_15774);
or U17751 (N_17751,N_14543,N_14929);
xnor U17752 (N_17752,N_15330,N_15053);
or U17753 (N_17753,N_15485,N_15634);
xnor U17754 (N_17754,N_14980,N_14523);
nor U17755 (N_17755,N_15849,N_15485);
or U17756 (N_17756,N_15309,N_15900);
nand U17757 (N_17757,N_15818,N_14740);
or U17758 (N_17758,N_14803,N_15503);
and U17759 (N_17759,N_15671,N_15572);
xor U17760 (N_17760,N_14113,N_15909);
nor U17761 (N_17761,N_14310,N_15246);
nor U17762 (N_17762,N_15816,N_14108);
and U17763 (N_17763,N_15985,N_14782);
and U17764 (N_17764,N_14879,N_15844);
xnor U17765 (N_17765,N_15603,N_15987);
nand U17766 (N_17766,N_15958,N_14201);
nor U17767 (N_17767,N_14914,N_15080);
nand U17768 (N_17768,N_14833,N_14688);
nand U17769 (N_17769,N_15910,N_15355);
nand U17770 (N_17770,N_15920,N_14624);
and U17771 (N_17771,N_15634,N_15346);
nand U17772 (N_17772,N_14012,N_15646);
xnor U17773 (N_17773,N_14409,N_15876);
or U17774 (N_17774,N_14036,N_15971);
and U17775 (N_17775,N_15244,N_15830);
nor U17776 (N_17776,N_15413,N_14864);
nand U17777 (N_17777,N_15208,N_14975);
xnor U17778 (N_17778,N_14669,N_15666);
nor U17779 (N_17779,N_15221,N_14909);
xor U17780 (N_17780,N_14513,N_14128);
and U17781 (N_17781,N_15074,N_14887);
nor U17782 (N_17782,N_14351,N_14047);
or U17783 (N_17783,N_14257,N_15145);
nand U17784 (N_17784,N_15911,N_15687);
xor U17785 (N_17785,N_15473,N_14731);
nor U17786 (N_17786,N_15227,N_14679);
nand U17787 (N_17787,N_14696,N_15390);
or U17788 (N_17788,N_14880,N_15276);
or U17789 (N_17789,N_14010,N_15290);
and U17790 (N_17790,N_15417,N_14528);
nand U17791 (N_17791,N_15646,N_14285);
or U17792 (N_17792,N_14863,N_14240);
and U17793 (N_17793,N_14439,N_14849);
or U17794 (N_17794,N_15300,N_14322);
and U17795 (N_17795,N_14882,N_14097);
and U17796 (N_17796,N_14949,N_15691);
xnor U17797 (N_17797,N_14527,N_15908);
and U17798 (N_17798,N_14759,N_15406);
nand U17799 (N_17799,N_15613,N_14741);
nor U17800 (N_17800,N_15792,N_15825);
nor U17801 (N_17801,N_15013,N_14643);
or U17802 (N_17802,N_15631,N_15869);
nor U17803 (N_17803,N_14269,N_14561);
or U17804 (N_17804,N_14750,N_15022);
and U17805 (N_17805,N_15111,N_15703);
and U17806 (N_17806,N_14487,N_15055);
or U17807 (N_17807,N_14854,N_14354);
xnor U17808 (N_17808,N_14096,N_15542);
or U17809 (N_17809,N_15953,N_15692);
and U17810 (N_17810,N_15624,N_14242);
or U17811 (N_17811,N_14996,N_15240);
nand U17812 (N_17812,N_15896,N_14172);
nor U17813 (N_17813,N_14929,N_15335);
xor U17814 (N_17814,N_14757,N_14814);
nor U17815 (N_17815,N_14806,N_15664);
nand U17816 (N_17816,N_15506,N_14969);
nor U17817 (N_17817,N_15051,N_15714);
xor U17818 (N_17818,N_14657,N_14516);
xnor U17819 (N_17819,N_14907,N_15840);
nand U17820 (N_17820,N_14146,N_15161);
xor U17821 (N_17821,N_15289,N_15076);
xor U17822 (N_17822,N_14390,N_14938);
or U17823 (N_17823,N_15222,N_15595);
xor U17824 (N_17824,N_15582,N_14098);
xnor U17825 (N_17825,N_15207,N_15494);
xnor U17826 (N_17826,N_15413,N_14448);
or U17827 (N_17827,N_15501,N_14451);
nand U17828 (N_17828,N_15819,N_14411);
nand U17829 (N_17829,N_15832,N_14744);
xnor U17830 (N_17830,N_15911,N_15673);
xor U17831 (N_17831,N_14455,N_14020);
nand U17832 (N_17832,N_14681,N_15841);
or U17833 (N_17833,N_15377,N_15742);
and U17834 (N_17834,N_15513,N_14695);
and U17835 (N_17835,N_14049,N_14793);
nor U17836 (N_17836,N_14602,N_15448);
nand U17837 (N_17837,N_14311,N_15024);
and U17838 (N_17838,N_14093,N_14694);
nor U17839 (N_17839,N_15565,N_15171);
and U17840 (N_17840,N_15657,N_14634);
or U17841 (N_17841,N_14231,N_15725);
nand U17842 (N_17842,N_15455,N_15902);
or U17843 (N_17843,N_14236,N_14413);
and U17844 (N_17844,N_15378,N_14135);
nor U17845 (N_17845,N_15614,N_14412);
or U17846 (N_17846,N_15041,N_15959);
nand U17847 (N_17847,N_14360,N_14110);
or U17848 (N_17848,N_15493,N_14626);
or U17849 (N_17849,N_14621,N_15469);
and U17850 (N_17850,N_15375,N_15541);
and U17851 (N_17851,N_14994,N_14526);
nand U17852 (N_17852,N_14088,N_14965);
or U17853 (N_17853,N_14797,N_14452);
nand U17854 (N_17854,N_15818,N_15506);
xnor U17855 (N_17855,N_15238,N_14035);
xor U17856 (N_17856,N_14772,N_15160);
nand U17857 (N_17857,N_15748,N_15208);
xor U17858 (N_17858,N_15105,N_14557);
nor U17859 (N_17859,N_14754,N_15249);
nand U17860 (N_17860,N_14617,N_15025);
xnor U17861 (N_17861,N_15967,N_14311);
xor U17862 (N_17862,N_15775,N_14112);
or U17863 (N_17863,N_14190,N_14181);
or U17864 (N_17864,N_14786,N_15256);
nand U17865 (N_17865,N_15119,N_15954);
xnor U17866 (N_17866,N_14773,N_15606);
nand U17867 (N_17867,N_15604,N_14701);
or U17868 (N_17868,N_15233,N_14174);
and U17869 (N_17869,N_14162,N_14968);
nand U17870 (N_17870,N_15802,N_14053);
or U17871 (N_17871,N_15934,N_14081);
xor U17872 (N_17872,N_15229,N_15163);
nor U17873 (N_17873,N_15471,N_14432);
xor U17874 (N_17874,N_14208,N_15902);
or U17875 (N_17875,N_15020,N_14118);
xnor U17876 (N_17876,N_15474,N_14174);
nor U17877 (N_17877,N_14613,N_14672);
nand U17878 (N_17878,N_14804,N_15628);
nand U17879 (N_17879,N_14767,N_15199);
and U17880 (N_17880,N_15932,N_14092);
nand U17881 (N_17881,N_14231,N_14796);
nor U17882 (N_17882,N_14182,N_15357);
or U17883 (N_17883,N_14042,N_14741);
or U17884 (N_17884,N_14923,N_15678);
and U17885 (N_17885,N_14066,N_14560);
and U17886 (N_17886,N_14059,N_15690);
or U17887 (N_17887,N_15449,N_14712);
or U17888 (N_17888,N_15649,N_15929);
or U17889 (N_17889,N_14161,N_14778);
or U17890 (N_17890,N_15795,N_15176);
xnor U17891 (N_17891,N_15075,N_15458);
xor U17892 (N_17892,N_14025,N_14036);
or U17893 (N_17893,N_15991,N_15276);
nand U17894 (N_17894,N_15456,N_14950);
or U17895 (N_17895,N_15933,N_14633);
and U17896 (N_17896,N_15811,N_15109);
xnor U17897 (N_17897,N_14237,N_15154);
and U17898 (N_17898,N_15887,N_15371);
nand U17899 (N_17899,N_15066,N_14108);
xnor U17900 (N_17900,N_15157,N_14507);
xor U17901 (N_17901,N_15102,N_14640);
xnor U17902 (N_17902,N_15736,N_15115);
xor U17903 (N_17903,N_15194,N_15760);
and U17904 (N_17904,N_14829,N_15020);
nor U17905 (N_17905,N_14192,N_14319);
nand U17906 (N_17906,N_14670,N_15001);
xnor U17907 (N_17907,N_14725,N_14332);
xor U17908 (N_17908,N_15834,N_15972);
nor U17909 (N_17909,N_14952,N_14207);
or U17910 (N_17910,N_14019,N_14579);
nand U17911 (N_17911,N_14682,N_15540);
and U17912 (N_17912,N_15763,N_15037);
or U17913 (N_17913,N_14322,N_14154);
or U17914 (N_17914,N_14951,N_14314);
and U17915 (N_17915,N_14492,N_14505);
or U17916 (N_17916,N_15637,N_14966);
xnor U17917 (N_17917,N_14622,N_15357);
nor U17918 (N_17918,N_15517,N_15044);
nor U17919 (N_17919,N_15696,N_14922);
or U17920 (N_17920,N_15428,N_15626);
or U17921 (N_17921,N_15910,N_14556);
and U17922 (N_17922,N_15904,N_14500);
nand U17923 (N_17923,N_14586,N_14176);
nor U17924 (N_17924,N_15410,N_15702);
or U17925 (N_17925,N_14692,N_15521);
or U17926 (N_17926,N_15226,N_14540);
nand U17927 (N_17927,N_15883,N_15549);
or U17928 (N_17928,N_14759,N_14347);
or U17929 (N_17929,N_15770,N_15114);
or U17930 (N_17930,N_14328,N_14442);
nand U17931 (N_17931,N_14670,N_14268);
xnor U17932 (N_17932,N_14011,N_14389);
or U17933 (N_17933,N_15858,N_14658);
nor U17934 (N_17934,N_14084,N_15955);
and U17935 (N_17935,N_14423,N_14020);
and U17936 (N_17936,N_15892,N_15470);
and U17937 (N_17937,N_14431,N_14543);
xor U17938 (N_17938,N_15749,N_15809);
nand U17939 (N_17939,N_15827,N_14192);
nand U17940 (N_17940,N_14165,N_14463);
and U17941 (N_17941,N_14309,N_15726);
or U17942 (N_17942,N_15769,N_15445);
nand U17943 (N_17943,N_14790,N_14051);
xor U17944 (N_17944,N_15656,N_14653);
xor U17945 (N_17945,N_14102,N_15383);
xor U17946 (N_17946,N_14159,N_15120);
nor U17947 (N_17947,N_15257,N_14856);
or U17948 (N_17948,N_14407,N_15464);
nor U17949 (N_17949,N_14453,N_14579);
or U17950 (N_17950,N_14994,N_14150);
or U17951 (N_17951,N_15798,N_15965);
nor U17952 (N_17952,N_14977,N_15097);
or U17953 (N_17953,N_14764,N_15692);
and U17954 (N_17954,N_14260,N_14550);
nand U17955 (N_17955,N_14690,N_14521);
or U17956 (N_17956,N_14845,N_14015);
nand U17957 (N_17957,N_14564,N_14874);
and U17958 (N_17958,N_15155,N_15737);
nand U17959 (N_17959,N_14636,N_15473);
and U17960 (N_17960,N_14346,N_14826);
nor U17961 (N_17961,N_14640,N_15585);
and U17962 (N_17962,N_15164,N_14462);
xor U17963 (N_17963,N_15895,N_15262);
xnor U17964 (N_17964,N_15406,N_15254);
and U17965 (N_17965,N_15928,N_14532);
and U17966 (N_17966,N_15239,N_14384);
xnor U17967 (N_17967,N_14685,N_14557);
nor U17968 (N_17968,N_15017,N_14418);
nor U17969 (N_17969,N_15380,N_14725);
xnor U17970 (N_17970,N_15642,N_15297);
nand U17971 (N_17971,N_15236,N_15400);
and U17972 (N_17972,N_15560,N_15061);
xnor U17973 (N_17973,N_15411,N_14031);
nand U17974 (N_17974,N_15202,N_14833);
xnor U17975 (N_17975,N_15954,N_15446);
nand U17976 (N_17976,N_15727,N_14155);
xor U17977 (N_17977,N_15221,N_15313);
nor U17978 (N_17978,N_15664,N_15932);
nand U17979 (N_17979,N_14499,N_14565);
and U17980 (N_17980,N_14284,N_15751);
nor U17981 (N_17981,N_14459,N_14989);
or U17982 (N_17982,N_15316,N_15706);
or U17983 (N_17983,N_15943,N_14384);
nor U17984 (N_17984,N_15048,N_14081);
nand U17985 (N_17985,N_14335,N_14020);
or U17986 (N_17986,N_15741,N_14863);
nor U17987 (N_17987,N_15597,N_14592);
nor U17988 (N_17988,N_15479,N_15338);
nand U17989 (N_17989,N_15107,N_14070);
and U17990 (N_17990,N_15797,N_15685);
nor U17991 (N_17991,N_14523,N_15110);
nand U17992 (N_17992,N_14474,N_14272);
and U17993 (N_17993,N_15175,N_15929);
or U17994 (N_17994,N_15628,N_15949);
and U17995 (N_17995,N_15685,N_14071);
nand U17996 (N_17996,N_15467,N_15444);
or U17997 (N_17997,N_15973,N_15011);
and U17998 (N_17998,N_14097,N_15067);
or U17999 (N_17999,N_14885,N_14134);
nor U18000 (N_18000,N_16654,N_17609);
nand U18001 (N_18001,N_16304,N_17713);
nor U18002 (N_18002,N_16671,N_17048);
nor U18003 (N_18003,N_16232,N_16025);
nor U18004 (N_18004,N_16582,N_17465);
nor U18005 (N_18005,N_16114,N_17475);
nor U18006 (N_18006,N_17354,N_17917);
and U18007 (N_18007,N_17988,N_16925);
or U18008 (N_18008,N_17066,N_17258);
nor U18009 (N_18009,N_17247,N_16010);
or U18010 (N_18010,N_17709,N_17278);
and U18011 (N_18011,N_17968,N_16225);
xor U18012 (N_18012,N_16073,N_17766);
or U18013 (N_18013,N_17426,N_17922);
xor U18014 (N_18014,N_16665,N_16086);
xor U18015 (N_18015,N_17040,N_16013);
xnor U18016 (N_18016,N_16873,N_16329);
and U18017 (N_18017,N_17757,N_17277);
nor U18018 (N_18018,N_17820,N_17320);
or U18019 (N_18019,N_16126,N_16479);
xnor U18020 (N_18020,N_17152,N_17849);
nor U18021 (N_18021,N_17555,N_17305);
or U18022 (N_18022,N_16138,N_17297);
nand U18023 (N_18023,N_16029,N_16685);
xnor U18024 (N_18024,N_17747,N_17759);
and U18025 (N_18025,N_16402,N_16041);
or U18026 (N_18026,N_17754,N_16170);
nor U18027 (N_18027,N_17742,N_17474);
nor U18028 (N_18028,N_17301,N_16326);
xor U18029 (N_18029,N_16901,N_16717);
nor U18030 (N_18030,N_16031,N_16005);
nor U18031 (N_18031,N_16392,N_16442);
or U18032 (N_18032,N_17865,N_17964);
nor U18033 (N_18033,N_17983,N_16719);
nand U18034 (N_18034,N_16516,N_17955);
xnor U18035 (N_18035,N_17398,N_16739);
nand U18036 (N_18036,N_17150,N_16848);
nor U18037 (N_18037,N_16491,N_17827);
and U18038 (N_18038,N_16471,N_17892);
nand U18039 (N_18039,N_16103,N_16815);
xnor U18040 (N_18040,N_17839,N_17431);
or U18041 (N_18041,N_17346,N_17452);
nor U18042 (N_18042,N_17542,N_16911);
and U18043 (N_18043,N_17401,N_16905);
xor U18044 (N_18044,N_17296,N_17280);
nand U18045 (N_18045,N_17038,N_16722);
xor U18046 (N_18046,N_17109,N_17873);
nand U18047 (N_18047,N_17574,N_16494);
nor U18048 (N_18048,N_17114,N_16229);
nand U18049 (N_18049,N_16180,N_16607);
xnor U18050 (N_18050,N_17908,N_17439);
or U18051 (N_18051,N_16288,N_17343);
nand U18052 (N_18052,N_16732,N_16259);
or U18053 (N_18053,N_16865,N_17599);
xor U18054 (N_18054,N_16880,N_17731);
nand U18055 (N_18055,N_16369,N_17058);
and U18056 (N_18056,N_17110,N_17261);
xor U18057 (N_18057,N_17479,N_17721);
nor U18058 (N_18058,N_17868,N_17680);
nand U18059 (N_18059,N_17081,N_16861);
and U18060 (N_18060,N_16580,N_17722);
nand U18061 (N_18061,N_17852,N_17959);
or U18062 (N_18062,N_16661,N_16769);
and U18063 (N_18063,N_16330,N_16287);
or U18064 (N_18064,N_16548,N_16622);
and U18065 (N_18065,N_17992,N_16166);
nand U18066 (N_18066,N_16443,N_16712);
and U18067 (N_18067,N_17457,N_16129);
and U18068 (N_18068,N_17537,N_17386);
and U18069 (N_18069,N_17860,N_17590);
nor U18070 (N_18070,N_16211,N_17324);
xor U18071 (N_18071,N_17635,N_17604);
and U18072 (N_18072,N_16547,N_16459);
xnor U18073 (N_18073,N_16590,N_17553);
or U18074 (N_18074,N_16648,N_17944);
nand U18075 (N_18075,N_16813,N_16976);
nand U18076 (N_18076,N_17734,N_16894);
nand U18077 (N_18077,N_17226,N_16387);
xor U18078 (N_18078,N_17684,N_17823);
or U18079 (N_18079,N_16958,N_16988);
xnor U18080 (N_18080,N_17941,N_17801);
xor U18081 (N_18081,N_16178,N_17877);
xor U18082 (N_18082,N_16694,N_17685);
and U18083 (N_18083,N_17028,N_16595);
nand U18084 (N_18084,N_17142,N_17436);
nand U18085 (N_18085,N_16718,N_16787);
nor U18086 (N_18086,N_17990,N_17629);
nand U18087 (N_18087,N_16151,N_16361);
xor U18088 (N_18088,N_16250,N_16721);
nand U18089 (N_18089,N_16597,N_16726);
nand U18090 (N_18090,N_16461,N_17595);
and U18091 (N_18091,N_17210,N_17156);
or U18092 (N_18092,N_16521,N_16952);
and U18093 (N_18093,N_16946,N_16983);
or U18094 (N_18094,N_16798,N_16950);
nand U18095 (N_18095,N_17331,N_16682);
or U18096 (N_18096,N_17520,N_16155);
xor U18097 (N_18097,N_16856,N_17923);
and U18098 (N_18098,N_16673,N_17135);
nor U18099 (N_18099,N_16328,N_17172);
or U18100 (N_18100,N_17377,N_17087);
nand U18101 (N_18101,N_16055,N_17915);
nor U18102 (N_18102,N_16113,N_16408);
xor U18103 (N_18103,N_17121,N_16604);
and U18104 (N_18104,N_16131,N_17306);
and U18105 (N_18105,N_16761,N_17031);
or U18106 (N_18106,N_16574,N_17022);
and U18107 (N_18107,N_17503,N_16945);
xnor U18108 (N_18108,N_16543,N_16474);
or U18109 (N_18109,N_17390,N_17687);
xor U18110 (N_18110,N_16697,N_16603);
or U18111 (N_18111,N_17803,N_16062);
or U18112 (N_18112,N_17111,N_16209);
xnor U18113 (N_18113,N_16744,N_16751);
or U18114 (N_18114,N_17429,N_16359);
nand U18115 (N_18115,N_17670,N_17032);
nand U18116 (N_18116,N_16450,N_16036);
xor U18117 (N_18117,N_16678,N_17522);
and U18118 (N_18118,N_17769,N_17833);
or U18119 (N_18119,N_16478,N_16281);
nand U18120 (N_18120,N_16220,N_17067);
nand U18121 (N_18121,N_16885,N_16285);
or U18122 (N_18122,N_17207,N_17554);
xnor U18123 (N_18123,N_17189,N_17191);
nor U18124 (N_18124,N_17487,N_16421);
or U18125 (N_18125,N_16923,N_16121);
nand U18126 (N_18126,N_17259,N_16143);
nand U18127 (N_18127,N_17034,N_17441);
and U18128 (N_18128,N_16072,N_16572);
and U18129 (N_18129,N_17644,N_17395);
nand U18130 (N_18130,N_17420,N_16782);
or U18131 (N_18131,N_16137,N_17989);
nor U18132 (N_18132,N_16818,N_16406);
xnor U18133 (N_18133,N_17242,N_17184);
or U18134 (N_18134,N_17244,N_17593);
xnor U18135 (N_18135,N_16438,N_16404);
and U18136 (N_18136,N_17530,N_16579);
or U18137 (N_18137,N_17003,N_16650);
or U18138 (N_18138,N_16437,N_16323);
or U18139 (N_18139,N_16305,N_16752);
nor U18140 (N_18140,N_17693,N_16422);
and U18141 (N_18141,N_17101,N_17788);
or U18142 (N_18142,N_16048,N_17037);
xnor U18143 (N_18143,N_16645,N_17541);
and U18144 (N_18144,N_17107,N_16506);
nand U18145 (N_18145,N_17671,N_17389);
and U18146 (N_18146,N_17136,N_17634);
nand U18147 (N_18147,N_17559,N_17625);
and U18148 (N_18148,N_16104,N_16948);
and U18149 (N_18149,N_17473,N_17737);
nand U18150 (N_18150,N_17516,N_16705);
xnor U18151 (N_18151,N_16997,N_16168);
nand U18152 (N_18152,N_16327,N_17043);
or U18153 (N_18153,N_16240,N_16069);
nand U18154 (N_18154,N_17815,N_16102);
xor U18155 (N_18155,N_17977,N_17648);
and U18156 (N_18156,N_16568,N_17112);
and U18157 (N_18157,N_17914,N_17491);
or U18158 (N_18158,N_16325,N_16979);
and U18159 (N_18159,N_17026,N_17500);
xor U18160 (N_18160,N_17761,N_16020);
and U18161 (N_18161,N_16293,N_17981);
and U18162 (N_18162,N_16337,N_17238);
nor U18163 (N_18163,N_17570,N_16345);
nor U18164 (N_18164,N_17164,N_16354);
xor U18165 (N_18165,N_16156,N_17883);
xor U18166 (N_18166,N_17578,N_16630);
xnor U18167 (N_18167,N_17281,N_17073);
or U18168 (N_18168,N_16116,N_17646);
xor U18169 (N_18169,N_16004,N_17698);
or U18170 (N_18170,N_16897,N_17196);
xor U18171 (N_18171,N_17518,N_17738);
or U18172 (N_18172,N_16162,N_17148);
or U18173 (N_18173,N_17750,N_17367);
or U18174 (N_18174,N_16331,N_17504);
or U18175 (N_18175,N_16247,N_16098);
xor U18176 (N_18176,N_17682,N_17155);
and U18177 (N_18177,N_16206,N_17997);
xnor U18178 (N_18178,N_17539,N_17468);
xor U18179 (N_18179,N_16655,N_16517);
nand U18180 (N_18180,N_17422,N_16540);
and U18181 (N_18181,N_17811,N_17963);
nor U18182 (N_18182,N_16870,N_16356);
nor U18183 (N_18183,N_16056,N_17300);
nand U18184 (N_18184,N_16881,N_16236);
and U18185 (N_18185,N_17779,N_17912);
or U18186 (N_18186,N_16231,N_17361);
and U18187 (N_18187,N_17176,N_16944);
nand U18188 (N_18188,N_17817,N_17802);
xnor U18189 (N_18189,N_17456,N_16342);
nor U18190 (N_18190,N_17869,N_16941);
nand U18191 (N_18191,N_17115,N_17130);
xnor U18192 (N_18192,N_16388,N_17837);
xor U18193 (N_18193,N_17621,N_16627);
nand U18194 (N_18194,N_17460,N_16068);
nand U18195 (N_18195,N_17239,N_16064);
or U18196 (N_18196,N_17834,N_17579);
or U18197 (N_18197,N_17774,N_16199);
xnor U18198 (N_18198,N_16451,N_16188);
xor U18199 (N_18199,N_17167,N_17064);
nor U18200 (N_18200,N_16039,N_17919);
nand U18201 (N_18201,N_16079,N_17667);
nor U18202 (N_18202,N_16564,N_16306);
nand U18203 (N_18203,N_17001,N_16044);
and U18204 (N_18204,N_17544,N_17220);
and U18205 (N_18205,N_16315,N_16115);
nor U18206 (N_18206,N_17700,N_17360);
nor U18207 (N_18207,N_16393,N_16176);
nand U18208 (N_18208,N_16576,N_16688);
nor U18209 (N_18209,N_17146,N_16942);
and U18210 (N_18210,N_16686,N_17939);
or U18211 (N_18211,N_17985,N_17848);
and U18212 (N_18212,N_16775,N_16303);
and U18213 (N_18213,N_17724,N_16350);
nand U18214 (N_18214,N_16740,N_17495);
or U18215 (N_18215,N_16058,N_17723);
and U18216 (N_18216,N_16184,N_16186);
and U18217 (N_18217,N_17074,N_16418);
xor U18218 (N_18218,N_17257,N_17949);
and U18219 (N_18219,N_16872,N_16360);
nand U18220 (N_18220,N_16358,N_17248);
nand U18221 (N_18221,N_17708,N_17119);
xor U18222 (N_18222,N_16571,N_17316);
nand U18223 (N_18223,N_17783,N_17195);
nor U18224 (N_18224,N_17661,N_16009);
or U18225 (N_18225,N_16123,N_17462);
and U18226 (N_18226,N_17828,N_17996);
and U18227 (N_18227,N_16581,N_16081);
or U18228 (N_18228,N_16675,N_17020);
nand U18229 (N_18229,N_17190,N_16251);
and U18230 (N_18230,N_17746,N_16801);
nand U18231 (N_18231,N_16618,N_17569);
and U18232 (N_18232,N_17694,N_17232);
or U18233 (N_18233,N_16641,N_17274);
nor U18234 (N_18234,N_16222,N_17973);
and U18235 (N_18235,N_16710,N_16702);
nor U18236 (N_18236,N_16898,N_16253);
or U18237 (N_18237,N_16525,N_16531);
nor U18238 (N_18238,N_16299,N_17986);
nand U18239 (N_18239,N_16120,N_16140);
nand U18240 (N_18240,N_17870,N_16614);
and U18241 (N_18241,N_17911,N_16819);
nand U18242 (N_18242,N_16834,N_16057);
nor U18243 (N_18243,N_17753,N_16218);
nor U18244 (N_18244,N_16959,N_17225);
xnor U18245 (N_18245,N_16753,N_16776);
or U18246 (N_18246,N_17933,N_17088);
nand U18247 (N_18247,N_17572,N_17206);
nand U18248 (N_18248,N_17467,N_17851);
xnor U18249 (N_18249,N_16527,N_16864);
and U18250 (N_18250,N_17607,N_16984);
xnor U18251 (N_18251,N_17931,N_17733);
and U18252 (N_18252,N_16669,N_17960);
and U18253 (N_18253,N_16532,N_17421);
nand U18254 (N_18254,N_16965,N_17948);
and U18255 (N_18255,N_16727,N_17231);
and U18256 (N_18256,N_16747,N_16953);
nand U18257 (N_18257,N_16700,N_17805);
nor U18258 (N_18258,N_17652,N_16074);
or U18259 (N_18259,N_16492,N_16847);
xor U18260 (N_18260,N_17089,N_16758);
and U18261 (N_18261,N_16239,N_17565);
nor U18262 (N_18262,N_17645,N_17012);
and U18263 (N_18263,N_16185,N_16110);
xnor U18264 (N_18264,N_16987,N_16106);
and U18265 (N_18265,N_16275,N_16508);
xnor U18266 (N_18266,N_16605,N_16080);
nor U18267 (N_18267,N_16460,N_17104);
and U18268 (N_18268,N_16366,N_16533);
or U18269 (N_18269,N_16696,N_17854);
nand U18270 (N_18270,N_17194,N_17942);
nor U18271 (N_18271,N_17351,N_17606);
or U18272 (N_18272,N_17924,N_16854);
nor U18273 (N_18273,N_17042,N_17732);
xor U18274 (N_18274,N_17276,N_17615);
nor U18275 (N_18275,N_16664,N_17647);
nor U18276 (N_18276,N_17719,N_16241);
xor U18277 (N_18277,N_17438,N_16951);
xor U18278 (N_18278,N_16071,N_17419);
xor U18279 (N_18279,N_16542,N_17643);
nor U18280 (N_18280,N_17245,N_17434);
nor U18281 (N_18281,N_16875,N_17295);
xor U18282 (N_18282,N_17617,N_17131);
xor U18283 (N_18283,N_17273,N_17529);
nand U18284 (N_18284,N_16411,N_17054);
nand U18285 (N_18285,N_17303,N_17889);
nand U18286 (N_18286,N_17366,N_17707);
nor U18287 (N_18287,N_16528,N_16981);
nand U18288 (N_18288,N_16197,N_16078);
nand U18289 (N_18289,N_16059,N_16820);
xnor U18290 (N_18290,N_16809,N_16016);
or U18291 (N_18291,N_17057,N_17484);
xor U18292 (N_18292,N_17430,N_16311);
xnor U18293 (N_18293,N_16196,N_17494);
nand U18294 (N_18294,N_16487,N_17106);
xor U18295 (N_18295,N_17006,N_16373);
or U18296 (N_18296,N_17151,N_16216);
or U18297 (N_18297,N_16619,N_17501);
nor U18298 (N_18298,N_16554,N_16998);
or U18299 (N_18299,N_17077,N_16558);
nor U18300 (N_18300,N_17459,N_17197);
and U18301 (N_18301,N_17029,N_17777);
nor U18302 (N_18302,N_17971,N_16573);
nor U18303 (N_18303,N_16376,N_17493);
and U18304 (N_18304,N_17138,N_17283);
xnor U18305 (N_18305,N_16280,N_16978);
and U18306 (N_18306,N_16108,N_16692);
nor U18307 (N_18307,N_16481,N_17214);
nand U18308 (N_18308,N_16006,N_17449);
nand U18309 (N_18309,N_16122,N_16458);
nand U18310 (N_18310,N_17512,N_16723);
and U18311 (N_18311,N_16884,N_17594);
nor U18312 (N_18312,N_17640,N_16507);
or U18313 (N_18313,N_16886,N_17177);
xor U18314 (N_18314,N_17143,N_17928);
nand U18315 (N_18315,N_16955,N_17192);
xor U18316 (N_18316,N_16523,N_16991);
xnor U18317 (N_18317,N_17790,N_17075);
nor U18318 (N_18318,N_17897,N_16101);
nor U18319 (N_18319,N_16264,N_17653);
nand U18320 (N_18320,N_17433,N_17978);
nand U18321 (N_18321,N_16125,N_17144);
xor U18322 (N_18322,N_17381,N_16628);
and U18323 (N_18323,N_17096,N_16099);
or U18324 (N_18324,N_17263,N_17443);
or U18325 (N_18325,N_17730,N_17383);
nor U18326 (N_18326,N_17266,N_17061);
nor U18327 (N_18327,N_16386,N_17881);
and U18328 (N_18328,N_16050,N_17342);
nand U18329 (N_18329,N_17329,N_16846);
nor U18330 (N_18330,N_17937,N_16845);
or U18331 (N_18331,N_16172,N_16545);
xnor U18332 (N_18332,N_17370,N_16445);
nor U18333 (N_18333,N_16907,N_16670);
nor U18334 (N_18334,N_16483,N_16498);
nand U18335 (N_18335,N_16157,N_17841);
and U18336 (N_18336,N_17764,N_17650);
and U18337 (N_18337,N_17781,N_16804);
nand U18338 (N_18338,N_17352,N_17410);
and U18339 (N_18339,N_17053,N_17677);
nor U18340 (N_18340,N_16488,N_16183);
or U18341 (N_18341,N_16428,N_16967);
nor U18342 (N_18342,N_16158,N_17587);
nand U18343 (N_18343,N_16254,N_17365);
and U18344 (N_18344,N_16038,N_16606);
nand U18345 (N_18345,N_16903,N_17952);
nand U18346 (N_18346,N_16466,N_17450);
and U18347 (N_18347,N_17536,N_17548);
nor U18348 (N_18348,N_17271,N_17378);
and U18349 (N_18349,N_16947,N_16943);
and U18350 (N_18350,N_16267,N_16118);
and U18351 (N_18351,N_16175,N_16772);
xor U18352 (N_18352,N_16189,N_17666);
nand U18353 (N_18353,N_17962,N_16312);
and U18354 (N_18354,N_17349,N_17379);
nor U18355 (N_18355,N_17065,N_17186);
and U18356 (N_18356,N_17691,N_17129);
nor U18357 (N_18357,N_16524,N_16193);
nor U18358 (N_18358,N_16921,N_17336);
nor U18359 (N_18359,N_16720,N_17141);
or U18360 (N_18360,N_17710,N_17725);
xor U18361 (N_18361,N_17899,N_17086);
or U18362 (N_18362,N_16235,N_16883);
nor U18363 (N_18363,N_17432,N_16920);
xor U18364 (N_18364,N_17562,N_17773);
xnor U18365 (N_18365,N_17162,N_16889);
nand U18366 (N_18366,N_17230,N_17113);
and U18367 (N_18367,N_16035,N_16139);
or U18368 (N_18368,N_16154,N_16486);
nor U18369 (N_18369,N_16570,N_16840);
nor U18370 (N_18370,N_17662,N_17372);
nor U18371 (N_18371,N_17669,N_17592);
nand U18372 (N_18372,N_16960,N_16629);
nor U18373 (N_18373,N_17575,N_17183);
xnor U18374 (N_18374,N_16476,N_17918);
and U18375 (N_18375,N_16511,N_16770);
nor U18376 (N_18376,N_16403,N_17649);
or U18377 (N_18377,N_17886,N_17181);
or U18378 (N_18378,N_16832,N_17478);
and U18379 (N_18379,N_16412,N_16119);
xor U18380 (N_18380,N_17882,N_16565);
or U18381 (N_18381,N_16933,N_17798);
or U18382 (N_18382,N_17165,N_16419);
nand U18383 (N_18383,N_16851,N_17673);
and U18384 (N_18384,N_16456,N_16742);
and U18385 (N_18385,N_17319,N_17749);
nand U18386 (N_18386,N_17613,N_16938);
nand U18387 (N_18387,N_17385,N_17158);
or U18388 (N_18388,N_17123,N_16262);
xor U18389 (N_18389,N_16931,N_17880);
nor U18390 (N_18390,N_17464,N_17526);
and U18391 (N_18391,N_16844,N_16030);
and U18392 (N_18392,N_16900,N_16750);
or U18393 (N_18393,N_17313,N_17581);
xnor U18394 (N_18394,N_16741,N_17292);
xnor U18395 (N_18395,N_17356,N_16874);
xnor U18396 (N_18396,N_17591,N_16759);
xnor U18397 (N_18397,N_16260,N_16643);
and U18398 (N_18398,N_16384,N_17577);
xnor U18399 (N_18399,N_16668,N_16142);
and U18400 (N_18400,N_17561,N_17770);
nand U18401 (N_18401,N_16993,N_16462);
nor U18402 (N_18402,N_17134,N_17596);
nand U18403 (N_18403,N_16519,N_17808);
or U18404 (N_18404,N_16130,N_17741);
and U18405 (N_18405,N_16169,N_17315);
nor U18406 (N_18406,N_17894,N_16584);
nand U18407 (N_18407,N_16937,N_17913);
nor U18408 (N_18408,N_17476,N_17905);
or U18409 (N_18409,N_16245,N_16141);
nor U18410 (N_18410,N_16802,N_16490);
and U18411 (N_18411,N_17163,N_17090);
and U18412 (N_18412,N_16213,N_17954);
or U18413 (N_18413,N_17369,N_17523);
xnor U18414 (N_18414,N_17347,N_16765);
nand U18415 (N_18415,N_17446,N_17224);
nor U18416 (N_18416,N_17223,N_17085);
nand U18417 (N_18417,N_17496,N_17157);
nor U18418 (N_18418,N_17287,N_17407);
xnor U18419 (N_18419,N_16957,N_16313);
nor U18420 (N_18420,N_16555,N_16857);
and U18421 (N_18421,N_17619,N_16733);
nand U18422 (N_18422,N_16349,N_16939);
and U18423 (N_18423,N_17884,N_16660);
nor U18424 (N_18424,N_16616,N_16469);
or U18425 (N_18425,N_16263,N_16257);
nand U18426 (N_18426,N_16283,N_17819);
and U18427 (N_18427,N_16994,N_16647);
or U18428 (N_18428,N_16868,N_17227);
or U18429 (N_18429,N_16805,N_17515);
nand U18430 (N_18430,N_16755,N_16177);
or U18431 (N_18431,N_16270,N_16746);
nand U18432 (N_18432,N_16191,N_17782);
xor U18433 (N_18433,N_17252,N_16763);
xnor U18434 (N_18434,N_16018,N_16277);
nand U18435 (N_18435,N_17816,N_17327);
nor U18436 (N_18436,N_17282,N_16786);
and U18437 (N_18437,N_17208,N_16567);
nand U18438 (N_18438,N_16019,N_17584);
nand U18439 (N_18439,N_16014,N_17505);
nor U18440 (N_18440,N_16536,N_16888);
or U18441 (N_18441,N_17703,N_16502);
nand U18442 (N_18442,N_16633,N_17657);
or U18443 (N_18443,N_16017,N_16452);
or U18444 (N_18444,N_17175,N_16539);
nor U18445 (N_18445,N_17062,N_17004);
or U18446 (N_18446,N_17626,N_16708);
nor U18447 (N_18447,N_17100,N_16663);
nor U18448 (N_18448,N_16698,N_16207);
and U18449 (N_18449,N_16493,N_16788);
xnor U18450 (N_18450,N_16195,N_17551);
nand U18451 (N_18451,N_17250,N_17083);
or U18452 (N_18452,N_17404,N_17580);
or U18453 (N_18453,N_17744,N_16695);
nand U18454 (N_18454,N_17966,N_17907);
and U18455 (N_18455,N_16215,N_17974);
nor U18456 (N_18456,N_17217,N_17965);
nand U18457 (N_18457,N_16145,N_17084);
or U18458 (N_18458,N_17128,N_17133);
or U18459 (N_18459,N_16893,N_16147);
nand U18460 (N_18460,N_16002,N_17799);
xor U18461 (N_18461,N_16396,N_17235);
nor U18462 (N_18462,N_17867,N_16632);
and U18463 (N_18463,N_16745,N_16027);
nand U18464 (N_18464,N_17916,N_17831);
nor U18465 (N_18465,N_16500,N_16454);
nor U18466 (N_18466,N_17472,N_16954);
xnor U18467 (N_18467,N_16256,N_17448);
and U18468 (N_18468,N_16707,N_17205);
nor U18469 (N_18469,N_17818,N_17209);
nand U18470 (N_18470,N_16586,N_17758);
nor U18471 (N_18471,N_17307,N_17938);
and U18472 (N_18472,N_17170,N_16778);
xor U18473 (N_18473,N_16082,N_16310);
or U18474 (N_18474,N_17984,N_16766);
nor U18475 (N_18475,N_16588,N_16961);
xor U18476 (N_18476,N_17998,N_17469);
or U18477 (N_18477,N_16594,N_16427);
nand U18478 (N_18478,N_16296,N_17507);
and U18479 (N_18479,N_17118,N_17014);
nand U18480 (N_18480,N_17338,N_17784);
or U18481 (N_18481,N_16187,N_16160);
xor U18482 (N_18482,N_16985,N_16292);
and U18483 (N_18483,N_17076,N_16174);
nand U18484 (N_18484,N_16284,N_16111);
and U18485 (N_18485,N_17601,N_16405);
and U18486 (N_18486,N_17308,N_16441);
xnor U18487 (N_18487,N_17658,N_16909);
nor U18488 (N_18488,N_17863,N_16575);
or U18489 (N_18489,N_17154,N_16703);
or U18490 (N_18490,N_17987,N_16447);
and U18491 (N_18491,N_16715,N_17080);
nand U18492 (N_18492,N_16754,N_16912);
and U18493 (N_18493,N_17202,N_16076);
xnor U18494 (N_18494,N_17980,N_17806);
and U18495 (N_18495,N_17702,N_17480);
xor U18496 (N_18496,N_16871,N_16996);
and U18497 (N_18497,N_17408,N_17674);
or U18498 (N_18498,N_16690,N_16252);
or U18499 (N_18499,N_16192,N_16194);
nor U18500 (N_18500,N_17284,N_17182);
or U18501 (N_18501,N_16075,N_16658);
nor U18502 (N_18502,N_16796,N_16926);
and U18503 (N_18503,N_17760,N_17940);
nor U18504 (N_18504,N_16455,N_17236);
or U18505 (N_18505,N_16591,N_17906);
xor U18506 (N_18506,N_16242,N_16593);
nand U18507 (N_18507,N_16320,N_17326);
and U18508 (N_18508,N_16977,N_17005);
and U18509 (N_18509,N_16266,N_17814);
or U18510 (N_18510,N_17879,N_16522);
and U18511 (N_18511,N_16302,N_17910);
nor U18512 (N_18512,N_16652,N_17127);
or U18513 (N_18513,N_16223,N_16375);
nor U18514 (N_18514,N_17525,N_17967);
xnor U18515 (N_18515,N_17015,N_17023);
xnor U18516 (N_18516,N_16133,N_17427);
and U18517 (N_18517,N_17729,N_16598);
or U18518 (N_18518,N_16672,N_16843);
nor U18519 (N_18519,N_17102,N_17743);
and U18520 (N_18520,N_17835,N_16365);
or U18521 (N_18521,N_16915,N_16348);
or U18522 (N_18522,N_17027,N_17160);
or U18523 (N_18523,N_16297,N_17564);
xnor U18524 (N_18524,N_17030,N_16749);
and U18525 (N_18525,N_17812,N_16850);
nand U18526 (N_18526,N_16837,N_17387);
xor U18527 (N_18527,N_16096,N_16756);
or U18528 (N_18528,N_17116,N_17796);
nor U18529 (N_18529,N_16489,N_17639);
or U18530 (N_18530,N_17763,N_16105);
xnor U18531 (N_18531,N_17103,N_17829);
or U18532 (N_18532,N_16771,N_17598);
xor U18533 (N_18533,N_16608,N_17686);
xnor U18534 (N_18534,N_17246,N_16891);
nand U18535 (N_18535,N_16100,N_16866);
nand U18536 (N_18536,N_17728,N_17161);
xor U18537 (N_18537,N_17715,N_16910);
nor U18538 (N_18538,N_16968,N_16321);
and U18539 (N_18539,N_17251,N_16282);
nor U18540 (N_18540,N_17211,N_17382);
and U18541 (N_18541,N_16268,N_17762);
or U18542 (N_18542,N_17809,N_17891);
and U18543 (N_18543,N_16735,N_16876);
and U18544 (N_18544,N_17991,N_16693);
nor U18545 (N_18545,N_17011,N_16762);
or U18546 (N_18546,N_16171,N_17126);
xnor U18547 (N_18547,N_17392,N_16307);
xor U18548 (N_18548,N_17995,N_17333);
xnor U18549 (N_18549,N_17380,N_17363);
xnor U18550 (N_18550,N_17692,N_17335);
nor U18551 (N_18551,N_16117,N_17424);
nand U18552 (N_18552,N_17795,N_16877);
nand U18553 (N_18553,N_17871,N_17836);
xor U18554 (N_18554,N_16791,N_16612);
nand U18555 (N_18555,N_16482,N_17310);
xor U18556 (N_18556,N_17558,N_16779);
or U18557 (N_18557,N_16092,N_16730);
nor U18558 (N_18558,N_17149,N_17676);
xnor U18559 (N_18559,N_16731,N_17060);
or U18560 (N_18560,N_16557,N_16821);
nand U18561 (N_18561,N_16684,N_16040);
nand U18562 (N_18562,N_16007,N_17663);
or U18563 (N_18563,N_16496,N_17498);
nor U18564 (N_18564,N_16344,N_16265);
and U18565 (N_18565,N_17290,N_16269);
nor U18566 (N_18566,N_16635,N_16409);
and U18567 (N_18567,N_17399,N_17659);
nand U18568 (N_18568,N_17632,N_16463);
or U18569 (N_18569,N_17117,N_17376);
nand U18570 (N_18570,N_16714,N_16803);
nand U18571 (N_18571,N_16070,N_16806);
or U18572 (N_18572,N_17481,N_16914);
xnor U18573 (N_18573,N_17628,N_16047);
xor U18574 (N_18574,N_17999,N_16012);
xnor U18575 (N_18575,N_17550,N_16298);
and U18576 (N_18576,N_16999,N_17935);
or U18577 (N_18577,N_16975,N_17780);
or U18578 (N_18578,N_16091,N_17355);
nor U18579 (N_18579,N_16849,N_16852);
xor U18580 (N_18580,N_17405,N_17069);
xor U18581 (N_18581,N_16357,N_16934);
nand U18582 (N_18582,N_17243,N_17188);
or U18583 (N_18583,N_16980,N_16918);
and U18584 (N_18584,N_16217,N_16084);
or U18585 (N_18585,N_16309,N_16895);
nand U18586 (N_18586,N_17630,N_16966);
and U18587 (N_18587,N_17341,N_17887);
xor U18588 (N_18588,N_17052,N_17885);
and U18589 (N_18589,N_16725,N_16601);
and U18590 (N_18590,N_16308,N_17254);
nand U18591 (N_18591,N_17610,N_17374);
xnor U18592 (N_18592,N_17547,N_16853);
nor U18593 (N_18593,N_17400,N_17950);
or U18594 (N_18594,N_17902,N_17497);
or U18595 (N_18595,N_16767,N_16680);
and U18596 (N_18596,N_16995,N_16385);
and U18597 (N_18597,N_16415,N_16435);
xor U18598 (N_18598,N_17875,N_17234);
xnor U18599 (N_18599,N_16468,N_17678);
or U18600 (N_18600,N_17945,N_16797);
xor U18601 (N_18601,N_16046,N_17193);
nor U18602 (N_18602,N_16773,N_17024);
nor U18603 (N_18603,N_17679,N_17016);
nor U18604 (N_18604,N_17605,N_16526);
or U18605 (N_18605,N_16066,N_16514);
xor U18606 (N_18606,N_17139,N_17482);
or U18607 (N_18607,N_16034,N_16136);
nor U18608 (N_18608,N_17402,N_16738);
nand U18609 (N_18609,N_17901,N_17265);
or U18610 (N_18610,N_17825,N_17614);
and U18611 (N_18611,N_17690,N_16879);
nand U18612 (N_18612,N_16089,N_17711);
nand U18613 (N_18613,N_16674,N_16553);
nor U18614 (N_18614,N_17583,N_16613);
nand U18615 (N_18615,N_17786,N_17508);
xor U18616 (N_18616,N_16230,N_16833);
nand U18617 (N_18617,N_17093,N_16512);
and U18618 (N_18618,N_17262,N_17576);
xor U18619 (N_18619,N_16609,N_17603);
xnor U18620 (N_18620,N_16916,N_16317);
and U18621 (N_18621,N_17822,N_17975);
xor U18622 (N_18622,N_16808,N_17846);
or U18623 (N_18623,N_17357,N_16153);
nand U18624 (N_18624,N_16649,N_17055);
nand U18625 (N_18625,N_17442,N_16475);
xor U18626 (N_18626,N_16592,N_16351);
nand U18627 (N_18627,N_16182,N_16274);
xor U18628 (N_18628,N_16318,N_17824);
nand U18629 (N_18629,N_16394,N_17041);
nand U18630 (N_18630,N_16430,N_17332);
nor U18631 (N_18631,N_17411,N_17253);
nor U18632 (N_18632,N_16777,N_16656);
nand U18633 (N_18633,N_16286,N_16546);
xnor U18634 (N_18634,N_17221,N_16828);
and U18635 (N_18635,N_17344,N_16294);
nor U18636 (N_18636,N_16340,N_16343);
xnor U18637 (N_18637,N_17701,N_16426);
or U18638 (N_18638,N_16637,N_16332);
nand U18639 (N_18639,N_16538,N_17772);
or U18640 (N_18640,N_16127,N_17483);
xnor U18641 (N_18641,N_17321,N_17862);
and U18642 (N_18642,N_16061,N_16676);
nor U18643 (N_18643,N_16552,N_16503);
or U18644 (N_18644,N_16173,N_16589);
or U18645 (N_18645,N_16817,N_16052);
or U18646 (N_18646,N_16760,N_16908);
and U18647 (N_18647,N_17716,N_17364);
nor U18648 (N_18648,N_16513,N_16624);
xnor U18649 (N_18649,N_17531,N_16090);
nand U18650 (N_18650,N_17445,N_17477);
or U18651 (N_18651,N_16858,N_17009);
nor U18652 (N_18652,N_17859,N_16465);
or U18653 (N_18653,N_17409,N_16882);
nor U18654 (N_18654,N_16003,N_17855);
nor U18655 (N_18655,N_17826,N_17216);
nor U18656 (N_18656,N_16748,N_16233);
xnor U18657 (N_18657,N_16198,N_17654);
and U18658 (N_18658,N_16646,N_16962);
nand U18659 (N_18659,N_17035,N_17993);
nor U18660 (N_18660,N_16144,N_16862);
xor U18661 (N_18661,N_17789,N_16887);
nor U18662 (N_18662,N_17388,N_16221);
xnor U18663 (N_18663,N_17222,N_17309);
nor U18664 (N_18664,N_16276,N_16699);
xnor U18665 (N_18665,N_17545,N_16830);
nand U18666 (N_18666,N_16472,N_16577);
nand U18667 (N_18667,N_16501,N_17771);
or U18668 (N_18668,N_16109,N_17068);
xor U18669 (N_18669,N_17045,N_16550);
nand U18670 (N_18670,N_16210,N_17312);
and U18671 (N_18671,N_16799,N_17631);
and U18672 (N_18672,N_16370,N_17314);
or U18673 (N_18673,N_17437,N_17132);
or U18674 (N_18674,N_17519,N_17304);
nor U18675 (N_18675,N_17920,N_16431);
nand U18676 (N_18676,N_16831,N_17633);
and U18677 (N_18677,N_17864,N_17423);
or U18678 (N_18678,N_16397,N_17173);
xor U18679 (N_18679,N_16768,N_16860);
or U18680 (N_18680,N_17059,N_17269);
nor U18681 (N_18681,N_16341,N_17797);
nand U18682 (N_18682,N_17095,N_17078);
nor U18683 (N_18683,N_17008,N_17140);
or U18684 (N_18684,N_17898,N_17108);
nand U18685 (N_18685,N_16518,N_17396);
and U18686 (N_18686,N_16401,N_17137);
and U18687 (N_18687,N_17237,N_16319);
nor U18688 (N_18688,N_17435,N_17768);
xnor U18689 (N_18689,N_16781,N_16636);
or U18690 (N_18690,N_16687,N_16273);
nand U18691 (N_18691,N_16556,N_16509);
nor U18692 (N_18692,N_16378,N_17755);
xor U18693 (N_18693,N_16666,N_16432);
xor U18694 (N_18694,N_17838,N_17444);
nor U18695 (N_18695,N_17348,N_16410);
nor U18696 (N_18696,N_17925,N_16927);
and U18697 (N_18697,N_16204,N_17642);
and U18698 (N_18698,N_17417,N_17776);
nor U18699 (N_18699,N_16163,N_16023);
or U18700 (N_18700,N_17071,N_16214);
nor U18701 (N_18701,N_17455,N_17813);
and U18702 (N_18702,N_16161,N_16424);
and U18703 (N_18703,N_16970,N_17393);
or U18704 (N_18704,N_16611,N_17890);
or U18705 (N_18705,N_16737,N_17018);
nor U18706 (N_18706,N_16651,N_17740);
xnor U18707 (N_18707,N_17804,N_16085);
nor U18708 (N_18708,N_17120,N_17521);
xor U18709 (N_18709,N_17588,N_16149);
nand U18710 (N_18710,N_16505,N_17416);
nand U18711 (N_18711,N_16261,N_17976);
and U18712 (N_18712,N_16610,N_17286);
and U18713 (N_18713,N_16716,N_16416);
xor U18714 (N_18714,N_17874,N_16200);
or U18715 (N_18715,N_17791,N_17302);
xor U18716 (N_18716,N_16711,N_17672);
nor U18717 (N_18717,N_17453,N_16679);
or U18718 (N_18718,N_16659,N_16063);
and U18719 (N_18719,N_17735,N_17982);
xor U18720 (N_18720,N_16367,N_16549);
nand U18721 (N_18721,N_16578,N_16790);
nand U18722 (N_18722,N_16701,N_16022);
xnor U18723 (N_18723,N_16380,N_16347);
or U18724 (N_18724,N_17514,N_16436);
xnor U18725 (N_18725,N_16060,N_16255);
or U18726 (N_18726,N_16510,N_17492);
xor U18727 (N_18727,N_17794,N_16936);
and U18728 (N_18728,N_17036,N_17169);
nand U18729 (N_18729,N_17488,N_16067);
nand U18730 (N_18730,N_16992,N_16499);
or U18731 (N_18731,N_17159,N_16982);
nor U18732 (N_18732,N_17844,N_17021);
xor U18733 (N_18733,N_17895,N_16899);
xor U18734 (N_18734,N_16585,N_17375);
nand U18735 (N_18735,N_17291,N_16811);
nand U18736 (N_18736,N_17618,N_17656);
or U18737 (N_18737,N_16827,N_17204);
xnor U18738 (N_18738,N_17622,N_17543);
xnor U18739 (N_18739,N_17418,N_17517);
nor U18740 (N_18740,N_17705,N_16822);
nor U18741 (N_18741,N_16146,N_17178);
xor U18742 (N_18742,N_16935,N_16464);
nand U18743 (N_18743,N_17602,N_16420);
nor U18744 (N_18744,N_16932,N_17056);
nand U18745 (N_18745,N_16623,N_17489);
xor U18746 (N_18746,N_17858,N_17958);
nand U18747 (N_18747,N_16065,N_17272);
or U18748 (N_18748,N_17972,N_17706);
nand U18749 (N_18749,N_17063,N_17748);
xor U18750 (N_18750,N_16444,N_16053);
nor U18751 (N_18751,N_16795,N_17739);
nand U18752 (N_18752,N_17368,N_16338);
nand U18753 (N_18753,N_16537,N_17091);
xnor U18754 (N_18754,N_17888,N_16272);
and U18755 (N_18755,N_17311,N_16278);
or U18756 (N_18756,N_16634,N_16964);
xor U18757 (N_18757,N_16956,N_16681);
nor U18758 (N_18758,N_16704,N_16364);
nand U18759 (N_18759,N_17527,N_17775);
or U18760 (N_18760,N_16520,N_16800);
or U18761 (N_18761,N_17124,N_16368);
nor U18762 (N_18762,N_16203,N_16638);
and U18763 (N_18763,N_16774,N_16973);
xor U18764 (N_18764,N_17627,N_17185);
xor U18765 (N_18765,N_16477,N_16051);
or U18766 (N_18766,N_16642,N_17792);
or U18767 (N_18767,N_17403,N_16353);
or U18768 (N_18768,N_17260,N_16448);
xor U18769 (N_18769,N_16867,N_17549);
nor U18770 (N_18770,N_16045,N_17122);
nor U18771 (N_18771,N_17168,N_17334);
xnor U18772 (N_18772,N_16346,N_16201);
nor U18773 (N_18773,N_17299,N_17861);
nor U18774 (N_18774,N_16026,N_16390);
nand U18775 (N_18775,N_17540,N_16301);
nand U18776 (N_18776,N_17934,N_17007);
nand U18777 (N_18777,N_17451,N_16227);
nor U18778 (N_18778,N_16838,N_16566);
xnor U18779 (N_18779,N_17793,N_16620);
nor U18780 (N_18780,N_16322,N_16757);
nand U18781 (N_18781,N_16400,N_16824);
nor U18782 (N_18782,N_16208,N_16135);
or U18783 (N_18783,N_17270,N_16202);
or U18784 (N_18784,N_16249,N_17876);
xnor U18785 (N_18785,N_16399,N_17174);
xor U18786 (N_18786,N_17904,N_17688);
nor U18787 (N_18787,N_16495,N_17756);
nand U18788 (N_18788,N_16639,N_16024);
or U18789 (N_18789,N_17830,N_16713);
nor U18790 (N_18790,N_16001,N_16433);
or U18791 (N_18791,N_16917,N_17322);
and U18792 (N_18792,N_17612,N_17720);
nor U18793 (N_18793,N_16429,N_17072);
nor U18794 (N_18794,N_17125,N_17490);
nor U18795 (N_18795,N_16449,N_16246);
nand U18796 (N_18796,N_16279,N_17800);
xnor U18797 (N_18797,N_16334,N_17339);
xnor U18798 (N_18798,N_16087,N_16363);
and U18799 (N_18799,N_16544,N_17535);
or U18800 (N_18800,N_17994,N_17203);
xor U18801 (N_18801,N_17832,N_16371);
or U18802 (N_18802,N_16640,N_17179);
and U18803 (N_18803,N_17546,N_16825);
xor U18804 (N_18804,N_16869,N_16922);
or U18805 (N_18805,N_16839,N_17509);
or U18806 (N_18806,N_17415,N_16563);
nor U18807 (N_18807,N_16314,N_16562);
and U18808 (N_18808,N_17406,N_17358);
and U18809 (N_18809,N_16124,N_17533);
and U18810 (N_18810,N_17017,N_17199);
xnor U18811 (N_18811,N_16238,N_16599);
nand U18812 (N_18812,N_17099,N_17847);
or U18813 (N_18813,N_17608,N_17019);
or U18814 (N_18814,N_17552,N_16823);
nor U18815 (N_18815,N_17714,N_16906);
or U18816 (N_18816,N_16398,N_16602);
xnor U18817 (N_18817,N_16355,N_16497);
xor U18818 (N_18818,N_17200,N_17318);
nand U18819 (N_18819,N_16736,N_17414);
xor U18820 (N_18820,N_17471,N_17359);
xor U18821 (N_18821,N_17219,N_16667);
and U18822 (N_18822,N_17689,N_17736);
or U18823 (N_18823,N_17921,N_17664);
nor U18824 (N_18824,N_16890,N_16190);
nand U18825 (N_18825,N_17699,N_17767);
or U18826 (N_18826,N_17082,N_17936);
and U18827 (N_18827,N_16535,N_16407);
nand U18828 (N_18828,N_17857,N_17636);
and U18829 (N_18829,N_17499,N_16551);
nand U18830 (N_18830,N_17458,N_16855);
nor U18831 (N_18831,N_16088,N_16226);
nor U18832 (N_18832,N_16504,N_16243);
xor U18833 (N_18833,N_16336,N_16615);
nand U18834 (N_18834,N_16878,N_16764);
or U18835 (N_18835,N_16033,N_16896);
and U18836 (N_18836,N_16785,N_16352);
or U18837 (N_18837,N_17013,N_17105);
nand U18838 (N_18838,N_16440,N_16008);
and U18839 (N_18839,N_17616,N_17293);
and U18840 (N_18840,N_16814,N_16224);
nor U18841 (N_18841,N_17440,N_16784);
or U18842 (N_18842,N_16150,N_17956);
and U18843 (N_18843,N_17362,N_16244);
or U18844 (N_18844,N_17033,N_16289);
xor U18845 (N_18845,N_16382,N_16794);
nand U18846 (N_18846,N_17275,N_17166);
or U18847 (N_18847,N_17511,N_17092);
nor U18848 (N_18848,N_16094,N_16439);
nand U18849 (N_18849,N_16728,N_16587);
xnor U18850 (N_18850,N_17000,N_16028);
nand U18851 (N_18851,N_16095,N_16569);
or U18852 (N_18852,N_16011,N_17582);
xnor U18853 (N_18853,N_16729,N_17896);
nor U18854 (N_18854,N_17264,N_16485);
nand U18855 (N_18855,N_17751,N_17668);
xor U18856 (N_18856,N_16389,N_16295);
nor U18857 (N_18857,N_16159,N_17187);
xor U18858 (N_18858,N_16810,N_17413);
and U18859 (N_18859,N_17198,N_17373);
nor U18860 (N_18860,N_17218,N_16434);
or U18861 (N_18861,N_17842,N_17201);
nor U18862 (N_18862,N_16237,N_17556);
nor U18863 (N_18863,N_17586,N_16248);
and U18864 (N_18864,N_16617,N_16892);
nor U18865 (N_18865,N_16042,N_16689);
nor U18866 (N_18866,N_16626,N_17943);
or U18867 (N_18867,N_16316,N_16467);
nand U18868 (N_18868,N_17872,N_17094);
and U18869 (N_18869,N_17538,N_16940);
or U18870 (N_18870,N_16835,N_17425);
xor U18871 (N_18871,N_17624,N_16743);
nand U18872 (N_18872,N_17778,N_16596);
nor U18873 (N_18873,N_17845,N_17240);
and U18874 (N_18874,N_17900,N_16093);
and U18875 (N_18875,N_17145,N_17171);
nand U18876 (N_18876,N_16530,N_17298);
or U18877 (N_18877,N_16395,N_17325);
nor U18878 (N_18878,N_16423,N_16043);
or U18879 (N_18879,N_16683,N_16037);
or U18880 (N_18880,N_16859,N_16148);
and U18881 (N_18881,N_16205,N_17215);
and U18882 (N_18882,N_16706,N_16473);
nor U18883 (N_18883,N_16377,N_17285);
nand U18884 (N_18884,N_17428,N_16971);
nor U18885 (N_18885,N_17532,N_16128);
nor U18886 (N_18886,N_16258,N_17932);
nand U18887 (N_18887,N_17524,N_16807);
nor U18888 (N_18888,N_17821,N_17153);
nand U18889 (N_18889,N_17470,N_16015);
nand U18890 (N_18890,N_16339,N_16812);
nand U18891 (N_18891,N_17279,N_17961);
xnor U18892 (N_18892,N_17337,N_16112);
nand U18893 (N_18893,N_17726,N_17502);
and U18894 (N_18894,N_16561,N_17893);
nor U18895 (N_18895,N_17785,N_17212);
and U18896 (N_18896,N_16974,N_16379);
and U18897 (N_18897,N_17213,N_16734);
and U18898 (N_18898,N_17002,N_16453);
and U18899 (N_18899,N_17466,N_17294);
nor U18900 (N_18900,N_16924,N_16290);
and U18901 (N_18901,N_17249,N_17039);
or U18902 (N_18902,N_17787,N_17463);
nand U18903 (N_18903,N_16989,N_17765);
and U18904 (N_18904,N_16972,N_17391);
xor U18905 (N_18905,N_16333,N_16374);
nand U18906 (N_18906,N_16152,N_17340);
and U18907 (N_18907,N_16446,N_17571);
or U18908 (N_18908,N_16372,N_17704);
nand U18909 (N_18909,N_17047,N_17180);
and U18910 (N_18910,N_16417,N_17317);
nand U18911 (N_18911,N_17727,N_17485);
xor U18912 (N_18912,N_16657,N_17454);
and U18913 (N_18913,N_17745,N_16457);
nor U18914 (N_18914,N_17717,N_17147);
or U18915 (N_18915,N_17345,N_16625);
and U18916 (N_18916,N_17853,N_16032);
and U18917 (N_18917,N_17528,N_17079);
xor U18918 (N_18918,N_16816,N_17638);
and U18919 (N_18919,N_16783,N_16963);
nor U18920 (N_18920,N_16841,N_17665);
xor U18921 (N_18921,N_17049,N_17712);
xnor U18922 (N_18922,N_16470,N_17909);
and U18923 (N_18923,N_17025,N_16644);
nand U18924 (N_18924,N_16054,N_17255);
nand U18925 (N_18925,N_16021,N_16600);
nor U18926 (N_18926,N_17573,N_16083);
nor U18927 (N_18927,N_17856,N_17807);
nand U18928 (N_18928,N_16793,N_17695);
nand U18929 (N_18929,N_16653,N_17510);
xor U18930 (N_18930,N_16986,N_17840);
nor U18931 (N_18931,N_17098,N_16691);
and U18932 (N_18932,N_16863,N_16077);
nor U18933 (N_18933,N_17597,N_16836);
nand U18934 (N_18934,N_16271,N_17560);
nor U18935 (N_18935,N_17397,N_17566);
and U18936 (N_18936,N_17486,N_16631);
nor U18937 (N_18937,N_17568,N_17323);
xor U18938 (N_18938,N_17600,N_17946);
xnor U18939 (N_18939,N_17655,N_16362);
and U18940 (N_18940,N_17070,N_16621);
nor U18941 (N_18941,N_16391,N_17970);
nor U18942 (N_18942,N_17330,N_16930);
xor U18943 (N_18943,N_16949,N_16480);
nor U18944 (N_18944,N_16212,N_17044);
nor U18945 (N_18945,N_16534,N_17660);
xnor U18946 (N_18946,N_17611,N_16165);
nor U18947 (N_18947,N_17752,N_16132);
nand U18948 (N_18948,N_17585,N_16383);
nor U18949 (N_18949,N_17589,N_17930);
and U18950 (N_18950,N_16919,N_16724);
and U18951 (N_18951,N_17697,N_17563);
or U18952 (N_18952,N_17681,N_16425);
and U18953 (N_18953,N_16780,N_16913);
nor U18954 (N_18954,N_17843,N_16662);
nor U18955 (N_18955,N_17513,N_17947);
nand U18956 (N_18956,N_17637,N_16134);
and U18957 (N_18957,N_16902,N_17350);
or U18958 (N_18958,N_17718,N_17256);
nand U18959 (N_18959,N_16792,N_16300);
nand U18960 (N_18960,N_17969,N_16000);
or U18961 (N_18961,N_17289,N_16167);
nand U18962 (N_18962,N_16324,N_17384);
or U18963 (N_18963,N_16107,N_16829);
xnor U18964 (N_18964,N_16049,N_17951);
nor U18965 (N_18965,N_17696,N_17927);
nand U18966 (N_18966,N_17046,N_16335);
or U18967 (N_18967,N_17353,N_17267);
nand U18968 (N_18968,N_17641,N_17371);
or U18969 (N_18969,N_16842,N_16529);
nor U18970 (N_18970,N_17288,N_16928);
xnor U18971 (N_18971,N_17328,N_16515);
and U18972 (N_18972,N_17929,N_17903);
nor U18973 (N_18973,N_17979,N_16789);
nand U18974 (N_18974,N_17878,N_17651);
xnor U18975 (N_18975,N_17675,N_17447);
nor U18976 (N_18976,N_16826,N_17623);
nor U18977 (N_18977,N_17810,N_17268);
nor U18978 (N_18978,N_16929,N_17534);
nand U18979 (N_18979,N_17557,N_16164);
xnor U18980 (N_18980,N_17953,N_16484);
nor U18981 (N_18981,N_17050,N_17233);
nand U18982 (N_18982,N_16583,N_17683);
and U18983 (N_18983,N_16709,N_17097);
or U18984 (N_18984,N_17957,N_16541);
xnor U18985 (N_18985,N_17051,N_16381);
nor U18986 (N_18986,N_17926,N_16677);
xor U18987 (N_18987,N_17412,N_16990);
nand U18988 (N_18988,N_17010,N_17620);
or U18989 (N_18989,N_17229,N_16413);
xor U18990 (N_18990,N_16559,N_17461);
or U18991 (N_18991,N_16228,N_16560);
nand U18992 (N_18992,N_16969,N_17567);
nor U18993 (N_18993,N_16181,N_16097);
nor U18994 (N_18994,N_16219,N_17228);
and U18995 (N_18995,N_17506,N_16414);
nor U18996 (N_18996,N_17241,N_17394);
or U18997 (N_18997,N_16291,N_16904);
nor U18998 (N_18998,N_17866,N_16234);
or U18999 (N_18999,N_17850,N_16179);
and U19000 (N_19000,N_16387,N_17844);
or U19001 (N_19001,N_17801,N_17511);
nand U19002 (N_19002,N_16292,N_16113);
or U19003 (N_19003,N_16613,N_17628);
nand U19004 (N_19004,N_17874,N_17188);
nand U19005 (N_19005,N_16093,N_17222);
nor U19006 (N_19006,N_17348,N_16975);
or U19007 (N_19007,N_17727,N_16735);
or U19008 (N_19008,N_16139,N_16371);
nor U19009 (N_19009,N_17975,N_17664);
xnor U19010 (N_19010,N_16237,N_17639);
xor U19011 (N_19011,N_16286,N_17721);
nand U19012 (N_19012,N_17606,N_16841);
nor U19013 (N_19013,N_17393,N_17066);
xnor U19014 (N_19014,N_16016,N_17914);
or U19015 (N_19015,N_17327,N_16066);
and U19016 (N_19016,N_17595,N_16331);
nor U19017 (N_19017,N_16369,N_16154);
nand U19018 (N_19018,N_17276,N_17904);
or U19019 (N_19019,N_16946,N_17330);
nor U19020 (N_19020,N_16395,N_17262);
and U19021 (N_19021,N_16776,N_16155);
and U19022 (N_19022,N_17072,N_17732);
xor U19023 (N_19023,N_16176,N_17348);
nand U19024 (N_19024,N_16903,N_17755);
and U19025 (N_19025,N_17465,N_16310);
or U19026 (N_19026,N_17233,N_17725);
or U19027 (N_19027,N_16301,N_17228);
xnor U19028 (N_19028,N_17346,N_17831);
nor U19029 (N_19029,N_16953,N_17642);
nand U19030 (N_19030,N_16369,N_16800);
or U19031 (N_19031,N_16992,N_16058);
or U19032 (N_19032,N_16706,N_17494);
or U19033 (N_19033,N_17056,N_16989);
xor U19034 (N_19034,N_17087,N_16473);
or U19035 (N_19035,N_17889,N_16807);
and U19036 (N_19036,N_16135,N_17256);
or U19037 (N_19037,N_16657,N_17564);
and U19038 (N_19038,N_16687,N_17980);
xor U19039 (N_19039,N_16112,N_16887);
or U19040 (N_19040,N_16437,N_16849);
or U19041 (N_19041,N_16381,N_16066);
nand U19042 (N_19042,N_16291,N_16334);
xnor U19043 (N_19043,N_16984,N_16730);
or U19044 (N_19044,N_17922,N_16676);
xor U19045 (N_19045,N_17697,N_16737);
nor U19046 (N_19046,N_16879,N_17744);
xor U19047 (N_19047,N_17074,N_16891);
or U19048 (N_19048,N_16734,N_16433);
or U19049 (N_19049,N_17633,N_17575);
nand U19050 (N_19050,N_16858,N_17869);
nor U19051 (N_19051,N_16009,N_17137);
nand U19052 (N_19052,N_17830,N_17856);
xor U19053 (N_19053,N_16659,N_16349);
nor U19054 (N_19054,N_16456,N_17882);
or U19055 (N_19055,N_17218,N_16862);
and U19056 (N_19056,N_16760,N_16383);
or U19057 (N_19057,N_16222,N_16360);
nand U19058 (N_19058,N_17803,N_16045);
or U19059 (N_19059,N_16755,N_16479);
xnor U19060 (N_19060,N_17804,N_17062);
xnor U19061 (N_19061,N_16488,N_16075);
nand U19062 (N_19062,N_17120,N_17104);
or U19063 (N_19063,N_17310,N_16340);
and U19064 (N_19064,N_17145,N_16271);
nand U19065 (N_19065,N_16013,N_16852);
xor U19066 (N_19066,N_16531,N_17734);
xor U19067 (N_19067,N_16094,N_17395);
nor U19068 (N_19068,N_16413,N_16199);
xor U19069 (N_19069,N_16378,N_16158);
nor U19070 (N_19070,N_16027,N_16628);
and U19071 (N_19071,N_17923,N_17811);
nand U19072 (N_19072,N_16856,N_17526);
xnor U19073 (N_19073,N_17575,N_16764);
nand U19074 (N_19074,N_16124,N_16920);
and U19075 (N_19075,N_16417,N_17766);
and U19076 (N_19076,N_16468,N_17773);
and U19077 (N_19077,N_17065,N_16576);
nand U19078 (N_19078,N_17618,N_16494);
xor U19079 (N_19079,N_16476,N_16689);
nor U19080 (N_19080,N_16371,N_17857);
nand U19081 (N_19081,N_16088,N_16663);
and U19082 (N_19082,N_17655,N_16915);
nand U19083 (N_19083,N_17029,N_17637);
and U19084 (N_19084,N_16264,N_17078);
and U19085 (N_19085,N_16466,N_17852);
or U19086 (N_19086,N_17599,N_16564);
nor U19087 (N_19087,N_16576,N_16721);
nand U19088 (N_19088,N_17381,N_16076);
or U19089 (N_19089,N_17338,N_17926);
nor U19090 (N_19090,N_16995,N_17177);
or U19091 (N_19091,N_17582,N_16967);
nand U19092 (N_19092,N_17940,N_17006);
nor U19093 (N_19093,N_17154,N_17300);
and U19094 (N_19094,N_17895,N_16539);
and U19095 (N_19095,N_17107,N_17898);
nand U19096 (N_19096,N_16622,N_17475);
nand U19097 (N_19097,N_17027,N_16777);
nor U19098 (N_19098,N_16183,N_16050);
and U19099 (N_19099,N_16681,N_16393);
and U19100 (N_19100,N_17014,N_16529);
and U19101 (N_19101,N_16151,N_16902);
nand U19102 (N_19102,N_16413,N_16244);
or U19103 (N_19103,N_16563,N_17174);
and U19104 (N_19104,N_17135,N_16270);
or U19105 (N_19105,N_16861,N_17664);
and U19106 (N_19106,N_17945,N_16488);
xnor U19107 (N_19107,N_17893,N_16518);
and U19108 (N_19108,N_16108,N_16479);
nand U19109 (N_19109,N_16582,N_17407);
nand U19110 (N_19110,N_17930,N_17881);
and U19111 (N_19111,N_17114,N_16957);
nand U19112 (N_19112,N_17462,N_16888);
or U19113 (N_19113,N_17573,N_17592);
xnor U19114 (N_19114,N_16278,N_16374);
nor U19115 (N_19115,N_16279,N_17143);
and U19116 (N_19116,N_17851,N_17838);
and U19117 (N_19117,N_17422,N_17210);
xnor U19118 (N_19118,N_17736,N_16905);
and U19119 (N_19119,N_16837,N_16799);
xor U19120 (N_19120,N_16463,N_16903);
and U19121 (N_19121,N_17289,N_16017);
nand U19122 (N_19122,N_17313,N_16288);
xor U19123 (N_19123,N_17374,N_17582);
and U19124 (N_19124,N_16899,N_17139);
nor U19125 (N_19125,N_16880,N_17808);
xnor U19126 (N_19126,N_17843,N_16303);
nor U19127 (N_19127,N_16889,N_17148);
or U19128 (N_19128,N_17249,N_16659);
or U19129 (N_19129,N_17613,N_17468);
or U19130 (N_19130,N_16792,N_16659);
nor U19131 (N_19131,N_17865,N_16364);
xor U19132 (N_19132,N_17882,N_16796);
and U19133 (N_19133,N_17608,N_17537);
nor U19134 (N_19134,N_16353,N_16988);
and U19135 (N_19135,N_16556,N_17154);
nand U19136 (N_19136,N_17557,N_17169);
and U19137 (N_19137,N_17761,N_16878);
and U19138 (N_19138,N_16874,N_17131);
nor U19139 (N_19139,N_16844,N_16769);
nand U19140 (N_19140,N_17605,N_17091);
nand U19141 (N_19141,N_16780,N_16519);
and U19142 (N_19142,N_16610,N_17451);
nand U19143 (N_19143,N_17386,N_16952);
nor U19144 (N_19144,N_16569,N_17102);
or U19145 (N_19145,N_16076,N_16691);
nor U19146 (N_19146,N_17930,N_16432);
and U19147 (N_19147,N_16263,N_17136);
nor U19148 (N_19148,N_17632,N_17743);
xnor U19149 (N_19149,N_16144,N_16098);
or U19150 (N_19150,N_17431,N_16430);
or U19151 (N_19151,N_17422,N_17323);
nand U19152 (N_19152,N_17909,N_17699);
nand U19153 (N_19153,N_17586,N_17272);
and U19154 (N_19154,N_17410,N_17617);
or U19155 (N_19155,N_17048,N_16047);
or U19156 (N_19156,N_16773,N_16680);
or U19157 (N_19157,N_17385,N_17831);
and U19158 (N_19158,N_17787,N_16822);
nand U19159 (N_19159,N_16309,N_16407);
nor U19160 (N_19160,N_17031,N_16048);
or U19161 (N_19161,N_16706,N_17117);
nor U19162 (N_19162,N_17984,N_17010);
nor U19163 (N_19163,N_16442,N_17557);
or U19164 (N_19164,N_16760,N_17368);
nor U19165 (N_19165,N_17903,N_16116);
xnor U19166 (N_19166,N_17763,N_16077);
xor U19167 (N_19167,N_16582,N_17947);
xnor U19168 (N_19168,N_16812,N_16051);
and U19169 (N_19169,N_17615,N_16350);
or U19170 (N_19170,N_16303,N_16527);
or U19171 (N_19171,N_16842,N_17423);
nand U19172 (N_19172,N_17189,N_16903);
or U19173 (N_19173,N_16593,N_16955);
and U19174 (N_19174,N_16878,N_17174);
or U19175 (N_19175,N_16011,N_17310);
nor U19176 (N_19176,N_17089,N_17329);
xor U19177 (N_19177,N_17563,N_16798);
nor U19178 (N_19178,N_17860,N_17822);
and U19179 (N_19179,N_17797,N_16662);
and U19180 (N_19180,N_16941,N_17213);
nor U19181 (N_19181,N_16438,N_17818);
or U19182 (N_19182,N_17459,N_16525);
and U19183 (N_19183,N_17677,N_17020);
or U19184 (N_19184,N_16913,N_17614);
xnor U19185 (N_19185,N_16896,N_16232);
xnor U19186 (N_19186,N_17176,N_17128);
nor U19187 (N_19187,N_17716,N_17628);
or U19188 (N_19188,N_16942,N_16539);
nor U19189 (N_19189,N_16331,N_16911);
and U19190 (N_19190,N_17802,N_16950);
and U19191 (N_19191,N_16820,N_16445);
or U19192 (N_19192,N_17207,N_17462);
or U19193 (N_19193,N_16011,N_16249);
xor U19194 (N_19194,N_17542,N_16693);
or U19195 (N_19195,N_16463,N_17115);
nor U19196 (N_19196,N_17492,N_16440);
xnor U19197 (N_19197,N_17329,N_16435);
nor U19198 (N_19198,N_16944,N_17535);
xor U19199 (N_19199,N_17435,N_17214);
and U19200 (N_19200,N_16192,N_17855);
nor U19201 (N_19201,N_16967,N_17559);
nand U19202 (N_19202,N_17294,N_17586);
and U19203 (N_19203,N_17794,N_16631);
nor U19204 (N_19204,N_16335,N_16485);
nand U19205 (N_19205,N_16844,N_17442);
xor U19206 (N_19206,N_16636,N_17337);
nor U19207 (N_19207,N_17887,N_16651);
nor U19208 (N_19208,N_17392,N_17690);
nor U19209 (N_19209,N_17055,N_16153);
or U19210 (N_19210,N_16296,N_16659);
nor U19211 (N_19211,N_17957,N_17486);
or U19212 (N_19212,N_16497,N_16674);
and U19213 (N_19213,N_16013,N_16380);
nand U19214 (N_19214,N_16041,N_16518);
and U19215 (N_19215,N_17360,N_16906);
xnor U19216 (N_19216,N_17948,N_17920);
nand U19217 (N_19217,N_16773,N_16767);
xnor U19218 (N_19218,N_16581,N_16519);
and U19219 (N_19219,N_16862,N_16181);
nor U19220 (N_19220,N_17360,N_16627);
and U19221 (N_19221,N_16169,N_16105);
and U19222 (N_19222,N_16560,N_17295);
or U19223 (N_19223,N_17274,N_17381);
nand U19224 (N_19224,N_17899,N_16213);
nor U19225 (N_19225,N_17161,N_16683);
xor U19226 (N_19226,N_16364,N_16461);
xnor U19227 (N_19227,N_16293,N_16820);
xor U19228 (N_19228,N_17090,N_17444);
or U19229 (N_19229,N_17954,N_16135);
and U19230 (N_19230,N_17019,N_16319);
or U19231 (N_19231,N_16077,N_17727);
or U19232 (N_19232,N_16707,N_17799);
nand U19233 (N_19233,N_17146,N_16202);
and U19234 (N_19234,N_17961,N_17651);
or U19235 (N_19235,N_16008,N_17906);
nor U19236 (N_19236,N_17410,N_17418);
and U19237 (N_19237,N_16408,N_17883);
and U19238 (N_19238,N_17393,N_17175);
and U19239 (N_19239,N_17745,N_16829);
nand U19240 (N_19240,N_16164,N_16359);
or U19241 (N_19241,N_16657,N_17674);
and U19242 (N_19242,N_17389,N_17403);
xnor U19243 (N_19243,N_17256,N_16422);
and U19244 (N_19244,N_16382,N_17208);
and U19245 (N_19245,N_16088,N_16485);
or U19246 (N_19246,N_16961,N_16984);
nor U19247 (N_19247,N_17487,N_17853);
nand U19248 (N_19248,N_16241,N_17965);
nor U19249 (N_19249,N_16989,N_17510);
nor U19250 (N_19250,N_17401,N_16196);
nand U19251 (N_19251,N_17338,N_17374);
or U19252 (N_19252,N_16029,N_16596);
or U19253 (N_19253,N_16513,N_17815);
or U19254 (N_19254,N_16608,N_16146);
or U19255 (N_19255,N_17575,N_17103);
nor U19256 (N_19256,N_16549,N_16303);
or U19257 (N_19257,N_16347,N_16733);
and U19258 (N_19258,N_16601,N_17872);
and U19259 (N_19259,N_17298,N_16867);
nor U19260 (N_19260,N_16254,N_17460);
and U19261 (N_19261,N_17731,N_16773);
and U19262 (N_19262,N_16348,N_16188);
nand U19263 (N_19263,N_16551,N_17617);
nand U19264 (N_19264,N_17443,N_16634);
xor U19265 (N_19265,N_16791,N_17702);
nand U19266 (N_19266,N_17595,N_16587);
nor U19267 (N_19267,N_16404,N_16820);
and U19268 (N_19268,N_16224,N_16128);
nand U19269 (N_19269,N_17652,N_16536);
and U19270 (N_19270,N_16749,N_16998);
xor U19271 (N_19271,N_17808,N_16388);
nand U19272 (N_19272,N_17952,N_17651);
nand U19273 (N_19273,N_16023,N_17651);
or U19274 (N_19274,N_17457,N_17525);
xor U19275 (N_19275,N_17099,N_17891);
nand U19276 (N_19276,N_17982,N_16385);
or U19277 (N_19277,N_17138,N_17507);
nor U19278 (N_19278,N_16846,N_16932);
nand U19279 (N_19279,N_17928,N_17386);
nand U19280 (N_19280,N_17281,N_17195);
and U19281 (N_19281,N_17225,N_16112);
or U19282 (N_19282,N_17236,N_16147);
nand U19283 (N_19283,N_17398,N_17380);
xor U19284 (N_19284,N_16267,N_17285);
nand U19285 (N_19285,N_17624,N_17804);
and U19286 (N_19286,N_17909,N_17143);
nor U19287 (N_19287,N_16072,N_17965);
and U19288 (N_19288,N_17845,N_17555);
and U19289 (N_19289,N_16153,N_17405);
and U19290 (N_19290,N_16774,N_17299);
or U19291 (N_19291,N_17079,N_16271);
or U19292 (N_19292,N_16902,N_16682);
and U19293 (N_19293,N_16697,N_17715);
or U19294 (N_19294,N_17369,N_17556);
nand U19295 (N_19295,N_16307,N_17948);
nor U19296 (N_19296,N_16001,N_16571);
and U19297 (N_19297,N_17706,N_17388);
nand U19298 (N_19298,N_16841,N_17633);
xor U19299 (N_19299,N_16427,N_17411);
nor U19300 (N_19300,N_17721,N_17567);
nor U19301 (N_19301,N_17205,N_16567);
xor U19302 (N_19302,N_17689,N_17110);
xor U19303 (N_19303,N_17208,N_17517);
xor U19304 (N_19304,N_17080,N_16809);
nand U19305 (N_19305,N_17538,N_16509);
nor U19306 (N_19306,N_16988,N_17674);
or U19307 (N_19307,N_17877,N_16174);
xor U19308 (N_19308,N_16879,N_16561);
and U19309 (N_19309,N_17437,N_16567);
nor U19310 (N_19310,N_16312,N_16916);
nand U19311 (N_19311,N_16046,N_16146);
nor U19312 (N_19312,N_16552,N_17320);
or U19313 (N_19313,N_16648,N_16632);
nand U19314 (N_19314,N_17672,N_16707);
and U19315 (N_19315,N_17393,N_17106);
or U19316 (N_19316,N_16923,N_17431);
nand U19317 (N_19317,N_17810,N_17917);
xor U19318 (N_19318,N_17573,N_17376);
and U19319 (N_19319,N_17850,N_17631);
nor U19320 (N_19320,N_17468,N_17875);
xor U19321 (N_19321,N_16495,N_17782);
xor U19322 (N_19322,N_17783,N_16109);
xnor U19323 (N_19323,N_16407,N_16345);
xor U19324 (N_19324,N_17116,N_17595);
nor U19325 (N_19325,N_17058,N_16032);
nand U19326 (N_19326,N_17023,N_17609);
and U19327 (N_19327,N_17997,N_16797);
xor U19328 (N_19328,N_16358,N_17394);
and U19329 (N_19329,N_16564,N_17958);
xor U19330 (N_19330,N_17366,N_17046);
and U19331 (N_19331,N_17583,N_16128);
and U19332 (N_19332,N_17910,N_17019);
xor U19333 (N_19333,N_17959,N_16110);
and U19334 (N_19334,N_17602,N_16160);
and U19335 (N_19335,N_16572,N_16441);
or U19336 (N_19336,N_16229,N_17613);
xnor U19337 (N_19337,N_17795,N_16518);
nor U19338 (N_19338,N_16935,N_16332);
and U19339 (N_19339,N_16121,N_17104);
nand U19340 (N_19340,N_17656,N_16984);
nor U19341 (N_19341,N_17076,N_17734);
nand U19342 (N_19342,N_16308,N_17956);
or U19343 (N_19343,N_16910,N_17091);
nand U19344 (N_19344,N_17598,N_17576);
xnor U19345 (N_19345,N_17419,N_17083);
and U19346 (N_19346,N_16008,N_17127);
nand U19347 (N_19347,N_16027,N_16573);
xnor U19348 (N_19348,N_16240,N_17880);
xnor U19349 (N_19349,N_17277,N_17874);
or U19350 (N_19350,N_16346,N_16768);
nand U19351 (N_19351,N_16167,N_16740);
nor U19352 (N_19352,N_16245,N_16653);
nand U19353 (N_19353,N_16984,N_16126);
and U19354 (N_19354,N_16470,N_16089);
xor U19355 (N_19355,N_16962,N_16338);
or U19356 (N_19356,N_16418,N_17939);
or U19357 (N_19357,N_17030,N_17083);
nand U19358 (N_19358,N_17650,N_17860);
or U19359 (N_19359,N_17668,N_17081);
xor U19360 (N_19360,N_16365,N_17277);
or U19361 (N_19361,N_16972,N_16101);
or U19362 (N_19362,N_17333,N_16440);
xor U19363 (N_19363,N_17861,N_16535);
nand U19364 (N_19364,N_16189,N_16937);
nand U19365 (N_19365,N_17737,N_16355);
nand U19366 (N_19366,N_16751,N_16648);
nor U19367 (N_19367,N_17348,N_16117);
nor U19368 (N_19368,N_17723,N_17757);
or U19369 (N_19369,N_17238,N_17397);
nand U19370 (N_19370,N_16833,N_17123);
nand U19371 (N_19371,N_16924,N_16932);
nand U19372 (N_19372,N_17865,N_16357);
nand U19373 (N_19373,N_16307,N_16719);
nor U19374 (N_19374,N_17515,N_16307);
and U19375 (N_19375,N_17877,N_16302);
nor U19376 (N_19376,N_17080,N_16901);
or U19377 (N_19377,N_16236,N_16779);
or U19378 (N_19378,N_17864,N_17261);
xor U19379 (N_19379,N_17337,N_17487);
nand U19380 (N_19380,N_17323,N_16335);
xor U19381 (N_19381,N_16399,N_17345);
nand U19382 (N_19382,N_17768,N_16024);
nor U19383 (N_19383,N_17199,N_17702);
nor U19384 (N_19384,N_16602,N_17190);
nor U19385 (N_19385,N_17895,N_16650);
and U19386 (N_19386,N_17891,N_16678);
xnor U19387 (N_19387,N_17713,N_17064);
nor U19388 (N_19388,N_16111,N_16486);
nor U19389 (N_19389,N_16404,N_16358);
nor U19390 (N_19390,N_16617,N_16351);
nor U19391 (N_19391,N_16347,N_17709);
or U19392 (N_19392,N_17684,N_17770);
nand U19393 (N_19393,N_17953,N_17890);
nor U19394 (N_19394,N_16224,N_16591);
or U19395 (N_19395,N_17803,N_17569);
and U19396 (N_19396,N_16036,N_17807);
xor U19397 (N_19397,N_16494,N_17854);
xnor U19398 (N_19398,N_17652,N_16692);
nand U19399 (N_19399,N_17000,N_17009);
nor U19400 (N_19400,N_16387,N_16095);
xnor U19401 (N_19401,N_17686,N_16990);
and U19402 (N_19402,N_16473,N_17697);
or U19403 (N_19403,N_16939,N_17934);
xnor U19404 (N_19404,N_17606,N_17265);
or U19405 (N_19405,N_17587,N_16397);
nand U19406 (N_19406,N_17412,N_16897);
and U19407 (N_19407,N_16843,N_16157);
nand U19408 (N_19408,N_17135,N_16458);
or U19409 (N_19409,N_17582,N_16484);
xor U19410 (N_19410,N_17446,N_17922);
xor U19411 (N_19411,N_17266,N_17611);
or U19412 (N_19412,N_16406,N_17218);
and U19413 (N_19413,N_17642,N_16237);
and U19414 (N_19414,N_17607,N_16393);
or U19415 (N_19415,N_17112,N_17089);
and U19416 (N_19416,N_16906,N_17979);
nand U19417 (N_19417,N_17581,N_17894);
or U19418 (N_19418,N_16124,N_16718);
or U19419 (N_19419,N_17653,N_17420);
nand U19420 (N_19420,N_16768,N_16582);
and U19421 (N_19421,N_16924,N_17995);
xnor U19422 (N_19422,N_17809,N_16582);
nand U19423 (N_19423,N_16244,N_16118);
xor U19424 (N_19424,N_17372,N_17714);
nand U19425 (N_19425,N_16721,N_17531);
xnor U19426 (N_19426,N_17257,N_17292);
nand U19427 (N_19427,N_17260,N_17178);
xor U19428 (N_19428,N_16455,N_17430);
nor U19429 (N_19429,N_16802,N_17712);
and U19430 (N_19430,N_17138,N_17752);
and U19431 (N_19431,N_17024,N_16604);
nor U19432 (N_19432,N_17386,N_17851);
or U19433 (N_19433,N_16556,N_16339);
nand U19434 (N_19434,N_16140,N_16977);
nor U19435 (N_19435,N_16995,N_16787);
nand U19436 (N_19436,N_16788,N_17959);
xnor U19437 (N_19437,N_17416,N_17080);
or U19438 (N_19438,N_16865,N_17409);
or U19439 (N_19439,N_16198,N_16502);
and U19440 (N_19440,N_17633,N_16478);
nor U19441 (N_19441,N_16202,N_16438);
xor U19442 (N_19442,N_17575,N_16818);
or U19443 (N_19443,N_16436,N_17723);
nor U19444 (N_19444,N_17375,N_17671);
xor U19445 (N_19445,N_17164,N_16073);
nand U19446 (N_19446,N_16671,N_17215);
nand U19447 (N_19447,N_16160,N_17286);
xnor U19448 (N_19448,N_17678,N_16085);
xor U19449 (N_19449,N_17459,N_17084);
or U19450 (N_19450,N_16622,N_16554);
xor U19451 (N_19451,N_17366,N_16451);
and U19452 (N_19452,N_16189,N_16106);
or U19453 (N_19453,N_17919,N_16106);
xor U19454 (N_19454,N_17659,N_17069);
or U19455 (N_19455,N_16651,N_17737);
or U19456 (N_19456,N_16492,N_16876);
or U19457 (N_19457,N_16897,N_16599);
nand U19458 (N_19458,N_17169,N_17810);
nor U19459 (N_19459,N_17056,N_16213);
or U19460 (N_19460,N_16976,N_16031);
nor U19461 (N_19461,N_17076,N_17354);
nand U19462 (N_19462,N_16103,N_17425);
or U19463 (N_19463,N_16962,N_17536);
and U19464 (N_19464,N_17878,N_17604);
and U19465 (N_19465,N_16582,N_17394);
xnor U19466 (N_19466,N_16491,N_17037);
or U19467 (N_19467,N_16055,N_17419);
nor U19468 (N_19468,N_16532,N_17748);
nor U19469 (N_19469,N_17441,N_17956);
xnor U19470 (N_19470,N_16803,N_17286);
xor U19471 (N_19471,N_17398,N_16534);
nand U19472 (N_19472,N_16879,N_16988);
xnor U19473 (N_19473,N_17553,N_16648);
nor U19474 (N_19474,N_17115,N_17802);
nor U19475 (N_19475,N_17204,N_16159);
and U19476 (N_19476,N_17109,N_16541);
xor U19477 (N_19477,N_17038,N_17941);
nand U19478 (N_19478,N_16968,N_17232);
nand U19479 (N_19479,N_17878,N_17150);
or U19480 (N_19480,N_16920,N_16912);
nor U19481 (N_19481,N_16865,N_17663);
xor U19482 (N_19482,N_16981,N_16853);
or U19483 (N_19483,N_16175,N_17494);
xnor U19484 (N_19484,N_17004,N_17397);
nor U19485 (N_19485,N_17423,N_17799);
nor U19486 (N_19486,N_16110,N_16287);
or U19487 (N_19487,N_16876,N_16992);
nor U19488 (N_19488,N_16654,N_16726);
xor U19489 (N_19489,N_16917,N_16561);
xor U19490 (N_19490,N_17909,N_16870);
nor U19491 (N_19491,N_17398,N_17096);
and U19492 (N_19492,N_16677,N_17521);
nand U19493 (N_19493,N_16783,N_16448);
xnor U19494 (N_19494,N_16391,N_16573);
nand U19495 (N_19495,N_16365,N_16764);
and U19496 (N_19496,N_16240,N_16557);
xnor U19497 (N_19497,N_17380,N_17358);
nand U19498 (N_19498,N_17437,N_16147);
nor U19499 (N_19499,N_16746,N_16548);
or U19500 (N_19500,N_16544,N_16044);
nor U19501 (N_19501,N_16635,N_17869);
and U19502 (N_19502,N_17714,N_17208);
and U19503 (N_19503,N_17388,N_16839);
nor U19504 (N_19504,N_17343,N_17060);
or U19505 (N_19505,N_17772,N_16122);
nand U19506 (N_19506,N_17245,N_17099);
nand U19507 (N_19507,N_16366,N_17522);
nand U19508 (N_19508,N_16598,N_16209);
nand U19509 (N_19509,N_16156,N_17722);
or U19510 (N_19510,N_16959,N_17929);
and U19511 (N_19511,N_17665,N_17451);
xor U19512 (N_19512,N_16475,N_17942);
xor U19513 (N_19513,N_16853,N_17432);
xnor U19514 (N_19514,N_16387,N_16825);
xor U19515 (N_19515,N_16797,N_16088);
or U19516 (N_19516,N_17381,N_16467);
or U19517 (N_19517,N_16737,N_17126);
xor U19518 (N_19518,N_16488,N_16596);
or U19519 (N_19519,N_17951,N_16427);
xnor U19520 (N_19520,N_17972,N_17997);
xnor U19521 (N_19521,N_16712,N_17534);
nand U19522 (N_19522,N_16708,N_16229);
nand U19523 (N_19523,N_16157,N_16534);
nor U19524 (N_19524,N_17269,N_17425);
nand U19525 (N_19525,N_16985,N_17736);
nand U19526 (N_19526,N_17418,N_16388);
nand U19527 (N_19527,N_16159,N_17032);
xor U19528 (N_19528,N_17101,N_17747);
nand U19529 (N_19529,N_16692,N_16097);
nand U19530 (N_19530,N_17644,N_16461);
nand U19531 (N_19531,N_17852,N_16911);
nand U19532 (N_19532,N_16152,N_16925);
nand U19533 (N_19533,N_16827,N_16123);
and U19534 (N_19534,N_17150,N_16288);
and U19535 (N_19535,N_17317,N_16173);
or U19536 (N_19536,N_16130,N_16538);
or U19537 (N_19537,N_16138,N_16459);
xor U19538 (N_19538,N_17527,N_17433);
or U19539 (N_19539,N_16027,N_16020);
and U19540 (N_19540,N_16031,N_16370);
nor U19541 (N_19541,N_16172,N_16687);
nor U19542 (N_19542,N_16209,N_16163);
nor U19543 (N_19543,N_16383,N_17469);
or U19544 (N_19544,N_17496,N_16667);
and U19545 (N_19545,N_16059,N_17353);
and U19546 (N_19546,N_16265,N_16496);
or U19547 (N_19547,N_17818,N_17361);
nor U19548 (N_19548,N_16666,N_17728);
xor U19549 (N_19549,N_17947,N_16342);
or U19550 (N_19550,N_17906,N_17670);
and U19551 (N_19551,N_16748,N_17453);
or U19552 (N_19552,N_16361,N_17906);
or U19553 (N_19553,N_17094,N_17935);
nor U19554 (N_19554,N_17655,N_17477);
xnor U19555 (N_19555,N_17341,N_17486);
or U19556 (N_19556,N_17234,N_17320);
and U19557 (N_19557,N_17394,N_17897);
and U19558 (N_19558,N_17318,N_17881);
and U19559 (N_19559,N_16380,N_17977);
and U19560 (N_19560,N_16839,N_17549);
nor U19561 (N_19561,N_17456,N_17175);
nor U19562 (N_19562,N_16279,N_16286);
xor U19563 (N_19563,N_17606,N_16436);
xor U19564 (N_19564,N_16639,N_17436);
nand U19565 (N_19565,N_16307,N_17490);
and U19566 (N_19566,N_16381,N_17186);
nor U19567 (N_19567,N_17073,N_17420);
nand U19568 (N_19568,N_17381,N_16566);
nor U19569 (N_19569,N_16335,N_16087);
or U19570 (N_19570,N_17159,N_16175);
nor U19571 (N_19571,N_16560,N_17136);
and U19572 (N_19572,N_16318,N_16634);
nand U19573 (N_19573,N_16578,N_16011);
and U19574 (N_19574,N_16348,N_16130);
or U19575 (N_19575,N_16423,N_17678);
or U19576 (N_19576,N_17880,N_16584);
nor U19577 (N_19577,N_17425,N_16905);
or U19578 (N_19578,N_17129,N_17606);
or U19579 (N_19579,N_17039,N_16729);
xor U19580 (N_19580,N_16285,N_17153);
and U19581 (N_19581,N_17543,N_17369);
and U19582 (N_19582,N_16010,N_16332);
nor U19583 (N_19583,N_17273,N_16342);
nand U19584 (N_19584,N_16046,N_16686);
xor U19585 (N_19585,N_16864,N_16429);
nor U19586 (N_19586,N_16321,N_16374);
xnor U19587 (N_19587,N_17489,N_17991);
xor U19588 (N_19588,N_16631,N_17789);
nor U19589 (N_19589,N_17208,N_17399);
and U19590 (N_19590,N_17339,N_16897);
xor U19591 (N_19591,N_17175,N_17849);
xor U19592 (N_19592,N_16879,N_17215);
xnor U19593 (N_19593,N_16246,N_17445);
nand U19594 (N_19594,N_17735,N_16790);
nor U19595 (N_19595,N_17533,N_17357);
xor U19596 (N_19596,N_16818,N_17778);
xor U19597 (N_19597,N_16307,N_16418);
or U19598 (N_19598,N_17015,N_17146);
xnor U19599 (N_19599,N_16282,N_17811);
or U19600 (N_19600,N_16996,N_16026);
and U19601 (N_19601,N_16547,N_17890);
xor U19602 (N_19602,N_17677,N_17743);
or U19603 (N_19603,N_17147,N_17352);
xnor U19604 (N_19604,N_16137,N_16368);
xnor U19605 (N_19605,N_16085,N_17569);
nor U19606 (N_19606,N_16945,N_17111);
nor U19607 (N_19607,N_17409,N_17090);
and U19608 (N_19608,N_17495,N_16679);
xnor U19609 (N_19609,N_16320,N_16433);
nor U19610 (N_19610,N_16297,N_16137);
xor U19611 (N_19611,N_16696,N_16305);
xnor U19612 (N_19612,N_16605,N_16446);
and U19613 (N_19613,N_16402,N_16812);
nand U19614 (N_19614,N_16740,N_16927);
and U19615 (N_19615,N_16594,N_17511);
xnor U19616 (N_19616,N_17769,N_16570);
nand U19617 (N_19617,N_17433,N_16899);
nor U19618 (N_19618,N_17901,N_16798);
xor U19619 (N_19619,N_16298,N_16260);
or U19620 (N_19620,N_16438,N_16397);
or U19621 (N_19621,N_17049,N_16045);
and U19622 (N_19622,N_16486,N_17883);
nor U19623 (N_19623,N_16609,N_17777);
nand U19624 (N_19624,N_16206,N_16675);
and U19625 (N_19625,N_17759,N_16406);
or U19626 (N_19626,N_17631,N_16646);
nand U19627 (N_19627,N_16789,N_17157);
or U19628 (N_19628,N_17572,N_17962);
or U19629 (N_19629,N_17284,N_17210);
nor U19630 (N_19630,N_17373,N_17947);
or U19631 (N_19631,N_17613,N_16787);
or U19632 (N_19632,N_17125,N_16955);
or U19633 (N_19633,N_17094,N_17881);
and U19634 (N_19634,N_16176,N_17278);
nor U19635 (N_19635,N_16620,N_16163);
nand U19636 (N_19636,N_17736,N_17732);
nand U19637 (N_19637,N_17795,N_17523);
xnor U19638 (N_19638,N_16215,N_16496);
nor U19639 (N_19639,N_16193,N_16939);
nand U19640 (N_19640,N_17016,N_17756);
nand U19641 (N_19641,N_16320,N_16996);
xnor U19642 (N_19642,N_17947,N_17786);
or U19643 (N_19643,N_17113,N_17526);
nor U19644 (N_19644,N_16577,N_17252);
nand U19645 (N_19645,N_16228,N_17486);
or U19646 (N_19646,N_17598,N_17522);
nor U19647 (N_19647,N_16685,N_17882);
or U19648 (N_19648,N_16877,N_17436);
nand U19649 (N_19649,N_17142,N_17633);
and U19650 (N_19650,N_17755,N_17117);
nand U19651 (N_19651,N_17427,N_17185);
and U19652 (N_19652,N_17642,N_17671);
xnor U19653 (N_19653,N_17463,N_17437);
and U19654 (N_19654,N_16109,N_16486);
nand U19655 (N_19655,N_17601,N_16995);
and U19656 (N_19656,N_16769,N_17045);
or U19657 (N_19657,N_17276,N_17968);
nor U19658 (N_19658,N_16308,N_16182);
nand U19659 (N_19659,N_16909,N_17068);
nand U19660 (N_19660,N_16936,N_16531);
nand U19661 (N_19661,N_17146,N_16989);
nand U19662 (N_19662,N_16475,N_17094);
and U19663 (N_19663,N_17617,N_16615);
or U19664 (N_19664,N_16359,N_16203);
nand U19665 (N_19665,N_17856,N_17132);
xnor U19666 (N_19666,N_17738,N_17496);
or U19667 (N_19667,N_17702,N_16710);
nor U19668 (N_19668,N_16844,N_16273);
nor U19669 (N_19669,N_16379,N_16227);
nor U19670 (N_19670,N_17877,N_17643);
nor U19671 (N_19671,N_17573,N_16458);
and U19672 (N_19672,N_17012,N_16112);
or U19673 (N_19673,N_17769,N_17707);
and U19674 (N_19674,N_16997,N_17313);
and U19675 (N_19675,N_17488,N_16065);
nor U19676 (N_19676,N_16471,N_17685);
xnor U19677 (N_19677,N_16893,N_16212);
nand U19678 (N_19678,N_17643,N_17473);
nand U19679 (N_19679,N_16921,N_17710);
or U19680 (N_19680,N_16655,N_17502);
xnor U19681 (N_19681,N_16658,N_16273);
nor U19682 (N_19682,N_16083,N_17848);
xnor U19683 (N_19683,N_17838,N_16611);
and U19684 (N_19684,N_17991,N_16317);
or U19685 (N_19685,N_17549,N_16715);
nand U19686 (N_19686,N_16080,N_17366);
xnor U19687 (N_19687,N_17538,N_16600);
xnor U19688 (N_19688,N_17427,N_17566);
xor U19689 (N_19689,N_17571,N_16908);
nor U19690 (N_19690,N_17737,N_16611);
xor U19691 (N_19691,N_16595,N_16480);
nand U19692 (N_19692,N_17806,N_16702);
xnor U19693 (N_19693,N_17398,N_17110);
nand U19694 (N_19694,N_17875,N_17377);
nor U19695 (N_19695,N_17364,N_17406);
nor U19696 (N_19696,N_16094,N_17403);
xnor U19697 (N_19697,N_16731,N_17199);
nor U19698 (N_19698,N_16780,N_17904);
nand U19699 (N_19699,N_16963,N_16667);
nand U19700 (N_19700,N_16748,N_16282);
and U19701 (N_19701,N_17845,N_17962);
nor U19702 (N_19702,N_16465,N_16119);
or U19703 (N_19703,N_17503,N_17681);
or U19704 (N_19704,N_16531,N_16553);
nand U19705 (N_19705,N_16472,N_16759);
nand U19706 (N_19706,N_16812,N_16973);
or U19707 (N_19707,N_17157,N_16082);
nand U19708 (N_19708,N_17209,N_17495);
nor U19709 (N_19709,N_17852,N_17112);
nor U19710 (N_19710,N_16369,N_16105);
xnor U19711 (N_19711,N_16121,N_16342);
nor U19712 (N_19712,N_17891,N_17777);
or U19713 (N_19713,N_17433,N_17060);
xor U19714 (N_19714,N_16935,N_16555);
nand U19715 (N_19715,N_16884,N_17558);
nand U19716 (N_19716,N_16931,N_17624);
nor U19717 (N_19717,N_17690,N_16163);
and U19718 (N_19718,N_16149,N_17461);
xnor U19719 (N_19719,N_17194,N_17454);
nand U19720 (N_19720,N_16328,N_17440);
and U19721 (N_19721,N_16546,N_16014);
nand U19722 (N_19722,N_16211,N_17765);
and U19723 (N_19723,N_16770,N_16055);
or U19724 (N_19724,N_16625,N_16957);
xor U19725 (N_19725,N_17294,N_16725);
or U19726 (N_19726,N_17395,N_17783);
nor U19727 (N_19727,N_17904,N_17593);
or U19728 (N_19728,N_16142,N_16755);
nand U19729 (N_19729,N_16697,N_17791);
nor U19730 (N_19730,N_16781,N_16135);
nor U19731 (N_19731,N_17088,N_16117);
nor U19732 (N_19732,N_16219,N_16186);
or U19733 (N_19733,N_16641,N_17545);
nor U19734 (N_19734,N_17369,N_16204);
nand U19735 (N_19735,N_17182,N_17323);
xnor U19736 (N_19736,N_16301,N_16247);
and U19737 (N_19737,N_17540,N_16114);
nor U19738 (N_19738,N_16298,N_17212);
or U19739 (N_19739,N_16269,N_17933);
and U19740 (N_19740,N_16350,N_17179);
and U19741 (N_19741,N_17208,N_17785);
and U19742 (N_19742,N_17958,N_17669);
xnor U19743 (N_19743,N_16974,N_16635);
and U19744 (N_19744,N_17927,N_17972);
and U19745 (N_19745,N_17087,N_16718);
or U19746 (N_19746,N_17852,N_16374);
xor U19747 (N_19747,N_16899,N_16670);
xnor U19748 (N_19748,N_17007,N_17714);
xor U19749 (N_19749,N_17857,N_17315);
nand U19750 (N_19750,N_17980,N_17136);
nor U19751 (N_19751,N_16296,N_16149);
xor U19752 (N_19752,N_16529,N_16154);
nor U19753 (N_19753,N_17185,N_17606);
nand U19754 (N_19754,N_17906,N_17325);
nor U19755 (N_19755,N_17417,N_16371);
or U19756 (N_19756,N_17995,N_16131);
and U19757 (N_19757,N_17370,N_17260);
nand U19758 (N_19758,N_17277,N_17945);
nand U19759 (N_19759,N_17312,N_17751);
and U19760 (N_19760,N_17392,N_17855);
and U19761 (N_19761,N_16710,N_17468);
or U19762 (N_19762,N_17260,N_17049);
nor U19763 (N_19763,N_17355,N_17803);
and U19764 (N_19764,N_16709,N_17362);
or U19765 (N_19765,N_17848,N_16104);
nor U19766 (N_19766,N_17550,N_17810);
or U19767 (N_19767,N_16444,N_16979);
nand U19768 (N_19768,N_16477,N_16974);
and U19769 (N_19769,N_16523,N_17189);
or U19770 (N_19770,N_16955,N_16911);
and U19771 (N_19771,N_16118,N_17243);
and U19772 (N_19772,N_17842,N_16664);
and U19773 (N_19773,N_16253,N_16332);
nor U19774 (N_19774,N_17161,N_17106);
xor U19775 (N_19775,N_16890,N_16615);
nor U19776 (N_19776,N_17425,N_17211);
or U19777 (N_19777,N_16671,N_16294);
nand U19778 (N_19778,N_16395,N_16891);
nand U19779 (N_19779,N_17648,N_16968);
nor U19780 (N_19780,N_16702,N_17543);
nor U19781 (N_19781,N_17248,N_16301);
xnor U19782 (N_19782,N_16113,N_17047);
xor U19783 (N_19783,N_17691,N_17554);
xor U19784 (N_19784,N_17486,N_16074);
nand U19785 (N_19785,N_17832,N_16604);
xnor U19786 (N_19786,N_16089,N_16771);
nand U19787 (N_19787,N_17972,N_16341);
and U19788 (N_19788,N_17872,N_16557);
or U19789 (N_19789,N_17910,N_17194);
xor U19790 (N_19790,N_16892,N_17108);
and U19791 (N_19791,N_17620,N_16388);
or U19792 (N_19792,N_16057,N_16656);
or U19793 (N_19793,N_16438,N_16542);
or U19794 (N_19794,N_16615,N_17711);
or U19795 (N_19795,N_17760,N_17044);
nand U19796 (N_19796,N_17679,N_16329);
and U19797 (N_19797,N_17498,N_16197);
or U19798 (N_19798,N_16451,N_16370);
and U19799 (N_19799,N_17829,N_17225);
nor U19800 (N_19800,N_16107,N_16952);
or U19801 (N_19801,N_16455,N_16690);
xor U19802 (N_19802,N_16621,N_16501);
nand U19803 (N_19803,N_16362,N_16946);
nand U19804 (N_19804,N_17003,N_16858);
and U19805 (N_19805,N_17208,N_16501);
nor U19806 (N_19806,N_17099,N_16833);
nand U19807 (N_19807,N_17947,N_16213);
or U19808 (N_19808,N_17625,N_17681);
nand U19809 (N_19809,N_17257,N_16889);
or U19810 (N_19810,N_17032,N_16684);
nand U19811 (N_19811,N_17297,N_16610);
nand U19812 (N_19812,N_17465,N_17167);
or U19813 (N_19813,N_16684,N_16630);
nand U19814 (N_19814,N_17879,N_16400);
xor U19815 (N_19815,N_16001,N_16354);
and U19816 (N_19816,N_17918,N_17244);
or U19817 (N_19817,N_16691,N_17978);
nor U19818 (N_19818,N_17272,N_17386);
xnor U19819 (N_19819,N_16403,N_17201);
xor U19820 (N_19820,N_17244,N_17386);
xor U19821 (N_19821,N_16194,N_16829);
or U19822 (N_19822,N_17104,N_16404);
xor U19823 (N_19823,N_16954,N_17254);
or U19824 (N_19824,N_17734,N_17338);
nor U19825 (N_19825,N_16699,N_16605);
xnor U19826 (N_19826,N_17207,N_17577);
nor U19827 (N_19827,N_17426,N_17892);
nand U19828 (N_19828,N_17037,N_16511);
or U19829 (N_19829,N_16985,N_16789);
nand U19830 (N_19830,N_16102,N_17592);
and U19831 (N_19831,N_16289,N_16366);
nor U19832 (N_19832,N_16956,N_17305);
and U19833 (N_19833,N_17912,N_17692);
nand U19834 (N_19834,N_17198,N_17158);
nor U19835 (N_19835,N_17676,N_16444);
and U19836 (N_19836,N_16776,N_16159);
xor U19837 (N_19837,N_16704,N_16429);
or U19838 (N_19838,N_17702,N_16298);
and U19839 (N_19839,N_16964,N_16986);
nor U19840 (N_19840,N_16195,N_17715);
and U19841 (N_19841,N_16732,N_17050);
xor U19842 (N_19842,N_17307,N_16253);
xor U19843 (N_19843,N_16180,N_17069);
or U19844 (N_19844,N_17772,N_17351);
or U19845 (N_19845,N_17741,N_17752);
and U19846 (N_19846,N_17336,N_16175);
or U19847 (N_19847,N_16493,N_16471);
or U19848 (N_19848,N_16798,N_17547);
and U19849 (N_19849,N_16916,N_16892);
nand U19850 (N_19850,N_16000,N_17037);
and U19851 (N_19851,N_16081,N_16332);
nand U19852 (N_19852,N_16532,N_16921);
and U19853 (N_19853,N_16518,N_17047);
xnor U19854 (N_19854,N_16846,N_16239);
or U19855 (N_19855,N_16872,N_16909);
nand U19856 (N_19856,N_17244,N_17322);
or U19857 (N_19857,N_16550,N_16512);
nand U19858 (N_19858,N_16465,N_16232);
nand U19859 (N_19859,N_17213,N_16093);
nor U19860 (N_19860,N_17417,N_17987);
or U19861 (N_19861,N_17761,N_16382);
xor U19862 (N_19862,N_16767,N_17316);
or U19863 (N_19863,N_16221,N_16209);
or U19864 (N_19864,N_17956,N_16304);
or U19865 (N_19865,N_17555,N_16078);
nand U19866 (N_19866,N_16657,N_17076);
and U19867 (N_19867,N_16572,N_17337);
or U19868 (N_19868,N_16110,N_17736);
nor U19869 (N_19869,N_17250,N_17364);
and U19870 (N_19870,N_16596,N_17943);
nand U19871 (N_19871,N_16667,N_17090);
and U19872 (N_19872,N_16905,N_16257);
or U19873 (N_19873,N_16464,N_17865);
and U19874 (N_19874,N_17079,N_17392);
nor U19875 (N_19875,N_17742,N_17303);
and U19876 (N_19876,N_17179,N_16371);
nor U19877 (N_19877,N_17978,N_17630);
xor U19878 (N_19878,N_17111,N_16421);
nor U19879 (N_19879,N_16850,N_17926);
or U19880 (N_19880,N_16227,N_17232);
nor U19881 (N_19881,N_17399,N_17033);
nor U19882 (N_19882,N_16972,N_17825);
xnor U19883 (N_19883,N_17939,N_17463);
or U19884 (N_19884,N_16706,N_17662);
nor U19885 (N_19885,N_17606,N_17371);
xnor U19886 (N_19886,N_17215,N_16524);
and U19887 (N_19887,N_16374,N_16461);
and U19888 (N_19888,N_16065,N_16371);
or U19889 (N_19889,N_17932,N_16312);
and U19890 (N_19890,N_16131,N_16632);
nand U19891 (N_19891,N_17165,N_16748);
xnor U19892 (N_19892,N_16866,N_16522);
nand U19893 (N_19893,N_17433,N_16126);
and U19894 (N_19894,N_16519,N_17170);
xnor U19895 (N_19895,N_16255,N_16372);
or U19896 (N_19896,N_16663,N_16189);
xor U19897 (N_19897,N_16003,N_16420);
xor U19898 (N_19898,N_17206,N_17403);
and U19899 (N_19899,N_17883,N_16139);
nand U19900 (N_19900,N_17314,N_16194);
nor U19901 (N_19901,N_16851,N_17273);
or U19902 (N_19902,N_16148,N_16215);
xor U19903 (N_19903,N_16305,N_16179);
xor U19904 (N_19904,N_17830,N_17375);
and U19905 (N_19905,N_17442,N_16572);
nor U19906 (N_19906,N_17336,N_17906);
and U19907 (N_19907,N_17746,N_16331);
nand U19908 (N_19908,N_17604,N_17886);
and U19909 (N_19909,N_16690,N_16229);
or U19910 (N_19910,N_16205,N_16006);
xor U19911 (N_19911,N_16833,N_16350);
xnor U19912 (N_19912,N_17144,N_16545);
or U19913 (N_19913,N_16781,N_17476);
or U19914 (N_19914,N_17250,N_16350);
and U19915 (N_19915,N_17271,N_16441);
xnor U19916 (N_19916,N_17727,N_17813);
nand U19917 (N_19917,N_16026,N_17781);
nor U19918 (N_19918,N_17529,N_16861);
xor U19919 (N_19919,N_16215,N_16274);
xnor U19920 (N_19920,N_17594,N_16809);
nor U19921 (N_19921,N_17924,N_17182);
and U19922 (N_19922,N_17767,N_17239);
and U19923 (N_19923,N_17313,N_16947);
or U19924 (N_19924,N_17661,N_16720);
nor U19925 (N_19925,N_17395,N_16886);
or U19926 (N_19926,N_17823,N_16939);
nand U19927 (N_19927,N_16548,N_16584);
xor U19928 (N_19928,N_17902,N_16293);
xnor U19929 (N_19929,N_17181,N_16909);
and U19930 (N_19930,N_17751,N_17519);
nor U19931 (N_19931,N_16569,N_17248);
nor U19932 (N_19932,N_17242,N_17794);
nand U19933 (N_19933,N_17463,N_17066);
and U19934 (N_19934,N_16744,N_17352);
xor U19935 (N_19935,N_16056,N_16036);
or U19936 (N_19936,N_17531,N_16937);
nor U19937 (N_19937,N_17817,N_17211);
or U19938 (N_19938,N_17312,N_17647);
or U19939 (N_19939,N_17211,N_17961);
or U19940 (N_19940,N_16288,N_17633);
and U19941 (N_19941,N_16576,N_17819);
xor U19942 (N_19942,N_17382,N_17379);
and U19943 (N_19943,N_16382,N_16724);
and U19944 (N_19944,N_16778,N_16478);
xnor U19945 (N_19945,N_17405,N_16341);
nand U19946 (N_19946,N_16885,N_17372);
nand U19947 (N_19947,N_17443,N_16667);
or U19948 (N_19948,N_17572,N_16910);
or U19949 (N_19949,N_16471,N_17333);
nand U19950 (N_19950,N_16112,N_16506);
nor U19951 (N_19951,N_16385,N_16730);
and U19952 (N_19952,N_16350,N_17172);
and U19953 (N_19953,N_16423,N_16984);
xor U19954 (N_19954,N_17287,N_17361);
nor U19955 (N_19955,N_16326,N_16422);
nand U19956 (N_19956,N_17333,N_16965);
or U19957 (N_19957,N_16563,N_17110);
and U19958 (N_19958,N_16151,N_16020);
and U19959 (N_19959,N_16587,N_17760);
or U19960 (N_19960,N_17910,N_16704);
nand U19961 (N_19961,N_16302,N_16324);
nand U19962 (N_19962,N_17547,N_16260);
nand U19963 (N_19963,N_17344,N_16992);
nor U19964 (N_19964,N_17757,N_16058);
xor U19965 (N_19965,N_16097,N_17015);
xor U19966 (N_19966,N_16027,N_16137);
nand U19967 (N_19967,N_17809,N_17589);
xnor U19968 (N_19968,N_17838,N_16722);
and U19969 (N_19969,N_16521,N_17373);
nor U19970 (N_19970,N_17233,N_16771);
xor U19971 (N_19971,N_17795,N_16981);
nor U19972 (N_19972,N_17124,N_16352);
and U19973 (N_19973,N_16024,N_17728);
and U19974 (N_19974,N_17071,N_17700);
nor U19975 (N_19975,N_17330,N_16256);
or U19976 (N_19976,N_17481,N_16983);
xor U19977 (N_19977,N_17887,N_17921);
or U19978 (N_19978,N_17333,N_17275);
nand U19979 (N_19979,N_17111,N_17185);
or U19980 (N_19980,N_17923,N_16910);
nand U19981 (N_19981,N_16098,N_17090);
and U19982 (N_19982,N_16405,N_16375);
nor U19983 (N_19983,N_17388,N_16801);
xor U19984 (N_19984,N_17916,N_16565);
nor U19985 (N_19985,N_16989,N_17353);
and U19986 (N_19986,N_16549,N_16128);
xor U19987 (N_19987,N_16569,N_16658);
and U19988 (N_19988,N_17004,N_17239);
and U19989 (N_19989,N_17748,N_17926);
or U19990 (N_19990,N_16083,N_17807);
and U19991 (N_19991,N_16117,N_17483);
nor U19992 (N_19992,N_16452,N_16370);
and U19993 (N_19993,N_16398,N_16007);
nand U19994 (N_19994,N_16865,N_16106);
xor U19995 (N_19995,N_16898,N_17016);
nor U19996 (N_19996,N_17514,N_17582);
nand U19997 (N_19997,N_16900,N_16028);
xnor U19998 (N_19998,N_16039,N_16873);
nand U19999 (N_19999,N_16190,N_16730);
xnor U20000 (N_20000,N_19728,N_18297);
or U20001 (N_20001,N_19180,N_18737);
nor U20002 (N_20002,N_18025,N_19595);
xor U20003 (N_20003,N_18186,N_18829);
nor U20004 (N_20004,N_19489,N_19476);
nor U20005 (N_20005,N_18927,N_18484);
or U20006 (N_20006,N_18434,N_18385);
nand U20007 (N_20007,N_18997,N_18991);
nor U20008 (N_20008,N_19474,N_19130);
and U20009 (N_20009,N_18042,N_19245);
or U20010 (N_20010,N_18220,N_18052);
xnor U20011 (N_20011,N_18516,N_19919);
nor U20012 (N_20012,N_18761,N_18617);
and U20013 (N_20013,N_19676,N_19109);
nor U20014 (N_20014,N_18800,N_18314);
or U20015 (N_20015,N_18588,N_19215);
xnor U20016 (N_20016,N_19636,N_18090);
or U20017 (N_20017,N_18245,N_19920);
nor U20018 (N_20018,N_18543,N_18106);
or U20019 (N_20019,N_18794,N_18177);
nor U20020 (N_20020,N_18027,N_18232);
or U20021 (N_20021,N_18460,N_18615);
or U20022 (N_20022,N_18426,N_18011);
nand U20023 (N_20023,N_19306,N_18571);
and U20024 (N_20024,N_19999,N_18867);
and U20025 (N_20025,N_18518,N_18185);
nand U20026 (N_20026,N_18868,N_18407);
xnor U20027 (N_20027,N_18221,N_18978);
nand U20028 (N_20028,N_19827,N_18870);
nand U20029 (N_20029,N_18631,N_18344);
or U20030 (N_20030,N_18359,N_18203);
xnor U20031 (N_20031,N_18134,N_18113);
xnor U20032 (N_20032,N_18575,N_19663);
and U20033 (N_20033,N_19094,N_19318);
nor U20034 (N_20034,N_19485,N_19962);
nor U20035 (N_20035,N_18764,N_19235);
xnor U20036 (N_20036,N_19185,N_19913);
nand U20037 (N_20037,N_18713,N_18288);
nand U20038 (N_20038,N_19203,N_19621);
and U20039 (N_20039,N_19517,N_19570);
and U20040 (N_20040,N_19272,N_18662);
or U20041 (N_20041,N_18551,N_18914);
or U20042 (N_20042,N_19986,N_18009);
nor U20043 (N_20043,N_19241,N_19335);
or U20044 (N_20044,N_18023,N_18087);
xnor U20045 (N_20045,N_19284,N_18539);
xor U20046 (N_20046,N_19882,N_18380);
xnor U20047 (N_20047,N_19340,N_18055);
and U20048 (N_20048,N_18020,N_18751);
nor U20049 (N_20049,N_19044,N_19724);
nand U20050 (N_20050,N_19769,N_19101);
nor U20051 (N_20051,N_18554,N_19220);
nor U20052 (N_20052,N_18367,N_19043);
or U20053 (N_20053,N_18133,N_19504);
nand U20054 (N_20054,N_18273,N_19680);
and U20055 (N_20055,N_19146,N_19748);
nor U20056 (N_20056,N_19062,N_18392);
nand U20057 (N_20057,N_19839,N_18897);
xnor U20058 (N_20058,N_19816,N_19231);
or U20059 (N_20059,N_19890,N_19701);
or U20060 (N_20060,N_18387,N_18029);
and U20061 (N_20061,N_18792,N_18907);
or U20062 (N_20062,N_18092,N_19973);
nor U20063 (N_20063,N_18108,N_19509);
nand U20064 (N_20064,N_19179,N_19520);
xnor U20065 (N_20065,N_18796,N_19332);
nand U20066 (N_20066,N_19689,N_19707);
or U20067 (N_20067,N_18293,N_18146);
or U20068 (N_20068,N_18188,N_18101);
or U20069 (N_20069,N_18022,N_18114);
or U20070 (N_20070,N_19206,N_19449);
or U20071 (N_20071,N_18136,N_18584);
nand U20072 (N_20072,N_18175,N_19696);
xor U20073 (N_20073,N_19899,N_18199);
nand U20074 (N_20074,N_19568,N_19149);
xnor U20075 (N_20075,N_19237,N_18975);
nand U20076 (N_20076,N_19246,N_18995);
nand U20077 (N_20077,N_18316,N_19699);
and U20078 (N_20078,N_19177,N_18266);
nand U20079 (N_20079,N_19114,N_18472);
and U20080 (N_20080,N_19585,N_18937);
nand U20081 (N_20081,N_18305,N_18406);
or U20082 (N_20082,N_19744,N_19995);
and U20083 (N_20083,N_19435,N_18876);
xor U20084 (N_20084,N_19194,N_18632);
and U20085 (N_20085,N_18856,N_19645);
or U20086 (N_20086,N_18140,N_18323);
nor U20087 (N_20087,N_19354,N_19025);
nor U20088 (N_20088,N_19071,N_19672);
nor U20089 (N_20089,N_19775,N_19771);
xnor U20090 (N_20090,N_18531,N_19971);
xnor U20091 (N_20091,N_19869,N_19331);
and U20092 (N_20092,N_18828,N_18289);
or U20093 (N_20093,N_19420,N_18373);
nand U20094 (N_20094,N_18393,N_19317);
or U20095 (N_20095,N_19813,N_19048);
or U20096 (N_20096,N_18283,N_18083);
and U20097 (N_20097,N_18299,N_19873);
nor U20098 (N_20098,N_19821,N_19761);
xnor U20099 (N_20099,N_19438,N_18920);
nand U20100 (N_20100,N_19455,N_18497);
and U20101 (N_20101,N_18007,N_18161);
or U20102 (N_20102,N_18388,N_19406);
nor U20103 (N_20103,N_18972,N_18681);
nor U20104 (N_20104,N_19577,N_18804);
xnor U20105 (N_20105,N_19028,N_18946);
and U20106 (N_20106,N_19785,N_18854);
and U20107 (N_20107,N_18335,N_19082);
nor U20108 (N_20108,N_19720,N_18770);
or U20109 (N_20109,N_18589,N_19429);
nor U20110 (N_20110,N_19947,N_19603);
nor U20111 (N_20111,N_19107,N_18461);
nor U20112 (N_20112,N_18673,N_18629);
xnor U20113 (N_20113,N_18481,N_19563);
nor U20114 (N_20114,N_19310,N_19549);
and U20115 (N_20115,N_18502,N_18157);
nand U20116 (N_20116,N_18984,N_19682);
nand U20117 (N_20117,N_18669,N_18532);
nand U20118 (N_20118,N_18791,N_19548);
and U20119 (N_20119,N_19214,N_18605);
or U20120 (N_20120,N_19358,N_18372);
and U20121 (N_20121,N_18331,N_19615);
or U20122 (N_20122,N_18965,N_19322);
or U20123 (N_20123,N_19841,N_19047);
or U20124 (N_20124,N_19295,N_19299);
nor U20125 (N_20125,N_18565,N_18158);
nand U20126 (N_20126,N_19679,N_19122);
nor U20127 (N_20127,N_18433,N_18892);
and U20128 (N_20128,N_19832,N_19385);
and U20129 (N_20129,N_18364,N_18477);
or U20130 (N_20130,N_19970,N_18059);
nand U20131 (N_20131,N_19933,N_19483);
and U20132 (N_20132,N_19730,N_19014);
nor U20133 (N_20133,N_18592,N_18495);
or U20134 (N_20134,N_19977,N_18882);
or U20135 (N_20135,N_18611,N_18742);
nor U20136 (N_20136,N_18895,N_18684);
xor U20137 (N_20137,N_19436,N_19802);
nand U20138 (N_20138,N_19768,N_19812);
nand U20139 (N_20139,N_18480,N_18228);
and U20140 (N_20140,N_19997,N_18853);
and U20141 (N_20141,N_19804,N_19844);
or U20142 (N_20142,N_18733,N_18339);
xnor U20143 (N_20143,N_18979,N_18390);
xor U20144 (N_20144,N_18046,N_19725);
nand U20145 (N_20145,N_19232,N_19068);
and U20146 (N_20146,N_19702,N_18465);
nand U20147 (N_20147,N_18845,N_18745);
or U20148 (N_20148,N_18744,N_18138);
nor U20149 (N_20149,N_18094,N_19265);
and U20150 (N_20150,N_19099,N_19319);
or U20151 (N_20151,N_19152,N_19355);
nand U20152 (N_20152,N_19700,N_19447);
or U20153 (N_20153,N_18568,N_18977);
and U20154 (N_20154,N_19077,N_19510);
xnor U20155 (N_20155,N_18425,N_19535);
nand U20156 (N_20156,N_19746,N_18780);
or U20157 (N_20157,N_18578,N_18529);
xnor U20158 (N_20158,N_18179,N_19249);
nor U20159 (N_20159,N_19404,N_18685);
xnor U20160 (N_20160,N_18125,N_18097);
xor U20161 (N_20161,N_19296,N_19498);
and U20162 (N_20162,N_19715,N_19770);
or U20163 (N_20163,N_19871,N_19528);
and U20164 (N_20164,N_19927,N_19872);
or U20165 (N_20165,N_18128,N_18811);
nor U20166 (N_20166,N_19974,N_18576);
or U20167 (N_20167,N_19393,N_19116);
or U20168 (N_20168,N_18889,N_19740);
and U20169 (N_20169,N_19137,N_18126);
xnor U20170 (N_20170,N_18274,N_19088);
and U20171 (N_20171,N_18064,N_19667);
nand U20172 (N_20172,N_19719,N_18071);
or U20173 (N_20173,N_18085,N_18814);
nor U20174 (N_20174,N_19642,N_18049);
or U20175 (N_20175,N_18490,N_18521);
nand U20176 (N_20176,N_18298,N_19522);
xor U20177 (N_20177,N_19566,N_19451);
nand U20178 (N_20178,N_18296,N_18812);
nand U20179 (N_20179,N_19278,N_19030);
nor U20180 (N_20180,N_19210,N_18378);
or U20181 (N_20181,N_18012,N_19035);
nor U20182 (N_20182,N_18766,N_18194);
xor U20183 (N_20183,N_19285,N_18139);
nand U20184 (N_20184,N_18900,N_19131);
xor U20185 (N_20185,N_18084,N_18201);
nand U20186 (N_20186,N_19234,N_19091);
xor U20187 (N_20187,N_18640,N_19533);
nand U20188 (N_20188,N_18835,N_18675);
nand U20189 (N_20189,N_19349,N_19789);
xor U20190 (N_20190,N_18725,N_18100);
nand U20191 (N_20191,N_19665,N_18476);
or U20192 (N_20192,N_18485,N_19594);
nand U20193 (N_20193,N_18523,N_18346);
nor U20194 (N_20194,N_19760,N_18703);
nand U20195 (N_20195,N_19968,N_19714);
and U20196 (N_20196,N_18902,N_18256);
xnor U20197 (N_20197,N_19302,N_19641);
and U20198 (N_20198,N_18430,N_18915);
xnor U20199 (N_20199,N_18533,N_19193);
or U20200 (N_20200,N_18005,N_18421);
nand U20201 (N_20201,N_18614,N_18779);
xnor U20202 (N_20202,N_19468,N_18604);
and U20203 (N_20203,N_19159,N_19567);
xor U20204 (N_20204,N_19726,N_19932);
xor U20205 (N_20205,N_19450,N_18229);
nand U20206 (N_20206,N_19481,N_18176);
or U20207 (N_20207,N_18479,N_19684);
xor U20208 (N_20208,N_18707,N_18351);
xor U20209 (N_20209,N_19323,N_18843);
nand U20210 (N_20210,N_18034,N_19041);
nor U20211 (N_20211,N_18165,N_18511);
or U20212 (N_20212,N_19938,N_18410);
nor U20213 (N_20213,N_19395,N_19316);
nor U20214 (N_20214,N_19855,N_19884);
and U20215 (N_20215,N_19542,N_18386);
or U20216 (N_20216,N_18369,N_19327);
xor U20217 (N_20217,N_19713,N_18226);
or U20218 (N_20218,N_18941,N_19524);
xnor U20219 (N_20219,N_18866,N_18603);
and U20220 (N_20220,N_18449,N_19902);
nor U20221 (N_20221,N_19826,N_18307);
and U20222 (N_20222,N_19321,N_19515);
nand U20223 (N_20223,N_19457,N_19396);
nand U20224 (N_20224,N_19743,N_18253);
nor U20225 (N_20225,N_19134,N_19367);
xor U20226 (N_20226,N_18998,N_19791);
and U20227 (N_20227,N_18024,N_19795);
nand U20228 (N_20228,N_18272,N_18704);
nor U20229 (N_20229,N_18916,N_18248);
nand U20230 (N_20230,N_18549,N_18374);
nand U20231 (N_20231,N_19007,N_18315);
xor U20232 (N_20232,N_19571,N_19192);
and U20233 (N_20233,N_19550,N_18819);
and U20234 (N_20234,N_18607,N_19410);
and U20235 (N_20235,N_18008,N_18858);
and U20236 (N_20236,N_19000,N_19664);
xnor U20237 (N_20237,N_18732,N_19247);
xnor U20238 (N_20238,N_19562,N_19338);
nand U20239 (N_20239,N_18899,N_19678);
nand U20240 (N_20240,N_18648,N_19733);
or U20241 (N_20241,N_18208,N_18738);
and U20242 (N_20242,N_19914,N_18688);
nand U20243 (N_20243,N_18381,N_18021);
nor U20244 (N_20244,N_18871,N_19484);
nor U20245 (N_20245,N_18017,N_19212);
or U20246 (N_20246,N_18382,N_19135);
nor U20247 (N_20247,N_19892,N_19300);
or U20248 (N_20248,N_19023,N_19688);
or U20249 (N_20249,N_18718,N_18668);
and U20250 (N_20250,N_18394,N_19492);
or U20251 (N_20251,N_18635,N_18187);
xnor U20252 (N_20252,N_19671,N_19691);
xor U20253 (N_20253,N_18261,N_18301);
or U20254 (N_20254,N_18620,N_18658);
and U20255 (N_20255,N_18141,N_18123);
or U20256 (N_20256,N_18864,N_18099);
and U20257 (N_20257,N_18467,N_19925);
nor U20258 (N_20258,N_19661,N_18817);
nand U20259 (N_20259,N_18417,N_18775);
or U20260 (N_20260,N_19390,N_18384);
nand U20261 (N_20261,N_19654,N_18061);
nor U20262 (N_20262,N_19467,N_18445);
or U20263 (N_20263,N_19473,N_19462);
or U20264 (N_20264,N_19494,N_18994);
xor U20265 (N_20265,N_19307,N_18127);
nor U20266 (N_20266,N_19197,N_18353);
nand U20267 (N_20267,N_18147,N_19461);
or U20268 (N_20268,N_18670,N_19526);
nand U20269 (N_20269,N_18728,N_18822);
nor U20270 (N_20270,N_19786,N_19312);
nand U20271 (N_20271,N_19787,N_19058);
or U20272 (N_20272,N_19590,N_19619);
xnor U20273 (N_20273,N_18646,N_18767);
nand U20274 (N_20274,N_19191,N_19546);
nand U20275 (N_20275,N_18526,N_19909);
or U20276 (N_20276,N_19084,N_19095);
and U20277 (N_20277,N_19065,N_18428);
nand U20278 (N_20278,N_19453,N_19334);
or U20279 (N_20279,N_18933,N_18330);
nand U20280 (N_20280,N_19710,N_18599);
xor U20281 (N_20281,N_19281,N_19779);
nor U20282 (N_20282,N_19380,N_19511);
or U20283 (N_20283,N_19994,N_18500);
nor U20284 (N_20284,N_18921,N_18789);
nor U20285 (N_20285,N_18028,N_19944);
nor U20286 (N_20286,N_19273,N_19426);
or U20287 (N_20287,N_18470,N_19421);
and U20288 (N_20288,N_18429,N_19118);
nor U20289 (N_20289,N_19709,N_19293);
nor U20290 (N_20290,N_19370,N_18156);
nor U20291 (N_20291,N_19239,N_19754);
or U20292 (N_20292,N_18820,N_18420);
nor U20293 (N_20293,N_19110,N_18016);
nor U20294 (N_20294,N_18039,N_19930);
nor U20295 (N_20295,N_19750,N_18370);
xnor U20296 (N_20296,N_19374,N_18135);
or U20297 (N_20297,N_18251,N_19963);
and U20298 (N_20298,N_19432,N_19456);
xor U20299 (N_20299,N_18486,N_18683);
xnor U20300 (N_20300,N_18045,N_19955);
or U20301 (N_20301,N_19274,N_18709);
nand U20302 (N_20302,N_19218,N_18677);
or U20303 (N_20303,N_19534,N_19958);
nand U20304 (N_20304,N_19069,N_19623);
and U20305 (N_20305,N_18983,N_19264);
or U20306 (N_20306,N_18002,N_18026);
xnor U20307 (N_20307,N_19514,N_19657);
and U20308 (N_20308,N_19252,N_19036);
or U20309 (N_20309,N_19856,N_19583);
or U20310 (N_20310,N_19998,N_18929);
xnor U20311 (N_20311,N_19064,N_19011);
nor U20312 (N_20312,N_18409,N_19989);
nand U20313 (N_20313,N_19207,N_18641);
nor U20314 (N_20314,N_18888,N_18115);
or U20315 (N_20315,N_18068,N_18333);
nand U20316 (N_20316,N_18212,N_18043);
or U20317 (N_20317,N_19482,N_19845);
and U20318 (N_20318,N_19172,N_19610);
nand U20319 (N_20319,N_18173,N_19379);
xnor U20320 (N_20320,N_18031,N_18196);
or U20321 (N_20321,N_19874,N_19433);
nand U20322 (N_20322,N_18065,N_18343);
nor U20323 (N_20323,N_19694,N_18956);
nand U20324 (N_20324,N_18698,N_19126);
or U20325 (N_20325,N_19747,N_18841);
nand U20326 (N_20326,N_18689,N_19488);
and U20327 (N_20327,N_19862,N_19924);
xnor U20328 (N_20328,N_19681,N_18679);
or U20329 (N_20329,N_18583,N_18836);
xor U20330 (N_20330,N_19120,N_18926);
xnor U20331 (N_20331,N_18540,N_18124);
or U20332 (N_20332,N_18649,N_18184);
nor U20333 (N_20333,N_18758,N_19555);
or U20334 (N_20334,N_19228,N_19383);
or U20335 (N_20335,N_18561,N_19038);
nor U20336 (N_20336,N_19002,N_18752);
nor U20337 (N_20337,N_19860,N_19151);
xnor U20338 (N_20338,N_18553,N_18708);
and U20339 (N_20339,N_18569,N_19034);
nand U20340 (N_20340,N_18881,N_18118);
nand U20341 (N_20341,N_19136,N_19407);
xnor U20342 (N_20342,N_19263,N_18719);
nand U20343 (N_20343,N_18475,N_18653);
nand U20344 (N_20344,N_19348,N_18545);
and U20345 (N_20345,N_19829,N_18803);
nor U20346 (N_20346,N_18070,N_18863);
or U20347 (N_20347,N_19105,N_18909);
and U20348 (N_20348,N_18210,N_18967);
nand U20349 (N_20349,N_19428,N_18924);
nor U20350 (N_20350,N_19119,N_19660);
nand U20351 (N_20351,N_18038,N_19092);
nor U20352 (N_20352,N_19073,N_19497);
and U20353 (N_20353,N_18181,N_19063);
or U20354 (N_20354,N_18341,N_18847);
and U20355 (N_20355,N_18504,N_18325);
nor U20356 (N_20356,N_19113,N_19153);
or U20357 (N_20357,N_18944,N_18722);
nand U20358 (N_20358,N_18556,N_18195);
xor U20359 (N_20359,N_18150,N_18285);
nor U20360 (N_20360,N_19183,N_19588);
nor U20361 (N_20361,N_18759,N_19521);
nand U20362 (N_20362,N_18348,N_19934);
nand U20363 (N_20363,N_18260,N_19276);
or U20364 (N_20364,N_19767,N_18117);
nor U20365 (N_20365,N_19818,N_19311);
xor U20366 (N_20366,N_19411,N_19764);
or U20367 (N_20367,N_19799,N_19557);
nor U20368 (N_20368,N_19801,N_18427);
xnor U20369 (N_20369,N_18659,N_19778);
or U20370 (N_20370,N_18633,N_18252);
nor U20371 (N_20371,N_18939,N_18522);
or U20372 (N_20372,N_18934,N_19441);
nand U20373 (N_20373,N_19591,N_18730);
nor U20374 (N_20374,N_18075,N_18352);
xor U20375 (N_20375,N_18174,N_18626);
nand U20376 (N_20376,N_18950,N_19267);
xnor U20377 (N_20377,N_19811,N_18699);
or U20378 (N_20378,N_19868,N_19144);
nor U20379 (N_20379,N_18906,N_18238);
xor U20380 (N_20380,N_18415,N_18838);
nor U20381 (N_20381,N_19403,N_18957);
or U20382 (N_20382,N_19951,N_19916);
nand U20383 (N_20383,N_19190,N_18462);
and U20384 (N_20384,N_19042,N_19551);
and U20385 (N_20385,N_18163,N_18999);
nor U20386 (N_20386,N_18701,N_19798);
nor U20387 (N_20387,N_18802,N_19257);
and U20388 (N_20388,N_18981,N_19851);
and U20389 (N_20389,N_19056,N_18337);
nor U20390 (N_20390,N_19347,N_19527);
xnor U20391 (N_20391,N_18785,N_19260);
and U20392 (N_20392,N_18474,N_19169);
and U20393 (N_20393,N_18078,N_18250);
nor U20394 (N_20394,N_18391,N_19202);
nor U20395 (N_20395,N_19271,N_19901);
nand U20396 (N_20396,N_18874,N_19132);
nor U20397 (N_20397,N_19060,N_19647);
nor U20398 (N_20398,N_19478,N_18538);
xor U20399 (N_20399,N_18182,N_18807);
and U20400 (N_20400,N_18851,N_19400);
and U20401 (N_20401,N_18143,N_19518);
nand U20402 (N_20402,N_18437,N_18326);
or U20403 (N_20403,N_19722,N_18682);
nand U20404 (N_20404,N_18625,N_18102);
nor U20405 (N_20405,N_18306,N_19121);
nor U20406 (N_20406,N_19343,N_19634);
and U20407 (N_20407,N_18862,N_19125);
nor U20408 (N_20408,N_18993,N_18643);
nor U20409 (N_20409,N_18989,N_18609);
and U20410 (N_20410,N_19824,N_19112);
and U20411 (N_20411,N_18690,N_19953);
nor U20412 (N_20412,N_19303,N_18441);
and U20413 (N_20413,N_18573,N_18636);
or U20414 (N_20414,N_18754,N_19875);
and U20415 (N_20415,N_19990,N_18593);
nor U20416 (N_20416,N_18786,N_19275);
nor U20417 (N_20417,N_18855,N_19376);
nand U20418 (N_20418,N_19941,N_18623);
or U20419 (N_20419,N_18268,N_19157);
xor U20420 (N_20420,N_18379,N_18755);
nand U20421 (N_20421,N_18990,N_19597);
and U20422 (N_20422,N_19578,N_19602);
xor U20423 (N_20423,N_19359,N_18627);
or U20424 (N_20424,N_18000,N_19848);
nor U20425 (N_20425,N_19800,N_19793);
and U20426 (N_20426,N_19238,N_18799);
nand U20427 (N_20427,N_19176,N_18107);
xor U20428 (N_20428,N_18763,N_19943);
nand U20429 (N_20429,N_19859,N_18507);
xnor U20430 (N_20430,N_18471,N_18564);
nand U20431 (N_20431,N_18726,N_19499);
xor U20432 (N_20432,N_19732,N_19516);
nor U20433 (N_20433,N_19115,N_19020);
nand U20434 (N_20434,N_19434,N_18715);
xnor U20435 (N_20435,N_18204,N_18563);
nand U20436 (N_20436,N_18439,N_18801);
or U20437 (N_20437,N_18618,N_19731);
or U20438 (N_20438,N_19059,N_18765);
xor U20439 (N_20439,N_18422,N_19049);
nand U20440 (N_20440,N_18198,N_19967);
xnor U20441 (N_20441,N_18654,N_18089);
nand U20442 (N_20442,N_19031,N_19586);
nor U20443 (N_20443,N_18456,N_19547);
xor U20444 (N_20444,N_18879,N_18413);
and U20445 (N_20445,N_19894,N_19513);
xnor U20446 (N_20446,N_19928,N_18714);
or U20447 (N_20447,N_18448,N_18041);
xor U20448 (N_20448,N_18361,N_18001);
nand U20449 (N_20449,N_19500,N_19051);
nor U20450 (N_20450,N_19329,N_19108);
or U20451 (N_20451,N_18963,N_19965);
or U20452 (N_20452,N_19074,N_19344);
xnor U20453 (N_20453,N_19838,N_18395);
nor U20454 (N_20454,N_19454,N_19541);
or U20455 (N_20455,N_19337,N_19032);
nand U20456 (N_20456,N_18674,N_19600);
nor U20457 (N_20457,N_19250,N_18606);
nand U20458 (N_20458,N_19258,N_19530);
nor U20459 (N_20459,N_19553,N_18727);
xnor U20460 (N_20460,N_18865,N_18162);
xnor U20461 (N_20461,N_19906,N_19632);
and U20462 (N_20462,N_19244,N_18520);
xor U20463 (N_20463,N_18458,N_19606);
xor U20464 (N_20464,N_18541,N_18711);
nor U20465 (N_20465,N_19262,N_18197);
and U20466 (N_20466,N_18544,N_19360);
nor U20467 (N_20467,N_18572,N_18294);
xor U20468 (N_20468,N_18825,N_18696);
or U20469 (N_20469,N_19897,N_19341);
or U20470 (N_20470,N_19749,N_19001);
or U20471 (N_20471,N_19050,N_19774);
and U20472 (N_20472,N_18214,N_18033);
xor U20473 (N_20473,N_19537,N_19415);
xnor U20474 (N_20474,N_19822,N_19877);
nand U20475 (N_20475,N_18355,N_18885);
or U20476 (N_20476,N_18769,N_18922);
or U20477 (N_20477,N_18290,N_19090);
nand U20478 (N_20478,N_19219,N_19718);
nor U20479 (N_20479,N_18190,N_19282);
or U20480 (N_20480,N_19605,N_18336);
or U20481 (N_20481,N_18040,N_19904);
xnor U20482 (N_20482,N_18300,N_18079);
nor U20483 (N_20483,N_19269,N_18067);
nor U20484 (N_20484,N_19846,N_19430);
nand U20485 (N_20485,N_19425,N_19666);
nand U20486 (N_20486,N_18400,N_18567);
and U20487 (N_20487,N_18846,N_19926);
nand U20488 (N_20488,N_19805,N_19614);
nand U20489 (N_20489,N_18356,N_19782);
or U20490 (N_20490,N_19458,N_19387);
or U20491 (N_20491,N_19066,N_19626);
nor U20492 (N_20492,N_18697,N_18557);
nor U20493 (N_20493,N_18438,N_19369);
or U20494 (N_20494,N_18757,N_19708);
nor U20495 (N_20495,N_18741,N_19022);
nor U20496 (N_20496,N_18656,N_19532);
nand U20497 (N_20497,N_18239,N_19723);
and U20498 (N_20498,N_19189,N_19501);
nand U20499 (N_20499,N_18524,N_19604);
or U20500 (N_20500,N_19196,N_19921);
nor U20501 (N_20501,N_19652,N_18911);
xor U20502 (N_20502,N_19756,N_18269);
nand U20503 (N_20503,N_18154,N_18246);
and U20504 (N_20504,N_19229,N_19394);
and U20505 (N_20505,N_18235,N_18223);
and U20506 (N_20506,N_18231,N_19290);
and U20507 (N_20507,N_18932,N_18886);
xor U20508 (N_20508,N_19147,N_19599);
or U20509 (N_20509,N_18267,N_19683);
and U20510 (N_20510,N_19784,N_18377);
nand U20511 (N_20511,N_18837,N_19009);
or U20512 (N_20512,N_19111,N_18263);
and U20513 (N_20513,N_19883,N_18287);
and U20514 (N_20514,N_19399,N_19163);
xor U20515 (N_20515,N_18959,N_19737);
and U20516 (N_20516,N_18418,N_18974);
xnor U20517 (N_20517,N_19620,N_19964);
or U20518 (N_20518,N_19674,N_18284);
nand U20519 (N_20519,N_19187,N_19423);
nand U20520 (N_20520,N_19093,N_18376);
and U20521 (N_20521,N_19992,N_19685);
xnor U20522 (N_20522,N_19029,N_19849);
or U20523 (N_20523,N_19825,N_18350);
or U20524 (N_20524,N_19475,N_19646);
nor U20525 (N_20525,N_19611,N_19757);
and U20526 (N_20526,N_18058,N_19503);
nand U20527 (N_20527,N_18202,N_19167);
and U20528 (N_20528,N_18686,N_18663);
nor U20529 (N_20529,N_18310,N_19216);
xor U20530 (N_20530,N_18896,N_19649);
xor U20531 (N_20531,N_18574,N_19978);
xnor U20532 (N_20532,N_18652,N_18015);
nor U20533 (N_20533,N_18612,N_19070);
xnor U20534 (N_20534,N_19294,N_18651);
and U20535 (N_20535,N_19096,N_19922);
and U20536 (N_20536,N_19917,N_18710);
nand U20537 (N_20537,N_18706,N_19418);
or U20538 (N_20538,N_19138,N_19937);
nand U20539 (N_20539,N_19479,N_19975);
nand U20540 (N_20540,N_18601,N_19170);
and U20541 (N_20541,N_18322,N_19704);
nor U20542 (N_20542,N_19046,N_19133);
nor U20543 (N_20543,N_19956,N_19419);
or U20544 (N_20544,N_18051,N_18227);
or U20545 (N_20545,N_18816,N_19079);
and U20546 (N_20546,N_18517,N_19286);
nand U20547 (N_20547,N_19377,N_18166);
nor U20548 (N_20548,N_19309,N_19414);
xor U20549 (N_20549,N_19445,N_19512);
and U20550 (N_20550,N_18443,N_18328);
or U20551 (N_20551,N_19324,N_18209);
xnor U20552 (N_20552,N_18905,N_18105);
xor U20553 (N_20553,N_18295,N_18230);
xor U20554 (N_20554,N_18717,N_19424);
nor U20555 (N_20555,N_18469,N_18840);
nand U20556 (N_20556,N_19543,N_18729);
or U20557 (N_20557,N_19427,N_18151);
xnor U20558 (N_20558,N_19466,N_18170);
nand U20559 (N_20559,N_18037,N_18875);
or U20560 (N_20560,N_18233,N_19560);
nand U20561 (N_20561,N_18596,N_19356);
and U20562 (N_20562,N_18657,N_19658);
nor U20563 (N_20563,N_18363,N_18528);
nand U20564 (N_20564,N_18189,N_18970);
nand U20565 (N_20565,N_19662,N_19174);
xnor U20566 (N_20566,N_19182,N_18806);
and U20567 (N_20567,N_18705,N_18961);
nor U20568 (N_20568,N_18442,N_19315);
nor U20569 (N_20569,N_19631,N_19195);
nor U20570 (N_20570,N_18960,N_19227);
xnor U20571 (N_20571,N_19879,N_18436);
and U20572 (N_20572,N_18692,N_19040);
or U20573 (N_20573,N_18622,N_18947);
or U20574 (N_20574,N_18508,N_18120);
nor U20575 (N_20575,N_18243,N_19507);
or U20576 (N_20576,N_19398,N_18942);
and U20577 (N_20577,N_18219,N_19005);
and U20578 (N_20578,N_19397,N_19729);
nand U20579 (N_20579,N_19470,N_19142);
or U20580 (N_20580,N_18968,N_19444);
and U20581 (N_20581,N_18548,N_19876);
nor U20582 (N_20582,N_19006,N_19721);
and U20583 (N_20583,N_19165,N_19352);
xnor U20584 (N_20584,N_19717,N_19854);
and U20585 (N_20585,N_18810,N_18530);
nor U20586 (N_20586,N_19361,N_19261);
nand U20587 (N_20587,N_18602,N_19129);
nand U20588 (N_20588,N_18945,N_19186);
nand U20589 (N_20589,N_19008,N_18503);
nand U20590 (N_20590,N_19253,N_19128);
nand U20591 (N_20591,N_18349,N_19103);
and U20592 (N_20592,N_18488,N_19828);
and U20593 (N_20593,N_18416,N_18778);
nand U20594 (N_20594,N_18506,N_19493);
or U20595 (N_20595,N_18671,N_19582);
nand U20596 (N_20596,N_18137,N_19712);
and U20597 (N_20597,N_19243,N_19745);
or U20598 (N_20598,N_19648,N_18224);
and U20599 (N_20599,N_19984,N_19305);
xor U20600 (N_20600,N_18076,N_18869);
nand U20601 (N_20601,N_18457,N_18424);
and U20602 (N_20602,N_18590,N_19201);
and U20603 (N_20603,N_18047,N_18702);
or U20604 (N_20604,N_18489,N_19918);
nor U20605 (N_20605,N_18958,N_19505);
xor U20606 (N_20606,N_18397,N_18795);
or U20607 (N_20607,N_19233,N_18639);
xnor U20608 (N_20608,N_19353,N_18036);
nor U20609 (N_20609,N_19181,N_18756);
and U20610 (N_20610,N_19842,N_19659);
nand U20611 (N_20611,N_18303,N_18672);
nor U20612 (N_20612,N_19788,N_18772);
nand U20613 (N_20613,N_19477,N_18057);
xnor U20614 (N_20614,N_18493,N_19819);
xor U20615 (N_20615,N_19288,N_19373);
nand U20616 (N_20616,N_19575,N_18452);
nand U20617 (N_20617,N_18976,N_18514);
or U20618 (N_20618,N_19959,N_18857);
or U20619 (N_20619,N_19929,N_19004);
or U20620 (N_20620,N_19437,N_18292);
xor U20621 (N_20621,N_19810,N_19205);
or U20622 (N_20622,N_18271,N_18628);
or U20623 (N_20623,N_19858,N_18890);
nand U20624 (N_20624,N_18798,N_19536);
nor U20625 (N_20625,N_18095,N_18172);
xnor U20626 (N_20626,N_18582,N_18581);
xnor U20627 (N_20627,N_18784,N_18168);
and U20628 (N_20628,N_18423,N_19375);
nand U20629 (N_20629,N_18142,N_18444);
nand U20630 (N_20630,N_19495,N_18093);
nand U20631 (N_20631,N_19703,N_19053);
or U20632 (N_20632,N_19753,N_19766);
and U20633 (N_20633,N_19490,N_18213);
and U20634 (N_20634,N_19166,N_18585);
nor U20635 (N_20635,N_19817,N_19148);
and U20636 (N_20636,N_18739,N_18122);
nand U20637 (N_20637,N_18537,N_18734);
nor U20638 (N_20638,N_18859,N_19382);
nor U20639 (N_20639,N_18808,N_19581);
and U20640 (N_20640,N_18365,N_18073);
nand U20641 (N_20641,N_18414,N_19037);
nand U20642 (N_20642,N_18345,N_19808);
nor U20643 (N_20643,N_18969,N_19448);
xnor U20644 (N_20644,N_19836,N_19886);
and U20645 (N_20645,N_19900,N_19706);
nand U20646 (N_20646,N_19629,N_19378);
xor U20647 (N_20647,N_18144,N_18237);
nor U20648 (N_20648,N_19178,N_19673);
xnor U20649 (N_20649,N_18404,N_19351);
and U20650 (N_20650,N_18178,N_19628);
or U20651 (N_20651,N_18498,N_18192);
nor U20652 (N_20652,N_19173,N_19698);
nand U20653 (N_20653,N_19052,N_18389);
nand U20654 (N_20654,N_19559,N_18566);
xnor U20655 (N_20655,N_18119,N_18048);
or U20656 (N_20656,N_19465,N_18340);
nand U20657 (N_20657,N_18700,N_18996);
or U20658 (N_20658,N_19638,N_19291);
and U20659 (N_20659,N_18987,N_19806);
nand U20660 (N_20660,N_18304,N_19055);
xnor U20661 (N_20661,N_19230,N_19017);
nand U20662 (N_20662,N_19388,N_19452);
nor U20663 (N_20663,N_19102,N_18383);
nor U20664 (N_20664,N_18749,N_18281);
nand U20665 (N_20665,N_18399,N_19942);
and U20666 (N_20666,N_19814,N_18275);
or U20667 (N_20667,N_19283,N_19607);
or U20668 (N_20668,N_19168,N_18234);
nor U20669 (N_20669,N_18823,N_19019);
and U20670 (N_20670,N_19308,N_18155);
or U20671 (N_20671,N_19695,N_18160);
and U20672 (N_20672,N_19083,N_19416);
and U20673 (N_20673,N_19155,N_19950);
xor U20674 (N_20674,N_18748,N_18586);
xor U20675 (N_20675,N_18953,N_19217);
or U20676 (N_20676,N_19630,N_19736);
nand U20677 (N_20677,N_18884,N_19655);
xnor U20678 (N_20678,N_18743,N_19865);
nand U20679 (N_20679,N_19716,N_18225);
or U20680 (N_20680,N_19891,N_19863);
nor U20681 (N_20681,N_19259,N_18447);
and U20682 (N_20682,N_19143,N_19803);
and U20683 (N_20683,N_19045,N_18952);
nand U20684 (N_20684,N_18562,N_18839);
and U20685 (N_20685,N_18054,N_18809);
nor U20686 (N_20686,N_18215,N_18247);
or U20687 (N_20687,N_19896,N_19616);
or U20688 (N_20688,N_19459,N_19643);
nor U20689 (N_20689,N_19670,N_19690);
and U20690 (N_20690,N_18018,N_19739);
or U20691 (N_20691,N_18004,N_19952);
nor U20692 (N_20692,N_19076,N_19248);
xor U20693 (N_20693,N_19080,N_18903);
nand U20694 (N_20694,N_19003,N_19980);
and U20695 (N_20695,N_19371,N_18494);
xnor U20696 (N_20696,N_19907,N_18193);
or U20697 (N_20697,N_19668,N_18830);
xnor U20698 (N_20698,N_18091,N_18624);
nand U20699 (N_20699,N_18419,N_18478);
xor U20700 (N_20700,N_18110,N_18962);
nand U20701 (N_20701,N_18638,N_19589);
or U20702 (N_20702,N_19540,N_19491);
nor U20703 (N_20703,N_19408,N_19580);
nor U20704 (N_20704,N_19391,N_18510);
or U20705 (N_20705,N_19364,N_19463);
and U20706 (N_20706,N_18276,N_19640);
or U20707 (N_20707,N_18129,N_19852);
or U20708 (N_20708,N_18716,N_18600);
nor U20709 (N_20709,N_18312,N_19413);
nand U20710 (N_20710,N_19443,N_18329);
xor U20711 (N_20711,N_19081,N_18948);
and U20712 (N_20712,N_19389,N_19790);
xnor U20713 (N_20713,N_18555,N_19328);
xnor U20714 (N_20714,N_19752,N_19912);
xor U20715 (N_20715,N_18608,N_18883);
xnor U20716 (N_20716,N_18736,N_18720);
nand U20717 (N_20717,N_18619,N_18262);
and U20718 (N_20718,N_18955,N_19297);
and U20719 (N_20719,N_18216,N_19574);
xnor U20720 (N_20720,N_19837,N_18964);
nand U20721 (N_20721,N_18797,N_19277);
nand U20722 (N_20722,N_18667,N_19117);
nand U20723 (N_20723,N_18793,N_18781);
nor U20724 (N_20724,N_18398,N_18111);
or U20725 (N_20725,N_19987,N_18912);
or U20726 (N_20726,N_19573,N_18824);
nor U20727 (N_20727,N_19089,N_19758);
xor U20728 (N_20728,N_18446,N_19976);
and U20729 (N_20729,N_18255,N_19368);
nand U20730 (N_20730,N_18762,N_18525);
or U20731 (N_20731,N_18342,N_19996);
or U20732 (N_20732,N_18826,N_18318);
xnor U20733 (N_20733,N_18616,N_19339);
and U20734 (N_20734,N_18116,N_19693);
nor U20735 (N_20735,N_19268,N_18412);
and U20736 (N_20736,N_18286,N_18062);
or U20737 (N_20737,N_18773,N_18860);
xor U20738 (N_20738,N_19697,N_19075);
and U20739 (N_20739,N_18935,N_19439);
nand U20740 (N_20740,N_18130,N_19830);
nor U20741 (N_20741,N_19960,N_18153);
nand U20742 (N_20742,N_18848,N_18450);
nand U20743 (N_20743,N_19139,N_18753);
nor U20744 (N_20744,N_19392,N_19106);
or U20745 (N_20745,N_18030,N_18032);
nor U20746 (N_20746,N_19910,N_19908);
nor U20747 (N_20747,N_18973,N_18077);
or U20748 (N_20748,N_19508,N_18191);
nor U20749 (N_20749,N_18180,N_18200);
nor U20750 (N_20750,N_18695,N_18842);
or U20751 (N_20751,N_19864,N_19027);
or U20752 (N_20752,N_18731,N_19773);
and U20753 (N_20753,N_19936,N_18676);
nand U20754 (N_20754,N_18904,N_18887);
nand U20755 (N_20755,N_19985,N_19538);
nand U20756 (N_20756,N_19336,N_18171);
or U20757 (N_20757,N_18455,N_19204);
nand U20758 (N_20758,N_19572,N_19422);
xor U20759 (N_20759,N_19923,N_18003);
nor U20760 (N_20760,N_19981,N_18453);
and U20761 (N_20761,N_18347,N_19893);
or U20762 (N_20762,N_18519,N_18279);
or U20763 (N_20763,N_19991,N_19781);
and U20764 (N_20764,N_19363,N_19677);
nand U20765 (N_20765,N_18362,N_19471);
or U20766 (N_20766,N_19150,N_19417);
xnor U20767 (N_20767,N_18546,N_19067);
xor U20768 (N_20768,N_18930,N_19866);
or U20769 (N_20769,N_19292,N_18815);
xnor U20770 (N_20770,N_19366,N_18918);
or U20771 (N_20771,N_19222,N_18496);
nor U20772 (N_20772,N_18735,N_18159);
and U20773 (N_20773,N_18149,N_19372);
xor U20774 (N_20774,N_18534,N_18901);
xor U20775 (N_20775,N_18844,N_19539);
or U20776 (N_20776,N_18321,N_18332);
xnor U20777 (N_20777,N_19010,N_19525);
xnor U20778 (N_20778,N_18282,N_18435);
nor U20779 (N_20779,N_18597,N_19885);
or U20780 (N_20780,N_19644,N_18645);
xnor U20781 (N_20781,N_19792,N_19759);
and U20782 (N_20782,N_18207,N_19911);
or U20783 (N_20783,N_19350,N_19487);
xor U20784 (N_20784,N_18121,N_19561);
nor U20785 (N_20785,N_18081,N_19738);
nand U20786 (N_20786,N_19381,N_18550);
nor U20787 (N_20787,N_19870,N_19320);
nor U20788 (N_20788,N_18264,N_19776);
nor U20789 (N_20789,N_19325,N_18938);
xor U20790 (N_20790,N_19145,N_19598);
nand U20791 (N_20791,N_19840,N_18894);
nand U20792 (N_20792,N_18587,N_18813);
or U20793 (N_20793,N_18069,N_19780);
nor U20794 (N_20794,N_18291,N_18872);
and U20795 (N_20795,N_18459,N_18831);
or U20796 (N_20796,N_18145,N_18919);
nand U20797 (N_20797,N_19236,N_18463);
nor U20798 (N_20798,N_19887,N_19794);
or U20799 (N_20799,N_19496,N_18499);
and U20800 (N_20800,N_18072,N_18661);
nand U20801 (N_20801,N_19815,N_18878);
xor U20802 (N_20802,N_19531,N_19905);
and U20803 (N_20803,N_19915,N_18760);
nor U20804 (N_20804,N_19564,N_18552);
nand U20805 (N_20805,N_18746,N_18783);
nor U20806 (N_20806,N_19097,N_18971);
nor U20807 (N_20807,N_19835,N_18877);
nor U20808 (N_20808,N_19624,N_18594);
xor U20809 (N_20809,N_18320,N_18723);
xor U20810 (N_20810,N_18169,N_19617);
nor U20811 (N_20811,N_19446,N_18308);
nand U20812 (N_20812,N_18908,N_18368);
and U20813 (N_20813,N_18610,N_19656);
nand U20814 (N_20814,N_19405,N_19633);
and U20815 (N_20815,N_18923,N_19519);
or U20816 (N_20816,N_18647,N_18805);
or U20817 (N_20817,N_18265,N_18992);
xnor U20818 (N_20818,N_19669,N_19625);
xor U20819 (N_20819,N_18103,N_18244);
xor U20820 (N_20820,N_18491,N_19160);
xor U20821 (N_20821,N_19592,N_18660);
or U20822 (N_20822,N_18466,N_18066);
nand U20823 (N_20823,N_18613,N_18982);
xor U20824 (N_20824,N_19061,N_19280);
or U20825 (N_20825,N_19587,N_18112);
xnor U20826 (N_20826,N_18249,N_18013);
xnor U20827 (N_20827,N_18019,N_19796);
nand U20828 (N_20828,N_19225,N_18010);
nor U20829 (N_20829,N_18790,N_19221);
nand U20830 (N_20830,N_19878,N_19650);
nand U20831 (N_20831,N_19523,N_18724);
or U20832 (N_20832,N_18691,N_19946);
nand U20833 (N_20833,N_18634,N_18771);
xnor U20834 (N_20834,N_19188,N_18050);
xnor U20835 (N_20835,N_18371,N_19940);
xor U20836 (N_20836,N_19544,N_19705);
and U20837 (N_20837,N_19431,N_19584);
xor U20838 (N_20838,N_18468,N_18309);
nor U20839 (N_20839,N_19464,N_18403);
and U20840 (N_20840,N_19289,N_19057);
nor U20841 (N_20841,N_19881,N_18666);
and U20842 (N_20842,N_18056,N_18747);
xnor U20843 (N_20843,N_18319,N_18893);
nor U20844 (N_20844,N_18818,N_19240);
nor U20845 (N_20845,N_18650,N_19270);
nor U20846 (N_20846,N_19140,N_18082);
or U20847 (N_20847,N_18236,N_19472);
and U20848 (N_20848,N_18547,N_19460);
or U20849 (N_20849,N_19156,N_18402);
xnor U20850 (N_20850,N_18454,N_18088);
or U20851 (N_20851,N_18985,N_19569);
and U20852 (N_20852,N_19033,N_18483);
and U20853 (N_20853,N_19558,N_18501);
nor U20854 (N_20854,N_18360,N_19330);
nand U20855 (N_20855,N_19618,N_18577);
or U20856 (N_20856,N_19301,N_18850);
xor U20857 (N_20857,N_19861,N_18152);
nor U20858 (N_20858,N_18687,N_19637);
and U20859 (N_20859,N_18943,N_19969);
nand U20860 (N_20860,N_18925,N_18988);
xnor U20861 (N_20861,N_19104,N_19409);
or U20862 (N_20862,N_18642,N_18375);
nor U20863 (N_20863,N_19021,N_19087);
nand U20864 (N_20864,N_19675,N_19098);
and U20865 (N_20865,N_18313,N_18664);
or U20866 (N_20866,N_18183,N_19256);
nor U20867 (N_20867,N_19013,N_18913);
and U20868 (N_20868,N_18401,N_19741);
nand U20869 (N_20869,N_18579,N_19026);
xor U20870 (N_20870,N_18954,N_19949);
nor U20871 (N_20871,N_18655,N_18536);
nand U20872 (N_20872,N_19164,N_19820);
and U20873 (N_20873,N_18951,N_19545);
nand U20874 (N_20874,N_18311,N_19442);
nand U20875 (N_20875,N_19898,N_18560);
nand U20876 (N_20876,N_18740,N_18240);
nor U20877 (N_20877,N_18431,N_19653);
and U20878 (N_20878,N_19935,N_19762);
xnor U20879 (N_20879,N_18473,N_18411);
and U20880 (N_20880,N_18542,N_18928);
or U20881 (N_20881,N_18637,N_18317);
nor U20882 (N_20882,N_18324,N_19209);
nor U20883 (N_20883,N_19154,N_19601);
nand U20884 (N_20884,N_18949,N_19651);
and U20885 (N_20885,N_18148,N_18852);
nor U20886 (N_20886,N_18630,N_18891);
nand U20887 (N_20887,N_18750,N_19171);
or U20888 (N_20888,N_18211,N_18665);
and U20889 (N_20889,N_18777,N_18832);
or U20890 (N_20890,N_18512,N_18132);
nand U20891 (N_20891,N_19386,N_18074);
and U20892 (N_20892,N_18241,N_18060);
and U20893 (N_20893,N_18513,N_19612);
nor U20894 (N_20894,N_18861,N_18131);
and U20895 (N_20895,N_19831,N_19018);
nand U20896 (N_20896,N_18257,N_18492);
xnor U20897 (N_20897,N_19486,N_19198);
and U20898 (N_20898,N_18254,N_19184);
xnor U20899 (N_20899,N_18787,N_19401);
or U20900 (N_20900,N_19735,N_18598);
or U20901 (N_20901,N_19734,N_19357);
nor U20902 (N_20902,N_19304,N_18910);
or U20903 (N_20903,N_18405,N_18086);
and U20904 (N_20904,N_19834,N_19298);
or U20905 (N_20905,N_18206,N_18898);
nor U20906 (N_20906,N_18833,N_18006);
and U20907 (N_20907,N_19480,N_19554);
nor U20908 (N_20908,N_18821,N_18440);
and U20909 (N_20909,N_18164,N_19502);
or U20910 (N_20910,N_19012,N_19809);
nor U20911 (N_20911,N_18354,N_18644);
nor U20912 (N_20912,N_18580,N_19015);
nor U20913 (N_20913,N_18986,N_18776);
nor U20914 (N_20914,N_18505,N_19161);
or U20915 (N_20915,N_18768,N_18044);
nor U20916 (N_20916,N_19333,N_19850);
xor U20917 (N_20917,N_19345,N_19469);
and U20918 (N_20918,N_19072,N_19823);
nand U20919 (N_20919,N_18408,N_18218);
nand U20920 (N_20920,N_19251,N_19847);
and U20921 (N_20921,N_18259,N_18558);
and U20922 (N_20922,N_19843,N_19402);
nor U20923 (N_20923,N_18096,N_18931);
and U20924 (N_20924,N_19162,N_19211);
nand U20925 (N_20925,N_18270,N_19867);
nand U20926 (N_20926,N_18222,N_18327);
or U20927 (N_20927,N_19954,N_18880);
nor U20928 (N_20928,N_19895,N_18535);
xnor U20929 (N_20929,N_19889,N_19124);
and U20930 (N_20930,N_18482,N_19686);
xnor U20931 (N_20931,N_18827,N_19777);
nand U20932 (N_20932,N_19226,N_19635);
or U20933 (N_20933,N_19727,N_18432);
and U20934 (N_20934,N_18966,N_18680);
nand U20935 (N_20935,N_19313,N_19765);
xnor U20936 (N_20936,N_18774,N_19552);
nor U20937 (N_20937,N_19127,N_18035);
and U20938 (N_20938,N_19242,N_18509);
or U20939 (N_20939,N_18834,N_19158);
nor U20940 (N_20940,N_19593,N_19565);
nor U20941 (N_20941,N_19888,N_19711);
or U20942 (N_20942,N_19853,N_18366);
nor U20943 (N_20943,N_19199,N_18053);
nand U20944 (N_20944,N_19807,N_19983);
xor U20945 (N_20945,N_19751,N_18334);
and U20946 (N_20946,N_18782,N_19979);
and U20947 (N_20947,N_18338,N_19342);
and U20948 (N_20948,N_19556,N_18849);
or U20949 (N_20949,N_18712,N_19100);
nand U20950 (N_20950,N_18464,N_19287);
and U20951 (N_20951,N_19880,N_19506);
or U20952 (N_20952,N_18217,N_19200);
nand U20953 (N_20953,N_18621,N_18721);
and U20954 (N_20954,N_19326,N_19783);
and U20955 (N_20955,N_19224,N_19939);
and U20956 (N_20956,N_18940,N_19988);
nor U20957 (N_20957,N_19255,N_18980);
nand U20958 (N_20958,N_19123,N_18167);
nor U20959 (N_20959,N_19609,N_19039);
nor U20960 (N_20960,N_18278,N_19223);
nor U20961 (N_20961,N_19365,N_18451);
or U20962 (N_20962,N_18515,N_19579);
xnor U20963 (N_20963,N_19931,N_19608);
or U20964 (N_20964,N_19639,N_18357);
xor U20965 (N_20965,N_19622,N_19208);
nand U20966 (N_20966,N_19613,N_19384);
and U20967 (N_20967,N_18917,N_18205);
and U20968 (N_20968,N_19078,N_19857);
nor U20969 (N_20969,N_18063,N_19213);
or U20970 (N_20970,N_18570,N_18014);
and U20971 (N_20971,N_19362,N_19687);
or U20972 (N_20972,N_18109,N_19833);
and U20973 (N_20973,N_19529,N_19972);
or U20974 (N_20974,N_18595,N_19266);
nand U20975 (N_20975,N_19692,N_19440);
xnor U20976 (N_20976,N_19254,N_19085);
nor U20977 (N_20977,N_18358,N_19175);
nand U20978 (N_20978,N_19961,N_19346);
and U20979 (N_20979,N_19797,N_19742);
xnor U20980 (N_20980,N_18242,N_19596);
or U20981 (N_20981,N_19993,N_18302);
nor U20982 (N_20982,N_19903,N_19966);
xnor U20983 (N_20983,N_19314,N_19016);
nor U20984 (N_20984,N_19755,N_18487);
nor U20985 (N_20985,N_19279,N_19054);
nor U20986 (N_20986,N_19772,N_18693);
or U20987 (N_20987,N_18280,N_18559);
or U20988 (N_20988,N_18788,N_19024);
nand U20989 (N_20989,N_18873,N_18396);
nor U20990 (N_20990,N_18277,N_19086);
or U20991 (N_20991,N_19957,N_18080);
xnor U20992 (N_20992,N_18527,N_19948);
and U20993 (N_20993,N_18098,N_18678);
and U20994 (N_20994,N_19576,N_18591);
nor U20995 (N_20995,N_18694,N_19141);
nand U20996 (N_20996,N_19627,N_19945);
and U20997 (N_20997,N_19412,N_18258);
nand U20998 (N_20998,N_18936,N_18104);
nand U20999 (N_20999,N_19763,N_19982);
or U21000 (N_21000,N_19282,N_19515);
xnor U21001 (N_21001,N_19835,N_18272);
nand U21002 (N_21002,N_18722,N_19256);
nor U21003 (N_21003,N_19726,N_18602);
nand U21004 (N_21004,N_19419,N_18344);
and U21005 (N_21005,N_19164,N_19165);
and U21006 (N_21006,N_19236,N_18138);
nand U21007 (N_21007,N_18727,N_19846);
or U21008 (N_21008,N_18140,N_19974);
xnor U21009 (N_21009,N_19141,N_19186);
nor U21010 (N_21010,N_18165,N_19218);
nor U21011 (N_21011,N_18306,N_18471);
or U21012 (N_21012,N_18212,N_19997);
and U21013 (N_21013,N_18232,N_19606);
or U21014 (N_21014,N_19664,N_19827);
and U21015 (N_21015,N_18013,N_19280);
or U21016 (N_21016,N_18667,N_19202);
nor U21017 (N_21017,N_18348,N_19557);
nand U21018 (N_21018,N_18802,N_18120);
xor U21019 (N_21019,N_19631,N_18392);
xor U21020 (N_21020,N_19868,N_18436);
nor U21021 (N_21021,N_19088,N_18392);
and U21022 (N_21022,N_18530,N_18342);
nor U21023 (N_21023,N_19101,N_18419);
nor U21024 (N_21024,N_19192,N_19436);
xnor U21025 (N_21025,N_19251,N_18998);
nor U21026 (N_21026,N_18665,N_19438);
xor U21027 (N_21027,N_19201,N_18625);
and U21028 (N_21028,N_18665,N_19623);
or U21029 (N_21029,N_19063,N_18221);
nor U21030 (N_21030,N_19379,N_18394);
or U21031 (N_21031,N_19933,N_19320);
xnor U21032 (N_21032,N_18709,N_19587);
nor U21033 (N_21033,N_18428,N_18452);
and U21034 (N_21034,N_18085,N_19725);
nand U21035 (N_21035,N_18581,N_18911);
xor U21036 (N_21036,N_19262,N_18841);
xnor U21037 (N_21037,N_18478,N_18578);
and U21038 (N_21038,N_19375,N_18688);
xor U21039 (N_21039,N_19347,N_19353);
nor U21040 (N_21040,N_19898,N_19902);
or U21041 (N_21041,N_19715,N_19709);
xnor U21042 (N_21042,N_19876,N_19711);
nand U21043 (N_21043,N_19455,N_19795);
xnor U21044 (N_21044,N_18232,N_18526);
nand U21045 (N_21045,N_19030,N_18554);
or U21046 (N_21046,N_19102,N_18815);
and U21047 (N_21047,N_18048,N_19268);
or U21048 (N_21048,N_18675,N_18402);
nor U21049 (N_21049,N_18793,N_19270);
nor U21050 (N_21050,N_18352,N_18765);
nand U21051 (N_21051,N_18217,N_19754);
xor U21052 (N_21052,N_18914,N_18935);
or U21053 (N_21053,N_18518,N_19382);
and U21054 (N_21054,N_18745,N_18240);
nor U21055 (N_21055,N_19221,N_19760);
nand U21056 (N_21056,N_19950,N_19002);
xor U21057 (N_21057,N_18773,N_18764);
xnor U21058 (N_21058,N_19318,N_19517);
or U21059 (N_21059,N_19504,N_18714);
nor U21060 (N_21060,N_19997,N_18014);
xor U21061 (N_21061,N_19968,N_19478);
or U21062 (N_21062,N_18112,N_18894);
nand U21063 (N_21063,N_18637,N_19721);
and U21064 (N_21064,N_19627,N_18768);
nor U21065 (N_21065,N_19860,N_18872);
or U21066 (N_21066,N_18171,N_18822);
and U21067 (N_21067,N_18555,N_19966);
and U21068 (N_21068,N_19426,N_18333);
and U21069 (N_21069,N_19355,N_19806);
nor U21070 (N_21070,N_18051,N_19516);
nor U21071 (N_21071,N_19569,N_18768);
or U21072 (N_21072,N_19568,N_19583);
and U21073 (N_21073,N_19712,N_19286);
nand U21074 (N_21074,N_18939,N_18374);
xor U21075 (N_21075,N_19684,N_18453);
and U21076 (N_21076,N_18278,N_19395);
xor U21077 (N_21077,N_19210,N_18783);
nor U21078 (N_21078,N_19474,N_18851);
nand U21079 (N_21079,N_18157,N_19723);
nor U21080 (N_21080,N_19491,N_19513);
and U21081 (N_21081,N_19467,N_18561);
nand U21082 (N_21082,N_18098,N_18642);
and U21083 (N_21083,N_19176,N_18455);
nand U21084 (N_21084,N_18214,N_18118);
nand U21085 (N_21085,N_18747,N_18669);
xor U21086 (N_21086,N_19104,N_18408);
xnor U21087 (N_21087,N_19595,N_18218);
nand U21088 (N_21088,N_19328,N_18037);
xor U21089 (N_21089,N_19939,N_19829);
xor U21090 (N_21090,N_18670,N_18738);
and U21091 (N_21091,N_19198,N_18081);
nand U21092 (N_21092,N_18315,N_19450);
nor U21093 (N_21093,N_19762,N_18150);
and U21094 (N_21094,N_19449,N_19322);
nor U21095 (N_21095,N_18668,N_18845);
and U21096 (N_21096,N_18255,N_19091);
xor U21097 (N_21097,N_19623,N_19417);
xor U21098 (N_21098,N_18412,N_18109);
or U21099 (N_21099,N_18888,N_18065);
or U21100 (N_21100,N_18850,N_19855);
or U21101 (N_21101,N_18971,N_19403);
nor U21102 (N_21102,N_19749,N_18183);
and U21103 (N_21103,N_19239,N_18840);
nor U21104 (N_21104,N_19236,N_18952);
and U21105 (N_21105,N_19818,N_19483);
xor U21106 (N_21106,N_19015,N_18257);
xnor U21107 (N_21107,N_19387,N_18810);
nor U21108 (N_21108,N_19436,N_19113);
nand U21109 (N_21109,N_19245,N_18108);
nor U21110 (N_21110,N_19705,N_19189);
xor U21111 (N_21111,N_18278,N_18113);
nand U21112 (N_21112,N_18302,N_18673);
xor U21113 (N_21113,N_18608,N_18845);
nor U21114 (N_21114,N_18977,N_18701);
nor U21115 (N_21115,N_19277,N_19844);
nand U21116 (N_21116,N_18480,N_19742);
nand U21117 (N_21117,N_18894,N_19329);
xnor U21118 (N_21118,N_18116,N_18713);
nand U21119 (N_21119,N_19653,N_18499);
nor U21120 (N_21120,N_19334,N_18989);
or U21121 (N_21121,N_19183,N_19882);
and U21122 (N_21122,N_19316,N_19429);
or U21123 (N_21123,N_19735,N_18883);
xnor U21124 (N_21124,N_18966,N_19792);
nor U21125 (N_21125,N_18263,N_18091);
nand U21126 (N_21126,N_19895,N_18352);
and U21127 (N_21127,N_18802,N_18582);
and U21128 (N_21128,N_19455,N_18237);
nor U21129 (N_21129,N_19503,N_19527);
xnor U21130 (N_21130,N_18670,N_19186);
xor U21131 (N_21131,N_18487,N_19073);
xor U21132 (N_21132,N_19053,N_19747);
or U21133 (N_21133,N_19803,N_19580);
or U21134 (N_21134,N_19503,N_18669);
nor U21135 (N_21135,N_18086,N_19307);
nor U21136 (N_21136,N_19551,N_18231);
nand U21137 (N_21137,N_19993,N_19384);
nand U21138 (N_21138,N_19270,N_19214);
xnor U21139 (N_21139,N_19227,N_18226);
or U21140 (N_21140,N_18297,N_19247);
and U21141 (N_21141,N_18780,N_18440);
nor U21142 (N_21142,N_18869,N_19780);
or U21143 (N_21143,N_19587,N_18006);
nor U21144 (N_21144,N_19150,N_18476);
or U21145 (N_21145,N_18028,N_18915);
xor U21146 (N_21146,N_19222,N_19961);
and U21147 (N_21147,N_19607,N_19520);
nor U21148 (N_21148,N_19961,N_19617);
or U21149 (N_21149,N_19327,N_18761);
xor U21150 (N_21150,N_18904,N_18956);
xor U21151 (N_21151,N_18459,N_19352);
xnor U21152 (N_21152,N_19577,N_18045);
xor U21153 (N_21153,N_19623,N_18586);
and U21154 (N_21154,N_18190,N_19557);
or U21155 (N_21155,N_19350,N_19053);
and U21156 (N_21156,N_19700,N_18417);
or U21157 (N_21157,N_18805,N_18695);
and U21158 (N_21158,N_18803,N_19133);
xor U21159 (N_21159,N_19794,N_18978);
xnor U21160 (N_21160,N_19403,N_19968);
and U21161 (N_21161,N_19688,N_18690);
nor U21162 (N_21162,N_18935,N_19636);
xnor U21163 (N_21163,N_18232,N_18544);
and U21164 (N_21164,N_19487,N_18947);
nor U21165 (N_21165,N_18967,N_19215);
nor U21166 (N_21166,N_19127,N_18020);
nor U21167 (N_21167,N_18557,N_18918);
and U21168 (N_21168,N_18226,N_19639);
xor U21169 (N_21169,N_19559,N_18772);
nand U21170 (N_21170,N_18289,N_19776);
nor U21171 (N_21171,N_19590,N_18099);
or U21172 (N_21172,N_19700,N_19499);
nor U21173 (N_21173,N_18513,N_19949);
and U21174 (N_21174,N_18788,N_19520);
nand U21175 (N_21175,N_18870,N_18481);
and U21176 (N_21176,N_18068,N_18254);
and U21177 (N_21177,N_19599,N_18996);
and U21178 (N_21178,N_18117,N_18870);
xnor U21179 (N_21179,N_18229,N_18794);
and U21180 (N_21180,N_18072,N_18121);
and U21181 (N_21181,N_18402,N_18285);
and U21182 (N_21182,N_19940,N_19951);
and U21183 (N_21183,N_19307,N_18922);
nor U21184 (N_21184,N_18871,N_18693);
nand U21185 (N_21185,N_19182,N_19435);
xnor U21186 (N_21186,N_18025,N_19529);
and U21187 (N_21187,N_19904,N_19900);
and U21188 (N_21188,N_18512,N_19285);
nor U21189 (N_21189,N_18484,N_19039);
or U21190 (N_21190,N_19670,N_18503);
xnor U21191 (N_21191,N_18786,N_19732);
xor U21192 (N_21192,N_18632,N_19460);
nand U21193 (N_21193,N_18954,N_19967);
nor U21194 (N_21194,N_19855,N_19164);
nand U21195 (N_21195,N_18509,N_19602);
nor U21196 (N_21196,N_18134,N_19241);
nor U21197 (N_21197,N_18155,N_19450);
nand U21198 (N_21198,N_18211,N_19068);
and U21199 (N_21199,N_18304,N_19220);
and U21200 (N_21200,N_18113,N_19527);
or U21201 (N_21201,N_18940,N_18507);
nand U21202 (N_21202,N_19897,N_19872);
or U21203 (N_21203,N_18434,N_19814);
xnor U21204 (N_21204,N_18464,N_18317);
xnor U21205 (N_21205,N_19009,N_18461);
xnor U21206 (N_21206,N_18761,N_19593);
nand U21207 (N_21207,N_18241,N_18279);
nand U21208 (N_21208,N_18687,N_19563);
xor U21209 (N_21209,N_19973,N_19584);
or U21210 (N_21210,N_19458,N_18047);
xor U21211 (N_21211,N_18067,N_19094);
nand U21212 (N_21212,N_18786,N_18810);
nor U21213 (N_21213,N_18913,N_18388);
and U21214 (N_21214,N_19469,N_18798);
nand U21215 (N_21215,N_18029,N_19381);
nand U21216 (N_21216,N_19545,N_18408);
and U21217 (N_21217,N_19376,N_18171);
nand U21218 (N_21218,N_18759,N_19139);
nor U21219 (N_21219,N_19555,N_18570);
or U21220 (N_21220,N_19820,N_19199);
or U21221 (N_21221,N_18792,N_19813);
and U21222 (N_21222,N_19990,N_18207);
xnor U21223 (N_21223,N_18834,N_19712);
or U21224 (N_21224,N_19655,N_19953);
nor U21225 (N_21225,N_19940,N_18579);
nand U21226 (N_21226,N_18639,N_19766);
xnor U21227 (N_21227,N_18576,N_18218);
and U21228 (N_21228,N_19908,N_19702);
xor U21229 (N_21229,N_18602,N_19809);
nand U21230 (N_21230,N_18797,N_18168);
xor U21231 (N_21231,N_18155,N_18272);
or U21232 (N_21232,N_18966,N_18087);
xnor U21233 (N_21233,N_19657,N_19804);
nor U21234 (N_21234,N_19451,N_19584);
and U21235 (N_21235,N_19795,N_19124);
and U21236 (N_21236,N_18479,N_19386);
nand U21237 (N_21237,N_19783,N_18911);
or U21238 (N_21238,N_18582,N_18344);
xnor U21239 (N_21239,N_19373,N_19767);
and U21240 (N_21240,N_19137,N_19808);
or U21241 (N_21241,N_18818,N_19937);
and U21242 (N_21242,N_19854,N_19650);
nand U21243 (N_21243,N_18972,N_18903);
or U21244 (N_21244,N_19753,N_19165);
nand U21245 (N_21245,N_18194,N_19753);
nor U21246 (N_21246,N_18536,N_18157);
xnor U21247 (N_21247,N_19934,N_19119);
nor U21248 (N_21248,N_19553,N_19364);
and U21249 (N_21249,N_19011,N_18480);
nor U21250 (N_21250,N_18413,N_18594);
xor U21251 (N_21251,N_19117,N_19683);
nor U21252 (N_21252,N_18099,N_18942);
nand U21253 (N_21253,N_19905,N_18771);
nand U21254 (N_21254,N_18306,N_19792);
nor U21255 (N_21255,N_18597,N_18412);
xor U21256 (N_21256,N_18580,N_18187);
nor U21257 (N_21257,N_19236,N_18430);
or U21258 (N_21258,N_18697,N_18733);
nand U21259 (N_21259,N_19599,N_18936);
and U21260 (N_21260,N_18008,N_18930);
and U21261 (N_21261,N_19320,N_18409);
xor U21262 (N_21262,N_18331,N_18157);
or U21263 (N_21263,N_19462,N_19176);
and U21264 (N_21264,N_18584,N_19683);
xor U21265 (N_21265,N_19245,N_19966);
nand U21266 (N_21266,N_19948,N_19318);
nor U21267 (N_21267,N_19857,N_19004);
nor U21268 (N_21268,N_19337,N_19625);
nor U21269 (N_21269,N_18703,N_18869);
nor U21270 (N_21270,N_18721,N_19028);
nand U21271 (N_21271,N_18604,N_18499);
and U21272 (N_21272,N_18520,N_19599);
xor U21273 (N_21273,N_19612,N_18740);
or U21274 (N_21274,N_18425,N_19434);
xnor U21275 (N_21275,N_19415,N_19646);
nor U21276 (N_21276,N_19300,N_19897);
or U21277 (N_21277,N_18624,N_18504);
and U21278 (N_21278,N_18389,N_19982);
nor U21279 (N_21279,N_18935,N_19571);
and U21280 (N_21280,N_19142,N_18967);
or U21281 (N_21281,N_18800,N_18863);
or U21282 (N_21282,N_18744,N_18948);
nand U21283 (N_21283,N_19107,N_19864);
and U21284 (N_21284,N_19078,N_18888);
xnor U21285 (N_21285,N_18965,N_18153);
or U21286 (N_21286,N_19829,N_19542);
and U21287 (N_21287,N_19086,N_19133);
or U21288 (N_21288,N_18304,N_18212);
and U21289 (N_21289,N_18415,N_19547);
and U21290 (N_21290,N_18388,N_18924);
nor U21291 (N_21291,N_19045,N_19981);
or U21292 (N_21292,N_18451,N_18686);
and U21293 (N_21293,N_18133,N_18447);
and U21294 (N_21294,N_19719,N_18432);
and U21295 (N_21295,N_19506,N_19524);
or U21296 (N_21296,N_18942,N_18491);
and U21297 (N_21297,N_18231,N_18356);
and U21298 (N_21298,N_18519,N_18175);
nand U21299 (N_21299,N_18336,N_18296);
nor U21300 (N_21300,N_19911,N_19596);
nand U21301 (N_21301,N_19440,N_18120);
nand U21302 (N_21302,N_18223,N_19079);
nand U21303 (N_21303,N_18581,N_18654);
nor U21304 (N_21304,N_19641,N_19161);
nand U21305 (N_21305,N_18611,N_18491);
xnor U21306 (N_21306,N_18872,N_18877);
xnor U21307 (N_21307,N_18394,N_19828);
nor U21308 (N_21308,N_19687,N_19619);
or U21309 (N_21309,N_18813,N_19788);
or U21310 (N_21310,N_19022,N_19488);
nor U21311 (N_21311,N_19118,N_19437);
or U21312 (N_21312,N_19580,N_18618);
xor U21313 (N_21313,N_19985,N_19617);
and U21314 (N_21314,N_18429,N_18141);
nor U21315 (N_21315,N_18919,N_19034);
and U21316 (N_21316,N_19679,N_18852);
nor U21317 (N_21317,N_19893,N_18297);
xor U21318 (N_21318,N_19594,N_18987);
or U21319 (N_21319,N_19636,N_18021);
or U21320 (N_21320,N_19532,N_18120);
xnor U21321 (N_21321,N_18395,N_19609);
and U21322 (N_21322,N_18607,N_19593);
nor U21323 (N_21323,N_19347,N_19646);
nor U21324 (N_21324,N_18121,N_18047);
nor U21325 (N_21325,N_18153,N_19738);
nor U21326 (N_21326,N_18259,N_18438);
nand U21327 (N_21327,N_19691,N_18828);
or U21328 (N_21328,N_18149,N_18220);
and U21329 (N_21329,N_19688,N_18138);
or U21330 (N_21330,N_19795,N_18581);
nor U21331 (N_21331,N_19231,N_19715);
xor U21332 (N_21332,N_18126,N_18303);
nand U21333 (N_21333,N_18909,N_19634);
or U21334 (N_21334,N_18269,N_19641);
nand U21335 (N_21335,N_18082,N_18681);
nand U21336 (N_21336,N_19854,N_18247);
xor U21337 (N_21337,N_19218,N_18787);
xnor U21338 (N_21338,N_18333,N_19594);
or U21339 (N_21339,N_19108,N_19557);
xor U21340 (N_21340,N_19334,N_19282);
and U21341 (N_21341,N_18106,N_19180);
and U21342 (N_21342,N_18477,N_18949);
nand U21343 (N_21343,N_19236,N_18003);
or U21344 (N_21344,N_18564,N_18692);
or U21345 (N_21345,N_18678,N_19253);
or U21346 (N_21346,N_19821,N_19895);
and U21347 (N_21347,N_19846,N_19906);
or U21348 (N_21348,N_18345,N_19608);
xor U21349 (N_21349,N_19284,N_18888);
and U21350 (N_21350,N_18808,N_18292);
and U21351 (N_21351,N_19338,N_18406);
xor U21352 (N_21352,N_19862,N_19149);
nor U21353 (N_21353,N_18248,N_18966);
or U21354 (N_21354,N_18699,N_18364);
or U21355 (N_21355,N_19536,N_18431);
and U21356 (N_21356,N_18345,N_19488);
xor U21357 (N_21357,N_19480,N_19470);
nor U21358 (N_21358,N_18348,N_19130);
nand U21359 (N_21359,N_18423,N_18831);
nand U21360 (N_21360,N_19761,N_18706);
and U21361 (N_21361,N_18454,N_18647);
nand U21362 (N_21362,N_19866,N_19815);
xor U21363 (N_21363,N_18003,N_18816);
and U21364 (N_21364,N_18464,N_19218);
xor U21365 (N_21365,N_19888,N_19989);
nand U21366 (N_21366,N_19433,N_18349);
xor U21367 (N_21367,N_18397,N_19099);
and U21368 (N_21368,N_19413,N_18305);
nand U21369 (N_21369,N_19814,N_19365);
or U21370 (N_21370,N_19319,N_19275);
nor U21371 (N_21371,N_19317,N_18488);
nand U21372 (N_21372,N_18478,N_18189);
or U21373 (N_21373,N_19632,N_18475);
nor U21374 (N_21374,N_19337,N_18040);
xor U21375 (N_21375,N_19051,N_18572);
or U21376 (N_21376,N_18191,N_18028);
xnor U21377 (N_21377,N_18340,N_18170);
nor U21378 (N_21378,N_19999,N_18410);
xor U21379 (N_21379,N_18459,N_18216);
nand U21380 (N_21380,N_19576,N_18732);
or U21381 (N_21381,N_18187,N_19549);
and U21382 (N_21382,N_19272,N_19553);
nor U21383 (N_21383,N_19810,N_19013);
and U21384 (N_21384,N_18797,N_18194);
and U21385 (N_21385,N_19696,N_19774);
nor U21386 (N_21386,N_18413,N_18682);
and U21387 (N_21387,N_19119,N_18891);
or U21388 (N_21388,N_18816,N_19009);
or U21389 (N_21389,N_18435,N_19332);
nand U21390 (N_21390,N_18288,N_18020);
nor U21391 (N_21391,N_19129,N_19986);
or U21392 (N_21392,N_18730,N_19357);
and U21393 (N_21393,N_19163,N_18868);
nor U21394 (N_21394,N_19268,N_19368);
and U21395 (N_21395,N_18021,N_18451);
or U21396 (N_21396,N_18028,N_18613);
nand U21397 (N_21397,N_18603,N_18677);
or U21398 (N_21398,N_19257,N_18873);
or U21399 (N_21399,N_19359,N_19523);
and U21400 (N_21400,N_19197,N_18678);
xor U21401 (N_21401,N_18183,N_18542);
and U21402 (N_21402,N_18768,N_18655);
xnor U21403 (N_21403,N_18638,N_18564);
xnor U21404 (N_21404,N_19844,N_19576);
nor U21405 (N_21405,N_18223,N_18890);
xor U21406 (N_21406,N_19581,N_18078);
or U21407 (N_21407,N_19109,N_18517);
nand U21408 (N_21408,N_18483,N_19525);
and U21409 (N_21409,N_19954,N_18105);
xor U21410 (N_21410,N_18617,N_18945);
xor U21411 (N_21411,N_18088,N_18515);
xor U21412 (N_21412,N_19533,N_18471);
nand U21413 (N_21413,N_19505,N_18065);
nand U21414 (N_21414,N_19774,N_18036);
nor U21415 (N_21415,N_18074,N_19063);
or U21416 (N_21416,N_18444,N_19650);
nor U21417 (N_21417,N_19339,N_19879);
or U21418 (N_21418,N_19885,N_18695);
or U21419 (N_21419,N_19498,N_18927);
xor U21420 (N_21420,N_18363,N_19654);
nand U21421 (N_21421,N_18668,N_19027);
nand U21422 (N_21422,N_19459,N_18770);
or U21423 (N_21423,N_19775,N_19618);
and U21424 (N_21424,N_18116,N_18268);
xor U21425 (N_21425,N_19694,N_18668);
nor U21426 (N_21426,N_19906,N_19629);
xnor U21427 (N_21427,N_19225,N_19756);
nor U21428 (N_21428,N_19289,N_18050);
xor U21429 (N_21429,N_18669,N_18703);
and U21430 (N_21430,N_19561,N_19597);
or U21431 (N_21431,N_18942,N_18972);
or U21432 (N_21432,N_19006,N_19098);
xnor U21433 (N_21433,N_18062,N_18549);
and U21434 (N_21434,N_18298,N_19404);
or U21435 (N_21435,N_19477,N_19290);
and U21436 (N_21436,N_18594,N_19005);
nand U21437 (N_21437,N_18488,N_18023);
nor U21438 (N_21438,N_18603,N_18531);
and U21439 (N_21439,N_18526,N_19653);
nor U21440 (N_21440,N_19322,N_18994);
nand U21441 (N_21441,N_18761,N_18609);
nor U21442 (N_21442,N_18137,N_19971);
nand U21443 (N_21443,N_18405,N_18118);
nand U21444 (N_21444,N_19064,N_18713);
and U21445 (N_21445,N_18947,N_18991);
and U21446 (N_21446,N_19417,N_18970);
and U21447 (N_21447,N_18459,N_19213);
and U21448 (N_21448,N_18702,N_18260);
or U21449 (N_21449,N_18805,N_18331);
nor U21450 (N_21450,N_18787,N_18838);
xnor U21451 (N_21451,N_19274,N_19298);
and U21452 (N_21452,N_19741,N_19465);
nor U21453 (N_21453,N_18297,N_18554);
or U21454 (N_21454,N_18016,N_18390);
xor U21455 (N_21455,N_18884,N_19516);
xor U21456 (N_21456,N_19899,N_18722);
xor U21457 (N_21457,N_19398,N_18643);
nand U21458 (N_21458,N_19853,N_18259);
nor U21459 (N_21459,N_18932,N_18426);
or U21460 (N_21460,N_19664,N_19571);
xnor U21461 (N_21461,N_19349,N_18000);
nor U21462 (N_21462,N_19533,N_18713);
nor U21463 (N_21463,N_19442,N_18871);
xor U21464 (N_21464,N_18690,N_19446);
or U21465 (N_21465,N_19149,N_19369);
xnor U21466 (N_21466,N_19364,N_18221);
or U21467 (N_21467,N_19260,N_19620);
nor U21468 (N_21468,N_19809,N_19122);
xor U21469 (N_21469,N_19697,N_19346);
nand U21470 (N_21470,N_19833,N_18570);
or U21471 (N_21471,N_19934,N_19162);
nor U21472 (N_21472,N_19949,N_19306);
nand U21473 (N_21473,N_19073,N_19712);
nand U21474 (N_21474,N_19933,N_19794);
xor U21475 (N_21475,N_18580,N_19375);
or U21476 (N_21476,N_18825,N_18301);
xnor U21477 (N_21477,N_18389,N_19325);
xnor U21478 (N_21478,N_18306,N_18824);
xnor U21479 (N_21479,N_19006,N_19481);
nor U21480 (N_21480,N_19988,N_19737);
nor U21481 (N_21481,N_19919,N_18190);
xor U21482 (N_21482,N_18308,N_19069);
xnor U21483 (N_21483,N_18094,N_18794);
and U21484 (N_21484,N_19302,N_18274);
nand U21485 (N_21485,N_19029,N_19721);
xor U21486 (N_21486,N_18995,N_19792);
or U21487 (N_21487,N_19286,N_18957);
or U21488 (N_21488,N_18182,N_19240);
nand U21489 (N_21489,N_18791,N_18389);
or U21490 (N_21490,N_18358,N_18090);
nor U21491 (N_21491,N_18393,N_19074);
and U21492 (N_21492,N_19481,N_19754);
xor U21493 (N_21493,N_19345,N_18851);
or U21494 (N_21494,N_19309,N_19298);
or U21495 (N_21495,N_18521,N_18640);
nor U21496 (N_21496,N_19241,N_19765);
nor U21497 (N_21497,N_18742,N_18448);
and U21498 (N_21498,N_19196,N_18128);
nand U21499 (N_21499,N_18470,N_18223);
nor U21500 (N_21500,N_19817,N_18292);
xor U21501 (N_21501,N_19606,N_19778);
nand U21502 (N_21502,N_19908,N_19893);
xnor U21503 (N_21503,N_19776,N_18105);
nand U21504 (N_21504,N_18209,N_18701);
nor U21505 (N_21505,N_18802,N_18818);
and U21506 (N_21506,N_19151,N_19338);
nand U21507 (N_21507,N_18975,N_18822);
and U21508 (N_21508,N_18885,N_19776);
nor U21509 (N_21509,N_19695,N_19525);
nand U21510 (N_21510,N_18753,N_18016);
nor U21511 (N_21511,N_19547,N_19844);
xnor U21512 (N_21512,N_18862,N_19943);
xnor U21513 (N_21513,N_19533,N_19906);
nand U21514 (N_21514,N_18694,N_18842);
xnor U21515 (N_21515,N_18280,N_18809);
nor U21516 (N_21516,N_18278,N_19340);
and U21517 (N_21517,N_19860,N_19639);
or U21518 (N_21518,N_18428,N_19000);
nor U21519 (N_21519,N_18854,N_18800);
and U21520 (N_21520,N_19812,N_19093);
or U21521 (N_21521,N_18386,N_19671);
nand U21522 (N_21522,N_19371,N_18632);
xor U21523 (N_21523,N_18559,N_18931);
or U21524 (N_21524,N_18644,N_18277);
nand U21525 (N_21525,N_18566,N_18193);
xor U21526 (N_21526,N_19800,N_18116);
nor U21527 (N_21527,N_19852,N_18510);
or U21528 (N_21528,N_19103,N_19268);
nor U21529 (N_21529,N_18768,N_19764);
nand U21530 (N_21530,N_18083,N_19220);
nor U21531 (N_21531,N_18302,N_18632);
nand U21532 (N_21532,N_19037,N_19879);
nand U21533 (N_21533,N_19393,N_18337);
nand U21534 (N_21534,N_18239,N_18595);
or U21535 (N_21535,N_18700,N_18293);
nor U21536 (N_21536,N_19775,N_19347);
or U21537 (N_21537,N_19008,N_18989);
or U21538 (N_21538,N_19670,N_19802);
nor U21539 (N_21539,N_19084,N_19897);
and U21540 (N_21540,N_19348,N_19001);
nor U21541 (N_21541,N_19435,N_19253);
xor U21542 (N_21542,N_18304,N_18708);
nor U21543 (N_21543,N_18886,N_19389);
xnor U21544 (N_21544,N_18637,N_18620);
nand U21545 (N_21545,N_18184,N_19620);
nand U21546 (N_21546,N_18845,N_18304);
xor U21547 (N_21547,N_18721,N_19006);
or U21548 (N_21548,N_18984,N_19690);
xor U21549 (N_21549,N_18877,N_19557);
nor U21550 (N_21550,N_18343,N_18383);
nor U21551 (N_21551,N_19859,N_18366);
nor U21552 (N_21552,N_19812,N_19289);
and U21553 (N_21553,N_18715,N_18279);
or U21554 (N_21554,N_18234,N_18049);
or U21555 (N_21555,N_19927,N_18834);
or U21556 (N_21556,N_19694,N_19740);
nand U21557 (N_21557,N_19397,N_18967);
nor U21558 (N_21558,N_19551,N_18502);
or U21559 (N_21559,N_19983,N_19729);
nand U21560 (N_21560,N_18147,N_19054);
or U21561 (N_21561,N_18014,N_19594);
and U21562 (N_21562,N_19673,N_18408);
or U21563 (N_21563,N_18732,N_18086);
nor U21564 (N_21564,N_18689,N_18156);
xor U21565 (N_21565,N_18319,N_18754);
and U21566 (N_21566,N_19683,N_18095);
or U21567 (N_21567,N_19721,N_19513);
nand U21568 (N_21568,N_18804,N_19460);
or U21569 (N_21569,N_19030,N_18440);
or U21570 (N_21570,N_19634,N_18885);
xnor U21571 (N_21571,N_18917,N_19188);
nor U21572 (N_21572,N_18841,N_18779);
xor U21573 (N_21573,N_18692,N_19423);
and U21574 (N_21574,N_18670,N_19651);
xor U21575 (N_21575,N_18929,N_19856);
or U21576 (N_21576,N_18565,N_18853);
or U21577 (N_21577,N_19711,N_18538);
nand U21578 (N_21578,N_19504,N_19161);
nor U21579 (N_21579,N_18988,N_18342);
nor U21580 (N_21580,N_18137,N_18124);
nor U21581 (N_21581,N_19344,N_18215);
and U21582 (N_21582,N_18136,N_18668);
xor U21583 (N_21583,N_18023,N_19240);
or U21584 (N_21584,N_18948,N_19917);
xor U21585 (N_21585,N_19298,N_19525);
nand U21586 (N_21586,N_19857,N_19772);
or U21587 (N_21587,N_18979,N_18164);
and U21588 (N_21588,N_19861,N_19454);
xor U21589 (N_21589,N_18650,N_18290);
and U21590 (N_21590,N_18168,N_19976);
nand U21591 (N_21591,N_19978,N_18832);
nand U21592 (N_21592,N_19259,N_18986);
and U21593 (N_21593,N_18641,N_19154);
or U21594 (N_21594,N_18874,N_18457);
and U21595 (N_21595,N_19860,N_19886);
or U21596 (N_21596,N_18486,N_18798);
xor U21597 (N_21597,N_19593,N_18339);
or U21598 (N_21598,N_19327,N_18565);
and U21599 (N_21599,N_18285,N_19826);
nor U21600 (N_21600,N_18963,N_18267);
nand U21601 (N_21601,N_19347,N_18410);
nor U21602 (N_21602,N_18666,N_18078);
nand U21603 (N_21603,N_18340,N_18665);
or U21604 (N_21604,N_19007,N_18256);
nand U21605 (N_21605,N_19059,N_19749);
nand U21606 (N_21606,N_19804,N_18985);
nor U21607 (N_21607,N_19923,N_18664);
or U21608 (N_21608,N_19584,N_19812);
nor U21609 (N_21609,N_18228,N_18666);
nor U21610 (N_21610,N_18474,N_18944);
or U21611 (N_21611,N_18585,N_18777);
or U21612 (N_21612,N_19824,N_18103);
xor U21613 (N_21613,N_18452,N_18369);
xor U21614 (N_21614,N_18553,N_18587);
and U21615 (N_21615,N_19897,N_18562);
or U21616 (N_21616,N_18821,N_19403);
nor U21617 (N_21617,N_19217,N_18032);
nor U21618 (N_21618,N_18228,N_18752);
or U21619 (N_21619,N_18329,N_18220);
xnor U21620 (N_21620,N_19922,N_19531);
or U21621 (N_21621,N_19713,N_18355);
or U21622 (N_21622,N_19671,N_18167);
nor U21623 (N_21623,N_19312,N_18892);
and U21624 (N_21624,N_18093,N_19347);
nand U21625 (N_21625,N_19276,N_18356);
xnor U21626 (N_21626,N_18531,N_19765);
nand U21627 (N_21627,N_18302,N_18930);
nand U21628 (N_21628,N_19790,N_19585);
nand U21629 (N_21629,N_19502,N_19397);
nor U21630 (N_21630,N_19565,N_19239);
nor U21631 (N_21631,N_18288,N_19638);
and U21632 (N_21632,N_18118,N_18669);
or U21633 (N_21633,N_18162,N_18359);
xnor U21634 (N_21634,N_19833,N_19937);
nand U21635 (N_21635,N_18465,N_19653);
xnor U21636 (N_21636,N_19228,N_19605);
or U21637 (N_21637,N_19865,N_19672);
or U21638 (N_21638,N_19710,N_18267);
nor U21639 (N_21639,N_18758,N_18458);
and U21640 (N_21640,N_18257,N_18104);
nor U21641 (N_21641,N_19709,N_18389);
nor U21642 (N_21642,N_19809,N_19619);
or U21643 (N_21643,N_19315,N_19945);
nand U21644 (N_21644,N_18884,N_19650);
xor U21645 (N_21645,N_19687,N_19970);
nand U21646 (N_21646,N_18091,N_19378);
nand U21647 (N_21647,N_18005,N_19023);
nor U21648 (N_21648,N_18204,N_19070);
nor U21649 (N_21649,N_18357,N_19379);
xnor U21650 (N_21650,N_19460,N_19949);
nor U21651 (N_21651,N_18158,N_19281);
nor U21652 (N_21652,N_19535,N_19123);
and U21653 (N_21653,N_19437,N_18848);
nor U21654 (N_21654,N_18528,N_19976);
and U21655 (N_21655,N_18035,N_18753);
nor U21656 (N_21656,N_19858,N_18333);
nor U21657 (N_21657,N_18806,N_18652);
nor U21658 (N_21658,N_18202,N_19543);
and U21659 (N_21659,N_19180,N_19518);
and U21660 (N_21660,N_18958,N_18702);
nor U21661 (N_21661,N_19634,N_19129);
or U21662 (N_21662,N_18773,N_19072);
and U21663 (N_21663,N_19150,N_19705);
or U21664 (N_21664,N_19104,N_19631);
nand U21665 (N_21665,N_19355,N_18674);
nor U21666 (N_21666,N_18232,N_18582);
and U21667 (N_21667,N_19161,N_19999);
xor U21668 (N_21668,N_18237,N_19873);
nand U21669 (N_21669,N_18011,N_19667);
or U21670 (N_21670,N_18303,N_18409);
and U21671 (N_21671,N_19004,N_18270);
and U21672 (N_21672,N_18963,N_18274);
and U21673 (N_21673,N_19466,N_18326);
or U21674 (N_21674,N_19457,N_19528);
or U21675 (N_21675,N_19735,N_18448);
nand U21676 (N_21676,N_18384,N_19828);
nand U21677 (N_21677,N_18846,N_18767);
nor U21678 (N_21678,N_18825,N_18216);
and U21679 (N_21679,N_18590,N_19028);
and U21680 (N_21680,N_19090,N_19398);
xnor U21681 (N_21681,N_19787,N_19351);
nor U21682 (N_21682,N_18009,N_19894);
nor U21683 (N_21683,N_19215,N_18738);
nor U21684 (N_21684,N_19325,N_19034);
nand U21685 (N_21685,N_18373,N_18740);
and U21686 (N_21686,N_18262,N_18501);
xor U21687 (N_21687,N_19828,N_18795);
xnor U21688 (N_21688,N_19798,N_19259);
or U21689 (N_21689,N_18500,N_18952);
or U21690 (N_21690,N_19780,N_18520);
and U21691 (N_21691,N_18009,N_18274);
xnor U21692 (N_21692,N_19752,N_19175);
or U21693 (N_21693,N_19242,N_19088);
nand U21694 (N_21694,N_18792,N_18552);
and U21695 (N_21695,N_18754,N_19661);
nand U21696 (N_21696,N_18501,N_18429);
nand U21697 (N_21697,N_19049,N_19196);
nor U21698 (N_21698,N_19990,N_19385);
xnor U21699 (N_21699,N_19786,N_18839);
or U21700 (N_21700,N_18404,N_18682);
nor U21701 (N_21701,N_18253,N_19913);
or U21702 (N_21702,N_19858,N_18861);
or U21703 (N_21703,N_19350,N_18433);
or U21704 (N_21704,N_19258,N_19430);
xnor U21705 (N_21705,N_18820,N_18246);
and U21706 (N_21706,N_19139,N_18991);
and U21707 (N_21707,N_18356,N_19587);
and U21708 (N_21708,N_19453,N_19889);
and U21709 (N_21709,N_18461,N_18503);
xor U21710 (N_21710,N_18542,N_19547);
and U21711 (N_21711,N_18255,N_19544);
xnor U21712 (N_21712,N_19290,N_19003);
or U21713 (N_21713,N_18656,N_19928);
nand U21714 (N_21714,N_18747,N_19829);
and U21715 (N_21715,N_18003,N_18421);
or U21716 (N_21716,N_19112,N_19320);
nor U21717 (N_21717,N_18552,N_18315);
nor U21718 (N_21718,N_19130,N_19093);
or U21719 (N_21719,N_18910,N_19261);
or U21720 (N_21720,N_18013,N_18755);
nor U21721 (N_21721,N_18166,N_19133);
nand U21722 (N_21722,N_18233,N_19072);
or U21723 (N_21723,N_18396,N_19528);
xor U21724 (N_21724,N_19299,N_19154);
nand U21725 (N_21725,N_19121,N_18303);
and U21726 (N_21726,N_19469,N_18055);
or U21727 (N_21727,N_19067,N_19164);
or U21728 (N_21728,N_19665,N_19245);
nor U21729 (N_21729,N_19555,N_19955);
nand U21730 (N_21730,N_18265,N_18592);
or U21731 (N_21731,N_18002,N_18776);
nand U21732 (N_21732,N_19569,N_19664);
nand U21733 (N_21733,N_19922,N_19595);
nor U21734 (N_21734,N_19756,N_18284);
and U21735 (N_21735,N_19729,N_18349);
nand U21736 (N_21736,N_18035,N_18652);
or U21737 (N_21737,N_19508,N_18573);
and U21738 (N_21738,N_18033,N_18158);
and U21739 (N_21739,N_18144,N_19226);
or U21740 (N_21740,N_19649,N_18995);
and U21741 (N_21741,N_19952,N_18156);
xnor U21742 (N_21742,N_19854,N_19554);
and U21743 (N_21743,N_18766,N_19238);
xnor U21744 (N_21744,N_18032,N_18533);
nor U21745 (N_21745,N_19328,N_19864);
nand U21746 (N_21746,N_18116,N_19916);
xnor U21747 (N_21747,N_18442,N_19185);
xnor U21748 (N_21748,N_18921,N_19801);
or U21749 (N_21749,N_19351,N_18774);
xor U21750 (N_21750,N_19783,N_18369);
xnor U21751 (N_21751,N_18468,N_18598);
nand U21752 (N_21752,N_19139,N_19669);
nand U21753 (N_21753,N_19981,N_18047);
xor U21754 (N_21754,N_18131,N_19421);
nand U21755 (N_21755,N_19649,N_18584);
xnor U21756 (N_21756,N_19122,N_18160);
or U21757 (N_21757,N_19086,N_18383);
or U21758 (N_21758,N_18545,N_19374);
or U21759 (N_21759,N_19785,N_18708);
nor U21760 (N_21760,N_19625,N_19382);
or U21761 (N_21761,N_18250,N_18738);
xor U21762 (N_21762,N_18232,N_19509);
and U21763 (N_21763,N_18931,N_19924);
and U21764 (N_21764,N_19407,N_19283);
or U21765 (N_21765,N_18013,N_18719);
or U21766 (N_21766,N_19449,N_18968);
or U21767 (N_21767,N_19794,N_19716);
xnor U21768 (N_21768,N_18114,N_18792);
nor U21769 (N_21769,N_18281,N_19075);
or U21770 (N_21770,N_18888,N_18509);
nor U21771 (N_21771,N_18595,N_19715);
nor U21772 (N_21772,N_19391,N_18102);
or U21773 (N_21773,N_19901,N_19352);
nand U21774 (N_21774,N_19772,N_19110);
or U21775 (N_21775,N_18347,N_18563);
and U21776 (N_21776,N_18993,N_18466);
nand U21777 (N_21777,N_19185,N_19590);
xnor U21778 (N_21778,N_18967,N_19689);
nor U21779 (N_21779,N_19268,N_18361);
nand U21780 (N_21780,N_18092,N_18954);
or U21781 (N_21781,N_19856,N_18336);
nor U21782 (N_21782,N_18170,N_18132);
or U21783 (N_21783,N_18660,N_19314);
or U21784 (N_21784,N_19729,N_19421);
nand U21785 (N_21785,N_18608,N_19496);
xor U21786 (N_21786,N_19412,N_18404);
nand U21787 (N_21787,N_18089,N_18357);
nand U21788 (N_21788,N_18545,N_18821);
nand U21789 (N_21789,N_18296,N_18244);
or U21790 (N_21790,N_18884,N_18889);
xnor U21791 (N_21791,N_18678,N_19006);
xnor U21792 (N_21792,N_19209,N_19720);
xnor U21793 (N_21793,N_18409,N_19334);
or U21794 (N_21794,N_19666,N_18395);
and U21795 (N_21795,N_18340,N_19970);
or U21796 (N_21796,N_19081,N_18884);
nor U21797 (N_21797,N_19766,N_19217);
or U21798 (N_21798,N_19403,N_19495);
xnor U21799 (N_21799,N_18878,N_19558);
and U21800 (N_21800,N_19282,N_19131);
nor U21801 (N_21801,N_19701,N_19485);
or U21802 (N_21802,N_19540,N_19737);
nor U21803 (N_21803,N_18828,N_19932);
and U21804 (N_21804,N_19639,N_19740);
and U21805 (N_21805,N_18037,N_18923);
xnor U21806 (N_21806,N_18722,N_19073);
or U21807 (N_21807,N_19143,N_18095);
nand U21808 (N_21808,N_19049,N_18008);
xnor U21809 (N_21809,N_18695,N_18064);
xnor U21810 (N_21810,N_19486,N_19307);
and U21811 (N_21811,N_18560,N_18741);
or U21812 (N_21812,N_18392,N_19318);
nand U21813 (N_21813,N_19613,N_18782);
or U21814 (N_21814,N_19040,N_19904);
xnor U21815 (N_21815,N_19481,N_19789);
and U21816 (N_21816,N_18219,N_19014);
nor U21817 (N_21817,N_18507,N_19368);
and U21818 (N_21818,N_19793,N_19243);
xnor U21819 (N_21819,N_18456,N_18158);
and U21820 (N_21820,N_18714,N_19581);
xnor U21821 (N_21821,N_18218,N_18286);
xor U21822 (N_21822,N_19065,N_19396);
or U21823 (N_21823,N_18547,N_19145);
nand U21824 (N_21824,N_18673,N_19636);
or U21825 (N_21825,N_19792,N_19211);
and U21826 (N_21826,N_18561,N_18219);
or U21827 (N_21827,N_19938,N_19512);
and U21828 (N_21828,N_18708,N_18997);
and U21829 (N_21829,N_19010,N_19666);
or U21830 (N_21830,N_18874,N_19950);
and U21831 (N_21831,N_18048,N_19540);
nor U21832 (N_21832,N_18494,N_19408);
xnor U21833 (N_21833,N_18001,N_18073);
nor U21834 (N_21834,N_18663,N_18073);
or U21835 (N_21835,N_19389,N_19339);
or U21836 (N_21836,N_19183,N_18001);
nand U21837 (N_21837,N_18109,N_18535);
and U21838 (N_21838,N_18235,N_19126);
xor U21839 (N_21839,N_18206,N_19475);
nand U21840 (N_21840,N_18092,N_18207);
or U21841 (N_21841,N_18406,N_18112);
and U21842 (N_21842,N_18485,N_18755);
nand U21843 (N_21843,N_18382,N_18027);
nor U21844 (N_21844,N_18871,N_19137);
nand U21845 (N_21845,N_19066,N_19672);
or U21846 (N_21846,N_18599,N_19775);
nand U21847 (N_21847,N_18915,N_18284);
and U21848 (N_21848,N_19702,N_19759);
and U21849 (N_21849,N_18506,N_19744);
and U21850 (N_21850,N_18213,N_18287);
nand U21851 (N_21851,N_19024,N_19872);
nand U21852 (N_21852,N_18507,N_18641);
nand U21853 (N_21853,N_19943,N_19552);
nand U21854 (N_21854,N_18602,N_18481);
xnor U21855 (N_21855,N_19812,N_18576);
and U21856 (N_21856,N_19582,N_19860);
nor U21857 (N_21857,N_18938,N_19596);
or U21858 (N_21858,N_18403,N_18419);
or U21859 (N_21859,N_18453,N_19388);
xor U21860 (N_21860,N_18080,N_19188);
nor U21861 (N_21861,N_19873,N_19288);
nor U21862 (N_21862,N_18569,N_19141);
and U21863 (N_21863,N_19766,N_18219);
xor U21864 (N_21864,N_19779,N_18770);
and U21865 (N_21865,N_19991,N_18176);
or U21866 (N_21866,N_19678,N_19966);
nor U21867 (N_21867,N_18009,N_19825);
nor U21868 (N_21868,N_18359,N_19035);
xor U21869 (N_21869,N_19650,N_19703);
nand U21870 (N_21870,N_19301,N_19251);
nor U21871 (N_21871,N_19652,N_18351);
nor U21872 (N_21872,N_19900,N_19570);
and U21873 (N_21873,N_19023,N_19705);
xor U21874 (N_21874,N_18947,N_19962);
xnor U21875 (N_21875,N_18338,N_19175);
and U21876 (N_21876,N_19591,N_18968);
or U21877 (N_21877,N_18472,N_18730);
nor U21878 (N_21878,N_19176,N_19972);
or U21879 (N_21879,N_19911,N_19972);
nand U21880 (N_21880,N_18781,N_19668);
or U21881 (N_21881,N_19912,N_18684);
nor U21882 (N_21882,N_18269,N_18228);
xnor U21883 (N_21883,N_19377,N_19378);
nand U21884 (N_21884,N_19609,N_19852);
and U21885 (N_21885,N_18301,N_19992);
or U21886 (N_21886,N_18803,N_19176);
nor U21887 (N_21887,N_19889,N_19675);
xor U21888 (N_21888,N_18354,N_18413);
and U21889 (N_21889,N_18308,N_18919);
nand U21890 (N_21890,N_18102,N_18631);
or U21891 (N_21891,N_19169,N_19216);
and U21892 (N_21892,N_19772,N_18666);
nor U21893 (N_21893,N_18766,N_18022);
and U21894 (N_21894,N_19584,N_19907);
nor U21895 (N_21895,N_19019,N_19397);
and U21896 (N_21896,N_19710,N_18365);
nand U21897 (N_21897,N_18340,N_19600);
nor U21898 (N_21898,N_18583,N_19880);
and U21899 (N_21899,N_19233,N_18778);
nor U21900 (N_21900,N_19686,N_19377);
and U21901 (N_21901,N_18860,N_19636);
xor U21902 (N_21902,N_19234,N_18389);
nor U21903 (N_21903,N_18276,N_19565);
xnor U21904 (N_21904,N_19286,N_18537);
nor U21905 (N_21905,N_19842,N_19688);
and U21906 (N_21906,N_18795,N_18267);
or U21907 (N_21907,N_19491,N_19214);
nor U21908 (N_21908,N_18233,N_19286);
nand U21909 (N_21909,N_18843,N_18596);
or U21910 (N_21910,N_19718,N_19852);
nand U21911 (N_21911,N_19903,N_19461);
and U21912 (N_21912,N_19796,N_18726);
and U21913 (N_21913,N_18102,N_18499);
or U21914 (N_21914,N_19645,N_19741);
and U21915 (N_21915,N_19262,N_19854);
or U21916 (N_21916,N_18697,N_19399);
nand U21917 (N_21917,N_19983,N_19692);
xnor U21918 (N_21918,N_19130,N_18043);
xor U21919 (N_21919,N_19100,N_18824);
and U21920 (N_21920,N_19172,N_18446);
nand U21921 (N_21921,N_18661,N_18364);
nor U21922 (N_21922,N_18499,N_18157);
nand U21923 (N_21923,N_19347,N_18532);
or U21924 (N_21924,N_18303,N_18330);
or U21925 (N_21925,N_19631,N_19429);
and U21926 (N_21926,N_18816,N_18136);
and U21927 (N_21927,N_19227,N_18783);
nor U21928 (N_21928,N_19583,N_19483);
nand U21929 (N_21929,N_18912,N_19391);
xor U21930 (N_21930,N_19054,N_19079);
nand U21931 (N_21931,N_19408,N_18486);
and U21932 (N_21932,N_19652,N_18345);
or U21933 (N_21933,N_19887,N_18242);
xor U21934 (N_21934,N_18755,N_19798);
xor U21935 (N_21935,N_19528,N_18341);
nor U21936 (N_21936,N_19312,N_18400);
nand U21937 (N_21937,N_19304,N_19806);
nand U21938 (N_21938,N_19776,N_18947);
and U21939 (N_21939,N_19412,N_18973);
nor U21940 (N_21940,N_18534,N_19730);
nand U21941 (N_21941,N_19070,N_18737);
and U21942 (N_21942,N_18355,N_18338);
and U21943 (N_21943,N_19321,N_19080);
nor U21944 (N_21944,N_19860,N_19349);
nor U21945 (N_21945,N_18100,N_18265);
or U21946 (N_21946,N_19467,N_18800);
xor U21947 (N_21947,N_19233,N_19343);
nand U21948 (N_21948,N_18129,N_19112);
and U21949 (N_21949,N_19785,N_19934);
xor U21950 (N_21950,N_19821,N_19413);
nand U21951 (N_21951,N_18757,N_18429);
and U21952 (N_21952,N_18541,N_19246);
or U21953 (N_21953,N_19262,N_19679);
or U21954 (N_21954,N_19661,N_18371);
xor U21955 (N_21955,N_19299,N_18476);
nand U21956 (N_21956,N_19014,N_19928);
nor U21957 (N_21957,N_18521,N_18507);
or U21958 (N_21958,N_19422,N_19703);
nor U21959 (N_21959,N_18226,N_18591);
xor U21960 (N_21960,N_19878,N_19596);
nand U21961 (N_21961,N_19521,N_18408);
nand U21962 (N_21962,N_18340,N_19275);
nand U21963 (N_21963,N_19640,N_18791);
nor U21964 (N_21964,N_18458,N_18388);
nor U21965 (N_21965,N_19281,N_19769);
nor U21966 (N_21966,N_18178,N_18795);
nand U21967 (N_21967,N_18808,N_18598);
nand U21968 (N_21968,N_19369,N_18706);
nor U21969 (N_21969,N_19536,N_19183);
and U21970 (N_21970,N_18249,N_19858);
or U21971 (N_21971,N_18091,N_19554);
and U21972 (N_21972,N_19673,N_18318);
or U21973 (N_21973,N_18446,N_18275);
xnor U21974 (N_21974,N_19092,N_19748);
xor U21975 (N_21975,N_18595,N_19717);
nand U21976 (N_21976,N_19049,N_18883);
nand U21977 (N_21977,N_19847,N_19665);
nor U21978 (N_21978,N_18721,N_19597);
and U21979 (N_21979,N_18343,N_18606);
nor U21980 (N_21980,N_18813,N_18283);
or U21981 (N_21981,N_18596,N_19495);
and U21982 (N_21982,N_19092,N_19256);
nor U21983 (N_21983,N_19471,N_18092);
and U21984 (N_21984,N_19368,N_19677);
xor U21985 (N_21985,N_18648,N_18728);
xor U21986 (N_21986,N_18920,N_19067);
and U21987 (N_21987,N_19758,N_18567);
xor U21988 (N_21988,N_19369,N_18262);
nand U21989 (N_21989,N_18047,N_18815);
or U21990 (N_21990,N_18044,N_18743);
xor U21991 (N_21991,N_19191,N_18707);
and U21992 (N_21992,N_18118,N_18070);
or U21993 (N_21993,N_19154,N_19435);
xnor U21994 (N_21994,N_18031,N_18407);
xnor U21995 (N_21995,N_18622,N_18667);
xor U21996 (N_21996,N_19721,N_19792);
xor U21997 (N_21997,N_18809,N_19968);
nand U21998 (N_21998,N_19292,N_18510);
xor U21999 (N_21999,N_19040,N_19099);
xnor U22000 (N_22000,N_21530,N_21147);
nor U22001 (N_22001,N_20445,N_20094);
nor U22002 (N_22002,N_20735,N_21304);
or U22003 (N_22003,N_21712,N_21048);
and U22004 (N_22004,N_21829,N_21312);
and U22005 (N_22005,N_20521,N_21746);
xor U22006 (N_22006,N_20157,N_21945);
or U22007 (N_22007,N_21768,N_21191);
and U22008 (N_22008,N_20655,N_20064);
nor U22009 (N_22009,N_20344,N_21799);
and U22010 (N_22010,N_20612,N_21810);
nand U22011 (N_22011,N_21627,N_21558);
nor U22012 (N_22012,N_20252,N_21729);
and U22013 (N_22013,N_20328,N_21473);
or U22014 (N_22014,N_20163,N_21106);
xnor U22015 (N_22015,N_20600,N_20489);
or U22016 (N_22016,N_21672,N_20678);
nor U22017 (N_22017,N_20817,N_20305);
nor U22018 (N_22018,N_21371,N_21244);
xnor U22019 (N_22019,N_21287,N_20066);
xor U22020 (N_22020,N_21347,N_20824);
nand U22021 (N_22021,N_20485,N_21600);
nor U22022 (N_22022,N_21130,N_20090);
or U22023 (N_22023,N_20581,N_20029);
xnor U22024 (N_22024,N_21029,N_21008);
nor U22025 (N_22025,N_20730,N_21210);
xor U22026 (N_22026,N_20766,N_20729);
or U22027 (N_22027,N_20725,N_20870);
and U22028 (N_22028,N_20342,N_21784);
or U22029 (N_22029,N_20892,N_21777);
nand U22030 (N_22030,N_20403,N_21960);
or U22031 (N_22031,N_21961,N_20830);
nand U22032 (N_22032,N_20625,N_20452);
nor U22033 (N_22033,N_20933,N_20013);
or U22034 (N_22034,N_20851,N_21930);
nor U22035 (N_22035,N_20818,N_21767);
nor U22036 (N_22036,N_21441,N_20126);
nor U22037 (N_22037,N_21389,N_20578);
or U22038 (N_22038,N_21061,N_20311);
nand U22039 (N_22039,N_20137,N_20756);
and U22040 (N_22040,N_21384,N_21894);
and U22041 (N_22041,N_21741,N_20596);
nor U22042 (N_22042,N_21516,N_21397);
nand U22043 (N_22043,N_20535,N_21694);
nand U22044 (N_22044,N_21276,N_21895);
or U22045 (N_22045,N_21013,N_21332);
xnor U22046 (N_22046,N_20855,N_21149);
xnor U22047 (N_22047,N_20147,N_21495);
or U22048 (N_22048,N_21203,N_20886);
and U22049 (N_22049,N_20303,N_20865);
and U22050 (N_22050,N_21725,N_21719);
nor U22051 (N_22051,N_21436,N_21372);
and U22052 (N_22052,N_21947,N_21797);
or U22053 (N_22053,N_20666,N_20661);
nand U22054 (N_22054,N_21238,N_21080);
and U22055 (N_22055,N_20041,N_21185);
xor U22056 (N_22056,N_20691,N_21569);
nand U22057 (N_22057,N_20832,N_20911);
xor U22058 (N_22058,N_20574,N_20503);
nand U22059 (N_22059,N_20474,N_21306);
nor U22060 (N_22060,N_21630,N_20772);
or U22061 (N_22061,N_21584,N_20367);
xor U22062 (N_22062,N_21903,N_21907);
xnor U22063 (N_22063,N_20968,N_21990);
and U22064 (N_22064,N_20940,N_21366);
xnor U22065 (N_22065,N_20358,N_21124);
nand U22066 (N_22066,N_20821,N_21370);
and U22067 (N_22067,N_20261,N_20633);
xnor U22068 (N_22068,N_20123,N_20321);
xor U22069 (N_22069,N_21993,N_21419);
nor U22070 (N_22070,N_21261,N_20250);
nand U22071 (N_22071,N_20944,N_20917);
and U22072 (N_22072,N_20055,N_20942);
xor U22073 (N_22073,N_21740,N_21240);
or U22074 (N_22074,N_21406,N_20042);
nand U22075 (N_22075,N_20547,N_20369);
or U22076 (N_22076,N_21074,N_21009);
and U22077 (N_22077,N_21246,N_21489);
and U22078 (N_22078,N_20693,N_21771);
nand U22079 (N_22079,N_21103,N_21085);
nand U22080 (N_22080,N_20816,N_20466);
xnor U22081 (N_22081,N_21598,N_20400);
and U22082 (N_22082,N_20105,N_20254);
and U22083 (N_22083,N_21296,N_20120);
xnor U22084 (N_22084,N_21926,N_21293);
or U22085 (N_22085,N_20195,N_21423);
or U22086 (N_22086,N_20523,N_21802);
nor U22087 (N_22087,N_21125,N_20813);
xnor U22088 (N_22088,N_20896,N_21579);
nand U22089 (N_22089,N_21018,N_21588);
xnor U22090 (N_22090,N_20138,N_21565);
xnor U22091 (N_22091,N_20615,N_20337);
and U22092 (N_22092,N_21105,N_21886);
xor U22093 (N_22093,N_20753,N_21157);
nand U22094 (N_22094,N_20316,N_21973);
or U22095 (N_22095,N_20179,N_21482);
and U22096 (N_22096,N_21405,N_21677);
nand U22097 (N_22097,N_21290,N_21450);
xor U22098 (N_22098,N_21718,N_20672);
nor U22099 (N_22099,N_21914,N_21484);
or U22100 (N_22100,N_20679,N_21316);
or U22101 (N_22101,N_21115,N_21796);
xnor U22102 (N_22102,N_21302,N_21390);
nand U22103 (N_22103,N_20270,N_21593);
or U22104 (N_22104,N_21064,N_20178);
nor U22105 (N_22105,N_21636,N_20026);
or U22106 (N_22106,N_21197,N_20376);
nand U22107 (N_22107,N_20675,N_21288);
nand U22108 (N_22108,N_21228,N_20515);
xnor U22109 (N_22109,N_21354,N_20021);
and U22110 (N_22110,N_20738,N_20276);
nor U22111 (N_22111,N_21911,N_20632);
nand U22112 (N_22112,N_21644,N_21214);
or U22113 (N_22113,N_20409,N_20775);
and U22114 (N_22114,N_20101,N_21083);
or U22115 (N_22115,N_21402,N_20461);
and U22116 (N_22116,N_20458,N_20765);
and U22117 (N_22117,N_21297,N_21568);
or U22118 (N_22118,N_21683,N_20031);
xor U22119 (N_22119,N_20361,N_20573);
or U22120 (N_22120,N_21252,N_21003);
and U22121 (N_22121,N_20304,N_21820);
and U22122 (N_22122,N_21749,N_20080);
nor U22123 (N_22123,N_20099,N_21684);
xnor U22124 (N_22124,N_21005,N_21359);
xor U22125 (N_22125,N_21036,N_21325);
xnor U22126 (N_22126,N_21910,N_20785);
nand U22127 (N_22127,N_20468,N_21078);
and U22128 (N_22128,N_21414,N_20692);
nand U22129 (N_22129,N_21351,N_20324);
xnor U22130 (N_22130,N_21873,N_20752);
nor U22131 (N_22131,N_21176,N_20302);
xnor U22132 (N_22132,N_21623,N_21700);
nor U22133 (N_22133,N_20008,N_20935);
nand U22134 (N_22134,N_21478,N_21500);
nand U22135 (N_22135,N_21842,N_21427);
nor U22136 (N_22136,N_21539,N_20273);
and U22137 (N_22137,N_21396,N_20780);
xor U22138 (N_22138,N_20519,N_21686);
and U22139 (N_22139,N_21985,N_21632);
or U22140 (N_22140,N_21616,N_21072);
or U22141 (N_22141,N_20091,N_21837);
xnor U22142 (N_22142,N_20564,N_20750);
or U22143 (N_22143,N_20487,N_20185);
nand U22144 (N_22144,N_20806,N_20603);
or U22145 (N_22145,N_20847,N_21338);
or U22146 (N_22146,N_20805,N_20132);
and U22147 (N_22147,N_21697,N_20259);
nand U22148 (N_22148,N_21890,N_21215);
nor U22149 (N_22149,N_20300,N_20015);
and U22150 (N_22150,N_20642,N_20397);
and U22151 (N_22151,N_21222,N_20443);
xor U22152 (N_22152,N_21497,N_20207);
xor U22153 (N_22153,N_20634,N_21146);
xnor U22154 (N_22154,N_21791,N_20501);
or U22155 (N_22155,N_21904,N_20315);
and U22156 (N_22156,N_20011,N_20526);
xor U22157 (N_22157,N_20719,N_20903);
and U22158 (N_22158,N_20505,N_20128);
or U22159 (N_22159,N_21273,N_21274);
or U22160 (N_22160,N_21765,N_20556);
or U22161 (N_22161,N_21650,N_20113);
nor U22162 (N_22162,N_20139,N_20647);
nor U22163 (N_22163,N_20966,N_21870);
xor U22164 (N_22164,N_20597,N_21094);
nor U22165 (N_22165,N_20715,N_20495);
nor U22166 (N_22166,N_21662,N_21174);
nand U22167 (N_22167,N_20538,N_21839);
xor U22168 (N_22168,N_20546,N_20133);
nor U22169 (N_22169,N_20580,N_21286);
nor U22170 (N_22170,N_21145,N_20670);
or U22171 (N_22171,N_21225,N_20525);
and U22172 (N_22172,N_21544,N_20943);
or U22173 (N_22173,N_20859,N_21902);
and U22174 (N_22174,N_20622,N_21832);
nand U22175 (N_22175,N_21126,N_21193);
nor U22176 (N_22176,N_20057,N_21192);
nor U22177 (N_22177,N_21950,N_21508);
nor U22178 (N_22178,N_20938,N_21709);
or U22179 (N_22179,N_21122,N_21320);
and U22180 (N_22180,N_20219,N_21975);
or U22181 (N_22181,N_20524,N_20238);
nand U22182 (N_22182,N_21242,N_20076);
nand U22183 (N_22183,N_20433,N_20203);
nor U22184 (N_22184,N_20319,N_21701);
nor U22185 (N_22185,N_20140,N_20548);
nand U22186 (N_22186,N_20370,N_21685);
and U22187 (N_22187,N_21531,N_20954);
nor U22188 (N_22188,N_20618,N_20994);
nor U22189 (N_22189,N_20230,N_21391);
and U22190 (N_22190,N_21514,N_21378);
and U22191 (N_22191,N_21457,N_21807);
and U22192 (N_22192,N_21437,N_21962);
nand U22193 (N_22193,N_21736,N_20012);
nor U22194 (N_22194,N_21368,N_21816);
and U22195 (N_22195,N_21693,N_21571);
nor U22196 (N_22196,N_20814,N_21303);
xor U22197 (N_22197,N_21407,N_21060);
xor U22198 (N_22198,N_20191,N_20770);
nand U22199 (N_22199,N_20795,N_21032);
and U22200 (N_22200,N_20767,N_20484);
or U22201 (N_22201,N_20595,N_21916);
xor U22202 (N_22202,N_21143,N_21294);
nand U22203 (N_22203,N_21594,N_20018);
nand U22204 (N_22204,N_20346,N_20507);
and U22205 (N_22205,N_21804,N_21045);
xnor U22206 (N_22206,N_20986,N_20957);
and U22207 (N_22207,N_20016,N_20669);
nand U22208 (N_22208,N_21862,N_21277);
nand U22209 (N_22209,N_21876,N_20408);
nor U22210 (N_22210,N_20084,N_20798);
and U22211 (N_22211,N_21570,N_21590);
or U22212 (N_22212,N_20286,N_21705);
or U22213 (N_22213,N_21267,N_20671);
xor U22214 (N_22214,N_21324,N_21559);
nor U22215 (N_22215,N_21847,N_20048);
or U22216 (N_22216,N_20266,N_20410);
nor U22217 (N_22217,N_21706,N_21449);
or U22218 (N_22218,N_21451,N_21442);
and U22219 (N_22219,N_21922,N_20350);
nor U22220 (N_22220,N_21076,N_20593);
and U22221 (N_22221,N_20629,N_21505);
and U22222 (N_22222,N_20656,N_20694);
xor U22223 (N_22223,N_20835,N_21166);
nand U22224 (N_22224,N_20292,N_21827);
and U22225 (N_22225,N_20224,N_21139);
nor U22226 (N_22226,N_21526,N_20586);
and U22227 (N_22227,N_20876,N_21538);
nor U22228 (N_22228,N_21443,N_20079);
or U22229 (N_22229,N_20697,N_21666);
or U22230 (N_22230,N_20293,N_20379);
nor U22231 (N_22231,N_20929,N_20437);
nand U22232 (N_22232,N_21738,N_21984);
nor U22233 (N_22233,N_20565,N_21560);
xor U22234 (N_22234,N_21178,N_21387);
or U22235 (N_22235,N_20274,N_20116);
xor U22236 (N_22236,N_20283,N_20477);
and U22237 (N_22237,N_21844,N_21168);
nor U22238 (N_22238,N_21855,N_21853);
or U22239 (N_22239,N_20757,N_21260);
and U22240 (N_22240,N_20450,N_21513);
nand U22241 (N_22241,N_21535,N_21349);
nor U22242 (N_22242,N_21806,N_21188);
nand U22243 (N_22243,N_20528,N_21780);
nand U22244 (N_22244,N_20038,N_21155);
or U22245 (N_22245,N_21187,N_21021);
nor U22246 (N_22246,N_21055,N_20861);
nand U22247 (N_22247,N_21369,N_20059);
and U22248 (N_22248,N_20150,N_21507);
nor U22249 (N_22249,N_20242,N_21580);
or U22250 (N_22250,N_20589,N_21793);
nor U22251 (N_22251,N_20343,N_20416);
nand U22252 (N_22252,N_20914,N_20068);
or U22253 (N_22253,N_20610,N_21050);
nor U22254 (N_22254,N_20871,N_20002);
xnor U22255 (N_22255,N_21458,N_20201);
nor U22256 (N_22256,N_21756,N_20313);
xnor U22257 (N_22257,N_20243,N_20115);
or U22258 (N_22258,N_20188,N_20160);
or U22259 (N_22259,N_21119,N_20990);
xnor U22260 (N_22260,N_21207,N_21781);
nor U22261 (N_22261,N_21722,N_20052);
or U22262 (N_22262,N_20513,N_20420);
xnor U22263 (N_22263,N_21172,N_21511);
and U22264 (N_22264,N_20184,N_21335);
nand U22265 (N_22265,N_21206,N_20648);
and U22266 (N_22266,N_20202,N_21248);
nand U22267 (N_22267,N_20383,N_20958);
nand U22268 (N_22268,N_21621,N_20268);
and U22269 (N_22269,N_20659,N_20844);
nor U22270 (N_22270,N_20599,N_20620);
and U22271 (N_22271,N_21762,N_21789);
or U22272 (N_22272,N_20457,N_21093);
nand U22273 (N_22273,N_21501,N_20024);
or U22274 (N_22274,N_21091,N_20754);
and U22275 (N_22275,N_20037,N_20989);
nor U22276 (N_22276,N_20186,N_20637);
and U22277 (N_22277,N_21994,N_20454);
nand U22278 (N_22278,N_20882,N_20034);
xnor U22279 (N_22279,N_20801,N_20340);
xor U22280 (N_22280,N_20924,N_21088);
and U22281 (N_22281,N_21269,N_21691);
nand U22282 (N_22282,N_20193,N_21480);
xor U22283 (N_22283,N_20272,N_21747);
xnor U22284 (N_22284,N_20036,N_21628);
xor U22285 (N_22285,N_21239,N_20345);
and U22286 (N_22286,N_21936,N_20479);
or U22287 (N_22287,N_21624,N_21026);
or U22288 (N_22288,N_21880,N_20658);
or U22289 (N_22289,N_21107,N_20159);
and U22290 (N_22290,N_20510,N_21417);
or U22291 (N_22291,N_21743,N_21609);
and U22292 (N_22292,N_20857,N_20728);
xnor U22293 (N_22293,N_21708,N_20893);
and U22294 (N_22294,N_20368,N_20288);
or U22295 (N_22295,N_20934,N_20331);
xnor U22296 (N_22296,N_20061,N_20907);
or U22297 (N_22297,N_21703,N_20349);
nand U22298 (N_22298,N_20743,N_21790);
nor U22299 (N_22299,N_21589,N_21334);
nand U22300 (N_22300,N_20469,N_21079);
or U22301 (N_22301,N_21220,N_20963);
or U22302 (N_22302,N_20295,N_20077);
and U22303 (N_22303,N_21398,N_20617);
or U22304 (N_22304,N_20182,N_21613);
or U22305 (N_22305,N_20774,N_21183);
xnor U22306 (N_22306,N_20755,N_21152);
nor U22307 (N_22307,N_20047,N_21424);
nor U22308 (N_22308,N_21929,N_21144);
and U22309 (N_22309,N_20396,N_21092);
xor U22310 (N_22310,N_20257,N_20145);
and U22311 (N_22311,N_21445,N_20987);
nor U22312 (N_22312,N_20950,N_20668);
xnor U22313 (N_22313,N_21657,N_21023);
xnor U22314 (N_22314,N_21135,N_20787);
and U22315 (N_22315,N_20192,N_21913);
and U22316 (N_22316,N_21615,N_20190);
and U22317 (N_22317,N_21834,N_21314);
nor U22318 (N_22318,N_20413,N_21217);
nor U22319 (N_22319,N_21127,N_20741);
nand U22320 (N_22320,N_20135,N_21476);
or U22321 (N_22321,N_21483,N_20621);
and U22322 (N_22322,N_21067,N_21553);
nor U22323 (N_22323,N_20791,N_21861);
xor U22324 (N_22324,N_21042,N_21561);
nand U22325 (N_22325,N_21141,N_20962);
and U22326 (N_22326,N_20335,N_21552);
nand U22327 (N_22327,N_20152,N_21953);
or U22328 (N_22328,N_20928,N_20699);
xnor U22329 (N_22329,N_21788,N_20594);
nand U22330 (N_22330,N_21081,N_21151);
or U22331 (N_22331,N_21825,N_21030);
or U22332 (N_22332,N_20210,N_20043);
nor U22333 (N_22333,N_21380,N_21748);
nand U22334 (N_22334,N_20241,N_20462);
and U22335 (N_22335,N_20583,N_20472);
nand U22336 (N_22336,N_20971,N_21692);
xor U22337 (N_22337,N_21957,N_20759);
and U22338 (N_22338,N_20710,N_21229);
nor U22339 (N_22339,N_21235,N_21035);
xnor U22340 (N_22340,N_21710,N_20246);
xnor U22341 (N_22341,N_21068,N_21651);
nand U22342 (N_22342,N_20054,N_20972);
and U22343 (N_22343,N_20590,N_20499);
or U22344 (N_22344,N_20863,N_21969);
xnor U22345 (N_22345,N_20554,N_20631);
and U22346 (N_22346,N_20153,N_20394);
and U22347 (N_22347,N_21100,N_20998);
nor U22348 (N_22348,N_21818,N_21573);
and U22349 (N_22349,N_21841,N_20262);
and U22350 (N_22350,N_20306,N_20912);
and U22351 (N_22351,N_21227,N_21935);
or U22352 (N_22352,N_21046,N_20213);
xor U22353 (N_22353,N_21585,N_21670);
and U22354 (N_22354,N_21728,N_20168);
and U22355 (N_22355,N_21699,N_21329);
and U22356 (N_22356,N_21150,N_20004);
nor U22357 (N_22357,N_21583,N_20339);
xnor U22358 (N_22358,N_20354,N_21365);
nand U22359 (N_22359,N_21564,N_21101);
xor U22360 (N_22360,N_20776,N_21943);
nor U22361 (N_22361,N_20260,N_21272);
or U22362 (N_22362,N_21874,N_21869);
or U22363 (N_22363,N_21646,N_20959);
nand U22364 (N_22364,N_20365,N_20901);
and U22365 (N_22365,N_20852,N_20271);
nand U22366 (N_22366,N_20406,N_21318);
nor U22367 (N_22367,N_21204,N_21720);
xnor U22368 (N_22368,N_20952,N_21941);
nor U22369 (N_22369,N_21012,N_21899);
or U22370 (N_22370,N_20236,N_21528);
or U22371 (N_22371,N_20181,N_20913);
and U22372 (N_22372,N_20742,N_21493);
nand U22373 (N_22373,N_20000,N_20904);
and U22374 (N_22374,N_21412,N_21388);
and U22375 (N_22375,N_21956,N_21872);
xor U22376 (N_22376,N_20716,N_20144);
or U22377 (N_22377,N_21459,N_21216);
or U22378 (N_22378,N_20700,N_21038);
xor U22379 (N_22379,N_20696,N_20464);
nand U22380 (N_22380,N_20837,N_20701);
or U22381 (N_22381,N_20541,N_21022);
and U22382 (N_22382,N_21305,N_20733);
or U22383 (N_22383,N_20431,N_21906);
and U22384 (N_22384,N_20172,N_20352);
or U22385 (N_22385,N_21271,N_21866);
xnor U22386 (N_22386,N_20177,N_20558);
nand U22387 (N_22387,N_20639,N_20652);
nand U22388 (N_22388,N_20112,N_20664);
nor U22389 (N_22389,N_21908,N_20045);
or U22390 (N_22390,N_21011,N_20840);
or U22391 (N_22391,N_21631,N_20623);
or U22392 (N_22392,N_20204,N_20627);
nand U22393 (N_22393,N_20404,N_21311);
nor U22394 (N_22394,N_20681,N_20455);
xnor U22395 (N_22395,N_20117,N_20398);
or U22396 (N_22396,N_21753,N_21537);
nor U22397 (N_22397,N_21852,N_20909);
xnor U22398 (N_22398,N_20975,N_21958);
or U22399 (N_22399,N_21939,N_20758);
nor U22400 (N_22400,N_21897,N_20299);
or U22401 (N_22401,N_20407,N_21291);
or U22402 (N_22402,N_20511,N_21017);
or U22403 (N_22403,N_20164,N_21724);
nor U22404 (N_22404,N_21612,N_21433);
or U22405 (N_22405,N_20856,N_21602);
nor U22406 (N_22406,N_20098,N_20984);
and U22407 (N_22407,N_20646,N_20014);
and U22408 (N_22408,N_21828,N_21606);
or U22409 (N_22409,N_20703,N_20685);
nor U22410 (N_22410,N_20786,N_21444);
nor U22411 (N_22411,N_20711,N_20850);
or U22412 (N_22412,N_20804,N_20736);
nand U22413 (N_22413,N_20439,N_20083);
or U22414 (N_22414,N_21470,N_20559);
or U22415 (N_22415,N_20211,N_20423);
nand U22416 (N_22416,N_20377,N_20312);
or U22417 (N_22417,N_21477,N_21170);
and U22418 (N_22418,N_20405,N_21915);
nor U22419 (N_22419,N_20289,N_21782);
or U22420 (N_22420,N_21704,N_20561);
and U22421 (N_22421,N_21475,N_20001);
and U22422 (N_22422,N_20320,N_20389);
nor U22423 (N_22423,N_21084,N_20417);
nor U22424 (N_22424,N_21610,N_21967);
nand U22425 (N_22425,N_20931,N_21439);
xor U22426 (N_22426,N_21040,N_21805);
or U22427 (N_22427,N_20500,N_20130);
and U22428 (N_22428,N_21498,N_20712);
and U22429 (N_22429,N_21757,N_21353);
and U22430 (N_22430,N_21472,N_21361);
or U22431 (N_22431,N_20284,N_20644);
nand U22432 (N_22432,N_21833,N_20682);
nand U22433 (N_22433,N_20930,N_21566);
or U22434 (N_22434,N_21070,N_21010);
nor U22435 (N_22435,N_21597,N_21004);
nor U22436 (N_22436,N_20866,N_21676);
and U22437 (N_22437,N_20605,N_21464);
or U22438 (N_22438,N_21669,N_20562);
nor U22439 (N_22439,N_21900,N_20430);
nand U22440 (N_22440,N_20749,N_20811);
and U22441 (N_22441,N_20571,N_20136);
nand U22442 (N_22442,N_20351,N_20149);
nand U22443 (N_22443,N_20082,N_20421);
nand U22444 (N_22444,N_21456,N_20297);
and U22445 (N_22445,N_20636,N_21859);
xor U22446 (N_22446,N_21491,N_20601);
or U22447 (N_22447,N_21099,N_20713);
nor U22448 (N_22448,N_20253,N_20778);
or U22449 (N_22449,N_21416,N_21803);
xnor U22450 (N_22450,N_20118,N_21376);
nand U22451 (N_22451,N_20926,N_21110);
nor U22452 (N_22452,N_21317,N_20764);
nand U22453 (N_22453,N_20799,N_20033);
nand U22454 (N_22454,N_21980,N_20974);
or U22455 (N_22455,N_20086,N_20566);
xnor U22456 (N_22456,N_21352,N_20060);
and U22457 (N_22457,N_20539,N_21158);
nor U22458 (N_22458,N_20820,N_20645);
or U22459 (N_22459,N_20208,N_21108);
nand U22460 (N_22460,N_21340,N_21428);
nand U22461 (N_22461,N_20362,N_21751);
xnor U22462 (N_22462,N_20854,N_20826);
xor U22463 (N_22463,N_20154,N_20602);
xor U22464 (N_22464,N_20517,N_21754);
and U22465 (N_22465,N_21732,N_20706);
nor U22466 (N_22466,N_20310,N_21132);
xnor U22467 (N_22467,N_21946,N_21678);
nor U22468 (N_22468,N_20829,N_21660);
nor U22469 (N_22469,N_20894,N_20378);
and U22470 (N_22470,N_20216,N_21851);
and U22471 (N_22471,N_21772,N_21626);
nand U22472 (N_22472,N_21292,N_21575);
or U22473 (N_22473,N_20322,N_20333);
xor U22474 (N_22474,N_20165,N_21041);
and U22475 (N_22475,N_21882,N_20684);
or U22476 (N_22476,N_21383,N_20482);
xor U22477 (N_22477,N_20807,N_21421);
or U22478 (N_22478,N_20418,N_20783);
and U22479 (N_22479,N_21256,N_21171);
xnor U22480 (N_22480,N_21393,N_20518);
nor U22481 (N_22481,N_21452,N_20747);
or U22482 (N_22482,N_20019,N_21205);
nand U22483 (N_22483,N_20991,N_21711);
or U22484 (N_22484,N_21044,N_20264);
or U22485 (N_22485,N_21307,N_21937);
and U22486 (N_22486,N_20874,N_21881);
xnor U22487 (N_22487,N_20078,N_20889);
and U22488 (N_22488,N_21965,N_21065);
xnor U22489 (N_22489,N_21607,N_20318);
and U22490 (N_22490,N_21438,N_21731);
nand U22491 (N_22491,N_20705,N_20973);
xnor U22492 (N_22492,N_20879,N_20608);
nand U22493 (N_22493,N_20784,N_20142);
nand U22494 (N_22494,N_21988,N_21879);
and U22495 (N_22495,N_21374,N_21154);
nor U22496 (N_22496,N_20453,N_21202);
and U22497 (N_22497,N_21576,N_21696);
or U22498 (N_22498,N_21582,N_20545);
or U22499 (N_22499,N_21053,N_20939);
xnor U22500 (N_22500,N_20222,N_20827);
nor U22501 (N_22501,N_21466,N_20819);
xnor U22502 (N_22502,N_20003,N_20411);
or U22503 (N_22503,N_20997,N_20332);
nor U22504 (N_22504,N_20143,N_21840);
nor U22505 (N_22505,N_21846,N_21194);
xor U22506 (N_22506,N_20745,N_20496);
or U22507 (N_22507,N_20356,N_20237);
or U22508 (N_22508,N_20611,N_20643);
nand U22509 (N_22509,N_20977,N_21547);
and U22510 (N_22510,N_21136,N_21453);
or U22511 (N_22511,N_21690,N_21448);
xnor U22512 (N_22512,N_21759,N_20570);
and U22513 (N_22513,N_21114,N_20531);
nor U22514 (N_22514,N_21715,N_21619);
xnor U22515 (N_22515,N_21730,N_21614);
or U22516 (N_22516,N_20414,N_21411);
or U22517 (N_22517,N_20232,N_21871);
and U22518 (N_22518,N_21865,N_20739);
nor U22519 (N_22519,N_21190,N_20792);
nor U22520 (N_22520,N_21891,N_21625);
nor U22521 (N_22521,N_20158,N_20072);
nand U22522 (N_22522,N_21095,N_20088);
and U22523 (N_22523,N_20591,N_21386);
and U22524 (N_22524,N_20471,N_21549);
and U22525 (N_22525,N_21663,N_20872);
and U22526 (N_22526,N_21679,N_20920);
xor U22527 (N_22527,N_20584,N_21479);
or U22528 (N_22528,N_21605,N_21315);
or U22529 (N_22529,N_20478,N_21826);
and U22530 (N_22530,N_20945,N_21364);
and U22531 (N_22531,N_21322,N_20393);
nor U22532 (N_22532,N_20228,N_21086);
nor U22533 (N_22533,N_21801,N_20746);
nor U22534 (N_22534,N_20869,N_20265);
nand U22535 (N_22535,N_21336,N_20050);
nand U22536 (N_22536,N_20360,N_21087);
nand U22537 (N_22537,N_20155,N_20822);
nand U22538 (N_22538,N_20125,N_20183);
and U22539 (N_22539,N_20231,N_21821);
nor U22540 (N_22540,N_20380,N_21800);
nor U22541 (N_22541,N_20301,N_21581);
or U22542 (N_22542,N_20727,N_20189);
nor U22543 (N_22543,N_21763,N_20442);
and U22544 (N_22544,N_20751,N_20263);
or U22545 (N_22545,N_21661,N_20095);
nand U22546 (N_22546,N_21454,N_20686);
nor U22547 (N_22547,N_21742,N_20247);
nor U22548 (N_22548,N_20044,N_21664);
or U22549 (N_22549,N_21682,N_21280);
nor U22550 (N_22550,N_20862,N_21752);
xnor U22551 (N_22551,N_20395,N_21221);
xor U22552 (N_22552,N_21051,N_21447);
xor U22553 (N_22553,N_21733,N_21066);
nand U22554 (N_22554,N_20768,N_21572);
and U22555 (N_22555,N_21330,N_20782);
and U22556 (N_22556,N_20111,N_20726);
nor U22557 (N_22557,N_21343,N_21485);
and U22558 (N_22558,N_20880,N_21656);
xor U22559 (N_22559,N_21062,N_20109);
nor U22560 (N_22560,N_20900,N_21481);
xor U22561 (N_22561,N_20373,N_20689);
nand U22562 (N_22562,N_20512,N_21779);
and U22563 (N_22563,N_21434,N_21928);
xor U22564 (N_22564,N_21721,N_21109);
nand U22565 (N_22565,N_20592,N_21918);
xor U22566 (N_22566,N_20460,N_21838);
or U22567 (N_22567,N_21494,N_20173);
nor U22568 (N_22568,N_21140,N_20717);
and U22569 (N_22569,N_21617,N_21512);
or U22570 (N_22570,N_20956,N_21681);
xnor U22571 (N_22571,N_21313,N_20883);
nand U22572 (N_22572,N_21964,N_21356);
or U22573 (N_22573,N_21640,N_21131);
nand U22574 (N_22574,N_20290,N_20877);
xor U22575 (N_22575,N_21236,N_21319);
and U22576 (N_22576,N_20803,N_21787);
nor U22577 (N_22577,N_20023,N_21554);
or U22578 (N_22578,N_21382,N_20577);
nand U22579 (N_22579,N_21758,N_20587);
and U22580 (N_22580,N_21394,N_21262);
or U22581 (N_22581,N_20129,N_21887);
nor U22582 (N_22582,N_21420,N_20279);
nor U22583 (N_22583,N_20074,N_20248);
and U22584 (N_22584,N_20674,N_21652);
xor U22585 (N_22585,N_21653,N_20946);
xor U22586 (N_22586,N_21925,N_20364);
nand U22587 (N_22587,N_20549,N_21995);
xor U22588 (N_22588,N_21342,N_20467);
or U22589 (N_22589,N_20156,N_20868);
and U22590 (N_22590,N_20895,N_21885);
nor U22591 (N_22591,N_21253,N_20428);
and U22592 (N_22592,N_20267,N_21463);
and U22593 (N_22593,N_21815,N_21510);
nand U22594 (N_22594,N_21927,N_20506);
nor U22595 (N_22595,N_20285,N_21199);
or U22596 (N_22596,N_21830,N_20317);
or U22597 (N_22597,N_20983,N_20017);
or U22598 (N_22598,N_21399,N_20280);
nor U22599 (N_22599,N_20049,N_21153);
nor U22600 (N_22600,N_21817,N_20081);
nor U22601 (N_22601,N_20563,N_21137);
or U22602 (N_22602,N_20056,N_21924);
and U22603 (N_22603,N_20353,N_20769);
nor U22604 (N_22604,N_20992,N_21245);
nand U22605 (N_22605,N_21592,N_21982);
nor U22606 (N_22606,N_21959,N_20215);
and U22607 (N_22607,N_21019,N_21998);
and U22608 (N_22608,N_20906,N_21808);
and U22609 (N_22609,N_20448,N_20823);
xnor U22610 (N_22610,N_20384,N_20897);
nor U22611 (N_22611,N_20240,N_20955);
nor U22612 (N_22612,N_21854,N_20732);
nor U22613 (N_22613,N_21785,N_21823);
or U22614 (N_22614,N_20709,N_20555);
nand U22615 (N_22615,N_21121,N_21987);
or U22616 (N_22616,N_20771,N_20551);
or U22617 (N_22617,N_20960,N_21795);
nand U22618 (N_22618,N_21275,N_21002);
nand U22619 (N_22619,N_21243,N_20881);
nor U22620 (N_22620,N_20206,N_21599);
or U22621 (N_22621,N_20386,N_20520);
nor U22622 (N_22622,N_20221,N_20226);
and U22623 (N_22623,N_20249,N_20527);
or U22624 (N_22624,N_21047,N_21917);
nand U22625 (N_22625,N_21028,N_20662);
nor U22626 (N_22626,N_21545,N_21360);
or U22627 (N_22627,N_20834,N_21892);
nand U22628 (N_22628,N_20124,N_20575);
and U22629 (N_22629,N_20579,N_21249);
xor U22630 (N_22630,N_21586,N_21931);
and U22631 (N_22631,N_20680,N_21542);
or U22632 (N_22632,N_21819,N_21523);
or U22633 (N_22633,N_21637,N_21440);
nor U22634 (N_22634,N_21460,N_20970);
and U22635 (N_22635,N_20382,N_21836);
nor U22636 (N_22636,N_21113,N_21655);
nand U22637 (N_22637,N_21608,N_21798);
xor U22638 (N_22638,N_20492,N_21082);
or U22639 (N_22639,N_21877,N_20277);
or U22640 (N_22640,N_21344,N_21289);
xnor U22641 (N_22641,N_20842,N_20529);
xor U22642 (N_22642,N_20217,N_21133);
nor U22643 (N_22643,N_21555,N_20588);
and U22644 (N_22644,N_21054,N_20884);
nor U22645 (N_22645,N_21521,N_21996);
nand U22646 (N_22646,N_20122,N_21735);
or U22647 (N_22647,N_20638,N_20677);
or U22648 (N_22648,N_21173,N_20020);
nor U22649 (N_22649,N_20441,N_20723);
or U22650 (N_22650,N_20773,N_21016);
nor U22651 (N_22651,N_21716,N_20695);
and U22652 (N_22652,N_21919,N_20258);
and U22653 (N_22653,N_21695,N_21849);
xnor U22654 (N_22654,N_21213,N_20982);
nand U22655 (N_22655,N_20761,N_20649);
nor U22656 (N_22656,N_20447,N_21971);
xor U22657 (N_22657,N_20102,N_20781);
nor U22658 (N_22658,N_21486,N_20878);
nand U22659 (N_22659,N_21212,N_21461);
or U22660 (N_22660,N_21309,N_21301);
nor U22661 (N_22661,N_20812,N_20106);
nor U22662 (N_22662,N_20665,N_21940);
and U22663 (N_22663,N_20281,N_21604);
or U22664 (N_22664,N_21226,N_20309);
nor U22665 (N_22665,N_20902,N_21200);
xnor U22666 (N_22666,N_21401,N_20606);
xor U22667 (N_22667,N_21413,N_21533);
nor U22668 (N_22668,N_21223,N_20167);
nor U22669 (N_22669,N_21431,N_20087);
and U22670 (N_22670,N_21642,N_20327);
nor U22671 (N_22671,N_21680,N_20085);
and U22672 (N_22672,N_20948,N_21014);
nor U22673 (N_22673,N_21257,N_20925);
nor U22674 (N_22674,N_20490,N_21075);
nor U22675 (N_22675,N_21425,N_21955);
xor U22676 (N_22676,N_20890,N_21770);
or U22677 (N_22677,N_21896,N_21551);
nor U22678 (N_22678,N_21786,N_20763);
nor U22679 (N_22679,N_21208,N_20831);
nor U22680 (N_22680,N_20220,N_21649);
xnor U22681 (N_22681,N_20800,N_20198);
and U22682 (N_22682,N_21156,N_20899);
xor U22683 (N_22683,N_20860,N_21857);
nand U22684 (N_22684,N_21951,N_20040);
or U22685 (N_22685,N_20391,N_21487);
and U22686 (N_22686,N_21346,N_21112);
nand U22687 (N_22687,N_20988,N_21949);
and U22688 (N_22688,N_20141,N_21641);
nor U22689 (N_22689,N_21426,N_21522);
or U22690 (N_22690,N_20802,N_20022);
nor U22691 (N_22691,N_20504,N_21266);
nand U22692 (N_22692,N_20516,N_20488);
or U22693 (N_22693,N_20100,N_21337);
xor U22694 (N_22694,N_20867,N_20522);
xor U22695 (N_22695,N_21667,N_21702);
or U22696 (N_22696,N_21822,N_20790);
xor U22697 (N_22697,N_20205,N_21001);
nor U22698 (N_22698,N_20550,N_21645);
xnor U22699 (N_22699,N_21905,N_21263);
xnor U22700 (N_22700,N_21546,N_20923);
and U22701 (N_22701,N_20287,N_20891);
xnor U22702 (N_22702,N_21578,N_20568);
or U22703 (N_22703,N_20916,N_20440);
xnor U22704 (N_22704,N_21160,N_21529);
xnor U22705 (N_22705,N_20196,N_21744);
nor U22706 (N_22706,N_20721,N_20793);
xnor U22707 (N_22707,N_20737,N_20218);
and U22708 (N_22708,N_20654,N_20839);
or U22709 (N_22709,N_20436,N_21348);
nand U22710 (N_22710,N_21247,N_20444);
and U22711 (N_22711,N_20334,N_20810);
xor U22712 (N_22712,N_21889,N_21750);
and U22713 (N_22713,N_21860,N_21134);
and U22714 (N_22714,N_21232,N_20731);
nand U22715 (N_22715,N_20338,N_20200);
and U22716 (N_22716,N_21775,N_20169);
and U22717 (N_22717,N_20483,N_20915);
and U22718 (N_22718,N_21015,N_21888);
xnor U22719 (N_22719,N_20567,N_20707);
xor U22720 (N_22720,N_21224,N_20427);
or U22721 (N_22721,N_21638,N_21404);
xnor U22722 (N_22722,N_21167,N_20127);
and U22723 (N_22723,N_20375,N_21893);
and U22724 (N_22724,N_20969,N_20569);
nor U22725 (N_22725,N_20278,N_21455);
nor U22726 (N_22726,N_20626,N_20005);
nor U22727 (N_22727,N_20459,N_20582);
xor U22728 (N_22728,N_20291,N_21333);
and U22729 (N_22729,N_20937,N_20614);
and U22730 (N_22730,N_20470,N_21310);
nor U22731 (N_22731,N_21270,N_20062);
nand U22732 (N_22732,N_21499,N_21218);
and U22733 (N_22733,N_21321,N_20096);
nand U22734 (N_22734,N_20808,N_20108);
nand U22735 (N_22735,N_20619,N_21327);
xnor U22736 (N_22736,N_21671,N_21233);
xor U22737 (N_22737,N_21323,N_20708);
and U22738 (N_22738,N_20336,N_21952);
nand U22739 (N_22739,N_21488,N_21773);
or U22740 (N_22740,N_21326,N_21116);
and U22741 (N_22741,N_21097,N_21367);
and U22742 (N_22742,N_20298,N_20256);
nand U22743 (N_22743,N_21794,N_20838);
and U22744 (N_22744,N_20097,N_21698);
or U22745 (N_22745,N_20922,N_21848);
nor U22746 (N_22746,N_21983,N_21831);
nand U22747 (N_22747,N_21255,N_20543);
nand U22748 (N_22748,N_21258,N_20294);
or U22749 (N_22749,N_21377,N_21182);
or U22750 (N_22750,N_21933,N_21633);
nand U22751 (N_22751,N_21587,N_20239);
and U22752 (N_22752,N_20624,N_20537);
nand U22753 (N_22753,N_21400,N_20995);
nand U22754 (N_22754,N_21355,N_21196);
and U22755 (N_22755,N_21811,N_21373);
and U22756 (N_22756,N_21435,N_20967);
xnor U22757 (N_22757,N_21259,N_20908);
nor U22758 (N_22758,N_21635,N_20508);
and U22759 (N_22759,N_21284,N_20552);
nand U22760 (N_22760,N_20704,N_20993);
nor U22761 (N_22761,N_20481,N_20176);
nand U22762 (N_22762,N_20229,N_21179);
xnor U22763 (N_22763,N_21209,N_21979);
nand U22764 (N_22764,N_20628,N_21462);
or U22765 (N_22765,N_21843,N_21520);
xnor U22766 (N_22766,N_20843,N_21375);
nand U22767 (N_22767,N_20476,N_21492);
or U22768 (N_22768,N_21241,N_20419);
nand U22769 (N_22769,N_20039,N_20722);
and U22770 (N_22770,N_21999,N_20463);
nand U22771 (N_22771,N_21250,N_21923);
xor U22772 (N_22772,N_20604,N_21970);
and U22773 (N_22773,N_21465,N_21165);
nor U22774 (N_22774,N_21536,N_20809);
nor U22775 (N_22775,N_20058,N_20720);
nand U22776 (N_22776,N_21175,N_20114);
nand U22777 (N_22777,N_21496,N_21659);
nand U22778 (N_22778,N_21673,N_21469);
nor U22779 (N_22779,N_20234,N_21506);
nand U22780 (N_22780,N_21977,N_20046);
and U22781 (N_22781,N_21418,N_20323);
nor U22782 (N_22782,N_20401,N_20572);
or U22783 (N_22783,N_21089,N_21944);
nand U22784 (N_22784,N_21997,N_20762);
xor U22785 (N_22785,N_21059,N_20366);
nand U22786 (N_22786,N_20363,N_21963);
xnor U22787 (N_22787,N_20166,N_21557);
nand U22788 (N_22788,N_21978,N_20424);
nor U22789 (N_22789,N_21524,N_21300);
or U22790 (N_22790,N_20534,N_20927);
or U22791 (N_22791,N_21611,N_21563);
or U22792 (N_22792,N_20104,N_20740);
xnor U22793 (N_22793,N_21909,N_21446);
nor U22794 (N_22794,N_20010,N_20683);
nor U22795 (N_22795,N_21298,N_21921);
or U22796 (N_22796,N_21540,N_21517);
or U22797 (N_22797,N_20557,N_20702);
or U22798 (N_22798,N_21195,N_21577);
and U22799 (N_22799,N_20326,N_21863);
or U22800 (N_22800,N_21737,N_21992);
nor U22801 (N_22801,N_20875,N_21177);
and U22802 (N_22802,N_20888,N_21783);
and U22803 (N_22803,N_21467,N_20607);
nand U22804 (N_22804,N_21968,N_20348);
nand U22805 (N_22805,N_21934,N_21503);
nor U22806 (N_22806,N_20953,N_20092);
nor U22807 (N_22807,N_20932,N_20374);
and U22808 (N_22808,N_21976,N_20497);
or U22809 (N_22809,N_20532,N_20905);
or U22810 (N_22810,N_21755,N_21104);
nor U22811 (N_22811,N_21687,N_20779);
or U22812 (N_22812,N_21717,N_20399);
xor U22813 (N_22813,N_20667,N_20641);
nand U22814 (N_22814,N_20030,N_20825);
nor U22815 (N_22815,N_21490,N_20828);
nand U22816 (N_22816,N_21658,N_21098);
xor U22817 (N_22817,N_21620,N_20162);
or U22818 (N_22818,N_21766,N_21991);
nand U22819 (N_22819,N_20025,N_20698);
xnor U22820 (N_22820,N_21363,N_20146);
and U22821 (N_22821,N_20687,N_20560);
xor U22822 (N_22822,N_20498,N_21007);
xor U22823 (N_22823,N_21518,N_21792);
nand U22824 (N_22824,N_21071,N_20853);
nor U22825 (N_22825,N_20429,N_20251);
xnor U22826 (N_22826,N_21634,N_21761);
nor U22827 (N_22827,N_20949,N_21381);
nor U22828 (N_22828,N_20609,N_21295);
nand U22829 (N_22829,N_20848,N_21474);
nand U22830 (N_22830,N_21884,N_20426);
or U22831 (N_22831,N_21111,N_20544);
xor U22832 (N_22832,N_21813,N_21713);
xor U22833 (N_22833,N_20212,N_20744);
or U22834 (N_22834,N_21648,N_21707);
nor U22835 (N_22835,N_21049,N_21000);
or U22836 (N_22836,N_21058,N_21090);
nand U22837 (N_22837,N_21674,N_21814);
nor U22838 (N_22838,N_20235,N_21647);
nor U22839 (N_22839,N_20653,N_21056);
and U22840 (N_22840,N_21123,N_20650);
nand U22841 (N_22841,N_20789,N_20197);
nand U22842 (N_22842,N_21912,N_21198);
nor U22843 (N_22843,N_20845,N_21595);
nor U22844 (N_22844,N_20964,N_20777);
nand U22845 (N_22845,N_21809,N_20357);
and U22846 (N_22846,N_20214,N_21689);
xnor U22847 (N_22847,N_20941,N_21031);
nor U22848 (N_22848,N_21120,N_20432);
and U22849 (N_22849,N_21601,N_21812);
and U22850 (N_22850,N_20676,N_21283);
nand U22851 (N_22851,N_21723,N_21509);
nand U22852 (N_22852,N_21358,N_20981);
or U22853 (N_22853,N_20325,N_20473);
nand U22854 (N_22854,N_20947,N_20307);
nor U22855 (N_22855,N_20598,N_21543);
or U22856 (N_22856,N_21385,N_21180);
nand U22857 (N_22857,N_20690,N_20425);
nand U22858 (N_22858,N_21989,N_21745);
nand U22859 (N_22859,N_20910,N_20388);
and U22860 (N_22860,N_21020,N_21858);
nor U22861 (N_22861,N_20223,N_20858);
nand U22862 (N_22862,N_21268,N_20613);
nor U22863 (N_22863,N_20390,N_20103);
nand U22864 (N_22864,N_21117,N_20412);
and U22865 (N_22865,N_21037,N_20244);
nor U22866 (N_22866,N_20985,N_20635);
nand U22867 (N_22867,N_21409,N_21328);
xor U22868 (N_22868,N_21415,N_20760);
xor U22869 (N_22869,N_21867,N_20663);
xor U22870 (N_22870,N_21006,N_21148);
and U22871 (N_22871,N_20075,N_21532);
or U22872 (N_22872,N_21668,N_21186);
nor U22873 (N_22873,N_21163,N_21341);
xor U22874 (N_22874,N_20225,N_21379);
nor U22875 (N_22875,N_20961,N_20381);
nand U22876 (N_22876,N_20308,N_21073);
nor U22877 (N_22877,N_21231,N_20480);
or U22878 (N_22878,N_21033,N_21966);
xor U22879 (N_22879,N_21281,N_21201);
xnor U22880 (N_22880,N_21688,N_20032);
nand U22881 (N_22881,N_21591,N_21556);
and U22882 (N_22882,N_21603,N_20514);
or U22883 (N_22883,N_21567,N_20475);
xnor U22884 (N_22884,N_21251,N_20296);
and U22885 (N_22885,N_20734,N_20965);
nor U22886 (N_22886,N_20509,N_21278);
nor U22887 (N_22887,N_20330,N_20836);
nor U22888 (N_22888,N_21986,N_21835);
nor U22889 (N_22889,N_20585,N_20815);
or U22890 (N_22890,N_20846,N_21574);
and U22891 (N_22891,N_21039,N_20657);
and U22892 (N_22892,N_21027,N_20435);
nand U22893 (N_22893,N_21345,N_20493);
nor U22894 (N_22894,N_21189,N_20035);
xor U22895 (N_22895,N_20233,N_21138);
and U22896 (N_22896,N_20918,N_21129);
xor U22897 (N_22897,N_20864,N_20887);
xnor U22898 (N_22898,N_21824,N_21403);
nor U22899 (N_22899,N_20797,N_20402);
xnor U22900 (N_22900,N_21726,N_20533);
nor U22901 (N_22901,N_21034,N_21395);
xor U22902 (N_22902,N_20885,N_20833);
and U22903 (N_22903,N_20093,N_21776);
xor U22904 (N_22904,N_21938,N_21920);
nand U22905 (N_22905,N_21883,N_20486);
nor U22906 (N_22906,N_20451,N_21410);
and U22907 (N_22907,N_21422,N_20385);
nor U22908 (N_22908,N_21299,N_20070);
xnor U22909 (N_22909,N_21622,N_20107);
and U22910 (N_22910,N_21898,N_21169);
or U22911 (N_22911,N_21519,N_21408);
nand U22912 (N_22912,N_20502,N_21429);
xnor U22913 (N_22913,N_21942,N_21159);
and U22914 (N_22914,N_20067,N_21392);
xnor U22915 (N_22915,N_21527,N_20976);
nand U22916 (N_22916,N_21350,N_21024);
nor U22917 (N_22917,N_20372,N_21471);
nor U22918 (N_22918,N_20921,N_20187);
nand U22919 (N_22919,N_20170,N_21282);
nand U22920 (N_22920,N_21675,N_21548);
and U22921 (N_22921,N_21525,N_20841);
and U22922 (N_22922,N_21774,N_20978);
and U22923 (N_22923,N_21954,N_21254);
and U22924 (N_22924,N_20161,N_21052);
and U22925 (N_22925,N_21901,N_21972);
or U22926 (N_22926,N_21102,N_20536);
or U22927 (N_22927,N_21868,N_21562);
nor U22928 (N_22928,N_21596,N_21981);
xnor U22929 (N_22929,N_20282,N_21430);
xnor U22930 (N_22930,N_20491,N_20053);
nor U22931 (N_22931,N_21219,N_20329);
and U22932 (N_22932,N_21432,N_20979);
or U22933 (N_22933,N_21308,N_21057);
or U22934 (N_22934,N_20227,N_20387);
xnor U22935 (N_22935,N_21362,N_20209);
nand U22936 (N_22936,N_20999,N_21128);
and U22937 (N_22937,N_21118,N_21096);
and U22938 (N_22938,N_20009,N_21639);
xor U22939 (N_22939,N_21727,N_20673);
nand U22940 (N_22940,N_20660,N_20119);
nand U22941 (N_22941,N_20456,N_20936);
nor U22942 (N_22942,N_20275,N_20171);
and U22943 (N_22943,N_20027,N_20542);
xor U22944 (N_22944,N_20028,N_21025);
and U22945 (N_22945,N_20980,N_21357);
nand U22946 (N_22946,N_20651,N_20194);
nand U22947 (N_22947,N_20131,N_20065);
or U22948 (N_22948,N_20796,N_20951);
xor U22949 (N_22949,N_20898,N_21164);
nor U22950 (N_22950,N_21764,N_20616);
xor U22951 (N_22951,N_20422,N_20465);
nor U22952 (N_22952,N_21161,N_20748);
and U22953 (N_22953,N_21974,N_20180);
and U22954 (N_22954,N_21043,N_20446);
and U22955 (N_22955,N_20415,N_20175);
nor U22956 (N_22956,N_21230,N_20121);
nor U22957 (N_22957,N_21948,N_21181);
and U22958 (N_22958,N_21339,N_21468);
nor U22959 (N_22959,N_21063,N_21856);
nor U22960 (N_22960,N_20530,N_21541);
nor U22961 (N_22961,N_20718,N_20174);
nand U22962 (N_22962,N_21504,N_21778);
and U22963 (N_22963,N_20576,N_21331);
or U22964 (N_22964,N_20073,N_20245);
or U22965 (N_22965,N_21237,N_20434);
nor U22966 (N_22966,N_21734,N_21234);
xor U22967 (N_22967,N_21932,N_20714);
xnor U22968 (N_22968,N_21502,N_20630);
and U22969 (N_22969,N_21665,N_20392);
nand U22970 (N_22970,N_20151,N_20788);
or U22971 (N_22971,N_20007,N_20355);
or U22972 (N_22972,N_20724,N_21515);
and U22973 (N_22973,N_20134,N_21878);
xnor U22974 (N_22974,N_21875,N_21264);
xnor U22975 (N_22975,N_20089,N_21285);
and U22976 (N_22976,N_21714,N_20449);
xnor U22977 (N_22977,N_20688,N_21279);
nand U22978 (N_22978,N_21077,N_21760);
xor U22979 (N_22979,N_21265,N_20063);
nor U22980 (N_22980,N_21534,N_20071);
nand U22981 (N_22981,N_20341,N_20255);
nor U22982 (N_22982,N_21845,N_20873);
nand U22983 (N_22983,N_20794,N_21142);
or U22984 (N_22984,N_21069,N_21769);
or U22985 (N_22985,N_20269,N_21618);
nor U22986 (N_22986,N_20996,N_20051);
and U22987 (N_22987,N_20359,N_20438);
nand U22988 (N_22988,N_21850,N_20494);
nor U22989 (N_22989,N_20371,N_20553);
xor U22990 (N_22990,N_21550,N_21211);
nor U22991 (N_22991,N_21162,N_21643);
and U22992 (N_22992,N_20919,N_20006);
nor U22993 (N_22993,N_20347,N_21739);
nand U22994 (N_22994,N_20199,N_21864);
or U22995 (N_22995,N_20314,N_21654);
nand U22996 (N_22996,N_20069,N_21629);
xor U22997 (N_22997,N_20148,N_21184);
xor U22998 (N_22998,N_20540,N_20640);
nor U22999 (N_22999,N_20110,N_20849);
and U23000 (N_23000,N_21456,N_21908);
and U23001 (N_23001,N_21006,N_20380);
xor U23002 (N_23002,N_20031,N_20193);
nand U23003 (N_23003,N_20716,N_20183);
and U23004 (N_23004,N_20414,N_20867);
or U23005 (N_23005,N_20421,N_21465);
and U23006 (N_23006,N_21158,N_20770);
and U23007 (N_23007,N_20164,N_21088);
xnor U23008 (N_23008,N_20776,N_21765);
xor U23009 (N_23009,N_20133,N_20549);
and U23010 (N_23010,N_21292,N_20266);
and U23011 (N_23011,N_20170,N_20144);
nor U23012 (N_23012,N_20550,N_21596);
and U23013 (N_23013,N_21448,N_21573);
nand U23014 (N_23014,N_20238,N_20426);
xor U23015 (N_23015,N_20936,N_20874);
and U23016 (N_23016,N_21717,N_21454);
xnor U23017 (N_23017,N_20550,N_20809);
nor U23018 (N_23018,N_21759,N_20628);
or U23019 (N_23019,N_21512,N_20970);
xnor U23020 (N_23020,N_20137,N_21117);
nor U23021 (N_23021,N_20237,N_21382);
nand U23022 (N_23022,N_21391,N_21734);
or U23023 (N_23023,N_21412,N_20172);
xor U23024 (N_23024,N_20107,N_21320);
xor U23025 (N_23025,N_21274,N_21535);
nand U23026 (N_23026,N_21016,N_20002);
nor U23027 (N_23027,N_21189,N_20431);
and U23028 (N_23028,N_21808,N_21641);
or U23029 (N_23029,N_21136,N_21095);
xnor U23030 (N_23030,N_20593,N_21558);
nor U23031 (N_23031,N_21347,N_20867);
and U23032 (N_23032,N_21402,N_21092);
or U23033 (N_23033,N_20801,N_21688);
and U23034 (N_23034,N_21565,N_20082);
nand U23035 (N_23035,N_21733,N_21875);
and U23036 (N_23036,N_20629,N_20085);
nor U23037 (N_23037,N_21299,N_21355);
xor U23038 (N_23038,N_20107,N_20217);
nor U23039 (N_23039,N_20396,N_21730);
xnor U23040 (N_23040,N_20475,N_21410);
nand U23041 (N_23041,N_20951,N_20946);
and U23042 (N_23042,N_21345,N_20237);
xnor U23043 (N_23043,N_21405,N_21883);
nor U23044 (N_23044,N_20923,N_20727);
nor U23045 (N_23045,N_21835,N_20638);
nand U23046 (N_23046,N_21631,N_21468);
xnor U23047 (N_23047,N_21152,N_21690);
or U23048 (N_23048,N_20463,N_21059);
or U23049 (N_23049,N_21977,N_21766);
and U23050 (N_23050,N_21928,N_20774);
nor U23051 (N_23051,N_20054,N_20796);
xor U23052 (N_23052,N_20846,N_21492);
or U23053 (N_23053,N_21036,N_20838);
or U23054 (N_23054,N_20393,N_20151);
nor U23055 (N_23055,N_21705,N_21025);
and U23056 (N_23056,N_20382,N_20194);
and U23057 (N_23057,N_20007,N_21032);
and U23058 (N_23058,N_20548,N_20724);
and U23059 (N_23059,N_21839,N_21756);
or U23060 (N_23060,N_21557,N_21898);
nand U23061 (N_23061,N_21469,N_21448);
or U23062 (N_23062,N_20049,N_20128);
or U23063 (N_23063,N_21368,N_20208);
xor U23064 (N_23064,N_21221,N_21805);
xnor U23065 (N_23065,N_20740,N_21489);
nor U23066 (N_23066,N_21347,N_21855);
or U23067 (N_23067,N_21310,N_21032);
xnor U23068 (N_23068,N_20630,N_20107);
nor U23069 (N_23069,N_21815,N_20565);
xnor U23070 (N_23070,N_20705,N_21688);
nand U23071 (N_23071,N_20623,N_20472);
nand U23072 (N_23072,N_20182,N_20636);
nor U23073 (N_23073,N_21671,N_20362);
or U23074 (N_23074,N_21873,N_20384);
or U23075 (N_23075,N_20696,N_20327);
nand U23076 (N_23076,N_21609,N_21042);
or U23077 (N_23077,N_20793,N_21772);
xor U23078 (N_23078,N_20838,N_21385);
nand U23079 (N_23079,N_20808,N_20493);
and U23080 (N_23080,N_20038,N_21846);
nand U23081 (N_23081,N_21899,N_20222);
and U23082 (N_23082,N_21048,N_21825);
xnor U23083 (N_23083,N_21171,N_21893);
nand U23084 (N_23084,N_20740,N_21548);
nor U23085 (N_23085,N_20191,N_21433);
xor U23086 (N_23086,N_20411,N_20378);
nor U23087 (N_23087,N_21613,N_21339);
xnor U23088 (N_23088,N_20225,N_21783);
xnor U23089 (N_23089,N_20892,N_20807);
xnor U23090 (N_23090,N_20335,N_20404);
or U23091 (N_23091,N_20192,N_21394);
nor U23092 (N_23092,N_21644,N_20636);
or U23093 (N_23093,N_21754,N_21575);
nand U23094 (N_23094,N_21412,N_21421);
and U23095 (N_23095,N_20891,N_20911);
nor U23096 (N_23096,N_21646,N_20811);
nand U23097 (N_23097,N_21983,N_21607);
nand U23098 (N_23098,N_20192,N_20980);
nand U23099 (N_23099,N_21714,N_20244);
and U23100 (N_23100,N_21267,N_20755);
xnor U23101 (N_23101,N_21511,N_20082);
nand U23102 (N_23102,N_20942,N_20549);
or U23103 (N_23103,N_21343,N_20556);
nand U23104 (N_23104,N_21024,N_20596);
nand U23105 (N_23105,N_21807,N_20961);
nor U23106 (N_23106,N_21242,N_20769);
xnor U23107 (N_23107,N_21292,N_20052);
nand U23108 (N_23108,N_21832,N_21401);
or U23109 (N_23109,N_21905,N_21508);
and U23110 (N_23110,N_20823,N_20122);
nand U23111 (N_23111,N_20868,N_20317);
or U23112 (N_23112,N_20040,N_21137);
nor U23113 (N_23113,N_20336,N_21162);
or U23114 (N_23114,N_20999,N_21516);
or U23115 (N_23115,N_21761,N_21333);
nand U23116 (N_23116,N_21937,N_21490);
nor U23117 (N_23117,N_21539,N_21647);
xnor U23118 (N_23118,N_20215,N_21411);
xor U23119 (N_23119,N_20443,N_21367);
nor U23120 (N_23120,N_21202,N_21534);
or U23121 (N_23121,N_20738,N_20179);
and U23122 (N_23122,N_20237,N_21714);
nor U23123 (N_23123,N_21758,N_21731);
xor U23124 (N_23124,N_21212,N_20082);
nand U23125 (N_23125,N_20678,N_21317);
xor U23126 (N_23126,N_20960,N_21133);
xnor U23127 (N_23127,N_21586,N_21775);
xor U23128 (N_23128,N_20931,N_21405);
nand U23129 (N_23129,N_21874,N_20806);
and U23130 (N_23130,N_21302,N_21349);
xor U23131 (N_23131,N_20641,N_21422);
and U23132 (N_23132,N_21228,N_20107);
or U23133 (N_23133,N_21437,N_21389);
and U23134 (N_23134,N_21440,N_20798);
or U23135 (N_23135,N_20353,N_20004);
xnor U23136 (N_23136,N_20914,N_21413);
xnor U23137 (N_23137,N_20289,N_20899);
nor U23138 (N_23138,N_21637,N_21811);
and U23139 (N_23139,N_20583,N_20996);
and U23140 (N_23140,N_20418,N_20945);
nor U23141 (N_23141,N_20592,N_21915);
or U23142 (N_23142,N_20139,N_20776);
or U23143 (N_23143,N_21326,N_20060);
nand U23144 (N_23144,N_21022,N_20594);
or U23145 (N_23145,N_20759,N_20161);
or U23146 (N_23146,N_20201,N_20440);
or U23147 (N_23147,N_21031,N_21167);
nand U23148 (N_23148,N_20036,N_20636);
or U23149 (N_23149,N_20759,N_20635);
xor U23150 (N_23150,N_20303,N_20091);
or U23151 (N_23151,N_21019,N_20711);
nor U23152 (N_23152,N_20950,N_21913);
nor U23153 (N_23153,N_21350,N_21013);
and U23154 (N_23154,N_21767,N_20082);
xnor U23155 (N_23155,N_20611,N_20631);
and U23156 (N_23156,N_20195,N_21089);
nand U23157 (N_23157,N_21637,N_21055);
nor U23158 (N_23158,N_20309,N_20535);
nand U23159 (N_23159,N_20812,N_21920);
nor U23160 (N_23160,N_21905,N_21493);
nand U23161 (N_23161,N_21817,N_20206);
and U23162 (N_23162,N_20402,N_21763);
xnor U23163 (N_23163,N_21238,N_21723);
and U23164 (N_23164,N_21083,N_20690);
or U23165 (N_23165,N_20129,N_20788);
xnor U23166 (N_23166,N_21432,N_20657);
nor U23167 (N_23167,N_21197,N_21909);
nand U23168 (N_23168,N_21841,N_21900);
or U23169 (N_23169,N_21404,N_20726);
xor U23170 (N_23170,N_21247,N_21306);
nor U23171 (N_23171,N_20611,N_20542);
or U23172 (N_23172,N_21341,N_20038);
nand U23173 (N_23173,N_21392,N_20078);
nor U23174 (N_23174,N_20084,N_21784);
or U23175 (N_23175,N_20645,N_21668);
or U23176 (N_23176,N_21858,N_20791);
or U23177 (N_23177,N_20031,N_20246);
nand U23178 (N_23178,N_21566,N_21663);
nand U23179 (N_23179,N_21392,N_21367);
nand U23180 (N_23180,N_21366,N_20944);
nor U23181 (N_23181,N_20299,N_20022);
nand U23182 (N_23182,N_20885,N_21026);
or U23183 (N_23183,N_20630,N_20555);
nand U23184 (N_23184,N_21244,N_20135);
xor U23185 (N_23185,N_21615,N_21755);
and U23186 (N_23186,N_20458,N_21769);
or U23187 (N_23187,N_20392,N_21762);
and U23188 (N_23188,N_21831,N_20269);
nand U23189 (N_23189,N_21903,N_21567);
nor U23190 (N_23190,N_20779,N_21020);
xnor U23191 (N_23191,N_20466,N_21275);
xnor U23192 (N_23192,N_20333,N_21486);
or U23193 (N_23193,N_20644,N_21874);
or U23194 (N_23194,N_21916,N_21979);
nor U23195 (N_23195,N_20632,N_21427);
nor U23196 (N_23196,N_20992,N_20241);
nor U23197 (N_23197,N_20893,N_21753);
and U23198 (N_23198,N_20409,N_21991);
and U23199 (N_23199,N_21765,N_21049);
nor U23200 (N_23200,N_21342,N_21634);
nand U23201 (N_23201,N_21115,N_20525);
nand U23202 (N_23202,N_21484,N_21093);
xor U23203 (N_23203,N_21525,N_20156);
nand U23204 (N_23204,N_20250,N_21498);
nor U23205 (N_23205,N_21504,N_21311);
xor U23206 (N_23206,N_21717,N_20733);
nor U23207 (N_23207,N_20534,N_20370);
xnor U23208 (N_23208,N_20742,N_20655);
or U23209 (N_23209,N_21657,N_21344);
nand U23210 (N_23210,N_21899,N_21643);
nand U23211 (N_23211,N_20069,N_20873);
xnor U23212 (N_23212,N_21801,N_21397);
and U23213 (N_23213,N_20567,N_21069);
or U23214 (N_23214,N_21208,N_20024);
or U23215 (N_23215,N_20704,N_20925);
and U23216 (N_23216,N_20580,N_20849);
nand U23217 (N_23217,N_20105,N_20323);
nor U23218 (N_23218,N_20885,N_20176);
xor U23219 (N_23219,N_20454,N_21913);
or U23220 (N_23220,N_21381,N_21818);
or U23221 (N_23221,N_21064,N_20722);
or U23222 (N_23222,N_20946,N_21915);
nand U23223 (N_23223,N_21595,N_21927);
nor U23224 (N_23224,N_21752,N_20143);
nand U23225 (N_23225,N_20208,N_20411);
and U23226 (N_23226,N_21116,N_21033);
nor U23227 (N_23227,N_20364,N_20903);
and U23228 (N_23228,N_20181,N_21695);
or U23229 (N_23229,N_20458,N_20105);
nand U23230 (N_23230,N_21744,N_20789);
and U23231 (N_23231,N_20270,N_20888);
nor U23232 (N_23232,N_21776,N_20488);
or U23233 (N_23233,N_21555,N_21164);
xor U23234 (N_23234,N_21637,N_21022);
nand U23235 (N_23235,N_21785,N_20617);
nor U23236 (N_23236,N_20955,N_21572);
nor U23237 (N_23237,N_21792,N_20506);
nor U23238 (N_23238,N_21229,N_21718);
xnor U23239 (N_23239,N_21897,N_21297);
and U23240 (N_23240,N_21974,N_21322);
or U23241 (N_23241,N_20366,N_20952);
nand U23242 (N_23242,N_20509,N_21019);
xnor U23243 (N_23243,N_20140,N_21277);
nor U23244 (N_23244,N_20866,N_20967);
nand U23245 (N_23245,N_21380,N_21639);
xnor U23246 (N_23246,N_20035,N_21033);
nor U23247 (N_23247,N_21680,N_20607);
and U23248 (N_23248,N_21759,N_21046);
nand U23249 (N_23249,N_20934,N_21869);
nor U23250 (N_23250,N_20707,N_20019);
xor U23251 (N_23251,N_21590,N_20327);
nand U23252 (N_23252,N_21114,N_20619);
nor U23253 (N_23253,N_21696,N_20121);
or U23254 (N_23254,N_21152,N_21283);
xor U23255 (N_23255,N_20309,N_21874);
and U23256 (N_23256,N_21024,N_21143);
or U23257 (N_23257,N_21919,N_20193);
xnor U23258 (N_23258,N_20400,N_21248);
or U23259 (N_23259,N_20603,N_20504);
nand U23260 (N_23260,N_20328,N_21673);
xnor U23261 (N_23261,N_20262,N_21150);
and U23262 (N_23262,N_20863,N_20487);
and U23263 (N_23263,N_20164,N_20293);
or U23264 (N_23264,N_21798,N_21413);
xnor U23265 (N_23265,N_20717,N_20348);
nand U23266 (N_23266,N_21057,N_21206);
and U23267 (N_23267,N_21185,N_20126);
or U23268 (N_23268,N_21937,N_21316);
and U23269 (N_23269,N_20038,N_21655);
xnor U23270 (N_23270,N_21010,N_21368);
nand U23271 (N_23271,N_20324,N_21849);
nor U23272 (N_23272,N_20337,N_21835);
nor U23273 (N_23273,N_21752,N_20675);
nor U23274 (N_23274,N_21893,N_21533);
xnor U23275 (N_23275,N_21650,N_20237);
nor U23276 (N_23276,N_20121,N_21861);
and U23277 (N_23277,N_20683,N_21916);
nor U23278 (N_23278,N_21555,N_20394);
and U23279 (N_23279,N_20498,N_20497);
and U23280 (N_23280,N_21216,N_21843);
nand U23281 (N_23281,N_21441,N_21843);
and U23282 (N_23282,N_21641,N_20249);
and U23283 (N_23283,N_20485,N_20492);
xnor U23284 (N_23284,N_20369,N_20569);
xor U23285 (N_23285,N_20150,N_20592);
xnor U23286 (N_23286,N_21203,N_20084);
nor U23287 (N_23287,N_20991,N_21188);
nand U23288 (N_23288,N_20830,N_20263);
nand U23289 (N_23289,N_21780,N_20185);
and U23290 (N_23290,N_21062,N_20277);
or U23291 (N_23291,N_21869,N_21775);
nand U23292 (N_23292,N_21538,N_21198);
xor U23293 (N_23293,N_21573,N_21815);
nand U23294 (N_23294,N_21785,N_20027);
nand U23295 (N_23295,N_21640,N_20583);
or U23296 (N_23296,N_21816,N_20227);
nand U23297 (N_23297,N_21818,N_20526);
xor U23298 (N_23298,N_21414,N_20232);
and U23299 (N_23299,N_21501,N_21834);
nand U23300 (N_23300,N_20569,N_20843);
nand U23301 (N_23301,N_21011,N_20965);
and U23302 (N_23302,N_20816,N_21010);
and U23303 (N_23303,N_21552,N_21001);
or U23304 (N_23304,N_20602,N_20655);
nor U23305 (N_23305,N_20451,N_20204);
nor U23306 (N_23306,N_20978,N_21295);
nor U23307 (N_23307,N_20501,N_20138);
nor U23308 (N_23308,N_20739,N_21949);
xnor U23309 (N_23309,N_21739,N_21025);
nor U23310 (N_23310,N_20442,N_20365);
xor U23311 (N_23311,N_20464,N_21690);
nand U23312 (N_23312,N_20001,N_21005);
nand U23313 (N_23313,N_21034,N_20507);
and U23314 (N_23314,N_21207,N_20116);
and U23315 (N_23315,N_20223,N_21534);
or U23316 (N_23316,N_20912,N_21380);
nand U23317 (N_23317,N_20910,N_21013);
nand U23318 (N_23318,N_20317,N_21306);
or U23319 (N_23319,N_20687,N_20316);
xor U23320 (N_23320,N_21480,N_20854);
or U23321 (N_23321,N_21184,N_21060);
xnor U23322 (N_23322,N_20053,N_20991);
or U23323 (N_23323,N_20258,N_20362);
xnor U23324 (N_23324,N_21125,N_20402);
nor U23325 (N_23325,N_20271,N_21907);
nor U23326 (N_23326,N_20043,N_21264);
and U23327 (N_23327,N_20634,N_20588);
nand U23328 (N_23328,N_21859,N_21134);
nor U23329 (N_23329,N_20298,N_21092);
and U23330 (N_23330,N_21828,N_20960);
or U23331 (N_23331,N_21951,N_20302);
xor U23332 (N_23332,N_21165,N_21990);
or U23333 (N_23333,N_20169,N_21030);
xor U23334 (N_23334,N_21499,N_20677);
and U23335 (N_23335,N_20630,N_21821);
xor U23336 (N_23336,N_20898,N_21443);
and U23337 (N_23337,N_20812,N_21036);
nor U23338 (N_23338,N_20660,N_20168);
or U23339 (N_23339,N_20850,N_20691);
nand U23340 (N_23340,N_20155,N_20066);
nand U23341 (N_23341,N_21460,N_20211);
or U23342 (N_23342,N_20100,N_20934);
nand U23343 (N_23343,N_20325,N_21221);
and U23344 (N_23344,N_20225,N_21459);
and U23345 (N_23345,N_20464,N_21817);
nor U23346 (N_23346,N_20420,N_20151);
or U23347 (N_23347,N_21271,N_20605);
nor U23348 (N_23348,N_21837,N_20974);
and U23349 (N_23349,N_20089,N_20947);
or U23350 (N_23350,N_20923,N_21643);
nor U23351 (N_23351,N_21856,N_20652);
xor U23352 (N_23352,N_21248,N_21667);
nand U23353 (N_23353,N_20115,N_21442);
and U23354 (N_23354,N_21290,N_20436);
or U23355 (N_23355,N_21536,N_20872);
nand U23356 (N_23356,N_21569,N_20295);
and U23357 (N_23357,N_21639,N_20056);
and U23358 (N_23358,N_20478,N_20684);
nor U23359 (N_23359,N_20993,N_20577);
nor U23360 (N_23360,N_20787,N_21339);
and U23361 (N_23361,N_21283,N_21638);
nor U23362 (N_23362,N_21436,N_20277);
and U23363 (N_23363,N_21067,N_20449);
xor U23364 (N_23364,N_20485,N_20621);
nor U23365 (N_23365,N_20951,N_20845);
and U23366 (N_23366,N_21541,N_20853);
nor U23367 (N_23367,N_20721,N_20853);
xnor U23368 (N_23368,N_20733,N_20384);
nand U23369 (N_23369,N_20515,N_21065);
and U23370 (N_23370,N_21169,N_20067);
or U23371 (N_23371,N_21097,N_20414);
and U23372 (N_23372,N_21415,N_21866);
xor U23373 (N_23373,N_20433,N_20766);
nor U23374 (N_23374,N_21540,N_21306);
xor U23375 (N_23375,N_21221,N_21461);
xnor U23376 (N_23376,N_21543,N_21132);
and U23377 (N_23377,N_21454,N_21989);
xor U23378 (N_23378,N_20594,N_21273);
xor U23379 (N_23379,N_21531,N_20919);
nand U23380 (N_23380,N_21392,N_21323);
and U23381 (N_23381,N_20740,N_20727);
nand U23382 (N_23382,N_21626,N_21541);
nand U23383 (N_23383,N_20343,N_21824);
nand U23384 (N_23384,N_21484,N_21593);
or U23385 (N_23385,N_20478,N_21498);
nor U23386 (N_23386,N_20718,N_21776);
nand U23387 (N_23387,N_21175,N_20341);
and U23388 (N_23388,N_20474,N_20604);
and U23389 (N_23389,N_20734,N_21579);
or U23390 (N_23390,N_20805,N_20234);
and U23391 (N_23391,N_21592,N_21804);
or U23392 (N_23392,N_21937,N_21742);
nor U23393 (N_23393,N_20741,N_20094);
xnor U23394 (N_23394,N_20347,N_21583);
xor U23395 (N_23395,N_20872,N_20354);
and U23396 (N_23396,N_21455,N_21155);
nand U23397 (N_23397,N_21436,N_21299);
nor U23398 (N_23398,N_20012,N_20831);
or U23399 (N_23399,N_20568,N_20430);
or U23400 (N_23400,N_20723,N_20338);
and U23401 (N_23401,N_21157,N_21576);
xnor U23402 (N_23402,N_20801,N_20545);
and U23403 (N_23403,N_21222,N_20983);
and U23404 (N_23404,N_21553,N_21111);
nand U23405 (N_23405,N_21567,N_20366);
or U23406 (N_23406,N_21696,N_20486);
nand U23407 (N_23407,N_21757,N_21800);
or U23408 (N_23408,N_20850,N_20134);
xnor U23409 (N_23409,N_20586,N_20982);
nand U23410 (N_23410,N_20273,N_20152);
and U23411 (N_23411,N_21618,N_20325);
and U23412 (N_23412,N_21157,N_21302);
nand U23413 (N_23413,N_21990,N_21656);
xor U23414 (N_23414,N_21684,N_21013);
nor U23415 (N_23415,N_21112,N_21252);
nor U23416 (N_23416,N_20881,N_21898);
or U23417 (N_23417,N_20092,N_20614);
nand U23418 (N_23418,N_21757,N_21370);
and U23419 (N_23419,N_20996,N_20338);
nor U23420 (N_23420,N_21774,N_21565);
xor U23421 (N_23421,N_20485,N_21203);
nor U23422 (N_23422,N_21196,N_20897);
or U23423 (N_23423,N_21183,N_21734);
and U23424 (N_23424,N_21023,N_20460);
and U23425 (N_23425,N_20222,N_20295);
nand U23426 (N_23426,N_21612,N_20038);
nor U23427 (N_23427,N_20388,N_21681);
or U23428 (N_23428,N_20266,N_20102);
or U23429 (N_23429,N_21464,N_20611);
xnor U23430 (N_23430,N_20381,N_20489);
and U23431 (N_23431,N_21829,N_21029);
xor U23432 (N_23432,N_20478,N_21825);
or U23433 (N_23433,N_20112,N_20940);
nand U23434 (N_23434,N_20552,N_20604);
xnor U23435 (N_23435,N_21559,N_20491);
and U23436 (N_23436,N_21783,N_21123);
nor U23437 (N_23437,N_21063,N_20149);
nor U23438 (N_23438,N_21736,N_21752);
nor U23439 (N_23439,N_21051,N_20387);
nand U23440 (N_23440,N_20010,N_20042);
xnor U23441 (N_23441,N_20182,N_20934);
or U23442 (N_23442,N_20677,N_20741);
nor U23443 (N_23443,N_20852,N_21799);
and U23444 (N_23444,N_20716,N_20904);
xnor U23445 (N_23445,N_21772,N_21719);
or U23446 (N_23446,N_21658,N_21705);
nor U23447 (N_23447,N_20749,N_21066);
nor U23448 (N_23448,N_21003,N_21105);
nor U23449 (N_23449,N_21027,N_20017);
nor U23450 (N_23450,N_21299,N_20989);
xor U23451 (N_23451,N_20446,N_20599);
nor U23452 (N_23452,N_20852,N_20390);
nor U23453 (N_23453,N_21074,N_21746);
and U23454 (N_23454,N_20323,N_21212);
nand U23455 (N_23455,N_20722,N_20460);
xnor U23456 (N_23456,N_20865,N_21527);
xor U23457 (N_23457,N_21109,N_20844);
and U23458 (N_23458,N_20966,N_20501);
xor U23459 (N_23459,N_20159,N_21971);
or U23460 (N_23460,N_20125,N_20431);
or U23461 (N_23461,N_21596,N_20809);
nand U23462 (N_23462,N_21814,N_21752);
nor U23463 (N_23463,N_21098,N_20764);
nor U23464 (N_23464,N_21761,N_21162);
and U23465 (N_23465,N_20230,N_21272);
xnor U23466 (N_23466,N_20419,N_21612);
or U23467 (N_23467,N_20820,N_20731);
nand U23468 (N_23468,N_20413,N_20264);
nand U23469 (N_23469,N_21298,N_20410);
or U23470 (N_23470,N_20240,N_20617);
and U23471 (N_23471,N_20923,N_21268);
or U23472 (N_23472,N_20576,N_21888);
nor U23473 (N_23473,N_20349,N_20812);
and U23474 (N_23474,N_20864,N_21830);
xnor U23475 (N_23475,N_21241,N_21067);
xnor U23476 (N_23476,N_21244,N_20493);
xor U23477 (N_23477,N_21915,N_20899);
xor U23478 (N_23478,N_21646,N_21333);
xnor U23479 (N_23479,N_20097,N_21128);
and U23480 (N_23480,N_21439,N_20190);
nor U23481 (N_23481,N_20768,N_21261);
nor U23482 (N_23482,N_20158,N_20313);
xnor U23483 (N_23483,N_21615,N_21984);
xnor U23484 (N_23484,N_21343,N_21477);
and U23485 (N_23485,N_20370,N_21663);
or U23486 (N_23486,N_20760,N_20160);
xnor U23487 (N_23487,N_21218,N_21823);
nand U23488 (N_23488,N_21594,N_20934);
nor U23489 (N_23489,N_20787,N_20585);
and U23490 (N_23490,N_20203,N_20617);
or U23491 (N_23491,N_20901,N_21245);
or U23492 (N_23492,N_20098,N_20032);
nor U23493 (N_23493,N_21855,N_20930);
nor U23494 (N_23494,N_21841,N_21552);
nand U23495 (N_23495,N_20880,N_20285);
and U23496 (N_23496,N_21763,N_21985);
or U23497 (N_23497,N_21500,N_21459);
and U23498 (N_23498,N_21752,N_20250);
xor U23499 (N_23499,N_21966,N_20915);
or U23500 (N_23500,N_20074,N_21882);
nand U23501 (N_23501,N_21254,N_21843);
nand U23502 (N_23502,N_20259,N_20015);
nor U23503 (N_23503,N_20311,N_21665);
xor U23504 (N_23504,N_20016,N_20357);
xor U23505 (N_23505,N_21822,N_21797);
nand U23506 (N_23506,N_21607,N_21655);
xor U23507 (N_23507,N_20839,N_20393);
xnor U23508 (N_23508,N_20906,N_21169);
nor U23509 (N_23509,N_20453,N_20305);
or U23510 (N_23510,N_20385,N_21555);
and U23511 (N_23511,N_20385,N_21082);
nor U23512 (N_23512,N_20972,N_21122);
xor U23513 (N_23513,N_21450,N_21975);
xnor U23514 (N_23514,N_20843,N_21533);
nand U23515 (N_23515,N_21052,N_20769);
or U23516 (N_23516,N_20363,N_20144);
or U23517 (N_23517,N_20515,N_21641);
xnor U23518 (N_23518,N_21241,N_21359);
or U23519 (N_23519,N_21748,N_20480);
or U23520 (N_23520,N_21079,N_21930);
or U23521 (N_23521,N_21940,N_20080);
nor U23522 (N_23522,N_20715,N_21771);
or U23523 (N_23523,N_20747,N_21343);
and U23524 (N_23524,N_21085,N_20611);
xor U23525 (N_23525,N_20080,N_20795);
xor U23526 (N_23526,N_21326,N_21331);
nand U23527 (N_23527,N_21099,N_20859);
nor U23528 (N_23528,N_20277,N_20864);
xnor U23529 (N_23529,N_20326,N_20956);
xnor U23530 (N_23530,N_20266,N_20800);
and U23531 (N_23531,N_20725,N_21586);
nor U23532 (N_23532,N_21442,N_20855);
or U23533 (N_23533,N_20643,N_20525);
xnor U23534 (N_23534,N_21089,N_20826);
or U23535 (N_23535,N_21129,N_20974);
or U23536 (N_23536,N_21327,N_21084);
xor U23537 (N_23537,N_21353,N_21065);
xor U23538 (N_23538,N_21479,N_21746);
or U23539 (N_23539,N_21622,N_21654);
or U23540 (N_23540,N_20072,N_20896);
nand U23541 (N_23541,N_20087,N_21057);
and U23542 (N_23542,N_21411,N_21086);
xnor U23543 (N_23543,N_21070,N_20740);
and U23544 (N_23544,N_20377,N_20553);
or U23545 (N_23545,N_20913,N_21309);
xnor U23546 (N_23546,N_20010,N_20513);
nor U23547 (N_23547,N_21270,N_20146);
nand U23548 (N_23548,N_20758,N_21453);
nor U23549 (N_23549,N_21561,N_20577);
or U23550 (N_23550,N_20002,N_21482);
nand U23551 (N_23551,N_20625,N_21862);
xnor U23552 (N_23552,N_21459,N_20203);
nor U23553 (N_23553,N_20993,N_21119);
or U23554 (N_23554,N_21537,N_20756);
or U23555 (N_23555,N_21395,N_21274);
nand U23556 (N_23556,N_21575,N_21307);
and U23557 (N_23557,N_20414,N_21898);
xnor U23558 (N_23558,N_21942,N_20501);
nor U23559 (N_23559,N_21538,N_21412);
or U23560 (N_23560,N_20910,N_21386);
and U23561 (N_23561,N_21615,N_20175);
or U23562 (N_23562,N_21710,N_20879);
nor U23563 (N_23563,N_20014,N_20690);
nor U23564 (N_23564,N_20471,N_20452);
or U23565 (N_23565,N_20863,N_21770);
nand U23566 (N_23566,N_21850,N_21095);
or U23567 (N_23567,N_20382,N_21281);
or U23568 (N_23568,N_21908,N_20768);
xor U23569 (N_23569,N_20948,N_20232);
nor U23570 (N_23570,N_21854,N_20877);
and U23571 (N_23571,N_21966,N_20794);
and U23572 (N_23572,N_20726,N_21999);
nor U23573 (N_23573,N_21264,N_21173);
or U23574 (N_23574,N_20095,N_21803);
and U23575 (N_23575,N_20235,N_21248);
and U23576 (N_23576,N_21665,N_21526);
and U23577 (N_23577,N_21658,N_20801);
and U23578 (N_23578,N_20046,N_20099);
and U23579 (N_23579,N_20544,N_21153);
nand U23580 (N_23580,N_21084,N_21993);
nor U23581 (N_23581,N_21801,N_21031);
or U23582 (N_23582,N_20016,N_21180);
nor U23583 (N_23583,N_20363,N_21881);
nand U23584 (N_23584,N_21429,N_21136);
and U23585 (N_23585,N_21215,N_20987);
nand U23586 (N_23586,N_21405,N_20990);
nand U23587 (N_23587,N_21535,N_21050);
and U23588 (N_23588,N_21212,N_21943);
and U23589 (N_23589,N_20407,N_21097);
xnor U23590 (N_23590,N_20004,N_21325);
nor U23591 (N_23591,N_21477,N_20192);
or U23592 (N_23592,N_21065,N_20208);
nor U23593 (N_23593,N_20228,N_21008);
xor U23594 (N_23594,N_21834,N_21254);
or U23595 (N_23595,N_20266,N_20196);
or U23596 (N_23596,N_20676,N_21852);
nor U23597 (N_23597,N_21039,N_20145);
nand U23598 (N_23598,N_21446,N_21033);
nand U23599 (N_23599,N_21465,N_20245);
xnor U23600 (N_23600,N_20757,N_21004);
or U23601 (N_23601,N_20379,N_21690);
nand U23602 (N_23602,N_21041,N_20365);
nor U23603 (N_23603,N_21590,N_21583);
xnor U23604 (N_23604,N_21448,N_21147);
or U23605 (N_23605,N_21371,N_20000);
nand U23606 (N_23606,N_21157,N_20285);
xnor U23607 (N_23607,N_21450,N_21277);
and U23608 (N_23608,N_21253,N_21382);
and U23609 (N_23609,N_20321,N_20531);
and U23610 (N_23610,N_20994,N_20213);
or U23611 (N_23611,N_21550,N_21047);
nand U23612 (N_23612,N_21561,N_20736);
or U23613 (N_23613,N_20780,N_20963);
nor U23614 (N_23614,N_20662,N_21235);
nand U23615 (N_23615,N_20070,N_20251);
nand U23616 (N_23616,N_21009,N_21430);
nor U23617 (N_23617,N_20807,N_21116);
or U23618 (N_23618,N_20317,N_21050);
nand U23619 (N_23619,N_20717,N_20269);
nor U23620 (N_23620,N_20564,N_21675);
or U23621 (N_23621,N_21205,N_20322);
nor U23622 (N_23622,N_21016,N_20791);
or U23623 (N_23623,N_21420,N_20712);
or U23624 (N_23624,N_21736,N_21937);
nand U23625 (N_23625,N_20114,N_20675);
and U23626 (N_23626,N_21650,N_21739);
nor U23627 (N_23627,N_21984,N_21183);
nand U23628 (N_23628,N_21090,N_20258);
nor U23629 (N_23629,N_20850,N_21173);
or U23630 (N_23630,N_20414,N_20038);
and U23631 (N_23631,N_20783,N_20904);
and U23632 (N_23632,N_20587,N_20689);
or U23633 (N_23633,N_20692,N_20583);
nor U23634 (N_23634,N_21529,N_21417);
or U23635 (N_23635,N_21173,N_21255);
and U23636 (N_23636,N_21696,N_21238);
nor U23637 (N_23637,N_21586,N_21929);
nor U23638 (N_23638,N_21450,N_21157);
nand U23639 (N_23639,N_20825,N_20594);
and U23640 (N_23640,N_21493,N_20768);
xor U23641 (N_23641,N_21418,N_21416);
and U23642 (N_23642,N_21307,N_21348);
nand U23643 (N_23643,N_21137,N_20864);
and U23644 (N_23644,N_20596,N_21979);
xnor U23645 (N_23645,N_21842,N_20981);
nand U23646 (N_23646,N_20591,N_21539);
and U23647 (N_23647,N_21945,N_20981);
nand U23648 (N_23648,N_21639,N_20965);
nor U23649 (N_23649,N_21168,N_21404);
and U23650 (N_23650,N_20679,N_20117);
nor U23651 (N_23651,N_20964,N_21835);
nand U23652 (N_23652,N_21530,N_21738);
xnor U23653 (N_23653,N_20036,N_21399);
nor U23654 (N_23654,N_21767,N_21513);
xor U23655 (N_23655,N_20449,N_21978);
or U23656 (N_23656,N_20421,N_21097);
or U23657 (N_23657,N_20462,N_20099);
xnor U23658 (N_23658,N_20810,N_20495);
and U23659 (N_23659,N_21592,N_20193);
and U23660 (N_23660,N_21520,N_20535);
or U23661 (N_23661,N_20040,N_21104);
nand U23662 (N_23662,N_21909,N_20866);
and U23663 (N_23663,N_21116,N_21497);
nor U23664 (N_23664,N_21868,N_21320);
nor U23665 (N_23665,N_20876,N_20808);
nand U23666 (N_23666,N_21082,N_20093);
and U23667 (N_23667,N_21111,N_21707);
nor U23668 (N_23668,N_21795,N_20916);
xor U23669 (N_23669,N_21301,N_21398);
xor U23670 (N_23670,N_20501,N_20503);
nor U23671 (N_23671,N_20301,N_20004);
and U23672 (N_23672,N_21471,N_21105);
and U23673 (N_23673,N_20331,N_21683);
xor U23674 (N_23674,N_20819,N_21021);
and U23675 (N_23675,N_20682,N_21521);
nor U23676 (N_23676,N_20534,N_20644);
nand U23677 (N_23677,N_21461,N_21274);
and U23678 (N_23678,N_21700,N_21601);
nor U23679 (N_23679,N_21119,N_20468);
or U23680 (N_23680,N_21320,N_21009);
xnor U23681 (N_23681,N_20572,N_20278);
or U23682 (N_23682,N_20165,N_20533);
xor U23683 (N_23683,N_20092,N_20454);
and U23684 (N_23684,N_21305,N_20856);
xnor U23685 (N_23685,N_21383,N_21951);
xnor U23686 (N_23686,N_20233,N_21140);
nor U23687 (N_23687,N_20364,N_20871);
nand U23688 (N_23688,N_21542,N_20075);
nand U23689 (N_23689,N_20125,N_20887);
nand U23690 (N_23690,N_20945,N_21029);
nand U23691 (N_23691,N_21054,N_20393);
or U23692 (N_23692,N_20293,N_21323);
nand U23693 (N_23693,N_20648,N_21665);
and U23694 (N_23694,N_20054,N_21351);
xnor U23695 (N_23695,N_21859,N_20831);
nor U23696 (N_23696,N_21788,N_20930);
xor U23697 (N_23697,N_20841,N_21872);
or U23698 (N_23698,N_21763,N_21719);
and U23699 (N_23699,N_20712,N_20497);
and U23700 (N_23700,N_20572,N_20157);
xor U23701 (N_23701,N_21656,N_20115);
or U23702 (N_23702,N_21071,N_20397);
and U23703 (N_23703,N_20603,N_21511);
or U23704 (N_23704,N_20929,N_20401);
and U23705 (N_23705,N_20065,N_21203);
nand U23706 (N_23706,N_20073,N_21699);
or U23707 (N_23707,N_20425,N_21343);
nand U23708 (N_23708,N_20995,N_21770);
nor U23709 (N_23709,N_21869,N_21898);
nor U23710 (N_23710,N_20558,N_21452);
xnor U23711 (N_23711,N_21164,N_21177);
nor U23712 (N_23712,N_20824,N_21233);
and U23713 (N_23713,N_21302,N_20120);
nor U23714 (N_23714,N_20868,N_21397);
xnor U23715 (N_23715,N_21664,N_20190);
nand U23716 (N_23716,N_21886,N_20058);
nor U23717 (N_23717,N_21217,N_21088);
xnor U23718 (N_23718,N_21087,N_21572);
nand U23719 (N_23719,N_20274,N_20546);
or U23720 (N_23720,N_21227,N_21677);
or U23721 (N_23721,N_20500,N_20755);
and U23722 (N_23722,N_20918,N_20545);
xnor U23723 (N_23723,N_21106,N_21166);
nand U23724 (N_23724,N_21874,N_20176);
nor U23725 (N_23725,N_20260,N_21921);
and U23726 (N_23726,N_21092,N_21935);
nand U23727 (N_23727,N_21351,N_20512);
or U23728 (N_23728,N_20886,N_21178);
or U23729 (N_23729,N_21509,N_20255);
nand U23730 (N_23730,N_20273,N_21854);
xor U23731 (N_23731,N_20822,N_21425);
xnor U23732 (N_23732,N_20561,N_21055);
nand U23733 (N_23733,N_21312,N_21647);
nand U23734 (N_23734,N_21908,N_21568);
nor U23735 (N_23735,N_20492,N_20530);
xnor U23736 (N_23736,N_21285,N_21719);
and U23737 (N_23737,N_21550,N_21775);
nand U23738 (N_23738,N_21895,N_21917);
nand U23739 (N_23739,N_21008,N_20100);
and U23740 (N_23740,N_20914,N_20501);
or U23741 (N_23741,N_21253,N_21007);
or U23742 (N_23742,N_20194,N_20307);
xor U23743 (N_23743,N_20608,N_20888);
nand U23744 (N_23744,N_20712,N_20918);
nand U23745 (N_23745,N_21242,N_20978);
nor U23746 (N_23746,N_21661,N_20000);
nand U23747 (N_23747,N_21934,N_21981);
or U23748 (N_23748,N_20280,N_20176);
nand U23749 (N_23749,N_21917,N_20287);
nor U23750 (N_23750,N_21536,N_21901);
and U23751 (N_23751,N_21246,N_21086);
nand U23752 (N_23752,N_21179,N_21255);
xor U23753 (N_23753,N_20693,N_20955);
and U23754 (N_23754,N_20994,N_21843);
xor U23755 (N_23755,N_21254,N_21430);
xor U23756 (N_23756,N_20259,N_20847);
or U23757 (N_23757,N_21147,N_20374);
or U23758 (N_23758,N_21113,N_20990);
and U23759 (N_23759,N_21324,N_21415);
and U23760 (N_23760,N_20741,N_20809);
nor U23761 (N_23761,N_21376,N_20842);
and U23762 (N_23762,N_21683,N_21585);
or U23763 (N_23763,N_20613,N_20855);
nor U23764 (N_23764,N_21012,N_21829);
nand U23765 (N_23765,N_21424,N_20807);
or U23766 (N_23766,N_21728,N_20893);
or U23767 (N_23767,N_20410,N_21345);
and U23768 (N_23768,N_21038,N_20561);
nor U23769 (N_23769,N_21825,N_20008);
and U23770 (N_23770,N_20413,N_20986);
or U23771 (N_23771,N_21872,N_21900);
xnor U23772 (N_23772,N_21664,N_21303);
nand U23773 (N_23773,N_21663,N_20666);
or U23774 (N_23774,N_20678,N_20104);
or U23775 (N_23775,N_21837,N_21252);
nand U23776 (N_23776,N_21939,N_21795);
nor U23777 (N_23777,N_20182,N_20945);
or U23778 (N_23778,N_21121,N_21001);
nor U23779 (N_23779,N_21777,N_20665);
and U23780 (N_23780,N_21539,N_21757);
or U23781 (N_23781,N_20382,N_20448);
nand U23782 (N_23782,N_20106,N_21960);
xnor U23783 (N_23783,N_21524,N_21625);
nand U23784 (N_23784,N_20492,N_21138);
xor U23785 (N_23785,N_21133,N_21713);
and U23786 (N_23786,N_21437,N_21550);
or U23787 (N_23787,N_21806,N_20311);
and U23788 (N_23788,N_21216,N_20956);
or U23789 (N_23789,N_21787,N_20402);
and U23790 (N_23790,N_21040,N_21740);
or U23791 (N_23791,N_21046,N_20369);
nand U23792 (N_23792,N_21810,N_21607);
nor U23793 (N_23793,N_21750,N_20667);
nor U23794 (N_23794,N_20099,N_21634);
nand U23795 (N_23795,N_20549,N_21900);
nor U23796 (N_23796,N_20388,N_21206);
and U23797 (N_23797,N_20175,N_20477);
and U23798 (N_23798,N_20522,N_21188);
nand U23799 (N_23799,N_20006,N_20322);
or U23800 (N_23800,N_21749,N_20099);
or U23801 (N_23801,N_20127,N_21931);
and U23802 (N_23802,N_21957,N_21416);
nor U23803 (N_23803,N_21158,N_21632);
and U23804 (N_23804,N_20974,N_20356);
or U23805 (N_23805,N_21019,N_21484);
and U23806 (N_23806,N_20473,N_21862);
and U23807 (N_23807,N_21236,N_21436);
and U23808 (N_23808,N_20397,N_21770);
nor U23809 (N_23809,N_20671,N_20446);
and U23810 (N_23810,N_21962,N_21631);
nand U23811 (N_23811,N_20965,N_20912);
nand U23812 (N_23812,N_21247,N_21865);
nor U23813 (N_23813,N_20154,N_21006);
xor U23814 (N_23814,N_21499,N_20183);
and U23815 (N_23815,N_20198,N_20630);
and U23816 (N_23816,N_21189,N_21295);
xor U23817 (N_23817,N_20135,N_21230);
and U23818 (N_23818,N_20605,N_20500);
nand U23819 (N_23819,N_21565,N_20033);
xnor U23820 (N_23820,N_20028,N_21379);
and U23821 (N_23821,N_21472,N_20820);
and U23822 (N_23822,N_21524,N_20889);
nor U23823 (N_23823,N_20103,N_20104);
and U23824 (N_23824,N_20061,N_21803);
and U23825 (N_23825,N_20989,N_21142);
nor U23826 (N_23826,N_21650,N_20212);
nor U23827 (N_23827,N_20843,N_21516);
nand U23828 (N_23828,N_21772,N_20241);
xor U23829 (N_23829,N_21774,N_20947);
nand U23830 (N_23830,N_21038,N_21373);
or U23831 (N_23831,N_21571,N_20309);
nand U23832 (N_23832,N_21477,N_20038);
nor U23833 (N_23833,N_21011,N_21583);
or U23834 (N_23834,N_21934,N_20416);
or U23835 (N_23835,N_20365,N_21037);
nor U23836 (N_23836,N_21046,N_21946);
nor U23837 (N_23837,N_20820,N_20985);
or U23838 (N_23838,N_21350,N_20137);
or U23839 (N_23839,N_20376,N_21812);
nand U23840 (N_23840,N_20298,N_20319);
xor U23841 (N_23841,N_21275,N_21397);
or U23842 (N_23842,N_20357,N_20682);
nand U23843 (N_23843,N_21523,N_20088);
xor U23844 (N_23844,N_21553,N_20179);
nand U23845 (N_23845,N_21998,N_21545);
nand U23846 (N_23846,N_21557,N_21617);
nor U23847 (N_23847,N_20546,N_21680);
nand U23848 (N_23848,N_20762,N_21380);
nand U23849 (N_23849,N_21365,N_21927);
nand U23850 (N_23850,N_21307,N_21276);
nand U23851 (N_23851,N_20750,N_21785);
nor U23852 (N_23852,N_21425,N_21640);
nor U23853 (N_23853,N_21489,N_21737);
nor U23854 (N_23854,N_20580,N_20897);
xor U23855 (N_23855,N_21242,N_20468);
or U23856 (N_23856,N_20651,N_20043);
and U23857 (N_23857,N_20164,N_21351);
nor U23858 (N_23858,N_21224,N_21749);
nand U23859 (N_23859,N_20130,N_20734);
nor U23860 (N_23860,N_21097,N_21663);
nand U23861 (N_23861,N_20237,N_21071);
or U23862 (N_23862,N_20978,N_21890);
nor U23863 (N_23863,N_21637,N_20154);
xor U23864 (N_23864,N_20075,N_20655);
nand U23865 (N_23865,N_20413,N_20907);
nand U23866 (N_23866,N_21349,N_21953);
nor U23867 (N_23867,N_20922,N_21308);
nor U23868 (N_23868,N_21515,N_20378);
nand U23869 (N_23869,N_21620,N_20844);
nor U23870 (N_23870,N_20217,N_20140);
nor U23871 (N_23871,N_20937,N_21966);
and U23872 (N_23872,N_20774,N_21188);
xnor U23873 (N_23873,N_21808,N_21374);
nor U23874 (N_23874,N_21575,N_20094);
nand U23875 (N_23875,N_20670,N_21793);
nand U23876 (N_23876,N_21912,N_21858);
nor U23877 (N_23877,N_21019,N_21421);
nor U23878 (N_23878,N_20794,N_21646);
and U23879 (N_23879,N_20999,N_20749);
nor U23880 (N_23880,N_20094,N_20170);
and U23881 (N_23881,N_21509,N_21155);
xor U23882 (N_23882,N_20959,N_21998);
or U23883 (N_23883,N_21307,N_21852);
or U23884 (N_23884,N_21615,N_20725);
xnor U23885 (N_23885,N_20663,N_20379);
or U23886 (N_23886,N_20908,N_21959);
or U23887 (N_23887,N_20360,N_20667);
nand U23888 (N_23888,N_20744,N_21120);
nor U23889 (N_23889,N_20783,N_21354);
nor U23890 (N_23890,N_21830,N_20059);
nand U23891 (N_23891,N_20998,N_20415);
and U23892 (N_23892,N_21450,N_20772);
nand U23893 (N_23893,N_20138,N_21021);
xor U23894 (N_23894,N_21859,N_21468);
or U23895 (N_23895,N_20911,N_21704);
xor U23896 (N_23896,N_20254,N_20564);
or U23897 (N_23897,N_21865,N_20331);
or U23898 (N_23898,N_21232,N_20390);
nor U23899 (N_23899,N_20892,N_21096);
and U23900 (N_23900,N_21826,N_20859);
xnor U23901 (N_23901,N_21951,N_21950);
or U23902 (N_23902,N_20172,N_21188);
or U23903 (N_23903,N_20138,N_20152);
or U23904 (N_23904,N_21616,N_20880);
nor U23905 (N_23905,N_21727,N_20414);
nand U23906 (N_23906,N_21734,N_21250);
xnor U23907 (N_23907,N_21486,N_20248);
nand U23908 (N_23908,N_21336,N_21718);
xor U23909 (N_23909,N_21438,N_20097);
nand U23910 (N_23910,N_20672,N_20338);
and U23911 (N_23911,N_21036,N_21765);
or U23912 (N_23912,N_21916,N_21240);
and U23913 (N_23913,N_21397,N_21848);
nor U23914 (N_23914,N_20775,N_20926);
xnor U23915 (N_23915,N_21715,N_20971);
xor U23916 (N_23916,N_20378,N_20753);
xor U23917 (N_23917,N_20821,N_20825);
or U23918 (N_23918,N_20736,N_20882);
and U23919 (N_23919,N_21628,N_21770);
and U23920 (N_23920,N_20836,N_21692);
or U23921 (N_23921,N_21300,N_20938);
and U23922 (N_23922,N_20698,N_21021);
and U23923 (N_23923,N_20916,N_21462);
or U23924 (N_23924,N_21949,N_20800);
nor U23925 (N_23925,N_21249,N_20738);
or U23926 (N_23926,N_20111,N_20128);
xor U23927 (N_23927,N_20402,N_21538);
xnor U23928 (N_23928,N_21590,N_21787);
nand U23929 (N_23929,N_20158,N_21162);
xnor U23930 (N_23930,N_21078,N_21330);
or U23931 (N_23931,N_21595,N_21651);
and U23932 (N_23932,N_21146,N_21408);
nor U23933 (N_23933,N_20821,N_21010);
xnor U23934 (N_23934,N_20924,N_21483);
or U23935 (N_23935,N_21344,N_20685);
nor U23936 (N_23936,N_20324,N_20234);
nor U23937 (N_23937,N_20676,N_20171);
and U23938 (N_23938,N_20130,N_21095);
nand U23939 (N_23939,N_20072,N_21478);
xnor U23940 (N_23940,N_21506,N_20811);
nand U23941 (N_23941,N_20423,N_21887);
nor U23942 (N_23942,N_21143,N_21404);
and U23943 (N_23943,N_21131,N_21136);
nand U23944 (N_23944,N_21189,N_20182);
or U23945 (N_23945,N_21056,N_20764);
and U23946 (N_23946,N_21157,N_20967);
nor U23947 (N_23947,N_20678,N_21415);
nand U23948 (N_23948,N_20321,N_20362);
nand U23949 (N_23949,N_21586,N_20021);
or U23950 (N_23950,N_20255,N_21343);
nor U23951 (N_23951,N_21127,N_20638);
nor U23952 (N_23952,N_20537,N_21304);
nor U23953 (N_23953,N_21217,N_21811);
nand U23954 (N_23954,N_21880,N_21584);
nor U23955 (N_23955,N_20461,N_21635);
nand U23956 (N_23956,N_20984,N_20133);
nor U23957 (N_23957,N_20746,N_20405);
nor U23958 (N_23958,N_20700,N_21871);
nor U23959 (N_23959,N_21921,N_21640);
or U23960 (N_23960,N_20827,N_21859);
and U23961 (N_23961,N_20988,N_21002);
or U23962 (N_23962,N_20839,N_20999);
and U23963 (N_23963,N_21812,N_20506);
and U23964 (N_23964,N_21341,N_21744);
nand U23965 (N_23965,N_20743,N_21902);
or U23966 (N_23966,N_21474,N_20195);
nor U23967 (N_23967,N_20283,N_20351);
or U23968 (N_23968,N_21903,N_20492);
xnor U23969 (N_23969,N_21129,N_21246);
or U23970 (N_23970,N_20739,N_21591);
nand U23971 (N_23971,N_21040,N_21790);
nand U23972 (N_23972,N_21924,N_21531);
nand U23973 (N_23973,N_20320,N_20768);
and U23974 (N_23974,N_21083,N_20931);
nand U23975 (N_23975,N_21284,N_20914);
or U23976 (N_23976,N_20409,N_21363);
xor U23977 (N_23977,N_20962,N_21191);
and U23978 (N_23978,N_20517,N_21179);
nor U23979 (N_23979,N_20986,N_21025);
xnor U23980 (N_23980,N_21850,N_20637);
or U23981 (N_23981,N_21839,N_21589);
nor U23982 (N_23982,N_20935,N_20499);
and U23983 (N_23983,N_20967,N_20222);
or U23984 (N_23984,N_20154,N_21789);
nand U23985 (N_23985,N_21652,N_20054);
or U23986 (N_23986,N_20180,N_21389);
xor U23987 (N_23987,N_21479,N_21449);
xnor U23988 (N_23988,N_20201,N_21034);
and U23989 (N_23989,N_21174,N_21876);
nor U23990 (N_23990,N_20265,N_21202);
xor U23991 (N_23991,N_21184,N_21138);
xor U23992 (N_23992,N_20839,N_21040);
xnor U23993 (N_23993,N_20792,N_21348);
nor U23994 (N_23994,N_20242,N_21060);
nor U23995 (N_23995,N_21663,N_20757);
and U23996 (N_23996,N_20340,N_21935);
xor U23997 (N_23997,N_20566,N_21420);
nand U23998 (N_23998,N_21261,N_21069);
or U23999 (N_23999,N_21512,N_20943);
nor U24000 (N_24000,N_23828,N_23067);
xor U24001 (N_24001,N_23405,N_22584);
xnor U24002 (N_24002,N_23306,N_22201);
xor U24003 (N_24003,N_22340,N_23732);
nor U24004 (N_24004,N_23330,N_23429);
and U24005 (N_24005,N_23111,N_23630);
nor U24006 (N_24006,N_23791,N_22695);
nor U24007 (N_24007,N_22539,N_23528);
and U24008 (N_24008,N_22650,N_22425);
nor U24009 (N_24009,N_23267,N_22687);
or U24010 (N_24010,N_22408,N_23259);
and U24011 (N_24011,N_22932,N_22752);
nor U24012 (N_24012,N_22352,N_22423);
xnor U24013 (N_24013,N_23491,N_22242);
xor U24014 (N_24014,N_23313,N_23045);
nor U24015 (N_24015,N_22249,N_23704);
and U24016 (N_24016,N_23304,N_22627);
xor U24017 (N_24017,N_22599,N_22476);
xor U24018 (N_24018,N_22371,N_23554);
or U24019 (N_24019,N_22037,N_22608);
nor U24020 (N_24020,N_22633,N_22648);
xor U24021 (N_24021,N_22130,N_23442);
nand U24022 (N_24022,N_22536,N_23492);
or U24023 (N_24023,N_22553,N_22422);
nand U24024 (N_24024,N_22732,N_23300);
and U24025 (N_24025,N_23724,N_23242);
nand U24026 (N_24026,N_23467,N_23290);
nand U24027 (N_24027,N_23224,N_23805);
nand U24028 (N_24028,N_22944,N_22898);
or U24029 (N_24029,N_22308,N_23503);
and U24030 (N_24030,N_22783,N_22176);
and U24031 (N_24031,N_22684,N_22796);
or U24032 (N_24032,N_23701,N_23777);
nand U24033 (N_24033,N_22670,N_22700);
and U24034 (N_24034,N_22400,N_22777);
nor U24035 (N_24035,N_22466,N_23591);
and U24036 (N_24036,N_22507,N_23870);
xor U24037 (N_24037,N_23678,N_22304);
and U24038 (N_24038,N_23628,N_22386);
or U24039 (N_24039,N_23097,N_23757);
or U24040 (N_24040,N_22624,N_23032);
xnor U24041 (N_24041,N_22985,N_23922);
and U24042 (N_24042,N_23855,N_23581);
xor U24043 (N_24043,N_22647,N_23090);
xor U24044 (N_24044,N_23022,N_22140);
or U24045 (N_24045,N_23472,N_22738);
or U24046 (N_24046,N_22078,N_22620);
nand U24047 (N_24047,N_23801,N_22988);
nand U24048 (N_24048,N_22026,N_22325);
nor U24049 (N_24049,N_22995,N_22157);
xnor U24050 (N_24050,N_23406,N_23399);
and U24051 (N_24051,N_23531,N_22493);
nor U24052 (N_24052,N_22162,N_22906);
nand U24053 (N_24053,N_23278,N_23241);
nor U24054 (N_24054,N_22012,N_23876);
and U24055 (N_24055,N_23138,N_22527);
and U24056 (N_24056,N_23151,N_23903);
xnor U24057 (N_24057,N_22188,N_22000);
xor U24058 (N_24058,N_23512,N_22896);
nand U24059 (N_24059,N_22744,N_23645);
nor U24060 (N_24060,N_23950,N_23066);
nand U24061 (N_24061,N_23793,N_23053);
nor U24062 (N_24062,N_23424,N_22150);
and U24063 (N_24063,N_23548,N_23599);
nor U24064 (N_24064,N_23122,N_23706);
and U24065 (N_24065,N_23418,N_23190);
nand U24066 (N_24066,N_22808,N_23946);
nor U24067 (N_24067,N_22879,N_23809);
xor U24068 (N_24068,N_23260,N_22893);
nand U24069 (N_24069,N_22267,N_23881);
and U24070 (N_24070,N_23089,N_22460);
and U24071 (N_24071,N_23532,N_22495);
xor U24072 (N_24072,N_22349,N_23525);
nor U24073 (N_24073,N_23507,N_23157);
nand U24074 (N_24074,N_22714,N_22745);
nor U24075 (N_24075,N_23380,N_23834);
and U24076 (N_24076,N_23981,N_22191);
nand U24077 (N_24077,N_23822,N_23667);
or U24078 (N_24078,N_23905,N_23520);
nor U24079 (N_24079,N_22285,N_23962);
and U24080 (N_24080,N_22913,N_23337);
xor U24081 (N_24081,N_23868,N_23617);
nor U24082 (N_24082,N_23501,N_23227);
and U24083 (N_24083,N_23314,N_23690);
and U24084 (N_24084,N_23573,N_23639);
or U24085 (N_24085,N_22617,N_23508);
nand U24086 (N_24086,N_23586,N_23686);
or U24087 (N_24087,N_23043,N_22543);
or U24088 (N_24088,N_23989,N_22046);
or U24089 (N_24089,N_23676,N_22256);
nand U24090 (N_24090,N_22595,N_22830);
or U24091 (N_24091,N_22215,N_22389);
xor U24092 (N_24092,N_23101,N_22924);
xor U24093 (N_24093,N_22917,N_23129);
nor U24094 (N_24094,N_23647,N_23450);
or U24095 (N_24095,N_23245,N_22148);
nor U24096 (N_24096,N_23545,N_22210);
xnor U24097 (N_24097,N_22071,N_23068);
or U24098 (N_24098,N_22982,N_23128);
or U24099 (N_24099,N_22205,N_23847);
and U24100 (N_24100,N_23863,N_22644);
and U24101 (N_24101,N_22713,N_23329);
and U24102 (N_24102,N_23017,N_23236);
xnor U24103 (N_24103,N_22014,N_23557);
nor U24104 (N_24104,N_23447,N_23204);
nor U24105 (N_24105,N_22383,N_22724);
and U24106 (N_24106,N_22002,N_22698);
or U24107 (N_24107,N_23749,N_23299);
nand U24108 (N_24108,N_23020,N_23815);
or U24109 (N_24109,N_22222,N_22113);
or U24110 (N_24110,N_23770,N_23028);
or U24111 (N_24111,N_22185,N_23481);
nand U24112 (N_24112,N_23265,N_22962);
nor U24113 (N_24113,N_23784,N_22231);
and U24114 (N_24114,N_22921,N_22846);
nand U24115 (N_24115,N_22861,N_22834);
and U24116 (N_24116,N_23535,N_23635);
nor U24117 (N_24117,N_23619,N_22845);
xor U24118 (N_24118,N_22407,N_22132);
nand U24119 (N_24119,N_23803,N_23490);
nand U24120 (N_24120,N_23445,N_23182);
or U24121 (N_24121,N_22709,N_22359);
and U24122 (N_24122,N_22467,N_22192);
xnor U24123 (N_24123,N_23268,N_22385);
and U24124 (N_24124,N_22935,N_23670);
and U24125 (N_24125,N_22248,N_22200);
nand U24126 (N_24126,N_23247,N_23335);
nor U24127 (N_24127,N_22520,N_22297);
xor U24128 (N_24128,N_22957,N_22811);
xor U24129 (N_24129,N_23297,N_23287);
nand U24130 (N_24130,N_23167,N_23195);
nor U24131 (N_24131,N_22060,N_22946);
or U24132 (N_24132,N_23907,N_22636);
or U24133 (N_24133,N_22265,N_23371);
and U24134 (N_24134,N_23911,N_22473);
xor U24135 (N_24135,N_22376,N_22426);
nand U24136 (N_24136,N_23715,N_23381);
and U24137 (N_24137,N_23956,N_23713);
nor U24138 (N_24138,N_23602,N_23483);
or U24139 (N_24139,N_22266,N_22331);
and U24140 (N_24140,N_23453,N_23438);
xor U24141 (N_24141,N_22427,N_23835);
or U24142 (N_24142,N_23369,N_23506);
nand U24143 (N_24143,N_22785,N_22829);
nor U24144 (N_24144,N_23428,N_22947);
and U24145 (N_24145,N_23149,N_22734);
or U24146 (N_24146,N_23585,N_22776);
xor U24147 (N_24147,N_22578,N_22848);
nor U24148 (N_24148,N_22526,N_22406);
nor U24149 (N_24149,N_22311,N_23353);
and U24150 (N_24150,N_22199,N_23363);
and U24151 (N_24151,N_22187,N_22902);
nand U24152 (N_24152,N_22051,N_23804);
xnor U24153 (N_24153,N_23159,N_23572);
nor U24154 (N_24154,N_22121,N_23885);
xor U24155 (N_24155,N_23720,N_22173);
and U24156 (N_24156,N_23192,N_22500);
and U24157 (N_24157,N_22807,N_23848);
nand U24158 (N_24158,N_22716,N_22914);
nand U24159 (N_24159,N_23347,N_22851);
and U24160 (N_24160,N_22705,N_22430);
and U24161 (N_24161,N_23158,N_22283);
or U24162 (N_24162,N_22496,N_22416);
xor U24163 (N_24163,N_22784,N_22490);
and U24164 (N_24164,N_22895,N_23637);
and U24165 (N_24165,N_23473,N_22803);
or U24166 (N_24166,N_22565,N_22293);
or U24167 (N_24167,N_23040,N_22577);
nand U24168 (N_24168,N_23030,N_23321);
and U24169 (N_24169,N_23431,N_22213);
and U24170 (N_24170,N_23665,N_23056);
nand U24171 (N_24171,N_22854,N_22429);
nand U24172 (N_24172,N_22263,N_22591);
and U24173 (N_24173,N_22609,N_23789);
nor U24174 (N_24174,N_22208,N_23048);
xnor U24175 (N_24175,N_22155,N_22890);
nand U24176 (N_24176,N_23331,N_22384);
nor U24177 (N_24177,N_23654,N_22125);
nand U24178 (N_24178,N_23634,N_23610);
and U24179 (N_24179,N_22262,N_22115);
nand U24180 (N_24180,N_23462,N_23559);
and U24181 (N_24181,N_23915,N_22072);
and U24182 (N_24182,N_23196,N_23609);
xnor U24183 (N_24183,N_22952,N_23705);
or U24184 (N_24184,N_23474,N_22719);
xnor U24185 (N_24185,N_22235,N_22598);
or U24186 (N_24186,N_23175,N_23824);
and U24187 (N_24187,N_23843,N_22382);
or U24188 (N_24188,N_22393,N_22418);
nand U24189 (N_24189,N_23294,N_22502);
xnor U24190 (N_24190,N_23739,N_22518);
nand U24191 (N_24191,N_23240,N_23320);
or U24192 (N_24192,N_22657,N_22669);
xor U24193 (N_24193,N_22509,N_23887);
nor U24194 (N_24194,N_22643,N_23046);
nor U24195 (N_24195,N_23465,N_22116);
nand U24196 (N_24196,N_22380,N_22471);
nor U24197 (N_24197,N_22540,N_23026);
xnor U24198 (N_24198,N_22711,N_22124);
or U24199 (N_24199,N_22552,N_22751);
and U24200 (N_24200,N_23312,N_22177);
nor U24201 (N_24201,N_23471,N_22064);
nand U24202 (N_24202,N_23711,N_23712);
xor U24203 (N_24203,N_23016,N_22750);
or U24204 (N_24204,N_22038,N_23833);
nand U24205 (N_24205,N_23451,N_22521);
nand U24206 (N_24206,N_22193,N_23727);
nor U24207 (N_24207,N_22146,N_22402);
nor U24208 (N_24208,N_23614,N_22542);
xnor U24209 (N_24209,N_22126,N_23914);
xnor U24210 (N_24210,N_23126,N_22198);
nand U24211 (N_24211,N_23475,N_23979);
nor U24212 (N_24212,N_22017,N_23194);
nor U24213 (N_24213,N_23376,N_23541);
nor U24214 (N_24214,N_23271,N_23695);
or U24215 (N_24215,N_22216,N_23315);
xor U24216 (N_24216,N_23094,N_23152);
or U24217 (N_24217,N_22619,N_23737);
nor U24218 (N_24218,N_22550,N_23011);
or U24219 (N_24219,N_22899,N_22149);
or U24220 (N_24220,N_22969,N_23041);
and U24221 (N_24221,N_23596,N_22922);
or U24222 (N_24222,N_22438,N_22301);
and U24223 (N_24223,N_22868,N_23656);
xor U24224 (N_24224,N_22761,N_22409);
xor U24225 (N_24225,N_23085,N_23411);
xor U24226 (N_24226,N_23936,N_23825);
or U24227 (N_24227,N_22703,N_23393);
and U24228 (N_24228,N_23958,N_23971);
nor U24229 (N_24229,N_22197,N_22976);
or U24230 (N_24230,N_23891,N_23487);
nand U24231 (N_24231,N_23064,N_23296);
nor U24232 (N_24232,N_23964,N_22747);
xor U24233 (N_24233,N_22101,N_23029);
and U24234 (N_24234,N_22175,N_23574);
or U24235 (N_24235,N_23781,N_22306);
nor U24236 (N_24236,N_23721,N_23975);
or U24237 (N_24237,N_23141,N_23199);
nand U24238 (N_24238,N_23148,N_22592);
or U24239 (N_24239,N_23857,N_22883);
and U24240 (N_24240,N_22322,N_23218);
xnor U24241 (N_24241,N_22091,N_23530);
nand U24242 (N_24242,N_23364,N_23529);
and U24243 (N_24243,N_22077,N_23555);
nor U24244 (N_24244,N_22887,N_22299);
or U24245 (N_24245,N_22978,N_23155);
or U24246 (N_24246,N_23957,N_23116);
xor U24247 (N_24247,N_22827,N_23864);
nand U24248 (N_24248,N_22907,N_22966);
xor U24249 (N_24249,N_23773,N_23622);
nor U24250 (N_24250,N_23323,N_22746);
or U24251 (N_24251,N_22601,N_23760);
nand U24252 (N_24252,N_22111,N_22492);
nor U24253 (N_24253,N_23896,N_23222);
nand U24254 (N_24254,N_23498,N_23049);
nor U24255 (N_24255,N_23980,N_23485);
and U24256 (N_24256,N_22207,N_22775);
nand U24257 (N_24257,N_22470,N_22920);
nor U24258 (N_24258,N_23435,N_22374);
and U24259 (N_24259,N_23354,N_22963);
xnor U24260 (N_24260,N_23894,N_22434);
and U24261 (N_24261,N_23550,N_23838);
or U24262 (N_24262,N_23093,N_22856);
and U24263 (N_24263,N_22128,N_23070);
and U24264 (N_24264,N_22459,N_22770);
nor U24265 (N_24265,N_22522,N_22945);
nand U24266 (N_24266,N_22481,N_23031);
nor U24267 (N_24267,N_23821,N_23303);
and U24268 (N_24268,N_23400,N_22779);
nor U24269 (N_24269,N_23687,N_22658);
nand U24270 (N_24270,N_23854,N_22998);
nand U24271 (N_24271,N_22715,N_22329);
nand U24272 (N_24272,N_22513,N_23493);
and U24273 (N_24273,N_22082,N_22478);
nand U24274 (N_24274,N_22635,N_22432);
nand U24275 (N_24275,N_22955,N_23496);
and U24276 (N_24276,N_23725,N_22833);
xnor U24277 (N_24277,N_23916,N_22821);
nand U24278 (N_24278,N_22264,N_22850);
nand U24279 (N_24279,N_23219,N_22597);
nor U24280 (N_24280,N_23792,N_23171);
nor U24281 (N_24281,N_23410,N_22606);
and U24282 (N_24282,N_23576,N_23307);
xor U24283 (N_24283,N_22160,N_22318);
and U24284 (N_24284,N_23547,N_23543);
xnor U24285 (N_24285,N_23909,N_23553);
or U24286 (N_24286,N_23302,N_23057);
or U24287 (N_24287,N_22449,N_22225);
nor U24288 (N_24288,N_23566,N_22270);
nor U24289 (N_24289,N_22277,N_22572);
or U24290 (N_24290,N_22835,N_23900);
and U24291 (N_24291,N_22486,N_22062);
nand U24292 (N_24292,N_23808,N_23598);
xor U24293 (N_24293,N_23753,N_23856);
nor U24294 (N_24294,N_23004,N_22673);
xnor U24295 (N_24295,N_23186,N_22036);
or U24296 (N_24296,N_22164,N_22085);
nor U24297 (N_24297,N_23154,N_23796);
nand U24298 (N_24298,N_22723,N_22656);
nor U24299 (N_24299,N_22344,N_22488);
nand U24300 (N_24300,N_22043,N_22630);
or U24301 (N_24301,N_22109,N_22491);
xnor U24302 (N_24302,N_22623,N_22610);
nand U24303 (N_24303,N_23193,N_22873);
and U24304 (N_24304,N_23800,N_22241);
nand U24305 (N_24305,N_22247,N_23918);
nand U24306 (N_24306,N_22039,N_22838);
xnor U24307 (N_24307,N_23270,N_22147);
nor U24308 (N_24308,N_22836,N_22424);
nand U24309 (N_24309,N_23412,N_22901);
and U24310 (N_24310,N_23849,N_23426);
nand U24311 (N_24311,N_22530,N_23661);
and U24312 (N_24312,N_22118,N_22613);
nand U24313 (N_24313,N_22871,N_23273);
xor U24314 (N_24314,N_23144,N_22886);
or U24315 (N_24315,N_23814,N_22433);
or U24316 (N_24316,N_23836,N_22787);
nor U24317 (N_24317,N_22568,N_23966);
nor U24318 (N_24318,N_22370,N_22279);
and U24319 (N_24319,N_22390,N_22455);
nand U24320 (N_24320,N_23858,N_22638);
or U24321 (N_24321,N_22720,N_22439);
nand U24322 (N_24322,N_22250,N_22992);
nand U24323 (N_24323,N_22693,N_23147);
or U24324 (N_24324,N_23209,N_23682);
xnor U24325 (N_24325,N_22727,N_22255);
and U24326 (N_24326,N_23624,N_22472);
nand U24327 (N_24327,N_22395,N_22120);
or U24328 (N_24328,N_22762,N_22204);
and U24329 (N_24329,N_22625,N_23044);
nor U24330 (N_24330,N_22240,N_23886);
xor U24331 (N_24331,N_22369,N_23456);
and U24332 (N_24332,N_23457,N_22135);
or U24333 (N_24333,N_22206,N_23762);
and U24334 (N_24334,N_23652,N_22928);
and U24335 (N_24335,N_23092,N_22379);
nand U24336 (N_24336,N_23142,N_23708);
xnor U24337 (N_24337,N_22748,N_23088);
and U24338 (N_24338,N_23134,N_23873);
nand U24339 (N_24339,N_22646,N_23850);
nor U24340 (N_24340,N_23375,N_22622);
nand U24341 (N_24341,N_23787,N_23767);
nand U24342 (N_24342,N_23461,N_22044);
nor U24343 (N_24343,N_22034,N_22866);
or U24344 (N_24344,N_23488,N_23365);
or U24345 (N_24345,N_23477,N_23058);
nand U24346 (N_24346,N_23276,N_23899);
nor U24347 (N_24347,N_23582,N_23379);
or U24348 (N_24348,N_23414,N_23208);
xnor U24349 (N_24349,N_22212,N_23441);
and U24350 (N_24350,N_22954,N_23766);
xor U24351 (N_24351,N_22765,N_23875);
and U24352 (N_24352,N_23370,N_23707);
nor U24353 (N_24353,N_22575,N_23763);
and U24354 (N_24354,N_22602,N_23683);
nand U24355 (N_24355,N_23594,N_22671);
and U24356 (N_24356,N_23898,N_22327);
and U24357 (N_24357,N_23003,N_22863);
xor U24358 (N_24358,N_23693,N_22964);
nor U24359 (N_24359,N_23829,N_23216);
xnor U24360 (N_24360,N_23967,N_23575);
or U24361 (N_24361,N_23060,N_23206);
nor U24362 (N_24362,N_23169,N_22942);
nand U24363 (N_24363,N_22021,N_23564);
xnor U24364 (N_24364,N_22537,N_22637);
xnor U24365 (N_24365,N_22755,N_22020);
xor U24366 (N_24366,N_22586,N_23768);
nor U24367 (N_24367,N_22431,N_23357);
nand U24368 (N_24368,N_22708,N_23166);
xor U24369 (N_24369,N_22313,N_22566);
nor U24370 (N_24370,N_23389,N_22047);
and U24371 (N_24371,N_22563,N_22826);
and U24372 (N_24372,N_22812,N_23377);
or U24373 (N_24373,N_23181,N_23785);
and U24374 (N_24374,N_23926,N_22639);
and U24375 (N_24375,N_23565,N_23524);
nand U24376 (N_24376,N_22234,N_22391);
or U24377 (N_24377,N_23225,N_22025);
and U24378 (N_24378,N_22166,N_23317);
xnor U24379 (N_24379,N_23051,N_23062);
nor U24380 (N_24380,N_22011,N_23927);
and U24381 (N_24381,N_22084,N_23065);
nand U24382 (N_24382,N_23510,N_23755);
nor U24383 (N_24383,N_22579,N_23742);
nand U24384 (N_24384,N_23925,N_23336);
xor U24385 (N_24385,N_23819,N_23679);
or U24386 (N_24386,N_23231,N_23769);
and U24387 (N_24387,N_22981,N_23761);
nor U24388 (N_24388,N_23215,N_22736);
nand U24389 (N_24389,N_22079,N_22678);
or U24390 (N_24390,N_22681,N_22223);
nor U24391 (N_24391,N_22209,N_22345);
xor U24392 (N_24392,N_22098,N_23527);
xnor U24393 (N_24393,N_23648,N_23923);
nor U24394 (N_24394,N_22768,N_22810);
and U24395 (N_24395,N_23251,N_22063);
nor U24396 (N_24396,N_23845,N_23396);
or U24397 (N_24397,N_23098,N_22066);
nor U24398 (N_24398,N_22224,N_22324);
and U24399 (N_24399,N_22652,N_22645);
nand U24400 (N_24400,N_23908,N_22961);
or U24401 (N_24401,N_22663,N_22479);
xor U24402 (N_24402,N_22501,N_22702);
or U24403 (N_24403,N_23608,N_22372);
nor U24404 (N_24404,N_23672,N_22328);
and U24405 (N_24405,N_23807,N_22824);
and U24406 (N_24406,N_23253,N_22517);
nand U24407 (N_24407,N_22603,N_22320);
nand U24408 (N_24408,N_23741,N_22589);
or U24409 (N_24409,N_22287,N_23746);
nor U24410 (N_24410,N_22106,N_22254);
xor U24411 (N_24411,N_23673,N_23425);
or U24412 (N_24412,N_22972,N_22554);
nor U24413 (N_24413,N_23588,N_23963);
or U24414 (N_24414,N_22960,N_23621);
nor U24415 (N_24415,N_22641,N_23050);
nand U24416 (N_24416,N_22366,N_23165);
xnor U24417 (N_24417,N_23282,N_22070);
and U24418 (N_24418,N_22864,N_23878);
xnor U24419 (N_24419,N_23612,N_22076);
nand U24420 (N_24420,N_22401,N_23174);
and U24421 (N_24421,N_23580,N_22660);
xor U24422 (N_24422,N_22143,N_22823);
or U24423 (N_24423,N_22278,N_23865);
nor U24424 (N_24424,N_22381,N_22685);
nand U24425 (N_24425,N_22778,N_23099);
and U24426 (N_24426,N_23655,N_22243);
nand U24427 (N_24427,N_23366,N_22356);
and U24428 (N_24428,N_23178,N_23110);
nand U24429 (N_24429,N_23832,N_22281);
nand U24430 (N_24430,N_23201,N_23131);
nand U24431 (N_24431,N_23817,N_23019);
nand U24432 (N_24432,N_22233,N_23616);
nand U24433 (N_24433,N_23620,N_22769);
xor U24434 (N_24434,N_23327,N_23696);
or U24435 (N_24435,N_22558,N_23145);
nand U24436 (N_24436,N_22154,N_22798);
xnor U24437 (N_24437,N_23860,N_23538);
nor U24438 (N_24438,N_23626,N_23324);
nor U24439 (N_24439,N_23162,N_22487);
or U24440 (N_24440,N_23593,N_23284);
nor U24441 (N_24441,N_23096,N_23592);
xnor U24442 (N_24442,N_22268,N_22549);
or U24443 (N_24443,N_23042,N_22582);
nor U24444 (N_24444,N_22252,N_22108);
or U24445 (N_24445,N_23177,N_22979);
nor U24446 (N_24446,N_22018,N_23434);
nand U24447 (N_24447,N_23984,N_23904);
xor U24448 (N_24448,N_23292,N_23942);
xnor U24449 (N_24449,N_22689,N_23458);
nand U24450 (N_24450,N_23500,N_23782);
xor U24451 (N_24451,N_23286,N_23797);
and U24452 (N_24452,N_22688,N_23205);
nand U24453 (N_24453,N_22911,N_22457);
and U24454 (N_24454,N_23944,N_22607);
nor U24455 (N_24455,N_23349,N_22008);
nand U24456 (N_24456,N_22035,N_22936);
xnor U24457 (N_24457,N_22544,N_22789);
nor U24458 (N_24458,N_22943,N_23680);
nor U24459 (N_24459,N_22334,N_23298);
nand U24460 (N_24460,N_23932,N_22837);
nor U24461 (N_24461,N_22123,N_23862);
or U24462 (N_24462,N_23289,N_23168);
nor U24463 (N_24463,N_23584,N_23571);
xor U24464 (N_24464,N_23308,N_23669);
nor U24465 (N_24465,N_22999,N_22326);
and U24466 (N_24466,N_22802,N_22170);
and U24467 (N_24467,N_22659,N_22525);
or U24468 (N_24468,N_23136,N_22184);
nor U24469 (N_24469,N_23879,N_22312);
xor U24470 (N_24470,N_23776,N_23627);
or U24471 (N_24471,N_23361,N_23484);
nand U24472 (N_24472,N_23750,N_22753);
xor U24473 (N_24473,N_23595,N_23256);
nand U24474 (N_24474,N_23470,N_22015);
nor U24475 (N_24475,N_22332,N_23124);
and U24476 (N_24476,N_22881,N_23851);
nor U24477 (N_24477,N_22341,N_22145);
or U24478 (N_24478,N_23035,N_23008);
and U24479 (N_24479,N_22168,N_23479);
or U24480 (N_24480,N_22977,N_23469);
or U24481 (N_24481,N_22891,N_22441);
or U24482 (N_24482,N_22712,N_23244);
xor U24483 (N_24483,N_23384,N_23318);
or U24484 (N_24484,N_23466,N_22953);
nand U24485 (N_24485,N_23600,N_23277);
nor U24486 (N_24486,N_22730,N_23698);
and U24487 (N_24487,N_22844,N_23691);
xnor U24488 (N_24488,N_23643,N_23937);
or U24489 (N_24489,N_23023,N_22217);
nand U24490 (N_24490,N_23988,N_22498);
xor U24491 (N_24491,N_22033,N_22559);
nand U24492 (N_24492,N_22004,N_22512);
nor U24493 (N_24493,N_23499,N_23568);
nor U24494 (N_24494,N_23059,N_22194);
nand U24495 (N_24495,N_22468,N_23104);
or U24496 (N_24496,N_23301,N_22594);
nor U24497 (N_24497,N_22323,N_23334);
xor U24498 (N_24498,N_23113,N_23478);
nor U24499 (N_24499,N_22667,N_22403);
nor U24500 (N_24500,N_22114,N_22272);
or U24501 (N_24501,N_22245,N_23589);
and U24502 (N_24502,N_22852,N_23120);
or U24503 (N_24503,N_23841,N_23081);
or U24504 (N_24504,N_22300,N_22909);
nor U24505 (N_24505,N_22528,N_22499);
and U24506 (N_24506,N_22878,N_22144);
nand U24507 (N_24507,N_23625,N_23671);
xor U24508 (N_24508,N_23125,N_23397);
xor U24509 (N_24509,N_22271,N_22075);
nor U24510 (N_24510,N_22275,N_23082);
or U24511 (N_24511,N_23272,N_22195);
nor U24512 (N_24512,N_22704,N_23869);
xnor U24513 (N_24513,N_22640,N_22339);
xnor U24514 (N_24514,N_22941,N_23108);
nand U24515 (N_24515,N_22590,N_23751);
and U24516 (N_24516,N_23709,N_23037);
or U24517 (N_24517,N_23533,N_22073);
nand U24518 (N_24518,N_23255,N_22174);
or U24519 (N_24519,N_23262,N_23788);
nor U24520 (N_24520,N_22997,N_22662);
xnor U24521 (N_24521,N_22048,N_22096);
nand U24522 (N_24522,N_22587,N_22806);
xor U24523 (N_24523,N_22127,N_22042);
nor U24524 (N_24524,N_22089,N_23987);
or U24525 (N_24525,N_22253,N_23552);
nand U24526 (N_24526,N_22503,N_23526);
nand U24527 (N_24527,N_23518,N_23722);
nor U24528 (N_24528,N_22182,N_23316);
or U24529 (N_24529,N_22355,N_22236);
nor U24530 (N_24530,N_22440,N_23080);
and U24531 (N_24531,N_22876,N_23119);
or U24532 (N_24532,N_22387,N_22417);
or U24533 (N_24533,N_23883,N_22869);
and U24534 (N_24534,N_23901,N_22405);
or U24535 (N_24535,N_22284,N_22413);
nand U24536 (N_24536,N_23605,N_22351);
or U24537 (N_24537,N_23074,N_22933);
nand U24538 (N_24538,N_22855,N_22691);
or U24539 (N_24539,N_22228,N_22158);
and U24540 (N_24540,N_22462,N_22083);
or U24541 (N_24541,N_22937,N_23332);
or U24542 (N_24542,N_23419,N_22560);
nand U24543 (N_24543,N_23997,N_22975);
xnor U24544 (N_24544,N_22364,N_22302);
nor U24545 (N_24545,N_22742,N_23563);
nand U24546 (N_24546,N_22749,N_22257);
nor U24547 (N_24547,N_23107,N_22202);
and U24548 (N_24548,N_23928,N_23994);
nor U24549 (N_24549,N_22001,N_23091);
nor U24550 (N_24550,N_22842,N_23095);
or U24551 (N_24551,N_23786,N_23266);
xor U24552 (N_24552,N_23223,N_23443);
nand U24553 (N_24553,N_22274,N_22843);
xor U24554 (N_24554,N_23038,N_22030);
xnor U24555 (N_24555,N_22515,N_23955);
xor U24556 (N_24556,N_23895,N_23859);
and U24557 (N_24557,N_23387,N_22136);
xnor U24558 (N_24558,N_22442,N_23748);
or U24559 (N_24559,N_23433,N_22485);
xor U24560 (N_24560,N_22122,N_23651);
nor U24561 (N_24561,N_22628,N_22682);
nor U24562 (N_24562,N_23516,N_23404);
or U24563 (N_24563,N_23021,N_23511);
nand U24564 (N_24564,N_22465,N_22831);
or U24565 (N_24565,N_23823,N_23745);
and U24566 (N_24566,N_23534,N_23360);
or U24567 (N_24567,N_22524,N_23577);
nor U24568 (N_24568,N_23826,N_22112);
nand U24569 (N_24569,N_23509,N_23954);
or U24570 (N_24570,N_22905,N_22056);
xnor U24571 (N_24571,N_22023,N_22100);
nand U24572 (N_24572,N_23146,N_23629);
xnor U24573 (N_24573,N_23250,N_23867);
and U24574 (N_24574,N_23567,N_22119);
xnor U24575 (N_24575,N_23562,N_22576);
nand U24576 (N_24576,N_22452,N_23756);
xnor U24577 (N_24577,N_23139,N_22103);
xnor U24578 (N_24578,N_23344,N_23912);
xor U24579 (N_24579,N_22631,N_23949);
xnor U24580 (N_24580,N_22925,N_22068);
nor U24581 (N_24581,N_23084,N_23115);
xor U24582 (N_24582,N_22161,N_22354);
and U24583 (N_24583,N_22022,N_23351);
or U24584 (N_24584,N_22475,N_23402);
nor U24585 (N_24585,N_22330,N_22419);
nand U24586 (N_24586,N_23644,N_22790);
or U24587 (N_24587,N_22548,N_23999);
nor U24588 (N_24588,N_22317,N_23214);
and U24589 (N_24589,N_23714,N_23390);
nand U24590 (N_24590,N_22319,N_23662);
or U24591 (N_24591,N_23114,N_22642);
xnor U24592 (N_24592,N_23010,N_23570);
and U24593 (N_24593,N_23338,N_23423);
or U24594 (N_24594,N_23965,N_23281);
nor U24595 (N_24595,N_22289,N_22221);
xor U24596 (N_24596,N_22701,N_22360);
xnor U24597 (N_24597,N_23853,N_22629);
nor U24598 (N_24598,N_23938,N_22564);
and U24599 (N_24599,N_22138,N_23888);
and U24600 (N_24600,N_23100,N_23005);
nor U24601 (N_24601,N_23340,N_22596);
nand U24602 (N_24602,N_23723,N_22183);
xnor U24603 (N_24603,N_23319,N_22930);
or U24604 (N_24604,N_22916,N_22203);
or U24605 (N_24605,N_22310,N_23395);
nor U24606 (N_24606,N_23325,N_22099);
nand U24607 (N_24607,N_23960,N_22276);
or U24608 (N_24608,N_23459,N_22804);
nand U24609 (N_24609,N_23675,N_22551);
xnor U24610 (N_24610,N_23816,N_23117);
or U24611 (N_24611,N_23546,N_22923);
nor U24612 (N_24612,N_22974,N_23697);
nand U24613 (N_24613,N_22996,N_23539);
and U24614 (N_24614,N_22984,N_22338);
and U24615 (N_24615,N_23674,N_22238);
and U24616 (N_24616,N_22726,N_22722);
or U24617 (N_24617,N_23772,N_22316);
nand U24618 (N_24618,N_23221,N_23969);
nor U24619 (N_24619,N_22196,N_22420);
xor U24620 (N_24620,N_23027,N_23073);
nor U24621 (N_24621,N_23127,N_22931);
or U24622 (N_24622,N_22692,N_23995);
nor U24623 (N_24623,N_22482,N_23719);
xor U24624 (N_24624,N_23210,N_23309);
nor U24625 (N_24625,N_22585,N_22546);
nand U24626 (N_24626,N_22514,N_22280);
or U24627 (N_24627,N_22259,N_23185);
xnor U24628 (N_24628,N_22904,N_22882);
or U24629 (N_24629,N_22394,N_23846);
nand U24630 (N_24630,N_23359,N_23646);
or U24631 (N_24631,N_22858,N_22729);
and U24632 (N_24632,N_22414,N_22875);
nor U24633 (N_24633,N_23861,N_23386);
nor U24634 (N_24634,N_23449,N_23497);
and U24635 (N_24635,N_23794,N_23735);
nand U24636 (N_24636,N_22665,N_22815);
or U24637 (N_24637,N_23852,N_23920);
nor U24638 (N_24638,N_22378,N_23383);
nand U24639 (N_24639,N_22246,N_23974);
nand U24640 (N_24640,N_22616,N_23398);
nand U24641 (N_24641,N_23759,N_23558);
and U24642 (N_24642,N_22358,N_22786);
nor U24643 (N_24643,N_23355,N_22437);
or U24644 (N_24644,N_22093,N_23176);
nand U24645 (N_24645,N_22840,N_23729);
nor U24646 (N_24646,N_22910,N_23352);
xor U24647 (N_24647,N_23054,N_23409);
nor U24648 (N_24648,N_22733,N_23504);
or U24649 (N_24649,N_23519,N_22461);
nor U24650 (N_24650,N_23258,N_23105);
and U24651 (N_24651,N_23700,N_23212);
or U24652 (N_24652,N_22448,N_23452);
xor U24653 (N_24653,N_22237,N_23311);
and U24654 (N_24654,N_22052,N_23328);
or U24655 (N_24655,N_23374,N_23494);
nor U24656 (N_24656,N_23140,N_23123);
or U24657 (N_24657,N_23156,N_22721);
xnor U24658 (N_24658,N_23657,N_23413);
and U24659 (N_24659,N_22117,N_22435);
nor U24660 (N_24660,N_22741,N_23839);
or U24661 (N_24661,N_23917,N_22973);
xnor U24662 (N_24662,N_22653,N_22346);
or U24663 (N_24663,N_22839,N_22680);
or U24664 (N_24664,N_22874,N_23229);
xor U24665 (N_24665,N_23133,N_22444);
xor U24666 (N_24666,N_23172,N_22814);
nor U24667 (N_24667,N_23269,N_23420);
nand U24668 (N_24668,N_22605,N_23468);
or U24669 (N_24669,N_22567,N_22226);
xnor U24670 (N_24670,N_22497,N_22156);
xnor U24671 (N_24671,N_22353,N_23106);
or U24672 (N_24672,N_23544,N_22809);
or U24673 (N_24673,N_22649,N_22820);
nor U24674 (N_24674,N_22805,N_22456);
and U24675 (N_24675,N_22940,N_23728);
xnor U24676 (N_24676,N_23668,N_23663);
nand U24677 (N_24677,N_22003,N_22919);
xnor U24678 (N_24678,N_22793,N_22801);
nor U24679 (N_24679,N_22069,N_22817);
or U24680 (N_24680,N_22489,N_23421);
or U24681 (N_24681,N_23684,N_22058);
and U24682 (N_24682,N_23579,N_23947);
nand U24683 (N_24683,N_23130,N_23392);
nor U24684 (N_24684,N_22580,N_23160);
nand U24685 (N_24685,N_23827,N_22010);
nor U24686 (N_24686,N_22451,N_23055);
nand U24687 (N_24687,N_22764,N_22987);
nor U24688 (N_24688,N_22545,N_23103);
and U24689 (N_24689,N_22519,N_22929);
or U24690 (N_24690,N_22672,N_22053);
nand U24691 (N_24691,N_22337,N_22092);
and U24692 (N_24692,N_23734,N_22396);
or U24693 (N_24693,N_22428,N_22927);
xor U24694 (N_24694,N_23358,N_22050);
nor U24695 (N_24695,N_23015,N_23924);
nand U24696 (N_24696,N_23132,N_22915);
nand U24697 (N_24697,N_22087,N_23342);
nand U24698 (N_24698,N_23505,N_22508);
nor U24699 (N_24699,N_23239,N_22794);
xor U24700 (N_24700,N_23872,N_22939);
nand U24701 (N_24701,N_22570,N_22897);
nand U24702 (N_24702,N_22951,N_23597);
and U24703 (N_24703,N_23235,N_23583);
and U24704 (N_24704,N_22888,N_23820);
nand U24705 (N_24705,N_22074,N_22445);
or U24706 (N_24706,N_22690,N_22792);
xor U24707 (N_24707,N_23343,N_22398);
and U24708 (N_24708,N_22841,N_23775);
nand U24709 (N_24709,N_23699,N_22095);
or U24710 (N_24710,N_23537,N_23341);
nand U24711 (N_24711,N_23771,N_23002);
and U24712 (N_24712,N_23941,N_23806);
xor U24713 (N_24713,N_22009,N_23889);
nand U24714 (N_24714,N_22361,N_23291);
or U24715 (N_24715,N_22860,N_23880);
and U24716 (N_24716,N_23077,N_23437);
and U24717 (N_24717,N_23959,N_23549);
nand U24718 (N_24718,N_23295,N_23346);
and U24719 (N_24719,N_22679,N_23890);
nand U24720 (N_24720,N_23203,N_23779);
xnor U24721 (N_24721,N_23052,N_23403);
xor U24722 (N_24722,N_22251,N_22065);
xnor U24723 (N_24723,N_23940,N_23877);
or U24724 (N_24724,N_22055,N_22614);
nand U24725 (N_24725,N_23992,N_23921);
and U24726 (N_24726,N_23495,N_22788);
nor U24727 (N_24727,N_22081,N_22436);
xor U24728 (N_24728,N_22728,N_22163);
and U24729 (N_24729,N_22818,N_23356);
nor U24730 (N_24730,N_23198,N_23249);
xnor U24731 (N_24731,N_22718,N_22737);
xnor U24732 (N_24732,N_23733,N_23939);
nand U24733 (N_24733,N_22134,N_23632);
or U24734 (N_24734,N_22970,N_22912);
xnor U24735 (N_24735,N_22696,N_22862);
and U24736 (N_24736,N_22604,N_22571);
nand U24737 (N_24737,N_23837,N_22918);
xor U24738 (N_24738,N_23717,N_22771);
or U24739 (N_24739,N_22291,N_23382);
nor U24740 (N_24740,N_22415,N_23934);
xnor U24741 (N_24741,N_23659,N_22024);
nand U24742 (N_24742,N_22260,N_22569);
and U24743 (N_24743,N_23274,N_22347);
nor U24744 (N_24744,N_22080,N_22261);
xnor U24745 (N_24745,N_22411,N_23640);
nand U24746 (N_24746,N_23427,N_22397);
xnor U24747 (N_24747,N_23952,N_23408);
nand U24748 (N_24748,N_23197,N_23018);
nor U24749 (N_24749,N_22133,N_23238);
nor U24750 (N_24750,N_22980,N_22538);
and U24751 (N_24751,N_23866,N_22950);
and U24752 (N_24752,N_22165,N_22028);
nand U24753 (N_24753,N_23978,N_22141);
or U24754 (N_24754,N_23279,N_23540);
nor U24755 (N_24755,N_23884,N_23071);
nand U24756 (N_24756,N_23230,N_23486);
nor U24757 (N_24757,N_23075,N_23943);
or U24758 (N_24758,N_22767,N_22463);
nand U24759 (N_24759,N_22634,N_22555);
nand U24760 (N_24760,N_23871,N_22230);
and U24761 (N_24761,N_22477,N_23986);
nand U24762 (N_24762,N_22813,N_23367);
or U24763 (N_24763,N_23283,N_22655);
and U24764 (N_24764,N_23455,N_23578);
nand U24765 (N_24765,N_23603,N_23970);
nand U24766 (N_24766,N_23280,N_22137);
xor U24767 (N_24767,N_23650,N_22227);
nor U24768 (N_24768,N_22534,N_23515);
xor U24769 (N_24769,N_23982,N_23432);
and U24770 (N_24770,N_23034,N_22169);
or U24771 (N_24771,N_22699,N_22766);
nor U24772 (N_24772,N_22336,N_22531);
or U24773 (N_24773,N_23079,N_22421);
or U24774 (N_24774,N_23618,N_23187);
nor U24775 (N_24775,N_23935,N_23953);
nor U24776 (N_24776,N_23560,N_23513);
xor U24777 (N_24777,N_22094,N_22086);
xor U24778 (N_24778,N_23811,N_22782);
or U24779 (N_24779,N_23556,N_23072);
and U24780 (N_24780,N_23372,N_23143);
nand U24781 (N_24781,N_23439,N_22031);
nand U24782 (N_24782,N_23137,N_23666);
xnor U24783 (N_24783,N_22731,N_22934);
nor U24784 (N_24784,N_22290,N_23388);
and U24785 (N_24785,N_23378,N_23844);
xnor U24786 (N_24786,N_22754,N_22872);
or U24787 (N_24787,N_23948,N_22877);
nand U24788 (N_24788,N_22697,N_22938);
and U24789 (N_24789,N_23417,N_23345);
and U24790 (N_24790,N_23754,N_22392);
nor U24791 (N_24791,N_22739,N_23747);
nor U24792 (N_24792,N_22363,N_23993);
nand U24793 (N_24793,N_23812,N_22894);
nand U24794 (N_24794,N_23783,N_23694);
or U24795 (N_24795,N_22377,N_22626);
nor U24796 (N_24796,N_23217,N_23780);
and U24797 (N_24797,N_23039,N_23118);
and U24798 (N_24798,N_23502,N_22088);
xor U24799 (N_24799,N_22828,N_23613);
and U24800 (N_24800,N_23188,N_22286);
xnor U24801 (N_24801,N_22615,N_22859);
or U24802 (N_24802,N_23394,N_23730);
nor U24803 (N_24803,N_22991,N_22666);
xor U24804 (N_24804,N_23211,N_23482);
xnor U24805 (N_24805,N_22239,N_22573);
nand U24806 (N_24806,N_22229,N_23373);
nand U24807 (N_24807,N_22506,N_22480);
nand U24808 (N_24808,N_22333,N_22314);
and U24809 (N_24809,N_23685,N_22107);
nand U24810 (N_24810,N_23189,N_23688);
and U24811 (N_24811,N_23902,N_23703);
or U24812 (N_24812,N_22218,N_22990);
and U24813 (N_24813,N_23758,N_22142);
or U24814 (N_24814,N_23951,N_22307);
xnor U24815 (N_24815,N_23436,N_23180);
xor U24816 (N_24816,N_22258,N_22303);
nor U24817 (N_24817,N_23401,N_22296);
nand U24818 (N_24818,N_22675,N_23184);
xor U24819 (N_24819,N_23063,N_22139);
or U24820 (N_24820,N_22756,N_22561);
xnor U24821 (N_24821,N_23454,N_23726);
nor U24822 (N_24822,N_23087,N_22740);
xnor U24823 (N_24823,N_22019,N_23161);
xnor U24824 (N_24824,N_22889,N_23795);
xnor U24825 (N_24825,N_23285,N_23996);
nand U24826 (N_24826,N_22800,N_23892);
nand U24827 (N_24827,N_22211,N_23874);
nor U24828 (N_24828,N_22795,N_23226);
nand U24829 (N_24829,N_23252,N_22892);
xor U24830 (N_24830,N_22825,N_22410);
xor U24831 (N_24831,N_23633,N_23220);
xor U24832 (N_24832,N_23968,N_23990);
or U24833 (N_24833,N_22446,N_22061);
or U24834 (N_24834,N_23587,N_23991);
nor U24835 (N_24835,N_22450,N_22760);
and U24836 (N_24836,N_22273,N_22547);
or U24837 (N_24837,N_23232,N_23257);
or U24838 (N_24838,N_22557,N_22335);
xnor U24839 (N_24839,N_23007,N_22097);
nor U24840 (N_24840,N_23536,N_23237);
nor U24841 (N_24841,N_22305,N_23333);
or U24842 (N_24842,N_22774,N_23014);
nand U24843 (N_24843,N_23882,N_22057);
nand U24844 (N_24844,N_22220,N_22674);
and U24845 (N_24845,N_23933,N_23069);
nor U24846 (N_24846,N_22129,N_22884);
and U24847 (N_24847,N_22971,N_23649);
xnor U24848 (N_24848,N_23813,N_22131);
and U24849 (N_24849,N_23636,N_22710);
and U24850 (N_24850,N_23973,N_23078);
and U24851 (N_24851,N_22049,N_22399);
nand U24852 (N_24852,N_23430,N_23322);
nand U24853 (N_24853,N_23604,N_23036);
and U24854 (N_24854,N_22956,N_23631);
nand U24855 (N_24855,N_22694,N_22593);
or U24856 (N_24856,N_22469,N_23945);
or U24857 (N_24857,N_23642,N_23551);
or U24858 (N_24858,N_22167,N_22581);
or U24859 (N_24859,N_22583,N_22105);
or U24860 (N_24860,N_22989,N_23368);
xnor U24861 (N_24861,N_23607,N_22853);
xnor U24862 (N_24862,N_22849,N_23275);
nand U24863 (N_24863,N_22110,N_22949);
nor U24864 (N_24864,N_22412,N_23444);
xnor U24865 (N_24865,N_22179,N_23692);
nand U24866 (N_24866,N_22819,N_22153);
nor U24867 (N_24867,N_23985,N_23293);
nor U24868 (N_24868,N_23542,N_22054);
and U24869 (N_24869,N_23233,N_22404);
nand U24870 (N_24870,N_23170,N_22375);
or U24871 (N_24871,N_22189,N_22006);
xor U24872 (N_24872,N_23326,N_23842);
nor U24873 (N_24873,N_23522,N_23983);
xnor U24874 (N_24874,N_22611,N_22799);
or U24875 (N_24875,N_22027,N_23744);
and U24876 (N_24876,N_22908,N_22903);
or U24877 (N_24877,N_23061,N_23658);
and U24878 (N_24878,N_22343,N_22454);
xnor U24879 (N_24879,N_23521,N_23339);
xor U24880 (N_24880,N_22367,N_23641);
nand U24881 (N_24881,N_22541,N_22797);
and U24882 (N_24882,N_22683,N_22171);
nand U24883 (N_24883,N_23150,N_23998);
and U24884 (N_24884,N_23561,N_22780);
xor U24885 (N_24885,N_22484,N_23569);
and U24886 (N_24886,N_22504,N_23460);
nand U24887 (N_24887,N_22926,N_22533);
xor U24888 (N_24888,N_22045,N_23765);
or U24889 (N_24889,N_22505,N_23590);
nand U24890 (N_24890,N_23179,N_22090);
nor U24891 (N_24891,N_23248,N_23228);
nand U24892 (N_24892,N_22483,N_23415);
and U24893 (N_24893,N_22309,N_22373);
and U24894 (N_24894,N_22151,N_23422);
xor U24895 (N_24895,N_23476,N_23480);
or U24896 (N_24896,N_23264,N_22269);
and U24897 (N_24897,N_23517,N_22214);
nand U24898 (N_24898,N_22865,N_22181);
nor U24899 (N_24899,N_22511,N_22885);
xnor U24900 (N_24900,N_23919,N_22219);
nor U24901 (N_24901,N_22706,N_23391);
and U24902 (N_24902,N_23738,N_22244);
nand U24903 (N_24903,N_22447,N_22832);
or U24904 (N_24904,N_22453,N_23752);
xnor U24905 (N_24905,N_23743,N_22321);
nand U24906 (N_24906,N_23790,N_22781);
nor U24907 (N_24907,N_22758,N_22295);
and U24908 (N_24908,N_23362,N_23798);
and U24909 (N_24909,N_23006,N_22556);
xnor U24910 (N_24910,N_22186,N_23109);
nor U24911 (N_24911,N_23623,N_22041);
nor U24912 (N_24912,N_22686,N_23893);
and U24913 (N_24913,N_23012,N_22464);
nor U24914 (N_24914,N_23202,N_22959);
or U24915 (N_24915,N_23350,N_23000);
nand U24916 (N_24916,N_22677,N_23731);
xnor U24917 (N_24917,N_23831,N_23929);
xnor U24918 (N_24918,N_22178,N_23086);
nand U24919 (N_24919,N_22759,N_23213);
nand U24920 (N_24920,N_22529,N_22986);
or U24921 (N_24921,N_22152,N_22190);
and U24922 (N_24922,N_22735,N_23164);
xor U24923 (N_24923,N_22232,N_22958);
and U24924 (N_24924,N_22172,N_23001);
nor U24925 (N_24925,N_22007,N_23254);
nor U24926 (N_24926,N_23243,N_22773);
nor U24927 (N_24927,N_23263,N_22005);
and U24928 (N_24928,N_22968,N_22743);
and U24929 (N_24929,N_22707,N_22159);
and U24930 (N_24930,N_22102,N_22725);
or U24931 (N_24931,N_23716,N_23448);
xnor U24932 (N_24932,N_23664,N_23710);
nor U24933 (N_24933,N_22676,N_23718);
nor U24934 (N_24934,N_22365,N_23523);
and U24935 (N_24935,N_22791,N_22350);
and U24936 (N_24936,N_22040,N_23906);
xnor U24937 (N_24937,N_23024,N_23310);
nand U24938 (N_24938,N_22948,N_23961);
and U24939 (N_24939,N_23764,N_22288);
nand U24940 (N_24940,N_23489,N_23840);
nor U24941 (N_24941,N_22870,N_23261);
nor U24942 (N_24942,N_22867,N_22717);
or U24943 (N_24943,N_22282,N_22523);
xnor U24944 (N_24944,N_23611,N_22816);
or U24945 (N_24945,N_22661,N_23013);
nand U24946 (N_24946,N_22880,N_22618);
xor U24947 (N_24947,N_22763,N_23153);
and U24948 (N_24948,N_23606,N_22104);
xnor U24949 (N_24949,N_23121,N_22013);
and U24950 (N_24950,N_23173,N_22298);
xnor U24951 (N_24951,N_23191,N_23810);
xor U24952 (N_24952,N_22180,N_23913);
xor U24953 (N_24953,N_23972,N_22600);
or U24954 (N_24954,N_23778,N_23135);
nand U24955 (N_24955,N_22562,N_22654);
nor U24956 (N_24956,N_23416,N_23112);
or U24957 (N_24957,N_23163,N_23200);
nand U24958 (N_24958,N_23677,N_22993);
nand U24959 (N_24959,N_23288,N_22362);
xor U24960 (N_24960,N_23076,N_22664);
nand U24961 (N_24961,N_23660,N_23740);
xnor U24962 (N_24962,N_22059,N_23407);
xor U24963 (N_24963,N_22016,N_23818);
or U24964 (N_24964,N_22621,N_23083);
and U24965 (N_24965,N_22757,N_22994);
nand U24966 (N_24966,N_22357,N_22510);
and U24967 (N_24967,N_22967,N_23976);
xor U24968 (N_24968,N_23615,N_23207);
nand U24969 (N_24969,N_23009,N_22348);
and U24970 (N_24970,N_23025,N_22315);
xor U24971 (N_24971,N_22847,N_23348);
or U24972 (N_24972,N_23047,N_23463);
or U24973 (N_24973,N_22612,N_23246);
or U24974 (N_24974,N_23464,N_22983);
and U24975 (N_24975,N_23910,N_23689);
or U24976 (N_24976,N_22342,N_22494);
or U24977 (N_24977,N_22292,N_22368);
and U24978 (N_24978,N_23638,N_23440);
nand U24979 (N_24979,N_22900,N_22029);
nand U24980 (N_24980,N_22032,N_22516);
and U24981 (N_24981,N_22535,N_22294);
and U24982 (N_24982,N_22588,N_23681);
xor U24983 (N_24983,N_22822,N_22772);
xnor U24984 (N_24984,N_23977,N_23102);
or U24985 (N_24985,N_23653,N_22458);
nor U24986 (N_24986,N_22474,N_23930);
and U24987 (N_24987,N_22632,N_22574);
and U24988 (N_24988,N_22067,N_23736);
nand U24989 (N_24989,N_23601,N_23234);
xor U24990 (N_24990,N_22857,N_23305);
nand U24991 (N_24991,N_23033,N_23931);
nor U24992 (N_24992,N_23830,N_23446);
or U24993 (N_24993,N_23802,N_23799);
and U24994 (N_24994,N_23514,N_23897);
xnor U24995 (N_24995,N_22532,N_22388);
xnor U24996 (N_24996,N_23702,N_23774);
and U24997 (N_24997,N_23183,N_22668);
or U24998 (N_24998,N_22965,N_23385);
nand U24999 (N_24999,N_22651,N_22443);
or U25000 (N_25000,N_22515,N_22908);
and U25001 (N_25001,N_23862,N_22555);
or U25002 (N_25002,N_23319,N_22722);
and U25003 (N_25003,N_23389,N_23322);
and U25004 (N_25004,N_23468,N_22410);
and U25005 (N_25005,N_23671,N_22518);
xor U25006 (N_25006,N_22441,N_22371);
nor U25007 (N_25007,N_22786,N_23315);
and U25008 (N_25008,N_23403,N_22933);
or U25009 (N_25009,N_22574,N_23863);
and U25010 (N_25010,N_22330,N_23307);
or U25011 (N_25011,N_22748,N_22876);
nor U25012 (N_25012,N_22911,N_23736);
and U25013 (N_25013,N_23889,N_22835);
nor U25014 (N_25014,N_23725,N_22628);
and U25015 (N_25015,N_22678,N_23260);
xnor U25016 (N_25016,N_23768,N_23617);
and U25017 (N_25017,N_22530,N_22207);
nor U25018 (N_25018,N_22577,N_22748);
and U25019 (N_25019,N_22064,N_22481);
and U25020 (N_25020,N_23418,N_22507);
nor U25021 (N_25021,N_22541,N_22885);
nand U25022 (N_25022,N_22066,N_23295);
and U25023 (N_25023,N_22225,N_23419);
nor U25024 (N_25024,N_22292,N_23204);
xor U25025 (N_25025,N_22265,N_22492);
xor U25026 (N_25026,N_23207,N_22718);
and U25027 (N_25027,N_22366,N_23209);
nor U25028 (N_25028,N_23514,N_23430);
nand U25029 (N_25029,N_22770,N_23571);
nand U25030 (N_25030,N_22211,N_23218);
xor U25031 (N_25031,N_23274,N_22143);
or U25032 (N_25032,N_22322,N_23252);
nor U25033 (N_25033,N_22482,N_23766);
or U25034 (N_25034,N_22622,N_22663);
xnor U25035 (N_25035,N_22023,N_23811);
and U25036 (N_25036,N_22138,N_23868);
or U25037 (N_25037,N_22524,N_22177);
xor U25038 (N_25038,N_22120,N_23783);
xor U25039 (N_25039,N_22769,N_23403);
or U25040 (N_25040,N_22474,N_23926);
xor U25041 (N_25041,N_23342,N_22152);
or U25042 (N_25042,N_23737,N_23539);
xnor U25043 (N_25043,N_22499,N_22805);
and U25044 (N_25044,N_22443,N_23599);
xor U25045 (N_25045,N_22503,N_22258);
nor U25046 (N_25046,N_22545,N_22744);
or U25047 (N_25047,N_23728,N_23843);
and U25048 (N_25048,N_22675,N_23042);
nor U25049 (N_25049,N_22180,N_22667);
and U25050 (N_25050,N_23226,N_23090);
nor U25051 (N_25051,N_23232,N_23209);
xnor U25052 (N_25052,N_22284,N_23717);
nand U25053 (N_25053,N_22753,N_23508);
and U25054 (N_25054,N_22975,N_22244);
or U25055 (N_25055,N_23284,N_23061);
nor U25056 (N_25056,N_22085,N_22027);
xnor U25057 (N_25057,N_23468,N_22617);
and U25058 (N_25058,N_23190,N_23787);
xnor U25059 (N_25059,N_22758,N_22214);
or U25060 (N_25060,N_22828,N_22895);
nor U25061 (N_25061,N_23687,N_23125);
nor U25062 (N_25062,N_22725,N_22688);
nand U25063 (N_25063,N_23305,N_23199);
nor U25064 (N_25064,N_23205,N_23350);
xor U25065 (N_25065,N_22875,N_23266);
or U25066 (N_25066,N_22014,N_22388);
xor U25067 (N_25067,N_22208,N_22214);
nor U25068 (N_25068,N_22995,N_23022);
nor U25069 (N_25069,N_22628,N_22615);
nor U25070 (N_25070,N_23706,N_22528);
nor U25071 (N_25071,N_23968,N_22207);
nand U25072 (N_25072,N_22404,N_22172);
nand U25073 (N_25073,N_22805,N_22075);
xnor U25074 (N_25074,N_23061,N_22783);
and U25075 (N_25075,N_22226,N_22589);
nor U25076 (N_25076,N_23662,N_22629);
or U25077 (N_25077,N_22871,N_23719);
xnor U25078 (N_25078,N_23977,N_22726);
nand U25079 (N_25079,N_23303,N_22286);
nor U25080 (N_25080,N_22526,N_23955);
and U25081 (N_25081,N_22501,N_22118);
nand U25082 (N_25082,N_22816,N_22046);
and U25083 (N_25083,N_23810,N_23566);
nor U25084 (N_25084,N_22836,N_23953);
nor U25085 (N_25085,N_22942,N_23459);
xnor U25086 (N_25086,N_23702,N_22331);
and U25087 (N_25087,N_22886,N_23555);
and U25088 (N_25088,N_22632,N_23705);
or U25089 (N_25089,N_23244,N_23233);
and U25090 (N_25090,N_22782,N_23896);
nor U25091 (N_25091,N_23868,N_22539);
nand U25092 (N_25092,N_23195,N_22958);
nor U25093 (N_25093,N_22116,N_23564);
nor U25094 (N_25094,N_23664,N_23466);
or U25095 (N_25095,N_23562,N_22793);
xor U25096 (N_25096,N_23046,N_23686);
nor U25097 (N_25097,N_22675,N_23821);
xor U25098 (N_25098,N_23652,N_22220);
and U25099 (N_25099,N_23529,N_22988);
nand U25100 (N_25100,N_23042,N_22319);
and U25101 (N_25101,N_23160,N_23700);
nor U25102 (N_25102,N_22528,N_23730);
nand U25103 (N_25103,N_23297,N_22850);
or U25104 (N_25104,N_22326,N_22549);
nor U25105 (N_25105,N_23289,N_23660);
nand U25106 (N_25106,N_22071,N_22229);
nor U25107 (N_25107,N_22828,N_22207);
nand U25108 (N_25108,N_22571,N_22758);
and U25109 (N_25109,N_22164,N_23439);
and U25110 (N_25110,N_23308,N_23325);
xor U25111 (N_25111,N_23990,N_22566);
or U25112 (N_25112,N_23457,N_22319);
nand U25113 (N_25113,N_23038,N_22824);
xnor U25114 (N_25114,N_22087,N_22512);
nand U25115 (N_25115,N_22355,N_23795);
nor U25116 (N_25116,N_23162,N_22596);
or U25117 (N_25117,N_22603,N_22946);
nand U25118 (N_25118,N_22449,N_23160);
nor U25119 (N_25119,N_23107,N_23610);
or U25120 (N_25120,N_23827,N_23905);
nor U25121 (N_25121,N_22609,N_22169);
nand U25122 (N_25122,N_23979,N_22269);
or U25123 (N_25123,N_22637,N_23639);
or U25124 (N_25124,N_23665,N_23315);
nand U25125 (N_25125,N_22676,N_22781);
nor U25126 (N_25126,N_23166,N_22493);
xnor U25127 (N_25127,N_23657,N_23629);
nand U25128 (N_25128,N_23036,N_22529);
nor U25129 (N_25129,N_22388,N_23485);
and U25130 (N_25130,N_22201,N_23691);
or U25131 (N_25131,N_22836,N_22304);
xnor U25132 (N_25132,N_23856,N_22053);
nor U25133 (N_25133,N_22072,N_22297);
nand U25134 (N_25134,N_22030,N_23313);
or U25135 (N_25135,N_22630,N_23223);
nor U25136 (N_25136,N_22286,N_22964);
or U25137 (N_25137,N_22810,N_22099);
xnor U25138 (N_25138,N_22144,N_23364);
nor U25139 (N_25139,N_23692,N_22422);
nor U25140 (N_25140,N_22277,N_22248);
and U25141 (N_25141,N_22128,N_22018);
nand U25142 (N_25142,N_23506,N_22921);
xnor U25143 (N_25143,N_22874,N_23380);
or U25144 (N_25144,N_22824,N_23466);
nand U25145 (N_25145,N_23546,N_23074);
and U25146 (N_25146,N_22248,N_23606);
and U25147 (N_25147,N_22934,N_22226);
or U25148 (N_25148,N_22986,N_22590);
xor U25149 (N_25149,N_22462,N_23381);
or U25150 (N_25150,N_23020,N_22014);
or U25151 (N_25151,N_22547,N_23689);
nor U25152 (N_25152,N_22662,N_22059);
and U25153 (N_25153,N_23824,N_23830);
and U25154 (N_25154,N_22319,N_22898);
nor U25155 (N_25155,N_23335,N_22982);
and U25156 (N_25156,N_22752,N_22623);
nor U25157 (N_25157,N_23732,N_23284);
or U25158 (N_25158,N_23797,N_22482);
nor U25159 (N_25159,N_22129,N_22329);
or U25160 (N_25160,N_22010,N_23218);
and U25161 (N_25161,N_22517,N_23067);
or U25162 (N_25162,N_22121,N_23919);
and U25163 (N_25163,N_22387,N_23768);
nor U25164 (N_25164,N_23861,N_22466);
and U25165 (N_25165,N_22455,N_22033);
xnor U25166 (N_25166,N_22140,N_23374);
nand U25167 (N_25167,N_23820,N_22814);
nand U25168 (N_25168,N_22721,N_23050);
and U25169 (N_25169,N_22969,N_23765);
xnor U25170 (N_25170,N_23015,N_22414);
and U25171 (N_25171,N_22790,N_22414);
xnor U25172 (N_25172,N_22460,N_22674);
and U25173 (N_25173,N_23762,N_22904);
and U25174 (N_25174,N_23297,N_23852);
and U25175 (N_25175,N_23152,N_23741);
nor U25176 (N_25176,N_22511,N_23595);
and U25177 (N_25177,N_22913,N_22588);
xor U25178 (N_25178,N_22870,N_22687);
xor U25179 (N_25179,N_22660,N_23463);
nor U25180 (N_25180,N_23078,N_22834);
and U25181 (N_25181,N_23034,N_23282);
nand U25182 (N_25182,N_22177,N_22539);
nand U25183 (N_25183,N_22400,N_22759);
nor U25184 (N_25184,N_23530,N_23187);
xor U25185 (N_25185,N_22669,N_23520);
or U25186 (N_25186,N_22578,N_23094);
nand U25187 (N_25187,N_23843,N_23172);
xor U25188 (N_25188,N_23465,N_23870);
xnor U25189 (N_25189,N_23260,N_23233);
xor U25190 (N_25190,N_23944,N_22517);
xnor U25191 (N_25191,N_23831,N_22804);
xor U25192 (N_25192,N_22295,N_23207);
or U25193 (N_25193,N_22146,N_22623);
nand U25194 (N_25194,N_22361,N_23713);
and U25195 (N_25195,N_22908,N_22213);
nand U25196 (N_25196,N_23462,N_23697);
nand U25197 (N_25197,N_23959,N_23416);
xnor U25198 (N_25198,N_22934,N_22445);
nor U25199 (N_25199,N_22661,N_23229);
and U25200 (N_25200,N_23819,N_22177);
nor U25201 (N_25201,N_22779,N_23699);
and U25202 (N_25202,N_23209,N_23936);
nor U25203 (N_25203,N_23235,N_23371);
or U25204 (N_25204,N_23180,N_22026);
and U25205 (N_25205,N_23553,N_22992);
nor U25206 (N_25206,N_22122,N_22045);
nand U25207 (N_25207,N_23981,N_22635);
or U25208 (N_25208,N_23928,N_23179);
nand U25209 (N_25209,N_22022,N_22676);
xor U25210 (N_25210,N_23206,N_22486);
nor U25211 (N_25211,N_22734,N_22602);
and U25212 (N_25212,N_23279,N_23889);
xnor U25213 (N_25213,N_23205,N_22920);
nor U25214 (N_25214,N_22887,N_22322);
nand U25215 (N_25215,N_23664,N_23039);
or U25216 (N_25216,N_23590,N_22790);
nor U25217 (N_25217,N_23231,N_23907);
or U25218 (N_25218,N_22890,N_23317);
xor U25219 (N_25219,N_23892,N_22332);
or U25220 (N_25220,N_23282,N_22284);
nor U25221 (N_25221,N_22605,N_23634);
or U25222 (N_25222,N_22826,N_23118);
nor U25223 (N_25223,N_23921,N_23805);
nand U25224 (N_25224,N_22914,N_22040);
xnor U25225 (N_25225,N_22947,N_22425);
nand U25226 (N_25226,N_22982,N_22112);
nand U25227 (N_25227,N_23571,N_23483);
and U25228 (N_25228,N_22523,N_23718);
nand U25229 (N_25229,N_22924,N_23328);
and U25230 (N_25230,N_23692,N_22438);
or U25231 (N_25231,N_23691,N_22801);
and U25232 (N_25232,N_23639,N_23081);
and U25233 (N_25233,N_22818,N_22873);
nand U25234 (N_25234,N_23170,N_22050);
or U25235 (N_25235,N_23336,N_22080);
nand U25236 (N_25236,N_22868,N_22770);
nand U25237 (N_25237,N_22570,N_23175);
nor U25238 (N_25238,N_22521,N_23267);
xnor U25239 (N_25239,N_22114,N_22646);
nand U25240 (N_25240,N_22595,N_22203);
or U25241 (N_25241,N_22703,N_23704);
or U25242 (N_25242,N_22859,N_22969);
xnor U25243 (N_25243,N_22576,N_22067);
and U25244 (N_25244,N_22773,N_22618);
or U25245 (N_25245,N_23814,N_22204);
nor U25246 (N_25246,N_22627,N_23576);
nor U25247 (N_25247,N_23164,N_22305);
or U25248 (N_25248,N_23666,N_22416);
nand U25249 (N_25249,N_22984,N_23968);
and U25250 (N_25250,N_22541,N_23208);
nand U25251 (N_25251,N_23691,N_22634);
nor U25252 (N_25252,N_23562,N_23662);
and U25253 (N_25253,N_23833,N_22113);
nand U25254 (N_25254,N_22845,N_22177);
xor U25255 (N_25255,N_23623,N_22306);
and U25256 (N_25256,N_23781,N_23291);
nor U25257 (N_25257,N_22933,N_22841);
nor U25258 (N_25258,N_23665,N_22362);
nand U25259 (N_25259,N_22532,N_23984);
nor U25260 (N_25260,N_22210,N_22639);
and U25261 (N_25261,N_22300,N_23065);
nor U25262 (N_25262,N_22314,N_22832);
nand U25263 (N_25263,N_22240,N_23532);
or U25264 (N_25264,N_22210,N_22972);
nand U25265 (N_25265,N_23793,N_23763);
nor U25266 (N_25266,N_22461,N_22900);
nor U25267 (N_25267,N_23845,N_22737);
or U25268 (N_25268,N_22368,N_23570);
xor U25269 (N_25269,N_23334,N_22397);
or U25270 (N_25270,N_23461,N_22176);
and U25271 (N_25271,N_23330,N_23313);
nor U25272 (N_25272,N_22310,N_23824);
xnor U25273 (N_25273,N_22268,N_22182);
nand U25274 (N_25274,N_23556,N_23980);
nor U25275 (N_25275,N_22539,N_22570);
xnor U25276 (N_25276,N_22451,N_23856);
nor U25277 (N_25277,N_22189,N_23266);
nand U25278 (N_25278,N_23296,N_22063);
nor U25279 (N_25279,N_23806,N_22993);
or U25280 (N_25280,N_22021,N_22257);
and U25281 (N_25281,N_22033,N_22180);
xnor U25282 (N_25282,N_22865,N_22595);
and U25283 (N_25283,N_23507,N_23653);
and U25284 (N_25284,N_23205,N_23315);
or U25285 (N_25285,N_23605,N_22376);
or U25286 (N_25286,N_23945,N_22676);
and U25287 (N_25287,N_22974,N_23488);
nand U25288 (N_25288,N_23149,N_23728);
and U25289 (N_25289,N_22085,N_23272);
nand U25290 (N_25290,N_22274,N_23280);
and U25291 (N_25291,N_23416,N_23949);
and U25292 (N_25292,N_22300,N_23962);
nand U25293 (N_25293,N_22654,N_23658);
nor U25294 (N_25294,N_22184,N_22836);
nor U25295 (N_25295,N_22777,N_23832);
or U25296 (N_25296,N_22768,N_23493);
and U25297 (N_25297,N_22926,N_22852);
nand U25298 (N_25298,N_23771,N_22242);
nand U25299 (N_25299,N_22791,N_22662);
xnor U25300 (N_25300,N_22438,N_22676);
or U25301 (N_25301,N_22472,N_22126);
or U25302 (N_25302,N_22893,N_23374);
or U25303 (N_25303,N_23637,N_22343);
nor U25304 (N_25304,N_22128,N_22852);
and U25305 (N_25305,N_23846,N_23718);
nand U25306 (N_25306,N_22555,N_23033);
nand U25307 (N_25307,N_22941,N_22509);
or U25308 (N_25308,N_23314,N_23817);
and U25309 (N_25309,N_23418,N_22072);
nand U25310 (N_25310,N_23917,N_23445);
or U25311 (N_25311,N_23478,N_23686);
xor U25312 (N_25312,N_22827,N_22563);
or U25313 (N_25313,N_23998,N_23282);
or U25314 (N_25314,N_22898,N_22444);
and U25315 (N_25315,N_22578,N_23902);
nand U25316 (N_25316,N_23179,N_23232);
and U25317 (N_25317,N_22219,N_23065);
and U25318 (N_25318,N_22930,N_23927);
nor U25319 (N_25319,N_23793,N_22660);
nand U25320 (N_25320,N_23906,N_22916);
or U25321 (N_25321,N_22086,N_23635);
or U25322 (N_25322,N_22347,N_22925);
nand U25323 (N_25323,N_23559,N_22300);
or U25324 (N_25324,N_23320,N_22347);
nand U25325 (N_25325,N_23377,N_22884);
or U25326 (N_25326,N_22056,N_22231);
xnor U25327 (N_25327,N_22619,N_23249);
and U25328 (N_25328,N_22846,N_22299);
and U25329 (N_25329,N_22253,N_22287);
or U25330 (N_25330,N_23642,N_22216);
nor U25331 (N_25331,N_22092,N_23118);
or U25332 (N_25332,N_23557,N_22895);
nor U25333 (N_25333,N_22496,N_22172);
and U25334 (N_25334,N_22551,N_23723);
nor U25335 (N_25335,N_22838,N_22830);
or U25336 (N_25336,N_23763,N_23830);
nor U25337 (N_25337,N_22347,N_22529);
and U25338 (N_25338,N_22324,N_23669);
xnor U25339 (N_25339,N_23644,N_23258);
or U25340 (N_25340,N_22556,N_23795);
nor U25341 (N_25341,N_23326,N_23570);
nand U25342 (N_25342,N_23627,N_23514);
nor U25343 (N_25343,N_22370,N_23097);
nor U25344 (N_25344,N_22726,N_22159);
or U25345 (N_25345,N_23914,N_23644);
nor U25346 (N_25346,N_23832,N_22788);
nor U25347 (N_25347,N_23535,N_22729);
or U25348 (N_25348,N_22198,N_23415);
or U25349 (N_25349,N_23876,N_22438);
and U25350 (N_25350,N_23299,N_23628);
nand U25351 (N_25351,N_22486,N_23699);
nor U25352 (N_25352,N_23721,N_22642);
nor U25353 (N_25353,N_23756,N_22604);
and U25354 (N_25354,N_23714,N_22144);
nand U25355 (N_25355,N_22179,N_22112);
and U25356 (N_25356,N_22057,N_23132);
and U25357 (N_25357,N_22180,N_22220);
xor U25358 (N_25358,N_23363,N_22175);
nor U25359 (N_25359,N_23545,N_22424);
nor U25360 (N_25360,N_22010,N_23478);
nor U25361 (N_25361,N_22375,N_23071);
or U25362 (N_25362,N_22500,N_22683);
xor U25363 (N_25363,N_22559,N_23759);
or U25364 (N_25364,N_23357,N_23083);
xnor U25365 (N_25365,N_22375,N_22448);
and U25366 (N_25366,N_22848,N_23991);
and U25367 (N_25367,N_23934,N_23775);
xor U25368 (N_25368,N_23232,N_23342);
nor U25369 (N_25369,N_22608,N_22070);
or U25370 (N_25370,N_23270,N_23152);
and U25371 (N_25371,N_23330,N_22451);
and U25372 (N_25372,N_22639,N_23035);
or U25373 (N_25373,N_22899,N_22634);
nor U25374 (N_25374,N_23481,N_23449);
nand U25375 (N_25375,N_23224,N_23884);
or U25376 (N_25376,N_23555,N_23694);
and U25377 (N_25377,N_23504,N_23061);
or U25378 (N_25378,N_22545,N_22434);
nand U25379 (N_25379,N_23874,N_22969);
nor U25380 (N_25380,N_22970,N_23998);
and U25381 (N_25381,N_22071,N_22546);
nor U25382 (N_25382,N_22785,N_22690);
xnor U25383 (N_25383,N_22677,N_22222);
nor U25384 (N_25384,N_22112,N_23935);
nor U25385 (N_25385,N_23926,N_22026);
nor U25386 (N_25386,N_22954,N_22646);
nor U25387 (N_25387,N_23002,N_22180);
nand U25388 (N_25388,N_23142,N_23234);
and U25389 (N_25389,N_22168,N_22766);
nor U25390 (N_25390,N_22657,N_22909);
nor U25391 (N_25391,N_22175,N_22567);
nor U25392 (N_25392,N_23002,N_22659);
nor U25393 (N_25393,N_22298,N_22762);
or U25394 (N_25394,N_23272,N_23394);
or U25395 (N_25395,N_23719,N_22847);
xnor U25396 (N_25396,N_22137,N_22778);
or U25397 (N_25397,N_22827,N_22070);
or U25398 (N_25398,N_22705,N_23507);
xor U25399 (N_25399,N_22621,N_23454);
or U25400 (N_25400,N_22101,N_23296);
nand U25401 (N_25401,N_23482,N_23957);
or U25402 (N_25402,N_23031,N_23085);
or U25403 (N_25403,N_22022,N_23387);
xor U25404 (N_25404,N_23458,N_22281);
xor U25405 (N_25405,N_22665,N_23362);
or U25406 (N_25406,N_22237,N_23204);
nor U25407 (N_25407,N_23613,N_23223);
or U25408 (N_25408,N_22281,N_22912);
and U25409 (N_25409,N_23419,N_22169);
nand U25410 (N_25410,N_22691,N_23177);
and U25411 (N_25411,N_23178,N_23526);
or U25412 (N_25412,N_22059,N_23931);
or U25413 (N_25413,N_23040,N_23378);
or U25414 (N_25414,N_23122,N_22170);
nand U25415 (N_25415,N_22167,N_23441);
and U25416 (N_25416,N_22874,N_22035);
or U25417 (N_25417,N_23711,N_22424);
or U25418 (N_25418,N_23412,N_23646);
xnor U25419 (N_25419,N_23816,N_23556);
xor U25420 (N_25420,N_23219,N_22544);
or U25421 (N_25421,N_23696,N_22014);
nand U25422 (N_25422,N_23821,N_23079);
and U25423 (N_25423,N_23701,N_23651);
and U25424 (N_25424,N_22942,N_23648);
xor U25425 (N_25425,N_23925,N_23567);
or U25426 (N_25426,N_22028,N_22502);
nor U25427 (N_25427,N_23596,N_23655);
nand U25428 (N_25428,N_23774,N_22009);
or U25429 (N_25429,N_23210,N_22718);
and U25430 (N_25430,N_23310,N_23454);
nor U25431 (N_25431,N_23956,N_23827);
nor U25432 (N_25432,N_23918,N_22585);
or U25433 (N_25433,N_23453,N_22722);
nor U25434 (N_25434,N_23299,N_23270);
xor U25435 (N_25435,N_22666,N_22372);
nand U25436 (N_25436,N_23126,N_22993);
and U25437 (N_25437,N_23488,N_22292);
and U25438 (N_25438,N_23584,N_22644);
or U25439 (N_25439,N_22325,N_22241);
nor U25440 (N_25440,N_23982,N_22002);
xnor U25441 (N_25441,N_22089,N_23637);
nand U25442 (N_25442,N_22918,N_22789);
xnor U25443 (N_25443,N_23478,N_23556);
nand U25444 (N_25444,N_22713,N_22040);
or U25445 (N_25445,N_22062,N_22139);
nor U25446 (N_25446,N_23577,N_23927);
nor U25447 (N_25447,N_23364,N_23640);
and U25448 (N_25448,N_23570,N_23130);
nor U25449 (N_25449,N_23480,N_22102);
xnor U25450 (N_25450,N_22702,N_23728);
xnor U25451 (N_25451,N_23059,N_23701);
or U25452 (N_25452,N_22421,N_22597);
or U25453 (N_25453,N_22726,N_23442);
or U25454 (N_25454,N_23013,N_23983);
or U25455 (N_25455,N_23954,N_23744);
or U25456 (N_25456,N_23542,N_22298);
or U25457 (N_25457,N_22114,N_22431);
and U25458 (N_25458,N_22016,N_22064);
xor U25459 (N_25459,N_23769,N_22434);
or U25460 (N_25460,N_22269,N_22755);
or U25461 (N_25461,N_23028,N_23010);
nor U25462 (N_25462,N_22636,N_23607);
or U25463 (N_25463,N_22271,N_23779);
or U25464 (N_25464,N_22560,N_22469);
xnor U25465 (N_25465,N_22967,N_23143);
nand U25466 (N_25466,N_23628,N_22346);
nor U25467 (N_25467,N_23642,N_22420);
or U25468 (N_25468,N_23580,N_22989);
xnor U25469 (N_25469,N_22693,N_23192);
xnor U25470 (N_25470,N_22661,N_23432);
nand U25471 (N_25471,N_23955,N_23864);
or U25472 (N_25472,N_23204,N_22548);
xor U25473 (N_25473,N_23201,N_23965);
nor U25474 (N_25474,N_23101,N_23610);
and U25475 (N_25475,N_23212,N_23240);
nor U25476 (N_25476,N_22111,N_22576);
xor U25477 (N_25477,N_23983,N_22597);
and U25478 (N_25478,N_22683,N_22467);
nor U25479 (N_25479,N_22206,N_23797);
xor U25480 (N_25480,N_22184,N_22577);
nand U25481 (N_25481,N_23862,N_22319);
and U25482 (N_25482,N_22095,N_23719);
or U25483 (N_25483,N_23740,N_23375);
xnor U25484 (N_25484,N_22251,N_22936);
and U25485 (N_25485,N_23641,N_22854);
xnor U25486 (N_25486,N_23215,N_23256);
nor U25487 (N_25487,N_22374,N_22717);
xor U25488 (N_25488,N_22914,N_22334);
and U25489 (N_25489,N_22456,N_23830);
nand U25490 (N_25490,N_23898,N_22898);
and U25491 (N_25491,N_22566,N_23573);
and U25492 (N_25492,N_22955,N_23176);
nor U25493 (N_25493,N_23089,N_23597);
and U25494 (N_25494,N_22022,N_22165);
and U25495 (N_25495,N_22090,N_22461);
and U25496 (N_25496,N_22734,N_23490);
nor U25497 (N_25497,N_22148,N_23449);
nand U25498 (N_25498,N_23641,N_22929);
xnor U25499 (N_25499,N_23524,N_22040);
or U25500 (N_25500,N_22086,N_23678);
xnor U25501 (N_25501,N_23973,N_23706);
nor U25502 (N_25502,N_23850,N_23704);
nor U25503 (N_25503,N_22650,N_22724);
xnor U25504 (N_25504,N_23909,N_23252);
nand U25505 (N_25505,N_23595,N_23715);
or U25506 (N_25506,N_22453,N_22474);
nor U25507 (N_25507,N_22221,N_23114);
xor U25508 (N_25508,N_22626,N_22372);
nor U25509 (N_25509,N_22019,N_22660);
nor U25510 (N_25510,N_22069,N_22480);
nor U25511 (N_25511,N_22948,N_23167);
or U25512 (N_25512,N_23660,N_23899);
or U25513 (N_25513,N_22860,N_22745);
nor U25514 (N_25514,N_23264,N_23948);
xor U25515 (N_25515,N_22222,N_22626);
nand U25516 (N_25516,N_23481,N_23255);
nor U25517 (N_25517,N_22949,N_23607);
nor U25518 (N_25518,N_22683,N_23570);
or U25519 (N_25519,N_22115,N_22366);
or U25520 (N_25520,N_22027,N_22491);
or U25521 (N_25521,N_23726,N_22517);
nand U25522 (N_25522,N_22968,N_23574);
and U25523 (N_25523,N_23486,N_23431);
xnor U25524 (N_25524,N_22473,N_22528);
or U25525 (N_25525,N_23580,N_23826);
and U25526 (N_25526,N_22766,N_23730);
or U25527 (N_25527,N_22156,N_22467);
xor U25528 (N_25528,N_23008,N_23155);
xnor U25529 (N_25529,N_23854,N_22090);
nand U25530 (N_25530,N_23563,N_22153);
nand U25531 (N_25531,N_23884,N_23387);
xor U25532 (N_25532,N_23758,N_23138);
xnor U25533 (N_25533,N_22094,N_23260);
nor U25534 (N_25534,N_23436,N_23718);
or U25535 (N_25535,N_22610,N_22858);
and U25536 (N_25536,N_22316,N_22551);
or U25537 (N_25537,N_22153,N_22474);
and U25538 (N_25538,N_23961,N_23163);
and U25539 (N_25539,N_23310,N_23381);
nor U25540 (N_25540,N_22637,N_22645);
nand U25541 (N_25541,N_23300,N_22346);
xor U25542 (N_25542,N_23326,N_23644);
xnor U25543 (N_25543,N_23166,N_22479);
xor U25544 (N_25544,N_22276,N_22501);
xnor U25545 (N_25545,N_22073,N_22299);
xor U25546 (N_25546,N_22897,N_22020);
or U25547 (N_25547,N_22107,N_22919);
and U25548 (N_25548,N_22472,N_22601);
and U25549 (N_25549,N_23337,N_22763);
and U25550 (N_25550,N_22750,N_22254);
and U25551 (N_25551,N_23151,N_22028);
nor U25552 (N_25552,N_23526,N_22340);
or U25553 (N_25553,N_22694,N_23547);
or U25554 (N_25554,N_23585,N_22709);
nor U25555 (N_25555,N_23158,N_22297);
xor U25556 (N_25556,N_23640,N_23670);
nand U25557 (N_25557,N_23302,N_22073);
or U25558 (N_25558,N_23110,N_22456);
nand U25559 (N_25559,N_22009,N_23293);
nor U25560 (N_25560,N_23590,N_23576);
nor U25561 (N_25561,N_23623,N_23971);
nand U25562 (N_25562,N_22592,N_22181);
or U25563 (N_25563,N_23672,N_23614);
nand U25564 (N_25564,N_23946,N_23896);
and U25565 (N_25565,N_22740,N_23733);
xor U25566 (N_25566,N_22464,N_23952);
and U25567 (N_25567,N_22089,N_22491);
nor U25568 (N_25568,N_23968,N_22209);
xnor U25569 (N_25569,N_22141,N_23107);
and U25570 (N_25570,N_22991,N_23567);
xor U25571 (N_25571,N_22296,N_22844);
nor U25572 (N_25572,N_23217,N_23867);
nand U25573 (N_25573,N_22732,N_23408);
or U25574 (N_25574,N_22989,N_23759);
and U25575 (N_25575,N_22456,N_22625);
and U25576 (N_25576,N_23404,N_23131);
and U25577 (N_25577,N_23073,N_22216);
nor U25578 (N_25578,N_22079,N_23438);
and U25579 (N_25579,N_23701,N_23103);
and U25580 (N_25580,N_23183,N_23989);
or U25581 (N_25581,N_23570,N_22497);
xor U25582 (N_25582,N_22380,N_23546);
nand U25583 (N_25583,N_23737,N_22038);
xnor U25584 (N_25584,N_23766,N_22007);
or U25585 (N_25585,N_22304,N_23530);
and U25586 (N_25586,N_22184,N_22927);
nand U25587 (N_25587,N_22185,N_22108);
and U25588 (N_25588,N_22805,N_23596);
or U25589 (N_25589,N_22305,N_22707);
xnor U25590 (N_25590,N_22653,N_22169);
and U25591 (N_25591,N_22639,N_23528);
xor U25592 (N_25592,N_23864,N_23131);
nand U25593 (N_25593,N_23029,N_23124);
and U25594 (N_25594,N_23490,N_22993);
or U25595 (N_25595,N_23791,N_23848);
and U25596 (N_25596,N_23237,N_23105);
and U25597 (N_25597,N_22451,N_23181);
xnor U25598 (N_25598,N_22281,N_23104);
xnor U25599 (N_25599,N_22096,N_23112);
xnor U25600 (N_25600,N_23380,N_23506);
or U25601 (N_25601,N_22892,N_22177);
or U25602 (N_25602,N_23119,N_23498);
xor U25603 (N_25603,N_23589,N_23370);
or U25604 (N_25604,N_23514,N_23093);
and U25605 (N_25605,N_23710,N_23181);
nor U25606 (N_25606,N_22108,N_22749);
and U25607 (N_25607,N_23019,N_23477);
or U25608 (N_25608,N_22945,N_22928);
xor U25609 (N_25609,N_22154,N_22408);
and U25610 (N_25610,N_22042,N_23095);
nand U25611 (N_25611,N_23920,N_23072);
nor U25612 (N_25612,N_23961,N_22683);
or U25613 (N_25613,N_23972,N_23045);
or U25614 (N_25614,N_22500,N_23766);
xnor U25615 (N_25615,N_22269,N_22587);
nand U25616 (N_25616,N_22767,N_22000);
nand U25617 (N_25617,N_22965,N_22723);
or U25618 (N_25618,N_23196,N_22450);
or U25619 (N_25619,N_23770,N_23618);
xnor U25620 (N_25620,N_22816,N_22557);
nor U25621 (N_25621,N_22723,N_22053);
and U25622 (N_25622,N_23558,N_22448);
or U25623 (N_25623,N_23460,N_23120);
and U25624 (N_25624,N_22424,N_22647);
or U25625 (N_25625,N_22867,N_22157);
xor U25626 (N_25626,N_22775,N_23245);
nand U25627 (N_25627,N_22540,N_22545);
nor U25628 (N_25628,N_23098,N_23555);
nor U25629 (N_25629,N_23724,N_22994);
and U25630 (N_25630,N_23873,N_22899);
nand U25631 (N_25631,N_23897,N_23707);
or U25632 (N_25632,N_22713,N_22137);
or U25633 (N_25633,N_23361,N_22201);
nor U25634 (N_25634,N_22990,N_22908);
nor U25635 (N_25635,N_23480,N_23182);
or U25636 (N_25636,N_23658,N_22281);
nand U25637 (N_25637,N_23954,N_22856);
and U25638 (N_25638,N_23414,N_23499);
nand U25639 (N_25639,N_22972,N_23492);
nor U25640 (N_25640,N_22436,N_22407);
or U25641 (N_25641,N_22287,N_23498);
or U25642 (N_25642,N_23028,N_23198);
nand U25643 (N_25643,N_22677,N_22192);
or U25644 (N_25644,N_23041,N_23021);
and U25645 (N_25645,N_23201,N_23030);
nand U25646 (N_25646,N_22156,N_22572);
nand U25647 (N_25647,N_23347,N_23877);
nand U25648 (N_25648,N_22905,N_23669);
or U25649 (N_25649,N_22075,N_23884);
nor U25650 (N_25650,N_22211,N_23608);
xor U25651 (N_25651,N_22276,N_23043);
nand U25652 (N_25652,N_23189,N_22618);
or U25653 (N_25653,N_22001,N_23470);
and U25654 (N_25654,N_23314,N_22087);
xor U25655 (N_25655,N_23562,N_22993);
nand U25656 (N_25656,N_23707,N_23650);
nor U25657 (N_25657,N_22085,N_23207);
xnor U25658 (N_25658,N_22149,N_23862);
or U25659 (N_25659,N_22775,N_22545);
and U25660 (N_25660,N_23658,N_23974);
nor U25661 (N_25661,N_23814,N_22878);
nand U25662 (N_25662,N_23292,N_22931);
nand U25663 (N_25663,N_22964,N_22743);
nor U25664 (N_25664,N_22898,N_23066);
and U25665 (N_25665,N_23279,N_22471);
or U25666 (N_25666,N_23040,N_22151);
xor U25667 (N_25667,N_23523,N_22642);
or U25668 (N_25668,N_23537,N_22255);
xor U25669 (N_25669,N_23322,N_22168);
nor U25670 (N_25670,N_22092,N_23253);
and U25671 (N_25671,N_23013,N_23436);
nor U25672 (N_25672,N_22084,N_22173);
or U25673 (N_25673,N_23898,N_23675);
xnor U25674 (N_25674,N_22257,N_22423);
nor U25675 (N_25675,N_22426,N_23603);
nor U25676 (N_25676,N_23913,N_23146);
and U25677 (N_25677,N_22476,N_22320);
or U25678 (N_25678,N_23748,N_22484);
or U25679 (N_25679,N_23884,N_22060);
nand U25680 (N_25680,N_22612,N_22134);
or U25681 (N_25681,N_23639,N_23107);
nand U25682 (N_25682,N_23642,N_22564);
xor U25683 (N_25683,N_22605,N_22388);
nand U25684 (N_25684,N_23066,N_22138);
or U25685 (N_25685,N_22117,N_22683);
nand U25686 (N_25686,N_22614,N_22236);
or U25687 (N_25687,N_23131,N_23281);
nor U25688 (N_25688,N_22827,N_23674);
or U25689 (N_25689,N_22704,N_22930);
or U25690 (N_25690,N_22351,N_22293);
nor U25691 (N_25691,N_22210,N_22511);
xor U25692 (N_25692,N_23918,N_23422);
or U25693 (N_25693,N_22318,N_23049);
or U25694 (N_25694,N_22549,N_22144);
or U25695 (N_25695,N_22570,N_22823);
and U25696 (N_25696,N_23972,N_22957);
nand U25697 (N_25697,N_22277,N_23874);
nand U25698 (N_25698,N_23966,N_22365);
or U25699 (N_25699,N_22459,N_22683);
xnor U25700 (N_25700,N_23474,N_23130);
nand U25701 (N_25701,N_23587,N_22762);
nor U25702 (N_25702,N_22447,N_22969);
nor U25703 (N_25703,N_23599,N_23892);
nor U25704 (N_25704,N_23148,N_22583);
or U25705 (N_25705,N_23751,N_23447);
nand U25706 (N_25706,N_22865,N_23062);
or U25707 (N_25707,N_22798,N_23516);
and U25708 (N_25708,N_22276,N_23637);
or U25709 (N_25709,N_22871,N_23426);
xor U25710 (N_25710,N_22790,N_23965);
nand U25711 (N_25711,N_22277,N_23705);
or U25712 (N_25712,N_22174,N_22914);
or U25713 (N_25713,N_23577,N_22983);
or U25714 (N_25714,N_23493,N_23139);
or U25715 (N_25715,N_22555,N_23772);
or U25716 (N_25716,N_22652,N_23510);
and U25717 (N_25717,N_22298,N_23381);
nor U25718 (N_25718,N_22282,N_23956);
and U25719 (N_25719,N_23185,N_22553);
nand U25720 (N_25720,N_22324,N_22297);
and U25721 (N_25721,N_23158,N_22714);
and U25722 (N_25722,N_23694,N_22125);
xnor U25723 (N_25723,N_23127,N_23540);
nand U25724 (N_25724,N_22081,N_23146);
and U25725 (N_25725,N_22342,N_23168);
and U25726 (N_25726,N_23140,N_22030);
nand U25727 (N_25727,N_23357,N_23926);
nand U25728 (N_25728,N_22901,N_23799);
xnor U25729 (N_25729,N_23648,N_23480);
or U25730 (N_25730,N_22031,N_22785);
nand U25731 (N_25731,N_22398,N_22762);
xor U25732 (N_25732,N_23323,N_23428);
nand U25733 (N_25733,N_22521,N_22360);
nand U25734 (N_25734,N_23654,N_23554);
nor U25735 (N_25735,N_22473,N_23149);
nor U25736 (N_25736,N_22375,N_22097);
xnor U25737 (N_25737,N_22515,N_23619);
nor U25738 (N_25738,N_23590,N_23195);
or U25739 (N_25739,N_22986,N_23201);
or U25740 (N_25740,N_23479,N_22340);
or U25741 (N_25741,N_22356,N_23168);
and U25742 (N_25742,N_23118,N_23555);
or U25743 (N_25743,N_23756,N_22012);
or U25744 (N_25744,N_23224,N_23555);
and U25745 (N_25745,N_22404,N_23685);
xor U25746 (N_25746,N_22186,N_23536);
and U25747 (N_25747,N_23591,N_23789);
nor U25748 (N_25748,N_23842,N_22555);
xnor U25749 (N_25749,N_22249,N_23388);
xor U25750 (N_25750,N_23730,N_23788);
xor U25751 (N_25751,N_23554,N_23475);
nor U25752 (N_25752,N_22503,N_22994);
and U25753 (N_25753,N_23869,N_22225);
xor U25754 (N_25754,N_22409,N_22870);
and U25755 (N_25755,N_23173,N_22306);
xor U25756 (N_25756,N_22189,N_22283);
nand U25757 (N_25757,N_23927,N_22108);
nand U25758 (N_25758,N_23907,N_23870);
and U25759 (N_25759,N_22499,N_22031);
and U25760 (N_25760,N_22645,N_23902);
or U25761 (N_25761,N_22946,N_22761);
xor U25762 (N_25762,N_22918,N_22782);
xor U25763 (N_25763,N_23268,N_23804);
and U25764 (N_25764,N_22752,N_23412);
nand U25765 (N_25765,N_22287,N_23451);
nor U25766 (N_25766,N_22426,N_23344);
nand U25767 (N_25767,N_23077,N_23817);
xor U25768 (N_25768,N_22864,N_22627);
nor U25769 (N_25769,N_23068,N_22404);
xor U25770 (N_25770,N_23304,N_22922);
nor U25771 (N_25771,N_23930,N_22875);
and U25772 (N_25772,N_23329,N_23858);
nor U25773 (N_25773,N_22212,N_22854);
and U25774 (N_25774,N_22935,N_22173);
or U25775 (N_25775,N_22966,N_22340);
or U25776 (N_25776,N_23418,N_22104);
nand U25777 (N_25777,N_23578,N_22272);
nor U25778 (N_25778,N_22684,N_23851);
xor U25779 (N_25779,N_22763,N_22741);
or U25780 (N_25780,N_22497,N_22013);
nor U25781 (N_25781,N_22764,N_23348);
and U25782 (N_25782,N_22809,N_23848);
xor U25783 (N_25783,N_23755,N_22998);
and U25784 (N_25784,N_23614,N_23092);
and U25785 (N_25785,N_23674,N_23390);
and U25786 (N_25786,N_23033,N_23160);
or U25787 (N_25787,N_22094,N_23327);
xnor U25788 (N_25788,N_23278,N_23072);
nor U25789 (N_25789,N_22482,N_22493);
xnor U25790 (N_25790,N_23396,N_23456);
nand U25791 (N_25791,N_22664,N_23521);
nand U25792 (N_25792,N_22453,N_22420);
and U25793 (N_25793,N_23059,N_23466);
nand U25794 (N_25794,N_22869,N_22347);
nor U25795 (N_25795,N_23601,N_23310);
or U25796 (N_25796,N_23676,N_22044);
and U25797 (N_25797,N_23616,N_22475);
or U25798 (N_25798,N_23019,N_23651);
or U25799 (N_25799,N_22957,N_22993);
or U25800 (N_25800,N_22795,N_22040);
nand U25801 (N_25801,N_22110,N_22125);
nor U25802 (N_25802,N_23156,N_22306);
nor U25803 (N_25803,N_22805,N_22877);
or U25804 (N_25804,N_22338,N_23672);
nor U25805 (N_25805,N_22047,N_23432);
and U25806 (N_25806,N_22438,N_23573);
xor U25807 (N_25807,N_22661,N_22933);
and U25808 (N_25808,N_22089,N_23946);
nand U25809 (N_25809,N_22584,N_23215);
and U25810 (N_25810,N_22873,N_22228);
nand U25811 (N_25811,N_22867,N_23113);
or U25812 (N_25812,N_22098,N_23105);
and U25813 (N_25813,N_22021,N_23847);
xor U25814 (N_25814,N_22215,N_23863);
and U25815 (N_25815,N_23137,N_22032);
nor U25816 (N_25816,N_22654,N_23180);
nand U25817 (N_25817,N_22193,N_22466);
nor U25818 (N_25818,N_22635,N_23689);
and U25819 (N_25819,N_23808,N_23107);
or U25820 (N_25820,N_22910,N_22444);
xnor U25821 (N_25821,N_23211,N_22550);
or U25822 (N_25822,N_22163,N_22477);
nand U25823 (N_25823,N_22458,N_22806);
or U25824 (N_25824,N_22776,N_22950);
nand U25825 (N_25825,N_22575,N_23530);
nand U25826 (N_25826,N_22305,N_22234);
and U25827 (N_25827,N_22220,N_22778);
and U25828 (N_25828,N_22387,N_23039);
or U25829 (N_25829,N_22804,N_23083);
nand U25830 (N_25830,N_22407,N_22168);
and U25831 (N_25831,N_23922,N_23359);
or U25832 (N_25832,N_23694,N_22688);
xnor U25833 (N_25833,N_23840,N_22365);
xnor U25834 (N_25834,N_23330,N_22966);
nor U25835 (N_25835,N_22616,N_22276);
and U25836 (N_25836,N_23782,N_22874);
and U25837 (N_25837,N_23949,N_22486);
and U25838 (N_25838,N_22737,N_22560);
or U25839 (N_25839,N_22957,N_22555);
nand U25840 (N_25840,N_22972,N_22812);
nand U25841 (N_25841,N_22227,N_22512);
or U25842 (N_25842,N_22608,N_22611);
nand U25843 (N_25843,N_23333,N_22731);
xnor U25844 (N_25844,N_22764,N_22847);
nor U25845 (N_25845,N_23085,N_23747);
and U25846 (N_25846,N_22853,N_22438);
nand U25847 (N_25847,N_23790,N_22505);
nor U25848 (N_25848,N_22888,N_22497);
nor U25849 (N_25849,N_22770,N_23362);
nand U25850 (N_25850,N_23210,N_22874);
nand U25851 (N_25851,N_22208,N_22655);
nand U25852 (N_25852,N_22428,N_22625);
and U25853 (N_25853,N_22705,N_22062);
xnor U25854 (N_25854,N_22576,N_23036);
or U25855 (N_25855,N_22479,N_23364);
nor U25856 (N_25856,N_23620,N_22964);
and U25857 (N_25857,N_22413,N_23880);
and U25858 (N_25858,N_22826,N_23331);
nand U25859 (N_25859,N_23446,N_23538);
nand U25860 (N_25860,N_22771,N_23311);
xor U25861 (N_25861,N_23968,N_22721);
and U25862 (N_25862,N_23454,N_23896);
nand U25863 (N_25863,N_22634,N_22740);
or U25864 (N_25864,N_23673,N_23923);
xor U25865 (N_25865,N_23596,N_22585);
nand U25866 (N_25866,N_23360,N_22491);
and U25867 (N_25867,N_23246,N_23134);
nand U25868 (N_25868,N_22843,N_22123);
or U25869 (N_25869,N_22023,N_22454);
nand U25870 (N_25870,N_22996,N_22497);
xnor U25871 (N_25871,N_22982,N_22628);
or U25872 (N_25872,N_22664,N_23745);
xor U25873 (N_25873,N_22395,N_22177);
xnor U25874 (N_25874,N_22229,N_23312);
and U25875 (N_25875,N_22289,N_23433);
and U25876 (N_25876,N_23185,N_22268);
nand U25877 (N_25877,N_22243,N_22956);
nor U25878 (N_25878,N_22863,N_23424);
xor U25879 (N_25879,N_23999,N_23011);
or U25880 (N_25880,N_22832,N_23274);
and U25881 (N_25881,N_22953,N_23740);
or U25882 (N_25882,N_22642,N_23666);
nor U25883 (N_25883,N_22597,N_23826);
or U25884 (N_25884,N_23032,N_23644);
and U25885 (N_25885,N_22015,N_23167);
or U25886 (N_25886,N_22393,N_22214);
nand U25887 (N_25887,N_23912,N_22374);
xor U25888 (N_25888,N_22632,N_22453);
or U25889 (N_25889,N_22018,N_22608);
nor U25890 (N_25890,N_22729,N_22376);
nand U25891 (N_25891,N_23591,N_23853);
and U25892 (N_25892,N_23888,N_23534);
nand U25893 (N_25893,N_22140,N_23761);
or U25894 (N_25894,N_22365,N_22609);
nor U25895 (N_25895,N_23584,N_22219);
nor U25896 (N_25896,N_22435,N_23846);
nand U25897 (N_25897,N_23049,N_22682);
nand U25898 (N_25898,N_23386,N_22228);
and U25899 (N_25899,N_23513,N_22913);
or U25900 (N_25900,N_23655,N_23574);
nand U25901 (N_25901,N_22028,N_23272);
nor U25902 (N_25902,N_22792,N_22752);
or U25903 (N_25903,N_22510,N_23853);
or U25904 (N_25904,N_23431,N_23302);
nor U25905 (N_25905,N_23106,N_22154);
nor U25906 (N_25906,N_23278,N_22373);
nand U25907 (N_25907,N_23165,N_22548);
nand U25908 (N_25908,N_23416,N_22375);
or U25909 (N_25909,N_23797,N_22984);
nor U25910 (N_25910,N_23364,N_22796);
nand U25911 (N_25911,N_22096,N_22795);
and U25912 (N_25912,N_23854,N_22945);
xor U25913 (N_25913,N_23986,N_22593);
xnor U25914 (N_25914,N_22366,N_23798);
nor U25915 (N_25915,N_22281,N_22865);
and U25916 (N_25916,N_23993,N_23315);
nor U25917 (N_25917,N_23001,N_23686);
nand U25918 (N_25918,N_22523,N_23921);
nor U25919 (N_25919,N_22148,N_22859);
nand U25920 (N_25920,N_22137,N_22676);
nor U25921 (N_25921,N_23498,N_22267);
xnor U25922 (N_25922,N_22251,N_22878);
and U25923 (N_25923,N_23918,N_23361);
nand U25924 (N_25924,N_23125,N_22125);
xor U25925 (N_25925,N_22976,N_23200);
and U25926 (N_25926,N_23030,N_22986);
and U25927 (N_25927,N_22382,N_23693);
xnor U25928 (N_25928,N_22783,N_23182);
nor U25929 (N_25929,N_23569,N_23272);
nor U25930 (N_25930,N_22675,N_23866);
nand U25931 (N_25931,N_23106,N_23042);
or U25932 (N_25932,N_22503,N_23327);
nand U25933 (N_25933,N_23091,N_23409);
and U25934 (N_25934,N_22240,N_23179);
or U25935 (N_25935,N_23437,N_23119);
and U25936 (N_25936,N_23031,N_23559);
and U25937 (N_25937,N_22421,N_23741);
xor U25938 (N_25938,N_22171,N_22495);
nand U25939 (N_25939,N_23419,N_22474);
and U25940 (N_25940,N_23017,N_22901);
xnor U25941 (N_25941,N_22278,N_23144);
nor U25942 (N_25942,N_23301,N_23181);
xor U25943 (N_25943,N_23680,N_23187);
and U25944 (N_25944,N_22039,N_23613);
and U25945 (N_25945,N_22404,N_23031);
and U25946 (N_25946,N_23943,N_23784);
nand U25947 (N_25947,N_22002,N_22875);
or U25948 (N_25948,N_22270,N_23415);
or U25949 (N_25949,N_22399,N_22294);
and U25950 (N_25950,N_22414,N_22489);
nand U25951 (N_25951,N_23511,N_22544);
nand U25952 (N_25952,N_22571,N_23924);
nor U25953 (N_25953,N_23674,N_22408);
or U25954 (N_25954,N_23253,N_22383);
and U25955 (N_25955,N_23053,N_22393);
and U25956 (N_25956,N_23514,N_23892);
xnor U25957 (N_25957,N_23357,N_22530);
xor U25958 (N_25958,N_23566,N_23155);
nand U25959 (N_25959,N_22422,N_22068);
xor U25960 (N_25960,N_23761,N_22410);
and U25961 (N_25961,N_22578,N_22563);
nand U25962 (N_25962,N_22529,N_22182);
and U25963 (N_25963,N_23347,N_22551);
and U25964 (N_25964,N_23038,N_23951);
xor U25965 (N_25965,N_23488,N_23135);
xor U25966 (N_25966,N_23778,N_22335);
or U25967 (N_25967,N_22500,N_22124);
xor U25968 (N_25968,N_23561,N_23374);
and U25969 (N_25969,N_22756,N_23189);
nor U25970 (N_25970,N_23558,N_23914);
and U25971 (N_25971,N_22251,N_22203);
nand U25972 (N_25972,N_22127,N_22087);
xnor U25973 (N_25973,N_22066,N_23567);
or U25974 (N_25974,N_23118,N_23727);
or U25975 (N_25975,N_23821,N_23479);
nand U25976 (N_25976,N_22312,N_23356);
nand U25977 (N_25977,N_22470,N_23706);
nor U25978 (N_25978,N_23841,N_23189);
nand U25979 (N_25979,N_23245,N_23501);
nor U25980 (N_25980,N_23662,N_23251);
nor U25981 (N_25981,N_23418,N_22876);
xnor U25982 (N_25982,N_22075,N_22309);
nand U25983 (N_25983,N_22822,N_22329);
or U25984 (N_25984,N_23245,N_23915);
xnor U25985 (N_25985,N_22939,N_22076);
nand U25986 (N_25986,N_22750,N_23732);
nor U25987 (N_25987,N_22854,N_22869);
nor U25988 (N_25988,N_23512,N_22722);
and U25989 (N_25989,N_23425,N_22437);
nor U25990 (N_25990,N_22435,N_22218);
nand U25991 (N_25991,N_22183,N_23012);
or U25992 (N_25992,N_22819,N_22518);
nand U25993 (N_25993,N_22095,N_22514);
xor U25994 (N_25994,N_22712,N_22137);
xnor U25995 (N_25995,N_22220,N_22078);
xnor U25996 (N_25996,N_22119,N_23392);
nor U25997 (N_25997,N_22878,N_22175);
xor U25998 (N_25998,N_23355,N_22921);
or U25999 (N_25999,N_22613,N_22489);
nor U26000 (N_26000,N_24143,N_25476);
and U26001 (N_26001,N_24852,N_25609);
nand U26002 (N_26002,N_25727,N_24174);
or U26003 (N_26003,N_25668,N_25745);
xnor U26004 (N_26004,N_25260,N_25485);
nand U26005 (N_26005,N_24823,N_24659);
and U26006 (N_26006,N_24171,N_25282);
nor U26007 (N_26007,N_25836,N_24597);
nand U26008 (N_26008,N_24731,N_25186);
or U26009 (N_26009,N_24432,N_25189);
and U26010 (N_26010,N_25439,N_24902);
xor U26011 (N_26011,N_25446,N_25837);
xnor U26012 (N_26012,N_24105,N_24637);
and U26013 (N_26013,N_24848,N_25240);
nor U26014 (N_26014,N_24720,N_24081);
nor U26015 (N_26015,N_25377,N_24818);
nor U26016 (N_26016,N_24967,N_24043);
or U26017 (N_26017,N_25208,N_24539);
xnor U26018 (N_26018,N_25433,N_25116);
xnor U26019 (N_26019,N_25110,N_25369);
and U26020 (N_26020,N_25529,N_25629);
nor U26021 (N_26021,N_25974,N_24390);
nand U26022 (N_26022,N_25098,N_24549);
and U26023 (N_26023,N_25472,N_25465);
and U26024 (N_26024,N_24221,N_24477);
and U26025 (N_26025,N_25852,N_25560);
or U26026 (N_26026,N_24610,N_24160);
nor U26027 (N_26027,N_24134,N_25569);
or U26028 (N_26028,N_24781,N_24186);
nor U26029 (N_26029,N_24794,N_24816);
nand U26030 (N_26030,N_24894,N_24126);
xor U26031 (N_26031,N_25677,N_24030);
nor U26032 (N_26032,N_25291,N_25811);
nand U26033 (N_26033,N_24669,N_25900);
xnor U26034 (N_26034,N_24488,N_25449);
or U26035 (N_26035,N_24328,N_25979);
xnor U26036 (N_26036,N_25955,N_24442);
and U26037 (N_26037,N_24289,N_24835);
or U26038 (N_26038,N_25583,N_25448);
and U26039 (N_26039,N_24276,N_24079);
nand U26040 (N_26040,N_24760,N_24972);
nor U26041 (N_26041,N_25849,N_24729);
nor U26042 (N_26042,N_24471,N_24920);
nand U26043 (N_26043,N_24080,N_24837);
or U26044 (N_26044,N_25588,N_24901);
and U26045 (N_26045,N_24849,N_24352);
nand U26046 (N_26046,N_25363,N_25872);
xor U26047 (N_26047,N_24560,N_25555);
xnor U26048 (N_26048,N_25058,N_24527);
nand U26049 (N_26049,N_25086,N_24485);
or U26050 (N_26050,N_24209,N_24065);
nor U26051 (N_26051,N_24858,N_24038);
nor U26052 (N_26052,N_25303,N_24426);
nor U26053 (N_26053,N_25776,N_24495);
and U26054 (N_26054,N_25273,N_25925);
and U26055 (N_26055,N_24064,N_24670);
nand U26056 (N_26056,N_24370,N_25532);
and U26057 (N_26057,N_24959,N_25311);
xor U26058 (N_26058,N_24569,N_25436);
or U26059 (N_26059,N_24071,N_24438);
and U26060 (N_26060,N_24592,N_25480);
nor U26061 (N_26061,N_25182,N_25494);
xor U26062 (N_26062,N_25873,N_24677);
xnor U26063 (N_26063,N_25349,N_25785);
nand U26064 (N_26064,N_25935,N_25947);
and U26065 (N_26065,N_24710,N_25982);
nor U26066 (N_26066,N_24286,N_25392);
nor U26067 (N_26067,N_25784,N_24227);
and U26068 (N_26068,N_24501,N_24980);
and U26069 (N_26069,N_25574,N_24354);
nand U26070 (N_26070,N_25561,N_24392);
xor U26071 (N_26071,N_25918,N_24253);
xnor U26072 (N_26072,N_24779,N_25562);
nand U26073 (N_26073,N_24784,N_25331);
xnor U26074 (N_26074,N_25624,N_24119);
nand U26075 (N_26075,N_24940,N_24383);
or U26076 (N_26076,N_25210,N_24019);
xnor U26077 (N_26077,N_25604,N_25597);
xor U26078 (N_26078,N_24575,N_24326);
nor U26079 (N_26079,N_24244,N_25773);
nand U26080 (N_26080,N_25959,N_25887);
nand U26081 (N_26081,N_25539,N_24210);
or U26082 (N_26082,N_24100,N_24884);
nand U26083 (N_26083,N_25570,N_25545);
and U26084 (N_26084,N_25358,N_24958);
nor U26085 (N_26085,N_25751,N_24216);
or U26086 (N_26086,N_25459,N_25805);
nand U26087 (N_26087,N_24861,N_25062);
or U26088 (N_26088,N_25807,N_24814);
or U26089 (N_26089,N_24552,N_24453);
and U26090 (N_26090,N_24054,N_25848);
and U26091 (N_26091,N_24195,N_24578);
and U26092 (N_26092,N_25664,N_25793);
nor U26093 (N_26093,N_25481,N_24003);
xnor U26094 (N_26094,N_25834,N_24605);
nand U26095 (N_26095,N_24376,N_24773);
nand U26096 (N_26096,N_25654,N_24374);
nand U26097 (N_26097,N_24742,N_25196);
xor U26098 (N_26098,N_25386,N_25989);
xor U26099 (N_26099,N_25296,N_25809);
nand U26100 (N_26100,N_24290,N_24821);
nand U26101 (N_26101,N_25783,N_25053);
and U26102 (N_26102,N_24255,N_24487);
xor U26103 (N_26103,N_25431,N_24166);
nand U26104 (N_26104,N_24943,N_25216);
or U26105 (N_26105,N_24184,N_24270);
xnor U26106 (N_26106,N_24006,N_25272);
xnor U26107 (N_26107,N_24481,N_24142);
and U26108 (N_26108,N_24014,N_25036);
xor U26109 (N_26109,N_25248,N_24306);
or U26110 (N_26110,N_24061,N_24050);
xnor U26111 (N_26111,N_24490,N_25922);
xor U26112 (N_26112,N_24051,N_25307);
nand U26113 (N_26113,N_24518,N_25401);
xnor U26114 (N_26114,N_24382,N_25359);
and U26115 (N_26115,N_24838,N_25200);
nand U26116 (N_26116,N_24904,N_24284);
nor U26117 (N_26117,N_25652,N_25141);
xnor U26118 (N_26118,N_24149,N_25402);
xor U26119 (N_26119,N_24145,N_25040);
nor U26120 (N_26120,N_24625,N_25841);
nand U26121 (N_26121,N_24748,N_24269);
nand U26122 (N_26122,N_25056,N_24070);
xnor U26123 (N_26123,N_24074,N_25398);
nand U26124 (N_26124,N_25428,N_25774);
and U26125 (N_26125,N_25600,N_24308);
nor U26126 (N_26126,N_24893,N_25888);
nand U26127 (N_26127,N_24090,N_24056);
nor U26128 (N_26128,N_24910,N_25142);
nor U26129 (N_26129,N_24939,N_25818);
xnor U26130 (N_26130,N_24235,N_25518);
nand U26131 (N_26131,N_25599,N_24346);
xnor U26132 (N_26132,N_25601,N_25970);
xor U26133 (N_26133,N_25031,N_25237);
xor U26134 (N_26134,N_25894,N_24220);
xnor U26135 (N_26135,N_25128,N_25558);
xor U26136 (N_26136,N_24329,N_25760);
nor U26137 (N_26137,N_24883,N_25091);
nor U26138 (N_26138,N_24749,N_24435);
and U26139 (N_26139,N_25394,N_24663);
nor U26140 (N_26140,N_24895,N_24368);
nand U26141 (N_26141,N_25080,N_25420);
and U26142 (N_26142,N_24826,N_25524);
xnor U26143 (N_26143,N_25670,N_24475);
nor U26144 (N_26144,N_25074,N_25525);
or U26145 (N_26145,N_25068,N_25645);
nor U26146 (N_26146,N_24176,N_24505);
or U26147 (N_26147,N_24387,N_25126);
nand U26148 (N_26148,N_25079,N_24443);
and U26149 (N_26149,N_24686,N_25218);
and U26150 (N_26150,N_25118,N_25617);
and U26151 (N_26151,N_24664,N_24215);
nor U26152 (N_26152,N_24257,N_24218);
nor U26153 (N_26153,N_25715,N_24259);
nand U26154 (N_26154,N_24363,N_24836);
xnor U26155 (N_26155,N_25637,N_25468);
nand U26156 (N_26156,N_24431,N_25350);
nor U26157 (N_26157,N_25180,N_25940);
or U26158 (N_26158,N_24500,N_24707);
nand U26159 (N_26159,N_25452,N_24408);
and U26160 (N_26160,N_25859,N_25860);
nand U26161 (N_26161,N_25926,N_25962);
xnor U26162 (N_26162,N_25846,N_25575);
xnor U26163 (N_26163,N_25564,N_25942);
or U26164 (N_26164,N_25214,N_24879);
or U26165 (N_26165,N_24036,N_24638);
xor U26166 (N_26166,N_24571,N_24639);
nor U26167 (N_26167,N_24744,N_24811);
nand U26168 (N_26168,N_24529,N_25422);
and U26169 (N_26169,N_24267,N_24470);
xnor U26170 (N_26170,N_24704,N_25330);
nor U26171 (N_26171,N_25150,N_25972);
or U26172 (N_26172,N_25673,N_24367);
or U26173 (N_26173,N_24224,N_24379);
nor U26174 (N_26174,N_25317,N_25647);
nand U26175 (N_26175,N_25626,N_24207);
nand U26176 (N_26176,N_24957,N_24878);
xor U26177 (N_26177,N_24199,N_25373);
and U26178 (N_26178,N_24628,N_24337);
or U26179 (N_26179,N_25703,N_25862);
nor U26180 (N_26180,N_25325,N_24551);
xnor U26181 (N_26181,N_25996,N_25538);
xnor U26182 (N_26182,N_24026,N_24076);
and U26183 (N_26183,N_25473,N_24737);
nand U26184 (N_26184,N_24619,N_25021);
xnor U26185 (N_26185,N_25801,N_25740);
nor U26186 (N_26186,N_25650,N_25364);
nand U26187 (N_26187,N_25915,N_24921);
xnor U26188 (N_26188,N_24839,N_24769);
xor U26189 (N_26189,N_24427,N_25850);
xnor U26190 (N_26190,N_25383,N_24110);
and U26191 (N_26191,N_25233,N_24538);
nand U26192 (N_26192,N_24787,N_24122);
nor U26193 (N_26193,N_24589,N_25457);
or U26194 (N_26194,N_24666,N_25826);
nand U26195 (N_26195,N_25298,N_24676);
and U26196 (N_26196,N_25345,N_24687);
nor U26197 (N_26197,N_25666,N_25884);
nor U26198 (N_26198,N_25059,N_25368);
and U26199 (N_26199,N_25840,N_25514);
and U26200 (N_26200,N_25965,N_24898);
or U26201 (N_26201,N_24870,N_25130);
or U26202 (N_26202,N_24739,N_25714);
nand U26203 (N_26203,N_24311,N_25725);
and U26204 (N_26204,N_24712,N_24891);
nor U26205 (N_26205,N_24260,N_25907);
and U26206 (N_26206,N_25831,N_24761);
and U26207 (N_26207,N_25642,N_24283);
nor U26208 (N_26208,N_25050,N_24928);
xor U26209 (N_26209,N_25566,N_25013);
and U26210 (N_26210,N_25313,N_25310);
nor U26211 (N_26211,N_25675,N_24371);
nor U26212 (N_26212,N_25799,N_24189);
xnor U26213 (N_26213,N_25423,N_24124);
nor U26214 (N_26214,N_25095,N_25391);
or U26215 (N_26215,N_25183,N_25354);
or U26216 (N_26216,N_25170,N_25513);
nor U26217 (N_26217,N_25553,N_24701);
and U26218 (N_26218,N_25897,N_25049);
and U26219 (N_26219,N_25447,N_24641);
and U26220 (N_26220,N_24911,N_24730);
nand U26221 (N_26221,N_24449,N_25474);
xor U26222 (N_26222,N_25615,N_25721);
nand U26223 (N_26223,N_25308,N_24468);
xor U26224 (N_26224,N_25206,N_25052);
xnor U26225 (N_26225,N_25691,N_25902);
nand U26226 (N_26226,N_25933,N_24421);
xor U26227 (N_26227,N_25632,N_25794);
nand U26228 (N_26228,N_24588,N_24440);
nor U26229 (N_26229,N_25572,N_25374);
nand U26230 (N_26230,N_24159,N_25334);
xor U26231 (N_26231,N_25226,N_25192);
nor U26232 (N_26232,N_24681,N_24250);
nand U26233 (N_26233,N_25608,N_25775);
xor U26234 (N_26234,N_24718,N_25875);
nand U26235 (N_26235,N_24579,N_25682);
xnor U26236 (N_26236,N_25093,N_25657);
xnor U26237 (N_26237,N_24310,N_24095);
xor U26238 (N_26238,N_25236,N_25026);
or U26239 (N_26239,N_24465,N_25285);
nor U26240 (N_26240,N_25385,N_25193);
or U26241 (N_26241,N_24626,N_25351);
and U26242 (N_26242,N_25415,N_24926);
nor U26243 (N_26243,N_25660,N_24570);
nand U26244 (N_26244,N_24157,N_24553);
nor U26245 (N_26245,N_24041,N_24632);
nor U26246 (N_26246,N_24684,N_25017);
and U26247 (N_26247,N_25782,N_24111);
nor U26248 (N_26248,N_24953,N_24970);
or U26249 (N_26249,N_24247,N_25343);
or U26250 (N_26250,N_25693,N_24585);
nor U26251 (N_26251,N_25618,N_24875);
nor U26252 (N_26252,N_25706,N_25360);
and U26253 (N_26253,N_25024,N_24312);
nor U26254 (N_26254,N_24607,N_25688);
nor U26255 (N_26255,N_25035,N_25424);
nand U26256 (N_26256,N_24966,N_25434);
and U26257 (N_26257,N_25713,N_25992);
and U26258 (N_26258,N_25695,N_25462);
xor U26259 (N_26259,N_25724,N_24219);
xor U26260 (N_26260,N_25766,N_24929);
xor U26261 (N_26261,N_24800,N_25055);
and U26262 (N_26262,N_25496,N_25081);
or U26263 (N_26263,N_24673,N_24073);
nor U26264 (N_26264,N_24042,N_25159);
and U26265 (N_26265,N_25824,N_25143);
and U26266 (N_26266,N_25864,N_24248);
nand U26267 (N_26267,N_24611,N_24001);
xnor U26268 (N_26268,N_24930,N_24600);
xor U26269 (N_26269,N_25270,N_24986);
or U26270 (N_26270,N_24716,N_25023);
nor U26271 (N_26271,N_25027,N_24275);
nand U26272 (N_26272,N_24708,N_24194);
and U26273 (N_26273,N_25039,N_24278);
nor U26274 (N_26274,N_24161,N_24411);
or U26275 (N_26275,N_24776,N_25157);
xnor U26276 (N_26276,N_25502,N_24567);
xnor U26277 (N_26277,N_24254,N_24565);
or U26278 (N_26278,N_25746,N_25295);
and U26279 (N_26279,N_24977,N_25104);
nor U26280 (N_26280,N_24581,N_25038);
nand U26281 (N_26281,N_24905,N_25919);
and U26282 (N_26282,N_24510,N_25771);
or U26283 (N_26283,N_24833,N_24168);
xor U26284 (N_26284,N_25442,N_24492);
and U26285 (N_26285,N_24293,N_24462);
xnor U26286 (N_26286,N_25580,N_25845);
or U26287 (N_26287,N_24546,N_24975);
nor U26288 (N_26288,N_25004,N_24604);
nor U26289 (N_26289,N_25011,N_24738);
xor U26290 (N_26290,N_25557,N_25440);
xnor U26291 (N_26291,N_24745,N_25728);
or U26292 (N_26292,N_25614,N_25758);
or U26293 (N_26293,N_24429,N_24532);
or U26294 (N_26294,N_24947,N_24522);
nand U26295 (N_26295,N_25578,N_24295);
nor U26296 (N_26296,N_24786,N_25762);
and U26297 (N_26297,N_24971,N_24192);
and U26298 (N_26298,N_25777,N_25239);
xor U26299 (N_26299,N_25515,N_24918);
nand U26300 (N_26300,N_25913,N_24706);
xnor U26301 (N_26301,N_24976,N_24467);
or U26302 (N_26302,N_24735,N_25851);
xor U26303 (N_26303,N_25865,N_25191);
nor U26304 (N_26304,N_25504,N_24175);
or U26305 (N_26305,N_24747,N_25981);
nand U26306 (N_26306,N_25261,N_24089);
and U26307 (N_26307,N_25175,N_25719);
nand U26308 (N_26308,N_25503,N_24034);
xnor U26309 (N_26309,N_24436,N_24647);
and U26310 (N_26310,N_25752,N_25347);
or U26311 (N_26311,N_25361,N_24069);
nor U26312 (N_26312,N_24989,N_25149);
xor U26313 (N_26313,N_25500,N_25366);
nand U26314 (N_26314,N_25726,N_24167);
xor U26315 (N_26315,N_24881,N_24242);
or U26316 (N_26316,N_24535,N_25867);
nand U26317 (N_26317,N_24212,N_24832);
or U26318 (N_26318,N_24999,N_24869);
nand U26319 (N_26319,N_25309,N_24507);
xnor U26320 (N_26320,N_24868,N_24562);
xor U26321 (N_26321,N_24923,N_25506);
nor U26322 (N_26322,N_25067,N_24683);
nand U26323 (N_26323,N_24088,N_24000);
nor U26324 (N_26324,N_25432,N_25938);
or U26325 (N_26325,N_25015,N_25305);
or U26326 (N_26326,N_24029,N_25340);
xnor U26327 (N_26327,N_24478,N_24596);
or U26328 (N_26328,N_25292,N_25579);
or U26329 (N_26329,N_24193,N_24951);
or U26330 (N_26330,N_25224,N_25546);
xnor U26331 (N_26331,N_25032,N_24154);
nor U26332 (N_26332,N_25117,N_25648);
nor U26333 (N_26333,N_24360,N_25946);
and U26334 (N_26334,N_25819,N_25491);
nor U26335 (N_26335,N_25978,N_25107);
nand U26336 (N_26336,N_24979,N_25892);
or U26337 (N_26337,N_24332,N_25927);
or U26338 (N_26338,N_24724,N_25679);
or U26339 (N_26339,N_25692,N_25328);
xor U26340 (N_26340,N_25672,N_24114);
and U26341 (N_26341,N_25808,N_24768);
or U26342 (N_26342,N_24452,N_24369);
and U26343 (N_26343,N_24287,N_24358);
and U26344 (N_26344,N_25530,N_25379);
or U26345 (N_26345,N_24827,N_24066);
nand U26346 (N_26346,N_24988,N_25797);
and U26347 (N_26347,N_24099,N_25934);
and U26348 (N_26348,N_24525,N_25533);
or U26349 (N_26349,N_24386,N_25581);
nand U26350 (N_26350,N_25202,N_24464);
or U26351 (N_26351,N_24316,N_24874);
nor U26352 (N_26352,N_24617,N_25611);
xor U26353 (N_26353,N_25968,N_24450);
nand U26354 (N_26354,N_24872,N_24807);
nand U26355 (N_26355,N_24851,N_25499);
nand U26356 (N_26356,N_25057,N_24506);
and U26357 (N_26357,N_25071,N_24262);
nand U26358 (N_26358,N_24646,N_24726);
and U26359 (N_26359,N_25390,N_25610);
nand U26360 (N_26360,N_25286,N_25871);
or U26361 (N_26361,N_24472,N_24795);
xor U26362 (N_26362,N_24648,N_24048);
and U26363 (N_26363,N_24946,N_25245);
or U26364 (N_26364,N_25928,N_25960);
nor U26365 (N_26365,N_24956,N_24335);
and U26366 (N_26366,N_25230,N_24927);
xnor U26367 (N_26367,N_25228,N_24954);
nor U26368 (N_26368,N_24138,N_24734);
or U26369 (N_26369,N_24547,N_25644);
nand U26370 (N_26370,N_24564,N_25522);
or U26371 (N_26371,N_25382,N_25041);
and U26372 (N_26372,N_25467,N_25352);
or U26373 (N_26373,N_25160,N_25847);
nand U26374 (N_26374,N_24780,N_24251);
nor U26375 (N_26375,N_24318,N_25607);
nand U26376 (N_26376,N_25399,N_24185);
xnor U26377 (N_26377,N_25000,N_24889);
or U26378 (N_26378,N_25283,N_25795);
or U26379 (N_26379,N_24533,N_24765);
or U26380 (N_26380,N_25620,N_24087);
nor U26381 (N_26381,N_25895,N_24645);
nor U26382 (N_26382,N_24256,N_25127);
nand U26383 (N_26383,N_24653,N_25696);
and U26384 (N_26384,N_24568,N_25221);
nand U26385 (N_26385,N_24615,N_24321);
nor U26386 (N_26386,N_24840,N_24294);
or U26387 (N_26387,N_24391,N_24350);
nand U26388 (N_26388,N_25507,N_24711);
xnor U26389 (N_26389,N_24595,N_24211);
and U26390 (N_26390,N_25855,N_25757);
or U26391 (N_26391,N_24530,N_24058);
nor U26392 (N_26392,N_24348,N_24356);
and U26393 (N_26393,N_25587,N_25028);
and U26394 (N_26394,N_24446,N_24300);
xnor U26395 (N_26395,N_25700,N_25112);
xor U26396 (N_26396,N_25199,N_25842);
nand U26397 (N_26397,N_24053,N_25323);
nand U26398 (N_26398,N_25014,N_24824);
nor U26399 (N_26399,N_24324,N_25077);
and U26400 (N_26400,N_25863,N_24609);
nor U26401 (N_26401,N_24480,N_25523);
and U26402 (N_26402,N_25950,N_25921);
nand U26403 (N_26403,N_24876,N_25250);
or U26404 (N_26404,N_25134,N_24912);
nor U26405 (N_26405,N_25742,N_24655);
and U26406 (N_26406,N_25162,N_24753);
nand U26407 (N_26407,N_24576,N_24743);
nor U26408 (N_26408,N_25698,N_25627);
nand U26409 (N_26409,N_24715,N_24937);
or U26410 (N_26410,N_25409,N_25042);
xor U26411 (N_26411,N_25516,N_24170);
nor U26412 (N_26412,N_25177,N_24799);
and U26413 (N_26413,N_25109,N_25763);
nor U26414 (N_26414,N_24112,N_25596);
and U26415 (N_26415,N_24936,N_24156);
nand U26416 (N_26416,N_24380,N_25262);
xor U26417 (N_26417,N_24320,N_25576);
nand U26418 (N_26418,N_24213,N_24005);
nor U26419 (N_26419,N_25490,N_25078);
xnor U26420 (N_26420,N_24841,N_24092);
nor U26421 (N_26421,N_24394,N_24016);
nor U26422 (N_26422,N_24430,N_24888);
or U26423 (N_26423,N_25868,N_25622);
and U26424 (N_26424,N_25806,N_25097);
or U26425 (N_26425,N_25945,N_24085);
or U26426 (N_26426,N_25563,N_24689);
or U26427 (N_26427,N_24123,N_25941);
or U26428 (N_26428,N_25289,N_24288);
nor U26429 (N_26429,N_25378,N_24031);
xor U26430 (N_26430,N_25461,N_25844);
xor U26431 (N_26431,N_24634,N_25591);
nand U26432 (N_26432,N_25293,N_24125);
nand U26433 (N_26433,N_25976,N_25075);
nand U26434 (N_26434,N_24855,N_24489);
and U26435 (N_26435,N_25621,N_25344);
or U26436 (N_26436,N_25280,N_24545);
and U26437 (N_26437,N_25710,N_24130);
and U26438 (N_26438,N_24407,N_25803);
nor U26439 (N_26439,N_25674,N_24860);
nor U26440 (N_26440,N_24766,N_24322);
or U26441 (N_26441,N_25048,N_25636);
nand U26442 (N_26442,N_24046,N_24828);
nand U26443 (N_26443,N_25163,N_25115);
and U26444 (N_26444,N_25426,N_24792);
and U26445 (N_26445,N_25619,N_25658);
xnor U26446 (N_26446,N_24059,N_25526);
nand U26447 (N_26447,N_24317,N_25069);
or U26448 (N_26448,N_24083,N_25786);
xor U26449 (N_26449,N_25967,N_24373);
or U26450 (N_26450,N_24230,N_25279);
nand U26451 (N_26451,N_24401,N_25635);
nor U26452 (N_26452,N_24830,N_25251);
or U26453 (N_26453,N_25764,N_24182);
nand U26454 (N_26454,N_24796,N_25554);
or U26455 (N_26455,N_25277,N_25899);
nor U26456 (N_26456,N_24002,N_24172);
nor U26457 (N_26457,N_24974,N_25005);
xnor U26458 (N_26458,N_25891,N_25090);
nor U26459 (N_26459,N_24118,N_25043);
nand U26460 (N_26460,N_25445,N_25723);
or U26461 (N_26461,N_25037,N_25737);
xor U26462 (N_26462,N_24150,N_24817);
nand U26463 (N_26463,N_24508,N_25625);
xor U26464 (N_26464,N_25889,N_25536);
nor U26465 (N_26465,N_25178,N_24528);
nor U26466 (N_26466,N_25137,N_25707);
xor U26467 (N_26467,N_25756,N_24397);
xnor U26468 (N_26468,N_25717,N_25393);
nor U26469 (N_26469,N_24035,N_25856);
nand U26470 (N_26470,N_24147,N_24829);
nand U26471 (N_26471,N_25821,N_25547);
xnor U26472 (N_26472,N_24187,N_25874);
nand U26473 (N_26473,N_24146,N_25264);
nor U26474 (N_26474,N_25898,N_24815);
nand U26475 (N_26475,N_25087,N_25744);
and U26476 (N_26476,N_24234,N_24691);
nand U26477 (N_26477,N_25092,N_24563);
and U26478 (N_26478,N_25788,N_25259);
xor U26479 (N_26479,N_24757,N_25920);
and U26480 (N_26480,N_24665,N_25991);
and U26481 (N_26481,N_25201,N_25094);
and U26482 (N_26482,N_24011,N_25132);
xnor U26483 (N_26483,N_24594,N_24128);
or U26484 (N_26484,N_24654,N_24094);
xor U26485 (N_26485,N_24789,N_24225);
or U26486 (N_26486,N_24107,N_25733);
and U26487 (N_26487,N_24762,N_24703);
nand U26488 (N_26488,N_24602,N_24273);
or U26489 (N_26489,N_25861,N_25400);
or U26490 (N_26490,N_24381,N_25640);
and U26491 (N_26491,N_24494,N_24351);
xor U26492 (N_26492,N_24217,N_24922);
nor U26493 (N_26493,N_25302,N_24614);
and U26494 (N_26494,N_24877,N_25893);
nor U26495 (N_26495,N_25505,N_25222);
nand U26496 (N_26496,N_25911,N_24345);
xnor U26497 (N_26497,N_25594,N_24709);
nand U26498 (N_26498,N_25438,N_24559);
and U26499 (N_26499,N_25930,N_24537);
nand U26500 (N_26500,N_24499,N_25829);
or U26501 (N_26501,N_24237,N_25969);
and U26502 (N_26502,N_24414,N_24997);
nor U26503 (N_26503,N_25906,N_25321);
or U26504 (N_26504,N_25407,N_24636);
xor U26505 (N_26505,N_25217,N_24424);
xnor U26506 (N_26506,N_24635,N_24025);
or U26507 (N_26507,N_25954,N_24844);
or U26508 (N_26508,N_25096,N_25255);
and U26509 (N_26509,N_25122,N_24004);
and U26510 (N_26510,N_24620,N_24842);
and U26511 (N_26511,N_24834,N_24422);
and U26512 (N_26512,N_25376,N_24469);
and U26513 (N_26513,N_25082,N_25729);
nor U26514 (N_26514,N_24583,N_24133);
and U26515 (N_26515,N_25616,N_24859);
xnor U26516 (N_26516,N_24330,N_24458);
or U26517 (N_26517,N_24153,N_25121);
or U26518 (N_26518,N_25275,N_24513);
or U26519 (N_26519,N_25164,N_24613);
xor U26520 (N_26520,N_24204,N_24987);
xnor U26521 (N_26521,N_24274,N_25337);
nor U26522 (N_26522,N_24882,N_24674);
or U26523 (N_26523,N_24733,N_25903);
or U26524 (N_26524,N_25019,N_25244);
nand U26525 (N_26525,N_25767,N_24266);
nor U26526 (N_26526,N_25252,N_24314);
nor U26527 (N_26527,N_25413,N_24077);
xor U26528 (N_26528,N_24309,N_25662);
xnor U26529 (N_26529,N_25661,N_24361);
nand U26530 (N_26530,N_24968,N_24804);
or U26531 (N_26531,N_24678,N_25129);
xor U26532 (N_26532,N_24845,N_25284);
nand U26533 (N_26533,N_24033,N_25215);
or U26534 (N_26534,N_24767,N_25810);
and U26535 (N_26535,N_24960,N_24866);
nor U26536 (N_26536,N_25478,N_25338);
and U26537 (N_26537,N_24517,N_24139);
xor U26538 (N_26538,N_25362,N_25550);
nand U26539 (N_26539,N_24023,N_25412);
and U26540 (N_26540,N_25663,N_25548);
xor U26541 (N_26541,N_24214,N_24694);
or U26542 (N_26542,N_25408,N_25983);
or U26543 (N_26543,N_24909,N_25381);
or U26544 (N_26544,N_25429,N_25731);
nor U26545 (N_26545,N_24479,N_25316);
nor U26546 (N_26546,N_25070,N_24203);
nor U26547 (N_26547,N_24498,N_25667);
or U26548 (N_26548,N_24873,N_24802);
and U26549 (N_26549,N_25741,N_25229);
and U26550 (N_26550,N_24657,N_25384);
xor U26551 (N_26551,N_25879,N_25489);
nand U26552 (N_26552,N_25089,N_24758);
xnor U26553 (N_26553,N_24086,N_25908);
or U26554 (N_26554,N_25995,N_24336);
xnor U26555 (N_26555,N_25312,N_25577);
or U26556 (N_26556,N_24245,N_24932);
nand U26557 (N_26557,N_24304,N_25455);
or U26558 (N_26558,N_24994,N_25441);
nor U26559 (N_26559,N_24075,N_24934);
nand U26560 (N_26560,N_24944,N_25531);
or U26561 (N_26561,N_24521,N_25194);
or U26562 (N_26562,N_24511,N_25167);
nand U26563 (N_26563,N_25593,N_24299);
or U26564 (N_26564,N_25589,N_25905);
and U26565 (N_26565,N_25778,N_25464);
xnor U26566 (N_26566,N_24591,N_24447);
and U26567 (N_26567,N_24378,N_25120);
xor U26568 (N_26568,N_25559,N_24141);
or U26569 (N_26569,N_24377,N_25508);
xor U26570 (N_26570,N_25443,N_24037);
xnor U26571 (N_26571,N_25348,N_24151);
and U26572 (N_26572,N_25007,N_24268);
or U26573 (N_26573,N_24406,N_25754);
and U26574 (N_26574,N_24136,N_24137);
xor U26575 (N_26575,N_24992,N_24696);
and U26576 (N_26576,N_24082,N_25697);
nand U26577 (N_26577,N_25483,N_25022);
or U26578 (N_26578,N_25813,N_25971);
and U26579 (N_26579,N_25155,N_25796);
nand U26580 (N_26580,N_25268,N_25100);
and U26581 (N_26581,N_24165,N_25397);
and U26582 (N_26582,N_24102,N_25169);
or U26583 (N_26583,N_24454,N_25866);
and U26584 (N_26584,N_24574,N_25147);
nand U26585 (N_26585,N_25403,N_25179);
nand U26586 (N_26586,N_25659,N_25790);
xor U26587 (N_26587,N_24612,N_25822);
nand U26588 (N_26588,N_25534,N_24423);
and U26589 (N_26589,N_25466,N_24996);
nand U26590 (N_26590,N_25498,N_24398);
nand U26591 (N_26591,N_25001,N_24177);
or U26592 (N_26592,N_25002,N_25463);
or U26593 (N_26593,N_25243,N_24652);
nor U26594 (N_26594,N_25009,N_25857);
nand U26595 (N_26595,N_25772,N_24365);
and U26596 (N_26596,N_25738,N_25712);
nor U26597 (N_26597,N_25044,N_25732);
nor U26598 (N_26598,N_24667,N_25683);
nand U26599 (N_26599,N_25314,N_24399);
or U26600 (N_26600,N_25495,N_25145);
nor U26601 (N_26601,N_24756,N_24417);
xor U26602 (N_26602,N_25598,N_24072);
xnor U26603 (N_26603,N_24364,N_24202);
nand U26604 (N_26604,N_25988,N_25300);
nand U26605 (N_26605,N_24344,N_24403);
or U26606 (N_26606,N_24343,N_24969);
or U26607 (N_26607,N_24948,N_25939);
nand U26608 (N_26608,N_24693,N_25643);
nand U26609 (N_26609,N_25628,N_25198);
and U26610 (N_26610,N_25932,N_24032);
nand U26611 (N_26611,N_25045,N_24445);
nor U26612 (N_26612,N_24846,N_24721);
xnor U26613 (N_26613,N_25568,N_24750);
xnor U26614 (N_26614,N_25247,N_25681);
xnor U26615 (N_26615,N_24272,N_24995);
or U26616 (N_26616,N_25084,N_24697);
nor U26617 (N_26617,N_25694,N_24764);
and U26618 (N_26618,N_25136,N_24109);
or U26619 (N_26619,N_24451,N_24949);
or U26620 (N_26620,N_25029,N_25389);
nor U26621 (N_26621,N_24319,N_24941);
or U26622 (N_26622,N_25185,N_24205);
nor U26623 (N_26623,N_24474,N_25114);
xor U26624 (N_26624,N_24323,N_24012);
nand U26625 (N_26625,N_25003,N_25356);
xor U26626 (N_26626,N_25460,N_25649);
or U26627 (N_26627,N_25235,N_25257);
nand U26628 (N_26628,N_25416,N_25838);
and U26629 (N_26629,N_24908,N_25421);
nor U26630 (N_26630,N_25319,N_24339);
nor U26631 (N_26631,N_24732,N_25488);
nor U26632 (N_26632,N_24950,N_24459);
and U26633 (N_26633,N_24722,N_25605);
nor U26634 (N_26634,N_24806,N_24942);
nor U26635 (N_26635,N_24463,N_24018);
xnor U26636 (N_26636,N_25006,N_24973);
or U26637 (N_26637,N_25065,N_25552);
or U26638 (N_26638,N_24935,N_24264);
or U26639 (N_26639,N_25105,N_25749);
nand U26640 (N_26640,N_24717,N_25975);
xor U26641 (N_26641,N_24754,N_25750);
and U26642 (N_26642,N_25238,N_25174);
and U26643 (N_26643,N_24650,N_25761);
xnor U26644 (N_26644,N_25511,N_24965);
and U26645 (N_26645,N_24627,N_25227);
nor U26646 (N_26646,N_25602,N_24593);
nand U26647 (N_26647,N_25102,N_24301);
xnor U26648 (N_26648,N_25549,N_25612);
nand U26649 (N_26649,N_25886,N_24907);
or U26650 (N_26650,N_25181,N_25395);
nor U26651 (N_26651,N_25025,N_24084);
nor U26652 (N_26652,N_24419,N_25073);
or U26653 (N_26653,N_24801,N_25521);
and U26654 (N_26654,N_24484,N_24491);
and U26655 (N_26655,N_25747,N_24808);
or U26656 (N_26656,N_25680,N_24180);
and U26657 (N_26657,N_25800,N_24790);
xor U26658 (N_26658,N_25917,N_25301);
xnor U26659 (N_26659,N_25492,N_25708);
or U26660 (N_26660,N_24384,N_24482);
and U26661 (N_26661,N_25770,N_24695);
and U26662 (N_26662,N_25371,N_25937);
and U26663 (N_26663,N_24347,N_25405);
and U26664 (N_26664,N_24978,N_25326);
nand U26665 (N_26665,N_24104,N_24353);
xor U26666 (N_26666,N_25220,N_24437);
nand U26667 (N_26667,N_24389,N_24728);
nand U26668 (N_26668,N_25595,N_24206);
nor U26669 (N_26669,N_25630,N_24961);
xor U26670 (N_26670,N_25336,N_24582);
and U26671 (N_26671,N_25205,N_24196);
nor U26672 (N_26672,N_25197,N_25276);
nand U26673 (N_26673,N_24007,N_24671);
and U26674 (N_26674,N_25791,N_25010);
and U26675 (N_26675,N_25685,N_24524);
and U26676 (N_26676,N_24982,N_24658);
and U26677 (N_26677,N_25711,N_25997);
or U26678 (N_26678,N_25702,N_25258);
xor U26679 (N_26679,N_25823,N_25173);
nand U26680 (N_26680,N_25961,N_24342);
xnor U26681 (N_26681,N_24777,N_25966);
nor U26682 (N_26682,N_24915,N_25669);
xor U26683 (N_26683,N_25520,N_25765);
xnor U26684 (N_26684,N_25869,N_24584);
xnor U26685 (N_26685,N_25139,N_24577);
or U26686 (N_26686,N_24865,N_24685);
or U26687 (N_26687,N_24413,N_25324);
and U26688 (N_26688,N_24404,N_25551);
nor U26689 (N_26689,N_24473,N_24534);
and U26690 (N_26690,N_24543,N_25063);
nor U26691 (N_26691,N_25166,N_25993);
nor U26692 (N_26692,N_25088,N_25380);
nand U26693 (N_26693,N_24113,N_25832);
or U26694 (N_26694,N_24621,N_25083);
xnor U26695 (N_26695,N_24420,N_25234);
xor U26696 (N_26696,N_25353,N_25542);
nand U26697 (N_26697,N_25209,N_25814);
xnor U26698 (N_26698,N_24772,N_25678);
nor U26699 (N_26699,N_24778,N_25211);
or U26700 (N_26700,N_25686,N_24410);
nand U26701 (N_26701,N_25843,N_25825);
and U26702 (N_26702,N_25963,N_24662);
nor U26703 (N_26703,N_24045,N_25299);
nor U26704 (N_26704,N_24412,N_25158);
nor U26705 (N_26705,N_25320,N_25603);
and U26706 (N_26706,N_25684,N_25064);
nor U26707 (N_26707,N_24013,N_24991);
xnor U26708 (N_26708,N_25290,N_24483);
xor U26709 (N_26709,N_24393,N_24331);
nand U26710 (N_26710,N_25676,N_24497);
nor U26711 (N_26711,N_24618,N_24243);
nand U26712 (N_26712,N_24572,N_25288);
nand U26713 (N_26713,N_25123,N_24587);
nor U26714 (N_26714,N_25047,N_24162);
or U26715 (N_26715,N_25051,N_25454);
nand U26716 (N_26716,N_24642,N_24751);
or U26717 (N_26717,N_25493,N_25820);
nor U26718 (N_26718,N_24516,N_25111);
nor U26719 (N_26719,N_25929,N_24871);
nand U26720 (N_26720,N_24372,N_24279);
nor U26721 (N_26721,N_25585,N_25878);
nor U26722 (N_26722,N_24121,N_25882);
nor U26723 (N_26723,N_25651,N_24897);
or U26724 (N_26724,N_24847,N_25722);
nand U26725 (N_26725,N_25901,N_24925);
xor U26726 (N_26726,N_25131,N_25914);
nor U26727 (N_26727,N_25339,N_24285);
nor U26728 (N_26728,N_24805,N_25225);
nor U26729 (N_26729,N_24763,N_25396);
xnor U26730 (N_26730,N_24850,N_25475);
nand U26731 (N_26731,N_24785,N_24233);
or U26732 (N_26732,N_25176,N_25453);
xor U26733 (N_26733,N_24558,N_25242);
nor U26734 (N_26734,N_25817,N_25709);
and U26735 (N_26735,N_24425,N_25430);
nor U26736 (N_26736,N_24906,N_24307);
or U26737 (N_26737,N_24190,N_25986);
nor U26738 (N_26738,N_24448,N_24962);
nand U26739 (N_26739,N_24238,N_25537);
or U26740 (N_26740,N_25753,N_24093);
nand U26741 (N_26741,N_24049,N_24357);
nor U26742 (N_26742,N_24554,N_25781);
xnor U26743 (N_26743,N_24649,N_24963);
xnor U26744 (N_26744,N_25987,N_24232);
or U26745 (N_26745,N_24998,N_24418);
nand U26746 (N_26746,N_24249,N_24362);
xor U26747 (N_26747,N_24556,N_24813);
nor U26748 (N_26748,N_24782,N_24240);
xnor U26749 (N_26749,N_25099,N_25964);
xor U26750 (N_26750,N_25318,N_25335);
and U26751 (N_26751,N_25948,N_24236);
nor U26752 (N_26752,N_25730,N_25444);
xor U26753 (N_26753,N_25287,N_25590);
xor U26754 (N_26754,N_24810,N_25406);
or U26755 (N_26755,N_25881,N_24017);
or U26756 (N_26756,N_25671,N_24178);
nand U26757 (N_26757,N_25567,N_24044);
nor U26758 (N_26758,N_25606,N_24129);
and U26759 (N_26759,N_24688,N_24366);
nor U26760 (N_26760,N_24981,N_25484);
nand U26761 (N_26761,N_25195,N_24740);
nor U26762 (N_26762,N_25736,N_24651);
or U26763 (N_26763,N_24444,N_24931);
and U26764 (N_26764,N_25512,N_24512);
or U26765 (N_26765,N_25207,N_24395);
nor U26766 (N_26766,N_25103,N_25066);
or U26767 (N_26767,N_25125,N_24705);
and U26768 (N_26768,N_24887,N_24015);
nor U26769 (N_26769,N_25154,N_24198);
nand U26770 (N_26770,N_25739,N_24867);
and U26771 (N_26771,N_25854,N_24900);
nor U26772 (N_26772,N_25748,N_25315);
nand U26773 (N_26773,N_24120,N_24258);
nor U26774 (N_26774,N_24163,N_24812);
or U26775 (N_26775,N_24280,N_25734);
or U26776 (N_26776,N_24021,N_24863);
and U26777 (N_26777,N_25486,N_25973);
xnor U26778 (N_26778,N_25171,N_24263);
xor U26779 (N_26779,N_24457,N_25980);
or U26780 (N_26780,N_24774,N_24598);
nand U26781 (N_26781,N_24252,N_25148);
nand U26782 (N_26782,N_24820,N_25858);
or U26783 (N_26783,N_24291,N_25151);
xnor U26784 (N_26784,N_25984,N_24057);
and U26785 (N_26785,N_25653,N_25135);
xnor U26786 (N_26786,N_24656,N_24679);
or U26787 (N_26787,N_25153,N_24544);
nand U26788 (N_26788,N_25184,N_24542);
and U26789 (N_26789,N_24913,N_25266);
or U26790 (N_26790,N_24886,N_25269);
xnor U26791 (N_26791,N_24690,N_24985);
or U26792 (N_26792,N_24952,N_24914);
nand U26793 (N_26793,N_24292,N_25720);
or U26794 (N_26794,N_25332,N_25885);
nor U26795 (N_26795,N_24573,N_25168);
and U26796 (N_26796,N_24783,N_25144);
xor U26797 (N_26797,N_24040,N_24327);
nor U26798 (N_26798,N_24550,N_24531);
or U26799 (N_26799,N_24561,N_24349);
xnor U26800 (N_26800,N_25418,N_24788);
or U26801 (N_26801,N_25718,N_24509);
nand U26802 (N_26802,N_25487,N_24200);
nand U26803 (N_26803,N_25477,N_25357);
nor U26804 (N_26804,N_25896,N_24144);
xor U26805 (N_26805,N_24271,N_24629);
or U26806 (N_26806,N_24885,N_24924);
nor U26807 (N_26807,N_24759,N_24132);
nor U26808 (N_26808,N_25953,N_24239);
nand U26809 (N_26809,N_25263,N_25203);
and U26810 (N_26810,N_25140,N_25076);
nand U26811 (N_26811,N_24340,N_24359);
or U26812 (N_26812,N_24298,N_24405);
and U26813 (N_26813,N_25528,N_25161);
nor U26814 (N_26814,N_25510,N_25699);
xnor U26815 (N_26815,N_24736,N_24938);
nand U26816 (N_26816,N_25519,N_25034);
or U26817 (N_26817,N_24723,N_25367);
nand U26818 (N_26818,N_25008,N_24179);
or U26819 (N_26819,N_25232,N_25815);
nor U26820 (N_26820,N_25410,N_24606);
or U26821 (N_26821,N_25880,N_24682);
nor U26822 (N_26822,N_24158,N_24557);
nand U26823 (N_26823,N_25769,N_25417);
and U26824 (N_26824,N_25517,N_24067);
nand U26825 (N_26825,N_25333,N_25877);
or U26826 (N_26826,N_25634,N_24188);
or U26827 (N_26827,N_24504,N_24131);
nand U26828 (N_26828,N_24890,N_24672);
or U26829 (N_26829,N_24402,N_25387);
and U26830 (N_26830,N_24140,N_25924);
nand U26831 (N_26831,N_25584,N_25437);
xor U26832 (N_26832,N_25018,N_24486);
nand U26833 (N_26833,N_24409,N_24098);
and U26834 (N_26834,N_24010,N_25952);
and U26835 (N_26835,N_24456,N_25172);
nand U26836 (N_26836,N_25271,N_25789);
xor U26837 (N_26837,N_24586,N_24831);
nor U26838 (N_26838,N_24461,N_24208);
xnor U26839 (N_26839,N_24039,N_25690);
or U26840 (N_26840,N_25957,N_24984);
nand U26841 (N_26841,N_24993,N_24155);
nand U26842 (N_26842,N_24590,N_25909);
and U26843 (N_26843,N_24009,N_24752);
or U26844 (N_26844,N_25212,N_24024);
and U26845 (N_26845,N_24265,N_25787);
or U26846 (N_26846,N_24630,N_24809);
xor U26847 (N_26847,N_24822,N_24428);
xor U26848 (N_26848,N_25456,N_25910);
nand U26849 (N_26849,N_25543,N_24434);
and U26850 (N_26850,N_24917,N_24455);
or U26851 (N_26851,N_24523,N_25916);
nand U26852 (N_26852,N_25241,N_24416);
nor U26853 (N_26853,N_24680,N_24644);
or U26854 (N_26854,N_25046,N_25743);
and U26855 (N_26855,N_24541,N_24164);
xnor U26856 (N_26856,N_25853,N_25944);
or U26857 (N_26857,N_24580,N_24027);
nand U26858 (N_26858,N_25213,N_24338);
xnor U26859 (N_26859,N_25998,N_25571);
xnor U26860 (N_26860,N_24746,N_25792);
nor U26861 (N_26861,N_24700,N_25471);
or U26862 (N_26862,N_25833,N_24315);
nor U26863 (N_26863,N_24183,N_24460);
nor U26864 (N_26864,N_24631,N_24548);
xnor U26865 (N_26865,N_24047,N_24222);
xnor U26866 (N_26866,N_25779,N_25704);
nor U26867 (N_26867,N_25119,N_24519);
nand U26868 (N_26868,N_24640,N_25327);
xor U26869 (N_26869,N_25586,N_25304);
or U26870 (N_26870,N_25951,N_24514);
nand U26871 (N_26871,N_25641,N_25306);
nor U26872 (N_26872,N_25501,N_24856);
nor U26873 (N_26873,N_25372,N_24843);
or U26874 (N_26874,N_24020,N_25994);
or U26875 (N_26875,N_25450,N_25535);
and U26876 (N_26876,N_24608,N_24060);
nor U26877 (N_26877,N_24116,N_24725);
nand U26878 (N_26878,N_25458,N_25482);
or U26879 (N_26879,N_24282,N_24466);
or U26880 (N_26880,N_24028,N_25613);
or U26881 (N_26881,N_24945,N_25278);
xnor U26882 (N_26882,N_25479,N_25254);
nand U26883 (N_26883,N_25509,N_24798);
nor U26884 (N_26884,N_24616,N_25999);
nand U26885 (N_26885,N_25812,N_25890);
nand U26886 (N_26886,N_24476,N_24229);
and U26887 (N_26887,N_25265,N_25020);
nor U26888 (N_26888,N_25219,N_24173);
nand U26889 (N_26889,N_25827,N_25828);
nor U26890 (N_26890,N_25322,N_25870);
and U26891 (N_26891,N_25931,N_24896);
nand U26892 (N_26892,N_25346,N_24668);
nor U26893 (N_26893,N_24008,N_24503);
nor U26894 (N_26894,N_25256,N_25294);
nor U26895 (N_26895,N_24117,N_25204);
nor U26896 (N_26896,N_24433,N_25267);
nand U26897 (N_26897,N_24296,N_25370);
xnor U26898 (N_26898,N_24864,N_25780);
or U26899 (N_26899,N_24334,N_24692);
nor U26900 (N_26900,N_25249,N_24068);
nand U26901 (N_26901,N_25689,N_25329);
and U26902 (N_26902,N_24990,N_25656);
nor U26903 (N_26903,N_24191,N_25124);
nand U26904 (N_26904,N_24853,N_25943);
nor U26905 (N_26905,N_24526,N_24964);
or U26906 (N_26906,N_24355,N_24983);
and U26907 (N_26907,N_24603,N_25541);
or U26908 (N_26908,N_24169,N_24281);
or U26909 (N_26909,N_25425,N_24152);
nor U26910 (N_26910,N_24228,N_24305);
and U26911 (N_26911,N_24226,N_24135);
nand U26912 (N_26912,N_24148,N_24727);
xnor U26913 (N_26913,N_24899,N_24297);
nor U26914 (N_26914,N_25904,N_24493);
and U26915 (N_26915,N_25977,N_24246);
or U26916 (N_26916,N_25231,N_24622);
or U26917 (N_26917,N_24223,N_25705);
nor U26918 (N_26918,N_24097,N_24063);
xor U26919 (N_26919,N_25341,N_24698);
nor U26920 (N_26920,N_25768,N_25106);
nor U26921 (N_26921,N_25469,N_25072);
xnor U26922 (N_26922,N_25016,N_25108);
or U26923 (N_26923,N_24496,N_25297);
and U26924 (N_26924,N_25190,N_24862);
and U26925 (N_26925,N_25152,N_25835);
nor U26926 (N_26926,N_24520,N_24333);
nor U26927 (N_26927,N_24277,N_25342);
or U26928 (N_26928,N_25138,N_25246);
xor U26929 (N_26929,N_25497,N_25365);
and U26930 (N_26930,N_25912,N_25527);
nand U26931 (N_26931,N_24633,N_24770);
nand U26932 (N_26932,N_24325,N_24303);
nand U26933 (N_26933,N_24719,N_25388);
xor U26934 (N_26934,N_24803,N_25631);
nor U26935 (N_26935,N_24675,N_24955);
nand U26936 (N_26936,N_24341,N_24903);
xor U26937 (N_26937,N_24540,N_25956);
nor U26938 (N_26938,N_24892,N_25556);
nand U26939 (N_26939,N_24825,N_25839);
nor U26940 (N_26940,N_24106,N_24201);
nand U26941 (N_26941,N_24566,N_25146);
xor U26942 (N_26942,N_25876,N_25427);
or U26943 (N_26943,N_25033,N_24919);
xnor U26944 (N_26944,N_24022,N_24755);
nand U26945 (N_26945,N_25883,N_24699);
or U26946 (N_26946,N_24771,N_24103);
nand U26947 (N_26947,N_24052,N_24660);
nand U26948 (N_26948,N_25165,N_24091);
or U26949 (N_26949,N_24127,N_24375);
or U26950 (N_26950,N_25633,N_24916);
nand U26951 (N_26951,N_25638,N_25936);
and U26952 (N_26952,N_25701,N_24096);
and U26953 (N_26953,N_25274,N_25802);
or U26954 (N_26954,N_25101,N_24108);
and U26955 (N_26955,N_24502,N_25623);
nor U26956 (N_26956,N_25816,N_24439);
nand U26957 (N_26957,N_25716,N_25544);
nand U26958 (N_26958,N_24797,N_25411);
nor U26959 (N_26959,N_25949,N_25565);
xor U26960 (N_26960,N_25404,N_25990);
xnor U26961 (N_26961,N_25451,N_24302);
xor U26962 (N_26962,N_24441,N_24599);
nor U26963 (N_26963,N_25375,N_25061);
or U26964 (N_26964,N_24115,N_25755);
and U26965 (N_26965,N_25923,N_25804);
nand U26966 (N_26966,N_25573,N_25592);
xnor U26967 (N_26967,N_25985,N_24400);
and U26968 (N_26968,N_24643,N_24396);
nand U26969 (N_26969,N_25156,N_24313);
nand U26970 (N_26970,N_25223,N_25639);
and U26971 (N_26971,N_24713,N_25060);
nand U26972 (N_26972,N_24555,N_24388);
nand U26973 (N_26973,N_24623,N_25759);
or U26974 (N_26974,N_25735,N_25798);
or U26975 (N_26975,N_24101,N_24854);
xnor U26976 (N_26976,N_25470,N_25414);
and U26977 (N_26977,N_24078,N_25687);
or U26978 (N_26978,N_24624,N_24181);
nand U26979 (N_26979,N_25113,N_25830);
or U26980 (N_26980,N_25435,N_24601);
nand U26981 (N_26981,N_25646,N_25958);
and U26982 (N_26982,N_24741,N_24933);
and U26983 (N_26983,N_24791,N_24515);
and U26984 (N_26984,N_25012,N_25355);
xor U26985 (N_26985,N_25253,N_24055);
nand U26986 (N_26986,N_25419,N_24062);
xnor U26987 (N_26987,N_25281,N_25054);
xnor U26988 (N_26988,N_25188,N_25655);
xor U26989 (N_26989,N_25030,N_24661);
nand U26990 (N_26990,N_24536,N_24714);
and U26991 (N_26991,N_25582,N_24197);
nand U26992 (N_26992,N_25540,N_24793);
xor U26993 (N_26993,N_24880,N_24415);
xnor U26994 (N_26994,N_25187,N_25665);
nor U26995 (N_26995,N_24775,N_24819);
or U26996 (N_26996,N_24241,N_24231);
xnor U26997 (N_26997,N_24385,N_24261);
or U26998 (N_26998,N_25085,N_24702);
xor U26999 (N_26999,N_24857,N_25133);
or U27000 (N_27000,N_24048,N_24644);
and U27001 (N_27001,N_24432,N_24807);
or U27002 (N_27002,N_24129,N_24008);
and U27003 (N_27003,N_25064,N_25345);
nand U27004 (N_27004,N_25578,N_25397);
nor U27005 (N_27005,N_25917,N_24617);
nor U27006 (N_27006,N_25949,N_25235);
and U27007 (N_27007,N_25562,N_24476);
and U27008 (N_27008,N_24170,N_25410);
and U27009 (N_27009,N_25401,N_24095);
nor U27010 (N_27010,N_25788,N_24979);
xor U27011 (N_27011,N_25921,N_24439);
nand U27012 (N_27012,N_25746,N_24040);
nor U27013 (N_27013,N_24804,N_24543);
and U27014 (N_27014,N_25759,N_24897);
nand U27015 (N_27015,N_25942,N_24165);
xnor U27016 (N_27016,N_25714,N_24607);
nand U27017 (N_27017,N_25739,N_25897);
xnor U27018 (N_27018,N_24943,N_24897);
nand U27019 (N_27019,N_25841,N_25611);
nor U27020 (N_27020,N_24282,N_24326);
nand U27021 (N_27021,N_25846,N_25006);
or U27022 (N_27022,N_25144,N_25308);
xor U27023 (N_27023,N_25472,N_25631);
and U27024 (N_27024,N_25395,N_25883);
nand U27025 (N_27025,N_25594,N_24853);
and U27026 (N_27026,N_24514,N_25317);
nor U27027 (N_27027,N_25999,N_24708);
xor U27028 (N_27028,N_25061,N_24794);
or U27029 (N_27029,N_24706,N_25494);
and U27030 (N_27030,N_24641,N_24339);
or U27031 (N_27031,N_25584,N_24495);
nor U27032 (N_27032,N_24565,N_25877);
nand U27033 (N_27033,N_25909,N_24563);
and U27034 (N_27034,N_25524,N_24958);
nor U27035 (N_27035,N_24774,N_24577);
nand U27036 (N_27036,N_25488,N_24158);
xnor U27037 (N_27037,N_25052,N_24306);
and U27038 (N_27038,N_24041,N_25416);
xor U27039 (N_27039,N_24068,N_24552);
nand U27040 (N_27040,N_24054,N_25274);
nand U27041 (N_27041,N_25440,N_25521);
and U27042 (N_27042,N_24548,N_25534);
nand U27043 (N_27043,N_25062,N_25381);
nand U27044 (N_27044,N_25420,N_25170);
and U27045 (N_27045,N_24612,N_24526);
xnor U27046 (N_27046,N_25294,N_24012);
nand U27047 (N_27047,N_25627,N_25542);
nor U27048 (N_27048,N_24879,N_25562);
xor U27049 (N_27049,N_24035,N_25424);
xnor U27050 (N_27050,N_24141,N_24648);
and U27051 (N_27051,N_25813,N_25103);
xnor U27052 (N_27052,N_24807,N_24033);
nor U27053 (N_27053,N_25099,N_25206);
xor U27054 (N_27054,N_25322,N_25614);
nand U27055 (N_27055,N_24276,N_24744);
and U27056 (N_27056,N_24414,N_25939);
nor U27057 (N_27057,N_24183,N_24241);
xnor U27058 (N_27058,N_24409,N_24197);
nor U27059 (N_27059,N_24277,N_24617);
nand U27060 (N_27060,N_25546,N_25726);
xnor U27061 (N_27061,N_25543,N_24034);
nor U27062 (N_27062,N_24230,N_24474);
or U27063 (N_27063,N_24093,N_24217);
and U27064 (N_27064,N_25931,N_24703);
nor U27065 (N_27065,N_25966,N_24751);
and U27066 (N_27066,N_24478,N_24405);
nand U27067 (N_27067,N_24506,N_25779);
and U27068 (N_27068,N_24688,N_25227);
and U27069 (N_27069,N_24823,N_25725);
nand U27070 (N_27070,N_25028,N_24721);
nor U27071 (N_27071,N_24138,N_24904);
nand U27072 (N_27072,N_25399,N_25875);
and U27073 (N_27073,N_24720,N_24936);
or U27074 (N_27074,N_25987,N_25237);
nor U27075 (N_27075,N_25373,N_25874);
or U27076 (N_27076,N_24204,N_25811);
nor U27077 (N_27077,N_24647,N_25771);
and U27078 (N_27078,N_25640,N_25975);
or U27079 (N_27079,N_24578,N_24069);
xnor U27080 (N_27080,N_24979,N_24007);
and U27081 (N_27081,N_24015,N_24775);
and U27082 (N_27082,N_25055,N_25780);
and U27083 (N_27083,N_24559,N_24310);
or U27084 (N_27084,N_25735,N_25822);
xor U27085 (N_27085,N_25795,N_24827);
or U27086 (N_27086,N_25165,N_25630);
xnor U27087 (N_27087,N_24969,N_24142);
xnor U27088 (N_27088,N_24886,N_25107);
or U27089 (N_27089,N_25323,N_24323);
and U27090 (N_27090,N_24892,N_24561);
and U27091 (N_27091,N_25589,N_24277);
and U27092 (N_27092,N_24454,N_24377);
nor U27093 (N_27093,N_25698,N_25080);
or U27094 (N_27094,N_25716,N_25514);
nor U27095 (N_27095,N_25469,N_25277);
nor U27096 (N_27096,N_25078,N_25994);
and U27097 (N_27097,N_25100,N_25897);
or U27098 (N_27098,N_24688,N_25613);
nand U27099 (N_27099,N_24771,N_24026);
or U27100 (N_27100,N_24695,N_25149);
or U27101 (N_27101,N_25849,N_25250);
and U27102 (N_27102,N_25812,N_24801);
or U27103 (N_27103,N_25452,N_25939);
xnor U27104 (N_27104,N_24414,N_24273);
xnor U27105 (N_27105,N_25925,N_25869);
nand U27106 (N_27106,N_24349,N_24288);
nor U27107 (N_27107,N_25389,N_24259);
xor U27108 (N_27108,N_24353,N_25307);
nand U27109 (N_27109,N_25344,N_25146);
xor U27110 (N_27110,N_24635,N_24768);
xor U27111 (N_27111,N_24972,N_25435);
nor U27112 (N_27112,N_25532,N_25563);
nor U27113 (N_27113,N_25772,N_25159);
or U27114 (N_27114,N_24876,N_25189);
or U27115 (N_27115,N_24325,N_24816);
xnor U27116 (N_27116,N_25331,N_25779);
nor U27117 (N_27117,N_25730,N_25797);
nand U27118 (N_27118,N_24406,N_24273);
nor U27119 (N_27119,N_24728,N_24450);
or U27120 (N_27120,N_25929,N_24604);
xor U27121 (N_27121,N_25047,N_25467);
xnor U27122 (N_27122,N_24970,N_25250);
or U27123 (N_27123,N_25011,N_24325);
or U27124 (N_27124,N_24412,N_24424);
nor U27125 (N_27125,N_24571,N_24385);
xor U27126 (N_27126,N_25614,N_25109);
nor U27127 (N_27127,N_24660,N_24754);
nand U27128 (N_27128,N_25001,N_24748);
nand U27129 (N_27129,N_24412,N_24987);
nand U27130 (N_27130,N_25432,N_24248);
nor U27131 (N_27131,N_25315,N_25531);
xor U27132 (N_27132,N_25329,N_25352);
nand U27133 (N_27133,N_24555,N_25710);
nand U27134 (N_27134,N_25686,N_25404);
and U27135 (N_27135,N_25691,N_24166);
and U27136 (N_27136,N_24283,N_25654);
nand U27137 (N_27137,N_24076,N_24157);
xnor U27138 (N_27138,N_24365,N_25192);
xor U27139 (N_27139,N_25982,N_25260);
or U27140 (N_27140,N_25072,N_24203);
xnor U27141 (N_27141,N_25892,N_25746);
nor U27142 (N_27142,N_25305,N_25684);
nor U27143 (N_27143,N_24691,N_25956);
and U27144 (N_27144,N_24624,N_24345);
nor U27145 (N_27145,N_24927,N_24849);
xnor U27146 (N_27146,N_24106,N_25779);
nand U27147 (N_27147,N_25743,N_25135);
nand U27148 (N_27148,N_25235,N_24342);
nor U27149 (N_27149,N_25594,N_24938);
nand U27150 (N_27150,N_25154,N_25078);
xnor U27151 (N_27151,N_25162,N_24275);
xor U27152 (N_27152,N_24798,N_25437);
or U27153 (N_27153,N_25492,N_25558);
or U27154 (N_27154,N_24657,N_24386);
or U27155 (N_27155,N_24793,N_24610);
nor U27156 (N_27156,N_25762,N_24864);
or U27157 (N_27157,N_24939,N_24525);
xnor U27158 (N_27158,N_25968,N_24432);
or U27159 (N_27159,N_24524,N_24903);
nor U27160 (N_27160,N_25337,N_25700);
nor U27161 (N_27161,N_24293,N_24890);
or U27162 (N_27162,N_24675,N_25822);
and U27163 (N_27163,N_25332,N_25506);
nor U27164 (N_27164,N_25167,N_25075);
xor U27165 (N_27165,N_25205,N_25332);
xor U27166 (N_27166,N_25919,N_25811);
and U27167 (N_27167,N_25042,N_25830);
nand U27168 (N_27168,N_25926,N_24413);
or U27169 (N_27169,N_25412,N_25889);
nor U27170 (N_27170,N_24941,N_24889);
nor U27171 (N_27171,N_25122,N_24655);
nor U27172 (N_27172,N_24835,N_25820);
nand U27173 (N_27173,N_24998,N_25201);
nor U27174 (N_27174,N_25519,N_24278);
nand U27175 (N_27175,N_24006,N_25842);
and U27176 (N_27176,N_24127,N_24969);
nand U27177 (N_27177,N_24138,N_24896);
or U27178 (N_27178,N_25219,N_25643);
nor U27179 (N_27179,N_25627,N_25693);
or U27180 (N_27180,N_24253,N_25294);
nand U27181 (N_27181,N_25251,N_25143);
nand U27182 (N_27182,N_24206,N_25639);
xnor U27183 (N_27183,N_25968,N_24469);
xnor U27184 (N_27184,N_25974,N_25655);
or U27185 (N_27185,N_24017,N_25613);
or U27186 (N_27186,N_25912,N_25505);
xnor U27187 (N_27187,N_24028,N_25269);
nor U27188 (N_27188,N_25640,N_25972);
xor U27189 (N_27189,N_24505,N_25912);
or U27190 (N_27190,N_25676,N_24130);
xor U27191 (N_27191,N_25750,N_24046);
nand U27192 (N_27192,N_25519,N_24221);
nor U27193 (N_27193,N_24130,N_25596);
nor U27194 (N_27194,N_24288,N_24025);
and U27195 (N_27195,N_24882,N_24146);
and U27196 (N_27196,N_25919,N_25653);
xor U27197 (N_27197,N_24446,N_24620);
or U27198 (N_27198,N_24918,N_24437);
or U27199 (N_27199,N_24948,N_24361);
xor U27200 (N_27200,N_24651,N_24449);
xor U27201 (N_27201,N_25829,N_25662);
and U27202 (N_27202,N_25347,N_25681);
nor U27203 (N_27203,N_25104,N_24041);
nand U27204 (N_27204,N_24882,N_25737);
nand U27205 (N_27205,N_25500,N_24923);
nor U27206 (N_27206,N_24111,N_24711);
and U27207 (N_27207,N_24564,N_25144);
and U27208 (N_27208,N_25824,N_24087);
or U27209 (N_27209,N_25628,N_24698);
and U27210 (N_27210,N_25911,N_25700);
nor U27211 (N_27211,N_25075,N_25640);
nand U27212 (N_27212,N_24924,N_24096);
or U27213 (N_27213,N_25683,N_24587);
and U27214 (N_27214,N_24107,N_25662);
nor U27215 (N_27215,N_25906,N_25411);
xor U27216 (N_27216,N_25097,N_25539);
nand U27217 (N_27217,N_25659,N_25305);
or U27218 (N_27218,N_25663,N_25993);
nor U27219 (N_27219,N_25744,N_25118);
nor U27220 (N_27220,N_24011,N_25950);
xor U27221 (N_27221,N_24338,N_24020);
nand U27222 (N_27222,N_24199,N_24332);
nand U27223 (N_27223,N_25467,N_24378);
xnor U27224 (N_27224,N_25892,N_25916);
and U27225 (N_27225,N_25777,N_24146);
or U27226 (N_27226,N_24073,N_24587);
and U27227 (N_27227,N_24015,N_24974);
nand U27228 (N_27228,N_24879,N_25929);
or U27229 (N_27229,N_25446,N_24536);
nand U27230 (N_27230,N_24549,N_25437);
xor U27231 (N_27231,N_24864,N_24585);
and U27232 (N_27232,N_25803,N_25614);
nand U27233 (N_27233,N_24295,N_24960);
and U27234 (N_27234,N_24754,N_24089);
or U27235 (N_27235,N_25867,N_24298);
nor U27236 (N_27236,N_25919,N_24562);
nor U27237 (N_27237,N_24801,N_24607);
nor U27238 (N_27238,N_25598,N_24143);
and U27239 (N_27239,N_24888,N_25140);
nor U27240 (N_27240,N_24819,N_24202);
or U27241 (N_27241,N_25838,N_25723);
or U27242 (N_27242,N_24568,N_24614);
nor U27243 (N_27243,N_24464,N_24463);
nor U27244 (N_27244,N_24377,N_24828);
or U27245 (N_27245,N_24935,N_24094);
xnor U27246 (N_27246,N_25944,N_24332);
nor U27247 (N_27247,N_24007,N_24183);
nor U27248 (N_27248,N_25227,N_24916);
nand U27249 (N_27249,N_24379,N_24646);
and U27250 (N_27250,N_25859,N_24533);
xor U27251 (N_27251,N_24958,N_24669);
nand U27252 (N_27252,N_24424,N_24390);
nand U27253 (N_27253,N_24762,N_25854);
or U27254 (N_27254,N_25548,N_25809);
and U27255 (N_27255,N_25907,N_24298);
xnor U27256 (N_27256,N_24268,N_24858);
and U27257 (N_27257,N_24000,N_25594);
nor U27258 (N_27258,N_24613,N_25410);
and U27259 (N_27259,N_25491,N_25537);
and U27260 (N_27260,N_24183,N_24619);
xnor U27261 (N_27261,N_25842,N_24290);
nand U27262 (N_27262,N_25463,N_25778);
or U27263 (N_27263,N_25554,N_24510);
or U27264 (N_27264,N_25389,N_25869);
nor U27265 (N_27265,N_25159,N_24907);
nand U27266 (N_27266,N_25863,N_24052);
nor U27267 (N_27267,N_24182,N_25281);
xor U27268 (N_27268,N_25017,N_24233);
or U27269 (N_27269,N_24531,N_25250);
and U27270 (N_27270,N_25250,N_25894);
and U27271 (N_27271,N_25984,N_25129);
and U27272 (N_27272,N_25691,N_25970);
nor U27273 (N_27273,N_24586,N_25747);
nor U27274 (N_27274,N_24984,N_25692);
xor U27275 (N_27275,N_24341,N_25572);
nor U27276 (N_27276,N_24353,N_25676);
nand U27277 (N_27277,N_25870,N_25165);
xor U27278 (N_27278,N_24724,N_24096);
nand U27279 (N_27279,N_25041,N_24053);
nor U27280 (N_27280,N_24191,N_24214);
or U27281 (N_27281,N_24742,N_25225);
or U27282 (N_27282,N_25441,N_25686);
nor U27283 (N_27283,N_25528,N_25062);
nor U27284 (N_27284,N_24848,N_25771);
xor U27285 (N_27285,N_25214,N_24070);
nor U27286 (N_27286,N_24501,N_24291);
nor U27287 (N_27287,N_24947,N_25922);
xnor U27288 (N_27288,N_24926,N_24451);
nand U27289 (N_27289,N_25079,N_25481);
xor U27290 (N_27290,N_24291,N_25420);
and U27291 (N_27291,N_25957,N_25595);
or U27292 (N_27292,N_25049,N_24993);
and U27293 (N_27293,N_25561,N_25763);
xnor U27294 (N_27294,N_24763,N_24271);
and U27295 (N_27295,N_25447,N_24689);
xnor U27296 (N_27296,N_24822,N_25778);
or U27297 (N_27297,N_25788,N_25835);
or U27298 (N_27298,N_25205,N_24905);
xnor U27299 (N_27299,N_25188,N_25636);
and U27300 (N_27300,N_24888,N_24565);
or U27301 (N_27301,N_24735,N_24828);
nor U27302 (N_27302,N_25915,N_24270);
or U27303 (N_27303,N_25765,N_24719);
nor U27304 (N_27304,N_24666,N_24541);
nand U27305 (N_27305,N_24411,N_25305);
nor U27306 (N_27306,N_25398,N_25712);
nor U27307 (N_27307,N_24855,N_24894);
xor U27308 (N_27308,N_24660,N_25187);
xnor U27309 (N_27309,N_24745,N_25685);
nand U27310 (N_27310,N_25949,N_25234);
nor U27311 (N_27311,N_25149,N_25109);
or U27312 (N_27312,N_25094,N_25723);
xnor U27313 (N_27313,N_24505,N_24433);
or U27314 (N_27314,N_25455,N_25843);
nand U27315 (N_27315,N_24219,N_25269);
or U27316 (N_27316,N_24088,N_24437);
or U27317 (N_27317,N_24966,N_24822);
nand U27318 (N_27318,N_24368,N_24701);
and U27319 (N_27319,N_25245,N_24092);
or U27320 (N_27320,N_25705,N_25506);
or U27321 (N_27321,N_25002,N_25564);
xor U27322 (N_27322,N_24385,N_24676);
nor U27323 (N_27323,N_24095,N_25774);
xnor U27324 (N_27324,N_24026,N_25035);
or U27325 (N_27325,N_24223,N_24724);
nor U27326 (N_27326,N_24803,N_25828);
and U27327 (N_27327,N_24491,N_25579);
and U27328 (N_27328,N_25393,N_24660);
or U27329 (N_27329,N_24049,N_24388);
and U27330 (N_27330,N_25823,N_24721);
or U27331 (N_27331,N_24481,N_24330);
and U27332 (N_27332,N_24702,N_25013);
xor U27333 (N_27333,N_25481,N_24468);
nor U27334 (N_27334,N_25313,N_24805);
and U27335 (N_27335,N_25669,N_25444);
nor U27336 (N_27336,N_24202,N_24660);
xnor U27337 (N_27337,N_25425,N_24392);
xor U27338 (N_27338,N_24864,N_25539);
nor U27339 (N_27339,N_24952,N_24751);
nand U27340 (N_27340,N_24290,N_25750);
nor U27341 (N_27341,N_25061,N_24435);
nor U27342 (N_27342,N_25066,N_24971);
nor U27343 (N_27343,N_25583,N_24898);
or U27344 (N_27344,N_24613,N_25889);
xor U27345 (N_27345,N_25960,N_24752);
nor U27346 (N_27346,N_24766,N_24029);
xor U27347 (N_27347,N_25944,N_24640);
nand U27348 (N_27348,N_25735,N_24924);
nand U27349 (N_27349,N_25958,N_25612);
nand U27350 (N_27350,N_25673,N_24386);
or U27351 (N_27351,N_25923,N_24305);
xor U27352 (N_27352,N_24709,N_25838);
xnor U27353 (N_27353,N_25024,N_24507);
or U27354 (N_27354,N_25928,N_25335);
nor U27355 (N_27355,N_25627,N_24640);
or U27356 (N_27356,N_24378,N_25491);
xor U27357 (N_27357,N_24821,N_24514);
or U27358 (N_27358,N_25992,N_24269);
and U27359 (N_27359,N_24384,N_25366);
and U27360 (N_27360,N_25775,N_25936);
nor U27361 (N_27361,N_24703,N_24002);
nor U27362 (N_27362,N_24036,N_25320);
nand U27363 (N_27363,N_25173,N_25177);
and U27364 (N_27364,N_24247,N_24697);
and U27365 (N_27365,N_25097,N_25821);
nor U27366 (N_27366,N_24941,N_24899);
nand U27367 (N_27367,N_24312,N_25218);
xnor U27368 (N_27368,N_25213,N_24337);
nand U27369 (N_27369,N_25559,N_25959);
or U27370 (N_27370,N_24079,N_24784);
or U27371 (N_27371,N_25815,N_24262);
nand U27372 (N_27372,N_24831,N_25235);
xnor U27373 (N_27373,N_25838,N_25268);
and U27374 (N_27374,N_25340,N_25514);
or U27375 (N_27375,N_24680,N_25026);
nor U27376 (N_27376,N_25510,N_25535);
nand U27377 (N_27377,N_24119,N_25109);
or U27378 (N_27378,N_25920,N_24028);
and U27379 (N_27379,N_25269,N_24959);
or U27380 (N_27380,N_24683,N_24495);
xor U27381 (N_27381,N_25772,N_25826);
and U27382 (N_27382,N_25284,N_24996);
or U27383 (N_27383,N_25207,N_25258);
xor U27384 (N_27384,N_25061,N_25037);
nand U27385 (N_27385,N_25729,N_24081);
xnor U27386 (N_27386,N_24314,N_25099);
or U27387 (N_27387,N_25191,N_25170);
nor U27388 (N_27388,N_25532,N_25836);
xnor U27389 (N_27389,N_24555,N_24883);
nand U27390 (N_27390,N_25648,N_24836);
or U27391 (N_27391,N_25484,N_25997);
xnor U27392 (N_27392,N_24971,N_25743);
or U27393 (N_27393,N_24908,N_24677);
nor U27394 (N_27394,N_25358,N_25331);
or U27395 (N_27395,N_24010,N_24746);
and U27396 (N_27396,N_25493,N_24073);
and U27397 (N_27397,N_24856,N_25455);
xnor U27398 (N_27398,N_25692,N_25952);
and U27399 (N_27399,N_24152,N_24863);
nor U27400 (N_27400,N_25260,N_24364);
nor U27401 (N_27401,N_24626,N_25996);
nor U27402 (N_27402,N_24075,N_25617);
or U27403 (N_27403,N_24786,N_25547);
xnor U27404 (N_27404,N_25006,N_25872);
nor U27405 (N_27405,N_25882,N_25078);
and U27406 (N_27406,N_25546,N_24560);
nand U27407 (N_27407,N_24622,N_24060);
nor U27408 (N_27408,N_25915,N_24505);
and U27409 (N_27409,N_24337,N_24134);
and U27410 (N_27410,N_25202,N_24126);
or U27411 (N_27411,N_25400,N_24478);
xnor U27412 (N_27412,N_24778,N_25094);
nand U27413 (N_27413,N_25979,N_25166);
nor U27414 (N_27414,N_24976,N_25711);
nor U27415 (N_27415,N_24112,N_24340);
nand U27416 (N_27416,N_25252,N_25242);
nor U27417 (N_27417,N_25506,N_24265);
nand U27418 (N_27418,N_25347,N_24429);
and U27419 (N_27419,N_25849,N_25199);
xnor U27420 (N_27420,N_25686,N_25770);
nand U27421 (N_27421,N_24643,N_24678);
or U27422 (N_27422,N_25561,N_25647);
or U27423 (N_27423,N_24214,N_24567);
nor U27424 (N_27424,N_25856,N_25489);
xor U27425 (N_27425,N_24224,N_24966);
or U27426 (N_27426,N_25797,N_25506);
nand U27427 (N_27427,N_25075,N_24139);
nor U27428 (N_27428,N_24058,N_24553);
or U27429 (N_27429,N_24339,N_25694);
nor U27430 (N_27430,N_25989,N_25232);
xor U27431 (N_27431,N_25567,N_24559);
xor U27432 (N_27432,N_24911,N_25138);
xnor U27433 (N_27433,N_25993,N_24026);
nand U27434 (N_27434,N_24204,N_24056);
nor U27435 (N_27435,N_24115,N_25710);
or U27436 (N_27436,N_24054,N_24481);
or U27437 (N_27437,N_25973,N_25440);
xnor U27438 (N_27438,N_24603,N_24332);
or U27439 (N_27439,N_24772,N_25855);
or U27440 (N_27440,N_25132,N_25477);
nand U27441 (N_27441,N_25861,N_25014);
and U27442 (N_27442,N_25636,N_25933);
or U27443 (N_27443,N_25038,N_25764);
or U27444 (N_27444,N_25676,N_24360);
or U27445 (N_27445,N_24620,N_24507);
nand U27446 (N_27446,N_25051,N_25327);
nor U27447 (N_27447,N_25189,N_24757);
xor U27448 (N_27448,N_24699,N_24743);
and U27449 (N_27449,N_24785,N_25536);
and U27450 (N_27450,N_24005,N_24881);
and U27451 (N_27451,N_24360,N_24717);
xnor U27452 (N_27452,N_25568,N_24074);
nor U27453 (N_27453,N_25831,N_25525);
or U27454 (N_27454,N_25757,N_24977);
nor U27455 (N_27455,N_25013,N_24049);
and U27456 (N_27456,N_24618,N_25753);
and U27457 (N_27457,N_25315,N_24249);
and U27458 (N_27458,N_25226,N_24789);
xnor U27459 (N_27459,N_25010,N_24221);
and U27460 (N_27460,N_24527,N_24441);
xnor U27461 (N_27461,N_25539,N_24887);
and U27462 (N_27462,N_25713,N_25457);
and U27463 (N_27463,N_24903,N_25147);
and U27464 (N_27464,N_25932,N_25385);
nand U27465 (N_27465,N_24165,N_25999);
and U27466 (N_27466,N_25357,N_25903);
xnor U27467 (N_27467,N_25578,N_25177);
nand U27468 (N_27468,N_25142,N_25336);
nand U27469 (N_27469,N_24396,N_24260);
and U27470 (N_27470,N_24743,N_24191);
nand U27471 (N_27471,N_25352,N_25596);
nand U27472 (N_27472,N_24299,N_25005);
and U27473 (N_27473,N_24316,N_25245);
nand U27474 (N_27474,N_24840,N_25105);
nand U27475 (N_27475,N_24778,N_24218);
and U27476 (N_27476,N_25469,N_25083);
or U27477 (N_27477,N_24947,N_24455);
nor U27478 (N_27478,N_24899,N_25627);
or U27479 (N_27479,N_25509,N_25931);
xnor U27480 (N_27480,N_24921,N_25142);
nand U27481 (N_27481,N_25100,N_24253);
nor U27482 (N_27482,N_25351,N_24427);
nor U27483 (N_27483,N_24061,N_24732);
nand U27484 (N_27484,N_25359,N_25293);
nand U27485 (N_27485,N_25935,N_25202);
nor U27486 (N_27486,N_24455,N_25359);
nor U27487 (N_27487,N_24875,N_24251);
nor U27488 (N_27488,N_25692,N_24887);
xnor U27489 (N_27489,N_25556,N_25263);
or U27490 (N_27490,N_25945,N_24954);
xnor U27491 (N_27491,N_25456,N_25361);
nand U27492 (N_27492,N_25709,N_24121);
or U27493 (N_27493,N_25925,N_24553);
and U27494 (N_27494,N_25788,N_24555);
or U27495 (N_27495,N_24980,N_25399);
xnor U27496 (N_27496,N_25093,N_24982);
nor U27497 (N_27497,N_25745,N_25349);
nor U27498 (N_27498,N_24881,N_25461);
or U27499 (N_27499,N_24302,N_24101);
and U27500 (N_27500,N_25738,N_25838);
or U27501 (N_27501,N_24346,N_25503);
or U27502 (N_27502,N_25977,N_25216);
nor U27503 (N_27503,N_24757,N_24349);
nor U27504 (N_27504,N_25749,N_24789);
nand U27505 (N_27505,N_25298,N_24111);
and U27506 (N_27506,N_25261,N_25262);
or U27507 (N_27507,N_25263,N_24527);
and U27508 (N_27508,N_25981,N_24080);
and U27509 (N_27509,N_25094,N_25740);
or U27510 (N_27510,N_25131,N_25287);
xor U27511 (N_27511,N_24399,N_25377);
or U27512 (N_27512,N_24302,N_25145);
and U27513 (N_27513,N_25320,N_24595);
xnor U27514 (N_27514,N_25979,N_25092);
nand U27515 (N_27515,N_25944,N_24688);
nor U27516 (N_27516,N_24931,N_25556);
nor U27517 (N_27517,N_25629,N_25373);
xor U27518 (N_27518,N_25721,N_25232);
nand U27519 (N_27519,N_24668,N_25129);
nand U27520 (N_27520,N_24083,N_24723);
nand U27521 (N_27521,N_24708,N_24964);
nand U27522 (N_27522,N_25156,N_24997);
and U27523 (N_27523,N_25008,N_24829);
and U27524 (N_27524,N_24755,N_25122);
and U27525 (N_27525,N_25983,N_24907);
xor U27526 (N_27526,N_25625,N_24530);
or U27527 (N_27527,N_25180,N_25728);
xor U27528 (N_27528,N_24230,N_25443);
nor U27529 (N_27529,N_25174,N_25698);
or U27530 (N_27530,N_25082,N_24045);
xor U27531 (N_27531,N_25782,N_24214);
nor U27532 (N_27532,N_24472,N_25255);
nor U27533 (N_27533,N_25714,N_25435);
nand U27534 (N_27534,N_24117,N_25413);
nor U27535 (N_27535,N_25887,N_25458);
nor U27536 (N_27536,N_25806,N_24320);
and U27537 (N_27537,N_24582,N_25600);
nor U27538 (N_27538,N_24925,N_25946);
and U27539 (N_27539,N_25569,N_24594);
nor U27540 (N_27540,N_24461,N_24785);
and U27541 (N_27541,N_24857,N_24582);
or U27542 (N_27542,N_25160,N_24470);
xor U27543 (N_27543,N_24320,N_25137);
or U27544 (N_27544,N_24423,N_24274);
nor U27545 (N_27545,N_25174,N_25480);
xnor U27546 (N_27546,N_24786,N_25102);
or U27547 (N_27547,N_24591,N_24255);
and U27548 (N_27548,N_25070,N_25287);
or U27549 (N_27549,N_24145,N_25038);
and U27550 (N_27550,N_24996,N_24217);
nor U27551 (N_27551,N_25868,N_24508);
nand U27552 (N_27552,N_24227,N_24453);
or U27553 (N_27553,N_25210,N_24657);
and U27554 (N_27554,N_25291,N_25854);
xor U27555 (N_27555,N_25179,N_24716);
nand U27556 (N_27556,N_25559,N_24022);
and U27557 (N_27557,N_24895,N_24632);
xnor U27558 (N_27558,N_24175,N_25483);
xor U27559 (N_27559,N_24217,N_25910);
xnor U27560 (N_27560,N_25280,N_25219);
or U27561 (N_27561,N_24044,N_25473);
nor U27562 (N_27562,N_25732,N_25798);
nand U27563 (N_27563,N_24445,N_24194);
nand U27564 (N_27564,N_24241,N_25690);
or U27565 (N_27565,N_25613,N_24177);
and U27566 (N_27566,N_25498,N_25869);
and U27567 (N_27567,N_25546,N_25970);
nand U27568 (N_27568,N_24830,N_25434);
or U27569 (N_27569,N_25213,N_25224);
or U27570 (N_27570,N_24358,N_24693);
nor U27571 (N_27571,N_24032,N_24163);
nand U27572 (N_27572,N_24982,N_25788);
xor U27573 (N_27573,N_25841,N_25891);
or U27574 (N_27574,N_25351,N_24739);
nand U27575 (N_27575,N_25635,N_25035);
and U27576 (N_27576,N_24447,N_25040);
or U27577 (N_27577,N_25436,N_25826);
nor U27578 (N_27578,N_25568,N_25314);
nand U27579 (N_27579,N_25361,N_25976);
and U27580 (N_27580,N_25378,N_25432);
nand U27581 (N_27581,N_25117,N_24597);
nor U27582 (N_27582,N_25280,N_24583);
nand U27583 (N_27583,N_25949,N_24346);
and U27584 (N_27584,N_25966,N_25213);
nor U27585 (N_27585,N_24932,N_25713);
nor U27586 (N_27586,N_25861,N_25381);
xor U27587 (N_27587,N_24087,N_24699);
xnor U27588 (N_27588,N_24296,N_24956);
or U27589 (N_27589,N_25417,N_25672);
and U27590 (N_27590,N_24046,N_25684);
and U27591 (N_27591,N_25827,N_24584);
nand U27592 (N_27592,N_24556,N_25248);
nor U27593 (N_27593,N_24496,N_24663);
or U27594 (N_27594,N_24417,N_25930);
xnor U27595 (N_27595,N_24044,N_25574);
nand U27596 (N_27596,N_25281,N_25187);
or U27597 (N_27597,N_24523,N_25155);
nor U27598 (N_27598,N_24509,N_24736);
or U27599 (N_27599,N_25728,N_25980);
nand U27600 (N_27600,N_25310,N_24043);
nand U27601 (N_27601,N_25499,N_24963);
or U27602 (N_27602,N_25967,N_25429);
nand U27603 (N_27603,N_25007,N_25714);
and U27604 (N_27604,N_24346,N_25207);
nor U27605 (N_27605,N_25693,N_25924);
nand U27606 (N_27606,N_24744,N_25702);
or U27607 (N_27607,N_25122,N_24516);
and U27608 (N_27608,N_25519,N_25066);
nor U27609 (N_27609,N_25816,N_25179);
xnor U27610 (N_27610,N_25716,N_24810);
nor U27611 (N_27611,N_25448,N_25794);
or U27612 (N_27612,N_24372,N_25064);
and U27613 (N_27613,N_25181,N_25157);
xor U27614 (N_27614,N_25910,N_24834);
xnor U27615 (N_27615,N_25970,N_24794);
or U27616 (N_27616,N_25308,N_25869);
or U27617 (N_27617,N_25456,N_25192);
xor U27618 (N_27618,N_25202,N_24074);
and U27619 (N_27619,N_25925,N_24644);
or U27620 (N_27620,N_24637,N_25344);
or U27621 (N_27621,N_25220,N_25109);
xor U27622 (N_27622,N_25714,N_25377);
or U27623 (N_27623,N_25782,N_24451);
nor U27624 (N_27624,N_24096,N_25047);
nor U27625 (N_27625,N_25358,N_25498);
nor U27626 (N_27626,N_24803,N_25217);
xnor U27627 (N_27627,N_24307,N_24100);
xor U27628 (N_27628,N_24404,N_24833);
nand U27629 (N_27629,N_25404,N_25053);
nand U27630 (N_27630,N_24768,N_24204);
or U27631 (N_27631,N_24024,N_25978);
nand U27632 (N_27632,N_24315,N_25886);
xor U27633 (N_27633,N_24701,N_24221);
or U27634 (N_27634,N_25190,N_25430);
nor U27635 (N_27635,N_24935,N_24192);
nand U27636 (N_27636,N_24586,N_24236);
and U27637 (N_27637,N_24827,N_24027);
or U27638 (N_27638,N_25342,N_25550);
and U27639 (N_27639,N_24942,N_24593);
nor U27640 (N_27640,N_25412,N_24427);
and U27641 (N_27641,N_24321,N_24026);
nor U27642 (N_27642,N_25136,N_25219);
or U27643 (N_27643,N_25242,N_25807);
nor U27644 (N_27644,N_25983,N_25428);
or U27645 (N_27645,N_24096,N_24638);
or U27646 (N_27646,N_24235,N_24570);
nand U27647 (N_27647,N_24194,N_25569);
nor U27648 (N_27648,N_24951,N_25038);
and U27649 (N_27649,N_25207,N_25931);
and U27650 (N_27650,N_24343,N_25429);
and U27651 (N_27651,N_24993,N_24661);
and U27652 (N_27652,N_24817,N_24440);
nor U27653 (N_27653,N_24505,N_25120);
or U27654 (N_27654,N_24117,N_25080);
or U27655 (N_27655,N_24461,N_25268);
and U27656 (N_27656,N_25831,N_25462);
or U27657 (N_27657,N_25772,N_24961);
or U27658 (N_27658,N_25581,N_25685);
xnor U27659 (N_27659,N_25759,N_25594);
nor U27660 (N_27660,N_25025,N_25405);
nand U27661 (N_27661,N_25622,N_24841);
or U27662 (N_27662,N_25157,N_24648);
nand U27663 (N_27663,N_24642,N_24762);
or U27664 (N_27664,N_25068,N_24869);
or U27665 (N_27665,N_24614,N_24709);
xnor U27666 (N_27666,N_25048,N_25286);
and U27667 (N_27667,N_25205,N_24411);
nor U27668 (N_27668,N_25544,N_24161);
and U27669 (N_27669,N_24989,N_24642);
nor U27670 (N_27670,N_24734,N_25783);
or U27671 (N_27671,N_24417,N_25180);
nor U27672 (N_27672,N_25199,N_25454);
and U27673 (N_27673,N_25693,N_25813);
xor U27674 (N_27674,N_25645,N_24437);
xor U27675 (N_27675,N_25951,N_24010);
or U27676 (N_27676,N_24412,N_24952);
xor U27677 (N_27677,N_25013,N_25630);
or U27678 (N_27678,N_24054,N_24727);
xnor U27679 (N_27679,N_25851,N_25817);
and U27680 (N_27680,N_24215,N_24328);
nor U27681 (N_27681,N_24027,N_25218);
nand U27682 (N_27682,N_25160,N_25888);
nand U27683 (N_27683,N_24411,N_25966);
xor U27684 (N_27684,N_25050,N_24149);
or U27685 (N_27685,N_25224,N_25873);
xor U27686 (N_27686,N_24619,N_25469);
xor U27687 (N_27687,N_24972,N_24776);
nand U27688 (N_27688,N_24422,N_25095);
xor U27689 (N_27689,N_24246,N_24722);
or U27690 (N_27690,N_25301,N_24303);
and U27691 (N_27691,N_25892,N_25223);
nand U27692 (N_27692,N_25712,N_24353);
nand U27693 (N_27693,N_24085,N_25874);
xnor U27694 (N_27694,N_24246,N_25662);
nor U27695 (N_27695,N_25612,N_24303);
or U27696 (N_27696,N_24068,N_24751);
nor U27697 (N_27697,N_25252,N_25304);
nor U27698 (N_27698,N_24787,N_25621);
xor U27699 (N_27699,N_24861,N_24300);
nor U27700 (N_27700,N_24474,N_25478);
xor U27701 (N_27701,N_24004,N_25666);
nor U27702 (N_27702,N_24400,N_24825);
nor U27703 (N_27703,N_25333,N_25144);
nand U27704 (N_27704,N_24723,N_24446);
nor U27705 (N_27705,N_25222,N_25651);
and U27706 (N_27706,N_25027,N_24764);
xnor U27707 (N_27707,N_24810,N_24228);
xnor U27708 (N_27708,N_24638,N_24422);
nand U27709 (N_27709,N_24083,N_24705);
nand U27710 (N_27710,N_24922,N_25277);
nand U27711 (N_27711,N_25150,N_24156);
nor U27712 (N_27712,N_24042,N_24924);
nand U27713 (N_27713,N_24898,N_25088);
xor U27714 (N_27714,N_24276,N_25861);
xor U27715 (N_27715,N_25807,N_24684);
or U27716 (N_27716,N_24462,N_25245);
xor U27717 (N_27717,N_24934,N_25798);
nor U27718 (N_27718,N_24821,N_24409);
xor U27719 (N_27719,N_24129,N_24107);
or U27720 (N_27720,N_25296,N_24245);
nand U27721 (N_27721,N_24441,N_24699);
and U27722 (N_27722,N_24895,N_25063);
xor U27723 (N_27723,N_24984,N_25580);
and U27724 (N_27724,N_24682,N_24958);
or U27725 (N_27725,N_24876,N_25516);
nor U27726 (N_27726,N_25087,N_24695);
nand U27727 (N_27727,N_24204,N_24879);
nor U27728 (N_27728,N_24184,N_24574);
and U27729 (N_27729,N_25026,N_24943);
or U27730 (N_27730,N_25877,N_24174);
or U27731 (N_27731,N_24720,N_24064);
nand U27732 (N_27732,N_24716,N_25417);
nor U27733 (N_27733,N_24637,N_25768);
xnor U27734 (N_27734,N_25005,N_24053);
or U27735 (N_27735,N_25649,N_25890);
nand U27736 (N_27736,N_24619,N_25392);
nand U27737 (N_27737,N_25202,N_24542);
xor U27738 (N_27738,N_24366,N_25549);
xnor U27739 (N_27739,N_24011,N_25661);
nand U27740 (N_27740,N_24635,N_25996);
or U27741 (N_27741,N_25138,N_24893);
nand U27742 (N_27742,N_25611,N_25238);
xnor U27743 (N_27743,N_25144,N_25638);
or U27744 (N_27744,N_24844,N_24720);
nor U27745 (N_27745,N_24385,N_24320);
xor U27746 (N_27746,N_24059,N_24890);
nand U27747 (N_27747,N_25902,N_24455);
nand U27748 (N_27748,N_24951,N_24247);
nand U27749 (N_27749,N_25307,N_25047);
and U27750 (N_27750,N_24530,N_25975);
xor U27751 (N_27751,N_25177,N_25655);
or U27752 (N_27752,N_24390,N_25291);
or U27753 (N_27753,N_25501,N_25202);
and U27754 (N_27754,N_24166,N_24909);
xnor U27755 (N_27755,N_25208,N_24293);
or U27756 (N_27756,N_24081,N_24980);
xor U27757 (N_27757,N_25927,N_25467);
xor U27758 (N_27758,N_25462,N_25429);
nor U27759 (N_27759,N_24319,N_25520);
and U27760 (N_27760,N_24142,N_25754);
and U27761 (N_27761,N_24017,N_25662);
xor U27762 (N_27762,N_25796,N_25319);
or U27763 (N_27763,N_24546,N_24422);
and U27764 (N_27764,N_25605,N_24968);
nor U27765 (N_27765,N_24908,N_25158);
nand U27766 (N_27766,N_24463,N_25498);
and U27767 (N_27767,N_24805,N_24962);
xnor U27768 (N_27768,N_25607,N_24041);
or U27769 (N_27769,N_25068,N_25010);
nor U27770 (N_27770,N_24161,N_25302);
or U27771 (N_27771,N_25179,N_25767);
nand U27772 (N_27772,N_24962,N_24270);
nor U27773 (N_27773,N_24985,N_24125);
xnor U27774 (N_27774,N_25204,N_25735);
or U27775 (N_27775,N_25304,N_24081);
nand U27776 (N_27776,N_24348,N_24515);
nor U27777 (N_27777,N_25410,N_25846);
nand U27778 (N_27778,N_24106,N_25562);
xnor U27779 (N_27779,N_25349,N_24466);
or U27780 (N_27780,N_25238,N_25242);
nand U27781 (N_27781,N_24349,N_25796);
nor U27782 (N_27782,N_25223,N_25585);
and U27783 (N_27783,N_24648,N_24723);
nand U27784 (N_27784,N_25998,N_24549);
and U27785 (N_27785,N_24649,N_25856);
xnor U27786 (N_27786,N_24220,N_24904);
and U27787 (N_27787,N_24643,N_25834);
or U27788 (N_27788,N_24607,N_25978);
and U27789 (N_27789,N_24278,N_24002);
or U27790 (N_27790,N_25689,N_24982);
and U27791 (N_27791,N_24755,N_25936);
or U27792 (N_27792,N_24083,N_24553);
nor U27793 (N_27793,N_25223,N_24680);
and U27794 (N_27794,N_25024,N_24078);
xnor U27795 (N_27795,N_24390,N_25831);
nor U27796 (N_27796,N_25793,N_24678);
and U27797 (N_27797,N_25590,N_25244);
xor U27798 (N_27798,N_24894,N_25330);
nor U27799 (N_27799,N_24617,N_24492);
or U27800 (N_27800,N_25037,N_25414);
nand U27801 (N_27801,N_24610,N_24192);
nand U27802 (N_27802,N_24972,N_24557);
nor U27803 (N_27803,N_25681,N_24843);
nand U27804 (N_27804,N_24166,N_24423);
xor U27805 (N_27805,N_24220,N_25886);
or U27806 (N_27806,N_24753,N_25052);
or U27807 (N_27807,N_24392,N_24429);
or U27808 (N_27808,N_25720,N_24165);
or U27809 (N_27809,N_25752,N_25600);
xor U27810 (N_27810,N_25465,N_25463);
nand U27811 (N_27811,N_25951,N_25828);
xor U27812 (N_27812,N_24268,N_25039);
or U27813 (N_27813,N_24056,N_25236);
and U27814 (N_27814,N_25411,N_24191);
and U27815 (N_27815,N_25547,N_25208);
nor U27816 (N_27816,N_25929,N_24588);
nand U27817 (N_27817,N_24431,N_25624);
or U27818 (N_27818,N_25465,N_24227);
or U27819 (N_27819,N_24609,N_24727);
or U27820 (N_27820,N_24739,N_24992);
xnor U27821 (N_27821,N_25089,N_25406);
and U27822 (N_27822,N_25061,N_24115);
or U27823 (N_27823,N_24352,N_24311);
nor U27824 (N_27824,N_24411,N_25324);
xnor U27825 (N_27825,N_24553,N_25976);
xor U27826 (N_27826,N_25894,N_24898);
and U27827 (N_27827,N_24677,N_25663);
and U27828 (N_27828,N_24397,N_24182);
and U27829 (N_27829,N_25664,N_25937);
nor U27830 (N_27830,N_24063,N_24244);
and U27831 (N_27831,N_24311,N_24039);
nand U27832 (N_27832,N_25167,N_25573);
nand U27833 (N_27833,N_25108,N_24918);
nand U27834 (N_27834,N_25237,N_25458);
and U27835 (N_27835,N_24652,N_24842);
and U27836 (N_27836,N_24014,N_24614);
nand U27837 (N_27837,N_24160,N_25885);
nor U27838 (N_27838,N_25811,N_25086);
nor U27839 (N_27839,N_25132,N_24532);
xnor U27840 (N_27840,N_25300,N_24444);
nor U27841 (N_27841,N_25137,N_24491);
and U27842 (N_27842,N_24504,N_25773);
nor U27843 (N_27843,N_24315,N_25977);
or U27844 (N_27844,N_25623,N_24017);
xnor U27845 (N_27845,N_24909,N_25346);
or U27846 (N_27846,N_24407,N_25163);
or U27847 (N_27847,N_25306,N_25288);
and U27848 (N_27848,N_25102,N_25150);
nor U27849 (N_27849,N_25562,N_25340);
and U27850 (N_27850,N_24121,N_25762);
or U27851 (N_27851,N_24193,N_24620);
or U27852 (N_27852,N_24201,N_24150);
nand U27853 (N_27853,N_25634,N_24289);
xnor U27854 (N_27854,N_25657,N_25365);
xnor U27855 (N_27855,N_24165,N_25793);
and U27856 (N_27856,N_25252,N_24630);
xor U27857 (N_27857,N_25050,N_25798);
and U27858 (N_27858,N_25408,N_25610);
or U27859 (N_27859,N_24455,N_25832);
and U27860 (N_27860,N_24849,N_25495);
xnor U27861 (N_27861,N_25940,N_25819);
nor U27862 (N_27862,N_25523,N_25498);
xnor U27863 (N_27863,N_24370,N_25071);
xnor U27864 (N_27864,N_24487,N_25874);
xnor U27865 (N_27865,N_24221,N_25230);
and U27866 (N_27866,N_25338,N_24322);
nor U27867 (N_27867,N_25135,N_24927);
and U27868 (N_27868,N_24083,N_25945);
xnor U27869 (N_27869,N_24012,N_24045);
or U27870 (N_27870,N_24704,N_24870);
and U27871 (N_27871,N_24095,N_24862);
xnor U27872 (N_27872,N_25050,N_25232);
and U27873 (N_27873,N_25151,N_25152);
nor U27874 (N_27874,N_24191,N_24696);
or U27875 (N_27875,N_25770,N_25654);
xnor U27876 (N_27876,N_24826,N_24311);
nor U27877 (N_27877,N_25098,N_25031);
and U27878 (N_27878,N_25879,N_24087);
xnor U27879 (N_27879,N_24751,N_24741);
or U27880 (N_27880,N_25823,N_25942);
xor U27881 (N_27881,N_24899,N_25815);
nor U27882 (N_27882,N_25891,N_25924);
and U27883 (N_27883,N_24301,N_24308);
xnor U27884 (N_27884,N_25976,N_25155);
xor U27885 (N_27885,N_25555,N_24830);
or U27886 (N_27886,N_24715,N_25533);
xor U27887 (N_27887,N_25423,N_24928);
xnor U27888 (N_27888,N_24421,N_24122);
xor U27889 (N_27889,N_24382,N_25697);
nor U27890 (N_27890,N_25726,N_25288);
nand U27891 (N_27891,N_24053,N_24356);
nor U27892 (N_27892,N_25287,N_24033);
xnor U27893 (N_27893,N_25722,N_24033);
xnor U27894 (N_27894,N_25586,N_25138);
nor U27895 (N_27895,N_25474,N_25891);
nand U27896 (N_27896,N_25512,N_24292);
nor U27897 (N_27897,N_24859,N_25883);
or U27898 (N_27898,N_25222,N_25919);
xor U27899 (N_27899,N_24201,N_24359);
or U27900 (N_27900,N_24583,N_24077);
xor U27901 (N_27901,N_25018,N_25915);
or U27902 (N_27902,N_25348,N_25534);
nand U27903 (N_27903,N_24972,N_25193);
xnor U27904 (N_27904,N_25164,N_24588);
nor U27905 (N_27905,N_24326,N_25324);
and U27906 (N_27906,N_25339,N_25750);
or U27907 (N_27907,N_25449,N_25119);
and U27908 (N_27908,N_25953,N_25647);
and U27909 (N_27909,N_25954,N_24148);
or U27910 (N_27910,N_24599,N_24367);
xnor U27911 (N_27911,N_25757,N_24483);
and U27912 (N_27912,N_25007,N_25385);
and U27913 (N_27913,N_24334,N_25787);
or U27914 (N_27914,N_24877,N_24861);
xnor U27915 (N_27915,N_25220,N_25970);
or U27916 (N_27916,N_24209,N_25943);
and U27917 (N_27917,N_24561,N_25955);
and U27918 (N_27918,N_25001,N_25174);
and U27919 (N_27919,N_25386,N_25709);
and U27920 (N_27920,N_25567,N_25610);
or U27921 (N_27921,N_25196,N_25195);
nor U27922 (N_27922,N_25974,N_24471);
nand U27923 (N_27923,N_24556,N_24577);
xnor U27924 (N_27924,N_24480,N_24453);
or U27925 (N_27925,N_25205,N_24031);
and U27926 (N_27926,N_25493,N_24471);
and U27927 (N_27927,N_25942,N_24359);
and U27928 (N_27928,N_24890,N_24211);
nor U27929 (N_27929,N_25080,N_24538);
and U27930 (N_27930,N_24651,N_24225);
nand U27931 (N_27931,N_25412,N_24941);
and U27932 (N_27932,N_24315,N_24350);
or U27933 (N_27933,N_25206,N_24556);
xnor U27934 (N_27934,N_25704,N_25573);
or U27935 (N_27935,N_24518,N_24985);
or U27936 (N_27936,N_24527,N_25260);
nand U27937 (N_27937,N_24379,N_25956);
and U27938 (N_27938,N_24513,N_24795);
and U27939 (N_27939,N_24911,N_24354);
or U27940 (N_27940,N_25369,N_25272);
xor U27941 (N_27941,N_25887,N_24216);
xor U27942 (N_27942,N_24400,N_24163);
or U27943 (N_27943,N_24349,N_25793);
nor U27944 (N_27944,N_25647,N_25584);
xor U27945 (N_27945,N_25428,N_24396);
xnor U27946 (N_27946,N_24324,N_25660);
xnor U27947 (N_27947,N_25085,N_24635);
or U27948 (N_27948,N_25895,N_25569);
nor U27949 (N_27949,N_24036,N_25227);
and U27950 (N_27950,N_25865,N_25337);
nor U27951 (N_27951,N_24278,N_24672);
or U27952 (N_27952,N_25695,N_25418);
or U27953 (N_27953,N_24797,N_24338);
nand U27954 (N_27954,N_25347,N_25183);
nor U27955 (N_27955,N_24983,N_24788);
and U27956 (N_27956,N_25051,N_24858);
nor U27957 (N_27957,N_24769,N_25999);
xnor U27958 (N_27958,N_25726,N_24968);
nand U27959 (N_27959,N_25620,N_24479);
nand U27960 (N_27960,N_24277,N_24751);
nand U27961 (N_27961,N_25872,N_25797);
and U27962 (N_27962,N_25389,N_25404);
xor U27963 (N_27963,N_25863,N_25101);
or U27964 (N_27964,N_25131,N_25055);
and U27965 (N_27965,N_24342,N_24336);
and U27966 (N_27966,N_25146,N_25362);
nor U27967 (N_27967,N_24835,N_24147);
nor U27968 (N_27968,N_25294,N_24043);
and U27969 (N_27969,N_24404,N_25357);
nand U27970 (N_27970,N_25375,N_24990);
xor U27971 (N_27971,N_25252,N_24240);
and U27972 (N_27972,N_24506,N_25131);
or U27973 (N_27973,N_25960,N_25214);
and U27974 (N_27974,N_24071,N_25087);
xor U27975 (N_27975,N_24892,N_25103);
nand U27976 (N_27976,N_25568,N_24108);
and U27977 (N_27977,N_24409,N_24030);
or U27978 (N_27978,N_24078,N_24346);
nor U27979 (N_27979,N_25266,N_24681);
xor U27980 (N_27980,N_24741,N_24299);
or U27981 (N_27981,N_24111,N_25340);
xnor U27982 (N_27982,N_25753,N_25583);
and U27983 (N_27983,N_24020,N_24536);
nand U27984 (N_27984,N_24273,N_25462);
nand U27985 (N_27985,N_25451,N_24289);
and U27986 (N_27986,N_25655,N_24472);
or U27987 (N_27987,N_25966,N_25536);
xor U27988 (N_27988,N_24995,N_24411);
or U27989 (N_27989,N_25082,N_25444);
nor U27990 (N_27990,N_24497,N_24865);
xor U27991 (N_27991,N_24526,N_24405);
nor U27992 (N_27992,N_24301,N_25680);
nand U27993 (N_27993,N_24686,N_25442);
nor U27994 (N_27994,N_25347,N_24392);
xor U27995 (N_27995,N_25104,N_24125);
xnor U27996 (N_27996,N_24304,N_24404);
or U27997 (N_27997,N_25952,N_25385);
nor U27998 (N_27998,N_25742,N_25045);
nand U27999 (N_27999,N_24421,N_24153);
nor U28000 (N_28000,N_26112,N_26709);
and U28001 (N_28001,N_27028,N_26947);
nor U28002 (N_28002,N_26756,N_27661);
nor U28003 (N_28003,N_26613,N_26820);
xor U28004 (N_28004,N_26462,N_27836);
and U28005 (N_28005,N_27831,N_26385);
nand U28006 (N_28006,N_26910,N_26353);
nand U28007 (N_28007,N_26582,N_27552);
and U28008 (N_28008,N_27789,N_27585);
nor U28009 (N_28009,N_27262,N_27628);
xnor U28010 (N_28010,N_27485,N_26817);
nand U28011 (N_28011,N_26030,N_27543);
nor U28012 (N_28012,N_27156,N_26854);
nand U28013 (N_28013,N_27581,N_27927);
or U28014 (N_28014,N_27302,N_27623);
or U28015 (N_28015,N_27551,N_26898);
nor U28016 (N_28016,N_26607,N_26453);
nor U28017 (N_28017,N_26873,N_27377);
xor U28018 (N_28018,N_26968,N_27700);
and U28019 (N_28019,N_26032,N_27645);
nor U28020 (N_28020,N_26598,N_27697);
and U28021 (N_28021,N_27422,N_27358);
nor U28022 (N_28022,N_27991,N_26215);
nor U28023 (N_28023,N_26704,N_27801);
or U28024 (N_28024,N_27383,N_27699);
nor U28025 (N_28025,N_27722,N_27056);
or U28026 (N_28026,N_27703,N_27394);
nand U28027 (N_28027,N_26605,N_26442);
nor U28028 (N_28028,N_27154,N_27362);
and U28029 (N_28029,N_26864,N_27388);
xor U28030 (N_28030,N_27077,N_26740);
nand U28031 (N_28031,N_26401,N_27178);
nor U28032 (N_28032,N_26714,N_27225);
nor U28033 (N_28033,N_26373,N_27640);
and U28034 (N_28034,N_26993,N_27355);
nor U28035 (N_28035,N_27762,N_27487);
and U28036 (N_28036,N_26603,N_26071);
nand U28037 (N_28037,N_27557,N_26339);
or U28038 (N_28038,N_26805,N_27881);
nor U28039 (N_28039,N_26166,N_26936);
nand U28040 (N_28040,N_27117,N_26776);
or U28041 (N_28041,N_27716,N_27080);
xor U28042 (N_28042,N_27042,N_27431);
or U28043 (N_28043,N_26037,N_27942);
and U28044 (N_28044,N_26865,N_27065);
xnor U28045 (N_28045,N_27064,N_26682);
nor U28046 (N_28046,N_27198,N_26432);
or U28047 (N_28047,N_27257,N_27228);
and U28048 (N_28048,N_26137,N_27610);
nor U28049 (N_28049,N_27639,N_27286);
nand U28050 (N_28050,N_27499,N_26945);
and U28051 (N_28051,N_27600,N_27146);
and U28052 (N_28052,N_27033,N_26702);
nor U28053 (N_28053,N_27644,N_27872);
and U28054 (N_28054,N_27111,N_27818);
nand U28055 (N_28055,N_27315,N_27773);
and U28056 (N_28056,N_26955,N_27405);
nor U28057 (N_28057,N_27994,N_26892);
nor U28058 (N_28058,N_26862,N_27239);
or U28059 (N_28059,N_27951,N_26349);
and U28060 (N_28060,N_27316,N_27312);
nor U28061 (N_28061,N_26157,N_27233);
and U28062 (N_28062,N_27106,N_26430);
and U28063 (N_28063,N_27588,N_26627);
and U28064 (N_28064,N_26930,N_27290);
or U28065 (N_28065,N_26724,N_27729);
nor U28066 (N_28066,N_27051,N_27322);
nand U28067 (N_28067,N_26122,N_27861);
nand U28068 (N_28068,N_27530,N_27977);
xor U28069 (N_28069,N_27775,N_27896);
and U28070 (N_28070,N_26590,N_27674);
nand U28071 (N_28071,N_27211,N_27886);
xor U28072 (N_28072,N_27569,N_26158);
or U28073 (N_28073,N_27075,N_26979);
or U28074 (N_28074,N_27741,N_26515);
nor U28075 (N_28075,N_27240,N_26549);
nor U28076 (N_28076,N_27196,N_26050);
nor U28077 (N_28077,N_27424,N_27113);
or U28078 (N_28078,N_27219,N_26725);
or U28079 (N_28079,N_26450,N_26942);
nor U28080 (N_28080,N_27010,N_27948);
and U28081 (N_28081,N_27331,N_26085);
xnor U28082 (N_28082,N_26665,N_26038);
nand U28083 (N_28083,N_26591,N_26212);
xnor U28084 (N_28084,N_27093,N_27371);
and U28085 (N_28085,N_27002,N_26683);
nor U28086 (N_28086,N_27491,N_27107);
nand U28087 (N_28087,N_27577,N_26490);
or U28088 (N_28088,N_26147,N_27918);
nor U28089 (N_28089,N_26036,N_26736);
xnor U28090 (N_28090,N_26352,N_27978);
xnor U28091 (N_28091,N_27755,N_26739);
nand U28092 (N_28092,N_26060,N_27528);
nand U28093 (N_28093,N_26668,N_27996);
and U28094 (N_28094,N_27205,N_26983);
xor U28095 (N_28095,N_26247,N_26843);
xor U28096 (N_28096,N_26869,N_27790);
xor U28097 (N_28097,N_26966,N_27335);
or U28098 (N_28098,N_27840,N_26513);
and U28099 (N_28099,N_27612,N_26960);
xor U28100 (N_28100,N_27970,N_26210);
nand U28101 (N_28101,N_26642,N_27008);
and U28102 (N_28102,N_26509,N_26584);
and U28103 (N_28103,N_26568,N_26191);
nor U28104 (N_28104,N_27369,N_27378);
nand U28105 (N_28105,N_26413,N_27309);
and U28106 (N_28106,N_26496,N_27791);
xor U28107 (N_28107,N_27462,N_26316);
xnor U28108 (N_28108,N_27475,N_26118);
or U28109 (N_28109,N_26408,N_26379);
and U28110 (N_28110,N_26610,N_26132);
and U28111 (N_28111,N_27698,N_26588);
nor U28112 (N_28112,N_27586,N_26559);
nor U28113 (N_28113,N_26715,N_26227);
nor U28114 (N_28114,N_26001,N_27825);
nor U28115 (N_28115,N_27745,N_26656);
and U28116 (N_28116,N_27438,N_26325);
and U28117 (N_28117,N_27862,N_26974);
nand U28118 (N_28118,N_27546,N_26851);
and U28119 (N_28119,N_26188,N_26802);
xor U28120 (N_28120,N_26689,N_26129);
or U28121 (N_28121,N_26197,N_27140);
nor U28122 (N_28122,N_27320,N_27602);
nand U28123 (N_28123,N_27120,N_26505);
or U28124 (N_28124,N_26972,N_26186);
nor U28125 (N_28125,N_26812,N_26622);
or U28126 (N_28126,N_27737,N_27165);
and U28127 (N_28127,N_26666,N_27838);
nand U28128 (N_28128,N_27769,N_27934);
nand U28129 (N_28129,N_26618,N_27134);
and U28130 (N_28130,N_26722,N_27772);
nor U28131 (N_28131,N_26435,N_26102);
or U28132 (N_28132,N_27964,N_26411);
xor U28133 (N_28133,N_27631,N_26612);
or U28134 (N_28134,N_26951,N_26276);
nor U28135 (N_28135,N_26289,N_26005);
and U28136 (N_28136,N_26209,N_27969);
nand U28137 (N_28137,N_26806,N_26954);
and U28138 (N_28138,N_27007,N_26346);
or U28139 (N_28139,N_27877,N_26192);
nor U28140 (N_28140,N_26141,N_26548);
nor U28141 (N_28141,N_26971,N_26069);
nand U28142 (N_28142,N_26818,N_26914);
xor U28143 (N_28143,N_27158,N_27516);
nand U28144 (N_28144,N_26597,N_26143);
xnor U28145 (N_28145,N_27784,N_27556);
nor U28146 (N_28146,N_27988,N_26285);
or U28147 (N_28147,N_26405,N_26308);
nor U28148 (N_28148,N_27465,N_26981);
xnor U28149 (N_28149,N_27962,N_26861);
and U28150 (N_28150,N_26008,N_27867);
nor U28151 (N_28151,N_27199,N_26671);
or U28152 (N_28152,N_27024,N_27856);
or U28153 (N_28153,N_26348,N_27005);
nor U28154 (N_28154,N_27453,N_27795);
or U28155 (N_28155,N_27116,N_27186);
nand U28156 (N_28156,N_27490,N_26727);
xor U28157 (N_28157,N_27448,N_27809);
nand U28158 (N_28158,N_27323,N_27232);
and U28159 (N_28159,N_27802,N_26090);
and U28160 (N_28160,N_27555,N_26524);
nor U28161 (N_28161,N_26335,N_26216);
xnor U28162 (N_28162,N_27899,N_27884);
nor U28163 (N_28163,N_27019,N_26378);
nor U28164 (N_28164,N_27376,N_26772);
and U28165 (N_28165,N_27882,N_27283);
xnor U28166 (N_28166,N_27293,N_26655);
and U28167 (N_28167,N_26204,N_26767);
xnor U28168 (N_28168,N_26437,N_27126);
nand U28169 (N_28169,N_26646,N_26661);
nor U28170 (N_28170,N_27979,N_26376);
xor U28171 (N_28171,N_26048,N_26305);
nor U28172 (N_28172,N_26717,N_27253);
xor U28173 (N_28173,N_26123,N_27379);
nand U28174 (N_28174,N_27003,N_26636);
xor U28175 (N_28175,N_26355,N_27169);
xnor U28176 (N_28176,N_27452,N_27786);
or U28177 (N_28177,N_27364,N_27161);
nor U28178 (N_28178,N_26784,N_27246);
or U28179 (N_28179,N_26110,N_27573);
nand U28180 (N_28180,N_26659,N_27777);
or U28181 (N_28181,N_27354,N_26798);
nor U28182 (N_28182,N_26878,N_27252);
xor U28183 (N_28183,N_26986,N_26575);
xnor U28184 (N_28184,N_27895,N_26708);
xnor U28185 (N_28185,N_27619,N_26630);
xor U28186 (N_28186,N_27396,N_26572);
nor U28187 (N_28187,N_27835,N_27855);
xnor U28188 (N_28188,N_26501,N_27039);
xor U28189 (N_28189,N_27606,N_26741);
nand U28190 (N_28190,N_26891,N_27869);
xnor U28191 (N_28191,N_27811,N_27193);
and U28192 (N_28192,N_27373,N_26231);
or U28193 (N_28193,N_26558,N_26078);
nor U28194 (N_28194,N_27300,N_27160);
nor U28195 (N_28195,N_26237,N_26456);
xor U28196 (N_28196,N_26587,N_27256);
xnor U28197 (N_28197,N_26097,N_27981);
and U28198 (N_28198,N_26043,N_27821);
xnor U28199 (N_28199,N_27101,N_27348);
or U28200 (N_28200,N_27724,N_26211);
and U28201 (N_28201,N_27764,N_26425);
nor U28202 (N_28202,N_27368,N_27215);
and U28203 (N_28203,N_27000,N_26059);
xnor U28204 (N_28204,N_26536,N_27030);
xnor U28205 (N_28205,N_27921,N_27036);
nand U28206 (N_28206,N_26713,N_26274);
and U28207 (N_28207,N_27616,N_26902);
nor U28208 (N_28208,N_27766,N_27542);
xor U28209 (N_28209,N_27952,N_27743);
nor U28210 (N_28210,N_27672,N_27128);
nor U28211 (N_28211,N_27758,N_26662);
and U28212 (N_28212,N_26874,N_26039);
nand U28213 (N_28213,N_26358,N_26912);
xor U28214 (N_28214,N_27421,N_26286);
or U28215 (N_28215,N_26354,N_27780);
and U28216 (N_28216,N_26466,N_27251);
or U28217 (N_28217,N_26415,N_26364);
and U28218 (N_28218,N_26821,N_27511);
and U28219 (N_28219,N_26270,N_27909);
or U28220 (N_28220,N_27541,N_27386);
nor U28221 (N_28221,N_26222,N_27387);
and U28222 (N_28222,N_27580,N_27400);
nor U28223 (N_28223,N_27014,N_27274);
or U28224 (N_28224,N_26206,N_26347);
or U28225 (N_28225,N_26007,N_26272);
nand U28226 (N_28226,N_26519,N_27812);
xnor U28227 (N_28227,N_27903,N_26243);
and U28228 (N_28228,N_27409,N_27187);
nand U28229 (N_28229,N_26620,N_26748);
and U28230 (N_28230,N_26952,N_26221);
xor U28231 (N_28231,N_26478,N_27598);
and U28232 (N_28232,N_27912,N_27695);
or U28233 (N_28233,N_26850,N_26455);
xnor U28234 (N_28234,N_27630,N_27566);
or U28235 (N_28235,N_27850,N_26919);
nor U28236 (N_28236,N_26135,N_27168);
xor U28237 (N_28237,N_27968,N_26755);
and U28238 (N_28238,N_27870,N_27365);
nor U28239 (N_28239,N_26762,N_27353);
nand U28240 (N_28240,N_27279,N_27684);
xnor U28241 (N_28241,N_27844,N_26908);
and U28242 (N_28242,N_27059,N_27428);
nor U28243 (N_28243,N_26583,N_27596);
xor U28244 (N_28244,N_26449,N_27078);
nor U28245 (N_28245,N_26336,N_26542);
xor U28246 (N_28246,N_26320,N_27306);
and U28247 (N_28247,N_27446,N_26306);
and U28248 (N_28248,N_27311,N_27534);
nor U28249 (N_28249,N_27461,N_27824);
and U28250 (N_28250,N_27793,N_27478);
xor U28251 (N_28251,N_26329,N_27174);
nor U28252 (N_28252,N_27998,N_26465);
and U28253 (N_28253,N_27670,N_26079);
xnor U28254 (N_28254,N_27052,N_27175);
xnor U28255 (N_28255,N_27009,N_26367);
nor U28256 (N_28256,N_26387,N_26905);
xnor U28257 (N_28257,N_27349,N_26394);
xnor U28258 (N_28258,N_26273,N_26626);
xor U28259 (N_28259,N_27691,N_27384);
nor U28260 (N_28260,N_27562,N_26390);
and U28261 (N_28261,N_26481,N_27627);
or U28262 (N_28262,N_26026,N_26980);
and U28263 (N_28263,N_26075,N_27561);
and U28264 (N_28264,N_27164,N_26365);
nand U28265 (N_28265,N_27121,N_26463);
or U28266 (N_28266,N_26239,N_26804);
or U28267 (N_28267,N_27216,N_27264);
and U28268 (N_28268,N_27820,N_27742);
nor U28269 (N_28269,N_27166,N_26021);
nand U28270 (N_28270,N_27294,N_26922);
xor U28271 (N_28271,N_26970,N_26538);
nor U28272 (N_28272,N_27518,N_27813);
and U28273 (N_28273,N_26235,N_27982);
or U28274 (N_28274,N_27454,N_26125);
xor U28275 (N_28275,N_26040,N_27292);
nor U28276 (N_28276,N_26576,N_26410);
or U28277 (N_28277,N_27271,N_27897);
and U28278 (N_28278,N_26091,N_26560);
nor U28279 (N_28279,N_27894,N_27040);
nand U28280 (N_28280,N_26600,N_27723);
xnor U28281 (N_28281,N_26863,N_26606);
nand U28282 (N_28282,N_27613,N_26637);
and U28283 (N_28283,N_26690,N_26380);
and U28284 (N_28284,N_27269,N_26396);
and U28285 (N_28285,N_27571,N_27129);
nand U28286 (N_28286,N_26472,N_27004);
or U28287 (N_28287,N_26976,N_27849);
and U28288 (N_28288,N_27221,N_26228);
nand U28289 (N_28289,N_26546,N_26096);
xnor U28290 (N_28290,N_27356,N_27920);
and U28291 (N_28291,N_26628,N_27427);
and U28292 (N_28292,N_26024,N_26962);
xor U28293 (N_28293,N_27466,N_27436);
or U28294 (N_28294,N_27984,N_27133);
xnor U28295 (N_28295,N_27071,N_27122);
nor U28296 (N_28296,N_27479,N_26343);
nor U28297 (N_28297,N_26115,N_27527);
and U28298 (N_28298,N_26594,N_27339);
nor U28299 (N_28299,N_27999,N_27765);
and U28300 (N_28300,N_27935,N_27288);
or U28301 (N_28301,N_26992,N_27460);
or U28302 (N_28302,N_27483,N_27489);
or U28303 (N_28303,N_27594,N_27137);
and U28304 (N_28304,N_27340,N_26058);
or U28305 (N_28305,N_26403,N_26187);
or U28306 (N_28306,N_27636,N_26807);
or U28307 (N_28307,N_26810,N_26081);
and U28308 (N_28308,N_27550,N_26232);
or U28309 (N_28309,N_26729,N_27761);
and U28310 (N_28310,N_27650,N_27188);
or U28311 (N_28311,N_27826,N_26883);
and U28312 (N_28312,N_27433,N_27798);
xnor U28313 (N_28313,N_26042,N_27980);
nor U28314 (N_28314,N_27370,N_27878);
or U28315 (N_28315,N_26476,N_27778);
nor U28316 (N_28316,N_27484,N_26545);
xnor U28317 (N_28317,N_26846,N_27827);
xnor U28318 (N_28318,N_27038,N_27863);
or U28319 (N_28319,N_26852,N_26492);
xor U28320 (N_28320,N_27564,N_27696);
and U28321 (N_28321,N_27522,N_27260);
nor U28322 (N_28322,N_27314,N_27704);
nor U28323 (N_28323,N_27709,N_26149);
xor U28324 (N_28324,N_27572,N_26046);
xnor U28325 (N_28325,N_27112,N_26652);
nor U28326 (N_28326,N_26426,N_26164);
nand U28327 (N_28327,N_26832,N_27480);
and U28328 (N_28328,N_27049,N_27443);
and U28329 (N_28329,N_26595,N_27091);
nand U28330 (N_28330,N_27099,N_26720);
and U28331 (N_28331,N_27105,N_26156);
and U28332 (N_28332,N_26291,N_26331);
nor U28333 (N_28333,N_27058,N_26161);
or U28334 (N_28334,N_26214,N_26881);
nand U28335 (N_28335,N_27702,N_27622);
xnor U28336 (N_28336,N_27083,N_26876);
xor U28337 (N_28337,N_26959,N_27265);
xnor U28338 (N_28338,N_26337,N_26448);
or U28339 (N_28339,N_26796,N_27347);
or U28340 (N_28340,N_27595,N_27015);
and U28341 (N_28341,N_26651,N_26314);
and U28342 (N_28342,N_26797,N_27304);
or U28343 (N_28343,N_26256,N_26480);
nand U28344 (N_28344,N_27313,N_26975);
and U28345 (N_28345,N_26633,N_26433);
xnor U28346 (N_28346,N_27395,N_26127);
nor U28347 (N_28347,N_27132,N_26567);
or U28348 (N_28348,N_26895,N_27297);
and U28349 (N_28349,N_26312,N_26064);
nand U28350 (N_28350,N_26025,N_26663);
or U28351 (N_28351,N_27570,N_27833);
or U28352 (N_28352,N_27108,N_26551);
nand U28353 (N_28353,N_27226,N_26497);
and U28354 (N_28354,N_27459,N_26643);
nand U28355 (N_28355,N_26816,N_27268);
nand U28356 (N_28356,N_27045,N_27705);
and U28357 (N_28357,N_26593,N_26200);
and U28358 (N_28358,N_26916,N_27675);
or U28359 (N_28359,N_26732,N_27237);
xor U28360 (N_28360,N_26067,N_27152);
nand U28361 (N_28361,N_26029,N_26566);
or U28362 (N_28362,N_26028,N_26944);
nand U28363 (N_28363,N_26800,N_27295);
and U28364 (N_28364,N_26829,N_27914);
and U28365 (N_28365,N_27060,N_27874);
nor U28366 (N_28366,N_27471,N_27756);
or U28367 (N_28367,N_26580,N_26053);
and U28368 (N_28368,N_27955,N_26140);
nor U28369 (N_28369,N_26332,N_27953);
nand U28370 (N_28370,N_27871,N_26317);
nand U28371 (N_28371,N_27263,N_26056);
or U28372 (N_28372,N_26307,N_26967);
nor U28373 (N_28373,N_27266,N_26742);
nor U28374 (N_28374,N_26988,N_27837);
and U28375 (N_28375,N_26615,N_27845);
xor U28376 (N_28376,N_26573,N_26106);
and U28377 (N_28377,N_26259,N_27653);
or U28378 (N_28378,N_26366,N_27513);
and U28379 (N_28379,N_26686,N_26330);
or U28380 (N_28380,N_27162,N_26089);
and U28381 (N_28381,N_27873,N_27603);
or U28382 (N_28382,N_27092,N_27554);
xnor U28383 (N_28383,N_27512,N_26342);
nand U28384 (N_28384,N_26504,N_26094);
or U28385 (N_28385,N_26823,N_26052);
and U28386 (N_28386,N_27496,N_26392);
nand U28387 (N_28387,N_26907,N_26639);
nor U28388 (N_28388,N_26326,N_27500);
and U28389 (N_28389,N_26837,N_26641);
xnor U28390 (N_28390,N_26840,N_27423);
and U28391 (N_28391,N_26836,N_26890);
nor U28392 (N_28392,N_27928,N_27343);
nand U28393 (N_28393,N_27734,N_26999);
or U28394 (N_28394,N_26427,N_26887);
or U28395 (N_28395,N_26015,N_27875);
nand U28396 (N_28396,N_26647,N_26194);
and U28397 (N_28397,N_27829,N_26645);
xnor U28398 (N_28398,N_27070,N_26080);
and U28399 (N_28399,N_27123,N_27718);
xor U28400 (N_28400,N_26266,N_26113);
nand U28401 (N_28401,N_27114,N_26570);
nor U28402 (N_28402,N_27391,N_26953);
nor U28403 (N_28403,N_26706,N_27177);
xnor U28404 (N_28404,N_26533,N_27848);
and U28405 (N_28405,N_26117,N_27148);
xnor U28406 (N_28406,N_26236,N_27389);
or U28407 (N_28407,N_27504,N_26774);
nor U28408 (N_28408,N_27966,N_26815);
xor U28409 (N_28409,N_26696,N_26002);
nor U28410 (N_28410,N_26268,N_26146);
nor U28411 (N_28411,N_26541,N_26019);
nand U28412 (N_28412,N_26913,N_26888);
nor U28413 (N_28413,N_26475,N_26402);
or U28414 (N_28414,N_26786,N_26733);
nor U28415 (N_28415,N_27692,N_26011);
and U28416 (N_28416,N_27757,N_26205);
or U28417 (N_28417,N_26092,N_26454);
xor U28418 (N_28418,N_27254,N_26879);
xor U28419 (N_28419,N_27375,N_26109);
nand U28420 (N_28420,N_26423,N_27851);
or U28421 (N_28421,N_26073,N_27416);
xor U28422 (N_28422,N_27710,N_26932);
and U28423 (N_28423,N_26899,N_26483);
nor U28424 (N_28424,N_26175,N_27933);
and U28425 (N_28425,N_27213,N_27191);
nor U28426 (N_28426,N_26531,N_27822);
nand U28427 (N_28427,N_27717,N_26023);
nor U28428 (N_28428,N_27046,N_27025);
xor U28429 (N_28429,N_26987,N_27497);
or U28430 (N_28430,N_26470,N_26163);
or U28431 (N_28431,N_26994,N_27136);
nand U28432 (N_28432,N_26867,N_27625);
or U28433 (N_28433,N_27218,N_27608);
and U28434 (N_28434,N_26609,N_27576);
xor U28435 (N_28435,N_26351,N_27053);
nand U28436 (N_28436,N_27214,N_27583);
or U28437 (N_28437,N_26518,N_27390);
and U28438 (N_28438,N_27751,N_26218);
nor U28439 (N_28439,N_27900,N_27929);
nor U28440 (N_28440,N_26340,N_26989);
nand U28441 (N_28441,N_26369,N_26128);
nand U28442 (N_28442,N_27632,N_27217);
xnor U28443 (N_28443,N_27965,N_26602);
or U28444 (N_28444,N_26429,N_27711);
nand U28445 (N_28445,N_27185,N_26281);
and U28446 (N_28446,N_27016,N_27308);
nand U28447 (N_28447,N_27195,N_26242);
nand U28448 (N_28448,N_27118,N_26083);
xnor U28449 (N_28449,N_27721,N_27001);
nand U28450 (N_28450,N_26710,N_26640);
nand U28451 (N_28451,N_26866,N_27651);
or U28452 (N_28452,N_27350,N_27498);
and U28453 (N_28453,N_26293,N_26278);
or U28454 (N_28454,N_26788,N_26982);
or U28455 (N_28455,N_27736,N_26770);
xor U28456 (N_28456,N_27915,N_26502);
nor U28457 (N_28457,N_26997,N_26554);
or U28458 (N_28458,N_27328,N_27707);
xnor U28459 (N_28459,N_27532,N_26139);
nand U28460 (N_28460,N_27860,N_27972);
or U28461 (N_28461,N_27455,N_26172);
and U28462 (N_28462,N_27022,N_26421);
and U28463 (N_28463,N_26420,N_26897);
nor U28464 (N_28464,N_27321,N_27701);
nor U28465 (N_28465,N_27342,N_26493);
and U28466 (N_28466,N_26016,N_27207);
and U28467 (N_28467,N_27887,N_26377);
nand U28468 (N_28468,N_27879,N_26949);
nand U28469 (N_28469,N_26917,N_26443);
and U28470 (N_28470,N_26787,N_26782);
xor U28471 (N_28471,N_26703,N_27209);
xnor U28472 (N_28472,N_26086,N_27731);
or U28473 (N_28473,N_27932,N_26669);
xor U28474 (N_28474,N_26150,N_27020);
xor U28475 (N_28475,N_26735,N_26957);
nor U28476 (N_28476,N_27469,N_26882);
and U28477 (N_28477,N_27507,N_26751);
or U28478 (N_28478,N_26857,N_27138);
or U28479 (N_28479,N_26875,N_26035);
or U28480 (N_28480,N_27486,N_27506);
nand U28481 (N_28481,N_27646,N_27797);
xnor U28482 (N_28482,N_27883,N_26051);
and U28483 (N_28483,N_27333,N_26077);
xnor U28484 (N_28484,N_26207,N_27441);
or U28485 (N_28485,N_26068,N_27006);
nand U28486 (N_28486,N_27482,N_27852);
or U28487 (N_28487,N_26240,N_27945);
nor U28488 (N_28488,N_27145,N_27495);
nand U28489 (N_28489,N_26900,N_27926);
and U28490 (N_28490,N_27591,N_27100);
xor U28491 (N_28491,N_26948,N_27247);
or U28492 (N_28492,N_26801,N_27830);
and U28493 (N_28493,N_27403,N_26880);
xnor U28494 (N_28494,N_27278,N_26745);
nor U28495 (N_28495,N_26956,N_27303);
and U28496 (N_28496,N_26672,N_26280);
nor U28497 (N_28497,N_26301,N_27167);
and U28498 (N_28498,N_27976,N_26532);
and U28499 (N_28499,N_27291,N_26477);
nor U28500 (N_28500,N_27468,N_26743);
xor U28501 (N_28501,N_26171,N_27202);
and U28502 (N_28502,N_27434,N_26100);
and U28503 (N_28503,N_26233,N_27553);
nor U28504 (N_28504,N_27567,N_26730);
or U28505 (N_28505,N_26484,N_26705);
xnor U28506 (N_28506,N_26495,N_27224);
and U28507 (N_28507,N_26847,N_27739);
and U28508 (N_28508,N_27243,N_27519);
and U28509 (N_28509,N_26749,N_27673);
nand U28510 (N_28510,N_27430,N_26154);
nor U28511 (N_28511,N_26061,N_27079);
xnor U28512 (N_28512,N_27919,N_27345);
xor U28513 (N_28513,N_27381,N_26738);
nand U28514 (N_28514,N_26131,N_27206);
nor U28515 (N_28515,N_27963,N_27086);
or U28516 (N_28516,N_27898,N_26287);
and U28517 (N_28517,N_26491,N_26292);
nor U28518 (N_28518,N_27938,N_27410);
and U28519 (N_28519,N_26500,N_27931);
nor U28520 (N_28520,N_27098,N_27141);
and U28521 (N_28521,N_26625,N_27437);
nor U28522 (N_28522,N_26265,N_26858);
or U28523 (N_28523,N_27330,N_26958);
nor U28524 (N_28524,N_26855,N_26066);
nor U28525 (N_28525,N_27449,N_26698);
or U28526 (N_28526,N_27961,N_27173);
or U28527 (N_28527,N_27317,N_26552);
or U28528 (N_28528,N_27287,N_26009);
nor U28529 (N_28529,N_27666,N_27748);
nand U28530 (N_28530,N_26623,N_26219);
and U28531 (N_28531,N_27714,N_26119);
and U28532 (N_28532,N_27760,N_26044);
or U28533 (N_28533,N_26924,N_27155);
and U28534 (N_28534,N_26255,N_26082);
and U28535 (N_28535,N_26973,N_26101);
xor U28536 (N_28536,N_26167,N_27859);
nand U28537 (N_28537,N_27885,N_27250);
or U28538 (N_28538,N_27284,N_26258);
nor U28539 (N_28539,N_26310,N_27074);
nand U28540 (N_28540,N_27604,N_27249);
and U28541 (N_28541,N_27135,N_26374);
xnor U28542 (N_28542,N_27259,N_27069);
or U28543 (N_28543,N_26747,N_26469);
xnor U28544 (N_28544,N_26350,N_26808);
and U28545 (N_28545,N_26599,N_26054);
nand U28546 (N_28546,N_27401,N_26834);
nor U28547 (N_28547,N_26412,N_26779);
and U28548 (N_28548,N_26868,N_26399);
nand U28549 (N_28549,N_26279,N_27172);
or U28550 (N_28550,N_27986,N_27864);
or U28551 (N_28551,N_27643,N_27911);
nor U28552 (N_28552,N_27943,N_27834);
or U28553 (N_28553,N_26783,N_27788);
nand U28554 (N_28554,N_27655,N_26409);
and U28555 (N_28555,N_26535,N_27289);
nor U28556 (N_28556,N_27688,N_26251);
xnor U28557 (N_28557,N_27800,N_27508);
or U28558 (N_28558,N_26694,N_27012);
and U28559 (N_28559,N_26414,N_27738);
xnor U28560 (N_28560,N_26257,N_27726);
or U28561 (N_28561,N_26547,N_27638);
nand U28562 (N_28562,N_27208,N_27067);
xor U28563 (N_28563,N_26931,N_26418);
xnor U28564 (N_28564,N_27993,N_27805);
nor U28565 (N_28565,N_26440,N_27037);
xor U28566 (N_28566,N_26526,N_27360);
or U28567 (N_28567,N_27607,N_27230);
nand U28568 (N_28568,N_27846,N_26726);
or U28569 (N_28569,N_27590,N_27280);
or U28570 (N_28570,N_27432,N_26539);
and U28571 (N_28571,N_26288,N_26589);
nor U28572 (N_28572,N_27244,N_26252);
xor U28573 (N_28573,N_27950,N_26693);
and U28574 (N_28574,N_26070,N_27525);
nor U28575 (N_28575,N_26830,N_27905);
nor U28576 (N_28576,N_26940,N_26381);
nor U28577 (N_28577,N_27298,N_27732);
nor U28578 (N_28578,N_26825,N_26438);
xnor U28579 (N_28579,N_27181,N_27361);
or U28580 (N_28580,N_27545,N_26202);
xor U28581 (N_28581,N_27398,N_27893);
nor U28582 (N_28582,N_27967,N_26752);
xor U28583 (N_28583,N_27338,N_26528);
nor U28584 (N_28584,N_26031,N_27648);
nand U28585 (N_28585,N_26764,N_26995);
xor U28586 (N_28586,N_26685,N_27916);
nor U28587 (N_28587,N_26616,N_27796);
and U28588 (N_28588,N_26111,N_27907);
and U28589 (N_28589,N_27346,N_27359);
xnor U28590 (N_28590,N_27066,N_26473);
xnor U28591 (N_28591,N_27753,N_27740);
or U28592 (N_28592,N_26296,N_26397);
or U28593 (N_28593,N_26673,N_27971);
or U28594 (N_28594,N_27810,N_26984);
xor U28595 (N_28595,N_27906,N_27799);
nand U28596 (N_28596,N_27954,N_26719);
xnor U28597 (N_28597,N_26543,N_26632);
nand U28598 (N_28598,N_26793,N_27085);
and U28599 (N_28599,N_26190,N_27062);
nor U28600 (N_28600,N_26664,N_27992);
xor U28601 (N_28601,N_26116,N_26262);
xnor U28602 (N_28602,N_26920,N_27735);
or U28603 (N_28603,N_27201,N_26884);
nor U28604 (N_28604,N_26168,N_26309);
nand U28605 (N_28605,N_27131,N_27605);
and U28606 (N_28606,N_27282,N_26189);
xnor U28607 (N_28607,N_26169,N_26393);
nor U28608 (N_28608,N_26275,N_26679);
nand U28609 (N_28609,N_26313,N_26778);
or U28610 (N_28610,N_26012,N_26124);
xor U28611 (N_28611,N_27270,N_26300);
nand U28612 (N_28612,N_27615,N_27679);
or U28613 (N_28613,N_26512,N_26220);
and U28614 (N_28614,N_27503,N_27248);
and U28615 (N_28615,N_26471,N_27517);
and U28616 (N_28616,N_26445,N_26699);
nand U28617 (N_28617,N_26926,N_27974);
and U28618 (N_28618,N_26277,N_27402);
xor U28619 (N_28619,N_26728,N_26675);
nand U28620 (N_28620,N_26180,N_26322);
xor U28621 (N_28621,N_26842,N_26697);
and U28622 (N_28622,N_27385,N_26871);
and U28623 (N_28623,N_27599,N_26489);
or U28624 (N_28624,N_27392,N_27277);
or U28625 (N_28625,N_26193,N_26785);
nand U28626 (N_28626,N_27200,N_27678);
and U28627 (N_28627,N_27474,N_26095);
and U28628 (N_28628,N_26178,N_26022);
nor U28629 (N_28629,N_27597,N_26213);
nor U28630 (N_28630,N_27635,N_26701);
and U28631 (N_28631,N_27858,N_26577);
nand U28632 (N_28632,N_27752,N_26723);
nor U28633 (N_28633,N_26142,N_26687);
and U28634 (N_28634,N_27663,N_26819);
nand U28635 (N_28635,N_26424,N_27267);
nor U28636 (N_28636,N_26822,N_27087);
nand U28637 (N_28637,N_27803,N_27593);
xnor U28638 (N_28638,N_26621,N_26055);
xnor U28639 (N_28639,N_27013,N_26224);
xnor U28640 (N_28640,N_26486,N_26334);
nor U28641 (N_28641,N_26596,N_27413);
nor U28642 (N_28642,N_26809,N_26634);
nor U28643 (N_28643,N_26737,N_27523);
and U28644 (N_28644,N_27559,N_26561);
or U28645 (N_28645,N_27686,N_27526);
nor U28646 (N_28646,N_26160,N_27669);
and U28647 (N_28647,N_27334,N_26467);
or U28648 (N_28648,N_27939,N_26758);
xnor U28649 (N_28649,N_27043,N_27073);
nand U28650 (N_28650,N_27026,N_26838);
nor U28651 (N_28651,N_26225,N_26937);
xor U28652 (N_28652,N_26534,N_26108);
or U28653 (N_28653,N_26441,N_26162);
xor U28654 (N_28654,N_27261,N_26813);
nand U28655 (N_28655,N_26153,N_27539);
and U28656 (N_28656,N_26406,N_26557);
xnor U28657 (N_28657,N_26375,N_27336);
nand U28658 (N_28658,N_26766,N_27411);
nand U28659 (N_28659,N_27642,N_26629);
or U28660 (N_28660,N_27804,N_26996);
or U28661 (N_28661,N_26773,N_27011);
and U28662 (N_28662,N_26911,N_26761);
and U28663 (N_28663,N_27127,N_27989);
nor U28664 (N_28664,N_26667,N_26853);
or U28665 (N_28665,N_26775,N_26511);
xor U28666 (N_28666,N_26198,N_26344);
and U28667 (N_28667,N_26181,N_26684);
or U28668 (N_28668,N_27689,N_26359);
xor U28669 (N_28669,N_27095,N_27404);
and U28670 (N_28670,N_27150,N_26099);
xnor U28671 (N_28671,N_27681,N_27913);
nand U28672 (N_28672,N_27930,N_27417);
nor U28673 (N_28673,N_27241,N_26203);
nand U28674 (N_28674,N_27072,N_26386);
nor U28675 (N_28675,N_26839,N_27445);
xnor U28676 (N_28676,N_27179,N_27842);
or U28677 (N_28677,N_26151,N_27235);
and U28678 (N_28678,N_26578,N_27944);
and U28679 (N_28679,N_26027,N_26638);
nor U28680 (N_28680,N_27494,N_27415);
or U28681 (N_28681,N_26447,N_26458);
xor U28682 (N_28682,N_27130,N_26833);
xnor U28683 (N_28683,N_26226,N_26184);
and U28684 (N_28684,N_26404,N_26915);
nor U28685 (N_28685,N_27451,N_26791);
nand U28686 (N_28686,N_26230,N_26522);
and U28687 (N_28687,N_26943,N_27589);
xor U28688 (N_28688,N_26479,N_27660);
nand U28689 (N_28689,N_27242,N_26260);
nand U28690 (N_28690,N_27876,N_26261);
nor U28691 (N_28691,N_27109,N_26649);
nand U28692 (N_28692,N_27720,N_27917);
xnor U28693 (N_28693,N_26939,N_26302);
and U28694 (N_28694,N_26925,N_26928);
and U28695 (N_28695,N_27668,N_27357);
nand U28696 (N_28696,N_27082,N_27151);
and U28697 (N_28697,N_27832,N_26311);
xnor U28698 (N_28698,N_27374,N_27582);
and U28699 (N_28699,N_27307,N_26461);
nor U28700 (N_28700,N_27521,N_26103);
xnor U28701 (N_28701,N_26608,N_27337);
xor U28702 (N_28702,N_26927,N_27234);
nand U28703 (N_28703,N_27922,N_26711);
and U28704 (N_28704,N_27547,N_27687);
nor U28705 (N_28705,N_26267,N_27924);
or U28706 (N_28706,N_26072,N_27031);
and U28707 (N_28707,N_26814,N_27892);
nand U28708 (N_28708,N_26765,N_26734);
and U28709 (N_28709,N_27096,N_27794);
xor U28710 (N_28710,N_26585,N_27776);
and U28711 (N_28711,N_27055,N_27212);
or U28712 (N_28712,N_26201,N_26562);
nand U28713 (N_28713,N_26831,N_26238);
and U28714 (N_28714,N_27634,N_27712);
nand U28715 (N_28715,N_27444,N_26282);
xor U28716 (N_28716,N_27412,N_26771);
xnor U28717 (N_28717,N_27204,N_26361);
xor U28718 (N_28718,N_26516,N_27332);
or U28719 (N_28719,N_27579,N_27094);
or U28720 (N_28720,N_27693,N_26248);
and U28721 (N_28721,N_27018,N_27393);
or U28722 (N_28722,N_27305,N_26731);
and U28723 (N_28723,N_26950,N_27620);
nand U28724 (N_28724,N_27866,N_27467);
or U28725 (N_28725,N_27032,N_27771);
nor U28726 (N_28726,N_26269,N_26196);
nand U28727 (N_28727,N_26503,N_27565);
xnor U28728 (N_28728,N_27637,N_27667);
or U28729 (N_28729,N_26676,N_26759);
xor U28730 (N_28730,N_26670,N_26592);
or U28731 (N_28731,N_26523,N_26208);
xnor U28732 (N_28732,N_26297,N_27367);
or U28733 (N_28733,N_26034,N_27502);
nor U28734 (N_28734,N_26827,N_27057);
and U28735 (N_28735,N_26338,N_26229);
nand U28736 (N_28736,N_26923,N_26107);
nand U28737 (N_28737,N_27578,N_27458);
xor U28738 (N_28738,N_26525,N_27808);
nor U28739 (N_28739,N_27767,N_27324);
or U28740 (N_28740,N_27035,N_26678);
and U28741 (N_28741,N_27868,N_27923);
nand U28742 (N_28742,N_27715,N_27192);
or U28743 (N_28743,N_26304,N_27774);
or U28744 (N_28744,N_26571,N_27190);
xor U28745 (N_28745,N_26904,N_27447);
and U28746 (N_28746,N_27654,N_27544);
xor U28747 (N_28747,N_27171,N_26356);
and U28748 (N_28748,N_26540,N_26581);
or U28749 (N_28749,N_27027,N_26794);
or U28750 (N_28750,N_27220,N_26965);
and U28751 (N_28751,N_26872,N_26315);
nand U28752 (N_28752,N_26177,N_27143);
xnor U28753 (N_28753,N_26688,N_26363);
or U28754 (N_28754,N_27050,N_27183);
nand U28755 (N_28755,N_26299,N_26555);
or U28756 (N_28756,N_27677,N_26795);
or U28757 (N_28757,N_26416,N_27407);
xor U28758 (N_28758,N_27144,N_27124);
or U28759 (N_28759,N_27957,N_27276);
and U28760 (N_28760,N_27725,N_27819);
nor U28761 (N_28761,N_27408,N_26253);
and U28762 (N_28762,N_27656,N_27450);
xnor U28763 (N_28763,N_27728,N_26138);
nor U28764 (N_28764,N_26104,N_26692);
nor U28765 (N_28765,N_26969,N_26753);
nor U28766 (N_28766,N_27694,N_26076);
nor U28767 (N_28767,N_27197,N_26978);
and U28768 (N_28768,N_27194,N_26017);
and U28769 (N_28769,N_26173,N_26565);
or U28770 (N_28770,N_27708,N_27329);
or U28771 (N_28771,N_27456,N_26327);
nand U28772 (N_28772,N_26563,N_27139);
xor U28773 (N_28773,N_27326,N_27296);
nor U28774 (N_28774,N_26065,N_27614);
xor U28775 (N_28775,N_27626,N_26657);
and U28776 (N_28776,N_26134,N_27783);
nand U28777 (N_28777,N_26195,N_26909);
and U28778 (N_28778,N_26417,N_26650);
and U28779 (N_28779,N_26389,N_27973);
or U28780 (N_28780,N_27792,N_26961);
or U28781 (N_28781,N_26382,N_26152);
xor U28782 (N_28782,N_27975,N_27182);
nand U28783 (N_28783,N_26004,N_27563);
xor U28784 (N_28784,N_27464,N_26844);
nor U28785 (N_28785,N_27733,N_27515);
and U28786 (N_28786,N_26199,N_27210);
xnor U28787 (N_28787,N_27960,N_26553);
xnor U28788 (N_28788,N_27514,N_27747);
or U28789 (N_28789,N_26114,N_26941);
or U28790 (N_28790,N_26341,N_27759);
or U28791 (N_28791,N_27925,N_26681);
nand U28792 (N_28792,N_26045,N_27425);
and U28793 (N_28793,N_27713,N_27891);
and U28794 (N_28794,N_27163,N_26136);
nor U28795 (N_28795,N_27488,N_26718);
and U28796 (N_28796,N_27352,N_27890);
nand U28797 (N_28797,N_26826,N_26569);
nand U28798 (N_28798,N_26611,N_27223);
nor U28799 (N_28799,N_27088,N_27746);
and U28800 (N_28800,N_26298,N_26328);
and U28801 (N_28801,N_27363,N_27685);
xnor U28802 (N_28802,N_27533,N_26294);
nor U28803 (N_28803,N_26517,N_26506);
xnor U28804 (N_28804,N_26754,N_27538);
and U28805 (N_28805,N_27501,N_27768);
nand U28806 (N_28806,N_27034,N_26485);
and U28807 (N_28807,N_26707,N_26249);
nor U28808 (N_28808,N_26537,N_26901);
nand U28809 (N_28809,N_27189,N_27958);
nor U28810 (N_28810,N_27568,N_26893);
nor U28811 (N_28811,N_27184,N_26977);
and U28812 (N_28812,N_26006,N_26244);
nand U28813 (N_28813,N_26886,N_26780);
nor U28814 (N_28814,N_27023,N_26619);
or U28815 (N_28815,N_26990,N_27624);
nand U28816 (N_28816,N_27492,N_26049);
nor U28817 (N_28817,N_27119,N_26093);
nand U28818 (N_28818,N_27536,N_26494);
and U28819 (N_28819,N_26991,N_26520);
and U28820 (N_28820,N_27081,N_26574);
xnor U28821 (N_28821,N_27601,N_27949);
nand U28822 (N_28822,N_26254,N_27901);
or U28823 (N_28823,N_27054,N_26617);
nand U28824 (N_28824,N_27947,N_27021);
xor U28825 (N_28825,N_27301,N_26020);
nor U28826 (N_28826,N_26088,N_26631);
nor U28827 (N_28827,N_26691,N_26234);
or U28828 (N_28828,N_26318,N_26985);
nand U28829 (N_28829,N_27318,N_26333);
and U28830 (N_28830,N_26824,N_27785);
xor U28831 (N_28831,N_27592,N_27865);
nor U28832 (N_28832,N_27327,N_27061);
nor U28833 (N_28833,N_27529,N_26057);
nand U28834 (N_28834,N_27380,N_26601);
or U28835 (N_28835,N_27258,N_26712);
xnor U28836 (N_28836,N_27236,N_27828);
or U28837 (N_28837,N_27520,N_27142);
nor U28838 (N_28838,N_26498,N_27611);
nor U28839 (N_28839,N_27621,N_27029);
xnor U28840 (N_28840,N_27157,N_27509);
xor U28841 (N_28841,N_26848,N_26658);
and U28842 (N_28842,N_27574,N_26062);
or U28843 (N_28843,N_26264,N_27524);
and U28844 (N_28844,N_27936,N_26105);
or U28845 (N_28845,N_27470,N_26896);
and U28846 (N_28846,N_27744,N_26695);
or U28847 (N_28847,N_26653,N_26384);
nand U28848 (N_28848,N_27418,N_27823);
and U28849 (N_28849,N_26284,N_26446);
xnor U28850 (N_28850,N_26488,N_27937);
xor U28851 (N_28851,N_26674,N_27816);
nor U28852 (N_28852,N_26010,N_26041);
xor U28853 (N_28853,N_26964,N_26290);
or U28854 (N_28854,N_27125,N_26644);
nor U28855 (N_28855,N_26126,N_26324);
xnor U28856 (N_28856,N_27366,N_26604);
and U28857 (N_28857,N_27531,N_27149);
nand U28858 (N_28858,N_27990,N_26514);
or U28859 (N_28859,N_27399,N_27956);
nor U28860 (N_28860,N_27652,N_27103);
or U28861 (N_28861,N_26323,N_27807);
nand U28862 (N_28862,N_27750,N_26860);
nand U28863 (N_28863,N_27068,N_27657);
nor U28864 (N_28864,N_26074,N_27779);
nor U28865 (N_28865,N_26148,N_27941);
nand U28866 (N_28866,N_26133,N_27787);
nand U28867 (N_28867,N_27558,N_27537);
and U28868 (N_28868,N_27047,N_27325);
nand U28869 (N_28869,N_27044,N_26660);
xnor U28870 (N_28870,N_26144,N_26013);
or U28871 (N_28871,N_27063,N_26998);
and U28872 (N_28872,N_27102,N_26903);
nand U28873 (N_28873,N_26018,N_26870);
xor U28874 (N_28874,N_27535,N_27439);
and U28875 (N_28875,N_26464,N_26529);
nand U28876 (N_28876,N_26963,N_26721);
and U28877 (N_28877,N_27940,N_26648);
or U28878 (N_28878,N_27281,N_26781);
and U28879 (N_28879,N_27782,N_27344);
or U28880 (N_28880,N_27180,N_26856);
nand U28881 (N_28881,N_26452,N_26319);
nor U28882 (N_28882,N_26174,N_26906);
nand U28883 (N_28883,N_27229,N_27397);
or U28884 (N_28884,N_27275,N_26400);
or U28885 (N_28885,N_27426,N_26789);
and U28886 (N_28886,N_27959,N_26245);
nand U28887 (N_28887,N_26487,N_26176);
nand U28888 (N_28888,N_26183,N_27440);
or U28889 (N_28889,N_26000,N_27104);
xnor U28890 (N_28890,N_27719,N_26792);
nand U28891 (N_28891,N_27419,N_27889);
nor U28892 (N_28892,N_27853,N_26803);
and U28893 (N_28893,N_26357,N_27727);
nand U28894 (N_28894,N_26744,N_27406);
or U28895 (N_28895,N_27770,N_26345);
or U28896 (N_28896,N_26250,N_27815);
nand U28897 (N_28897,N_27910,N_26769);
nor U28898 (N_28898,N_27227,N_26508);
or U28899 (N_28899,N_27908,N_27560);
nand U28900 (N_28900,N_26877,N_27090);
nor U28901 (N_28901,N_26677,N_27255);
and U28902 (N_28902,N_26084,N_26757);
nand U28903 (N_28903,N_27690,N_26368);
xor U28904 (N_28904,N_26428,N_26811);
and U28905 (N_28905,N_27097,N_26159);
nor U28906 (N_28906,N_27633,N_27351);
xor U28907 (N_28907,N_26918,N_27641);
xor U28908 (N_28908,N_27662,N_27176);
and U28909 (N_28909,N_26263,N_27847);
and U28910 (N_28910,N_26835,N_27041);
xor U28911 (N_28911,N_26398,N_27676);
xnor U28912 (N_28912,N_26321,N_26431);
nor U28913 (N_28913,N_27505,N_27147);
or U28914 (N_28914,N_27231,N_27510);
xnor U28915 (N_28915,N_26241,N_26527);
nand U28916 (N_28916,N_27170,N_27682);
nand U28917 (N_28917,N_26544,N_26422);
nand U28918 (N_28918,N_26654,N_27222);
nor U28919 (N_28919,N_26370,N_26894);
nand U28920 (N_28920,N_27414,N_26362);
nand U28921 (N_28921,N_26482,N_26436);
or U28922 (N_28922,N_27299,N_26383);
xor U28923 (N_28923,N_26223,N_26165);
or U28924 (N_28924,N_26371,N_26003);
nor U28925 (N_28925,N_26790,N_26182);
xnor U28926 (N_28926,N_26439,N_26360);
and U28927 (N_28927,N_27372,N_27476);
or U28928 (N_28928,N_26098,N_26841);
and U28929 (N_28929,N_27540,N_26474);
nor U28930 (N_28930,N_26388,N_26014);
nor U28931 (N_28931,N_27493,N_27987);
xor U28932 (N_28932,N_26680,N_26087);
and U28933 (N_28933,N_27084,N_27319);
or U28934 (N_28934,N_27429,N_26635);
xnor U28935 (N_28935,N_26750,N_27584);
nand U28936 (N_28936,N_26564,N_26246);
xnor U28937 (N_28937,N_27310,N_26033);
nor U28938 (N_28938,N_27473,N_26885);
or U28939 (N_28939,N_26063,N_27843);
or U28940 (N_28940,N_26444,N_27839);
or U28941 (N_28941,N_27110,N_27665);
xnor U28942 (N_28942,N_27153,N_26271);
and U28943 (N_28943,N_27649,N_27341);
and U28944 (N_28944,N_26777,N_26510);
xnor U28945 (N_28945,N_27983,N_27880);
xor U28946 (N_28946,N_27854,N_26145);
nand U28947 (N_28947,N_26845,N_26579);
nand U28948 (N_28948,N_26760,N_26550);
or U28949 (N_28949,N_26614,N_27549);
xnor U28950 (N_28950,N_26716,N_26459);
or U28951 (N_28951,N_27629,N_26768);
and U28952 (N_28952,N_27749,N_26938);
xnor U28953 (N_28953,N_27754,N_26946);
or U28954 (N_28954,N_26185,N_27472);
or U28955 (N_28955,N_26530,N_27902);
nand U28956 (N_28956,N_26451,N_26933);
nor U28957 (N_28957,N_27904,N_27763);
and U28958 (N_28958,N_26303,N_27817);
nand U28959 (N_28959,N_27048,N_26499);
nand U28960 (N_28960,N_27159,N_27658);
or U28961 (N_28961,N_26155,N_27442);
nor U28962 (N_28962,N_27647,N_27272);
nor U28963 (N_28963,N_26391,N_27575);
nor U28964 (N_28964,N_26889,N_27435);
and U28965 (N_28965,N_27420,N_26934);
nor U28966 (N_28966,N_26170,N_27382);
and U28967 (N_28967,N_26849,N_26395);
nor U28968 (N_28968,N_27841,N_27730);
and U28969 (N_28969,N_27285,N_27806);
xor U28970 (N_28970,N_26372,N_26921);
nand U28971 (N_28971,N_26929,N_26407);
nor U28972 (N_28972,N_26507,N_26746);
or U28973 (N_28973,N_27617,N_26179);
nor U28974 (N_28974,N_27587,N_27089);
or U28975 (N_28975,N_26859,N_27203);
nand U28976 (N_28976,N_27245,N_26700);
xnor U28977 (N_28977,N_27457,N_27618);
or U28978 (N_28978,N_27946,N_27548);
or U28979 (N_28979,N_27888,N_27664);
or U28980 (N_28980,N_26763,N_27076);
and U28981 (N_28981,N_27680,N_27477);
xor U28982 (N_28982,N_26828,N_26460);
nor U28983 (N_28983,N_26217,N_26521);
nor U28984 (N_28984,N_27683,N_27238);
nor U28985 (N_28985,N_26047,N_27997);
nand U28986 (N_28986,N_27814,N_26624);
nand U28987 (N_28987,N_26283,N_27481);
nand U28988 (N_28988,N_26295,N_26799);
nor U28989 (N_28989,N_27706,N_27609);
or U28990 (N_28990,N_27857,N_27273);
or U28991 (N_28991,N_27017,N_26457);
xor U28992 (N_28992,N_27659,N_26434);
nand U28993 (N_28993,N_27995,N_26120);
and U28994 (N_28994,N_27671,N_26130);
xnor U28995 (N_28995,N_27781,N_26121);
nor U28996 (N_28996,N_27115,N_26556);
nand U28997 (N_28997,N_27463,N_26468);
nand U28998 (N_28998,N_26586,N_26935);
xnor U28999 (N_28999,N_27985,N_26419);
xor U29000 (N_29000,N_26500,N_26690);
nor U29001 (N_29001,N_26534,N_27676);
nor U29002 (N_29002,N_26424,N_27724);
and U29003 (N_29003,N_27044,N_27450);
or U29004 (N_29004,N_26886,N_27131);
or U29005 (N_29005,N_26143,N_27956);
and U29006 (N_29006,N_26724,N_27038);
and U29007 (N_29007,N_27366,N_27606);
nor U29008 (N_29008,N_27082,N_27421);
xor U29009 (N_29009,N_26550,N_27963);
nand U29010 (N_29010,N_27452,N_27035);
nor U29011 (N_29011,N_26361,N_26263);
and U29012 (N_29012,N_27231,N_26338);
and U29013 (N_29013,N_27520,N_27059);
and U29014 (N_29014,N_26403,N_26526);
xnor U29015 (N_29015,N_26128,N_27676);
nor U29016 (N_29016,N_26930,N_27819);
and U29017 (N_29017,N_27343,N_27256);
and U29018 (N_29018,N_27441,N_26913);
nor U29019 (N_29019,N_26432,N_26258);
or U29020 (N_29020,N_27476,N_27565);
nand U29021 (N_29021,N_26921,N_26072);
xnor U29022 (N_29022,N_26874,N_26332);
xor U29023 (N_29023,N_27334,N_26407);
xor U29024 (N_29024,N_27919,N_26239);
xnor U29025 (N_29025,N_26458,N_27583);
nor U29026 (N_29026,N_26062,N_27141);
nand U29027 (N_29027,N_27074,N_26262);
and U29028 (N_29028,N_27117,N_26958);
nand U29029 (N_29029,N_27698,N_27330);
and U29030 (N_29030,N_26893,N_27557);
or U29031 (N_29031,N_26281,N_27894);
or U29032 (N_29032,N_27057,N_27478);
and U29033 (N_29033,N_27881,N_27766);
nor U29034 (N_29034,N_27020,N_27533);
and U29035 (N_29035,N_26953,N_26115);
and U29036 (N_29036,N_26680,N_27692);
nor U29037 (N_29037,N_27346,N_27181);
or U29038 (N_29038,N_27924,N_27426);
or U29039 (N_29039,N_26416,N_26627);
or U29040 (N_29040,N_26969,N_26414);
and U29041 (N_29041,N_27452,N_26477);
and U29042 (N_29042,N_27573,N_27467);
or U29043 (N_29043,N_26623,N_26506);
and U29044 (N_29044,N_26194,N_26318);
and U29045 (N_29045,N_27120,N_26818);
xnor U29046 (N_29046,N_27060,N_26146);
nand U29047 (N_29047,N_26672,N_26971);
nor U29048 (N_29048,N_26554,N_27460);
nor U29049 (N_29049,N_27597,N_26036);
nor U29050 (N_29050,N_27480,N_26109);
nand U29051 (N_29051,N_27931,N_27846);
and U29052 (N_29052,N_26398,N_26587);
nor U29053 (N_29053,N_26903,N_26541);
and U29054 (N_29054,N_26530,N_26630);
xnor U29055 (N_29055,N_26682,N_26646);
nand U29056 (N_29056,N_26226,N_27932);
nand U29057 (N_29057,N_27469,N_27836);
xnor U29058 (N_29058,N_26370,N_26576);
or U29059 (N_29059,N_27258,N_27728);
xor U29060 (N_29060,N_26090,N_27211);
xor U29061 (N_29061,N_26549,N_27031);
or U29062 (N_29062,N_26945,N_26443);
and U29063 (N_29063,N_27948,N_27193);
xor U29064 (N_29064,N_26524,N_27760);
or U29065 (N_29065,N_27397,N_27599);
nor U29066 (N_29066,N_27672,N_26525);
nand U29067 (N_29067,N_27270,N_27213);
xor U29068 (N_29068,N_27354,N_26843);
nor U29069 (N_29069,N_26970,N_27105);
nand U29070 (N_29070,N_27195,N_26552);
nor U29071 (N_29071,N_26554,N_27426);
nor U29072 (N_29072,N_26400,N_26043);
or U29073 (N_29073,N_27290,N_27520);
and U29074 (N_29074,N_26349,N_26338);
nor U29075 (N_29075,N_26459,N_26421);
or U29076 (N_29076,N_27159,N_27918);
or U29077 (N_29077,N_27440,N_27954);
or U29078 (N_29078,N_26614,N_27255);
nand U29079 (N_29079,N_26652,N_26956);
xnor U29080 (N_29080,N_26351,N_26011);
and U29081 (N_29081,N_27995,N_27626);
nor U29082 (N_29082,N_27117,N_27167);
nand U29083 (N_29083,N_26934,N_27731);
or U29084 (N_29084,N_27381,N_26401);
xor U29085 (N_29085,N_26257,N_26012);
or U29086 (N_29086,N_26830,N_26516);
or U29087 (N_29087,N_27608,N_27638);
and U29088 (N_29088,N_27719,N_26618);
nand U29089 (N_29089,N_26697,N_26044);
or U29090 (N_29090,N_27462,N_26171);
nand U29091 (N_29091,N_26677,N_26146);
and U29092 (N_29092,N_26805,N_27672);
xnor U29093 (N_29093,N_26657,N_27541);
nand U29094 (N_29094,N_27192,N_26428);
xor U29095 (N_29095,N_26464,N_26552);
and U29096 (N_29096,N_27535,N_26770);
nand U29097 (N_29097,N_26131,N_26170);
or U29098 (N_29098,N_26156,N_27869);
nor U29099 (N_29099,N_27712,N_26428);
and U29100 (N_29100,N_27191,N_26392);
or U29101 (N_29101,N_26368,N_27321);
nor U29102 (N_29102,N_26141,N_26535);
or U29103 (N_29103,N_27719,N_26797);
nand U29104 (N_29104,N_27659,N_27925);
xor U29105 (N_29105,N_26526,N_27668);
and U29106 (N_29106,N_26045,N_26519);
nor U29107 (N_29107,N_27575,N_26092);
xnor U29108 (N_29108,N_26710,N_27416);
xor U29109 (N_29109,N_27272,N_26604);
or U29110 (N_29110,N_26186,N_27934);
nand U29111 (N_29111,N_26468,N_26196);
xor U29112 (N_29112,N_26466,N_26214);
and U29113 (N_29113,N_27558,N_26260);
or U29114 (N_29114,N_27612,N_27270);
or U29115 (N_29115,N_27579,N_26007);
nor U29116 (N_29116,N_26140,N_27667);
and U29117 (N_29117,N_27237,N_26934);
and U29118 (N_29118,N_26945,N_27748);
and U29119 (N_29119,N_26084,N_27070);
nor U29120 (N_29120,N_26712,N_27031);
xnor U29121 (N_29121,N_27338,N_26498);
xnor U29122 (N_29122,N_27686,N_26177);
nor U29123 (N_29123,N_27981,N_27552);
xor U29124 (N_29124,N_27192,N_26311);
nor U29125 (N_29125,N_26038,N_26267);
and U29126 (N_29126,N_26841,N_26135);
or U29127 (N_29127,N_27242,N_26770);
and U29128 (N_29128,N_26094,N_26676);
nor U29129 (N_29129,N_26447,N_27235);
nor U29130 (N_29130,N_27016,N_27320);
nand U29131 (N_29131,N_26700,N_27920);
or U29132 (N_29132,N_27601,N_26386);
nor U29133 (N_29133,N_26651,N_27795);
or U29134 (N_29134,N_27611,N_26109);
nand U29135 (N_29135,N_26817,N_26325);
and U29136 (N_29136,N_27176,N_27304);
and U29137 (N_29137,N_27682,N_26226);
nor U29138 (N_29138,N_26951,N_27069);
nand U29139 (N_29139,N_27580,N_27441);
and U29140 (N_29140,N_27558,N_27492);
xnor U29141 (N_29141,N_26842,N_27975);
nand U29142 (N_29142,N_27848,N_27582);
nand U29143 (N_29143,N_27421,N_27049);
nand U29144 (N_29144,N_27504,N_27567);
and U29145 (N_29145,N_26244,N_26171);
or U29146 (N_29146,N_27319,N_26202);
nand U29147 (N_29147,N_26540,N_26663);
nor U29148 (N_29148,N_27622,N_27172);
and U29149 (N_29149,N_27907,N_27374);
nand U29150 (N_29150,N_26318,N_26756);
nand U29151 (N_29151,N_26453,N_26864);
and U29152 (N_29152,N_26444,N_26682);
xor U29153 (N_29153,N_27521,N_26281);
nand U29154 (N_29154,N_26267,N_27957);
and U29155 (N_29155,N_27691,N_26538);
nand U29156 (N_29156,N_27838,N_27463);
xnor U29157 (N_29157,N_27498,N_26176);
or U29158 (N_29158,N_27184,N_27769);
nand U29159 (N_29159,N_27008,N_26974);
or U29160 (N_29160,N_26814,N_27955);
or U29161 (N_29161,N_27362,N_27965);
nor U29162 (N_29162,N_27402,N_26191);
or U29163 (N_29163,N_27428,N_27977);
xor U29164 (N_29164,N_26653,N_26529);
xor U29165 (N_29165,N_27858,N_27097);
or U29166 (N_29166,N_26580,N_27940);
xnor U29167 (N_29167,N_26458,N_27043);
xnor U29168 (N_29168,N_27310,N_27009);
nand U29169 (N_29169,N_27949,N_26921);
or U29170 (N_29170,N_27318,N_27545);
and U29171 (N_29171,N_27903,N_26454);
xnor U29172 (N_29172,N_26845,N_26140);
or U29173 (N_29173,N_27749,N_27841);
and U29174 (N_29174,N_26596,N_26950);
and U29175 (N_29175,N_27426,N_26990);
nor U29176 (N_29176,N_27819,N_27839);
nand U29177 (N_29177,N_26204,N_27252);
and U29178 (N_29178,N_27379,N_27880);
nor U29179 (N_29179,N_26492,N_26425);
and U29180 (N_29180,N_27150,N_27436);
xnor U29181 (N_29181,N_26911,N_26084);
xnor U29182 (N_29182,N_26438,N_26988);
or U29183 (N_29183,N_26209,N_26988);
or U29184 (N_29184,N_26104,N_26520);
nand U29185 (N_29185,N_26687,N_26578);
or U29186 (N_29186,N_26874,N_27507);
nor U29187 (N_29187,N_27077,N_26268);
nor U29188 (N_29188,N_27497,N_27036);
nor U29189 (N_29189,N_27176,N_26233);
or U29190 (N_29190,N_27481,N_27387);
and U29191 (N_29191,N_27070,N_26871);
and U29192 (N_29192,N_27580,N_27861);
and U29193 (N_29193,N_27662,N_26212);
xor U29194 (N_29194,N_27566,N_26369);
nor U29195 (N_29195,N_27540,N_26966);
nor U29196 (N_29196,N_27536,N_26359);
nor U29197 (N_29197,N_27686,N_26729);
and U29198 (N_29198,N_26977,N_26139);
or U29199 (N_29199,N_26250,N_27154);
and U29200 (N_29200,N_27767,N_27370);
xnor U29201 (N_29201,N_27003,N_26972);
and U29202 (N_29202,N_26813,N_27736);
and U29203 (N_29203,N_26863,N_26354);
or U29204 (N_29204,N_26648,N_26913);
or U29205 (N_29205,N_26713,N_27519);
nand U29206 (N_29206,N_27227,N_26904);
nand U29207 (N_29207,N_26438,N_26515);
xor U29208 (N_29208,N_26135,N_27796);
nor U29209 (N_29209,N_26530,N_27087);
nand U29210 (N_29210,N_26668,N_26754);
xor U29211 (N_29211,N_27625,N_27666);
nor U29212 (N_29212,N_26225,N_27940);
nor U29213 (N_29213,N_26667,N_26937);
xor U29214 (N_29214,N_27271,N_27948);
or U29215 (N_29215,N_27242,N_26836);
xnor U29216 (N_29216,N_27977,N_26621);
nor U29217 (N_29217,N_26435,N_26338);
and U29218 (N_29218,N_26426,N_27389);
nor U29219 (N_29219,N_27398,N_27033);
or U29220 (N_29220,N_26584,N_27500);
xnor U29221 (N_29221,N_26524,N_27982);
xnor U29222 (N_29222,N_26728,N_26680);
nor U29223 (N_29223,N_26743,N_26728);
and U29224 (N_29224,N_27695,N_26435);
nand U29225 (N_29225,N_27269,N_26274);
and U29226 (N_29226,N_26471,N_26974);
and U29227 (N_29227,N_27210,N_26067);
or U29228 (N_29228,N_27165,N_27812);
nand U29229 (N_29229,N_27037,N_27761);
nand U29230 (N_29230,N_27729,N_26317);
or U29231 (N_29231,N_27018,N_26681);
and U29232 (N_29232,N_27774,N_26787);
xor U29233 (N_29233,N_27326,N_26322);
nand U29234 (N_29234,N_27064,N_27591);
xnor U29235 (N_29235,N_27794,N_26522);
xor U29236 (N_29236,N_26368,N_27373);
nor U29237 (N_29237,N_27859,N_27132);
nor U29238 (N_29238,N_27590,N_26568);
or U29239 (N_29239,N_27120,N_26248);
nor U29240 (N_29240,N_26979,N_26509);
and U29241 (N_29241,N_26666,N_26372);
nor U29242 (N_29242,N_26721,N_27914);
xnor U29243 (N_29243,N_26175,N_27864);
xor U29244 (N_29244,N_27221,N_26183);
nand U29245 (N_29245,N_26054,N_26313);
or U29246 (N_29246,N_26585,N_26378);
and U29247 (N_29247,N_26487,N_26659);
and U29248 (N_29248,N_27205,N_26691);
or U29249 (N_29249,N_27232,N_26149);
or U29250 (N_29250,N_26254,N_27165);
and U29251 (N_29251,N_26481,N_27874);
and U29252 (N_29252,N_26090,N_27254);
or U29253 (N_29253,N_27483,N_26848);
nor U29254 (N_29254,N_26882,N_26393);
nor U29255 (N_29255,N_27469,N_27688);
xor U29256 (N_29256,N_26577,N_27167);
nand U29257 (N_29257,N_27182,N_26272);
and U29258 (N_29258,N_26048,N_27345);
nand U29259 (N_29259,N_27719,N_27132);
nor U29260 (N_29260,N_26893,N_27538);
nand U29261 (N_29261,N_26084,N_27822);
or U29262 (N_29262,N_26543,N_27841);
and U29263 (N_29263,N_27149,N_26413);
nand U29264 (N_29264,N_26274,N_26261);
or U29265 (N_29265,N_27820,N_27927);
and U29266 (N_29266,N_27237,N_27756);
or U29267 (N_29267,N_26708,N_27156);
nor U29268 (N_29268,N_27938,N_27080);
nand U29269 (N_29269,N_27613,N_26114);
and U29270 (N_29270,N_27867,N_26223);
and U29271 (N_29271,N_27153,N_27114);
or U29272 (N_29272,N_27175,N_27253);
xnor U29273 (N_29273,N_26993,N_26358);
and U29274 (N_29274,N_26558,N_27682);
xor U29275 (N_29275,N_27416,N_26843);
nand U29276 (N_29276,N_26813,N_27126);
xnor U29277 (N_29277,N_26058,N_27145);
xor U29278 (N_29278,N_27214,N_26079);
or U29279 (N_29279,N_27626,N_27478);
and U29280 (N_29280,N_26846,N_26242);
nand U29281 (N_29281,N_27894,N_27702);
nand U29282 (N_29282,N_27952,N_27159);
xnor U29283 (N_29283,N_26293,N_27606);
or U29284 (N_29284,N_26556,N_27800);
nand U29285 (N_29285,N_26480,N_26772);
nand U29286 (N_29286,N_26763,N_27254);
and U29287 (N_29287,N_26368,N_27738);
nor U29288 (N_29288,N_27519,N_27008);
nand U29289 (N_29289,N_27097,N_27212);
and U29290 (N_29290,N_26599,N_26555);
nand U29291 (N_29291,N_26828,N_27234);
and U29292 (N_29292,N_26843,N_27227);
or U29293 (N_29293,N_26342,N_26575);
or U29294 (N_29294,N_27535,N_26476);
nand U29295 (N_29295,N_26248,N_26128);
xor U29296 (N_29296,N_26091,N_27426);
and U29297 (N_29297,N_26571,N_27688);
or U29298 (N_29298,N_27614,N_27406);
xor U29299 (N_29299,N_27910,N_27039);
xor U29300 (N_29300,N_26540,N_26491);
nor U29301 (N_29301,N_27625,N_27155);
or U29302 (N_29302,N_27942,N_26978);
xor U29303 (N_29303,N_26389,N_26211);
nor U29304 (N_29304,N_26620,N_27858);
xor U29305 (N_29305,N_26157,N_27203);
or U29306 (N_29306,N_27820,N_27924);
xor U29307 (N_29307,N_26138,N_26445);
xor U29308 (N_29308,N_26627,N_27963);
or U29309 (N_29309,N_27932,N_26377);
or U29310 (N_29310,N_26043,N_27045);
and U29311 (N_29311,N_27809,N_26224);
nand U29312 (N_29312,N_27206,N_27636);
and U29313 (N_29313,N_26390,N_26284);
or U29314 (N_29314,N_26244,N_27240);
or U29315 (N_29315,N_26988,N_26027);
nand U29316 (N_29316,N_27349,N_26627);
or U29317 (N_29317,N_26351,N_26132);
or U29318 (N_29318,N_26980,N_27539);
nand U29319 (N_29319,N_27190,N_27142);
nor U29320 (N_29320,N_27844,N_27769);
xnor U29321 (N_29321,N_27035,N_27333);
nand U29322 (N_29322,N_26324,N_26224);
and U29323 (N_29323,N_26145,N_27008);
or U29324 (N_29324,N_27831,N_27746);
nor U29325 (N_29325,N_27555,N_27532);
or U29326 (N_29326,N_26032,N_27501);
xnor U29327 (N_29327,N_27661,N_27466);
and U29328 (N_29328,N_27998,N_26399);
xnor U29329 (N_29329,N_26212,N_26270);
nor U29330 (N_29330,N_27500,N_27620);
and U29331 (N_29331,N_27619,N_26542);
and U29332 (N_29332,N_26824,N_26180);
and U29333 (N_29333,N_26443,N_27818);
nor U29334 (N_29334,N_26810,N_27237);
nand U29335 (N_29335,N_27466,N_27109);
or U29336 (N_29336,N_27810,N_27349);
nand U29337 (N_29337,N_27826,N_26420);
nor U29338 (N_29338,N_26663,N_26044);
nor U29339 (N_29339,N_26145,N_26257);
xor U29340 (N_29340,N_26382,N_27518);
or U29341 (N_29341,N_27823,N_26864);
nor U29342 (N_29342,N_26353,N_27873);
nor U29343 (N_29343,N_27596,N_26803);
or U29344 (N_29344,N_26454,N_27700);
nor U29345 (N_29345,N_26757,N_26507);
and U29346 (N_29346,N_27984,N_26911);
nor U29347 (N_29347,N_27597,N_27307);
nand U29348 (N_29348,N_27402,N_26679);
and U29349 (N_29349,N_27944,N_27012);
or U29350 (N_29350,N_26677,N_27412);
nor U29351 (N_29351,N_26235,N_26386);
xnor U29352 (N_29352,N_26947,N_27295);
nand U29353 (N_29353,N_27848,N_26721);
nand U29354 (N_29354,N_27339,N_26055);
nor U29355 (N_29355,N_27019,N_26300);
nand U29356 (N_29356,N_27909,N_26626);
or U29357 (N_29357,N_26038,N_26365);
nor U29358 (N_29358,N_26819,N_27455);
nor U29359 (N_29359,N_27465,N_27126);
or U29360 (N_29360,N_26061,N_26680);
nor U29361 (N_29361,N_27738,N_27558);
or U29362 (N_29362,N_27709,N_27328);
or U29363 (N_29363,N_26570,N_26276);
and U29364 (N_29364,N_27120,N_27673);
nand U29365 (N_29365,N_26238,N_26730);
nand U29366 (N_29366,N_26092,N_27323);
and U29367 (N_29367,N_26958,N_26708);
nand U29368 (N_29368,N_26769,N_26964);
nor U29369 (N_29369,N_27260,N_26568);
nor U29370 (N_29370,N_26563,N_27079);
or U29371 (N_29371,N_26487,N_27337);
nand U29372 (N_29372,N_26063,N_27830);
nand U29373 (N_29373,N_26064,N_26012);
xor U29374 (N_29374,N_27358,N_27993);
and U29375 (N_29375,N_27956,N_27767);
nand U29376 (N_29376,N_26618,N_27326);
or U29377 (N_29377,N_26364,N_26002);
nor U29378 (N_29378,N_26779,N_27686);
nand U29379 (N_29379,N_27489,N_27016);
xor U29380 (N_29380,N_26459,N_26191);
xor U29381 (N_29381,N_27987,N_26400);
nand U29382 (N_29382,N_26934,N_26091);
and U29383 (N_29383,N_27044,N_26875);
and U29384 (N_29384,N_26736,N_27718);
or U29385 (N_29385,N_26318,N_27894);
or U29386 (N_29386,N_27340,N_27259);
xnor U29387 (N_29387,N_27964,N_27427);
xnor U29388 (N_29388,N_26322,N_27657);
nor U29389 (N_29389,N_27791,N_26859);
xnor U29390 (N_29390,N_27931,N_26015);
or U29391 (N_29391,N_26840,N_27684);
or U29392 (N_29392,N_26191,N_27436);
and U29393 (N_29393,N_26169,N_27845);
nor U29394 (N_29394,N_27773,N_27689);
nand U29395 (N_29395,N_26749,N_27467);
and U29396 (N_29396,N_27988,N_27851);
or U29397 (N_29397,N_27699,N_27978);
and U29398 (N_29398,N_27432,N_26726);
and U29399 (N_29399,N_26080,N_26770);
and U29400 (N_29400,N_27235,N_27422);
and U29401 (N_29401,N_27966,N_26842);
and U29402 (N_29402,N_26380,N_27432);
and U29403 (N_29403,N_27163,N_27170);
or U29404 (N_29404,N_26010,N_27917);
nand U29405 (N_29405,N_26241,N_27482);
xnor U29406 (N_29406,N_26069,N_26364);
nor U29407 (N_29407,N_26459,N_26547);
xnor U29408 (N_29408,N_27853,N_27349);
and U29409 (N_29409,N_26574,N_26735);
or U29410 (N_29410,N_27140,N_26946);
and U29411 (N_29411,N_27889,N_27715);
xor U29412 (N_29412,N_27183,N_27214);
or U29413 (N_29413,N_26538,N_27856);
or U29414 (N_29414,N_27327,N_27392);
nand U29415 (N_29415,N_26557,N_26194);
or U29416 (N_29416,N_26250,N_27263);
or U29417 (N_29417,N_26973,N_27048);
nand U29418 (N_29418,N_26480,N_27809);
nand U29419 (N_29419,N_26694,N_26731);
xnor U29420 (N_29420,N_26315,N_27029);
xnor U29421 (N_29421,N_26157,N_26242);
xor U29422 (N_29422,N_27680,N_26960);
nand U29423 (N_29423,N_26817,N_26095);
and U29424 (N_29424,N_27479,N_27039);
or U29425 (N_29425,N_27150,N_26033);
or U29426 (N_29426,N_27842,N_27031);
nor U29427 (N_29427,N_27516,N_26516);
nor U29428 (N_29428,N_26901,N_26536);
nand U29429 (N_29429,N_26477,N_26691);
nor U29430 (N_29430,N_26041,N_26081);
nand U29431 (N_29431,N_27069,N_26000);
nand U29432 (N_29432,N_27961,N_26607);
and U29433 (N_29433,N_27670,N_26929);
or U29434 (N_29434,N_27582,N_27299);
nand U29435 (N_29435,N_26821,N_26469);
nor U29436 (N_29436,N_26794,N_26762);
nor U29437 (N_29437,N_26573,N_26255);
xnor U29438 (N_29438,N_27119,N_27313);
nor U29439 (N_29439,N_26114,N_27436);
nor U29440 (N_29440,N_26157,N_26826);
xnor U29441 (N_29441,N_26327,N_27050);
or U29442 (N_29442,N_27834,N_26202);
xnor U29443 (N_29443,N_27889,N_26057);
and U29444 (N_29444,N_27852,N_27491);
or U29445 (N_29445,N_26687,N_26349);
or U29446 (N_29446,N_26309,N_27294);
nand U29447 (N_29447,N_26444,N_26095);
and U29448 (N_29448,N_27389,N_26475);
xnor U29449 (N_29449,N_26039,N_26102);
and U29450 (N_29450,N_26159,N_26010);
nand U29451 (N_29451,N_26752,N_26386);
nand U29452 (N_29452,N_27694,N_27003);
or U29453 (N_29453,N_27010,N_27933);
or U29454 (N_29454,N_26399,N_26374);
and U29455 (N_29455,N_26603,N_26717);
nor U29456 (N_29456,N_27018,N_26136);
and U29457 (N_29457,N_26338,N_27083);
and U29458 (N_29458,N_26409,N_26268);
nor U29459 (N_29459,N_26721,N_26641);
nand U29460 (N_29460,N_26467,N_27372);
or U29461 (N_29461,N_27209,N_27350);
xnor U29462 (N_29462,N_26539,N_26522);
nand U29463 (N_29463,N_27929,N_26490);
xor U29464 (N_29464,N_27728,N_27497);
nand U29465 (N_29465,N_26897,N_26631);
xnor U29466 (N_29466,N_26297,N_26423);
nor U29467 (N_29467,N_26795,N_26442);
and U29468 (N_29468,N_26306,N_27055);
and U29469 (N_29469,N_27202,N_27992);
nor U29470 (N_29470,N_27546,N_27284);
or U29471 (N_29471,N_27424,N_27494);
xnor U29472 (N_29472,N_26326,N_27084);
nand U29473 (N_29473,N_26493,N_26834);
and U29474 (N_29474,N_27950,N_27241);
nand U29475 (N_29475,N_26448,N_27282);
nor U29476 (N_29476,N_27603,N_26331);
nand U29477 (N_29477,N_26995,N_26591);
or U29478 (N_29478,N_26998,N_26777);
or U29479 (N_29479,N_27512,N_26711);
and U29480 (N_29480,N_27099,N_26050);
and U29481 (N_29481,N_27997,N_26132);
xor U29482 (N_29482,N_26355,N_26236);
and U29483 (N_29483,N_26636,N_27127);
nor U29484 (N_29484,N_26434,N_27536);
xnor U29485 (N_29485,N_27162,N_27649);
and U29486 (N_29486,N_27284,N_27994);
and U29487 (N_29487,N_26727,N_26696);
nor U29488 (N_29488,N_27336,N_26595);
nor U29489 (N_29489,N_27718,N_27024);
or U29490 (N_29490,N_27226,N_27567);
nand U29491 (N_29491,N_27597,N_26971);
nand U29492 (N_29492,N_26863,N_26958);
or U29493 (N_29493,N_27617,N_26188);
nor U29494 (N_29494,N_26493,N_27084);
and U29495 (N_29495,N_27270,N_27628);
xnor U29496 (N_29496,N_27008,N_27554);
and U29497 (N_29497,N_27437,N_26102);
or U29498 (N_29498,N_27358,N_26140);
or U29499 (N_29499,N_27144,N_26940);
and U29500 (N_29500,N_27024,N_27872);
nand U29501 (N_29501,N_26250,N_26265);
or U29502 (N_29502,N_26985,N_26047);
nor U29503 (N_29503,N_27926,N_27577);
nand U29504 (N_29504,N_27111,N_27134);
and U29505 (N_29505,N_26026,N_26001);
xor U29506 (N_29506,N_26892,N_26167);
and U29507 (N_29507,N_26882,N_27773);
nor U29508 (N_29508,N_26884,N_27800);
xor U29509 (N_29509,N_27588,N_27808);
nand U29510 (N_29510,N_26829,N_26954);
xnor U29511 (N_29511,N_27856,N_26732);
nand U29512 (N_29512,N_26580,N_27441);
nand U29513 (N_29513,N_26479,N_26762);
xnor U29514 (N_29514,N_27246,N_26997);
and U29515 (N_29515,N_27304,N_26522);
or U29516 (N_29516,N_26214,N_26994);
nor U29517 (N_29517,N_27528,N_26883);
and U29518 (N_29518,N_27308,N_26104);
nand U29519 (N_29519,N_27679,N_26742);
xor U29520 (N_29520,N_27009,N_26429);
or U29521 (N_29521,N_26923,N_26786);
and U29522 (N_29522,N_27917,N_27347);
or U29523 (N_29523,N_27360,N_26838);
or U29524 (N_29524,N_27948,N_27484);
and U29525 (N_29525,N_26732,N_27985);
nand U29526 (N_29526,N_27549,N_26742);
nor U29527 (N_29527,N_26547,N_27386);
or U29528 (N_29528,N_26910,N_26245);
nor U29529 (N_29529,N_26109,N_26628);
and U29530 (N_29530,N_27787,N_26697);
xor U29531 (N_29531,N_27952,N_27619);
xnor U29532 (N_29532,N_27091,N_26784);
or U29533 (N_29533,N_27671,N_26849);
nor U29534 (N_29534,N_27782,N_26293);
xnor U29535 (N_29535,N_26597,N_27588);
xor U29536 (N_29536,N_26723,N_27749);
and U29537 (N_29537,N_26458,N_27706);
nand U29538 (N_29538,N_26043,N_26447);
and U29539 (N_29539,N_27244,N_27921);
or U29540 (N_29540,N_26787,N_26715);
nand U29541 (N_29541,N_26201,N_26707);
xor U29542 (N_29542,N_27566,N_26750);
xor U29543 (N_29543,N_27199,N_27402);
nor U29544 (N_29544,N_26420,N_26654);
or U29545 (N_29545,N_27188,N_27581);
xor U29546 (N_29546,N_27058,N_26486);
xor U29547 (N_29547,N_26096,N_26133);
xor U29548 (N_29548,N_26566,N_26669);
nand U29549 (N_29549,N_26045,N_27267);
nand U29550 (N_29550,N_27706,N_27418);
nand U29551 (N_29551,N_26647,N_27396);
xnor U29552 (N_29552,N_27438,N_27233);
nand U29553 (N_29553,N_26282,N_26884);
xor U29554 (N_29554,N_27503,N_27576);
nand U29555 (N_29555,N_26746,N_27414);
nor U29556 (N_29556,N_26178,N_26824);
xnor U29557 (N_29557,N_27852,N_27120);
nand U29558 (N_29558,N_26992,N_26967);
and U29559 (N_29559,N_26825,N_27280);
or U29560 (N_29560,N_27716,N_26472);
nor U29561 (N_29561,N_27190,N_26598);
or U29562 (N_29562,N_27307,N_26524);
nor U29563 (N_29563,N_27440,N_26635);
nand U29564 (N_29564,N_27652,N_27780);
nor U29565 (N_29565,N_27904,N_26523);
or U29566 (N_29566,N_26835,N_26771);
or U29567 (N_29567,N_26829,N_26147);
or U29568 (N_29568,N_26996,N_27888);
nor U29569 (N_29569,N_27797,N_27313);
xor U29570 (N_29570,N_26984,N_26249);
nor U29571 (N_29571,N_27964,N_27879);
and U29572 (N_29572,N_27028,N_27395);
xnor U29573 (N_29573,N_27916,N_27849);
nor U29574 (N_29574,N_26244,N_26599);
and U29575 (N_29575,N_27820,N_27500);
nand U29576 (N_29576,N_27418,N_27853);
or U29577 (N_29577,N_26331,N_27500);
xnor U29578 (N_29578,N_26752,N_26594);
xor U29579 (N_29579,N_27449,N_27150);
and U29580 (N_29580,N_27159,N_27419);
xor U29581 (N_29581,N_26204,N_27462);
nor U29582 (N_29582,N_27190,N_26287);
xor U29583 (N_29583,N_26026,N_27433);
nand U29584 (N_29584,N_27105,N_27432);
nor U29585 (N_29585,N_27944,N_26495);
nor U29586 (N_29586,N_27534,N_26095);
or U29587 (N_29587,N_27876,N_26745);
and U29588 (N_29588,N_26528,N_27765);
nand U29589 (N_29589,N_26170,N_26420);
and U29590 (N_29590,N_26143,N_27407);
and U29591 (N_29591,N_27146,N_27895);
and U29592 (N_29592,N_26265,N_26954);
nand U29593 (N_29593,N_26563,N_26622);
xnor U29594 (N_29594,N_27660,N_27882);
nand U29595 (N_29595,N_26555,N_27642);
xnor U29596 (N_29596,N_27144,N_27723);
nand U29597 (N_29597,N_27405,N_26272);
or U29598 (N_29598,N_27552,N_27773);
or U29599 (N_29599,N_26546,N_26833);
nand U29600 (N_29600,N_26825,N_26787);
nand U29601 (N_29601,N_26253,N_26662);
nand U29602 (N_29602,N_26416,N_26502);
or U29603 (N_29603,N_27358,N_27284);
xnor U29604 (N_29604,N_26176,N_27144);
nor U29605 (N_29605,N_27785,N_27504);
xor U29606 (N_29606,N_27403,N_26102);
and U29607 (N_29607,N_27852,N_26759);
nand U29608 (N_29608,N_27755,N_26152);
and U29609 (N_29609,N_27038,N_26087);
xnor U29610 (N_29610,N_26459,N_26315);
nor U29611 (N_29611,N_27163,N_26023);
and U29612 (N_29612,N_27920,N_27043);
and U29613 (N_29613,N_27626,N_27204);
xor U29614 (N_29614,N_27671,N_27240);
nand U29615 (N_29615,N_26326,N_26754);
or U29616 (N_29616,N_26019,N_26081);
or U29617 (N_29617,N_26713,N_26770);
nand U29618 (N_29618,N_27325,N_27640);
and U29619 (N_29619,N_27847,N_26376);
nand U29620 (N_29620,N_27450,N_27494);
nand U29621 (N_29621,N_26390,N_26686);
and U29622 (N_29622,N_27044,N_26260);
xor U29623 (N_29623,N_27750,N_27023);
and U29624 (N_29624,N_27494,N_27462);
or U29625 (N_29625,N_27977,N_26344);
nor U29626 (N_29626,N_27456,N_26227);
or U29627 (N_29627,N_27462,N_26039);
and U29628 (N_29628,N_26473,N_26298);
xnor U29629 (N_29629,N_26261,N_26607);
or U29630 (N_29630,N_26723,N_26052);
or U29631 (N_29631,N_27373,N_27535);
nor U29632 (N_29632,N_26416,N_26431);
and U29633 (N_29633,N_27946,N_26825);
or U29634 (N_29634,N_26432,N_27059);
or U29635 (N_29635,N_26249,N_27797);
nand U29636 (N_29636,N_26421,N_27994);
nand U29637 (N_29637,N_27546,N_26773);
nor U29638 (N_29638,N_26592,N_26449);
or U29639 (N_29639,N_27697,N_27706);
or U29640 (N_29640,N_26465,N_27478);
nand U29641 (N_29641,N_27103,N_26344);
xor U29642 (N_29642,N_26555,N_27133);
xor U29643 (N_29643,N_26217,N_27248);
nor U29644 (N_29644,N_27514,N_27595);
nor U29645 (N_29645,N_26210,N_27838);
xnor U29646 (N_29646,N_26392,N_26324);
or U29647 (N_29647,N_26304,N_27559);
nor U29648 (N_29648,N_26508,N_26186);
nand U29649 (N_29649,N_27191,N_27282);
nor U29650 (N_29650,N_27496,N_27377);
nand U29651 (N_29651,N_27925,N_27849);
nand U29652 (N_29652,N_27541,N_26816);
nor U29653 (N_29653,N_26631,N_27112);
nor U29654 (N_29654,N_27071,N_27822);
nor U29655 (N_29655,N_26166,N_27633);
or U29656 (N_29656,N_26506,N_27167);
or U29657 (N_29657,N_26602,N_27134);
nand U29658 (N_29658,N_27709,N_26046);
nor U29659 (N_29659,N_26735,N_26263);
nor U29660 (N_29660,N_26101,N_26211);
nor U29661 (N_29661,N_27961,N_26357);
or U29662 (N_29662,N_27766,N_27910);
xnor U29663 (N_29663,N_26380,N_26065);
and U29664 (N_29664,N_26485,N_27429);
nor U29665 (N_29665,N_26807,N_26460);
nor U29666 (N_29666,N_27568,N_27633);
nand U29667 (N_29667,N_27920,N_27581);
xnor U29668 (N_29668,N_26970,N_27025);
nor U29669 (N_29669,N_26277,N_26500);
nand U29670 (N_29670,N_26324,N_26025);
and U29671 (N_29671,N_26376,N_26586);
or U29672 (N_29672,N_27776,N_27604);
and U29673 (N_29673,N_27260,N_27611);
nand U29674 (N_29674,N_26727,N_27830);
and U29675 (N_29675,N_26202,N_27415);
or U29676 (N_29676,N_27912,N_27223);
and U29677 (N_29677,N_27729,N_27047);
or U29678 (N_29678,N_27156,N_26049);
and U29679 (N_29679,N_27029,N_27103);
or U29680 (N_29680,N_26643,N_27341);
and U29681 (N_29681,N_26410,N_27981);
nand U29682 (N_29682,N_27650,N_27693);
nand U29683 (N_29683,N_26250,N_26837);
xnor U29684 (N_29684,N_27577,N_27811);
xor U29685 (N_29685,N_26382,N_26878);
nor U29686 (N_29686,N_26488,N_27640);
nand U29687 (N_29687,N_26074,N_26672);
nor U29688 (N_29688,N_26015,N_27840);
and U29689 (N_29689,N_27175,N_26954);
nor U29690 (N_29690,N_27733,N_27303);
nor U29691 (N_29691,N_27320,N_27388);
xor U29692 (N_29692,N_26279,N_26134);
or U29693 (N_29693,N_26007,N_27073);
nor U29694 (N_29694,N_27478,N_27753);
nand U29695 (N_29695,N_26235,N_27974);
xor U29696 (N_29696,N_27036,N_26521);
nand U29697 (N_29697,N_27882,N_26688);
xnor U29698 (N_29698,N_27455,N_26301);
nand U29699 (N_29699,N_26894,N_26050);
xor U29700 (N_29700,N_27969,N_27824);
nand U29701 (N_29701,N_26603,N_27142);
nor U29702 (N_29702,N_26203,N_26838);
nor U29703 (N_29703,N_27792,N_26893);
or U29704 (N_29704,N_27341,N_26321);
or U29705 (N_29705,N_27465,N_26321);
nand U29706 (N_29706,N_26517,N_26237);
nor U29707 (N_29707,N_26140,N_27435);
or U29708 (N_29708,N_26600,N_27013);
and U29709 (N_29709,N_27364,N_26006);
and U29710 (N_29710,N_26463,N_27473);
nand U29711 (N_29711,N_26407,N_26444);
or U29712 (N_29712,N_27333,N_26792);
nor U29713 (N_29713,N_26356,N_27219);
or U29714 (N_29714,N_27629,N_26860);
nand U29715 (N_29715,N_26394,N_26088);
or U29716 (N_29716,N_27648,N_26356);
xnor U29717 (N_29717,N_27676,N_26235);
xor U29718 (N_29718,N_27214,N_27271);
xor U29719 (N_29719,N_26650,N_26522);
or U29720 (N_29720,N_27385,N_26133);
nor U29721 (N_29721,N_27833,N_27155);
xnor U29722 (N_29722,N_27528,N_27322);
nor U29723 (N_29723,N_27059,N_26956);
xnor U29724 (N_29724,N_27764,N_26833);
or U29725 (N_29725,N_27537,N_27835);
nand U29726 (N_29726,N_27636,N_26697);
or U29727 (N_29727,N_26741,N_26374);
xnor U29728 (N_29728,N_26433,N_26608);
and U29729 (N_29729,N_26774,N_27721);
xor U29730 (N_29730,N_27058,N_26532);
or U29731 (N_29731,N_27126,N_26177);
and U29732 (N_29732,N_27051,N_27272);
xor U29733 (N_29733,N_26094,N_27351);
nand U29734 (N_29734,N_26584,N_27832);
nor U29735 (N_29735,N_26947,N_26042);
or U29736 (N_29736,N_26398,N_27237);
xor U29737 (N_29737,N_26606,N_26180);
or U29738 (N_29738,N_26548,N_27463);
and U29739 (N_29739,N_26606,N_26440);
or U29740 (N_29740,N_26423,N_27270);
nor U29741 (N_29741,N_26300,N_26214);
nor U29742 (N_29742,N_27603,N_27715);
and U29743 (N_29743,N_26084,N_27418);
and U29744 (N_29744,N_26347,N_27537);
and U29745 (N_29745,N_26551,N_27687);
nand U29746 (N_29746,N_27384,N_27120);
nand U29747 (N_29747,N_27888,N_27555);
xor U29748 (N_29748,N_26203,N_26276);
nor U29749 (N_29749,N_26552,N_26475);
nand U29750 (N_29750,N_27205,N_27866);
or U29751 (N_29751,N_27073,N_27681);
nand U29752 (N_29752,N_26456,N_26590);
and U29753 (N_29753,N_26189,N_27670);
nand U29754 (N_29754,N_26119,N_26991);
or U29755 (N_29755,N_26500,N_26967);
and U29756 (N_29756,N_26513,N_27935);
and U29757 (N_29757,N_26693,N_27649);
nand U29758 (N_29758,N_26013,N_26791);
and U29759 (N_29759,N_26852,N_26603);
xor U29760 (N_29760,N_27125,N_26445);
nor U29761 (N_29761,N_27917,N_27913);
nor U29762 (N_29762,N_26912,N_26867);
nor U29763 (N_29763,N_26749,N_26965);
nand U29764 (N_29764,N_27650,N_27664);
or U29765 (N_29765,N_26802,N_26245);
nand U29766 (N_29766,N_26951,N_27627);
nand U29767 (N_29767,N_27689,N_27379);
nor U29768 (N_29768,N_27134,N_26752);
xnor U29769 (N_29769,N_27489,N_26503);
or U29770 (N_29770,N_27751,N_26570);
nand U29771 (N_29771,N_26391,N_27472);
or U29772 (N_29772,N_27553,N_26222);
or U29773 (N_29773,N_27100,N_26942);
or U29774 (N_29774,N_26475,N_26608);
nor U29775 (N_29775,N_26265,N_26761);
xor U29776 (N_29776,N_26200,N_27924);
or U29777 (N_29777,N_26331,N_26623);
xnor U29778 (N_29778,N_26722,N_26750);
xor U29779 (N_29779,N_27708,N_27919);
and U29780 (N_29780,N_27255,N_26031);
xor U29781 (N_29781,N_26317,N_27948);
xor U29782 (N_29782,N_27398,N_26777);
nor U29783 (N_29783,N_27253,N_27892);
xor U29784 (N_29784,N_27726,N_27858);
and U29785 (N_29785,N_27970,N_26482);
nand U29786 (N_29786,N_26641,N_26450);
or U29787 (N_29787,N_26698,N_26555);
nand U29788 (N_29788,N_27786,N_26708);
or U29789 (N_29789,N_27028,N_27296);
nor U29790 (N_29790,N_26060,N_26569);
nand U29791 (N_29791,N_27115,N_27099);
xnor U29792 (N_29792,N_27662,N_27425);
xnor U29793 (N_29793,N_26791,N_27788);
nand U29794 (N_29794,N_27803,N_26413);
nor U29795 (N_29795,N_26003,N_26487);
nand U29796 (N_29796,N_26683,N_27167);
or U29797 (N_29797,N_26353,N_26777);
nand U29798 (N_29798,N_27335,N_26962);
and U29799 (N_29799,N_26017,N_26045);
xor U29800 (N_29800,N_27088,N_26229);
nor U29801 (N_29801,N_27634,N_27743);
or U29802 (N_29802,N_27052,N_26270);
xnor U29803 (N_29803,N_26509,N_26064);
nor U29804 (N_29804,N_26180,N_27287);
nand U29805 (N_29805,N_26295,N_26331);
nand U29806 (N_29806,N_26970,N_26852);
or U29807 (N_29807,N_27168,N_27434);
or U29808 (N_29808,N_26247,N_26841);
nor U29809 (N_29809,N_26533,N_27666);
or U29810 (N_29810,N_27677,N_26445);
or U29811 (N_29811,N_27147,N_27252);
nand U29812 (N_29812,N_27825,N_26949);
nor U29813 (N_29813,N_26228,N_27920);
nor U29814 (N_29814,N_27591,N_27622);
nand U29815 (N_29815,N_26432,N_27539);
and U29816 (N_29816,N_27076,N_26924);
and U29817 (N_29817,N_27645,N_26789);
nor U29818 (N_29818,N_27392,N_26997);
xnor U29819 (N_29819,N_27218,N_26378);
and U29820 (N_29820,N_27171,N_26816);
and U29821 (N_29821,N_27728,N_26744);
nor U29822 (N_29822,N_27917,N_27715);
xnor U29823 (N_29823,N_26079,N_27662);
nor U29824 (N_29824,N_27416,N_26301);
and U29825 (N_29825,N_27549,N_26654);
nor U29826 (N_29826,N_26593,N_26887);
or U29827 (N_29827,N_27811,N_27923);
and U29828 (N_29828,N_27950,N_26837);
nor U29829 (N_29829,N_26804,N_26561);
nand U29830 (N_29830,N_27355,N_26835);
nor U29831 (N_29831,N_26770,N_27384);
xor U29832 (N_29832,N_26987,N_27162);
and U29833 (N_29833,N_26022,N_27331);
or U29834 (N_29834,N_26226,N_27086);
nor U29835 (N_29835,N_27384,N_26223);
and U29836 (N_29836,N_26531,N_27854);
and U29837 (N_29837,N_27387,N_26019);
and U29838 (N_29838,N_27223,N_26687);
or U29839 (N_29839,N_26574,N_26496);
nand U29840 (N_29840,N_26152,N_27344);
nor U29841 (N_29841,N_26369,N_27378);
nand U29842 (N_29842,N_26435,N_27771);
xnor U29843 (N_29843,N_26763,N_27529);
nand U29844 (N_29844,N_27870,N_27818);
xor U29845 (N_29845,N_26201,N_27475);
xnor U29846 (N_29846,N_26597,N_26089);
nand U29847 (N_29847,N_26829,N_26726);
and U29848 (N_29848,N_27956,N_27019);
or U29849 (N_29849,N_26736,N_26157);
nand U29850 (N_29850,N_27921,N_27979);
and U29851 (N_29851,N_27364,N_27904);
nand U29852 (N_29852,N_26184,N_26636);
xor U29853 (N_29853,N_27399,N_27735);
or U29854 (N_29854,N_26639,N_27012);
and U29855 (N_29855,N_26067,N_27155);
nand U29856 (N_29856,N_26401,N_27137);
xor U29857 (N_29857,N_26287,N_27153);
and U29858 (N_29858,N_26452,N_27088);
or U29859 (N_29859,N_26297,N_26646);
or U29860 (N_29860,N_26134,N_26074);
nand U29861 (N_29861,N_26024,N_27150);
or U29862 (N_29862,N_27749,N_26864);
and U29863 (N_29863,N_26383,N_27020);
or U29864 (N_29864,N_26436,N_27283);
nor U29865 (N_29865,N_27615,N_26723);
xnor U29866 (N_29866,N_27373,N_27485);
nor U29867 (N_29867,N_27222,N_26980);
and U29868 (N_29868,N_26833,N_27345);
and U29869 (N_29869,N_27493,N_27427);
and U29870 (N_29870,N_26739,N_27510);
nor U29871 (N_29871,N_27386,N_26449);
nand U29872 (N_29872,N_26819,N_27227);
xnor U29873 (N_29873,N_27981,N_26371);
nand U29874 (N_29874,N_27075,N_27977);
and U29875 (N_29875,N_26211,N_27194);
nand U29876 (N_29876,N_27436,N_27898);
nand U29877 (N_29877,N_26143,N_26274);
and U29878 (N_29878,N_26803,N_27129);
and U29879 (N_29879,N_26715,N_27958);
or U29880 (N_29880,N_26621,N_27391);
xor U29881 (N_29881,N_27933,N_27671);
xor U29882 (N_29882,N_26776,N_27524);
and U29883 (N_29883,N_27579,N_27736);
and U29884 (N_29884,N_26204,N_26457);
or U29885 (N_29885,N_26246,N_27066);
xnor U29886 (N_29886,N_26929,N_26473);
and U29887 (N_29887,N_26544,N_26761);
or U29888 (N_29888,N_27206,N_27082);
nand U29889 (N_29889,N_26509,N_27977);
xnor U29890 (N_29890,N_26544,N_27436);
xor U29891 (N_29891,N_27822,N_26126);
xnor U29892 (N_29892,N_27847,N_27787);
nor U29893 (N_29893,N_27592,N_27969);
nor U29894 (N_29894,N_27424,N_26449);
and U29895 (N_29895,N_26745,N_26441);
nand U29896 (N_29896,N_27185,N_27571);
or U29897 (N_29897,N_26962,N_27472);
nand U29898 (N_29898,N_27067,N_27624);
nor U29899 (N_29899,N_26755,N_26557);
nor U29900 (N_29900,N_27885,N_27714);
xnor U29901 (N_29901,N_26856,N_26239);
xnor U29902 (N_29902,N_26726,N_26613);
nor U29903 (N_29903,N_26843,N_26623);
nor U29904 (N_29904,N_26040,N_27479);
nand U29905 (N_29905,N_26204,N_27323);
and U29906 (N_29906,N_27285,N_27110);
nand U29907 (N_29907,N_27774,N_26515);
or U29908 (N_29908,N_27172,N_27317);
or U29909 (N_29909,N_26933,N_27302);
nand U29910 (N_29910,N_26148,N_26329);
nand U29911 (N_29911,N_26356,N_27962);
or U29912 (N_29912,N_27599,N_27331);
and U29913 (N_29913,N_27994,N_26163);
and U29914 (N_29914,N_26821,N_26220);
and U29915 (N_29915,N_27407,N_27357);
nand U29916 (N_29916,N_27905,N_27737);
and U29917 (N_29917,N_26208,N_27307);
and U29918 (N_29918,N_26458,N_26944);
xor U29919 (N_29919,N_26641,N_27538);
nand U29920 (N_29920,N_27102,N_27371);
nor U29921 (N_29921,N_26576,N_26465);
xnor U29922 (N_29922,N_27034,N_27054);
and U29923 (N_29923,N_26817,N_27875);
or U29924 (N_29924,N_27569,N_26525);
or U29925 (N_29925,N_26184,N_27325);
xnor U29926 (N_29926,N_26544,N_26547);
nor U29927 (N_29927,N_27291,N_26850);
and U29928 (N_29928,N_27934,N_26491);
nor U29929 (N_29929,N_27957,N_27895);
or U29930 (N_29930,N_27800,N_27588);
xnor U29931 (N_29931,N_27776,N_27080);
or U29932 (N_29932,N_27633,N_26842);
or U29933 (N_29933,N_26797,N_27117);
and U29934 (N_29934,N_27454,N_27412);
and U29935 (N_29935,N_27620,N_26760);
nand U29936 (N_29936,N_27623,N_26337);
or U29937 (N_29937,N_26033,N_27246);
nor U29938 (N_29938,N_27735,N_27821);
nor U29939 (N_29939,N_27020,N_27160);
and U29940 (N_29940,N_26886,N_27930);
and U29941 (N_29941,N_27483,N_27066);
nor U29942 (N_29942,N_27414,N_27967);
nor U29943 (N_29943,N_27271,N_27185);
xor U29944 (N_29944,N_26200,N_27252);
xor U29945 (N_29945,N_26323,N_27359);
or U29946 (N_29946,N_26997,N_27731);
and U29947 (N_29947,N_27844,N_26180);
or U29948 (N_29948,N_27052,N_26152);
or U29949 (N_29949,N_26592,N_27506);
or U29950 (N_29950,N_27404,N_27141);
and U29951 (N_29951,N_26119,N_27341);
or U29952 (N_29952,N_27677,N_27854);
nor U29953 (N_29953,N_26352,N_27638);
nand U29954 (N_29954,N_26280,N_26524);
xnor U29955 (N_29955,N_27438,N_26267);
or U29956 (N_29956,N_27546,N_27401);
nor U29957 (N_29957,N_26546,N_27196);
nor U29958 (N_29958,N_26124,N_26841);
and U29959 (N_29959,N_27667,N_27488);
nand U29960 (N_29960,N_27468,N_26271);
or U29961 (N_29961,N_27732,N_27961);
xor U29962 (N_29962,N_26565,N_26640);
nor U29963 (N_29963,N_27973,N_26348);
xor U29964 (N_29964,N_26488,N_27978);
and U29965 (N_29965,N_27055,N_27300);
or U29966 (N_29966,N_27570,N_27649);
nand U29967 (N_29967,N_26984,N_26256);
xor U29968 (N_29968,N_27579,N_26867);
or U29969 (N_29969,N_27436,N_27471);
xnor U29970 (N_29970,N_27472,N_27555);
nand U29971 (N_29971,N_26211,N_26367);
or U29972 (N_29972,N_27450,N_27265);
xor U29973 (N_29973,N_26160,N_27569);
nor U29974 (N_29974,N_27215,N_26936);
xnor U29975 (N_29975,N_27278,N_26960);
nand U29976 (N_29976,N_27419,N_27602);
or U29977 (N_29977,N_26480,N_26170);
xnor U29978 (N_29978,N_26151,N_27953);
xnor U29979 (N_29979,N_26851,N_26979);
nor U29980 (N_29980,N_26222,N_26160);
xnor U29981 (N_29981,N_26520,N_26965);
xor U29982 (N_29982,N_26540,N_27758);
nor U29983 (N_29983,N_27121,N_26499);
nor U29984 (N_29984,N_26458,N_26835);
nor U29985 (N_29985,N_27121,N_27557);
xor U29986 (N_29986,N_27687,N_26783);
and U29987 (N_29987,N_26886,N_27644);
nand U29988 (N_29988,N_26371,N_27791);
and U29989 (N_29989,N_26335,N_26463);
nor U29990 (N_29990,N_26723,N_26601);
nand U29991 (N_29991,N_26992,N_27671);
xor U29992 (N_29992,N_26179,N_27285);
or U29993 (N_29993,N_26669,N_27919);
nand U29994 (N_29994,N_26635,N_26539);
and U29995 (N_29995,N_26457,N_27657);
or U29996 (N_29996,N_27323,N_27275);
and U29997 (N_29997,N_27680,N_26697);
nor U29998 (N_29998,N_26707,N_27681);
nor U29999 (N_29999,N_26199,N_26590);
xor U30000 (N_30000,N_29616,N_29163);
nor U30001 (N_30001,N_28741,N_28474);
and U30002 (N_30002,N_28936,N_28857);
nor U30003 (N_30003,N_29674,N_28003);
or U30004 (N_30004,N_28994,N_29822);
or U30005 (N_30005,N_28191,N_28672);
and U30006 (N_30006,N_29361,N_28410);
xnor U30007 (N_30007,N_29853,N_28443);
or U30008 (N_30008,N_28385,N_28128);
xor U30009 (N_30009,N_29375,N_29942);
nand U30010 (N_30010,N_28331,N_29106);
and U30011 (N_30011,N_28275,N_28313);
xor U30012 (N_30012,N_28232,N_29390);
or U30013 (N_30013,N_28406,N_28924);
or U30014 (N_30014,N_28247,N_29657);
nand U30015 (N_30015,N_29964,N_29357);
nor U30016 (N_30016,N_28438,N_29571);
xnor U30017 (N_30017,N_28527,N_28584);
xor U30018 (N_30018,N_29648,N_29503);
and U30019 (N_30019,N_29977,N_29762);
xor U30020 (N_30020,N_29703,N_29140);
or U30021 (N_30021,N_28956,N_29034);
xnor U30022 (N_30022,N_28043,N_29982);
or U30023 (N_30023,N_29259,N_29475);
xor U30024 (N_30024,N_29702,N_28881);
xor U30025 (N_30025,N_29146,N_28951);
nor U30026 (N_30026,N_29180,N_29362);
or U30027 (N_30027,N_28530,N_29410);
or U30028 (N_30028,N_29195,N_29554);
xnor U30029 (N_30029,N_29654,N_29265);
xor U30030 (N_30030,N_29452,N_28214);
nor U30031 (N_30031,N_28758,N_28146);
and U30032 (N_30032,N_29930,N_29841);
nor U30033 (N_30033,N_29539,N_28476);
and U30034 (N_30034,N_28624,N_28234);
and U30035 (N_30035,N_29007,N_28168);
nand U30036 (N_30036,N_29083,N_29851);
nor U30037 (N_30037,N_29580,N_28616);
nand U30038 (N_30038,N_29679,N_28067);
nand U30039 (N_30039,N_29024,N_28787);
nand U30040 (N_30040,N_28903,N_28480);
nor U30041 (N_30041,N_29814,N_28482);
or U30042 (N_30042,N_29791,N_28337);
xnor U30043 (N_30043,N_29189,N_28386);
and U30044 (N_30044,N_29842,N_28017);
nand U30045 (N_30045,N_29209,N_29105);
nor U30046 (N_30046,N_29520,N_28177);
nand U30047 (N_30047,N_28535,N_28422);
nand U30048 (N_30048,N_29276,N_29377);
nand U30049 (N_30049,N_29243,N_28210);
xnor U30050 (N_30050,N_28200,N_29890);
and U30051 (N_30051,N_29584,N_29775);
and U30052 (N_30052,N_28435,N_28022);
nand U30053 (N_30053,N_28496,N_29834);
nand U30054 (N_30054,N_28811,N_28409);
or U30055 (N_30055,N_28548,N_28119);
or U30056 (N_30056,N_28380,N_28834);
xor U30057 (N_30057,N_28108,N_28689);
nand U30058 (N_30058,N_29168,N_29640);
nor U30059 (N_30059,N_28273,N_29714);
xnor U30060 (N_30060,N_28105,N_29301);
nand U30061 (N_30061,N_29774,N_29961);
nand U30062 (N_30062,N_29321,N_28823);
nor U30063 (N_30063,N_29351,N_29787);
or U30064 (N_30064,N_28302,N_29058);
nor U30065 (N_30065,N_28381,N_29049);
xnor U30066 (N_30066,N_28378,N_29417);
nand U30067 (N_30067,N_28363,N_28144);
xnor U30068 (N_30068,N_29673,N_29371);
or U30069 (N_30069,N_29393,N_28849);
xnor U30070 (N_30070,N_28416,N_28166);
and U30071 (N_30071,N_29000,N_28700);
nor U30072 (N_30072,N_28341,N_28668);
nand U30073 (N_30073,N_29583,N_28193);
or U30074 (N_30074,N_29710,N_29161);
nand U30075 (N_30075,N_29650,N_28803);
and U30076 (N_30076,N_29339,N_28892);
and U30077 (N_30077,N_29440,N_28263);
nor U30078 (N_30078,N_28559,N_28449);
or U30079 (N_30079,N_28074,N_29638);
nor U30080 (N_30080,N_28454,N_29072);
nand U30081 (N_30081,N_29380,N_28224);
and U30082 (N_30082,N_29993,N_28918);
nor U30083 (N_30083,N_28844,N_28150);
or U30084 (N_30084,N_29717,N_28483);
nor U30085 (N_30085,N_29818,N_29652);
nand U30086 (N_30086,N_28019,N_28110);
nor U30087 (N_30087,N_28688,N_28753);
and U30088 (N_30088,N_28259,N_29820);
or U30089 (N_30089,N_29167,N_28012);
and U30090 (N_30090,N_28901,N_29952);
or U30091 (N_30091,N_29767,N_28008);
and U30092 (N_30092,N_28455,N_29695);
or U30093 (N_30093,N_29668,N_29701);
nor U30094 (N_30094,N_29512,N_28942);
and U30095 (N_30095,N_29581,N_29789);
nor U30096 (N_30096,N_28537,N_29399);
and U30097 (N_30097,N_29332,N_29911);
nand U30098 (N_30098,N_29847,N_28967);
xor U30099 (N_30099,N_29606,N_28033);
xnor U30100 (N_30100,N_29576,N_28452);
xnor U30101 (N_30101,N_28458,N_28159);
and U30102 (N_30102,N_29279,N_28466);
nor U30103 (N_30103,N_28106,N_29719);
nand U30104 (N_30104,N_29198,N_28592);
nor U30105 (N_30105,N_29447,N_28189);
or U30106 (N_30106,N_29014,N_28032);
and U30107 (N_30107,N_28819,N_28220);
and U30108 (N_30108,N_28913,N_28622);
xor U30109 (N_30109,N_28478,N_28240);
and U30110 (N_30110,N_29839,N_28647);
and U30111 (N_30111,N_28368,N_29376);
and U30112 (N_30112,N_29886,N_29423);
and U30113 (N_30113,N_29223,N_29988);
nand U30114 (N_30114,N_28262,N_28899);
and U30115 (N_30115,N_29159,N_28948);
or U30116 (N_30116,N_29621,N_29460);
xor U30117 (N_30117,N_29813,N_29551);
nor U30118 (N_30118,N_29166,N_28068);
nand U30119 (N_30119,N_28506,N_28860);
or U30120 (N_30120,N_28692,N_29909);
nand U30121 (N_30121,N_29645,N_29500);
and U30122 (N_30122,N_29277,N_29006);
xnor U30123 (N_30123,N_29023,N_29045);
or U30124 (N_30124,N_28366,N_28077);
and U30125 (N_30125,N_29634,N_28195);
or U30126 (N_30126,N_29941,N_28101);
or U30127 (N_30127,N_29465,N_28223);
or U30128 (N_30128,N_28118,N_29972);
xnor U30129 (N_30129,N_28710,N_28151);
and U30130 (N_30130,N_29076,N_28549);
nor U30131 (N_30131,N_28423,N_29442);
nor U30132 (N_30132,N_28255,N_29592);
nor U30133 (N_30133,N_28827,N_29412);
and U30134 (N_30134,N_28864,N_28205);
nand U30135 (N_30135,N_29996,N_28276);
or U30136 (N_30136,N_28280,N_29372);
nand U30137 (N_30137,N_29112,N_29759);
xnor U30138 (N_30138,N_28136,N_29901);
nor U30139 (N_30139,N_29086,N_28870);
or U30140 (N_30140,N_28867,N_28078);
xor U30141 (N_30141,N_29385,N_28593);
nand U30142 (N_30142,N_28635,N_29492);
and U30143 (N_30143,N_29295,N_29833);
and U30144 (N_30144,N_28939,N_29685);
xnor U30145 (N_30145,N_28374,N_28338);
xor U30146 (N_30146,N_29887,N_29698);
xnor U30147 (N_30147,N_29478,N_29816);
and U30148 (N_30148,N_28174,N_28854);
and U30149 (N_30149,N_28733,N_29724);
or U30150 (N_30150,N_28408,N_28900);
and U30151 (N_30151,N_28243,N_28612);
and U30152 (N_30152,N_28469,N_28035);
and U30153 (N_30153,N_28201,N_28349);
and U30154 (N_30154,N_28590,N_28451);
or U30155 (N_30155,N_28459,N_28011);
and U30156 (N_30156,N_29080,N_28832);
nor U30157 (N_30157,N_28375,N_28132);
or U30158 (N_30158,N_28204,N_28991);
xnor U30159 (N_30159,N_28969,N_28283);
nor U30160 (N_30160,N_29625,N_28444);
or U30161 (N_30161,N_28034,N_29020);
xnor U30162 (N_30162,N_29360,N_28016);
nand U30163 (N_30163,N_29204,N_28712);
or U30164 (N_30164,N_29677,N_28487);
or U30165 (N_30165,N_29487,N_28573);
and U30166 (N_30166,N_28081,N_29974);
nor U30167 (N_30167,N_28853,N_29329);
or U30168 (N_30168,N_29473,N_29028);
nor U30169 (N_30169,N_28437,N_28520);
nor U30170 (N_30170,N_29975,N_29530);
nor U30171 (N_30171,N_28072,N_29733);
or U30172 (N_30172,N_28206,N_28037);
or U30173 (N_30173,N_29463,N_29121);
nand U30174 (N_30174,N_29236,N_28738);
and U30175 (N_30175,N_29699,N_29016);
nand U30176 (N_30176,N_29145,N_28976);
nand U30177 (N_30177,N_29835,N_28114);
xor U30178 (N_30178,N_29256,N_28493);
and U30179 (N_30179,N_29122,N_29792);
nand U30180 (N_30180,N_29519,N_29726);
xnor U30181 (N_30181,N_28937,N_29036);
nand U30182 (N_30182,N_28258,N_29751);
or U30183 (N_30183,N_29926,N_29591);
or U30184 (N_30184,N_28794,N_28543);
xor U30185 (N_30185,N_29437,N_28165);
xor U30186 (N_30186,N_29435,N_29210);
nor U30187 (N_30187,N_29405,N_28601);
xnor U30188 (N_30188,N_29918,N_29420);
and U30189 (N_30189,N_29597,N_29418);
and U30190 (N_30190,N_29931,N_29338);
xor U30191 (N_30191,N_28868,N_28638);
xor U30192 (N_30192,N_28477,N_28286);
xor U30193 (N_30193,N_28801,N_28776);
or U30194 (N_30194,N_29090,N_29139);
xnor U30195 (N_30195,N_29365,N_28009);
xor U30196 (N_30196,N_28359,N_29451);
xor U30197 (N_30197,N_29119,N_29297);
and U30198 (N_30198,N_28046,N_29817);
or U30199 (N_30199,N_29561,N_28063);
nand U30200 (N_30200,N_29828,N_29569);
and U30201 (N_30201,N_29075,N_28307);
or U30202 (N_30202,N_29311,N_28902);
xnor U30203 (N_30203,N_28891,N_29402);
or U30204 (N_30204,N_28556,N_28236);
xor U30205 (N_30205,N_28311,N_28926);
nand U30206 (N_30206,N_28694,N_29197);
xor U30207 (N_30207,N_28203,N_29644);
nand U30208 (N_30208,N_29866,N_28364);
nor U30209 (N_30209,N_28583,N_28566);
nand U30210 (N_30210,N_29077,N_28499);
nand U30211 (N_30211,N_29507,N_28998);
and U30212 (N_30212,N_29085,N_29199);
xor U30213 (N_30213,N_29194,N_28329);
and U30214 (N_30214,N_28851,N_28065);
and U30215 (N_30215,N_28387,N_29779);
xnor U30216 (N_30216,N_29323,N_28400);
and U30217 (N_30217,N_29030,N_29336);
nand U30218 (N_30218,N_29212,N_29535);
or U30219 (N_30219,N_28097,N_29862);
nor U30220 (N_30220,N_29722,N_28277);
and U30221 (N_30221,N_28898,N_28662);
and U30222 (N_30222,N_28836,N_28190);
nor U30223 (N_30223,N_28653,N_28895);
or U30224 (N_30224,N_28884,N_28257);
and U30225 (N_30225,N_29778,N_29617);
nand U30226 (N_30226,N_28878,N_29057);
xor U30227 (N_30227,N_29432,N_28326);
or U30228 (N_30228,N_29102,N_28197);
xnor U30229 (N_30229,N_29856,N_28578);
or U30230 (N_30230,N_29671,N_28815);
nor U30231 (N_30231,N_28606,N_29560);
and U30232 (N_30232,N_28085,N_28574);
or U30233 (N_30233,N_28419,N_28781);
nand U30234 (N_30234,N_28405,N_28555);
nor U30235 (N_30235,N_28595,N_29858);
or U30236 (N_30236,N_29469,N_29428);
nand U30237 (N_30237,N_28015,N_29441);
xor U30238 (N_30238,N_28539,N_28031);
and U30239 (N_30239,N_29298,N_28157);
nor U30240 (N_30240,N_29317,N_29620);
nor U30241 (N_30241,N_29244,N_29548);
xnor U30242 (N_30242,N_29579,N_29831);
xor U30243 (N_30243,N_29656,N_28248);
or U30244 (N_30244,N_28718,N_29157);
xor U30245 (N_30245,N_29949,N_29002);
nor U30246 (N_30246,N_28564,N_28585);
xor U30247 (N_30247,N_28352,N_29837);
nand U30248 (N_30248,N_29924,N_28111);
nand U30249 (N_30249,N_28489,N_29128);
xnor U30250 (N_30250,N_29552,N_28432);
nand U30251 (N_30251,N_28941,N_29411);
xor U30252 (N_30252,N_28757,N_28615);
nand U30253 (N_30253,N_28759,N_29306);
and U30254 (N_30254,N_28825,N_28066);
nand U30255 (N_30255,N_29871,N_28663);
nor U30256 (N_30256,N_29896,N_28199);
and U30257 (N_30257,N_28347,N_28030);
nor U30258 (N_30258,N_28271,N_28877);
nand U30259 (N_30259,N_29781,N_29610);
nand U30260 (N_30260,N_28344,N_29480);
xor U30261 (N_30261,N_28427,N_29136);
nor U30262 (N_30262,N_29995,N_29590);
nand U30263 (N_30263,N_28135,N_29730);
and U30264 (N_30264,N_29476,N_28350);
and U30265 (N_30265,N_29994,N_28355);
nor U30266 (N_30266,N_29630,N_28181);
nand U30267 (N_30267,N_29809,N_29663);
nand U30268 (N_30268,N_28743,N_29596);
or U30269 (N_30269,N_29516,N_28533);
nor U30270 (N_30270,N_28163,N_28793);
and U30271 (N_30271,N_29486,N_29148);
and U30272 (N_30272,N_29300,N_29282);
nor U30273 (N_30273,N_29387,N_28785);
xor U30274 (N_30274,N_28058,N_28295);
xnor U30275 (N_30275,N_28353,N_29096);
and U30276 (N_30276,N_29917,N_28553);
or U30277 (N_30277,N_28681,N_28728);
or U30278 (N_30278,N_29494,N_29193);
and U30279 (N_30279,N_28810,N_29984);
nand U30280 (N_30280,N_29400,N_28562);
nand U30281 (N_30281,N_29665,N_29690);
nor U30282 (N_30282,N_28253,N_28029);
nand U30283 (N_30283,N_28082,N_29234);
nor U30284 (N_30284,N_29288,N_28826);
nand U30285 (N_30285,N_28383,N_28652);
or U30286 (N_30286,N_28354,N_28861);
nor U30287 (N_30287,N_29935,N_28704);
nor U30288 (N_30288,N_28429,N_28550);
nand U30289 (N_30289,N_28183,N_29047);
nand U30290 (N_30290,N_29675,N_28795);
xnor U30291 (N_30291,N_28923,N_29213);
xor U30292 (N_30292,N_29706,N_28783);
and U30293 (N_30293,N_28270,N_28701);
or U30294 (N_30294,N_29578,N_29761);
or U30295 (N_30295,N_28122,N_28202);
nor U30296 (N_30296,N_29692,N_28634);
and U30297 (N_30297,N_29861,N_28833);
and U30298 (N_30298,N_28521,N_29299);
and U30299 (N_30299,N_28510,N_28522);
nand U30300 (N_30300,N_28494,N_29992);
or U30301 (N_30301,N_29811,N_28176);
xor U30302 (N_30302,N_28325,N_29651);
nand U30303 (N_30303,N_28238,N_28880);
or U30304 (N_30304,N_29458,N_29904);
nand U30305 (N_30305,N_29766,N_28184);
and U30306 (N_30306,N_29269,N_29358);
or U30307 (N_30307,N_29855,N_28091);
or U30308 (N_30308,N_28594,N_29543);
and U30309 (N_30309,N_28125,N_29178);
xnor U30310 (N_30310,N_28044,N_29783);
and U30311 (N_30311,N_29408,N_28848);
nand U30312 (N_30312,N_29344,N_29255);
and U30313 (N_30313,N_29230,N_29369);
nor U30314 (N_30314,N_29433,N_28523);
or U30315 (N_30315,N_29490,N_29882);
xnor U30316 (N_30316,N_28401,N_29865);
nand U30317 (N_30317,N_29922,N_28279);
nor U30318 (N_30318,N_28796,N_28720);
xor U30319 (N_30319,N_29455,N_28488);
nor U30320 (N_30320,N_29723,N_28467);
nand U30321 (N_30321,N_29114,N_29015);
xor U30322 (N_30322,N_28225,N_29107);
xnor U30323 (N_30323,N_29461,N_29327);
or U30324 (N_30324,N_28628,N_28933);
xnor U30325 (N_30325,N_29350,N_28389);
nand U30326 (N_30326,N_29716,N_28698);
and U30327 (N_30327,N_29768,N_29770);
xor U30328 (N_30328,N_28096,N_29836);
nand U30329 (N_30329,N_28312,N_29248);
nand U30330 (N_30330,N_29088,N_29564);
and U30331 (N_30331,N_29222,N_29595);
nor U30332 (N_30332,N_28361,N_29175);
nand U30333 (N_30333,N_29479,N_28830);
xor U30334 (N_30334,N_28515,N_29233);
xnor U30335 (N_30335,N_28431,N_29875);
nor U30336 (N_30336,N_28099,N_28673);
nor U30337 (N_30337,N_29852,N_28852);
nand U30338 (N_30338,N_29454,N_28666);
or U30339 (N_30339,N_29293,N_29672);
and U30340 (N_30340,N_29678,N_28300);
nor U30341 (N_30341,N_29544,N_29309);
xor U30342 (N_30342,N_29424,N_28175);
and U30343 (N_30343,N_28896,N_28552);
and U30344 (N_30344,N_29720,N_28943);
nor U30345 (N_30345,N_29043,N_28514);
nand U30346 (N_30346,N_29915,N_28565);
nand U30347 (N_30347,N_28670,N_28507);
xor U30348 (N_30348,N_28570,N_29141);
xnor U30349 (N_30349,N_29735,N_29664);
nand U30350 (N_30350,N_28862,N_28740);
xnor U30351 (N_30351,N_28588,N_28968);
or U30352 (N_30352,N_29513,N_29878);
xor U30353 (N_30353,N_28428,N_28036);
and U30354 (N_30354,N_28396,N_28726);
xnor U30355 (N_30355,N_29933,N_28468);
nand U30356 (N_30356,N_29518,N_29566);
and U30357 (N_30357,N_28702,N_29147);
nor U30358 (N_30358,N_29546,N_29704);
or U30359 (N_30359,N_29796,N_28742);
nand U30360 (N_30360,N_29079,N_28139);
and U30361 (N_30361,N_28876,N_29438);
xnor U30362 (N_30362,N_28953,N_29880);
and U30363 (N_30363,N_28842,N_28858);
nor U30364 (N_30364,N_28705,N_28920);
nor U30365 (N_30365,N_29721,N_29349);
and U30366 (N_30366,N_28308,N_28264);
xor U30367 (N_30367,N_29343,N_28007);
nand U30368 (N_30368,N_28045,N_29021);
xnor U30369 (N_30369,N_28379,N_28465);
or U30370 (N_30370,N_28774,N_28054);
xnor U30371 (N_30371,N_29421,N_28642);
and U30372 (N_30372,N_29748,N_29419);
or U30373 (N_30373,N_28235,N_28789);
nor U30374 (N_30374,N_29863,N_29939);
or U30375 (N_30375,N_28501,N_29976);
xnor U30376 (N_30376,N_28450,N_28216);
nand U30377 (N_30377,N_29981,N_28241);
nor U30378 (N_30378,N_29345,N_29819);
nand U30379 (N_30379,N_29764,N_28762);
nor U30380 (N_30380,N_28597,N_29618);
nor U30381 (N_30381,N_29954,N_28840);
and U30382 (N_30382,N_28805,N_28500);
nor U30383 (N_30383,N_28148,N_29626);
nand U30384 (N_30384,N_29803,N_28026);
xnor U30385 (N_30385,N_28974,N_29927);
or U30386 (N_30386,N_29290,N_29541);
xor U30387 (N_30387,N_28390,N_29403);
nor U30388 (N_30388,N_29352,N_29348);
or U30389 (N_30389,N_29202,N_29962);
or U30390 (N_30390,N_29908,N_29967);
nor U30391 (N_30391,N_28581,N_29547);
nand U30392 (N_30392,N_28780,N_29646);
nand U30393 (N_30393,N_29502,N_28242);
xor U30394 (N_30394,N_29250,N_29874);
xnor U30395 (N_30395,N_28886,N_28472);
xnor U30396 (N_30396,N_29054,N_28348);
and U30397 (N_30397,N_28439,N_28115);
or U30398 (N_30398,N_28281,N_29124);
nor U30399 (N_30399,N_29971,N_28336);
xor U30400 (N_30400,N_28342,N_29116);
xor U30401 (N_30401,N_29963,N_28996);
and U30402 (N_30402,N_28707,N_29050);
nand U30403 (N_30403,N_28691,N_28984);
or U30404 (N_30404,N_29005,N_28186);
or U30405 (N_30405,N_28440,N_29091);
nand U30406 (N_30406,N_28430,N_29131);
nand U30407 (N_30407,N_29434,N_28524);
or U30408 (N_30408,N_29484,N_29739);
or U30409 (N_30409,N_29588,N_29200);
or U30410 (N_30410,N_28442,N_28945);
nand U30411 (N_30411,N_29039,N_28293);
nor U30412 (N_30412,N_28665,N_29048);
nor U30413 (N_30413,N_28983,N_29565);
xnor U30414 (N_30414,N_28260,N_29888);
and U30415 (N_30415,N_28576,N_29331);
and U30416 (N_30416,N_28804,N_28471);
nand U30417 (N_30417,N_28988,N_29660);
nor U30418 (N_30418,N_29600,N_28822);
xor U30419 (N_30419,N_29756,N_28481);
nand U30420 (N_30420,N_28095,N_29374);
xnor U30421 (N_30421,N_28818,N_29824);
xor U30422 (N_30422,N_29326,N_29870);
or U30423 (N_30423,N_28182,N_29613);
nor U30424 (N_30424,N_28547,N_29413);
or U30425 (N_30425,N_28233,N_29308);
or U30426 (N_30426,N_28417,N_28211);
and U30427 (N_30427,N_28103,N_29997);
and U30428 (N_30428,N_29355,N_28960);
nand U30429 (N_30429,N_28505,N_29449);
nor U30430 (N_30430,N_28502,N_28332);
nor U30431 (N_30431,N_29806,N_28403);
nand U30432 (N_30432,N_29068,N_28964);
nor U30433 (N_30433,N_28706,N_29488);
nand U30434 (N_30434,N_28971,N_28315);
or U30435 (N_30435,N_29712,N_28914);
xnor U30436 (N_30436,N_28137,N_28231);
and U30437 (N_30437,N_28630,N_29691);
and U30438 (N_30438,N_29589,N_29776);
xnor U30439 (N_30439,N_28544,N_29353);
nand U30440 (N_30440,N_29208,N_29328);
or U30441 (N_30441,N_28167,N_29249);
nand U30442 (N_30442,N_28028,N_29092);
xnor U30443 (N_30443,N_29176,N_28546);
nor U30444 (N_30444,N_28152,N_29472);
xnor U30445 (N_30445,N_29582,N_28373);
nor U30446 (N_30446,N_28305,N_29549);
and U30447 (N_30447,N_29533,N_28143);
nand U30448 (N_30448,N_28059,N_28893);
nand U30449 (N_30449,N_29046,N_28875);
nor U30450 (N_30450,N_29587,N_28256);
and U30451 (N_30451,N_28027,N_28327);
and U30452 (N_30452,N_29523,N_29680);
nand U30453 (N_30453,N_29383,N_29214);
nor U30454 (N_30454,N_29123,N_28087);
nor U30455 (N_30455,N_28786,N_28069);
nand U30456 (N_30456,N_28536,N_29602);
nor U30457 (N_30457,N_28569,N_28418);
nor U30458 (N_30458,N_28598,N_29245);
xor U30459 (N_30459,N_28394,N_28226);
or U30460 (N_30460,N_28120,N_29773);
xor U30461 (N_30461,N_29563,N_28649);
xnor U30462 (N_30462,N_29396,N_28557);
nand U30463 (N_30463,N_28798,N_29171);
nand U30464 (N_30464,N_28112,N_28749);
nor U30465 (N_30465,N_28838,N_29263);
nor U30466 (N_30466,N_28907,N_29392);
and U30467 (N_30467,N_29430,N_28445);
xor U30468 (N_30468,N_29359,N_29335);
or U30469 (N_30469,N_29099,N_28792);
or U30470 (N_30470,N_29894,N_28021);
nand U30471 (N_30471,N_28042,N_29066);
nand U30472 (N_30472,N_29743,N_28970);
nor U30473 (N_30473,N_28497,N_28679);
nand U30474 (N_30474,N_28572,N_28145);
and U30475 (N_30475,N_29676,N_28051);
and U30476 (N_30476,N_28887,N_29164);
and U30477 (N_30477,N_29903,N_28062);
and U30478 (N_30478,N_28655,N_29378);
nor U30479 (N_30479,N_29741,N_29330);
xor U30480 (N_30480,N_29524,N_29026);
or U30481 (N_30481,N_29873,N_29260);
xnor U30482 (N_30482,N_28683,N_28957);
nor U30483 (N_30483,N_28623,N_29316);
and U30484 (N_30484,N_28109,N_29854);
nand U30485 (N_30485,N_29071,N_28563);
nand U30486 (N_30486,N_29499,N_29221);
or U30487 (N_30487,N_29823,N_28614);
or U30488 (N_30488,N_28282,N_28227);
xnor U30489 (N_30489,N_28575,N_28790);
or U30490 (N_30490,N_29594,N_28334);
xor U30491 (N_30491,N_29572,N_28310);
or U30492 (N_30492,N_29556,N_29070);
and U30493 (N_30493,N_28699,N_28763);
nor U30494 (N_30494,N_29914,N_28816);
nor U30495 (N_30495,N_29219,N_28265);
nor U30496 (N_30496,N_29989,N_29444);
and U30497 (N_30497,N_28599,N_28504);
or U30498 (N_30498,N_28140,N_29558);
and U30499 (N_30499,N_28185,N_28863);
nor U30500 (N_30500,N_28979,N_28660);
xnor U30501 (N_30501,N_29179,N_29872);
nand U30502 (N_30502,N_29832,N_28987);
xnor U30503 (N_30503,N_29060,N_29999);
xor U30504 (N_30504,N_29607,N_28813);
xnor U30505 (N_30505,N_28919,N_28369);
nand U30506 (N_30506,N_29509,N_29829);
and U30507 (N_30507,N_29517,N_29797);
or U30508 (N_30508,N_28346,N_28371);
nand U30509 (N_30509,N_28617,N_28731);
nor U30510 (N_30510,N_28645,N_29757);
or U30511 (N_30511,N_29528,N_28208);
and U30512 (N_30512,N_28073,N_29641);
xnor U30513 (N_30513,N_29718,N_28222);
or U30514 (N_30514,N_28828,N_28843);
nor U30515 (N_30515,N_28797,N_29187);
xnor U30516 (N_30516,N_28739,N_29537);
and U30517 (N_30517,N_28607,N_29041);
and U30518 (N_30518,N_29525,N_28291);
or U30519 (N_30519,N_29165,N_28024);
nor U30520 (N_30520,N_29240,N_29275);
xnor U30521 (N_30521,N_28534,N_29073);
or U30522 (N_30522,N_29598,N_29363);
nand U30523 (N_30523,N_28413,N_29170);
nand U30524 (N_30524,N_29270,N_28755);
nor U30525 (N_30525,N_28484,N_28296);
nor U30526 (N_30526,N_29056,N_28098);
or U30527 (N_30527,N_28142,N_28376);
or U30528 (N_30528,N_28126,N_28318);
xor U30529 (N_30529,N_28767,N_29884);
or U30530 (N_30530,N_28356,N_28048);
nor U30531 (N_30531,N_28782,N_29881);
or U30532 (N_30532,N_29746,N_28370);
nor U30533 (N_30533,N_29422,N_28324);
and U30534 (N_30534,N_28874,N_29897);
nand U30535 (N_30535,N_29707,N_28056);
nor U30536 (N_30536,N_29337,N_28847);
nand U30537 (N_30537,N_29906,N_28362);
xnor U30538 (N_30538,N_28060,N_29785);
nor U30539 (N_30539,N_28784,N_28212);
or U30540 (N_30540,N_28959,N_29237);
or U30541 (N_30541,N_29129,N_29394);
nand U30542 (N_30542,N_29958,N_29750);
and U30543 (N_30543,N_29913,N_29429);
nand U30544 (N_30544,N_28716,N_28932);
and U30545 (N_30545,N_29902,N_28407);
and U30546 (N_30546,N_28735,N_28961);
nor U30547 (N_30547,N_28526,N_29287);
or U30548 (N_30548,N_28686,N_28927);
and U30549 (N_30549,N_29315,N_29815);
or U30550 (N_30550,N_29700,N_28160);
and U30551 (N_30551,N_28722,N_28113);
and U30552 (N_30552,N_28274,N_28053);
nand U30553 (N_30553,N_29755,N_29760);
nor U30554 (N_30554,N_29605,N_29144);
xnor U30555 (N_30555,N_28005,N_29211);
xor U30556 (N_30556,N_28064,N_29983);
xor U30557 (N_30557,N_28639,N_28475);
nand U30558 (N_30558,N_28230,N_28448);
and U30559 (N_30559,N_29169,N_29215);
and U30560 (N_30560,N_28047,N_29150);
or U30561 (N_30561,N_29133,N_28769);
nor U30562 (N_30562,N_29409,N_29108);
xor U30563 (N_30563,N_29529,N_29575);
nand U30564 (N_30564,N_29919,N_28817);
nand U30565 (N_30565,N_29312,N_29688);
xnor U30566 (N_30566,N_29303,N_28917);
or U30567 (N_30567,N_29262,N_29973);
and U30568 (N_30568,N_28746,N_28820);
or U30569 (N_30569,N_29567,N_29373);
nor U30570 (N_30570,N_29184,N_28006);
xor U30571 (N_30571,N_28049,N_28955);
and U30572 (N_30572,N_28778,N_29749);
and U30573 (N_30573,N_28567,N_29267);
or U30574 (N_30574,N_28882,N_29426);
or U30575 (N_30575,N_29912,N_29001);
or U30576 (N_30576,N_29082,N_28761);
nor U30577 (N_30577,N_28252,N_29100);
or U30578 (N_30578,N_28905,N_28978);
or U30579 (N_30579,N_28654,N_29953);
nor U30580 (N_30580,N_28107,N_29482);
or U30581 (N_30581,N_29807,N_29174);
xor U30582 (N_30582,N_28675,N_28245);
xnor U30583 (N_30583,N_29526,N_29130);
xnor U30584 (N_30584,N_29540,N_28682);
nor U30585 (N_30585,N_29231,N_28169);
nand U30586 (N_30586,N_29278,N_29181);
and U30587 (N_30587,N_28102,N_29990);
xnor U30588 (N_30588,N_29574,N_29310);
and U30589 (N_30589,N_29916,N_28316);
or U30590 (N_30590,N_29521,N_29655);
or U30591 (N_30591,N_29948,N_28589);
and U30592 (N_30592,N_28540,N_28531);
and U30593 (N_30593,N_28001,N_28285);
xor U30594 (N_30594,N_28703,N_29078);
nand U30595 (N_30595,N_28775,N_29156);
nor U30596 (N_30596,N_29857,N_28412);
xnor U30597 (N_30597,N_28173,N_29562);
xor U30598 (N_30598,N_29970,N_29740);
xor U30599 (N_30599,N_28664,N_28736);
nand U30600 (N_30600,N_28687,N_28713);
and U30601 (N_30601,N_29850,N_28719);
and U30602 (N_30602,N_29736,N_29940);
or U30603 (N_30603,N_29334,N_28278);
nor U30604 (N_30604,N_28966,N_29868);
xnor U30605 (N_30605,N_29955,N_29731);
nand U30606 (N_30606,N_29381,N_28267);
nand U30607 (N_30607,N_28425,N_29101);
nor U30608 (N_30608,N_29771,N_28963);
nor U30609 (N_30609,N_28178,N_28298);
and U30610 (N_30610,N_29273,N_29531);
nand U30611 (N_30611,N_29728,N_28631);
xor U30612 (N_30612,N_29064,N_28490);
or U30613 (N_30613,N_28290,N_28711);
nor U30614 (N_30614,N_28754,N_29055);
nand U30615 (N_30615,N_28317,N_28982);
and U30616 (N_30616,N_28023,N_29633);
xnor U30617 (N_30617,N_29155,N_28246);
nand U30618 (N_30618,N_28855,N_29804);
nor U30619 (N_30619,N_28100,N_29937);
or U30620 (N_30620,N_29876,N_29031);
and U30621 (N_30621,N_28532,N_28491);
xnor U30622 (N_30622,N_28766,N_28619);
nand U30623 (N_30623,N_28727,N_28084);
or U30624 (N_30624,N_29110,N_28392);
nand U30625 (N_30625,N_28591,N_28821);
nand U30626 (N_30626,N_28462,N_29238);
and U30627 (N_30627,N_28164,N_28288);
or U30628 (N_30628,N_29004,N_29501);
nand U30629 (N_30629,N_28990,N_28117);
and U30630 (N_30630,N_29965,N_29784);
or U30631 (N_30631,N_28123,N_28732);
nor U30632 (N_30632,N_28912,N_28975);
xnor U30633 (N_30633,N_28411,N_28678);
or U30634 (N_30634,N_29037,N_29867);
or U30635 (N_30635,N_29830,N_28577);
nor U30636 (N_30636,N_28561,N_29205);
xor U30637 (N_30637,N_29481,N_28039);
xnor U30638 (N_30638,N_29235,N_28395);
or U30639 (N_30639,N_29966,N_28717);
nand U30640 (N_30640,N_28725,N_29883);
and U30641 (N_30641,N_28734,N_29367);
and U30642 (N_30642,N_28528,N_28972);
and U30643 (N_30643,N_29257,N_29619);
xor U30644 (N_30644,N_29786,N_29154);
xnor U30645 (N_30645,N_28129,N_28340);
and U30646 (N_30646,N_29609,N_28127);
xor U30647 (N_30647,N_29220,N_28218);
and U30648 (N_30648,N_29115,N_29859);
xor U30649 (N_30649,N_29772,N_28284);
nor U30650 (N_30650,N_29318,N_29693);
nor U30651 (N_30651,N_29468,N_29511);
nor U30652 (N_30652,N_28814,N_29160);
nand U30653 (N_30653,N_29800,N_28620);
nor U30654 (N_30654,N_28721,N_29553);
xnor U30655 (N_30655,N_29207,N_28986);
xnor U30656 (N_30656,N_29289,N_28627);
nor U30657 (N_30657,N_28608,N_29109);
and U30658 (N_30658,N_29217,N_28013);
and U30659 (N_30659,N_29687,N_29603);
or U30660 (N_30660,N_29812,N_29885);
xnor U30661 (N_30661,N_29667,N_29098);
xnor U30662 (N_30662,N_29067,N_29611);
nand U30663 (N_30663,N_29386,N_28958);
nor U30664 (N_30664,N_29577,N_28339);
nor U30665 (N_30665,N_29459,N_28981);
nor U30666 (N_30666,N_28251,N_28215);
xnor U30667 (N_30667,N_29810,N_29506);
nand U30668 (N_30668,N_29126,N_29158);
and U30669 (N_30669,N_29401,N_29642);
nor U30670 (N_30670,N_28517,N_28299);
nor U30671 (N_30671,N_29765,N_29860);
nor U30672 (N_30672,N_28441,N_29347);
nand U30673 (N_30673,N_29898,N_28808);
nor U30674 (N_30674,N_28156,N_29307);
and U30675 (N_30675,N_28773,N_28560);
nand U30676 (N_30676,N_28928,N_29138);
and U30677 (N_30677,N_29113,N_29557);
or U30678 (N_30678,N_28587,N_29497);
and U30679 (N_30679,N_29956,N_28685);
nand U30680 (N_30680,N_29087,N_28723);
nand U30681 (N_30681,N_28680,N_28424);
xnor U30682 (N_30682,N_28254,N_29261);
and U30683 (N_30683,N_29969,N_29846);
xnor U30684 (N_30684,N_28659,N_28269);
nand U30685 (N_30685,N_29991,N_28292);
and U30686 (N_30686,N_29464,N_29936);
xnor U30687 (N_30687,N_29943,N_29264);
nand U30688 (N_30688,N_29732,N_29637);
and U30689 (N_30689,N_28889,N_29769);
or U30690 (N_30690,N_29191,N_29986);
or U30691 (N_30691,N_28609,N_28464);
or U30692 (N_30692,N_29135,N_28365);
xnor U30693 (N_30693,N_29684,N_29011);
or U30694 (N_30694,N_28626,N_29094);
nor U30695 (N_30695,N_29527,N_29900);
nor U30696 (N_30696,N_28398,N_28693);
or U30697 (N_30697,N_29946,N_29799);
or U30698 (N_30698,N_29869,N_29923);
xor U30699 (N_30699,N_28426,N_28791);
nand U30700 (N_30700,N_29737,N_28519);
or U30701 (N_30701,N_28397,N_29763);
and U30702 (N_30702,N_28768,N_29593);
or U30703 (N_30703,N_28198,N_28856);
xnor U30704 (N_30704,N_29322,N_29510);
nand U30705 (N_30705,N_29132,N_28596);
nor U30706 (N_30706,N_29681,N_28089);
nand U30707 (N_30707,N_29729,N_29042);
and U30708 (N_30708,N_28306,N_28509);
or U30709 (N_30709,N_29398,N_28764);
xnor U30710 (N_30710,N_28946,N_28301);
xnor U30711 (N_30711,N_29305,N_28752);
nor U30712 (N_30712,N_29320,N_29084);
nand U30713 (N_30713,N_28657,N_29185);
and U30714 (N_30714,N_29379,N_29777);
or U30715 (N_30715,N_29027,N_28977);
xnor U30716 (N_30716,N_28871,N_28367);
xnor U30717 (N_30717,N_28708,N_28131);
nor U30718 (N_30718,N_29793,N_29522);
xor U30719 (N_30719,N_29062,N_29009);
or U30720 (N_30720,N_28525,N_28083);
xnor U30721 (N_30721,N_28498,N_28973);
nor U30722 (N_30722,N_28075,N_28737);
or U30723 (N_30723,N_29008,N_28954);
xor U30724 (N_30724,N_29089,N_28690);
and U30725 (N_30725,N_29742,N_29427);
nand U30726 (N_30726,N_29864,N_29356);
xor U30727 (N_30727,N_28360,N_29798);
or U30728 (N_30728,N_29794,N_28018);
nor U30729 (N_30729,N_28812,N_29947);
xor U30730 (N_30730,N_28343,N_28134);
or U30731 (N_30731,N_29097,N_29281);
or U30732 (N_30732,N_29694,N_29570);
nand U30733 (N_30733,N_29069,N_28436);
nand U30734 (N_30734,N_29251,N_28116);
nor U30735 (N_30735,N_29493,N_28104);
or U30736 (N_30736,N_29188,N_28571);
xor U30737 (N_30737,N_28010,N_29225);
xor U30738 (N_30738,N_29294,N_28992);
xor U30739 (N_30739,N_29683,N_28625);
and U30740 (N_30740,N_29253,N_28192);
nor U30741 (N_30741,N_29384,N_29615);
nand U30742 (N_30742,N_29696,N_28086);
or U30743 (N_30743,N_29232,N_28170);
and U30744 (N_30744,N_29653,N_28092);
or U30745 (N_30745,N_29239,N_28041);
and U30746 (N_30746,N_29845,N_28696);
xnor U30747 (N_30747,N_28745,N_29025);
or U30748 (N_30748,N_28133,N_28850);
and U30749 (N_30749,N_29550,N_29889);
and U30750 (N_30750,N_29456,N_29910);
nand U30751 (N_30751,N_29040,N_29491);
nor U30752 (N_30752,N_29177,N_29446);
and U30753 (N_30753,N_28516,N_28221);
nor U30754 (N_30754,N_28513,N_29905);
and U30755 (N_30755,N_28080,N_29018);
or U30756 (N_30756,N_29725,N_28586);
nand U30757 (N_30757,N_29891,N_28228);
nand U30758 (N_30758,N_29203,N_28962);
or U30759 (N_30759,N_28772,N_29246);
xnor U30760 (N_30760,N_29670,N_29614);
nor U30761 (N_30761,N_28799,N_29629);
or U30762 (N_30762,N_28940,N_28057);
nand U30763 (N_30763,N_29978,N_28809);
nand U30764 (N_30764,N_28421,N_29934);
nand U30765 (N_30765,N_28093,N_28415);
nor U30766 (N_30766,N_29364,N_28384);
or U30767 (N_30767,N_28545,N_28730);
or U30768 (N_30768,N_28651,N_28309);
nor U30769 (N_30769,N_28002,N_29051);
xnor U30770 (N_30770,N_28038,N_29555);
and U30771 (N_30771,N_28303,N_28931);
nand U30772 (N_30772,N_28807,N_28052);
nand U30773 (N_30773,N_29149,N_29286);
and U30774 (N_30774,N_29095,N_28025);
xor U30775 (N_30775,N_29998,N_29929);
nand U30776 (N_30776,N_29708,N_29843);
nor U30777 (N_30777,N_28879,N_29536);
and U30778 (N_30778,N_28000,N_29711);
or U30779 (N_30779,N_28929,N_29052);
xnor U30780 (N_30780,N_29585,N_28894);
xor U30781 (N_30781,N_29821,N_28076);
xor U30782 (N_30782,N_29782,N_28328);
xor U30783 (N_30783,N_28644,N_28050);
xnor U30784 (N_30784,N_28289,N_29987);
nand U30785 (N_30785,N_29838,N_28207);
nor U30786 (N_30786,N_28055,N_29254);
nand U30787 (N_30787,N_29498,N_29573);
nor U30788 (N_30788,N_29182,N_29825);
nand U30789 (N_30789,N_29292,N_29907);
nand U30790 (N_30790,N_28777,N_28888);
nor U30791 (N_30791,N_28724,N_29242);
nand U30792 (N_30792,N_28070,N_29627);
or U30793 (N_30793,N_29938,N_28503);
and U30794 (N_30794,N_29532,N_29032);
nor U30795 (N_30795,N_29407,N_28995);
and U30796 (N_30796,N_28669,N_28470);
nor U30797 (N_30797,N_28319,N_28153);
nor U30798 (N_30798,N_29319,N_28382);
nor U30799 (N_30799,N_29285,N_29601);
or U30800 (N_30800,N_28079,N_28453);
nor U30801 (N_30801,N_28839,N_28297);
nor U30802 (N_30802,N_28883,N_29515);
nor U30803 (N_30803,N_28580,N_28714);
and U30804 (N_30804,N_29790,N_28287);
nor U30805 (N_30805,N_28765,N_29635);
nor U30806 (N_30806,N_29445,N_28944);
xor U30807 (N_30807,N_29877,N_29879);
and U30808 (N_30808,N_29117,N_29143);
and U30809 (N_30809,N_29622,N_28650);
nor U30810 (N_30810,N_28321,N_28121);
xor U30811 (N_30811,N_29414,N_29436);
nor U30812 (N_30812,N_28602,N_29404);
nand U30813 (N_30813,N_29397,N_28771);
nor U30814 (N_30814,N_28377,N_29747);
or U30815 (N_30815,N_29120,N_29103);
and U30816 (N_30816,N_29632,N_29495);
or U30817 (N_30817,N_29074,N_28947);
xor U30818 (N_30818,N_28872,N_28071);
nand U30819 (N_30819,N_28420,N_28434);
nand U30820 (N_30820,N_28750,N_28779);
or U30821 (N_30821,N_28770,N_28294);
xnor U30822 (N_30822,N_29980,N_28949);
xnor U30823 (N_30823,N_29059,N_29945);
or U30824 (N_30824,N_28551,N_28219);
or U30825 (N_30825,N_28250,N_29508);
nor U30826 (N_30826,N_28149,N_29647);
xor U30827 (N_30827,N_29228,N_29623);
or U30828 (N_30828,N_29186,N_28632);
or U30829 (N_30829,N_29944,N_29928);
xnor U30830 (N_30830,N_28244,N_29183);
xnor U30831 (N_30831,N_28621,N_29346);
or U30832 (N_30832,N_28161,N_29448);
nand U30833 (N_30833,N_28333,N_28921);
xnor U30834 (N_30834,N_28916,N_29604);
or U30835 (N_30835,N_29324,N_28358);
nor U30836 (N_30836,N_28268,N_28646);
nor U30837 (N_30837,N_28909,N_28829);
or U30838 (N_30838,N_29932,N_28320);
or U30839 (N_30839,N_28677,N_28446);
xor U30840 (N_30840,N_28641,N_28715);
or U30841 (N_30841,N_29545,N_28094);
xnor U30842 (N_30842,N_29559,N_29957);
nor U30843 (N_30843,N_29416,N_28806);
and U30844 (N_30844,N_29662,N_29268);
xnor U30845 (N_30845,N_29968,N_28643);
nand U30846 (N_30846,N_29192,N_29142);
xnor U30847 (N_30847,N_28180,N_28217);
or U30848 (N_30848,N_28138,N_29354);
xnor U30849 (N_30849,N_28541,N_29752);
xnor U30850 (N_30850,N_29035,N_29457);
nand U30851 (N_30851,N_28697,N_29127);
nand U30852 (N_30852,N_28399,N_28473);
nand U30853 (N_30853,N_29669,N_28460);
xnor U30854 (N_30854,N_28061,N_29467);
and U30855 (N_30855,N_28800,N_29471);
xnor U30856 (N_30856,N_29284,N_28729);
or U30857 (N_30857,N_28187,N_28674);
or U30858 (N_30858,N_28610,N_29271);
nand U30859 (N_30859,N_28744,N_28512);
and U30860 (N_30860,N_29808,N_28304);
and U30861 (N_30861,N_29659,N_29477);
xor U30862 (N_30862,N_28846,N_29805);
or U30863 (N_30863,N_29780,N_29899);
nor U30864 (N_30864,N_29950,N_29489);
nor U30865 (N_30865,N_29848,N_28314);
or U30866 (N_30866,N_29104,N_28229);
nor U30867 (N_30867,N_29496,N_28636);
nor U30868 (N_30868,N_29542,N_29689);
nand U30869 (N_30869,N_28756,N_28004);
or U30870 (N_30870,N_29391,N_28463);
or U30871 (N_30871,N_29734,N_29340);
xnor U30872 (N_30872,N_29065,N_29802);
nor U30873 (N_30873,N_29093,N_29053);
and U30874 (N_30874,N_28158,N_28040);
xnor U30875 (N_30875,N_28910,N_28020);
or U30876 (N_30876,N_29826,N_29649);
xor U30877 (N_30877,N_29801,N_28456);
nor U30878 (N_30878,N_29272,N_29162);
nand U30879 (N_30879,N_28485,N_28249);
xor U30880 (N_30880,N_28709,N_28993);
nor U30881 (N_30881,N_28357,N_29247);
xnor U30882 (N_30882,N_29727,N_28479);
or U30883 (N_30883,N_28171,N_29125);
nor U30884 (N_30884,N_28558,N_29304);
nand U30885 (N_30885,N_28934,N_29061);
nor U30886 (N_30886,N_28618,N_28667);
nor U30887 (N_30887,N_29538,N_28486);
nor U30888 (N_30888,N_28088,N_29017);
nand U30889 (N_30889,N_28196,N_29134);
xor U30890 (N_30890,N_28457,N_28014);
nor U30891 (N_30891,N_29063,N_28658);
nor U30892 (N_30892,N_29382,N_29153);
and U30893 (N_30893,N_29631,N_28090);
and U30894 (N_30894,N_29624,N_29218);
nor U30895 (N_30895,N_29568,N_28172);
and U30896 (N_30896,N_28640,N_28323);
nand U30897 (N_30897,N_29206,N_29190);
nor U30898 (N_30898,N_28950,N_29709);
xnor U30899 (N_30899,N_28613,N_28209);
xor U30900 (N_30900,N_28582,N_28147);
nor U30901 (N_30901,N_29252,N_29960);
and U30902 (N_30902,N_28661,N_28897);
and U30903 (N_30903,N_28866,N_29474);
xnor U30904 (N_30904,N_29395,N_28965);
xor U30905 (N_30905,N_28511,N_29341);
and U30906 (N_30906,N_29241,N_28999);
or U30907 (N_30907,N_29504,N_28554);
nor U30908 (N_30908,N_29754,N_28845);
nand U30909 (N_30909,N_28873,N_28179);
nand U30910 (N_30910,N_29227,N_28461);
nand U30911 (N_30911,N_28414,N_29152);
nand U30912 (N_30912,N_28684,N_28637);
or U30913 (N_30913,N_29483,N_29019);
nor U30914 (N_30914,N_28841,N_28922);
and U30915 (N_30915,N_28402,N_28261);
nand U30916 (N_30916,N_29022,N_28433);
nor U30917 (N_30917,N_29368,N_28938);
nand U30918 (N_30918,N_29443,N_28788);
and U30919 (N_30919,N_28495,N_29111);
nand U30920 (N_30920,N_29505,N_29661);
nor U30921 (N_30921,N_28925,N_29370);
and U30922 (N_30922,N_28604,N_28760);
nand U30923 (N_30923,N_28508,N_28130);
nor U30924 (N_30924,N_29425,N_29745);
and U30925 (N_30925,N_29196,N_28869);
or U30926 (N_30926,N_29849,N_28188);
and U30927 (N_30927,N_29216,N_28906);
nand U30928 (N_30928,N_29283,N_29266);
and U30929 (N_30929,N_28930,N_28372);
nand U30930 (N_30930,N_29314,N_28529);
nand U30931 (N_30931,N_29296,N_28980);
nand U30932 (N_30932,N_29013,N_29959);
nand U30933 (N_30933,N_28600,N_28272);
nor U30934 (N_30934,N_28859,N_29686);
or U30935 (N_30935,N_29366,N_29599);
nor U30936 (N_30936,N_28648,N_28802);
and U30937 (N_30937,N_29895,N_28656);
or U30938 (N_30938,N_28824,N_28162);
xnor U30939 (N_30939,N_28579,N_29302);
and U30940 (N_30940,N_28542,N_29388);
nor U30941 (N_30941,N_29389,N_29118);
or U30942 (N_30942,N_28885,N_28611);
and U30943 (N_30943,N_29636,N_29951);
nand U30944 (N_30944,N_28997,N_28633);
and U30945 (N_30945,N_29485,N_29453);
or U30946 (N_30946,N_28911,N_29466);
and U30947 (N_30947,N_28518,N_29612);
and U30948 (N_30948,N_29586,N_29033);
nand U30949 (N_30949,N_29439,N_28237);
or U30950 (N_30950,N_29151,N_28915);
and U30951 (N_30951,N_28695,N_28393);
and U30952 (N_30952,N_29081,N_29003);
or U30953 (N_30953,N_28835,N_28751);
and U30954 (N_30954,N_28155,N_29892);
nand U30955 (N_30955,N_29313,N_28908);
xnor U30956 (N_30956,N_28538,N_29280);
nor U30957 (N_30957,N_28391,N_28831);
nor U30958 (N_30958,N_29715,N_29713);
and U30959 (N_30959,N_29628,N_29201);
xnor U30960 (N_30960,N_29840,N_29038);
or U30961 (N_30961,N_28952,N_29291);
and U30962 (N_30962,N_28447,N_29705);
and U30963 (N_30963,N_29666,N_28603);
xnor U30964 (N_30964,N_29333,N_29173);
and U30965 (N_30965,N_29226,N_29979);
nor U30966 (N_30966,N_28747,N_29985);
nand U30967 (N_30967,N_28989,N_29274);
and U30968 (N_30968,N_29029,N_28239);
or U30969 (N_30969,N_28568,N_28124);
or U30970 (N_30970,N_29844,N_29608);
nand U30971 (N_30971,N_29639,N_28985);
or U30972 (N_30972,N_29744,N_29258);
and U30973 (N_30973,N_28904,N_28194);
xnor U30974 (N_30974,N_29470,N_29172);
nand U30975 (N_30975,N_28676,N_29920);
and U30976 (N_30976,N_29012,N_28605);
and U30977 (N_30977,N_29788,N_29229);
xor U30978 (N_30978,N_29893,N_29462);
nor U30979 (N_30979,N_29753,N_29406);
nand U30980 (N_30980,N_29342,N_29643);
and U30981 (N_30981,N_28671,N_29325);
nand U30982 (N_30982,N_29921,N_28629);
and U30983 (N_30983,N_29738,N_29925);
and U30984 (N_30984,N_28388,N_29827);
and U30985 (N_30985,N_29682,N_28335);
and U30986 (N_30986,N_29697,N_29044);
and U30987 (N_30987,N_28322,N_29431);
nand U30988 (N_30988,N_28351,N_28837);
or U30989 (N_30989,N_29514,N_29450);
nand U30990 (N_30990,N_28492,N_28748);
xor U30991 (N_30991,N_29137,N_28935);
nor U30992 (N_30992,N_28154,N_28266);
and U30993 (N_30993,N_29758,N_29795);
and U30994 (N_30994,N_28404,N_28890);
and U30995 (N_30995,N_29658,N_29224);
nor U30996 (N_30996,N_29415,N_28141);
nand U30997 (N_30997,N_28330,N_28213);
nor U30998 (N_30998,N_29010,N_28865);
nand U30999 (N_30999,N_28345,N_29534);
or U31000 (N_31000,N_28902,N_29641);
xnor U31001 (N_31001,N_29461,N_29449);
or U31002 (N_31002,N_28162,N_28904);
nand U31003 (N_31003,N_29595,N_29651);
xnor U31004 (N_31004,N_29742,N_29911);
or U31005 (N_31005,N_28175,N_28815);
or U31006 (N_31006,N_28071,N_28587);
xor U31007 (N_31007,N_29762,N_28732);
or U31008 (N_31008,N_28038,N_28055);
and U31009 (N_31009,N_28120,N_28662);
nand U31010 (N_31010,N_29323,N_29955);
nand U31011 (N_31011,N_29763,N_29591);
and U31012 (N_31012,N_28913,N_29483);
nor U31013 (N_31013,N_29113,N_29014);
and U31014 (N_31014,N_29638,N_28428);
nand U31015 (N_31015,N_29715,N_28711);
xor U31016 (N_31016,N_28206,N_28337);
xnor U31017 (N_31017,N_28896,N_29351);
and U31018 (N_31018,N_28988,N_28226);
nor U31019 (N_31019,N_29922,N_28724);
nor U31020 (N_31020,N_29000,N_28609);
and U31021 (N_31021,N_29940,N_29226);
and U31022 (N_31022,N_28477,N_29891);
or U31023 (N_31023,N_28726,N_29202);
xnor U31024 (N_31024,N_28601,N_28016);
xor U31025 (N_31025,N_28762,N_29991);
or U31026 (N_31026,N_29323,N_29396);
or U31027 (N_31027,N_28849,N_28208);
xor U31028 (N_31028,N_28539,N_28669);
or U31029 (N_31029,N_29752,N_28712);
and U31030 (N_31030,N_28454,N_28042);
and U31031 (N_31031,N_28734,N_28072);
or U31032 (N_31032,N_28836,N_28813);
and U31033 (N_31033,N_29779,N_28788);
nor U31034 (N_31034,N_29866,N_28558);
nor U31035 (N_31035,N_29519,N_28893);
nor U31036 (N_31036,N_29218,N_28742);
or U31037 (N_31037,N_28893,N_29162);
nand U31038 (N_31038,N_28990,N_29037);
and U31039 (N_31039,N_28999,N_28594);
xor U31040 (N_31040,N_29628,N_29078);
nor U31041 (N_31041,N_29304,N_28669);
and U31042 (N_31042,N_28423,N_28920);
and U31043 (N_31043,N_28786,N_29924);
or U31044 (N_31044,N_28212,N_28838);
nor U31045 (N_31045,N_28276,N_28678);
nor U31046 (N_31046,N_28862,N_29731);
or U31047 (N_31047,N_28517,N_28806);
and U31048 (N_31048,N_29140,N_29446);
and U31049 (N_31049,N_28803,N_29360);
nand U31050 (N_31050,N_28091,N_29189);
xnor U31051 (N_31051,N_29170,N_28336);
and U31052 (N_31052,N_28171,N_29190);
and U31053 (N_31053,N_28793,N_29660);
nand U31054 (N_31054,N_28501,N_29209);
xor U31055 (N_31055,N_29177,N_28322);
xor U31056 (N_31056,N_29623,N_29320);
nand U31057 (N_31057,N_28996,N_29035);
xor U31058 (N_31058,N_29660,N_29266);
nor U31059 (N_31059,N_29738,N_29832);
and U31060 (N_31060,N_29202,N_29528);
and U31061 (N_31061,N_29869,N_29112);
and U31062 (N_31062,N_29965,N_28951);
nor U31063 (N_31063,N_28519,N_28168);
and U31064 (N_31064,N_29535,N_28367);
nand U31065 (N_31065,N_28261,N_29706);
or U31066 (N_31066,N_29333,N_29146);
xnor U31067 (N_31067,N_28577,N_28175);
nand U31068 (N_31068,N_29985,N_28084);
and U31069 (N_31069,N_29247,N_28984);
nor U31070 (N_31070,N_28217,N_28306);
or U31071 (N_31071,N_28232,N_29198);
xnor U31072 (N_31072,N_28074,N_28001);
nor U31073 (N_31073,N_28764,N_28983);
or U31074 (N_31074,N_29174,N_29384);
and U31075 (N_31075,N_29971,N_29142);
xor U31076 (N_31076,N_29963,N_28850);
nand U31077 (N_31077,N_28386,N_29186);
and U31078 (N_31078,N_28919,N_29662);
xor U31079 (N_31079,N_28501,N_28103);
nand U31080 (N_31080,N_28859,N_28973);
nor U31081 (N_31081,N_29022,N_29842);
xor U31082 (N_31082,N_28626,N_28324);
nand U31083 (N_31083,N_28413,N_29034);
and U31084 (N_31084,N_29334,N_28265);
nor U31085 (N_31085,N_28264,N_29436);
nand U31086 (N_31086,N_28393,N_29411);
nor U31087 (N_31087,N_29428,N_29569);
nor U31088 (N_31088,N_28496,N_29006);
and U31089 (N_31089,N_29220,N_29594);
nor U31090 (N_31090,N_28367,N_28142);
nor U31091 (N_31091,N_28436,N_29440);
nand U31092 (N_31092,N_28113,N_29356);
or U31093 (N_31093,N_29960,N_29924);
nor U31094 (N_31094,N_29572,N_29841);
xor U31095 (N_31095,N_28119,N_29147);
xnor U31096 (N_31096,N_28371,N_28852);
xnor U31097 (N_31097,N_28498,N_28226);
or U31098 (N_31098,N_29055,N_28768);
and U31099 (N_31099,N_28034,N_28546);
or U31100 (N_31100,N_29296,N_28255);
nand U31101 (N_31101,N_29133,N_29697);
nand U31102 (N_31102,N_28265,N_28740);
or U31103 (N_31103,N_29660,N_29597);
nor U31104 (N_31104,N_29754,N_28164);
xor U31105 (N_31105,N_29047,N_28255);
nand U31106 (N_31106,N_29649,N_29119);
xor U31107 (N_31107,N_29768,N_29510);
or U31108 (N_31108,N_28267,N_28760);
and U31109 (N_31109,N_28615,N_28910);
nor U31110 (N_31110,N_29833,N_28768);
nor U31111 (N_31111,N_28551,N_28738);
or U31112 (N_31112,N_29408,N_29387);
or U31113 (N_31113,N_28302,N_29008);
or U31114 (N_31114,N_28788,N_28134);
and U31115 (N_31115,N_29948,N_29953);
nor U31116 (N_31116,N_29081,N_28193);
xor U31117 (N_31117,N_28774,N_29481);
or U31118 (N_31118,N_28576,N_28507);
nor U31119 (N_31119,N_28120,N_29951);
nor U31120 (N_31120,N_29471,N_29672);
nand U31121 (N_31121,N_28467,N_29657);
nor U31122 (N_31122,N_29643,N_28795);
and U31123 (N_31123,N_29699,N_28803);
xnor U31124 (N_31124,N_28411,N_28948);
or U31125 (N_31125,N_28320,N_29521);
xnor U31126 (N_31126,N_28044,N_29224);
or U31127 (N_31127,N_28802,N_29820);
or U31128 (N_31128,N_28611,N_29211);
or U31129 (N_31129,N_28278,N_28651);
or U31130 (N_31130,N_28542,N_29566);
nand U31131 (N_31131,N_29810,N_29307);
nand U31132 (N_31132,N_29865,N_28865);
xnor U31133 (N_31133,N_28718,N_28775);
nand U31134 (N_31134,N_29414,N_29413);
nand U31135 (N_31135,N_29530,N_29901);
and U31136 (N_31136,N_28005,N_29720);
or U31137 (N_31137,N_28965,N_28831);
nand U31138 (N_31138,N_28519,N_28463);
and U31139 (N_31139,N_28565,N_28625);
and U31140 (N_31140,N_28302,N_29212);
and U31141 (N_31141,N_29333,N_28600);
nand U31142 (N_31142,N_29811,N_29639);
or U31143 (N_31143,N_28670,N_29239);
nand U31144 (N_31144,N_28143,N_28654);
nor U31145 (N_31145,N_28282,N_28071);
and U31146 (N_31146,N_28085,N_28122);
xor U31147 (N_31147,N_29970,N_28537);
and U31148 (N_31148,N_29669,N_28167);
or U31149 (N_31149,N_29933,N_29092);
nand U31150 (N_31150,N_29628,N_29210);
xor U31151 (N_31151,N_28578,N_28437);
xnor U31152 (N_31152,N_28055,N_28689);
xor U31153 (N_31153,N_28042,N_29610);
or U31154 (N_31154,N_28742,N_29390);
and U31155 (N_31155,N_28903,N_28677);
and U31156 (N_31156,N_29357,N_28285);
or U31157 (N_31157,N_28894,N_29892);
and U31158 (N_31158,N_28624,N_29734);
and U31159 (N_31159,N_29764,N_29747);
or U31160 (N_31160,N_28666,N_28787);
nand U31161 (N_31161,N_29260,N_29973);
or U31162 (N_31162,N_29165,N_28368);
nand U31163 (N_31163,N_29120,N_28669);
and U31164 (N_31164,N_28901,N_28921);
nand U31165 (N_31165,N_29415,N_29307);
nand U31166 (N_31166,N_28897,N_29059);
or U31167 (N_31167,N_28598,N_28925);
nor U31168 (N_31168,N_28104,N_28184);
and U31169 (N_31169,N_29292,N_28465);
and U31170 (N_31170,N_28437,N_29895);
xnor U31171 (N_31171,N_28105,N_29093);
nand U31172 (N_31172,N_29793,N_29332);
xnor U31173 (N_31173,N_29619,N_29363);
and U31174 (N_31174,N_29159,N_29296);
nor U31175 (N_31175,N_28421,N_28409);
or U31176 (N_31176,N_28306,N_29210);
or U31177 (N_31177,N_28898,N_28853);
and U31178 (N_31178,N_29940,N_29833);
nand U31179 (N_31179,N_29959,N_29931);
or U31180 (N_31180,N_28312,N_29927);
nand U31181 (N_31181,N_28863,N_29286);
or U31182 (N_31182,N_29293,N_29385);
and U31183 (N_31183,N_28801,N_28347);
nor U31184 (N_31184,N_29467,N_28480);
and U31185 (N_31185,N_28564,N_28342);
nand U31186 (N_31186,N_28114,N_28675);
and U31187 (N_31187,N_29097,N_29478);
xor U31188 (N_31188,N_28381,N_29885);
nand U31189 (N_31189,N_29643,N_29275);
nand U31190 (N_31190,N_29680,N_28901);
or U31191 (N_31191,N_28342,N_28381);
xor U31192 (N_31192,N_28161,N_29856);
nand U31193 (N_31193,N_28421,N_29637);
or U31194 (N_31194,N_29369,N_28234);
xor U31195 (N_31195,N_29227,N_28994);
nor U31196 (N_31196,N_29933,N_29519);
nor U31197 (N_31197,N_29108,N_28673);
and U31198 (N_31198,N_28928,N_29752);
and U31199 (N_31199,N_28502,N_29335);
nor U31200 (N_31200,N_28923,N_28483);
nor U31201 (N_31201,N_28535,N_29510);
and U31202 (N_31202,N_29291,N_28141);
or U31203 (N_31203,N_29700,N_29808);
or U31204 (N_31204,N_28679,N_28405);
nor U31205 (N_31205,N_29281,N_29428);
xnor U31206 (N_31206,N_29417,N_29833);
nor U31207 (N_31207,N_29177,N_28597);
and U31208 (N_31208,N_28745,N_29185);
and U31209 (N_31209,N_29496,N_29312);
or U31210 (N_31210,N_28345,N_28717);
or U31211 (N_31211,N_28732,N_29711);
and U31212 (N_31212,N_29799,N_28803);
and U31213 (N_31213,N_29082,N_29938);
nor U31214 (N_31214,N_28932,N_28320);
nor U31215 (N_31215,N_29276,N_29534);
and U31216 (N_31216,N_28677,N_28938);
nor U31217 (N_31217,N_29321,N_29828);
nor U31218 (N_31218,N_28260,N_28727);
or U31219 (N_31219,N_29851,N_29097);
or U31220 (N_31220,N_29123,N_29371);
or U31221 (N_31221,N_28985,N_28079);
or U31222 (N_31222,N_29256,N_28114);
xnor U31223 (N_31223,N_29993,N_28529);
or U31224 (N_31224,N_28861,N_28306);
and U31225 (N_31225,N_28574,N_29080);
and U31226 (N_31226,N_29455,N_29853);
or U31227 (N_31227,N_29748,N_29365);
and U31228 (N_31228,N_29846,N_29170);
or U31229 (N_31229,N_28452,N_29642);
or U31230 (N_31230,N_29466,N_29782);
or U31231 (N_31231,N_28042,N_29628);
xnor U31232 (N_31232,N_28848,N_29276);
nor U31233 (N_31233,N_28878,N_28782);
nand U31234 (N_31234,N_28817,N_28878);
xnor U31235 (N_31235,N_29877,N_29995);
nand U31236 (N_31236,N_28446,N_29761);
xnor U31237 (N_31237,N_28213,N_29384);
nor U31238 (N_31238,N_28935,N_28813);
xnor U31239 (N_31239,N_29875,N_29309);
or U31240 (N_31240,N_28620,N_29714);
nor U31241 (N_31241,N_28575,N_29435);
nand U31242 (N_31242,N_29739,N_28302);
nand U31243 (N_31243,N_28295,N_28859);
or U31244 (N_31244,N_28746,N_28719);
or U31245 (N_31245,N_28539,N_28084);
nand U31246 (N_31246,N_29794,N_29689);
xor U31247 (N_31247,N_28965,N_28844);
nor U31248 (N_31248,N_29814,N_29693);
nand U31249 (N_31249,N_28588,N_29571);
or U31250 (N_31250,N_29440,N_29542);
and U31251 (N_31251,N_28902,N_28672);
nor U31252 (N_31252,N_29651,N_29718);
xnor U31253 (N_31253,N_29724,N_29390);
nor U31254 (N_31254,N_29502,N_29948);
or U31255 (N_31255,N_28276,N_28791);
xor U31256 (N_31256,N_29327,N_29314);
xor U31257 (N_31257,N_28844,N_29557);
or U31258 (N_31258,N_29793,N_28957);
or U31259 (N_31259,N_28180,N_29657);
and U31260 (N_31260,N_28767,N_29705);
nor U31261 (N_31261,N_29863,N_29283);
or U31262 (N_31262,N_29923,N_28659);
or U31263 (N_31263,N_29733,N_28014);
xnor U31264 (N_31264,N_29150,N_28034);
and U31265 (N_31265,N_29058,N_29198);
or U31266 (N_31266,N_28123,N_28999);
and U31267 (N_31267,N_29553,N_29248);
xor U31268 (N_31268,N_29430,N_28567);
nand U31269 (N_31269,N_28440,N_29633);
nor U31270 (N_31270,N_28907,N_28133);
and U31271 (N_31271,N_28310,N_28529);
xnor U31272 (N_31272,N_29390,N_29957);
nor U31273 (N_31273,N_28798,N_28939);
xnor U31274 (N_31274,N_29918,N_29042);
xor U31275 (N_31275,N_29713,N_29824);
or U31276 (N_31276,N_29591,N_28215);
or U31277 (N_31277,N_29490,N_29101);
and U31278 (N_31278,N_28850,N_29887);
nand U31279 (N_31279,N_29548,N_29549);
or U31280 (N_31280,N_29791,N_29523);
nand U31281 (N_31281,N_28146,N_29387);
and U31282 (N_31282,N_28795,N_29022);
nor U31283 (N_31283,N_28079,N_29301);
and U31284 (N_31284,N_29848,N_28851);
and U31285 (N_31285,N_28462,N_28439);
and U31286 (N_31286,N_28541,N_28763);
nand U31287 (N_31287,N_28397,N_28271);
or U31288 (N_31288,N_28870,N_28632);
or U31289 (N_31289,N_28670,N_29964);
nor U31290 (N_31290,N_28903,N_29505);
nor U31291 (N_31291,N_28081,N_28557);
nand U31292 (N_31292,N_28661,N_29846);
or U31293 (N_31293,N_29208,N_28721);
or U31294 (N_31294,N_28803,N_29058);
and U31295 (N_31295,N_29156,N_28765);
and U31296 (N_31296,N_29163,N_28507);
nand U31297 (N_31297,N_28771,N_28993);
and U31298 (N_31298,N_28407,N_28836);
or U31299 (N_31299,N_28600,N_29745);
or U31300 (N_31300,N_28366,N_29620);
and U31301 (N_31301,N_28971,N_28838);
nor U31302 (N_31302,N_29701,N_28698);
nand U31303 (N_31303,N_28222,N_28460);
nand U31304 (N_31304,N_28930,N_28140);
nand U31305 (N_31305,N_29507,N_28063);
nor U31306 (N_31306,N_28565,N_28824);
nand U31307 (N_31307,N_29556,N_29079);
and U31308 (N_31308,N_28551,N_28029);
nor U31309 (N_31309,N_29251,N_28845);
or U31310 (N_31310,N_29986,N_29280);
and U31311 (N_31311,N_28157,N_29947);
nor U31312 (N_31312,N_28293,N_29922);
nand U31313 (N_31313,N_28516,N_29587);
xnor U31314 (N_31314,N_28738,N_28557);
and U31315 (N_31315,N_29273,N_28975);
and U31316 (N_31316,N_28521,N_29043);
nand U31317 (N_31317,N_29465,N_29263);
xor U31318 (N_31318,N_29051,N_29791);
nand U31319 (N_31319,N_29585,N_29858);
or U31320 (N_31320,N_29322,N_28266);
or U31321 (N_31321,N_29935,N_29631);
xor U31322 (N_31322,N_29800,N_28889);
nor U31323 (N_31323,N_28035,N_28120);
xnor U31324 (N_31324,N_29887,N_28810);
or U31325 (N_31325,N_28444,N_28319);
and U31326 (N_31326,N_28752,N_28938);
and U31327 (N_31327,N_29513,N_29377);
xnor U31328 (N_31328,N_28207,N_28225);
and U31329 (N_31329,N_28164,N_28710);
and U31330 (N_31330,N_28487,N_29315);
nor U31331 (N_31331,N_28944,N_29328);
nor U31332 (N_31332,N_28923,N_28421);
or U31333 (N_31333,N_28901,N_29759);
or U31334 (N_31334,N_29502,N_29350);
or U31335 (N_31335,N_29476,N_28237);
and U31336 (N_31336,N_28681,N_29237);
xnor U31337 (N_31337,N_28622,N_28813);
or U31338 (N_31338,N_28771,N_28349);
nand U31339 (N_31339,N_28041,N_28368);
and U31340 (N_31340,N_29051,N_29676);
and U31341 (N_31341,N_29310,N_29242);
nor U31342 (N_31342,N_28783,N_28630);
nand U31343 (N_31343,N_28360,N_29100);
or U31344 (N_31344,N_28923,N_29540);
and U31345 (N_31345,N_28646,N_29114);
or U31346 (N_31346,N_29139,N_28604);
nor U31347 (N_31347,N_28401,N_28771);
xor U31348 (N_31348,N_29031,N_28957);
nand U31349 (N_31349,N_28224,N_28426);
or U31350 (N_31350,N_28922,N_28694);
and U31351 (N_31351,N_28466,N_28542);
nand U31352 (N_31352,N_28392,N_29542);
and U31353 (N_31353,N_28994,N_29596);
or U31354 (N_31354,N_29674,N_29569);
nor U31355 (N_31355,N_29375,N_29363);
xor U31356 (N_31356,N_28828,N_29741);
and U31357 (N_31357,N_29560,N_28840);
nand U31358 (N_31358,N_29408,N_29403);
xnor U31359 (N_31359,N_28812,N_29337);
or U31360 (N_31360,N_28547,N_28596);
or U31361 (N_31361,N_29367,N_28446);
and U31362 (N_31362,N_28879,N_28209);
xor U31363 (N_31363,N_28392,N_28417);
and U31364 (N_31364,N_28938,N_29985);
or U31365 (N_31365,N_29926,N_28370);
nand U31366 (N_31366,N_28632,N_29277);
nand U31367 (N_31367,N_28731,N_29184);
nor U31368 (N_31368,N_28483,N_29710);
or U31369 (N_31369,N_28458,N_29899);
nand U31370 (N_31370,N_29221,N_29688);
xor U31371 (N_31371,N_28874,N_29596);
nand U31372 (N_31372,N_28769,N_28289);
nor U31373 (N_31373,N_29607,N_28323);
and U31374 (N_31374,N_28383,N_29613);
or U31375 (N_31375,N_29927,N_28397);
and U31376 (N_31376,N_28999,N_28304);
or U31377 (N_31377,N_29084,N_28111);
or U31378 (N_31378,N_29333,N_29410);
xnor U31379 (N_31379,N_28171,N_28134);
nor U31380 (N_31380,N_28094,N_28071);
xnor U31381 (N_31381,N_28636,N_28921);
or U31382 (N_31382,N_29421,N_29041);
nor U31383 (N_31383,N_29731,N_29143);
nand U31384 (N_31384,N_28273,N_28059);
nor U31385 (N_31385,N_28632,N_28789);
nand U31386 (N_31386,N_29454,N_28262);
nand U31387 (N_31387,N_29862,N_29991);
xor U31388 (N_31388,N_28724,N_29905);
nand U31389 (N_31389,N_28540,N_28628);
nand U31390 (N_31390,N_28274,N_28177);
nor U31391 (N_31391,N_28401,N_28460);
nor U31392 (N_31392,N_29118,N_29991);
nor U31393 (N_31393,N_28729,N_29902);
xnor U31394 (N_31394,N_29059,N_28893);
or U31395 (N_31395,N_29827,N_29514);
or U31396 (N_31396,N_29132,N_28975);
xor U31397 (N_31397,N_28733,N_28119);
nor U31398 (N_31398,N_29532,N_28211);
or U31399 (N_31399,N_28674,N_28312);
or U31400 (N_31400,N_28408,N_29438);
nand U31401 (N_31401,N_29674,N_28390);
nand U31402 (N_31402,N_29253,N_29007);
and U31403 (N_31403,N_29855,N_28466);
nand U31404 (N_31404,N_29882,N_28446);
and U31405 (N_31405,N_29393,N_28165);
nand U31406 (N_31406,N_29217,N_29467);
and U31407 (N_31407,N_29690,N_29180);
nor U31408 (N_31408,N_28901,N_28082);
or U31409 (N_31409,N_29796,N_29831);
or U31410 (N_31410,N_29202,N_29747);
nand U31411 (N_31411,N_29313,N_29751);
and U31412 (N_31412,N_28329,N_29934);
and U31413 (N_31413,N_29821,N_29518);
xnor U31414 (N_31414,N_29137,N_28858);
and U31415 (N_31415,N_28140,N_28495);
xor U31416 (N_31416,N_28162,N_28331);
nor U31417 (N_31417,N_29812,N_28969);
and U31418 (N_31418,N_29580,N_28748);
nor U31419 (N_31419,N_28001,N_28458);
and U31420 (N_31420,N_29268,N_29447);
nand U31421 (N_31421,N_29035,N_29245);
nor U31422 (N_31422,N_29964,N_28140);
nand U31423 (N_31423,N_29620,N_29278);
nand U31424 (N_31424,N_28972,N_28770);
nor U31425 (N_31425,N_28022,N_29838);
and U31426 (N_31426,N_29842,N_29923);
or U31427 (N_31427,N_29326,N_29747);
nor U31428 (N_31428,N_28846,N_29434);
or U31429 (N_31429,N_28992,N_28168);
nand U31430 (N_31430,N_28146,N_28076);
nand U31431 (N_31431,N_28928,N_29949);
nand U31432 (N_31432,N_28359,N_28779);
xor U31433 (N_31433,N_28230,N_28266);
and U31434 (N_31434,N_28454,N_28552);
nand U31435 (N_31435,N_28911,N_29953);
nor U31436 (N_31436,N_29331,N_29336);
nor U31437 (N_31437,N_28126,N_28750);
and U31438 (N_31438,N_29984,N_28779);
nor U31439 (N_31439,N_28101,N_28511);
nor U31440 (N_31440,N_29837,N_29719);
and U31441 (N_31441,N_28237,N_29610);
nor U31442 (N_31442,N_29631,N_29508);
nand U31443 (N_31443,N_29239,N_28375);
nor U31444 (N_31444,N_29188,N_28598);
nor U31445 (N_31445,N_29329,N_28362);
nor U31446 (N_31446,N_29558,N_29542);
or U31447 (N_31447,N_28898,N_29204);
or U31448 (N_31448,N_28232,N_28867);
nor U31449 (N_31449,N_28319,N_28613);
or U31450 (N_31450,N_29324,N_28148);
nor U31451 (N_31451,N_29642,N_28616);
xor U31452 (N_31452,N_28486,N_28843);
or U31453 (N_31453,N_29244,N_28001);
or U31454 (N_31454,N_28967,N_29601);
xor U31455 (N_31455,N_29328,N_28772);
and U31456 (N_31456,N_28370,N_29495);
and U31457 (N_31457,N_28120,N_28695);
nand U31458 (N_31458,N_29579,N_29602);
or U31459 (N_31459,N_29501,N_29805);
or U31460 (N_31460,N_28351,N_29429);
nand U31461 (N_31461,N_29087,N_29792);
xnor U31462 (N_31462,N_29208,N_28487);
nor U31463 (N_31463,N_28922,N_29748);
or U31464 (N_31464,N_28063,N_29896);
nand U31465 (N_31465,N_28753,N_28494);
or U31466 (N_31466,N_29358,N_29088);
or U31467 (N_31467,N_29686,N_29321);
xor U31468 (N_31468,N_28987,N_29527);
or U31469 (N_31469,N_28834,N_28409);
nor U31470 (N_31470,N_28376,N_29117);
and U31471 (N_31471,N_29754,N_28279);
nand U31472 (N_31472,N_29412,N_29614);
nand U31473 (N_31473,N_29829,N_28001);
nand U31474 (N_31474,N_29825,N_28942);
and U31475 (N_31475,N_29303,N_28666);
and U31476 (N_31476,N_28009,N_28575);
nand U31477 (N_31477,N_29614,N_28128);
nor U31478 (N_31478,N_29604,N_28962);
nand U31479 (N_31479,N_28590,N_29598);
nor U31480 (N_31480,N_28846,N_29021);
and U31481 (N_31481,N_28044,N_29113);
nand U31482 (N_31482,N_28731,N_28048);
nor U31483 (N_31483,N_28559,N_28366);
nor U31484 (N_31484,N_28983,N_28303);
nand U31485 (N_31485,N_29690,N_29326);
nor U31486 (N_31486,N_29595,N_28157);
nand U31487 (N_31487,N_28031,N_28105);
nand U31488 (N_31488,N_29624,N_29779);
or U31489 (N_31489,N_28859,N_29730);
and U31490 (N_31490,N_28270,N_28843);
or U31491 (N_31491,N_28580,N_28689);
and U31492 (N_31492,N_29400,N_28234);
xnor U31493 (N_31493,N_29666,N_28727);
nand U31494 (N_31494,N_28572,N_29345);
or U31495 (N_31495,N_28746,N_28206);
xnor U31496 (N_31496,N_28603,N_29872);
and U31497 (N_31497,N_28386,N_29449);
xor U31498 (N_31498,N_29374,N_29763);
or U31499 (N_31499,N_29342,N_29809);
xnor U31500 (N_31500,N_28690,N_28237);
or U31501 (N_31501,N_28326,N_28548);
or U31502 (N_31502,N_29692,N_28608);
xnor U31503 (N_31503,N_28938,N_28561);
or U31504 (N_31504,N_28361,N_28002);
nor U31505 (N_31505,N_29108,N_29373);
nor U31506 (N_31506,N_28191,N_28576);
nor U31507 (N_31507,N_28823,N_29835);
nor U31508 (N_31508,N_28385,N_28322);
nand U31509 (N_31509,N_29678,N_28781);
or U31510 (N_31510,N_29928,N_29664);
or U31511 (N_31511,N_28170,N_29942);
nand U31512 (N_31512,N_29534,N_28051);
or U31513 (N_31513,N_28081,N_29739);
xnor U31514 (N_31514,N_28486,N_29788);
or U31515 (N_31515,N_29021,N_28104);
nor U31516 (N_31516,N_28581,N_29158);
nor U31517 (N_31517,N_29393,N_29517);
nor U31518 (N_31518,N_29555,N_29001);
and U31519 (N_31519,N_29680,N_29193);
nand U31520 (N_31520,N_29378,N_29915);
nor U31521 (N_31521,N_29034,N_28003);
or U31522 (N_31522,N_29791,N_29720);
nand U31523 (N_31523,N_29622,N_28689);
and U31524 (N_31524,N_28497,N_28397);
or U31525 (N_31525,N_28491,N_29081);
and U31526 (N_31526,N_29475,N_28863);
and U31527 (N_31527,N_28555,N_28955);
nor U31528 (N_31528,N_28491,N_29578);
or U31529 (N_31529,N_29732,N_29808);
nor U31530 (N_31530,N_29492,N_28121);
nor U31531 (N_31531,N_29634,N_29442);
and U31532 (N_31532,N_29816,N_29984);
or U31533 (N_31533,N_28024,N_28881);
nor U31534 (N_31534,N_28056,N_29437);
or U31535 (N_31535,N_28861,N_29855);
nor U31536 (N_31536,N_28400,N_28150);
nand U31537 (N_31537,N_29091,N_29844);
and U31538 (N_31538,N_29973,N_28676);
nand U31539 (N_31539,N_29868,N_28751);
nand U31540 (N_31540,N_28242,N_28892);
xor U31541 (N_31541,N_28499,N_28040);
or U31542 (N_31542,N_28405,N_29351);
and U31543 (N_31543,N_28947,N_29742);
nor U31544 (N_31544,N_28564,N_29577);
or U31545 (N_31545,N_29973,N_29065);
xnor U31546 (N_31546,N_28570,N_28391);
nand U31547 (N_31547,N_28602,N_29936);
nand U31548 (N_31548,N_29980,N_28389);
nand U31549 (N_31549,N_28935,N_28803);
or U31550 (N_31550,N_28058,N_29915);
and U31551 (N_31551,N_29178,N_29453);
and U31552 (N_31552,N_28553,N_29870);
or U31553 (N_31553,N_28646,N_29481);
or U31554 (N_31554,N_28212,N_28150);
and U31555 (N_31555,N_28329,N_29774);
and U31556 (N_31556,N_29122,N_28346);
nor U31557 (N_31557,N_28315,N_28703);
or U31558 (N_31558,N_28419,N_29924);
or U31559 (N_31559,N_28444,N_29214);
xnor U31560 (N_31560,N_28835,N_28342);
or U31561 (N_31561,N_28571,N_29353);
nor U31562 (N_31562,N_29356,N_29226);
nor U31563 (N_31563,N_29244,N_29241);
or U31564 (N_31564,N_29201,N_28679);
nand U31565 (N_31565,N_28692,N_28260);
and U31566 (N_31566,N_28880,N_29411);
xnor U31567 (N_31567,N_29417,N_29098);
or U31568 (N_31568,N_29544,N_28979);
nor U31569 (N_31569,N_28478,N_29162);
nand U31570 (N_31570,N_28919,N_29234);
nand U31571 (N_31571,N_28331,N_29791);
nand U31572 (N_31572,N_29777,N_28470);
xor U31573 (N_31573,N_28916,N_28741);
nor U31574 (N_31574,N_28062,N_29542);
xnor U31575 (N_31575,N_28849,N_28733);
or U31576 (N_31576,N_29869,N_29925);
and U31577 (N_31577,N_28335,N_29542);
and U31578 (N_31578,N_29375,N_29202);
xor U31579 (N_31579,N_29528,N_28567);
nor U31580 (N_31580,N_29661,N_28547);
nor U31581 (N_31581,N_28192,N_29133);
and U31582 (N_31582,N_29096,N_29244);
xor U31583 (N_31583,N_29223,N_29103);
nand U31584 (N_31584,N_29105,N_29192);
nand U31585 (N_31585,N_28087,N_28214);
nor U31586 (N_31586,N_29204,N_29755);
nor U31587 (N_31587,N_29229,N_28772);
nor U31588 (N_31588,N_28442,N_29863);
nand U31589 (N_31589,N_29176,N_29402);
or U31590 (N_31590,N_28981,N_29667);
xor U31591 (N_31591,N_28543,N_29436);
xnor U31592 (N_31592,N_28008,N_28458);
nand U31593 (N_31593,N_28809,N_29948);
and U31594 (N_31594,N_29294,N_28313);
or U31595 (N_31595,N_28452,N_28180);
or U31596 (N_31596,N_29530,N_28275);
and U31597 (N_31597,N_28219,N_29076);
nor U31598 (N_31598,N_28178,N_28014);
xor U31599 (N_31599,N_29896,N_28766);
or U31600 (N_31600,N_29552,N_29809);
and U31601 (N_31601,N_29459,N_29608);
nand U31602 (N_31602,N_28104,N_29167);
xor U31603 (N_31603,N_29929,N_28349);
and U31604 (N_31604,N_28424,N_29844);
nand U31605 (N_31605,N_29893,N_29357);
nor U31606 (N_31606,N_28915,N_28370);
and U31607 (N_31607,N_29045,N_29413);
or U31608 (N_31608,N_28825,N_29835);
or U31609 (N_31609,N_29059,N_29783);
nand U31610 (N_31610,N_28853,N_28269);
nand U31611 (N_31611,N_29592,N_29623);
and U31612 (N_31612,N_29550,N_28788);
nor U31613 (N_31613,N_29280,N_29810);
nand U31614 (N_31614,N_29259,N_28249);
and U31615 (N_31615,N_29501,N_28293);
or U31616 (N_31616,N_28224,N_29418);
or U31617 (N_31617,N_28156,N_29142);
nand U31618 (N_31618,N_28661,N_29933);
and U31619 (N_31619,N_28100,N_28610);
or U31620 (N_31620,N_28208,N_28743);
xor U31621 (N_31621,N_29147,N_29211);
xor U31622 (N_31622,N_28198,N_29823);
or U31623 (N_31623,N_29843,N_28956);
xor U31624 (N_31624,N_28887,N_29542);
xnor U31625 (N_31625,N_28302,N_28268);
nor U31626 (N_31626,N_29782,N_28582);
nand U31627 (N_31627,N_29442,N_29872);
nor U31628 (N_31628,N_29537,N_28014);
and U31629 (N_31629,N_28256,N_28664);
and U31630 (N_31630,N_28668,N_29928);
xnor U31631 (N_31631,N_28092,N_29134);
nand U31632 (N_31632,N_29707,N_29645);
or U31633 (N_31633,N_28516,N_28673);
or U31634 (N_31634,N_28982,N_28230);
nand U31635 (N_31635,N_28453,N_29031);
and U31636 (N_31636,N_29686,N_28669);
and U31637 (N_31637,N_29431,N_29618);
nand U31638 (N_31638,N_28944,N_28111);
and U31639 (N_31639,N_29675,N_29395);
nand U31640 (N_31640,N_28877,N_28795);
nor U31641 (N_31641,N_29969,N_29654);
nor U31642 (N_31642,N_29817,N_28934);
and U31643 (N_31643,N_29662,N_28885);
or U31644 (N_31644,N_28950,N_29398);
nor U31645 (N_31645,N_28576,N_28356);
or U31646 (N_31646,N_28338,N_28870);
xnor U31647 (N_31647,N_29860,N_29350);
or U31648 (N_31648,N_28257,N_29693);
or U31649 (N_31649,N_29809,N_29716);
or U31650 (N_31650,N_29692,N_28249);
or U31651 (N_31651,N_29349,N_28565);
nand U31652 (N_31652,N_29475,N_29740);
nand U31653 (N_31653,N_28811,N_28923);
or U31654 (N_31654,N_28713,N_28143);
and U31655 (N_31655,N_29289,N_28262);
or U31656 (N_31656,N_29004,N_28153);
xnor U31657 (N_31657,N_28121,N_29047);
nor U31658 (N_31658,N_28173,N_29553);
or U31659 (N_31659,N_29575,N_29754);
nor U31660 (N_31660,N_28370,N_29729);
nand U31661 (N_31661,N_29049,N_28845);
xnor U31662 (N_31662,N_28013,N_29584);
nor U31663 (N_31663,N_29966,N_29816);
or U31664 (N_31664,N_29737,N_29497);
and U31665 (N_31665,N_29777,N_29982);
and U31666 (N_31666,N_28607,N_28945);
xor U31667 (N_31667,N_28997,N_28105);
and U31668 (N_31668,N_29778,N_28527);
xnor U31669 (N_31669,N_29595,N_29064);
and U31670 (N_31670,N_29051,N_29363);
xor U31671 (N_31671,N_29083,N_28930);
or U31672 (N_31672,N_28311,N_29876);
or U31673 (N_31673,N_29695,N_28784);
and U31674 (N_31674,N_29133,N_29946);
xnor U31675 (N_31675,N_28044,N_28604);
nand U31676 (N_31676,N_28389,N_29855);
nand U31677 (N_31677,N_28036,N_29717);
nand U31678 (N_31678,N_29955,N_28553);
nand U31679 (N_31679,N_28958,N_28955);
xor U31680 (N_31680,N_28493,N_29676);
nand U31681 (N_31681,N_28779,N_28170);
or U31682 (N_31682,N_28639,N_29832);
nand U31683 (N_31683,N_29056,N_29102);
nor U31684 (N_31684,N_28609,N_29476);
or U31685 (N_31685,N_28024,N_29547);
nand U31686 (N_31686,N_29353,N_29539);
or U31687 (N_31687,N_28835,N_29278);
or U31688 (N_31688,N_28346,N_28844);
nand U31689 (N_31689,N_28420,N_29877);
and U31690 (N_31690,N_29931,N_28563);
nor U31691 (N_31691,N_28437,N_29167);
nand U31692 (N_31692,N_29420,N_28142);
nor U31693 (N_31693,N_29780,N_28088);
nand U31694 (N_31694,N_28561,N_29921);
and U31695 (N_31695,N_28825,N_28646);
and U31696 (N_31696,N_28782,N_28812);
and U31697 (N_31697,N_28546,N_29104);
nor U31698 (N_31698,N_28952,N_29001);
nor U31699 (N_31699,N_29562,N_28510);
nand U31700 (N_31700,N_28245,N_29618);
or U31701 (N_31701,N_28982,N_28671);
and U31702 (N_31702,N_29854,N_28536);
nand U31703 (N_31703,N_28143,N_29889);
or U31704 (N_31704,N_29346,N_29287);
xor U31705 (N_31705,N_29281,N_28438);
xnor U31706 (N_31706,N_28791,N_28053);
and U31707 (N_31707,N_28484,N_28307);
and U31708 (N_31708,N_28727,N_29948);
or U31709 (N_31709,N_29267,N_28931);
or U31710 (N_31710,N_29426,N_28728);
xor U31711 (N_31711,N_29086,N_29568);
xnor U31712 (N_31712,N_28934,N_29690);
or U31713 (N_31713,N_29241,N_29859);
nand U31714 (N_31714,N_28386,N_28567);
or U31715 (N_31715,N_28191,N_29086);
and U31716 (N_31716,N_28573,N_28668);
nor U31717 (N_31717,N_29680,N_28643);
or U31718 (N_31718,N_28277,N_28411);
xnor U31719 (N_31719,N_29662,N_29179);
and U31720 (N_31720,N_29633,N_29880);
and U31721 (N_31721,N_28740,N_28566);
or U31722 (N_31722,N_29610,N_28461);
and U31723 (N_31723,N_28178,N_28768);
or U31724 (N_31724,N_29546,N_28204);
xnor U31725 (N_31725,N_29054,N_29724);
nand U31726 (N_31726,N_29999,N_29871);
nand U31727 (N_31727,N_29418,N_28980);
nand U31728 (N_31728,N_28667,N_29534);
nor U31729 (N_31729,N_28284,N_29004);
or U31730 (N_31730,N_28896,N_29709);
nor U31731 (N_31731,N_29695,N_29808);
or U31732 (N_31732,N_29807,N_28712);
or U31733 (N_31733,N_28140,N_29146);
xnor U31734 (N_31734,N_29735,N_28657);
nor U31735 (N_31735,N_28419,N_29414);
and U31736 (N_31736,N_29638,N_28974);
xnor U31737 (N_31737,N_29095,N_29763);
xnor U31738 (N_31738,N_29458,N_29761);
nand U31739 (N_31739,N_29174,N_29064);
xnor U31740 (N_31740,N_28688,N_28608);
or U31741 (N_31741,N_29421,N_28710);
or U31742 (N_31742,N_29882,N_29480);
xor U31743 (N_31743,N_28669,N_28918);
nor U31744 (N_31744,N_28459,N_28340);
nand U31745 (N_31745,N_28348,N_29782);
and U31746 (N_31746,N_28162,N_29976);
nand U31747 (N_31747,N_28590,N_29194);
or U31748 (N_31748,N_29832,N_28562);
and U31749 (N_31749,N_29337,N_28770);
nor U31750 (N_31750,N_28612,N_28562);
or U31751 (N_31751,N_29615,N_28465);
nand U31752 (N_31752,N_29587,N_29881);
and U31753 (N_31753,N_28025,N_28087);
xnor U31754 (N_31754,N_29775,N_28075);
nand U31755 (N_31755,N_29234,N_28077);
or U31756 (N_31756,N_28099,N_29412);
nor U31757 (N_31757,N_29100,N_29521);
xnor U31758 (N_31758,N_28615,N_28163);
and U31759 (N_31759,N_29432,N_28572);
xor U31760 (N_31760,N_28252,N_29001);
nor U31761 (N_31761,N_28080,N_29235);
or U31762 (N_31762,N_29159,N_28313);
nand U31763 (N_31763,N_29894,N_29697);
nor U31764 (N_31764,N_29839,N_29225);
and U31765 (N_31765,N_29872,N_29661);
and U31766 (N_31766,N_29268,N_29571);
nor U31767 (N_31767,N_29855,N_28365);
nand U31768 (N_31768,N_29204,N_28506);
and U31769 (N_31769,N_28345,N_29387);
or U31770 (N_31770,N_28019,N_29956);
xnor U31771 (N_31771,N_28235,N_29967);
nand U31772 (N_31772,N_29787,N_29484);
or U31773 (N_31773,N_29839,N_29963);
xnor U31774 (N_31774,N_29814,N_28820);
or U31775 (N_31775,N_29039,N_29557);
or U31776 (N_31776,N_28097,N_29949);
or U31777 (N_31777,N_28816,N_29012);
nand U31778 (N_31778,N_29755,N_28407);
and U31779 (N_31779,N_28682,N_28027);
or U31780 (N_31780,N_29110,N_29984);
xor U31781 (N_31781,N_28454,N_28186);
xor U31782 (N_31782,N_29268,N_29786);
nor U31783 (N_31783,N_28205,N_28073);
nor U31784 (N_31784,N_29621,N_28415);
nand U31785 (N_31785,N_29434,N_28621);
nor U31786 (N_31786,N_29108,N_28192);
xor U31787 (N_31787,N_28892,N_28495);
and U31788 (N_31788,N_28532,N_28696);
and U31789 (N_31789,N_29757,N_29218);
xor U31790 (N_31790,N_28912,N_29367);
xnor U31791 (N_31791,N_29397,N_29803);
or U31792 (N_31792,N_28199,N_29239);
nor U31793 (N_31793,N_29460,N_29646);
nor U31794 (N_31794,N_29303,N_29934);
nand U31795 (N_31795,N_28321,N_28667);
xor U31796 (N_31796,N_29963,N_28446);
nor U31797 (N_31797,N_28427,N_29781);
nand U31798 (N_31798,N_29241,N_28980);
xnor U31799 (N_31799,N_28974,N_29337);
or U31800 (N_31800,N_28668,N_29054);
nand U31801 (N_31801,N_28073,N_28272);
xor U31802 (N_31802,N_28274,N_29836);
xnor U31803 (N_31803,N_28566,N_28910);
or U31804 (N_31804,N_28816,N_28187);
or U31805 (N_31805,N_29579,N_28347);
xor U31806 (N_31806,N_29031,N_29554);
or U31807 (N_31807,N_28601,N_28168);
nand U31808 (N_31808,N_28682,N_28699);
or U31809 (N_31809,N_29679,N_29615);
xnor U31810 (N_31810,N_29002,N_29308);
and U31811 (N_31811,N_28076,N_28021);
xor U31812 (N_31812,N_28178,N_29473);
nor U31813 (N_31813,N_29666,N_28251);
or U31814 (N_31814,N_28843,N_28513);
or U31815 (N_31815,N_29575,N_28518);
xor U31816 (N_31816,N_28718,N_28748);
nand U31817 (N_31817,N_29872,N_28458);
xor U31818 (N_31818,N_28136,N_29603);
or U31819 (N_31819,N_28545,N_28237);
and U31820 (N_31820,N_28077,N_29236);
and U31821 (N_31821,N_29345,N_28568);
xor U31822 (N_31822,N_28371,N_29226);
xor U31823 (N_31823,N_29686,N_28233);
nor U31824 (N_31824,N_28421,N_29341);
and U31825 (N_31825,N_28620,N_28624);
nand U31826 (N_31826,N_29358,N_28111);
nand U31827 (N_31827,N_28070,N_29677);
and U31828 (N_31828,N_28462,N_29045);
xnor U31829 (N_31829,N_29493,N_29473);
nand U31830 (N_31830,N_28989,N_28741);
nor U31831 (N_31831,N_29117,N_28791);
or U31832 (N_31832,N_28798,N_29620);
xor U31833 (N_31833,N_29621,N_28880);
nor U31834 (N_31834,N_29357,N_29172);
and U31835 (N_31835,N_29277,N_29570);
and U31836 (N_31836,N_29775,N_28415);
nand U31837 (N_31837,N_28274,N_29140);
nand U31838 (N_31838,N_29019,N_29275);
and U31839 (N_31839,N_28232,N_29933);
xor U31840 (N_31840,N_29940,N_29752);
nand U31841 (N_31841,N_29553,N_29556);
nand U31842 (N_31842,N_29465,N_28358);
nor U31843 (N_31843,N_29744,N_28048);
and U31844 (N_31844,N_28368,N_28135);
xor U31845 (N_31845,N_29282,N_29090);
xnor U31846 (N_31846,N_29365,N_28913);
and U31847 (N_31847,N_29289,N_28410);
xnor U31848 (N_31848,N_29527,N_28947);
nand U31849 (N_31849,N_28294,N_28024);
nand U31850 (N_31850,N_28632,N_28119);
or U31851 (N_31851,N_28188,N_29825);
and U31852 (N_31852,N_29855,N_28373);
or U31853 (N_31853,N_28055,N_28427);
nor U31854 (N_31854,N_28489,N_29241);
nand U31855 (N_31855,N_28745,N_29373);
and U31856 (N_31856,N_29787,N_29479);
xor U31857 (N_31857,N_29441,N_29218);
nor U31858 (N_31858,N_28570,N_29067);
nand U31859 (N_31859,N_29828,N_28085);
nand U31860 (N_31860,N_28789,N_28935);
and U31861 (N_31861,N_28931,N_28250);
xor U31862 (N_31862,N_29936,N_29368);
nor U31863 (N_31863,N_29706,N_29758);
nand U31864 (N_31864,N_29405,N_29784);
xor U31865 (N_31865,N_28308,N_29564);
nand U31866 (N_31866,N_29070,N_29016);
and U31867 (N_31867,N_28708,N_29751);
nor U31868 (N_31868,N_28239,N_28815);
nor U31869 (N_31869,N_28704,N_29784);
nor U31870 (N_31870,N_28947,N_29814);
or U31871 (N_31871,N_28263,N_29602);
nor U31872 (N_31872,N_29135,N_28364);
xor U31873 (N_31873,N_28013,N_29030);
xnor U31874 (N_31874,N_28611,N_29422);
and U31875 (N_31875,N_29260,N_29634);
nor U31876 (N_31876,N_28804,N_28292);
nand U31877 (N_31877,N_28663,N_29080);
and U31878 (N_31878,N_29400,N_29589);
xnor U31879 (N_31879,N_28678,N_29760);
or U31880 (N_31880,N_28938,N_28648);
nor U31881 (N_31881,N_28360,N_28749);
or U31882 (N_31882,N_28993,N_29539);
and U31883 (N_31883,N_28956,N_28928);
nand U31884 (N_31884,N_28807,N_29384);
nor U31885 (N_31885,N_28662,N_29873);
nor U31886 (N_31886,N_29650,N_29335);
xnor U31887 (N_31887,N_29471,N_29026);
and U31888 (N_31888,N_28489,N_28328);
nor U31889 (N_31889,N_28043,N_29141);
nand U31890 (N_31890,N_29929,N_28893);
xor U31891 (N_31891,N_29149,N_28002);
xnor U31892 (N_31892,N_28725,N_29572);
xnor U31893 (N_31893,N_28075,N_29404);
nor U31894 (N_31894,N_28990,N_29036);
and U31895 (N_31895,N_29710,N_28545);
xnor U31896 (N_31896,N_29090,N_29162);
and U31897 (N_31897,N_28346,N_28991);
or U31898 (N_31898,N_28445,N_28810);
nor U31899 (N_31899,N_28215,N_28604);
and U31900 (N_31900,N_29499,N_28899);
or U31901 (N_31901,N_29253,N_29254);
nand U31902 (N_31902,N_28564,N_28119);
nor U31903 (N_31903,N_28804,N_29902);
xnor U31904 (N_31904,N_29835,N_29031);
and U31905 (N_31905,N_29728,N_29639);
nor U31906 (N_31906,N_29840,N_28945);
xnor U31907 (N_31907,N_29916,N_28974);
nand U31908 (N_31908,N_28239,N_29876);
xnor U31909 (N_31909,N_29692,N_28146);
xnor U31910 (N_31910,N_29773,N_28526);
xor U31911 (N_31911,N_28657,N_29687);
nor U31912 (N_31912,N_28129,N_29013);
nand U31913 (N_31913,N_29278,N_29853);
and U31914 (N_31914,N_28246,N_28206);
and U31915 (N_31915,N_28865,N_29114);
or U31916 (N_31916,N_29160,N_28358);
nor U31917 (N_31917,N_28438,N_29831);
nor U31918 (N_31918,N_28010,N_29537);
nor U31919 (N_31919,N_29390,N_28143);
nand U31920 (N_31920,N_28746,N_29847);
nor U31921 (N_31921,N_29574,N_29711);
nor U31922 (N_31922,N_29914,N_29466);
nor U31923 (N_31923,N_28337,N_29294);
and U31924 (N_31924,N_29972,N_29415);
and U31925 (N_31925,N_28516,N_29794);
and U31926 (N_31926,N_29656,N_28430);
nor U31927 (N_31927,N_29767,N_29425);
or U31928 (N_31928,N_28462,N_29863);
nor U31929 (N_31929,N_29054,N_29456);
nor U31930 (N_31930,N_28823,N_28279);
xnor U31931 (N_31931,N_28681,N_28484);
and U31932 (N_31932,N_28884,N_29400);
or U31933 (N_31933,N_29850,N_28188);
or U31934 (N_31934,N_29746,N_28331);
xor U31935 (N_31935,N_28835,N_29492);
and U31936 (N_31936,N_29879,N_29686);
nor U31937 (N_31937,N_29087,N_28848);
or U31938 (N_31938,N_28242,N_29266);
nor U31939 (N_31939,N_29100,N_29760);
nor U31940 (N_31940,N_28049,N_28675);
nor U31941 (N_31941,N_28573,N_29971);
nor U31942 (N_31942,N_28684,N_29335);
and U31943 (N_31943,N_28855,N_28180);
xor U31944 (N_31944,N_29586,N_29114);
xnor U31945 (N_31945,N_28397,N_28105);
or U31946 (N_31946,N_28544,N_28942);
or U31947 (N_31947,N_29426,N_28840);
or U31948 (N_31948,N_28094,N_29239);
and U31949 (N_31949,N_29991,N_28829);
or U31950 (N_31950,N_28075,N_29519);
nand U31951 (N_31951,N_29092,N_29209);
xor U31952 (N_31952,N_29540,N_28273);
and U31953 (N_31953,N_28779,N_28407);
or U31954 (N_31954,N_28511,N_28422);
nand U31955 (N_31955,N_28572,N_29313);
nand U31956 (N_31956,N_28303,N_29514);
nand U31957 (N_31957,N_29106,N_29811);
xor U31958 (N_31958,N_28993,N_28897);
and U31959 (N_31959,N_28774,N_29601);
xor U31960 (N_31960,N_28509,N_28412);
nand U31961 (N_31961,N_28921,N_28977);
or U31962 (N_31962,N_29314,N_29987);
nor U31963 (N_31963,N_29479,N_29952);
nor U31964 (N_31964,N_29480,N_28871);
nand U31965 (N_31965,N_28745,N_29311);
or U31966 (N_31966,N_28940,N_28250);
or U31967 (N_31967,N_28448,N_28060);
nor U31968 (N_31968,N_28675,N_28583);
nor U31969 (N_31969,N_29636,N_28067);
or U31970 (N_31970,N_28884,N_28348);
nand U31971 (N_31971,N_29260,N_28825);
nand U31972 (N_31972,N_29103,N_28643);
and U31973 (N_31973,N_29932,N_28428);
nor U31974 (N_31974,N_28045,N_28517);
nand U31975 (N_31975,N_29778,N_29753);
xor U31976 (N_31976,N_28795,N_29047);
xnor U31977 (N_31977,N_28568,N_29897);
and U31978 (N_31978,N_28581,N_29683);
and U31979 (N_31979,N_28732,N_28061);
nand U31980 (N_31980,N_28548,N_28491);
xnor U31981 (N_31981,N_29658,N_29299);
nor U31982 (N_31982,N_28052,N_29429);
or U31983 (N_31983,N_28387,N_29677);
or U31984 (N_31984,N_29160,N_29589);
nor U31985 (N_31985,N_29121,N_29208);
xnor U31986 (N_31986,N_28927,N_29406);
and U31987 (N_31987,N_29482,N_28729);
and U31988 (N_31988,N_29212,N_28052);
nor U31989 (N_31989,N_29568,N_28947);
and U31990 (N_31990,N_28848,N_29097);
nand U31991 (N_31991,N_29232,N_28125);
or U31992 (N_31992,N_28701,N_29575);
nand U31993 (N_31993,N_29433,N_29840);
nand U31994 (N_31994,N_28362,N_28554);
and U31995 (N_31995,N_29623,N_29347);
nor U31996 (N_31996,N_29565,N_29927);
or U31997 (N_31997,N_29556,N_29818);
or U31998 (N_31998,N_29859,N_29330);
or U31999 (N_31999,N_28600,N_29591);
and U32000 (N_32000,N_30633,N_31454);
xnor U32001 (N_32001,N_31946,N_30869);
and U32002 (N_32002,N_31987,N_30252);
xor U32003 (N_32003,N_30729,N_31111);
xnor U32004 (N_32004,N_30058,N_31093);
xnor U32005 (N_32005,N_30565,N_31033);
or U32006 (N_32006,N_30557,N_30552);
nor U32007 (N_32007,N_31301,N_30338);
nand U32008 (N_32008,N_31576,N_30891);
xnor U32009 (N_32009,N_31335,N_31386);
and U32010 (N_32010,N_31757,N_30900);
nand U32011 (N_32011,N_31603,N_31799);
nand U32012 (N_32012,N_30010,N_31903);
and U32013 (N_32013,N_30423,N_31518);
and U32014 (N_32014,N_31483,N_30330);
and U32015 (N_32015,N_30677,N_30518);
and U32016 (N_32016,N_30568,N_31068);
or U32017 (N_32017,N_31362,N_30420);
xor U32018 (N_32018,N_31546,N_30984);
nor U32019 (N_32019,N_30882,N_30656);
or U32020 (N_32020,N_30837,N_30777);
xnor U32021 (N_32021,N_31031,N_31183);
or U32022 (N_32022,N_31368,N_30881);
or U32023 (N_32023,N_31293,N_31707);
or U32024 (N_32024,N_30359,N_31389);
or U32025 (N_32025,N_30855,N_31783);
and U32026 (N_32026,N_31678,N_31871);
or U32027 (N_32027,N_31222,N_30017);
nor U32028 (N_32028,N_31807,N_31319);
nand U32029 (N_32029,N_30817,N_30657);
and U32030 (N_32030,N_31512,N_31457);
and U32031 (N_32031,N_30844,N_31276);
and U32032 (N_32032,N_30524,N_30339);
xor U32033 (N_32033,N_30705,N_30475);
xor U32034 (N_32034,N_30481,N_30024);
xor U32035 (N_32035,N_30030,N_30344);
nor U32036 (N_32036,N_30413,N_31689);
xnor U32037 (N_32037,N_30977,N_31211);
or U32038 (N_32038,N_30585,N_30722);
nand U32039 (N_32039,N_31806,N_30347);
or U32040 (N_32040,N_30778,N_30887);
and U32041 (N_32041,N_31417,N_31739);
nor U32042 (N_32042,N_31458,N_31261);
or U32043 (N_32043,N_31930,N_31556);
or U32044 (N_32044,N_30685,N_30211);
or U32045 (N_32045,N_31326,N_30516);
or U32046 (N_32046,N_30104,N_31575);
and U32047 (N_32047,N_30045,N_31342);
and U32048 (N_32048,N_30453,N_31565);
nand U32049 (N_32049,N_31046,N_31455);
and U32050 (N_32050,N_31882,N_30428);
nor U32051 (N_32051,N_31038,N_30749);
and U32052 (N_32052,N_31025,N_31352);
nor U32053 (N_32053,N_30609,N_30617);
xnor U32054 (N_32054,N_31192,N_31844);
xor U32055 (N_32055,N_30174,N_30526);
or U32056 (N_32056,N_30071,N_30971);
xor U32057 (N_32057,N_30590,N_30397);
nor U32058 (N_32058,N_31957,N_31879);
nor U32059 (N_32059,N_31670,N_31595);
nor U32060 (N_32060,N_31652,N_31085);
nand U32061 (N_32061,N_30287,N_31440);
nor U32062 (N_32062,N_30631,N_30219);
nor U32063 (N_32063,N_30506,N_30515);
nand U32064 (N_32064,N_31185,N_31938);
nor U32065 (N_32065,N_30035,N_30079);
nand U32066 (N_32066,N_31850,N_31558);
nor U32067 (N_32067,N_31126,N_30802);
nand U32068 (N_32068,N_30788,N_30871);
and U32069 (N_32069,N_30438,N_30675);
xor U32070 (N_32070,N_30694,N_31557);
nand U32071 (N_32071,N_30070,N_31538);
or U32072 (N_32072,N_31376,N_31515);
or U32073 (N_32073,N_30640,N_30502);
and U32074 (N_32074,N_31607,N_30576);
and U32075 (N_32075,N_31079,N_31717);
xnor U32076 (N_32076,N_31840,N_30091);
nor U32077 (N_32077,N_30872,N_30066);
or U32078 (N_32078,N_31856,N_31400);
and U32079 (N_32079,N_30425,N_31446);
or U32080 (N_32080,N_30402,N_30271);
nand U32081 (N_32081,N_31028,N_30944);
xor U32082 (N_32082,N_31304,N_31955);
nand U32083 (N_32083,N_30849,N_30263);
nor U32084 (N_32084,N_31470,N_31241);
or U32085 (N_32085,N_30150,N_30100);
nand U32086 (N_32086,N_30937,N_31469);
or U32087 (N_32087,N_31519,N_31263);
nand U32088 (N_32088,N_31026,N_31941);
and U32089 (N_32089,N_30845,N_30843);
or U32090 (N_32090,N_30600,N_31287);
and U32091 (N_32091,N_30779,N_30105);
xor U32092 (N_32092,N_30061,N_30088);
xnor U32093 (N_32093,N_31696,N_30093);
or U32094 (N_32094,N_30445,N_30447);
or U32095 (N_32095,N_30701,N_31655);
nand U32096 (N_32096,N_30716,N_30063);
xnor U32097 (N_32097,N_30369,N_30690);
nand U32098 (N_32098,N_30895,N_30492);
and U32099 (N_32099,N_30798,N_30121);
nor U32100 (N_32100,N_30567,N_30990);
nor U32101 (N_32101,N_30296,N_30825);
xnor U32102 (N_32102,N_31822,N_31665);
or U32103 (N_32103,N_30302,N_31220);
or U32104 (N_32104,N_30038,N_31718);
or U32105 (N_32105,N_30201,N_30771);
and U32106 (N_32106,N_30493,N_31180);
or U32107 (N_32107,N_31012,N_31249);
nor U32108 (N_32108,N_30514,N_30251);
nand U32109 (N_32109,N_30813,N_31204);
nand U32110 (N_32110,N_30435,N_31269);
and U32111 (N_32111,N_31825,N_31378);
xor U32112 (N_32112,N_31484,N_31507);
xnor U32113 (N_32113,N_30185,N_31349);
and U32114 (N_32114,N_31305,N_30549);
or U32115 (N_32115,N_30233,N_30225);
nor U32116 (N_32116,N_31870,N_30662);
or U32117 (N_32117,N_30665,N_30486);
or U32118 (N_32118,N_30786,N_30508);
and U32119 (N_32119,N_31845,N_30537);
and U32120 (N_32120,N_30653,N_30196);
or U32121 (N_32121,N_30950,N_31165);
nor U32122 (N_32122,N_30765,N_30520);
nand U32123 (N_32123,N_30449,N_30528);
nand U32124 (N_32124,N_30725,N_30897);
xor U32125 (N_32125,N_30189,N_31096);
and U32126 (N_32126,N_31555,N_30801);
nand U32127 (N_32127,N_30917,N_31169);
xor U32128 (N_32128,N_30069,N_30929);
nand U32129 (N_32129,N_30266,N_31090);
nand U32130 (N_32130,N_30822,N_30766);
nand U32131 (N_32131,N_30365,N_31059);
and U32132 (N_32132,N_30842,N_30139);
or U32133 (N_32133,N_31226,N_31816);
or U32134 (N_32134,N_30324,N_31864);
or U32135 (N_32135,N_31354,N_30868);
nand U32136 (N_32136,N_31920,N_30510);
xnor U32137 (N_32137,N_30215,N_30074);
xor U32138 (N_32138,N_30734,N_30394);
nor U32139 (N_32139,N_31874,N_30578);
nand U32140 (N_32140,N_30461,N_31766);
and U32141 (N_32141,N_30889,N_31243);
nand U32142 (N_32142,N_30229,N_31159);
xor U32143 (N_32143,N_31426,N_30404);
or U32144 (N_32144,N_31923,N_30446);
nor U32145 (N_32145,N_31753,N_31817);
nor U32146 (N_32146,N_31937,N_30561);
nand U32147 (N_32147,N_30239,N_30744);
and U32148 (N_32148,N_31441,N_31235);
or U32149 (N_32149,N_31466,N_31520);
or U32150 (N_32150,N_31917,N_31632);
and U32151 (N_32151,N_30148,N_30129);
nor U32152 (N_32152,N_30180,N_31307);
and U32153 (N_32153,N_30130,N_30337);
xor U32154 (N_32154,N_30328,N_31421);
or U32155 (N_32155,N_30770,N_31979);
nor U32156 (N_32156,N_31708,N_31171);
xnor U32157 (N_32157,N_30754,N_31786);
or U32158 (N_32158,N_31756,N_30336);
or U32159 (N_32159,N_31745,N_31819);
and U32160 (N_32160,N_31161,N_30213);
xnor U32161 (N_32161,N_30621,N_30382);
or U32162 (N_32162,N_30538,N_31212);
nand U32163 (N_32163,N_30313,N_31580);
nand U32164 (N_32164,N_30919,N_31311);
or U32165 (N_32165,N_31742,N_30673);
nand U32166 (N_32166,N_30742,N_30852);
nand U32167 (N_32167,N_31741,N_30769);
or U32168 (N_32168,N_30969,N_30946);
nand U32169 (N_32169,N_30441,N_30395);
nand U32170 (N_32170,N_31091,N_31526);
nor U32171 (N_32171,N_31474,N_31729);
and U32172 (N_32172,N_31824,N_31925);
and U32173 (N_32173,N_31495,N_30584);
or U32174 (N_32174,N_30949,N_30197);
or U32175 (N_32175,N_30941,N_30278);
or U32176 (N_32176,N_31251,N_31506);
nand U32177 (N_32177,N_30939,N_31338);
nor U32178 (N_32178,N_30473,N_31110);
and U32179 (N_32179,N_31744,N_30275);
or U32180 (N_32180,N_31069,N_30570);
or U32181 (N_32181,N_31115,N_31189);
or U32182 (N_32182,N_31160,N_31728);
or U32183 (N_32183,N_30859,N_31736);
and U32184 (N_32184,N_31430,N_31238);
nand U32185 (N_32185,N_31590,N_30226);
xor U32186 (N_32186,N_30907,N_30081);
or U32187 (N_32187,N_31501,N_31361);
or U32188 (N_32188,N_30361,N_31477);
or U32189 (N_32189,N_31401,N_31582);
xor U32190 (N_32190,N_30295,N_30522);
xnor U32191 (N_32191,N_30857,N_31567);
xnor U32192 (N_32192,N_30536,N_30638);
and U32193 (N_32193,N_30607,N_30102);
nor U32194 (N_32194,N_30647,N_30400);
xor U32195 (N_32195,N_30043,N_30052);
and U32196 (N_32196,N_30767,N_31107);
and U32197 (N_32197,N_31749,N_30434);
or U32198 (N_32198,N_31774,N_30998);
xor U32199 (N_32199,N_30676,N_30507);
and U32200 (N_32200,N_30965,N_31909);
and U32201 (N_32201,N_30957,N_31253);
or U32202 (N_32202,N_31569,N_30469);
xor U32203 (N_32203,N_30978,N_31347);
nand U32204 (N_32204,N_31480,N_30267);
and U32205 (N_32205,N_31605,N_30118);
and U32206 (N_32206,N_30926,N_30599);
xor U32207 (N_32207,N_30542,N_30529);
nor U32208 (N_32208,N_30468,N_31881);
nor U32209 (N_32209,N_30630,N_31945);
nor U32210 (N_32210,N_30214,N_31570);
nand U32211 (N_32211,N_30839,N_31773);
nor U32212 (N_32212,N_31700,N_30559);
nor U32213 (N_32213,N_31579,N_31043);
and U32214 (N_32214,N_31382,N_31995);
nor U32215 (N_32215,N_31018,N_31967);
nand U32216 (N_32216,N_31725,N_31921);
nand U32217 (N_32217,N_31999,N_31895);
nand U32218 (N_32218,N_31589,N_30471);
and U32219 (N_32219,N_31510,N_31529);
and U32220 (N_32220,N_30112,N_30745);
xnor U32221 (N_32221,N_30873,N_30586);
nand U32222 (N_32222,N_30426,N_31723);
nor U32223 (N_32223,N_30042,N_30184);
xnor U32224 (N_32224,N_31360,N_31146);
and U32225 (N_32225,N_30994,N_30146);
nand U32226 (N_32226,N_31981,N_30027);
and U32227 (N_32227,N_30790,N_30711);
or U32228 (N_32228,N_30979,N_31996);
nand U32229 (N_32229,N_30188,N_30316);
nor U32230 (N_32230,N_30132,N_30735);
or U32231 (N_32231,N_30671,N_30216);
xor U32232 (N_32232,N_30606,N_31587);
nand U32233 (N_32233,N_31064,N_30668);
or U32234 (N_32234,N_30244,N_30807);
and U32235 (N_32235,N_31794,N_31523);
xnor U32236 (N_32236,N_31420,N_31244);
and U32237 (N_32237,N_31542,N_30659);
nand U32238 (N_32238,N_30200,N_31563);
nor U32239 (N_32239,N_31394,N_30173);
and U32240 (N_32240,N_31657,N_31493);
and U32241 (N_32241,N_30564,N_30596);
or U32242 (N_32242,N_31887,N_30810);
or U32243 (N_32243,N_30488,N_31913);
xor U32244 (N_32244,N_31922,N_30370);
or U32245 (N_32245,N_30149,N_30667);
xor U32246 (N_32246,N_31828,N_30288);
and U32247 (N_32247,N_30966,N_31131);
and U32248 (N_32248,N_31298,N_30476);
nand U32249 (N_32249,N_31438,N_30953);
xor U32250 (N_32250,N_31366,N_31422);
and U32251 (N_32251,N_30658,N_30163);
nor U32252 (N_32252,N_30901,N_31734);
or U32253 (N_32253,N_30731,N_31133);
xnor U32254 (N_32254,N_31318,N_31695);
and U32255 (N_32255,N_31040,N_31528);
or U32256 (N_32256,N_31504,N_31129);
or U32257 (N_32257,N_31768,N_31897);
nand U32258 (N_32258,N_30545,N_30142);
nand U32259 (N_32259,N_30265,N_31927);
and U32260 (N_32260,N_30899,N_31746);
xor U32261 (N_32261,N_31596,N_30389);
and U32262 (N_32262,N_31434,N_30032);
nand U32263 (N_32263,N_30120,N_31296);
xor U32264 (N_32264,N_31142,N_31388);
nor U32265 (N_32265,N_31199,N_31503);
and U32266 (N_32266,N_31780,N_31508);
nor U32267 (N_32267,N_31083,N_31187);
and U32268 (N_32268,N_31312,N_31705);
nand U32269 (N_32269,N_31853,N_31796);
xor U32270 (N_32270,N_30925,N_31641);
nor U32271 (N_32271,N_30311,N_31174);
xnor U32272 (N_32272,N_30304,N_31292);
xnor U32273 (N_32273,N_31379,N_31445);
nand U32274 (N_32274,N_31343,N_31163);
or U32275 (N_32275,N_31924,N_30191);
and U32276 (N_32276,N_30885,N_30695);
and U32277 (N_32277,N_30409,N_31597);
xnor U32278 (N_32278,N_30748,N_31384);
xor U32279 (N_32279,N_30095,N_31811);
or U32280 (N_32280,N_30367,N_31099);
nor U32281 (N_32281,N_30172,N_31081);
nand U32282 (N_32282,N_31057,N_30624);
and U32283 (N_32283,N_31065,N_31140);
and U32284 (N_32284,N_31553,N_31153);
and U32285 (N_32285,N_30222,N_30718);
or U32286 (N_32286,N_31554,N_31274);
nor U32287 (N_32287,N_31016,N_31055);
or U32288 (N_32288,N_31186,N_30107);
or U32289 (N_32289,N_31341,N_31517);
nand U32290 (N_32290,N_30963,N_30416);
and U32291 (N_32291,N_30799,N_31502);
and U32292 (N_32292,N_31683,N_31615);
or U32293 (N_32293,N_30012,N_30574);
and U32294 (N_32294,N_30905,N_31252);
or U32295 (N_32295,N_30377,N_30831);
and U32296 (N_32296,N_30715,N_31315);
and U32297 (N_32297,N_30047,N_31968);
or U32298 (N_32298,N_31693,N_31948);
nor U32299 (N_32299,N_31203,N_31877);
xnor U32300 (N_32300,N_30106,N_30013);
nor U32301 (N_32301,N_30571,N_31884);
nor U32302 (N_32302,N_31541,N_30232);
nand U32303 (N_32303,N_30732,N_31795);
nand U32304 (N_32304,N_30562,N_31835);
nor U32305 (N_32305,N_31574,N_30041);
and U32306 (N_32306,N_31381,N_30448);
and U32307 (N_32307,N_30719,N_30613);
and U32308 (N_32308,N_30127,N_30487);
or U32309 (N_32309,N_30223,N_30593);
and U32310 (N_32310,N_31865,N_31713);
or U32311 (N_32311,N_31490,N_31722);
nor U32312 (N_32312,N_31758,N_31290);
nand U32313 (N_32313,N_31704,N_30764);
xor U32314 (N_32314,N_30997,N_30342);
nor U32315 (N_32315,N_31721,N_31888);
xor U32316 (N_32316,N_30955,N_31348);
or U32317 (N_32317,N_30605,N_30366);
xor U32318 (N_32318,N_31667,N_30273);
and U32319 (N_32319,N_30444,N_31339);
xor U32320 (N_32320,N_30323,N_31694);
nor U32321 (N_32321,N_31218,N_30752);
nor U32322 (N_32322,N_30406,N_31775);
xor U32323 (N_32323,N_30970,N_30616);
and U32324 (N_32324,N_30846,N_30283);
or U32325 (N_32325,N_31077,N_31798);
and U32326 (N_32326,N_30076,N_30332);
xnor U32327 (N_32327,N_31755,N_30085);
xnor U32328 (N_32328,N_31984,N_30833);
and U32329 (N_32329,N_31284,N_30649);
xor U32330 (N_32330,N_31566,N_30281);
xnor U32331 (N_32331,N_31697,N_30411);
nor U32332 (N_32332,N_31479,N_31215);
or U32333 (N_32333,N_30847,N_30721);
and U32334 (N_32334,N_31698,N_31939);
nand U32335 (N_32335,N_30577,N_30591);
nand U32336 (N_32336,N_30811,N_31061);
and U32337 (N_32337,N_30218,N_30333);
nand U32338 (N_32338,N_31393,N_31513);
nor U32339 (N_32339,N_31801,N_31971);
xnor U32340 (N_32340,N_31087,N_30485);
nand U32341 (N_32341,N_30405,N_31647);
and U32342 (N_32342,N_31210,N_31793);
or U32343 (N_32343,N_30916,N_30064);
and U32344 (N_32344,N_31256,N_31473);
and U32345 (N_32345,N_31158,N_30666);
or U32346 (N_32346,N_30964,N_31195);
nand U32347 (N_32347,N_30360,N_30987);
nor U32348 (N_32348,N_30375,N_30451);
nand U32349 (N_32349,N_30740,N_31358);
xnor U32350 (N_32350,N_31482,N_31308);
nand U32351 (N_32351,N_31359,N_30224);
or U32352 (N_32352,N_31150,N_31245);
xor U32353 (N_32353,N_30096,N_30153);
nor U32354 (N_32354,N_30472,N_30959);
nand U32355 (N_32355,N_30911,N_31001);
xor U32356 (N_32356,N_30164,N_31719);
nand U32357 (N_32357,N_30034,N_30741);
and U32358 (N_32358,N_30384,N_30220);
nor U32359 (N_32359,N_30388,N_30611);
nor U32360 (N_32360,N_30908,N_30724);
and U32361 (N_32361,N_31970,N_31521);
or U32362 (N_32362,N_31273,N_31547);
nand U32363 (N_32363,N_31154,N_31906);
or U32364 (N_32364,N_31965,N_31804);
and U32365 (N_32365,N_30175,N_31701);
xnor U32366 (N_32366,N_30457,N_31390);
nand U32367 (N_32367,N_30372,N_30761);
xor U32368 (N_32368,N_31021,N_30829);
or U32369 (N_32369,N_30083,N_31205);
and U32370 (N_32370,N_30254,N_30029);
nor U32371 (N_32371,N_31892,N_30592);
or U32372 (N_32372,N_30828,N_30354);
nand U32373 (N_32373,N_31522,N_31787);
and U32374 (N_32374,N_31498,N_31336);
nor U32375 (N_32375,N_30004,N_31385);
nand U32376 (N_32376,N_30422,N_30714);
xor U32377 (N_32377,N_31066,N_31200);
nor U32378 (N_32378,N_31280,N_30948);
or U32379 (N_32379,N_31139,N_31428);
and U32380 (N_32380,N_30892,N_31095);
or U32381 (N_32381,N_30835,N_30168);
or U32382 (N_32382,N_31690,N_30092);
nand U32383 (N_32383,N_31823,N_31000);
nor U32384 (N_32384,N_31890,N_31666);
and U32385 (N_32385,N_30904,N_30708);
nor U32386 (N_32386,N_31112,N_31092);
nor U32387 (N_32387,N_30221,N_31990);
and U32388 (N_32388,N_30020,N_30321);
or U32389 (N_32389,N_31188,N_31042);
xnor U32390 (N_32390,N_30235,N_30679);
xnor U32391 (N_32391,N_31184,N_31899);
nor U32392 (N_32392,N_30040,N_30875);
or U32393 (N_32393,N_31275,N_30080);
and U32394 (N_32394,N_30503,N_30597);
xnor U32395 (N_32395,N_31983,N_30031);
nor U32396 (N_32396,N_31489,N_30635);
and U32397 (N_32397,N_30099,N_30755);
nand U32398 (N_32398,N_31748,N_31964);
xnor U32399 (N_32399,N_31620,N_30583);
and U32400 (N_32400,N_31716,N_30260);
nand U32401 (N_32401,N_31377,N_31524);
xor U32402 (N_32402,N_31496,N_31475);
and U32403 (N_32403,N_30883,N_31432);
and U32404 (N_32404,N_31356,N_31859);
xnor U32405 (N_32405,N_31190,N_30644);
xnor U32406 (N_32406,N_31076,N_30182);
nand U32407 (N_32407,N_30856,N_30867);
nor U32408 (N_32408,N_31279,N_30812);
nand U32409 (N_32409,N_31265,N_30303);
nand U32410 (N_32410,N_31436,N_31991);
nor U32411 (N_32411,N_31340,N_30186);
xor U32412 (N_32412,N_30595,N_30016);
nand U32413 (N_32413,N_31317,N_31444);
or U32414 (N_32414,N_30037,N_31125);
nor U32415 (N_32415,N_31872,N_31600);
nand U32416 (N_32416,N_30376,N_31468);
nor U32417 (N_32417,N_30049,N_30103);
or U32418 (N_32418,N_31592,N_31942);
nand U32419 (N_32419,N_31050,N_30525);
and U32420 (N_32420,N_30785,N_31223);
and U32421 (N_32421,N_30230,N_30019);
or U32422 (N_32422,N_30128,N_31141);
nand U32423 (N_32423,N_31998,N_30758);
nand U32424 (N_32424,N_31571,N_30726);
nand U32425 (N_32425,N_30407,N_31300);
nor U32426 (N_32426,N_31910,N_31883);
nor U32427 (N_32427,N_31754,N_31041);
nor U32428 (N_32428,N_31487,N_31313);
xor U32429 (N_32429,N_30757,N_31494);
nor U32430 (N_32430,N_30880,N_31119);
or U32431 (N_32431,N_31413,N_30495);
and U32432 (N_32432,N_31649,N_30642);
nand U32433 (N_32433,N_30259,N_31854);
or U32434 (N_32434,N_31264,N_30650);
xor U32435 (N_32435,N_30157,N_31671);
or U32436 (N_32436,N_31969,N_30738);
or U32437 (N_32437,N_31973,N_31425);
or U32438 (N_32438,N_30165,N_31030);
xor U32439 (N_32439,N_31404,N_30888);
nand U32440 (N_32440,N_30484,N_30727);
or U32441 (N_32441,N_30961,N_31837);
or U32442 (N_32442,N_30933,N_30340);
nand U32443 (N_32443,N_30893,N_31443);
xnor U32444 (N_32444,N_31650,N_30101);
nor U32445 (N_32445,N_30439,N_30300);
and U32446 (N_32446,N_31581,N_31509);
or U32447 (N_32447,N_30906,N_30463);
nand U32448 (N_32448,N_30116,N_30532);
and U32449 (N_32449,N_30312,N_30289);
and U32450 (N_32450,N_31201,N_30379);
or U32451 (N_32451,N_31688,N_31550);
xnor U32452 (N_32452,N_31735,N_31833);
nor U32453 (N_32453,N_31992,N_30308);
xor U32454 (N_32454,N_31669,N_31216);
and U32455 (N_32455,N_30923,N_31789);
nor U32456 (N_32456,N_31486,N_31886);
nor U32457 (N_32457,N_31894,N_30494);
and U32458 (N_32458,N_30654,N_30498);
xnor U32459 (N_32459,N_31790,N_30381);
nand U32460 (N_32460,N_30417,N_31637);
and U32461 (N_32461,N_30298,N_30131);
nor U32462 (N_32462,N_30364,N_31548);
nand U32463 (N_32463,N_30410,N_30158);
xor U32464 (N_32464,N_31258,N_31060);
nor U32465 (N_32465,N_31453,N_30141);
and U32466 (N_32466,N_31023,N_31399);
or U32467 (N_32467,N_31624,N_30231);
nor U32468 (N_32468,N_31838,N_30238);
nand U32469 (N_32469,N_31534,N_31989);
xor U32470 (N_32470,N_30903,N_31949);
and U32471 (N_32471,N_31374,N_30432);
nand U32472 (N_32472,N_31875,N_30176);
or U32473 (N_32473,N_30992,N_31157);
or U32474 (N_32474,N_31631,N_31958);
or U32475 (N_32475,N_30806,N_30815);
and U32476 (N_32476,N_30315,N_31283);
and U32477 (N_32477,N_31411,N_30850);
xor U32478 (N_32478,N_30001,N_31063);
nand U32479 (N_32479,N_31488,N_30205);
nand U32480 (N_32480,N_31034,N_31588);
and U32481 (N_32481,N_30934,N_31709);
and U32482 (N_32482,N_30046,N_31640);
nand U32483 (N_32483,N_30009,N_30082);
or U32484 (N_32484,N_31659,N_30913);
or U32485 (N_32485,N_31772,N_30466);
or U32486 (N_32486,N_31395,N_31463);
or U32487 (N_32487,N_30918,N_30002);
nor U32488 (N_32488,N_30117,N_31306);
nor U32489 (N_32489,N_30632,N_31013);
nor U32490 (N_32490,N_30023,N_30479);
xor U32491 (N_32491,N_31198,N_30318);
nor U32492 (N_32492,N_30629,N_31584);
or U32493 (N_32493,N_31345,N_30145);
nand U32494 (N_32494,N_30044,N_30418);
xor U32495 (N_32495,N_31953,N_31599);
nand U32496 (N_32496,N_30728,N_30212);
nand U32497 (N_32497,N_31224,N_31685);
nor U32498 (N_32498,N_31834,N_30258);
nand U32499 (N_32499,N_31767,N_31295);
or U32500 (N_32500,N_31978,N_30928);
nand U32501 (N_32501,N_31233,N_30138);
or U32502 (N_32502,N_30309,N_30774);
or U32503 (N_32503,N_31726,N_31122);
and U32504 (N_32504,N_31086,N_31197);
and U32505 (N_32505,N_31610,N_31442);
xor U32506 (N_32506,N_30820,N_30670);
nand U32507 (N_32507,N_31648,N_31710);
nor U32508 (N_32508,N_30826,N_30137);
or U32509 (N_32509,N_30858,N_31578);
nor U32510 (N_32510,N_30912,N_31437);
nor U32511 (N_32511,N_30199,N_30166);
xor U32512 (N_32512,N_31858,N_30217);
nor U32513 (N_32513,N_30573,N_30527);
nand U32514 (N_32514,N_30115,N_30282);
xnor U32515 (N_32515,N_31147,N_31118);
nand U32516 (N_32516,N_31074,N_31947);
nor U32517 (N_32517,N_30830,N_30329);
nand U32518 (N_32518,N_30553,N_31408);
nor U32519 (N_32519,N_31977,N_30558);
xnor U32520 (N_32520,N_31672,N_30795);
and U32521 (N_32521,N_31478,N_31105);
and U32522 (N_32522,N_31075,N_30608);
xor U32523 (N_32523,N_31321,N_31471);
xnor U32524 (N_32524,N_31976,N_31836);
and U32525 (N_32525,N_30739,N_30203);
nand U32526 (N_32526,N_31070,N_30713);
and U32527 (N_32527,N_31214,N_31114);
and U32528 (N_32528,N_30179,N_31645);
nor U32529 (N_32529,N_30028,N_30119);
xor U32530 (N_32530,N_30976,N_30824);
nand U32531 (N_32531,N_31530,N_30094);
or U32532 (N_32532,N_31743,N_30930);
nand U32533 (N_32533,N_30022,N_30078);
nand U32534 (N_32534,N_31476,N_30261);
nand U32535 (N_32535,N_31863,N_31175);
or U32536 (N_32536,N_31164,N_31491);
and U32537 (N_32537,N_31418,N_31402);
and U32538 (N_32538,N_30202,N_31658);
nand U32539 (N_32539,N_31961,N_31309);
nand U32540 (N_32540,N_31009,N_30555);
nand U32541 (N_32541,N_31779,N_30927);
nor U32542 (N_32542,N_31573,N_31451);
or U32543 (N_32543,N_31896,N_31916);
nor U32544 (N_32544,N_30135,N_30458);
or U32545 (N_32545,N_30864,N_31851);
and U32546 (N_32546,N_30140,N_31277);
nand U32547 (N_32547,N_31559,N_31365);
or U32548 (N_32548,N_31350,N_30554);
nor U32549 (N_32549,N_31371,N_31691);
and U32550 (N_32550,N_31231,N_30227);
xnor U32551 (N_32551,N_30945,N_31120);
or U32552 (N_32552,N_31431,N_30972);
and U32553 (N_32553,N_30768,N_31706);
or U32554 (N_32554,N_30350,N_30902);
nand U32555 (N_32555,N_31738,N_30192);
or U32556 (N_32556,N_30335,N_30050);
or U32557 (N_32557,N_31409,N_31166);
xor U32558 (N_32558,N_31219,N_30533);
xor U32559 (N_32559,N_30712,N_30443);
nor U32560 (N_32560,N_31611,N_31435);
nor U32561 (N_32561,N_31960,N_30550);
xor U32562 (N_32562,N_30113,N_30293);
xor U32563 (N_32563,N_30007,N_30343);
nand U32564 (N_32564,N_31024,N_31633);
nand U32565 (N_32565,N_30787,N_30144);
nor U32566 (N_32566,N_31675,N_30651);
and U32567 (N_32567,N_31134,N_31673);
and U32568 (N_32568,N_30915,N_30393);
or U32569 (N_32569,N_31549,N_31213);
nor U32570 (N_32570,N_31831,N_30236);
nand U32571 (N_32571,N_30960,N_30053);
and U32572 (N_32572,N_31082,N_30143);
or U32573 (N_32573,N_30879,N_31143);
nor U32574 (N_32574,N_30264,N_30305);
and U32575 (N_32575,N_30284,N_30178);
or U32576 (N_32576,N_31533,N_30894);
nor U32577 (N_32577,N_30349,N_30467);
nand U32578 (N_32578,N_31037,N_30556);
nand U32579 (N_32579,N_31132,N_31208);
or U32580 (N_32580,N_30588,N_31450);
or U32581 (N_32581,N_31047,N_31137);
or U32582 (N_32582,N_30006,N_30643);
or U32583 (N_32583,N_31808,N_30794);
and U32584 (N_32584,N_30664,N_30598);
xnor U32585 (N_32585,N_31255,N_30776);
nand U32586 (N_32586,N_31067,N_30072);
or U32587 (N_32587,N_31940,N_31936);
or U32588 (N_32588,N_30272,N_31653);
nor U32589 (N_32589,N_31880,N_31123);
xnor U32590 (N_32590,N_31908,N_31869);
nor U32591 (N_32591,N_30090,N_30610);
or U32592 (N_32592,N_30865,N_30703);
nor U32593 (N_32593,N_30383,N_30832);
and U32594 (N_32594,N_31952,N_31406);
and U32595 (N_32595,N_30618,N_30942);
nor U32596 (N_32596,N_30954,N_30256);
nand U32597 (N_32597,N_30154,N_31170);
xnor U32598 (N_32598,N_31986,N_30772);
nor U32599 (N_32599,N_31155,N_30539);
nor U32600 (N_32600,N_30702,N_31572);
xor U32601 (N_32601,N_31259,N_31351);
and U32602 (N_32602,N_30424,N_30781);
nor U32603 (N_32603,N_31805,N_30497);
and U32604 (N_32604,N_30684,N_31015);
or U32605 (N_32605,N_31240,N_31639);
and U32606 (N_32606,N_31416,N_31380);
xnor U32607 (N_32607,N_30692,N_31156);
nor U32608 (N_32608,N_30460,N_31727);
or U32609 (N_32609,N_31813,N_30521);
or U32610 (N_32610,N_31329,N_31544);
xor U32611 (N_32611,N_30519,N_31237);
or U32612 (N_32612,N_30746,N_31623);
or U32613 (N_32613,N_30792,N_30177);
and U32614 (N_32614,N_31078,N_31364);
or U32615 (N_32615,N_31327,N_31959);
nor U32616 (N_32616,N_30750,N_30838);
nor U32617 (N_32617,N_31121,N_31752);
nand U32618 (N_32618,N_31621,N_31250);
nand U32619 (N_32619,N_31097,N_30747);
or U32620 (N_32620,N_31585,N_30804);
nand U32621 (N_32621,N_31985,N_30003);
xor U32622 (N_32622,N_30073,N_31124);
nor U32623 (N_32623,N_30816,N_31784);
nor U32624 (N_32624,N_30935,N_30981);
and U32625 (N_32625,N_30615,N_30014);
and U32626 (N_32626,N_31254,N_30986);
or U32627 (N_32627,N_30980,N_31651);
or U32628 (N_32628,N_31531,N_30534);
xnor U32629 (N_32629,N_31660,N_31839);
nor U32630 (N_32630,N_31230,N_30290);
nand U32631 (N_32631,N_30125,N_31089);
or U32632 (N_32632,N_30496,N_31181);
nand U32633 (N_32633,N_31545,N_30884);
nor U32634 (N_32634,N_30008,N_31634);
nor U32635 (N_32635,N_31601,N_30932);
or U32636 (N_32636,N_30110,N_31730);
xor U32637 (N_32637,N_30123,N_30159);
xor U32638 (N_32638,N_30974,N_31933);
or U32639 (N_32639,N_31681,N_30109);
and U32640 (N_32640,N_30408,N_30968);
or U32641 (N_32641,N_31472,N_30437);
nor U32642 (N_32642,N_30234,N_30371);
xor U32643 (N_32643,N_31322,N_30625);
nor U32644 (N_32644,N_31616,N_30505);
nand U32645 (N_32645,N_31278,N_30310);
and U32646 (N_32646,N_31262,N_31761);
or U32647 (N_32647,N_31027,N_30544);
nor U32648 (N_32648,N_31732,N_31325);
or U32649 (N_32649,N_30317,N_31646);
or U32650 (N_32650,N_31168,N_30604);
nand U32651 (N_32651,N_31367,N_31011);
nor U32652 (N_32652,N_31525,N_30431);
or U32653 (N_32653,N_30193,N_30572);
nor U32654 (N_32654,N_30385,N_31116);
nand U32655 (N_32655,N_30363,N_30257);
and U32656 (N_32656,N_30983,N_31412);
or U32657 (N_32657,N_31861,N_30841);
nor U32658 (N_32658,N_30678,N_31035);
or U32659 (N_32659,N_30943,N_30156);
nand U32660 (N_32660,N_30464,N_31677);
xnor U32661 (N_32661,N_30809,N_30669);
or U32662 (N_32662,N_31465,N_31135);
or U32663 (N_32663,N_31614,N_30433);
nor U32664 (N_32664,N_31847,N_31934);
nand U32665 (N_32665,N_30958,N_31172);
nor U32666 (N_32666,N_30075,N_31684);
xnor U32667 (N_32667,N_31668,N_31207);
nor U32668 (N_32668,N_30299,N_31720);
nand U32669 (N_32669,N_30840,N_31344);
xor U32670 (N_32670,N_30877,N_31625);
or U32671 (N_32671,N_31759,N_30878);
xnor U32672 (N_32672,N_30483,N_31485);
or U32673 (N_32673,N_31102,N_30991);
nor U32674 (N_32674,N_31048,N_30169);
xnor U32675 (N_32675,N_31053,N_30242);
nor U32676 (N_32676,N_31247,N_31227);
xnor U32677 (N_32677,N_31628,N_31333);
xor U32678 (N_32678,N_31848,N_31073);
xor U32679 (N_32679,N_31505,N_31369);
or U32680 (N_32680,N_30280,N_31656);
and U32681 (N_32681,N_30814,N_30255);
and U32682 (N_32682,N_30575,N_30736);
nor U32683 (N_32683,N_30614,N_30306);
or U32684 (N_32684,N_31403,N_30427);
xnor U32685 (N_32685,N_31149,N_30579);
xor U32686 (N_32686,N_30985,N_31827);
and U32687 (N_32687,N_31104,N_30641);
or U32688 (N_32688,N_31711,N_30414);
or U32689 (N_32689,N_30198,N_30415);
xnor U32690 (N_32690,N_31375,N_30511);
or U32691 (N_32691,N_31270,N_31357);
nor U32692 (N_32692,N_31733,N_30773);
nor U32693 (N_32693,N_31138,N_31591);
and U32694 (N_32694,N_30805,N_30962);
and U32695 (N_32695,N_30836,N_31337);
and U32696 (N_32696,N_30672,N_30853);
nor U32697 (N_32697,N_30477,N_31889);
and U32698 (N_32698,N_30866,N_31747);
nor U32699 (N_32699,N_30334,N_30380);
nand U32700 (N_32700,N_31391,N_31760);
nor U32701 (N_32701,N_30710,N_30504);
xor U32702 (N_32702,N_31228,N_31461);
xor U32703 (N_32703,N_30782,N_31257);
or U32704 (N_32704,N_31912,N_30697);
and U32705 (N_32705,N_31862,N_31931);
or U32706 (N_32706,N_31267,N_31291);
xnor U32707 (N_32707,N_30566,N_30373);
nor U32708 (N_32708,N_31907,N_31202);
nor U32709 (N_32709,N_31750,N_30967);
xnor U32710 (N_32710,N_30491,N_30548);
and U32711 (N_32711,N_31577,N_30733);
or U32712 (N_32712,N_30194,N_30462);
nor U32713 (N_32713,N_31452,N_31272);
and U32714 (N_32714,N_30207,N_30793);
xnor U32715 (N_32715,N_30399,N_31771);
nand U32716 (N_32716,N_30851,N_31017);
nand U32717 (N_32717,N_30026,N_31763);
and U32718 (N_32718,N_30000,N_30760);
xor U32719 (N_32719,N_30531,N_31448);
nor U32720 (N_32720,N_31331,N_30890);
or U32721 (N_32721,N_30478,N_30246);
and U32722 (N_32722,N_30569,N_31820);
nor U32723 (N_32723,N_31145,N_30645);
and U32724 (N_32724,N_30819,N_30183);
or U32725 (N_32725,N_30208,N_31370);
nor U32726 (N_32726,N_30691,N_31209);
or U32727 (N_32727,N_31674,N_31363);
or U32728 (N_32728,N_31609,N_31751);
nand U32729 (N_32729,N_31407,N_31537);
nor U32730 (N_32730,N_31643,N_30136);
or U32731 (N_32731,N_30294,N_31271);
nand U32732 (N_32732,N_31619,N_31962);
or U32733 (N_32733,N_31788,N_31564);
nand U32734 (N_32734,N_31682,N_31467);
nand U32735 (N_32735,N_30392,N_30663);
or U32736 (N_32736,N_30626,N_30560);
or U32737 (N_32737,N_30999,N_30619);
or U32738 (N_32738,N_31885,N_31239);
nand U32739 (N_32739,N_30301,N_31098);
nor U32740 (N_32740,N_30362,N_31841);
or U32741 (N_32741,N_31866,N_31818);
xor U32742 (N_32742,N_31980,N_31462);
or U32743 (N_32743,N_31330,N_30704);
or U32744 (N_32744,N_30783,N_30947);
nand U32745 (N_32745,N_31613,N_31324);
nor U32746 (N_32746,N_31842,N_30190);
and U32747 (N_32747,N_30648,N_31891);
or U32748 (N_32748,N_31943,N_30368);
nand U32749 (N_32749,N_31410,N_30720);
xnor U32750 (N_32750,N_30181,N_30346);
nor U32751 (N_32751,N_31221,N_30086);
nor U32752 (N_32752,N_30940,N_31288);
and U32753 (N_32753,N_30087,N_31935);
xor U32754 (N_32754,N_30910,N_30784);
or U32755 (N_32755,N_31229,N_31044);
and U32756 (N_32756,N_31612,N_31117);
nand U32757 (N_32757,N_30808,N_30114);
and U32758 (N_32758,N_30580,N_30587);
or U32759 (N_32759,N_30655,N_30274);
or U32760 (N_32760,N_31383,N_30834);
nor U32761 (N_32761,N_30036,N_31056);
or U32762 (N_32762,N_30253,N_31860);
nor U32763 (N_32763,N_30051,N_30124);
xnor U32764 (N_32764,N_30262,N_31911);
and U32765 (N_32765,N_30547,N_30450);
nand U32766 (N_32766,N_31148,N_30652);
or U32767 (N_32767,N_30111,N_30920);
and U32768 (N_32768,N_30351,N_31777);
and U32769 (N_32769,N_30403,N_31039);
and U32770 (N_32770,N_30622,N_31975);
and U32771 (N_32771,N_30456,N_30005);
and U32772 (N_32772,N_30250,N_30931);
nand U32773 (N_32773,N_30700,N_31058);
and U32774 (N_32774,N_30249,N_31178);
and U32775 (N_32775,N_30698,N_31113);
xnor U32776 (N_32776,N_31829,N_31429);
and U32777 (N_32777,N_31702,N_31826);
xor U32778 (N_32778,N_31234,N_31246);
nand U32779 (N_32779,N_30639,N_31598);
xnor U32780 (N_32780,N_30683,N_30240);
xor U32781 (N_32781,N_31106,N_30089);
xnor U32782 (N_32782,N_30270,N_31792);
nor U32783 (N_32783,N_30248,N_31692);
or U32784 (N_32784,N_30509,N_31323);
or U32785 (N_32785,N_31282,N_30325);
and U32786 (N_32786,N_31071,N_31868);
or U32787 (N_32787,N_31499,N_31447);
nor U32788 (N_32788,N_30057,N_30717);
and U32789 (N_32789,N_31497,N_31714);
nor U32790 (N_32790,N_31045,N_30546);
nand U32791 (N_32791,N_31353,N_31540);
xnor U32792 (N_32792,N_30848,N_31904);
xnor U32793 (N_32793,N_30541,N_31898);
xnor U32794 (N_32794,N_30681,N_31008);
or U32795 (N_32795,N_31527,N_30789);
xor U32796 (N_32796,N_31020,N_31928);
or U32797 (N_32797,N_30723,N_30048);
and U32798 (N_32798,N_30996,N_30098);
xor U32799 (N_32799,N_31419,N_31661);
or U32800 (N_32800,N_31932,N_30429);
nor U32801 (N_32801,N_30975,N_31679);
nor U32802 (N_32802,N_31414,N_30025);
xnor U32803 (N_32803,N_31003,N_31049);
xor U32804 (N_32804,N_31626,N_31206);
xnor U32805 (N_32805,N_31769,N_31128);
nand U32806 (N_32806,N_31355,N_31608);
xor U32807 (N_32807,N_30355,N_31006);
or U32808 (N_32808,N_31950,N_31873);
or U32809 (N_32809,N_31918,N_30818);
xor U32810 (N_32810,N_31583,N_31629);
xor U32811 (N_32811,N_30993,N_30055);
or U32812 (N_32812,N_31764,N_31815);
and U32813 (N_32813,N_31812,N_31602);
or U32814 (N_32814,N_31005,N_31830);
xor U32815 (N_32815,N_30523,N_31397);
nand U32816 (N_32816,N_31988,N_30170);
and U32817 (N_32817,N_31516,N_31993);
nor U32818 (N_32818,N_30059,N_31919);
and U32819 (N_32819,N_31332,N_30341);
xor U32820 (N_32820,N_31019,N_31855);
nand U32821 (N_32821,N_31809,N_31857);
nand U32822 (N_32822,N_30674,N_31072);
or U32823 (N_32823,N_31821,N_31770);
and U32824 (N_32824,N_31552,N_31686);
and U32825 (N_32825,N_31427,N_30602);
nand U32826 (N_32826,N_31644,N_30386);
or U32827 (N_32827,N_31791,N_31604);
or U32828 (N_32828,N_31781,N_31843);
and U32829 (N_32829,N_31088,N_30870);
xor U32830 (N_32830,N_30269,N_30015);
xor U32831 (N_32831,N_30292,N_30455);
and U32832 (N_32832,N_30686,N_30661);
xnor U32833 (N_32833,N_30470,N_31561);
and U32834 (N_32834,N_30374,N_30603);
nor U32835 (N_32835,N_31654,N_30513);
or U32836 (N_32836,N_30206,N_31303);
or U32837 (N_32837,N_30331,N_31176);
and U32838 (N_32838,N_31562,N_31715);
nand U32839 (N_32839,N_30854,N_31127);
or U32840 (N_32840,N_30696,N_30084);
nor U32841 (N_32841,N_30620,N_31007);
nor U32842 (N_32842,N_31014,N_31396);
nor U32843 (N_32843,N_30759,N_31136);
and U32844 (N_32844,N_31052,N_31776);
nand U32845 (N_32845,N_30018,N_31492);
nand U32846 (N_32846,N_31636,N_30039);
or U32847 (N_32847,N_31299,N_31982);
or U32848 (N_32848,N_31532,N_31511);
xnor U32849 (N_32849,N_30067,N_31680);
or U32850 (N_32850,N_30952,N_30876);
or U32851 (N_32851,N_30627,N_31424);
or U32852 (N_32852,N_30791,N_30730);
nor U32853 (N_32853,N_30938,N_30162);
nand U32854 (N_32854,N_30862,N_30540);
xnor U32855 (N_32855,N_31266,N_30898);
nor U32856 (N_32856,N_30682,N_30459);
and U32857 (N_32857,N_31663,N_30861);
or U32858 (N_32858,N_30482,N_30797);
nand U32859 (N_32859,N_30276,N_30011);
nor U32860 (N_32860,N_31248,N_31876);
nand U32861 (N_32861,N_30922,N_31778);
and U32862 (N_32862,N_31785,N_31109);
xor U32863 (N_32863,N_30951,N_30065);
nor U32864 (N_32864,N_30636,N_31285);
nor U32865 (N_32865,N_30314,N_30147);
xor U32866 (N_32866,N_30612,N_30860);
and U32867 (N_32867,N_31173,N_31398);
or U32868 (N_32868,N_30512,N_30751);
xnor U32869 (N_32869,N_31130,N_31814);
nand U32870 (N_32870,N_31914,N_30241);
and U32871 (N_32871,N_30155,N_30108);
nand U32872 (N_32872,N_30753,N_31320);
xor U32873 (N_32873,N_31535,N_31101);
and U32874 (N_32874,N_31144,N_30319);
or U32875 (N_32875,N_31152,N_30874);
nor U32876 (N_32876,N_30167,N_30419);
or U32877 (N_32877,N_31901,N_31177);
nand U32878 (N_32878,N_30821,N_30352);
xor U32879 (N_32879,N_30401,N_31423);
nor U32880 (N_32880,N_31703,N_30160);
nor U32881 (N_32881,N_30056,N_30126);
nand U32882 (N_32882,N_31731,N_30517);
xnor U32883 (N_32883,N_30077,N_31108);
or U32884 (N_32884,N_31103,N_31456);
and U32885 (N_32885,N_31481,N_30680);
and U32886 (N_32886,N_30780,N_31294);
xnor U32887 (N_32887,N_31893,N_31449);
nor U32888 (N_32888,N_30756,N_31100);
xnor U32889 (N_32889,N_30489,N_31606);
nor U32890 (N_32890,N_30737,N_31080);
or U32891 (N_32891,N_31994,N_30268);
nor U32892 (N_32892,N_31179,N_31635);
and U32893 (N_32893,N_31167,N_30396);
nor U32894 (N_32894,N_31182,N_30921);
xor U32895 (N_32895,N_30762,N_30245);
or U32896 (N_32896,N_30465,N_31974);
xnor U32897 (N_32897,N_30345,N_30062);
and U32898 (N_32898,N_31642,N_31051);
xnor U32899 (N_32899,N_31926,N_31373);
xor U32900 (N_32900,N_31268,N_30237);
or U32901 (N_32901,N_30693,N_31084);
xnor U32902 (N_32902,N_30204,N_30474);
nor U32903 (N_32903,N_31062,N_31803);
or U32904 (N_32904,N_30151,N_30989);
nand U32905 (N_32905,N_30763,N_30327);
xor U32906 (N_32906,N_30490,N_30709);
nand U32907 (N_32907,N_30982,N_30122);
nor U32908 (N_32908,N_30348,N_30707);
xnor U32909 (N_32909,N_31310,N_30358);
and U32910 (N_32910,N_30823,N_31944);
and U32911 (N_32911,N_30909,N_30279);
or U32912 (N_32912,N_31196,N_30247);
or U32913 (N_32913,N_31878,N_30297);
or U32914 (N_32914,N_31543,N_30243);
nand U32915 (N_32915,N_31852,N_31724);
and U32916 (N_32916,N_31191,N_30021);
or U32917 (N_32917,N_30581,N_30634);
or U32918 (N_32918,N_30688,N_31297);
or U32919 (N_32919,N_31194,N_31225);
nand U32920 (N_32920,N_31630,N_30452);
xor U32921 (N_32921,N_30356,N_31415);
nor U32922 (N_32922,N_30995,N_30440);
xor U32923 (N_32923,N_31800,N_31002);
and U32924 (N_32924,N_30660,N_30543);
nor U32925 (N_32925,N_31236,N_31316);
or U32926 (N_32926,N_31765,N_31560);
nand U32927 (N_32927,N_30097,N_30033);
and U32928 (N_32928,N_31551,N_31004);
nand U32929 (N_32929,N_30187,N_31915);
and U32930 (N_32930,N_31260,N_31568);
xnor U32931 (N_32931,N_30391,N_30480);
nor U32932 (N_32932,N_31334,N_30551);
and U32933 (N_32933,N_31281,N_30353);
xor U32934 (N_32934,N_30988,N_30171);
nor U32935 (N_32935,N_31232,N_30291);
and U32936 (N_32936,N_31712,N_31193);
xnor U32937 (N_32937,N_31036,N_30646);
nor U32938 (N_32938,N_31594,N_30628);
nand U32939 (N_32939,N_30687,N_30357);
and U32940 (N_32940,N_30601,N_31289);
and U32941 (N_32941,N_31392,N_30589);
nand U32942 (N_32942,N_31662,N_30134);
nor U32943 (N_32943,N_31627,N_31536);
xnor U32944 (N_32944,N_31439,N_31622);
or U32945 (N_32945,N_30775,N_31849);
and U32946 (N_32946,N_31539,N_31217);
nor U32947 (N_32947,N_31929,N_30796);
or U32948 (N_32948,N_31966,N_30060);
xnor U32949 (N_32949,N_30390,N_30914);
or U32950 (N_32950,N_30924,N_30210);
nor U32951 (N_32951,N_30896,N_31846);
and U32952 (N_32952,N_31433,N_31867);
nand U32953 (N_32953,N_30398,N_30195);
nor U32954 (N_32954,N_31586,N_31687);
nor U32955 (N_32955,N_31459,N_31054);
nor U32956 (N_32956,N_30530,N_31022);
xor U32957 (N_32957,N_30623,N_30412);
xor U32958 (N_32958,N_31029,N_31617);
or U32959 (N_32959,N_30378,N_30421);
nor U32960 (N_32960,N_30886,N_31500);
and U32961 (N_32961,N_30803,N_31302);
and U32962 (N_32962,N_31242,N_31664);
and U32963 (N_32963,N_30594,N_31676);
xor U32964 (N_32964,N_31972,N_31346);
xor U32965 (N_32965,N_31514,N_30706);
nor U32966 (N_32966,N_31782,N_30973);
and U32967 (N_32967,N_30637,N_30800);
nor U32968 (N_32968,N_31699,N_30430);
and U32969 (N_32969,N_31405,N_30326);
nand U32970 (N_32970,N_30068,N_31802);
or U32971 (N_32971,N_31464,N_30500);
and U32972 (N_32972,N_31372,N_31010);
or U32973 (N_32973,N_31638,N_31314);
or U32974 (N_32974,N_30320,N_31951);
xnor U32975 (N_32975,N_31094,N_30936);
xor U32976 (N_32976,N_31328,N_31162);
nand U32977 (N_32977,N_30454,N_30863);
and U32978 (N_32978,N_30535,N_30152);
nor U32979 (N_32979,N_31956,N_31810);
nand U32980 (N_32980,N_31902,N_30699);
nand U32981 (N_32981,N_31832,N_30436);
xor U32982 (N_32982,N_31997,N_30563);
and U32983 (N_32983,N_30307,N_31593);
nor U32984 (N_32984,N_30442,N_31618);
nand U32985 (N_32985,N_31737,N_30322);
or U32986 (N_32986,N_31387,N_30285);
nand U32987 (N_32987,N_30501,N_30133);
or U32988 (N_32988,N_31151,N_31032);
and U32989 (N_32989,N_30286,N_30827);
or U32990 (N_32990,N_31954,N_31460);
and U32991 (N_32991,N_30499,N_31762);
xor U32992 (N_32992,N_30209,N_30387);
and U32993 (N_32993,N_31905,N_30277);
xor U32994 (N_32994,N_30228,N_30956);
nand U32995 (N_32995,N_30161,N_31900);
or U32996 (N_32996,N_31286,N_30582);
xnor U32997 (N_32997,N_31963,N_30054);
nand U32998 (N_32998,N_30743,N_30689);
or U32999 (N_32999,N_31797,N_31740);
xor U33000 (N_33000,N_30660,N_30803);
nor U33001 (N_33001,N_30441,N_31337);
or U33002 (N_33002,N_31864,N_31315);
nor U33003 (N_33003,N_30912,N_30078);
nor U33004 (N_33004,N_31772,N_30158);
and U33005 (N_33005,N_30266,N_30827);
and U33006 (N_33006,N_30181,N_30990);
nand U33007 (N_33007,N_30270,N_31247);
xor U33008 (N_33008,N_30487,N_31960);
xor U33009 (N_33009,N_30097,N_30269);
xor U33010 (N_33010,N_31021,N_31731);
nor U33011 (N_33011,N_31130,N_30529);
xor U33012 (N_33012,N_31959,N_31351);
nor U33013 (N_33013,N_31369,N_31442);
nor U33014 (N_33014,N_30320,N_30051);
nand U33015 (N_33015,N_30546,N_30816);
and U33016 (N_33016,N_30302,N_30188);
xnor U33017 (N_33017,N_31822,N_31260);
nor U33018 (N_33018,N_30528,N_31875);
nor U33019 (N_33019,N_31696,N_31983);
xor U33020 (N_33020,N_30481,N_31947);
and U33021 (N_33021,N_31603,N_31851);
nand U33022 (N_33022,N_30123,N_30249);
and U33023 (N_33023,N_30378,N_31804);
or U33024 (N_33024,N_31130,N_31504);
xnor U33025 (N_33025,N_31693,N_30764);
nand U33026 (N_33026,N_30187,N_30834);
xor U33027 (N_33027,N_30718,N_30603);
nand U33028 (N_33028,N_30242,N_31510);
nand U33029 (N_33029,N_30502,N_31905);
and U33030 (N_33030,N_31553,N_31619);
xnor U33031 (N_33031,N_31971,N_31638);
xor U33032 (N_33032,N_31323,N_31306);
nand U33033 (N_33033,N_31108,N_30973);
or U33034 (N_33034,N_31769,N_30604);
nand U33035 (N_33035,N_30302,N_31775);
and U33036 (N_33036,N_31919,N_31033);
nand U33037 (N_33037,N_31943,N_30690);
and U33038 (N_33038,N_31615,N_31548);
and U33039 (N_33039,N_30578,N_30930);
xnor U33040 (N_33040,N_30760,N_31138);
nor U33041 (N_33041,N_30960,N_30718);
xor U33042 (N_33042,N_30045,N_30409);
nor U33043 (N_33043,N_30223,N_31556);
xor U33044 (N_33044,N_31794,N_31415);
nand U33045 (N_33045,N_31257,N_30423);
xor U33046 (N_33046,N_31610,N_30134);
nand U33047 (N_33047,N_30302,N_31203);
nor U33048 (N_33048,N_30711,N_31243);
xor U33049 (N_33049,N_30324,N_31768);
or U33050 (N_33050,N_31994,N_31144);
nor U33051 (N_33051,N_30002,N_31591);
xor U33052 (N_33052,N_31664,N_30669);
xnor U33053 (N_33053,N_31034,N_31963);
nand U33054 (N_33054,N_31474,N_31049);
and U33055 (N_33055,N_30374,N_30498);
nand U33056 (N_33056,N_31409,N_31840);
and U33057 (N_33057,N_30224,N_30859);
and U33058 (N_33058,N_30237,N_31359);
xor U33059 (N_33059,N_30994,N_31603);
nand U33060 (N_33060,N_30570,N_30211);
nand U33061 (N_33061,N_31099,N_30608);
and U33062 (N_33062,N_30372,N_31220);
nand U33063 (N_33063,N_31931,N_30313);
xor U33064 (N_33064,N_30434,N_31096);
nor U33065 (N_33065,N_30652,N_30696);
and U33066 (N_33066,N_30004,N_30299);
nor U33067 (N_33067,N_31704,N_30107);
or U33068 (N_33068,N_30910,N_31008);
nand U33069 (N_33069,N_30350,N_30584);
nand U33070 (N_33070,N_31634,N_30325);
or U33071 (N_33071,N_31748,N_31973);
nand U33072 (N_33072,N_30770,N_30722);
nand U33073 (N_33073,N_31892,N_30361);
or U33074 (N_33074,N_30637,N_30227);
xor U33075 (N_33075,N_31282,N_30634);
or U33076 (N_33076,N_31415,N_30934);
and U33077 (N_33077,N_31288,N_30447);
nand U33078 (N_33078,N_31281,N_31438);
and U33079 (N_33079,N_30303,N_30856);
xor U33080 (N_33080,N_30570,N_31555);
nand U33081 (N_33081,N_31112,N_31243);
xnor U33082 (N_33082,N_31862,N_31409);
nand U33083 (N_33083,N_31335,N_31561);
nor U33084 (N_33084,N_30845,N_30371);
nor U33085 (N_33085,N_30951,N_30352);
nand U33086 (N_33086,N_31736,N_30342);
nand U33087 (N_33087,N_31412,N_30285);
and U33088 (N_33088,N_30706,N_30178);
or U33089 (N_33089,N_31420,N_30666);
nor U33090 (N_33090,N_30683,N_31736);
nand U33091 (N_33091,N_31981,N_31008);
or U33092 (N_33092,N_30692,N_30167);
nand U33093 (N_33093,N_30716,N_31477);
nor U33094 (N_33094,N_30719,N_30466);
nand U33095 (N_33095,N_30631,N_30134);
xnor U33096 (N_33096,N_30648,N_31590);
nor U33097 (N_33097,N_31864,N_30183);
nor U33098 (N_33098,N_30402,N_31880);
xnor U33099 (N_33099,N_30062,N_31933);
nand U33100 (N_33100,N_31044,N_31186);
and U33101 (N_33101,N_30357,N_30353);
xnor U33102 (N_33102,N_31134,N_30270);
and U33103 (N_33103,N_31257,N_30400);
nor U33104 (N_33104,N_31043,N_30865);
and U33105 (N_33105,N_30569,N_31202);
nor U33106 (N_33106,N_31971,N_30072);
nor U33107 (N_33107,N_30780,N_30301);
nor U33108 (N_33108,N_31371,N_31140);
and U33109 (N_33109,N_30545,N_31189);
or U33110 (N_33110,N_31323,N_30901);
and U33111 (N_33111,N_30228,N_30859);
and U33112 (N_33112,N_30884,N_30318);
nor U33113 (N_33113,N_31621,N_30514);
nor U33114 (N_33114,N_30435,N_30521);
or U33115 (N_33115,N_30498,N_30331);
nand U33116 (N_33116,N_30045,N_30350);
or U33117 (N_33117,N_31954,N_31426);
xnor U33118 (N_33118,N_30764,N_31753);
xnor U33119 (N_33119,N_31281,N_31640);
or U33120 (N_33120,N_31203,N_30473);
nor U33121 (N_33121,N_30792,N_31291);
nor U33122 (N_33122,N_31853,N_31325);
xor U33123 (N_33123,N_31240,N_31412);
nor U33124 (N_33124,N_30539,N_31517);
or U33125 (N_33125,N_30286,N_30241);
xnor U33126 (N_33126,N_30237,N_30714);
nor U33127 (N_33127,N_31469,N_30023);
nor U33128 (N_33128,N_31242,N_31647);
nand U33129 (N_33129,N_30977,N_31651);
nor U33130 (N_33130,N_31664,N_30684);
nor U33131 (N_33131,N_31709,N_30469);
or U33132 (N_33132,N_31511,N_31819);
nor U33133 (N_33133,N_30958,N_30684);
and U33134 (N_33134,N_30685,N_30933);
or U33135 (N_33135,N_31561,N_30731);
nand U33136 (N_33136,N_31746,N_31034);
nor U33137 (N_33137,N_30328,N_30750);
xnor U33138 (N_33138,N_30755,N_30851);
nand U33139 (N_33139,N_30945,N_30381);
and U33140 (N_33140,N_30697,N_31886);
xor U33141 (N_33141,N_31777,N_30405);
and U33142 (N_33142,N_30921,N_30331);
or U33143 (N_33143,N_30382,N_30897);
or U33144 (N_33144,N_31589,N_31942);
or U33145 (N_33145,N_31382,N_31637);
nand U33146 (N_33146,N_30270,N_30102);
or U33147 (N_33147,N_30717,N_31602);
nand U33148 (N_33148,N_31198,N_30326);
or U33149 (N_33149,N_31065,N_31725);
xor U33150 (N_33150,N_31038,N_30770);
and U33151 (N_33151,N_31335,N_31371);
nand U33152 (N_33152,N_31888,N_31441);
or U33153 (N_33153,N_31920,N_30644);
nor U33154 (N_33154,N_31646,N_30642);
xor U33155 (N_33155,N_31806,N_30757);
xnor U33156 (N_33156,N_31632,N_31593);
and U33157 (N_33157,N_31168,N_30314);
and U33158 (N_33158,N_30555,N_31526);
xnor U33159 (N_33159,N_30138,N_31193);
and U33160 (N_33160,N_30243,N_30370);
nand U33161 (N_33161,N_31209,N_31664);
or U33162 (N_33162,N_31144,N_30163);
or U33163 (N_33163,N_31320,N_31707);
nand U33164 (N_33164,N_31131,N_30457);
or U33165 (N_33165,N_31729,N_30230);
or U33166 (N_33166,N_30857,N_30354);
xnor U33167 (N_33167,N_30259,N_30951);
or U33168 (N_33168,N_31211,N_31568);
or U33169 (N_33169,N_30185,N_31793);
and U33170 (N_33170,N_31775,N_30878);
xor U33171 (N_33171,N_30618,N_30586);
and U33172 (N_33172,N_30230,N_31481);
or U33173 (N_33173,N_31153,N_31282);
and U33174 (N_33174,N_31422,N_30589);
nor U33175 (N_33175,N_31115,N_30650);
or U33176 (N_33176,N_31767,N_30840);
nand U33177 (N_33177,N_30635,N_31524);
nand U33178 (N_33178,N_30999,N_31852);
or U33179 (N_33179,N_30208,N_30419);
nand U33180 (N_33180,N_31598,N_31163);
and U33181 (N_33181,N_30239,N_31105);
nand U33182 (N_33182,N_30292,N_30784);
or U33183 (N_33183,N_30775,N_30457);
nor U33184 (N_33184,N_31139,N_31750);
xnor U33185 (N_33185,N_30209,N_31457);
or U33186 (N_33186,N_31830,N_31716);
and U33187 (N_33187,N_30263,N_30409);
or U33188 (N_33188,N_30390,N_30011);
nand U33189 (N_33189,N_31496,N_31492);
or U33190 (N_33190,N_30905,N_31011);
xnor U33191 (N_33191,N_31764,N_30106);
or U33192 (N_33192,N_31884,N_30928);
or U33193 (N_33193,N_30137,N_31376);
nor U33194 (N_33194,N_30167,N_31550);
nor U33195 (N_33195,N_31147,N_30629);
nor U33196 (N_33196,N_31504,N_31642);
and U33197 (N_33197,N_31730,N_30850);
xnor U33198 (N_33198,N_31723,N_31770);
or U33199 (N_33199,N_30792,N_30444);
xnor U33200 (N_33200,N_30717,N_31993);
or U33201 (N_33201,N_30030,N_31179);
or U33202 (N_33202,N_31092,N_31884);
nor U33203 (N_33203,N_30176,N_31184);
nor U33204 (N_33204,N_30080,N_30957);
nand U33205 (N_33205,N_30995,N_30273);
and U33206 (N_33206,N_31549,N_31398);
and U33207 (N_33207,N_30488,N_31311);
or U33208 (N_33208,N_30313,N_31824);
and U33209 (N_33209,N_31167,N_31494);
or U33210 (N_33210,N_30501,N_31015);
or U33211 (N_33211,N_31516,N_31770);
nand U33212 (N_33212,N_31031,N_31500);
nor U33213 (N_33213,N_31485,N_30848);
and U33214 (N_33214,N_30960,N_31503);
nor U33215 (N_33215,N_31934,N_30206);
nand U33216 (N_33216,N_31807,N_31695);
and U33217 (N_33217,N_30506,N_30454);
nor U33218 (N_33218,N_31526,N_30404);
nor U33219 (N_33219,N_31914,N_31440);
xnor U33220 (N_33220,N_30669,N_30371);
nor U33221 (N_33221,N_30484,N_31074);
and U33222 (N_33222,N_31841,N_30201);
nand U33223 (N_33223,N_31717,N_31236);
or U33224 (N_33224,N_31807,N_30632);
xor U33225 (N_33225,N_30004,N_31861);
nand U33226 (N_33226,N_30792,N_31701);
and U33227 (N_33227,N_30350,N_30537);
xnor U33228 (N_33228,N_31342,N_31025);
xor U33229 (N_33229,N_30126,N_31156);
xor U33230 (N_33230,N_30381,N_31713);
nand U33231 (N_33231,N_30675,N_31168);
nor U33232 (N_33232,N_30163,N_30735);
nor U33233 (N_33233,N_30894,N_30360);
nand U33234 (N_33234,N_31921,N_31977);
nand U33235 (N_33235,N_31467,N_31567);
nand U33236 (N_33236,N_31410,N_31119);
or U33237 (N_33237,N_31697,N_30036);
nand U33238 (N_33238,N_31907,N_30274);
and U33239 (N_33239,N_30577,N_31135);
nor U33240 (N_33240,N_31130,N_31027);
and U33241 (N_33241,N_30983,N_31173);
and U33242 (N_33242,N_31379,N_31651);
or U33243 (N_33243,N_30793,N_31299);
xnor U33244 (N_33244,N_30508,N_30233);
or U33245 (N_33245,N_30419,N_30954);
and U33246 (N_33246,N_30679,N_31598);
xor U33247 (N_33247,N_30626,N_31155);
xnor U33248 (N_33248,N_31844,N_30739);
nor U33249 (N_33249,N_31734,N_30810);
xor U33250 (N_33250,N_31225,N_31749);
and U33251 (N_33251,N_30730,N_30705);
xor U33252 (N_33252,N_31081,N_30416);
or U33253 (N_33253,N_30042,N_30605);
or U33254 (N_33254,N_30635,N_30752);
and U33255 (N_33255,N_30337,N_30324);
nor U33256 (N_33256,N_31851,N_30723);
or U33257 (N_33257,N_31288,N_30749);
and U33258 (N_33258,N_30761,N_31375);
xnor U33259 (N_33259,N_30265,N_30755);
nand U33260 (N_33260,N_30904,N_31570);
nand U33261 (N_33261,N_30430,N_31275);
nor U33262 (N_33262,N_31322,N_31067);
or U33263 (N_33263,N_30837,N_31828);
xor U33264 (N_33264,N_31908,N_30560);
and U33265 (N_33265,N_31821,N_31900);
and U33266 (N_33266,N_31548,N_30849);
or U33267 (N_33267,N_30369,N_30020);
xor U33268 (N_33268,N_31963,N_31578);
nor U33269 (N_33269,N_30020,N_31014);
and U33270 (N_33270,N_30466,N_30663);
nand U33271 (N_33271,N_30685,N_30527);
and U33272 (N_33272,N_30532,N_31466);
nand U33273 (N_33273,N_31212,N_30117);
and U33274 (N_33274,N_31405,N_31924);
nor U33275 (N_33275,N_31620,N_31974);
nor U33276 (N_33276,N_30725,N_30786);
nor U33277 (N_33277,N_30534,N_30263);
nand U33278 (N_33278,N_30242,N_30249);
nor U33279 (N_33279,N_31247,N_30877);
or U33280 (N_33280,N_30363,N_30808);
nand U33281 (N_33281,N_31241,N_31446);
nand U33282 (N_33282,N_31163,N_31580);
nand U33283 (N_33283,N_31301,N_31278);
xnor U33284 (N_33284,N_30724,N_30726);
xnor U33285 (N_33285,N_30209,N_30277);
nor U33286 (N_33286,N_30979,N_30787);
nor U33287 (N_33287,N_31654,N_30971);
nand U33288 (N_33288,N_31271,N_30812);
or U33289 (N_33289,N_31264,N_30004);
xnor U33290 (N_33290,N_31518,N_31794);
nand U33291 (N_33291,N_30797,N_31893);
and U33292 (N_33292,N_31839,N_30943);
and U33293 (N_33293,N_31223,N_31947);
and U33294 (N_33294,N_30733,N_30856);
nand U33295 (N_33295,N_31316,N_31518);
nand U33296 (N_33296,N_30189,N_31766);
nor U33297 (N_33297,N_31439,N_31805);
and U33298 (N_33298,N_31354,N_31733);
xnor U33299 (N_33299,N_31655,N_30855);
nand U33300 (N_33300,N_31659,N_30214);
nor U33301 (N_33301,N_31397,N_31963);
xnor U33302 (N_33302,N_31507,N_31945);
or U33303 (N_33303,N_31288,N_30668);
xor U33304 (N_33304,N_31561,N_30206);
xnor U33305 (N_33305,N_31749,N_31817);
xor U33306 (N_33306,N_30186,N_31537);
nor U33307 (N_33307,N_31161,N_30942);
xor U33308 (N_33308,N_30981,N_30538);
nand U33309 (N_33309,N_30001,N_31007);
or U33310 (N_33310,N_30264,N_31909);
nor U33311 (N_33311,N_30344,N_30697);
and U33312 (N_33312,N_31564,N_31983);
and U33313 (N_33313,N_31666,N_30940);
nor U33314 (N_33314,N_30891,N_31880);
and U33315 (N_33315,N_30388,N_30241);
or U33316 (N_33316,N_31456,N_31949);
nand U33317 (N_33317,N_31728,N_30565);
and U33318 (N_33318,N_30784,N_31752);
and U33319 (N_33319,N_31159,N_30714);
and U33320 (N_33320,N_30864,N_30031);
nor U33321 (N_33321,N_30518,N_30845);
xnor U33322 (N_33322,N_31558,N_30965);
nand U33323 (N_33323,N_30236,N_31177);
nor U33324 (N_33324,N_30107,N_30157);
nand U33325 (N_33325,N_30310,N_31843);
nor U33326 (N_33326,N_31769,N_30292);
xnor U33327 (N_33327,N_31106,N_30575);
xnor U33328 (N_33328,N_31905,N_30574);
nor U33329 (N_33329,N_31579,N_30973);
xor U33330 (N_33330,N_31223,N_31587);
or U33331 (N_33331,N_30664,N_30404);
nor U33332 (N_33332,N_30269,N_30126);
and U33333 (N_33333,N_30890,N_31877);
or U33334 (N_33334,N_30149,N_31693);
nor U33335 (N_33335,N_31533,N_31366);
or U33336 (N_33336,N_31844,N_30400);
or U33337 (N_33337,N_30147,N_30439);
xor U33338 (N_33338,N_30008,N_31284);
xnor U33339 (N_33339,N_31685,N_30056);
nor U33340 (N_33340,N_30917,N_31096);
or U33341 (N_33341,N_31706,N_31056);
or U33342 (N_33342,N_30129,N_31821);
xnor U33343 (N_33343,N_31799,N_31281);
or U33344 (N_33344,N_30174,N_30508);
and U33345 (N_33345,N_30760,N_30753);
nand U33346 (N_33346,N_30099,N_31604);
or U33347 (N_33347,N_31370,N_30761);
nor U33348 (N_33348,N_31312,N_30081);
nand U33349 (N_33349,N_31095,N_30472);
xor U33350 (N_33350,N_31400,N_31282);
xor U33351 (N_33351,N_31807,N_30489);
nand U33352 (N_33352,N_30367,N_30186);
or U33353 (N_33353,N_30527,N_30251);
or U33354 (N_33354,N_30641,N_31095);
nand U33355 (N_33355,N_31789,N_31467);
or U33356 (N_33356,N_30511,N_31598);
and U33357 (N_33357,N_30994,N_30968);
nand U33358 (N_33358,N_30098,N_30481);
nor U33359 (N_33359,N_30284,N_30818);
and U33360 (N_33360,N_30741,N_31847);
and U33361 (N_33361,N_31775,N_31111);
xor U33362 (N_33362,N_31039,N_30217);
or U33363 (N_33363,N_31181,N_30327);
nor U33364 (N_33364,N_30799,N_30702);
xnor U33365 (N_33365,N_31955,N_30058);
xnor U33366 (N_33366,N_31909,N_31710);
and U33367 (N_33367,N_31173,N_30850);
nor U33368 (N_33368,N_30275,N_30370);
and U33369 (N_33369,N_30497,N_30718);
nand U33370 (N_33370,N_31375,N_31294);
nor U33371 (N_33371,N_31949,N_31218);
nor U33372 (N_33372,N_31564,N_30223);
and U33373 (N_33373,N_30619,N_30954);
nand U33374 (N_33374,N_31496,N_31553);
nor U33375 (N_33375,N_31573,N_31644);
nand U33376 (N_33376,N_30929,N_30922);
and U33377 (N_33377,N_30808,N_31638);
or U33378 (N_33378,N_30547,N_31522);
xnor U33379 (N_33379,N_31853,N_30621);
nand U33380 (N_33380,N_30950,N_31595);
xor U33381 (N_33381,N_31160,N_30823);
nand U33382 (N_33382,N_31651,N_31771);
xnor U33383 (N_33383,N_31149,N_31659);
nor U33384 (N_33384,N_31762,N_30296);
or U33385 (N_33385,N_30946,N_31464);
nor U33386 (N_33386,N_30551,N_30157);
xor U33387 (N_33387,N_31192,N_30611);
xor U33388 (N_33388,N_30764,N_30342);
nand U33389 (N_33389,N_30943,N_31688);
xnor U33390 (N_33390,N_30746,N_30516);
xnor U33391 (N_33391,N_31185,N_31647);
or U33392 (N_33392,N_31413,N_31292);
or U33393 (N_33393,N_30228,N_30484);
and U33394 (N_33394,N_30860,N_30544);
or U33395 (N_33395,N_31512,N_30919);
xnor U33396 (N_33396,N_30526,N_31388);
nor U33397 (N_33397,N_31235,N_31536);
or U33398 (N_33398,N_30972,N_30061);
and U33399 (N_33399,N_30801,N_30068);
nor U33400 (N_33400,N_30805,N_31176);
nand U33401 (N_33401,N_30744,N_31307);
nor U33402 (N_33402,N_31580,N_30257);
nand U33403 (N_33403,N_31733,N_31382);
xnor U33404 (N_33404,N_31102,N_30654);
nand U33405 (N_33405,N_31308,N_30082);
nor U33406 (N_33406,N_30033,N_30964);
nand U33407 (N_33407,N_30131,N_31222);
or U33408 (N_33408,N_31300,N_31353);
nand U33409 (N_33409,N_31214,N_31397);
or U33410 (N_33410,N_31233,N_30250);
nand U33411 (N_33411,N_31362,N_31747);
nand U33412 (N_33412,N_30074,N_31562);
xnor U33413 (N_33413,N_30433,N_31292);
nor U33414 (N_33414,N_30823,N_31763);
or U33415 (N_33415,N_31338,N_30153);
nor U33416 (N_33416,N_31037,N_31320);
nand U33417 (N_33417,N_30787,N_31786);
nand U33418 (N_33418,N_30503,N_30412);
nand U33419 (N_33419,N_30151,N_31635);
xor U33420 (N_33420,N_30560,N_31452);
or U33421 (N_33421,N_30809,N_30207);
xnor U33422 (N_33422,N_31009,N_31589);
xnor U33423 (N_33423,N_31362,N_30382);
xnor U33424 (N_33424,N_30082,N_30851);
and U33425 (N_33425,N_30166,N_30865);
or U33426 (N_33426,N_30306,N_31744);
nand U33427 (N_33427,N_31538,N_30087);
nor U33428 (N_33428,N_31849,N_30855);
or U33429 (N_33429,N_30717,N_30401);
xnor U33430 (N_33430,N_31023,N_31644);
or U33431 (N_33431,N_31204,N_31646);
nor U33432 (N_33432,N_30875,N_31588);
nor U33433 (N_33433,N_31505,N_31467);
xor U33434 (N_33434,N_30009,N_31753);
and U33435 (N_33435,N_30477,N_31381);
xnor U33436 (N_33436,N_31137,N_31446);
or U33437 (N_33437,N_31141,N_30930);
and U33438 (N_33438,N_31577,N_30572);
nand U33439 (N_33439,N_30133,N_31288);
and U33440 (N_33440,N_31241,N_30286);
nand U33441 (N_33441,N_31715,N_30784);
nor U33442 (N_33442,N_30928,N_30783);
and U33443 (N_33443,N_31815,N_30544);
or U33444 (N_33444,N_30112,N_31151);
nand U33445 (N_33445,N_30346,N_30929);
nor U33446 (N_33446,N_31887,N_30938);
nand U33447 (N_33447,N_31312,N_30010);
or U33448 (N_33448,N_31352,N_30022);
xor U33449 (N_33449,N_31206,N_30797);
xnor U33450 (N_33450,N_30293,N_30416);
nor U33451 (N_33451,N_30675,N_31575);
and U33452 (N_33452,N_30881,N_31223);
xnor U33453 (N_33453,N_31097,N_30983);
or U33454 (N_33454,N_30190,N_30679);
nand U33455 (N_33455,N_31339,N_30134);
nand U33456 (N_33456,N_31291,N_31723);
nor U33457 (N_33457,N_31532,N_30554);
nor U33458 (N_33458,N_31742,N_31455);
xnor U33459 (N_33459,N_30355,N_30811);
or U33460 (N_33460,N_31664,N_30651);
and U33461 (N_33461,N_31371,N_31117);
or U33462 (N_33462,N_31369,N_30350);
and U33463 (N_33463,N_30970,N_31991);
nand U33464 (N_33464,N_30949,N_31970);
nor U33465 (N_33465,N_30372,N_30391);
nand U33466 (N_33466,N_30183,N_30056);
xnor U33467 (N_33467,N_30760,N_30438);
and U33468 (N_33468,N_31068,N_30210);
xor U33469 (N_33469,N_31624,N_30087);
and U33470 (N_33470,N_31539,N_30679);
nor U33471 (N_33471,N_30384,N_30967);
and U33472 (N_33472,N_30226,N_30937);
nand U33473 (N_33473,N_30859,N_30274);
or U33474 (N_33474,N_30565,N_31391);
nand U33475 (N_33475,N_30193,N_31860);
nor U33476 (N_33476,N_31344,N_31444);
or U33477 (N_33477,N_31092,N_31143);
nor U33478 (N_33478,N_30393,N_31265);
or U33479 (N_33479,N_31379,N_30083);
and U33480 (N_33480,N_31959,N_30701);
and U33481 (N_33481,N_31838,N_30236);
nor U33482 (N_33482,N_30218,N_31753);
and U33483 (N_33483,N_30798,N_31633);
and U33484 (N_33484,N_31697,N_31164);
and U33485 (N_33485,N_31819,N_30808);
and U33486 (N_33486,N_31736,N_31702);
nor U33487 (N_33487,N_31525,N_31832);
or U33488 (N_33488,N_31155,N_31563);
nor U33489 (N_33489,N_30897,N_31328);
nand U33490 (N_33490,N_31664,N_31247);
and U33491 (N_33491,N_31207,N_31596);
and U33492 (N_33492,N_30102,N_30747);
and U33493 (N_33493,N_30896,N_30010);
and U33494 (N_33494,N_30934,N_30095);
or U33495 (N_33495,N_30545,N_30299);
or U33496 (N_33496,N_30939,N_30444);
nor U33497 (N_33497,N_31369,N_30633);
or U33498 (N_33498,N_30505,N_31102);
and U33499 (N_33499,N_31004,N_31864);
and U33500 (N_33500,N_31278,N_31774);
and U33501 (N_33501,N_30907,N_30220);
or U33502 (N_33502,N_30265,N_31416);
nor U33503 (N_33503,N_30112,N_30421);
and U33504 (N_33504,N_31290,N_30029);
nor U33505 (N_33505,N_30820,N_31180);
nor U33506 (N_33506,N_31235,N_31897);
and U33507 (N_33507,N_30417,N_30302);
or U33508 (N_33508,N_31846,N_30830);
or U33509 (N_33509,N_30768,N_30106);
or U33510 (N_33510,N_30774,N_30130);
nor U33511 (N_33511,N_31649,N_30651);
or U33512 (N_33512,N_31969,N_30191);
and U33513 (N_33513,N_30773,N_30537);
or U33514 (N_33514,N_30781,N_30861);
and U33515 (N_33515,N_31698,N_30987);
or U33516 (N_33516,N_31258,N_30092);
xnor U33517 (N_33517,N_30777,N_31798);
or U33518 (N_33518,N_31465,N_31085);
nor U33519 (N_33519,N_31110,N_31998);
nand U33520 (N_33520,N_30854,N_31128);
and U33521 (N_33521,N_31190,N_30282);
and U33522 (N_33522,N_31309,N_31050);
nor U33523 (N_33523,N_30886,N_30508);
nor U33524 (N_33524,N_30311,N_30276);
nand U33525 (N_33525,N_31016,N_30404);
or U33526 (N_33526,N_30582,N_30506);
nand U33527 (N_33527,N_30814,N_31573);
and U33528 (N_33528,N_30866,N_31817);
or U33529 (N_33529,N_30551,N_30747);
nand U33530 (N_33530,N_30059,N_30517);
or U33531 (N_33531,N_30743,N_30856);
nand U33532 (N_33532,N_31428,N_31992);
nand U33533 (N_33533,N_30370,N_30857);
or U33534 (N_33534,N_30015,N_30888);
or U33535 (N_33535,N_30633,N_31866);
nor U33536 (N_33536,N_31169,N_31705);
nor U33537 (N_33537,N_31353,N_31516);
nand U33538 (N_33538,N_31924,N_30366);
and U33539 (N_33539,N_31838,N_30545);
xor U33540 (N_33540,N_30491,N_31122);
nor U33541 (N_33541,N_31939,N_30222);
nor U33542 (N_33542,N_31872,N_31532);
nand U33543 (N_33543,N_31873,N_30360);
or U33544 (N_33544,N_31768,N_31184);
or U33545 (N_33545,N_31063,N_31552);
nor U33546 (N_33546,N_31487,N_31416);
nand U33547 (N_33547,N_31621,N_30429);
xnor U33548 (N_33548,N_31276,N_30167);
or U33549 (N_33549,N_30096,N_30367);
xnor U33550 (N_33550,N_30507,N_30810);
xor U33551 (N_33551,N_31154,N_31002);
nor U33552 (N_33552,N_31600,N_31597);
or U33553 (N_33553,N_30529,N_30640);
or U33554 (N_33554,N_30081,N_31964);
nand U33555 (N_33555,N_31598,N_30308);
or U33556 (N_33556,N_30178,N_31068);
or U33557 (N_33557,N_31149,N_31756);
xor U33558 (N_33558,N_30188,N_30406);
nor U33559 (N_33559,N_31009,N_30851);
nor U33560 (N_33560,N_30272,N_31567);
and U33561 (N_33561,N_31940,N_30060);
nor U33562 (N_33562,N_30599,N_30522);
or U33563 (N_33563,N_31531,N_30640);
or U33564 (N_33564,N_30553,N_31974);
and U33565 (N_33565,N_30459,N_30789);
and U33566 (N_33566,N_31081,N_30047);
and U33567 (N_33567,N_31583,N_31987);
xnor U33568 (N_33568,N_30199,N_31726);
and U33569 (N_33569,N_30077,N_31213);
nor U33570 (N_33570,N_31160,N_30076);
xor U33571 (N_33571,N_31168,N_30980);
and U33572 (N_33572,N_30547,N_30185);
nand U33573 (N_33573,N_31911,N_30962);
nand U33574 (N_33574,N_30104,N_31496);
nor U33575 (N_33575,N_31929,N_31075);
or U33576 (N_33576,N_30026,N_31004);
or U33577 (N_33577,N_30505,N_31916);
or U33578 (N_33578,N_30695,N_30050);
and U33579 (N_33579,N_30457,N_31822);
and U33580 (N_33580,N_31348,N_31241);
nor U33581 (N_33581,N_31612,N_31540);
nor U33582 (N_33582,N_30219,N_31410);
nand U33583 (N_33583,N_30927,N_31005);
or U33584 (N_33584,N_30501,N_31806);
xor U33585 (N_33585,N_31981,N_31582);
nand U33586 (N_33586,N_30942,N_31067);
xnor U33587 (N_33587,N_31011,N_30440);
nand U33588 (N_33588,N_30066,N_30496);
nand U33589 (N_33589,N_30836,N_31196);
nand U33590 (N_33590,N_31308,N_30765);
nand U33591 (N_33591,N_31806,N_31881);
nand U33592 (N_33592,N_31690,N_31681);
nor U33593 (N_33593,N_31233,N_30245);
nand U33594 (N_33594,N_31705,N_31829);
or U33595 (N_33595,N_30024,N_31561);
nor U33596 (N_33596,N_30140,N_31930);
or U33597 (N_33597,N_30804,N_30716);
nand U33598 (N_33598,N_31947,N_31046);
nand U33599 (N_33599,N_30889,N_31986);
xor U33600 (N_33600,N_30658,N_30309);
or U33601 (N_33601,N_30337,N_30629);
xor U33602 (N_33602,N_30181,N_31867);
xor U33603 (N_33603,N_30450,N_30801);
or U33604 (N_33604,N_31901,N_30570);
or U33605 (N_33605,N_31191,N_30894);
and U33606 (N_33606,N_31204,N_30453);
nor U33607 (N_33607,N_30558,N_31076);
xnor U33608 (N_33608,N_31342,N_31192);
xnor U33609 (N_33609,N_30600,N_30283);
nor U33610 (N_33610,N_31541,N_30391);
xor U33611 (N_33611,N_30937,N_31764);
nor U33612 (N_33612,N_30121,N_30117);
or U33613 (N_33613,N_30472,N_31496);
or U33614 (N_33614,N_31076,N_31334);
and U33615 (N_33615,N_30632,N_31422);
nand U33616 (N_33616,N_31088,N_31365);
nor U33617 (N_33617,N_31691,N_31414);
nor U33618 (N_33618,N_30947,N_31666);
xnor U33619 (N_33619,N_31764,N_31828);
nor U33620 (N_33620,N_30478,N_31612);
xnor U33621 (N_33621,N_30538,N_30548);
nand U33622 (N_33622,N_30312,N_30476);
xor U33623 (N_33623,N_31307,N_30141);
nor U33624 (N_33624,N_30540,N_31139);
xor U33625 (N_33625,N_30274,N_30760);
xnor U33626 (N_33626,N_31637,N_30095);
nand U33627 (N_33627,N_30901,N_30619);
or U33628 (N_33628,N_31235,N_30610);
or U33629 (N_33629,N_31363,N_31776);
nor U33630 (N_33630,N_30963,N_30347);
nand U33631 (N_33631,N_31970,N_31066);
nand U33632 (N_33632,N_30575,N_31467);
and U33633 (N_33633,N_31238,N_31273);
xor U33634 (N_33634,N_31243,N_31730);
nand U33635 (N_33635,N_30743,N_31847);
or U33636 (N_33636,N_30349,N_31776);
or U33637 (N_33637,N_31439,N_30630);
or U33638 (N_33638,N_31690,N_30470);
and U33639 (N_33639,N_31815,N_30685);
nand U33640 (N_33640,N_30729,N_30368);
nor U33641 (N_33641,N_31331,N_30569);
xnor U33642 (N_33642,N_31813,N_31852);
and U33643 (N_33643,N_31051,N_31985);
nand U33644 (N_33644,N_30482,N_30167);
or U33645 (N_33645,N_31770,N_31568);
xor U33646 (N_33646,N_31230,N_31909);
nand U33647 (N_33647,N_31981,N_31127);
and U33648 (N_33648,N_31509,N_31092);
nor U33649 (N_33649,N_30314,N_30460);
nor U33650 (N_33650,N_31783,N_31620);
nand U33651 (N_33651,N_30291,N_31704);
or U33652 (N_33652,N_31015,N_30380);
and U33653 (N_33653,N_31818,N_31858);
nand U33654 (N_33654,N_31497,N_31336);
xnor U33655 (N_33655,N_31656,N_30347);
or U33656 (N_33656,N_31284,N_30670);
xor U33657 (N_33657,N_30566,N_30514);
xor U33658 (N_33658,N_30840,N_31088);
and U33659 (N_33659,N_30018,N_30115);
nand U33660 (N_33660,N_31303,N_30438);
nor U33661 (N_33661,N_30482,N_30671);
nand U33662 (N_33662,N_31503,N_30061);
xor U33663 (N_33663,N_30594,N_31417);
nor U33664 (N_33664,N_30595,N_31309);
nand U33665 (N_33665,N_30144,N_31127);
nand U33666 (N_33666,N_30253,N_31909);
nor U33667 (N_33667,N_31679,N_31518);
xor U33668 (N_33668,N_31398,N_31943);
or U33669 (N_33669,N_31735,N_30430);
nand U33670 (N_33670,N_30640,N_31269);
or U33671 (N_33671,N_31221,N_31664);
xor U33672 (N_33672,N_31970,N_31440);
nand U33673 (N_33673,N_30987,N_30384);
xnor U33674 (N_33674,N_31729,N_30435);
nand U33675 (N_33675,N_31749,N_30651);
or U33676 (N_33676,N_31129,N_30792);
nor U33677 (N_33677,N_31170,N_31037);
and U33678 (N_33678,N_30280,N_30706);
nor U33679 (N_33679,N_30182,N_30890);
nand U33680 (N_33680,N_30269,N_30334);
nor U33681 (N_33681,N_30573,N_31159);
nand U33682 (N_33682,N_30773,N_30345);
and U33683 (N_33683,N_31831,N_31196);
nand U33684 (N_33684,N_30949,N_30970);
nor U33685 (N_33685,N_31564,N_30486);
xnor U33686 (N_33686,N_31536,N_30219);
and U33687 (N_33687,N_31966,N_31432);
nand U33688 (N_33688,N_30240,N_30746);
nor U33689 (N_33689,N_31066,N_31817);
nand U33690 (N_33690,N_31386,N_31346);
nor U33691 (N_33691,N_30080,N_30738);
and U33692 (N_33692,N_31776,N_31537);
nand U33693 (N_33693,N_31081,N_31678);
nand U33694 (N_33694,N_30637,N_30751);
nor U33695 (N_33695,N_31732,N_30143);
nand U33696 (N_33696,N_30475,N_30935);
or U33697 (N_33697,N_31295,N_31458);
and U33698 (N_33698,N_30066,N_30265);
nor U33699 (N_33699,N_31759,N_31704);
xor U33700 (N_33700,N_31145,N_30998);
nand U33701 (N_33701,N_30578,N_31147);
or U33702 (N_33702,N_30713,N_31887);
nand U33703 (N_33703,N_31913,N_31368);
and U33704 (N_33704,N_30242,N_31731);
nand U33705 (N_33705,N_31711,N_30997);
xnor U33706 (N_33706,N_31542,N_30015);
xor U33707 (N_33707,N_30508,N_31489);
xor U33708 (N_33708,N_30615,N_30905);
xor U33709 (N_33709,N_30231,N_31554);
or U33710 (N_33710,N_31981,N_31985);
or U33711 (N_33711,N_30636,N_31611);
nand U33712 (N_33712,N_31304,N_31414);
and U33713 (N_33713,N_30914,N_31975);
and U33714 (N_33714,N_31227,N_31418);
nor U33715 (N_33715,N_30519,N_31669);
or U33716 (N_33716,N_30662,N_30091);
nor U33717 (N_33717,N_30038,N_30178);
or U33718 (N_33718,N_31051,N_31973);
or U33719 (N_33719,N_30294,N_31806);
or U33720 (N_33720,N_31769,N_31524);
or U33721 (N_33721,N_30999,N_31866);
or U33722 (N_33722,N_31769,N_31869);
or U33723 (N_33723,N_30427,N_30597);
and U33724 (N_33724,N_30323,N_30544);
or U33725 (N_33725,N_31236,N_30847);
xor U33726 (N_33726,N_30707,N_30452);
xnor U33727 (N_33727,N_31853,N_30908);
xor U33728 (N_33728,N_30448,N_31506);
or U33729 (N_33729,N_30512,N_31110);
nor U33730 (N_33730,N_31371,N_31535);
and U33731 (N_33731,N_30315,N_31579);
nand U33732 (N_33732,N_30916,N_31095);
or U33733 (N_33733,N_31758,N_30815);
or U33734 (N_33734,N_30250,N_31575);
or U33735 (N_33735,N_31588,N_31281);
nor U33736 (N_33736,N_31796,N_30394);
nand U33737 (N_33737,N_30884,N_31454);
xnor U33738 (N_33738,N_30608,N_30674);
nor U33739 (N_33739,N_31770,N_31615);
or U33740 (N_33740,N_31789,N_31315);
or U33741 (N_33741,N_30675,N_31770);
or U33742 (N_33742,N_30561,N_31458);
and U33743 (N_33743,N_30192,N_31419);
and U33744 (N_33744,N_31932,N_30058);
and U33745 (N_33745,N_30237,N_30185);
or U33746 (N_33746,N_30146,N_31308);
or U33747 (N_33747,N_30822,N_31373);
xnor U33748 (N_33748,N_31478,N_30370);
nor U33749 (N_33749,N_30151,N_30387);
nor U33750 (N_33750,N_31069,N_31039);
xnor U33751 (N_33751,N_30379,N_31875);
xnor U33752 (N_33752,N_31928,N_31991);
nand U33753 (N_33753,N_30148,N_30835);
xnor U33754 (N_33754,N_31239,N_30770);
or U33755 (N_33755,N_31025,N_30034);
xnor U33756 (N_33756,N_30202,N_31901);
nor U33757 (N_33757,N_31613,N_31598);
xnor U33758 (N_33758,N_30262,N_30769);
and U33759 (N_33759,N_31542,N_31404);
or U33760 (N_33760,N_30540,N_30344);
or U33761 (N_33761,N_30499,N_30166);
nor U33762 (N_33762,N_30060,N_31989);
xor U33763 (N_33763,N_31572,N_30378);
and U33764 (N_33764,N_30734,N_30168);
xnor U33765 (N_33765,N_30238,N_31538);
nand U33766 (N_33766,N_30550,N_30694);
or U33767 (N_33767,N_30735,N_30161);
nand U33768 (N_33768,N_31383,N_31831);
or U33769 (N_33769,N_31961,N_31846);
xor U33770 (N_33770,N_30105,N_31330);
xnor U33771 (N_33771,N_31718,N_31845);
xnor U33772 (N_33772,N_30628,N_30326);
or U33773 (N_33773,N_30886,N_31610);
and U33774 (N_33774,N_30688,N_30457);
nand U33775 (N_33775,N_30528,N_31508);
or U33776 (N_33776,N_31477,N_31409);
or U33777 (N_33777,N_31893,N_30398);
nor U33778 (N_33778,N_30402,N_30305);
nand U33779 (N_33779,N_31487,N_31747);
and U33780 (N_33780,N_30847,N_31092);
or U33781 (N_33781,N_31558,N_31905);
nor U33782 (N_33782,N_31649,N_31903);
or U33783 (N_33783,N_31502,N_31845);
or U33784 (N_33784,N_31254,N_30339);
or U33785 (N_33785,N_30250,N_30717);
nor U33786 (N_33786,N_30702,N_30631);
xor U33787 (N_33787,N_31150,N_30830);
xnor U33788 (N_33788,N_31169,N_30841);
nor U33789 (N_33789,N_31897,N_31688);
nand U33790 (N_33790,N_30277,N_30759);
nor U33791 (N_33791,N_31339,N_31161);
and U33792 (N_33792,N_30636,N_30110);
nor U33793 (N_33793,N_30692,N_31177);
xnor U33794 (N_33794,N_31238,N_31808);
xnor U33795 (N_33795,N_31893,N_31845);
nor U33796 (N_33796,N_31566,N_31763);
and U33797 (N_33797,N_30274,N_31307);
xnor U33798 (N_33798,N_30916,N_31500);
or U33799 (N_33799,N_30866,N_30578);
xnor U33800 (N_33800,N_31890,N_31717);
or U33801 (N_33801,N_30308,N_30712);
nand U33802 (N_33802,N_31007,N_30126);
nand U33803 (N_33803,N_30048,N_30078);
and U33804 (N_33804,N_31737,N_31273);
nor U33805 (N_33805,N_31074,N_31440);
nand U33806 (N_33806,N_31588,N_30750);
or U33807 (N_33807,N_31920,N_31606);
nand U33808 (N_33808,N_30563,N_30212);
or U33809 (N_33809,N_30860,N_30732);
xor U33810 (N_33810,N_30846,N_31657);
xnor U33811 (N_33811,N_31538,N_31758);
nor U33812 (N_33812,N_31691,N_30540);
nor U33813 (N_33813,N_30553,N_31025);
nor U33814 (N_33814,N_30371,N_30414);
nand U33815 (N_33815,N_30718,N_30581);
and U33816 (N_33816,N_30295,N_31347);
and U33817 (N_33817,N_30538,N_30528);
and U33818 (N_33818,N_31673,N_31628);
or U33819 (N_33819,N_31953,N_31051);
or U33820 (N_33820,N_30420,N_31606);
nor U33821 (N_33821,N_31761,N_31815);
nor U33822 (N_33822,N_30226,N_31995);
or U33823 (N_33823,N_31619,N_31735);
nor U33824 (N_33824,N_31439,N_31087);
and U33825 (N_33825,N_31448,N_31462);
and U33826 (N_33826,N_31148,N_30471);
xor U33827 (N_33827,N_30529,N_31441);
and U33828 (N_33828,N_30386,N_31218);
xor U33829 (N_33829,N_30796,N_31308);
and U33830 (N_33830,N_31103,N_30693);
nor U33831 (N_33831,N_31535,N_31268);
and U33832 (N_33832,N_31092,N_31942);
nand U33833 (N_33833,N_30651,N_30304);
nand U33834 (N_33834,N_31023,N_30615);
xor U33835 (N_33835,N_30554,N_31178);
and U33836 (N_33836,N_30442,N_30317);
nor U33837 (N_33837,N_31300,N_30444);
nand U33838 (N_33838,N_30383,N_31172);
nor U33839 (N_33839,N_31734,N_30924);
xor U33840 (N_33840,N_31153,N_31836);
xor U33841 (N_33841,N_31235,N_31784);
xnor U33842 (N_33842,N_30594,N_30535);
xor U33843 (N_33843,N_31458,N_30558);
xor U33844 (N_33844,N_31790,N_31187);
or U33845 (N_33845,N_31297,N_30801);
nand U33846 (N_33846,N_31156,N_30975);
and U33847 (N_33847,N_31592,N_31619);
xor U33848 (N_33848,N_31286,N_31431);
nor U33849 (N_33849,N_31044,N_30000);
and U33850 (N_33850,N_31941,N_30907);
nand U33851 (N_33851,N_30085,N_30925);
xor U33852 (N_33852,N_30478,N_31082);
xnor U33853 (N_33853,N_30070,N_30915);
nand U33854 (N_33854,N_30797,N_30503);
nand U33855 (N_33855,N_31322,N_31949);
nand U33856 (N_33856,N_30215,N_30791);
nand U33857 (N_33857,N_30124,N_30118);
or U33858 (N_33858,N_31520,N_30210);
nand U33859 (N_33859,N_31898,N_31158);
or U33860 (N_33860,N_31510,N_31207);
nor U33861 (N_33861,N_31770,N_31773);
nor U33862 (N_33862,N_30537,N_31683);
and U33863 (N_33863,N_31259,N_31600);
nor U33864 (N_33864,N_30262,N_30360);
or U33865 (N_33865,N_30866,N_30656);
or U33866 (N_33866,N_30139,N_30456);
nand U33867 (N_33867,N_30313,N_30928);
or U33868 (N_33868,N_31484,N_30913);
and U33869 (N_33869,N_30008,N_30326);
nand U33870 (N_33870,N_30222,N_31851);
nor U33871 (N_33871,N_31475,N_30273);
and U33872 (N_33872,N_30040,N_30717);
or U33873 (N_33873,N_30065,N_31334);
and U33874 (N_33874,N_31851,N_30670);
or U33875 (N_33875,N_30888,N_30459);
xnor U33876 (N_33876,N_30641,N_30578);
and U33877 (N_33877,N_31491,N_31322);
and U33878 (N_33878,N_31499,N_30313);
and U33879 (N_33879,N_31334,N_30811);
xnor U33880 (N_33880,N_30269,N_30175);
xnor U33881 (N_33881,N_30229,N_31048);
or U33882 (N_33882,N_30127,N_31434);
and U33883 (N_33883,N_30824,N_31481);
xor U33884 (N_33884,N_30953,N_30414);
and U33885 (N_33885,N_31976,N_30375);
nor U33886 (N_33886,N_30128,N_31851);
nand U33887 (N_33887,N_31157,N_31574);
and U33888 (N_33888,N_30797,N_30446);
and U33889 (N_33889,N_31064,N_31958);
nand U33890 (N_33890,N_31012,N_31822);
nand U33891 (N_33891,N_30073,N_31989);
and U33892 (N_33892,N_31301,N_30649);
and U33893 (N_33893,N_30087,N_30353);
xnor U33894 (N_33894,N_30451,N_30379);
nor U33895 (N_33895,N_30573,N_30477);
and U33896 (N_33896,N_31498,N_31041);
xnor U33897 (N_33897,N_31634,N_30466);
nor U33898 (N_33898,N_31835,N_30306);
and U33899 (N_33899,N_30546,N_30271);
or U33900 (N_33900,N_30674,N_30365);
nand U33901 (N_33901,N_30753,N_31585);
and U33902 (N_33902,N_31568,N_31543);
nand U33903 (N_33903,N_30777,N_31305);
and U33904 (N_33904,N_31153,N_31389);
nor U33905 (N_33905,N_30808,N_31620);
nor U33906 (N_33906,N_31225,N_31109);
xor U33907 (N_33907,N_31440,N_31495);
nand U33908 (N_33908,N_30141,N_30178);
xnor U33909 (N_33909,N_31612,N_31079);
nor U33910 (N_33910,N_31822,N_30690);
nand U33911 (N_33911,N_31314,N_30981);
and U33912 (N_33912,N_30314,N_30121);
nand U33913 (N_33913,N_30872,N_31899);
xor U33914 (N_33914,N_30091,N_30453);
and U33915 (N_33915,N_30458,N_30072);
or U33916 (N_33916,N_30400,N_30816);
xnor U33917 (N_33917,N_31554,N_31997);
nor U33918 (N_33918,N_30351,N_31380);
xor U33919 (N_33919,N_30921,N_30454);
nand U33920 (N_33920,N_31056,N_31304);
or U33921 (N_33921,N_31495,N_31502);
nor U33922 (N_33922,N_30634,N_30419);
xnor U33923 (N_33923,N_31612,N_31174);
nor U33924 (N_33924,N_30921,N_31097);
and U33925 (N_33925,N_31143,N_30324);
nand U33926 (N_33926,N_31439,N_31219);
xnor U33927 (N_33927,N_30770,N_30920);
or U33928 (N_33928,N_30570,N_31543);
nand U33929 (N_33929,N_30162,N_31546);
or U33930 (N_33930,N_30855,N_31108);
nand U33931 (N_33931,N_30366,N_31832);
or U33932 (N_33932,N_31809,N_31905);
xnor U33933 (N_33933,N_30670,N_31512);
nor U33934 (N_33934,N_31737,N_31655);
and U33935 (N_33935,N_31475,N_30408);
nand U33936 (N_33936,N_31506,N_31677);
and U33937 (N_33937,N_31275,N_30428);
and U33938 (N_33938,N_30570,N_31363);
nor U33939 (N_33939,N_30277,N_30826);
nand U33940 (N_33940,N_31211,N_30737);
xor U33941 (N_33941,N_30884,N_30107);
xor U33942 (N_33942,N_31181,N_30642);
nand U33943 (N_33943,N_30434,N_30117);
or U33944 (N_33944,N_30253,N_30378);
nand U33945 (N_33945,N_30745,N_30254);
nand U33946 (N_33946,N_30140,N_30089);
nand U33947 (N_33947,N_30178,N_30809);
xnor U33948 (N_33948,N_31340,N_30208);
nor U33949 (N_33949,N_31448,N_30331);
nor U33950 (N_33950,N_31562,N_31429);
or U33951 (N_33951,N_31218,N_30239);
nor U33952 (N_33952,N_30599,N_30612);
and U33953 (N_33953,N_30424,N_30969);
nor U33954 (N_33954,N_31153,N_30950);
nor U33955 (N_33955,N_31948,N_31371);
or U33956 (N_33956,N_31460,N_31451);
xor U33957 (N_33957,N_31050,N_31784);
xor U33958 (N_33958,N_31003,N_30777);
xnor U33959 (N_33959,N_30440,N_30354);
and U33960 (N_33960,N_30108,N_30890);
or U33961 (N_33961,N_30500,N_30473);
or U33962 (N_33962,N_30054,N_30989);
nor U33963 (N_33963,N_31450,N_30222);
nand U33964 (N_33964,N_31383,N_30397);
or U33965 (N_33965,N_30812,N_31943);
or U33966 (N_33966,N_30689,N_30007);
and U33967 (N_33967,N_31558,N_30834);
xor U33968 (N_33968,N_30750,N_31344);
or U33969 (N_33969,N_31395,N_30614);
nor U33970 (N_33970,N_30174,N_31840);
xnor U33971 (N_33971,N_31820,N_31842);
or U33972 (N_33972,N_30530,N_30857);
nand U33973 (N_33973,N_31649,N_30842);
xor U33974 (N_33974,N_31985,N_30890);
nand U33975 (N_33975,N_31431,N_30321);
nand U33976 (N_33976,N_31537,N_31713);
and U33977 (N_33977,N_31163,N_30123);
or U33978 (N_33978,N_31753,N_31425);
or U33979 (N_33979,N_31526,N_30742);
nor U33980 (N_33980,N_30852,N_30758);
nor U33981 (N_33981,N_30749,N_31228);
xnor U33982 (N_33982,N_30885,N_31997);
nand U33983 (N_33983,N_31722,N_30532);
or U33984 (N_33984,N_31522,N_31034);
xnor U33985 (N_33985,N_30980,N_30734);
and U33986 (N_33986,N_31879,N_30082);
nand U33987 (N_33987,N_30363,N_31284);
nor U33988 (N_33988,N_31825,N_31350);
nand U33989 (N_33989,N_31669,N_30432);
nor U33990 (N_33990,N_30987,N_31406);
xnor U33991 (N_33991,N_30482,N_31457);
and U33992 (N_33992,N_31175,N_30403);
and U33993 (N_33993,N_31014,N_31046);
or U33994 (N_33994,N_30874,N_30435);
nor U33995 (N_33995,N_30352,N_30697);
and U33996 (N_33996,N_30474,N_31422);
nand U33997 (N_33997,N_31590,N_30405);
or U33998 (N_33998,N_31333,N_31818);
xnor U33999 (N_33999,N_31034,N_30567);
xnor U34000 (N_34000,N_33864,N_33268);
or U34001 (N_34001,N_33229,N_33859);
xor U34002 (N_34002,N_33944,N_33773);
xnor U34003 (N_34003,N_32731,N_33187);
or U34004 (N_34004,N_32776,N_32068);
xnor U34005 (N_34005,N_32429,N_32348);
xor U34006 (N_34006,N_33048,N_33263);
xnor U34007 (N_34007,N_33219,N_32524);
and U34008 (N_34008,N_32922,N_32054);
or U34009 (N_34009,N_32224,N_32093);
nor U34010 (N_34010,N_32114,N_33493);
nand U34011 (N_34011,N_33490,N_32080);
nor U34012 (N_34012,N_33200,N_32069);
nand U34013 (N_34013,N_32651,N_33030);
or U34014 (N_34014,N_32852,N_32896);
or U34015 (N_34015,N_32029,N_32109);
xor U34016 (N_34016,N_33081,N_32540);
xnor U34017 (N_34017,N_33166,N_33655);
nor U34018 (N_34018,N_33561,N_33999);
nand U34019 (N_34019,N_33651,N_33499);
xnor U34020 (N_34020,N_32799,N_32070);
nand U34021 (N_34021,N_32181,N_33188);
nor U34022 (N_34022,N_32211,N_32486);
or U34023 (N_34023,N_32479,N_32312);
or U34024 (N_34024,N_32753,N_33452);
or U34025 (N_34025,N_33280,N_33356);
nor U34026 (N_34026,N_32930,N_33389);
nand U34027 (N_34027,N_32280,N_33282);
or U34028 (N_34028,N_32763,N_33871);
nand U34029 (N_34029,N_32291,N_33050);
nand U34030 (N_34030,N_33421,N_32563);
nor U34031 (N_34031,N_33932,N_33772);
nand U34032 (N_34032,N_33752,N_33558);
nor U34033 (N_34033,N_32624,N_33956);
nor U34034 (N_34034,N_33982,N_33007);
or U34035 (N_34035,N_32106,N_33427);
nand U34036 (N_34036,N_32047,N_32640);
or U34037 (N_34037,N_33438,N_33748);
nor U34038 (N_34038,N_33235,N_33617);
and U34039 (N_34039,N_32172,N_33258);
nand U34040 (N_34040,N_33986,N_32285);
nand U34041 (N_34041,N_33112,N_33509);
nand U34042 (N_34042,N_32633,N_32391);
and U34043 (N_34043,N_32078,N_32893);
or U34044 (N_34044,N_32822,N_32977);
nand U34045 (N_34045,N_33082,N_32597);
nand U34046 (N_34046,N_33261,N_32673);
nor U34047 (N_34047,N_32081,N_33898);
nand U34048 (N_34048,N_32571,N_33766);
xor U34049 (N_34049,N_32733,N_33096);
nand U34050 (N_34050,N_33425,N_32694);
nor U34051 (N_34051,N_33878,N_33073);
nor U34052 (N_34052,N_32341,N_33259);
and U34053 (N_34053,N_32873,N_32046);
nor U34054 (N_34054,N_32842,N_32333);
and U34055 (N_34055,N_33355,N_33338);
and U34056 (N_34056,N_33315,N_32905);
or U34057 (N_34057,N_32750,N_33114);
and U34058 (N_34058,N_32838,N_32385);
and U34059 (N_34059,N_32553,N_32236);
nor U34060 (N_34060,N_32511,N_32064);
nor U34061 (N_34061,N_32695,N_33636);
or U34062 (N_34062,N_33309,N_32482);
nand U34063 (N_34063,N_33650,N_32796);
nand U34064 (N_34064,N_33819,N_33829);
and U34065 (N_34065,N_33202,N_33323);
nand U34066 (N_34066,N_32543,N_33199);
nor U34067 (N_34067,N_32184,N_33808);
nand U34068 (N_34068,N_33983,N_33256);
and U34069 (N_34069,N_32840,N_33845);
nor U34070 (N_34070,N_32092,N_33844);
nor U34071 (N_34071,N_33693,N_33092);
and U34072 (N_34072,N_33669,N_33093);
nand U34073 (N_34073,N_32743,N_33987);
xor U34074 (N_34074,N_33622,N_33977);
xnor U34075 (N_34075,N_33747,N_33190);
nor U34076 (N_34076,N_33423,N_33530);
or U34077 (N_34077,N_33086,N_33273);
or U34078 (N_34078,N_33821,N_32659);
or U34079 (N_34079,N_32661,N_32386);
xor U34080 (N_34080,N_33279,N_33002);
xnor U34081 (N_34081,N_32306,N_32336);
or U34082 (N_34082,N_33415,N_33457);
nand U34083 (N_34083,N_33569,N_33919);
nand U34084 (N_34084,N_33991,N_32805);
xor U34085 (N_34085,N_33632,N_32666);
nor U34086 (N_34086,N_32992,N_32042);
xnor U34087 (N_34087,N_32883,N_33573);
nor U34088 (N_34088,N_32084,N_32300);
xor U34089 (N_34089,N_32376,N_33441);
or U34090 (N_34090,N_33248,N_33550);
nand U34091 (N_34091,N_32574,N_33469);
nor U34092 (N_34092,N_32460,N_33284);
xor U34093 (N_34093,N_32755,N_33520);
and U34094 (N_34094,N_33948,N_32803);
xor U34095 (N_34095,N_32797,N_33954);
xor U34096 (N_34096,N_32589,N_32611);
nand U34097 (N_34097,N_32477,N_32710);
nor U34098 (N_34098,N_33385,N_32494);
or U34099 (N_34099,N_33619,N_32667);
nand U34100 (N_34100,N_32531,N_32798);
or U34101 (N_34101,N_33095,N_33787);
nand U34102 (N_34102,N_32990,N_33176);
xor U34103 (N_34103,N_33091,N_33465);
nand U34104 (N_34104,N_33146,N_32945);
or U34105 (N_34105,N_33137,N_32168);
nand U34106 (N_34106,N_32848,N_32706);
and U34107 (N_34107,N_32475,N_32235);
nor U34108 (N_34108,N_32186,N_33387);
nand U34109 (N_34109,N_32973,N_32968);
nand U34110 (N_34110,N_33697,N_33236);
nand U34111 (N_34111,N_32222,N_32095);
nor U34112 (N_34112,N_33475,N_32271);
or U34113 (N_34113,N_32427,N_33797);
xor U34114 (N_34114,N_33739,N_32630);
and U34115 (N_34115,N_32538,N_33957);
nand U34116 (N_34116,N_33147,N_32394);
nand U34117 (N_34117,N_32768,N_32950);
xor U34118 (N_34118,N_33156,N_32520);
or U34119 (N_34119,N_33910,N_33401);
and U34120 (N_34120,N_32578,N_32573);
or U34121 (N_34121,N_33927,N_32780);
nor U34122 (N_34122,N_33350,N_32588);
xnor U34123 (N_34123,N_33643,N_33313);
or U34124 (N_34124,N_33865,N_33684);
and U34125 (N_34125,N_32672,N_32503);
nor U34126 (N_34126,N_32396,N_32153);
or U34127 (N_34127,N_33471,N_33270);
nand U34128 (N_34128,N_33902,N_32119);
or U34129 (N_34129,N_33241,N_32432);
nor U34130 (N_34130,N_33311,N_33726);
and U34131 (N_34131,N_33319,N_33388);
xor U34132 (N_34132,N_33770,N_33064);
nor U34133 (N_34133,N_33782,N_33310);
and U34134 (N_34134,N_33790,N_32875);
nand U34135 (N_34135,N_32554,N_33394);
nand U34136 (N_34136,N_32652,N_32674);
xor U34137 (N_34137,N_32721,N_33897);
nor U34138 (N_34138,N_32227,N_32147);
and U34139 (N_34139,N_32980,N_32263);
nor U34140 (N_34140,N_33005,N_32898);
nor U34141 (N_34141,N_33379,N_33157);
xor U34142 (N_34142,N_32139,N_32193);
and U34143 (N_34143,N_32861,N_32966);
or U34144 (N_34144,N_32121,N_32491);
nor U34145 (N_34145,N_32827,N_32732);
nand U34146 (N_34146,N_33523,N_33283);
nor U34147 (N_34147,N_33195,N_32877);
or U34148 (N_34148,N_33209,N_32473);
xor U34149 (N_34149,N_32365,N_33646);
xor U34150 (N_34150,N_32997,N_33866);
nand U34151 (N_34151,N_33854,N_32602);
xor U34152 (N_34152,N_32343,N_33083);
xnor U34153 (N_34153,N_33160,N_32603);
xor U34154 (N_34154,N_32495,N_32577);
nand U34155 (N_34155,N_32202,N_32175);
and U34156 (N_34156,N_33227,N_33847);
xor U34157 (N_34157,N_33333,N_32485);
nor U34158 (N_34158,N_33447,N_32372);
and U34159 (N_34159,N_33481,N_33788);
or U34160 (N_34160,N_33049,N_32471);
nand U34161 (N_34161,N_33367,N_33488);
nand U34162 (N_34162,N_32065,N_32665);
or U34163 (N_34163,N_32041,N_32294);
xor U34164 (N_34164,N_33969,N_32606);
and U34165 (N_34165,N_33963,N_32819);
nand U34166 (N_34166,N_33408,N_33706);
or U34167 (N_34167,N_33761,N_32214);
xnor U34168 (N_34168,N_32981,N_32387);
and U34169 (N_34169,N_33217,N_33774);
xor U34170 (N_34170,N_32794,N_33721);
xor U34171 (N_34171,N_32051,N_33124);
nor U34172 (N_34172,N_32276,N_32252);
xor U34173 (N_34173,N_32159,N_32157);
or U34174 (N_34174,N_32982,N_32444);
xnor U34175 (N_34175,N_32539,N_32650);
or U34176 (N_34176,N_32496,N_32259);
and U34177 (N_34177,N_32585,N_32257);
xnor U34178 (N_34178,N_33103,N_33760);
or U34179 (N_34179,N_33640,N_33665);
nand U34180 (N_34180,N_32584,N_32632);
xnor U34181 (N_34181,N_33710,N_33216);
nor U34182 (N_34182,N_32105,N_33119);
and U34183 (N_34183,N_33541,N_33915);
nor U34184 (N_34184,N_33744,N_32392);
or U34185 (N_34185,N_33140,N_33574);
nand U34186 (N_34186,N_33317,N_33487);
nor U34187 (N_34187,N_32649,N_32789);
nand U34188 (N_34188,N_33123,N_32956);
or U34189 (N_34189,N_33153,N_32845);
xnor U34190 (N_34190,N_33508,N_32870);
and U34191 (N_34191,N_33841,N_32914);
and U34192 (N_34192,N_33476,N_33656);
and U34193 (N_34193,N_32298,N_33719);
nand U34194 (N_34194,N_33564,N_32761);
nand U34195 (N_34195,N_33567,N_33247);
nand U34196 (N_34196,N_33113,N_32498);
or U34197 (N_34197,N_32124,N_33330);
nand U34198 (N_34198,N_32442,N_33911);
and U34199 (N_34199,N_33513,N_33221);
nand U34200 (N_34200,N_32897,N_33627);
and U34201 (N_34201,N_32687,N_32366);
nand U34202 (N_34202,N_32424,N_33998);
nand U34203 (N_34203,N_32703,N_33712);
nand U34204 (N_34204,N_32150,N_33392);
or U34205 (N_34205,N_32804,N_33322);
and U34206 (N_34206,N_32003,N_33604);
or U34207 (N_34207,N_33725,N_33729);
xnor U34208 (N_34208,N_32836,N_32268);
xor U34209 (N_34209,N_32132,N_32036);
and U34210 (N_34210,N_33715,N_33295);
nand U34211 (N_34211,N_32087,N_33357);
nor U34212 (N_34212,N_33529,N_32638);
xor U34213 (N_34213,N_32868,N_32592);
and U34214 (N_34214,N_32621,N_33435);
nand U34215 (N_34215,N_33633,N_32851);
nand U34216 (N_34216,N_32828,N_33110);
nand U34217 (N_34217,N_33132,N_33758);
or U34218 (N_34218,N_33664,N_32814);
nand U34219 (N_34219,N_33439,N_32413);
and U34220 (N_34220,N_33934,N_33139);
or U34221 (N_34221,N_32729,N_32567);
nor U34222 (N_34222,N_33009,N_33131);
xnor U34223 (N_34223,N_32217,N_33560);
or U34224 (N_34224,N_33237,N_32024);
nor U34225 (N_34225,N_33344,N_32718);
nor U34226 (N_34226,N_32762,N_32209);
xnor U34227 (N_34227,N_32240,N_32648);
or U34228 (N_34228,N_32908,N_32942);
nor U34229 (N_34229,N_33728,N_32690);
xnor U34230 (N_34230,N_32233,N_33399);
xnor U34231 (N_34231,N_33533,N_32198);
or U34232 (N_34232,N_32337,N_32452);
xnor U34233 (N_34233,N_33659,N_33730);
nor U34234 (N_34234,N_33252,N_32140);
nand U34235 (N_34235,N_32936,N_32742);
and U34236 (N_34236,N_32253,N_32112);
nand U34237 (N_34237,N_32691,N_32944);
nor U34238 (N_34238,N_32974,N_32170);
nor U34239 (N_34239,N_32931,N_33716);
or U34240 (N_34240,N_32062,N_33159);
xnor U34241 (N_34241,N_33674,N_32351);
xor U34242 (N_34242,N_32408,N_32130);
nand U34243 (N_34243,N_33738,N_33046);
nor U34244 (N_34244,N_33945,N_33026);
nand U34245 (N_34245,N_32519,N_32142);
nand U34246 (N_34246,N_32484,N_32255);
xnor U34247 (N_34247,N_33035,N_32660);
or U34248 (N_34248,N_33965,N_33253);
xnor U34249 (N_34249,N_32244,N_33928);
nand U34250 (N_34250,N_32013,N_33211);
or U34251 (N_34251,N_32226,N_33691);
xnor U34252 (N_34252,N_32404,N_32704);
and U34253 (N_34253,N_33763,N_33873);
nor U34254 (N_34254,N_33565,N_33568);
xnor U34255 (N_34255,N_32515,N_33489);
xnor U34256 (N_34256,N_33653,N_32039);
and U34257 (N_34257,N_32894,N_33437);
or U34258 (N_34258,N_32456,N_33251);
xor U34259 (N_34259,N_32685,N_32018);
nand U34260 (N_34260,N_33833,N_33006);
and U34261 (N_34261,N_33740,N_32698);
or U34262 (N_34262,N_33352,N_33177);
nor U34263 (N_34263,N_33661,N_33305);
nor U34264 (N_34264,N_33792,N_32085);
nand U34265 (N_34265,N_33791,N_33862);
or U34266 (N_34266,N_32760,N_32215);
or U34267 (N_34267,N_32565,N_33224);
or U34268 (N_34268,N_32994,N_33807);
nand U34269 (N_34269,N_33714,N_33165);
nand U34270 (N_34270,N_32192,N_33364);
xnor U34271 (N_34271,N_33486,N_33491);
nand U34272 (N_34272,N_33825,N_32960);
xor U34273 (N_34273,N_33800,N_33215);
or U34274 (N_34274,N_32418,N_32537);
xor U34275 (N_34275,N_33801,N_32635);
nand U34276 (N_34276,N_33828,N_32608);
nor U34277 (N_34277,N_32216,N_33750);
and U34278 (N_34278,N_32869,N_33984);
or U34279 (N_34279,N_32247,N_32523);
and U34280 (N_34280,N_33585,N_33501);
and U34281 (N_34281,N_32979,N_33810);
or U34282 (N_34282,N_32824,N_33014);
or U34283 (N_34283,N_32714,N_32508);
xnor U34284 (N_34284,N_32900,N_33180);
nor U34285 (N_34285,N_33522,N_32162);
and U34286 (N_34286,N_33345,N_33542);
nor U34287 (N_34287,N_32110,N_33278);
nor U34288 (N_34288,N_32976,N_33053);
xor U34289 (N_34289,N_33056,N_33128);
or U34290 (N_34290,N_33966,N_33127);
xnor U34291 (N_34291,N_32127,N_33588);
and U34292 (N_34292,N_33074,N_33170);
and U34293 (N_34293,N_32670,N_32582);
or U34294 (N_34294,N_33802,N_33861);
or U34295 (N_34295,N_32034,N_33813);
nand U34296 (N_34296,N_33996,N_33886);
and U34297 (N_34297,N_32813,N_32111);
nand U34298 (N_34298,N_33168,N_32527);
nand U34299 (N_34299,N_32405,N_33985);
nand U34300 (N_34300,N_32658,N_33134);
nor U34301 (N_34301,N_33173,N_32746);
nor U34302 (N_34302,N_33855,N_32783);
nand U34303 (N_34303,N_32536,N_32361);
nand U34304 (N_34304,N_33135,N_32438);
or U34305 (N_34305,N_33548,N_33973);
nand U34306 (N_34306,N_33941,N_33610);
and U34307 (N_34307,N_32200,N_33608);
xor U34308 (N_34308,N_32604,N_32810);
nor U34309 (N_34309,N_33045,N_33938);
nor U34310 (N_34310,N_33296,N_33361);
nand U34311 (N_34311,N_32786,N_33746);
and U34312 (N_34312,N_33495,N_33018);
xnor U34313 (N_34313,N_33794,N_33250);
or U34314 (N_34314,N_32073,N_33198);
or U34315 (N_34315,N_32411,N_33600);
nor U34316 (N_34316,N_32628,N_33894);
xnor U34317 (N_34317,N_33276,N_33848);
or U34318 (N_34318,N_33578,N_33582);
and U34319 (N_34319,N_33875,N_32579);
and U34320 (N_34320,N_33901,N_32135);
or U34321 (N_34321,N_32448,N_32885);
xor U34322 (N_34322,N_33281,N_32481);
nand U34323 (N_34323,N_32711,N_33989);
xor U34324 (N_34324,N_33274,N_32229);
and U34325 (N_34325,N_33353,N_32008);
and U34326 (N_34326,N_33230,N_33926);
nand U34327 (N_34327,N_33196,N_32664);
nor U34328 (N_34328,N_32451,N_32656);
xor U34329 (N_34329,N_32251,N_33396);
nand U34330 (N_34330,N_32120,N_33803);
nor U34331 (N_34331,N_33857,N_32262);
nand U34332 (N_34332,N_33454,N_33593);
xnor U34333 (N_34333,N_33576,N_33930);
nand U34334 (N_34334,N_33020,N_32195);
xor U34335 (N_34335,N_32339,N_32561);
and U34336 (N_34336,N_32260,N_33868);
or U34337 (N_34337,N_32547,N_33637);
xor U34338 (N_34338,N_33406,N_32590);
or U34339 (N_34339,N_32097,N_32330);
nor U34340 (N_34340,N_32434,N_32359);
and U34341 (N_34341,N_33291,N_33806);
xnor U34342 (N_34342,N_33990,N_32360);
and U34343 (N_34343,N_32282,N_32188);
and U34344 (N_34344,N_33167,N_32915);
nand U34345 (N_34345,N_32014,N_33480);
nand U34346 (N_34346,N_33122,N_33683);
nand U34347 (N_34347,N_33887,N_32802);
xor U34348 (N_34348,N_32946,N_32518);
and U34349 (N_34349,N_33673,N_33070);
xor U34350 (N_34350,N_32199,N_32340);
xor U34351 (N_34351,N_32774,N_33470);
xor U34352 (N_34352,N_32548,N_32100);
and U34353 (N_34353,N_33613,N_32161);
nor U34354 (N_34354,N_33374,N_33877);
xor U34355 (N_34355,N_33440,N_32975);
nor U34356 (N_34356,N_32983,N_32472);
and U34357 (N_34357,N_32775,N_33347);
or U34358 (N_34358,N_32232,N_32395);
or U34359 (N_34359,N_33511,N_33144);
nand U34360 (N_34360,N_32772,N_32594);
and U34361 (N_34361,N_32220,N_33949);
or U34362 (N_34362,N_33223,N_33572);
or U34363 (N_34363,N_32788,N_32212);
nand U34364 (N_34364,N_32812,N_32962);
nor U34365 (N_34365,N_33702,N_32959);
nor U34366 (N_34366,N_32045,N_32735);
nand U34367 (N_34367,N_33366,N_32254);
and U34368 (N_34368,N_33312,N_32402);
xnor U34369 (N_34369,N_32927,N_33909);
xnor U34370 (N_34370,N_33449,N_33359);
nor U34371 (N_34371,N_33097,N_33734);
xor U34372 (N_34372,N_33880,N_32581);
or U34373 (N_34373,N_32430,N_32862);
xnor U34374 (N_34374,N_33753,N_33431);
nand U34375 (N_34375,N_32843,N_32249);
and U34376 (N_34376,N_32154,N_33072);
nand U34377 (N_34377,N_32952,N_32323);
or U34378 (N_34378,N_33686,N_33039);
nand U34379 (N_34379,N_33155,N_33556);
xnor U34380 (N_34380,N_33069,N_32194);
xor U34381 (N_34381,N_33946,N_32899);
nand U34382 (N_34382,N_32307,N_32301);
nor U34383 (N_34383,N_32693,N_33596);
or U34384 (N_34384,N_33913,N_33519);
and U34385 (N_34385,N_32368,N_32700);
nor U34386 (N_34386,N_32420,N_33587);
and U34387 (N_34387,N_32378,N_32598);
nor U34388 (N_34388,N_33321,N_32270);
nand U34389 (N_34389,N_32010,N_32474);
or U34390 (N_34390,N_33876,N_32770);
or U34391 (N_34391,N_32441,N_33436);
and U34392 (N_34392,N_32948,N_33755);
or U34393 (N_34393,N_33277,N_33300);
nor U34394 (N_34394,N_32855,N_33076);
nor U34395 (N_34395,N_32075,N_33346);
nor U34396 (N_34396,N_32492,N_33951);
or U34397 (N_34397,N_33759,N_33382);
and U34398 (N_34398,N_33444,N_32514);
nand U34399 (N_34399,N_33265,N_32910);
and U34400 (N_34400,N_33502,N_32144);
nand U34401 (N_34401,N_32071,N_33785);
or U34402 (N_34402,N_33171,N_33301);
nor U34403 (N_34403,N_33583,N_32723);
nand U34404 (N_34404,N_33955,N_33084);
or U34405 (N_34405,N_32933,N_32044);
or U34406 (N_34406,N_32532,N_33642);
nor U34407 (N_34407,N_33395,N_33022);
and U34408 (N_34408,N_33243,N_33192);
xnor U34409 (N_34409,N_33370,N_33889);
nand U34410 (N_34410,N_33872,N_32715);
and U34411 (N_34411,N_32911,N_33586);
nor U34412 (N_34412,N_32559,N_33013);
xor U34413 (N_34413,N_33334,N_33041);
nor U34414 (N_34414,N_33384,N_33733);
nor U34415 (N_34415,N_32586,N_33545);
or U34416 (N_34416,N_33667,N_32642);
xnor U34417 (N_34417,N_33240,N_33975);
xnor U34418 (N_34418,N_32857,N_32744);
nand U34419 (N_34419,N_32790,N_33818);
xnor U34420 (N_34420,N_33205,N_33138);
nand U34421 (N_34421,N_33834,N_33109);
nand U34422 (N_34422,N_32655,N_33704);
nand U34423 (N_34423,N_32679,N_32709);
nand U34424 (N_34424,N_33705,N_33724);
and U34425 (N_34425,N_33152,N_32439);
xnor U34426 (N_34426,N_33843,N_32208);
nand U34427 (N_34427,N_33443,N_32978);
nand U34428 (N_34428,N_32443,N_32072);
xor U34429 (N_34429,N_33467,N_32499);
nor U34430 (N_34430,N_32707,N_33019);
nand U34431 (N_34431,N_32191,N_33879);
xor U34432 (N_34432,N_33590,N_32066);
and U34433 (N_34433,N_32388,N_33094);
xnor U34434 (N_34434,N_33515,N_33078);
nand U34435 (N_34435,N_32516,N_33145);
xor U34436 (N_34436,N_33940,N_33777);
nand U34437 (N_34437,N_32015,N_33809);
or U34438 (N_34438,N_32461,N_33972);
and U34439 (N_34439,N_32422,N_33459);
or U34440 (N_34440,N_33722,N_32230);
nor U34441 (N_34441,N_33822,N_32128);
xor U34442 (N_34442,N_32767,N_33057);
nand U34443 (N_34443,N_32089,N_32412);
and U34444 (N_34444,N_32446,N_33290);
and U34445 (N_34445,N_33950,N_33668);
xnor U34446 (N_34446,N_33101,N_32844);
and U34447 (N_34447,N_33182,N_33654);
and U34448 (N_34448,N_33612,N_33105);
and U34449 (N_34449,N_32053,N_32273);
nand U34450 (N_34450,N_32146,N_33824);
and U34451 (N_34451,N_33472,N_32613);
or U34452 (N_34452,N_32326,N_33194);
and U34453 (N_34453,N_33837,N_32925);
nor U34454 (N_34454,N_32390,N_32784);
nand U34455 (N_34455,N_32304,N_32445);
nand U34456 (N_34456,N_33936,N_33121);
nor U34457 (N_34457,N_32712,N_33479);
nor U34458 (N_34458,N_32489,N_32309);
xnor U34459 (N_34459,N_32591,N_33689);
nor U34460 (N_34460,N_33430,N_32887);
nor U34461 (N_34461,N_32373,N_32688);
or U34462 (N_34462,N_33186,N_32795);
nand U34463 (N_34463,N_33115,N_33089);
nor U34464 (N_34464,N_32859,N_33641);
xor U34465 (N_34465,N_33918,N_33635);
and U34466 (N_34466,N_33553,N_32464);
or U34467 (N_34467,N_32345,N_32141);
nand U34468 (N_34468,N_32740,N_33796);
and U34469 (N_34469,N_33713,N_32916);
xnor U34470 (N_34470,N_32371,N_33197);
nand U34471 (N_34471,N_33061,N_32864);
and U34472 (N_34472,N_32699,N_32277);
or U34473 (N_34473,N_33671,N_33953);
nand U34474 (N_34474,N_33500,N_32004);
or U34475 (N_34475,N_32145,N_32826);
nand U34476 (N_34476,N_32171,N_33962);
xor U34477 (N_34477,N_32834,N_32937);
xor U34478 (N_34478,N_32808,N_32605);
or U34479 (N_34479,N_32654,N_33598);
xnor U34480 (N_34480,N_33781,N_32480);
nand U34481 (N_34481,N_32414,N_33212);
and U34482 (N_34482,N_33870,N_33085);
nor U34483 (N_34483,N_32169,N_32137);
or U34484 (N_34484,N_33660,N_32818);
nor U34485 (N_34485,N_33275,N_32022);
xnor U34486 (N_34486,N_33191,N_33151);
and U34487 (N_34487,N_32506,N_33011);
nor U34488 (N_34488,N_33831,N_33756);
nor U34489 (N_34489,N_32860,N_33566);
nand U34490 (N_34490,N_32028,N_33757);
or U34491 (N_34491,N_32399,N_32383);
nor U34492 (N_34492,N_32210,N_32256);
nor U34493 (N_34493,N_33997,N_33360);
or U34494 (N_34494,N_33980,N_33474);
and U34495 (N_34495,N_33368,N_33605);
nor U34496 (N_34496,N_33618,N_33043);
nand U34497 (N_34497,N_32196,N_32580);
or U34498 (N_34498,N_33647,N_33639);
xnor U34499 (N_34499,N_33099,N_32009);
and U34500 (N_34500,N_32149,N_32017);
xnor U34501 (N_34501,N_33891,N_33448);
or U34502 (N_34502,N_33851,N_32281);
nor U34503 (N_34503,N_32355,N_32926);
or U34504 (N_34504,N_33468,N_32040);
nor U34505 (N_34505,N_33771,N_33682);
or U34506 (N_34506,N_32689,N_33193);
and U34507 (N_34507,N_33414,N_33117);
and U34508 (N_34508,N_33850,N_32314);
xor U34509 (N_34509,N_32286,N_32421);
or U34510 (N_34510,N_33544,N_32874);
nor U34511 (N_34511,N_32542,N_33994);
or U34512 (N_34512,N_33885,N_32310);
nand U34513 (N_34513,N_32143,N_33412);
and U34514 (N_34514,N_32791,N_32048);
xnor U34515 (N_34515,N_33783,N_32639);
xor U34516 (N_34516,N_32940,N_33287);
or U34517 (N_34517,N_33342,N_33442);
and U34518 (N_34518,N_33185,N_33688);
and U34519 (N_34519,N_33775,N_32758);
nand U34520 (N_34520,N_33079,N_33884);
and U34521 (N_34521,N_33776,N_33979);
xor U34522 (N_34522,N_33547,N_33174);
nor U34523 (N_34523,N_33858,N_33225);
and U34524 (N_34524,N_33737,N_33521);
nor U34525 (N_34525,N_32025,N_33672);
nor U34526 (N_34526,N_32713,N_32002);
and U34527 (N_34527,N_32423,N_32043);
and U34528 (N_34528,N_32657,N_33175);
and U34529 (N_34529,N_33010,N_32830);
nand U34530 (N_34530,N_33077,N_32021);
or U34531 (N_34531,N_32264,N_32354);
or U34532 (N_34532,N_32030,N_33696);
and U34533 (N_34533,N_32165,N_32367);
xor U34534 (N_34534,N_33524,N_32705);
xnor U34535 (N_34535,N_32401,N_32500);
nor U34536 (N_34536,N_33937,N_32324);
and U34537 (N_34537,N_33267,N_33434);
and U34538 (N_34538,N_33246,N_33000);
or U34539 (N_34539,N_33687,N_33451);
or U34540 (N_34540,N_33213,N_33184);
and U34541 (N_34541,N_33410,N_33286);
nor U34542 (N_34542,N_33768,N_33708);
xnor U34543 (N_34543,N_32431,N_33549);
and U34544 (N_34544,N_33025,N_33554);
and U34545 (N_34545,N_32296,N_33559);
nor U34546 (N_34546,N_32237,N_32467);
and U34547 (N_34547,N_32677,N_33328);
xnor U34548 (N_34548,N_33518,N_32871);
nand U34549 (N_34549,N_32436,N_33609);
nand U34550 (N_34550,N_32878,N_32241);
and U34551 (N_34551,N_32569,N_32865);
xnor U34552 (N_34552,N_32278,N_32179);
or U34553 (N_34553,N_32912,N_33063);
and U34554 (N_34554,N_33133,N_33210);
nor U34555 (N_34555,N_32684,N_32468);
or U34556 (N_34556,N_32972,N_33228);
nor U34557 (N_34557,N_33988,N_33234);
or U34558 (N_34558,N_33266,N_32575);
or U34559 (N_34559,N_33343,N_32406);
nand U34560 (N_34560,N_32243,N_32697);
nor U34561 (N_34561,N_33921,N_32163);
nor U34562 (N_34562,N_33024,N_33817);
or U34563 (N_34563,N_33537,N_33255);
xnor U34564 (N_34564,N_32737,N_33658);
or U34565 (N_34565,N_33065,N_32060);
nand U34566 (N_34566,N_32939,N_33534);
and U34567 (N_34567,N_33336,N_32615);
xor U34568 (N_34568,N_32617,N_32736);
and U34569 (N_34569,N_32781,N_33130);
nor U34570 (N_34570,N_32338,N_32641);
or U34571 (N_34571,N_32816,N_32631);
xnor U34572 (N_34572,N_32701,N_33607);
nand U34573 (N_34573,N_33066,N_32447);
nor U34574 (N_34574,N_32205,N_32601);
nand U34575 (N_34575,N_33462,N_33786);
and U34576 (N_34576,N_32099,N_33874);
and U34577 (N_34577,N_33327,N_32102);
and U34578 (N_34578,N_32676,N_32610);
nand U34579 (N_34579,N_32476,N_32389);
and U34580 (N_34580,N_33233,N_33111);
or U34581 (N_34581,N_32653,N_32238);
or U34582 (N_34582,N_33749,N_32643);
or U34583 (N_34583,N_32525,N_33732);
xnor U34584 (N_34584,N_33446,N_33424);
xnor U34585 (N_34585,N_32152,N_32891);
nor U34586 (N_34586,N_32934,N_33398);
or U34587 (N_34587,N_33380,N_32941);
xnor U34588 (N_34588,N_32098,N_33571);
xnor U34589 (N_34589,N_32811,N_32815);
xor U34590 (N_34590,N_33047,N_32634);
nor U34591 (N_34591,N_33516,N_32138);
xnor U34592 (N_34592,N_33717,N_32782);
xor U34593 (N_34593,N_32918,N_33090);
nor U34594 (N_34594,N_32035,N_33765);
xor U34595 (N_34595,N_33037,N_32091);
or U34596 (N_34596,N_32397,N_32466);
nand U34597 (N_34597,N_32720,N_32331);
and U34598 (N_34598,N_32459,N_32435);
xnor U34599 (N_34599,N_32107,N_33562);
and U34600 (N_34600,N_32739,N_32541);
nor U34601 (N_34601,N_33484,N_32512);
nor U34602 (N_34602,N_32052,N_32557);
xnor U34603 (N_34603,N_32953,N_33751);
or U34604 (N_34604,N_32766,N_33418);
nand U34605 (N_34605,N_33743,N_33907);
nor U34606 (N_34606,N_33707,N_32678);
xnor U34607 (N_34607,N_33718,N_33591);
xor U34608 (N_34608,N_32349,N_32858);
nand U34609 (N_34609,N_32173,N_32166);
nand U34610 (N_34610,N_32283,N_33589);
nor U34611 (N_34611,N_32866,N_32101);
nand U34612 (N_34612,N_33816,N_33840);
and U34613 (N_34613,N_32437,N_32213);
nor U34614 (N_34614,N_32620,N_32023);
nand U34615 (N_34615,N_32993,N_33413);
nand U34616 (N_34616,N_32284,N_32800);
or U34617 (N_34617,N_33767,N_32528);
nand U34618 (N_34618,N_32356,N_33308);
and U34619 (N_34619,N_33207,N_32961);
xor U34620 (N_34620,N_32487,N_33860);
xnor U34621 (N_34621,N_32550,N_33625);
xor U34622 (N_34622,N_32627,N_32618);
nand U34623 (N_34623,N_33912,N_33028);
nand U34624 (N_34624,N_32967,N_32510);
nor U34625 (N_34625,N_33555,N_32134);
or U34626 (N_34626,N_32829,N_33546);
nor U34627 (N_34627,N_33784,N_33044);
xor U34628 (N_34628,N_32094,N_33245);
and U34629 (N_34629,N_33720,N_32245);
or U34630 (N_34630,N_32293,N_33381);
nor U34631 (N_34631,N_32458,N_32305);
nor U34632 (N_34632,N_32957,N_32164);
nor U34633 (N_34633,N_33376,N_33795);
nor U34634 (N_34634,N_33900,N_33054);
nor U34635 (N_34635,N_33021,N_32958);
xor U34636 (N_34636,N_32239,N_32507);
nor U34637 (N_34637,N_32088,N_32872);
or U34638 (N_34638,N_32288,N_32328);
xnor U34639 (N_34639,N_32505,N_33372);
xor U34640 (N_34640,N_33914,N_32409);
xnor U34641 (N_34641,N_33365,N_33034);
xnor U34642 (N_34642,N_32079,N_33629);
nand U34643 (N_34643,N_33038,N_33592);
nand U34644 (N_34644,N_32991,N_33062);
or U34645 (N_34645,N_33778,N_33922);
nand U34646 (N_34646,N_33551,N_32572);
xnor U34647 (N_34647,N_33680,N_32067);
or U34648 (N_34648,N_32258,N_32513);
or U34649 (N_34649,N_33970,N_33552);
and U34650 (N_34650,N_33992,N_33677);
xnor U34651 (N_34651,N_32148,N_32644);
and U34652 (N_34652,N_32129,N_33340);
nand U34653 (N_34653,N_32521,N_33842);
nand U34654 (N_34654,N_33830,N_33060);
and U34655 (N_34655,N_33029,N_33106);
or U34656 (N_34656,N_33172,N_33527);
and U34657 (N_34657,N_33584,N_33675);
nand U34658 (N_34658,N_32369,N_32880);
xor U34659 (N_34659,N_33594,N_33933);
or U34660 (N_34660,N_33645,N_32455);
or U34661 (N_34661,N_32686,N_32924);
nand U34662 (N_34662,N_33961,N_32483);
and U34663 (N_34663,N_33804,N_33445);
nand U34664 (N_34664,N_33917,N_32682);
or U34665 (N_34665,N_33580,N_32988);
and U34666 (N_34666,N_32969,N_33496);
nand U34667 (N_34667,N_32425,N_32886);
nor U34668 (N_34668,N_32320,N_32074);
nor U34669 (N_34669,N_32530,N_32879);
nand U34670 (N_34670,N_33428,N_33820);
nor U34671 (N_34671,N_33512,N_32526);
xor U34672 (N_34672,N_32619,N_32375);
nand U34673 (N_34673,N_32807,N_33485);
xnor U34674 (N_34674,N_32626,N_32668);
or U34675 (N_34675,N_33325,N_32463);
or U34676 (N_34676,N_32453,N_33239);
nor U34677 (N_34677,N_32504,N_33853);
and U34678 (N_34678,N_32839,N_33924);
nor U34679 (N_34679,N_33925,N_33288);
or U34680 (N_34680,N_32117,N_32955);
xor U34681 (N_34681,N_32400,N_32938);
xor U34682 (N_34682,N_32662,N_33455);
and U34683 (N_34683,N_32773,N_33606);
xor U34684 (N_34684,N_32488,N_32076);
and U34685 (N_34685,N_32747,N_32986);
xnor U34686 (N_34686,N_32546,N_33271);
or U34687 (N_34687,N_32850,N_32725);
nand U34688 (N_34688,N_32517,N_32225);
or U34689 (N_34689,N_33143,N_32847);
and U34690 (N_34690,N_32987,N_32964);
xor U34691 (N_34691,N_33838,N_33036);
nor U34692 (N_34692,N_33799,N_33222);
and U34693 (N_34693,N_33762,N_32380);
nand U34694 (N_34694,N_33638,N_32995);
or U34695 (N_34695,N_33390,N_33510);
nor U34696 (N_34696,N_32207,N_32749);
xor U34697 (N_34697,N_32856,N_33464);
xnor U34698 (N_34698,N_32265,N_32752);
and U34699 (N_34699,N_33709,N_32156);
or U34700 (N_34700,N_32551,N_32963);
nor U34701 (N_34701,N_33690,N_33304);
xor U34702 (N_34702,N_32311,N_32675);
and U34703 (N_34703,N_32764,N_32274);
or U34704 (N_34704,N_33206,N_33458);
xnor U34705 (N_34705,N_32221,N_32748);
nor U34706 (N_34706,N_32556,N_32629);
xnor U34707 (N_34707,N_32113,N_32545);
nand U34708 (N_34708,N_33163,N_33351);
nor U34709 (N_34709,N_33181,N_32001);
nand U34710 (N_34710,N_33272,N_32754);
or U34711 (N_34711,N_33648,N_32663);
nor U34712 (N_34712,N_32771,N_32892);
xnor U34713 (N_34713,N_32996,N_33042);
nand U34714 (N_34714,N_32037,N_32329);
and U34715 (N_34715,N_33107,N_33032);
and U34716 (N_34716,N_33735,N_33540);
and U34717 (N_34717,N_33742,N_33015);
nor U34718 (N_34718,N_33189,N_33071);
nand U34719 (N_34719,N_33249,N_33536);
xnor U34720 (N_34720,N_33626,N_33952);
and U34721 (N_34721,N_32544,N_32316);
nand U34722 (N_34722,N_33422,N_33307);
xnor U34723 (N_34723,N_33332,N_33971);
and U34724 (N_34724,N_32759,N_33974);
xor U34725 (N_34725,N_33403,N_32031);
xor U34726 (N_34726,N_33407,N_33896);
xor U34727 (N_34727,N_33383,N_33269);
xnor U34728 (N_34728,N_33678,N_33631);
xnor U34729 (N_34729,N_32344,N_32895);
xor U34730 (N_34730,N_33793,N_33397);
xor U34731 (N_34731,N_33892,N_32647);
nand U34732 (N_34732,N_32719,N_33460);
and U34733 (N_34733,N_33409,N_32125);
xnor U34734 (N_34734,N_33634,N_32057);
nor U34735 (N_34735,N_32623,N_32625);
and U34736 (N_34736,N_33178,N_33027);
or U34737 (N_34737,N_32809,N_33354);
or U34738 (N_34738,N_32248,N_32350);
and U34739 (N_34739,N_33419,N_32219);
xnor U34740 (N_34740,N_33098,N_32622);
nor U34741 (N_34741,N_32792,N_32363);
xnor U34742 (N_34742,N_33692,N_33023);
or U34743 (N_34743,N_33805,N_32921);
nor U34744 (N_34744,N_33630,N_32381);
and U34745 (N_34745,N_33432,N_33052);
and U34746 (N_34746,N_33507,N_33087);
xor U34747 (N_34747,N_33059,N_33482);
nor U34748 (N_34748,N_33492,N_33595);
and U34749 (N_34749,N_33827,N_33531);
xnor U34750 (N_34750,N_33741,N_33823);
and U34751 (N_34751,N_32319,N_32549);
or U34752 (N_34752,N_32353,N_33358);
nor U34753 (N_34753,N_33623,N_33254);
or U34754 (N_34754,N_32317,N_32231);
nand U34755 (N_34755,N_32379,N_32645);
nand U34756 (N_34756,N_32884,N_33404);
nand U34757 (N_34757,N_32832,N_33208);
or U34758 (N_34758,N_33349,N_32478);
or U34759 (N_34759,N_33494,N_32923);
or U34760 (N_34760,N_33108,N_32696);
and U34761 (N_34761,N_32449,N_33080);
or U34762 (N_34762,N_32292,N_32058);
and U34763 (N_34763,N_33375,N_33426);
xor U34764 (N_34764,N_33297,N_32269);
xnor U34765 (N_34765,N_32560,N_33906);
or U34766 (N_34766,N_32061,N_32261);
and U34767 (N_34767,N_32167,N_33003);
xor U34768 (N_34768,N_32279,N_33505);
nand U34769 (N_34769,N_32246,N_32867);
nand U34770 (N_34770,N_33292,N_32250);
nand U34771 (N_34771,N_33652,N_33104);
nor U34772 (N_34772,N_32454,N_33314);
xnor U34773 (N_34773,N_33882,N_33203);
xor U34774 (N_34774,N_32493,N_32178);
nand U34775 (N_34775,N_33736,N_32223);
or U34776 (N_34776,N_32702,N_33179);
nor U34777 (N_34777,N_33503,N_33294);
nor U34778 (N_34778,N_32228,N_33597);
nor U34779 (N_34779,N_32778,N_32917);
nor U34780 (N_34780,N_32609,N_32063);
xnor U34781 (N_34781,N_32158,N_32299);
nor U34782 (N_34782,N_32943,N_32854);
nor U34783 (N_34783,N_33477,N_32555);
xor U34784 (N_34784,N_33450,N_33326);
nor U34785 (N_34785,N_33183,N_33543);
or U34786 (N_34786,N_32863,N_32377);
and U34787 (N_34787,N_32322,N_32738);
and U34788 (N_34788,N_32342,N_32734);
xnor U34789 (N_34789,N_32050,N_32717);
or U34790 (N_34790,N_32190,N_33899);
nand U34791 (N_34791,N_32115,N_32646);
xor U34792 (N_34792,N_32382,N_32090);
or U34793 (N_34793,N_33378,N_32019);
and U34794 (N_34794,N_32825,N_32984);
or U34795 (N_34795,N_32059,N_33402);
and U34796 (N_34796,N_32998,N_33815);
and U34797 (N_34797,N_33162,N_32416);
and U34798 (N_34798,N_33429,N_33670);
nand U34799 (N_34799,N_32835,N_32522);
xnor U34800 (N_34800,N_32841,N_32853);
or U34801 (N_34801,N_32126,N_33628);
nand U34802 (N_34802,N_33575,N_32971);
xnor U34803 (N_34803,N_33754,N_32182);
xnor U34804 (N_34804,N_33881,N_33244);
and U34805 (N_34805,N_32751,N_33417);
and U34806 (N_34806,N_32616,N_33068);
nor U34807 (N_34807,N_32032,N_32607);
nand U34808 (N_34808,N_33141,N_32683);
or U34809 (N_34809,N_32593,N_33400);
nor U34810 (N_34810,N_33895,N_33923);
xnor U34811 (N_34811,N_32779,N_33118);
and U34812 (N_34812,N_32903,N_33960);
or U34813 (N_34813,N_32600,N_33731);
or U34814 (N_34814,N_32308,N_33993);
and U34815 (N_34815,N_33169,N_33769);
and U34816 (N_34816,N_33257,N_33603);
xnor U34817 (N_34817,N_33700,N_33517);
nor U34818 (N_34818,N_33033,N_33463);
xnor U34819 (N_34819,N_32297,N_33863);
and U34820 (N_34820,N_32785,N_33067);
nor U34821 (N_34821,N_32005,N_33150);
nand U34822 (N_34822,N_32787,N_33016);
nor U34823 (N_34823,N_32680,N_33433);
nand U34824 (N_34824,N_32077,N_32793);
nor U34825 (N_34825,N_32833,N_32118);
nor U34826 (N_34826,N_32932,N_32906);
or U34827 (N_34827,N_33557,N_32470);
nor U34828 (N_34828,N_32901,N_33204);
nand U34829 (N_34829,N_32398,N_32837);
xnor U34830 (N_34830,N_33602,N_32562);
nor U34831 (N_34831,N_33369,N_33201);
and U34832 (N_34832,N_32335,N_33514);
nor U34833 (N_34833,N_33100,N_32122);
nor U34834 (N_34834,N_33040,N_32000);
nor U34835 (N_34835,N_32450,N_32083);
nand U34836 (N_34836,N_32313,N_33681);
nor U34837 (N_34837,N_32849,N_32203);
xor U34838 (N_34838,N_33318,N_32806);
and U34839 (N_34839,N_33764,N_33959);
nand U34840 (N_34840,N_33473,N_32636);
xnor U34841 (N_34841,N_33298,N_33888);
xor U34842 (N_34842,N_33711,N_32929);
nor U34843 (N_34843,N_33264,N_33832);
xnor U34844 (N_34844,N_33164,N_32614);
and U34845 (N_34845,N_33614,N_33393);
and U34846 (N_34846,N_32204,N_33242);
nor U34847 (N_34847,N_33779,N_32055);
and U34848 (N_34848,N_32947,N_33621);
nor U34849 (N_34849,N_32716,N_33483);
nor U34850 (N_34850,N_33968,N_33663);
nand U34851 (N_34851,N_33867,N_33939);
nand U34852 (N_34852,N_33535,N_32346);
nand U34853 (N_34853,N_32954,N_32907);
nand U34854 (N_34854,N_33289,N_32889);
nand U34855 (N_34855,N_33411,N_33120);
and U34856 (N_34856,N_33978,N_33905);
xor U34857 (N_34857,N_32289,N_32103);
xor U34858 (N_34858,N_32108,N_33539);
and U34859 (N_34859,N_33136,N_32935);
nand U34860 (N_34860,N_32177,N_33055);
nand U34861 (N_34861,N_33466,N_33995);
and U34862 (N_34862,N_32777,N_33362);
nor U34863 (N_34863,N_32347,N_33335);
xor U34864 (N_34864,N_32730,N_32295);
xnor U34865 (N_34865,N_33812,N_32501);
and U34866 (N_34866,N_32928,N_32599);
xor U34867 (N_34867,N_32407,N_32096);
or U34868 (N_34868,N_33856,N_33386);
nor U34869 (N_34869,N_33420,N_33226);
or U34870 (N_34870,N_32890,N_33644);
or U34871 (N_34871,N_32287,N_33008);
nor U34872 (N_34872,N_33890,N_32920);
and U34873 (N_34873,N_32133,N_33088);
or U34874 (N_34874,N_32587,N_33012);
or U34875 (N_34875,N_33148,N_33947);
and U34876 (N_34876,N_33161,N_33836);
nor U34877 (N_34877,N_32185,N_33694);
nand U34878 (N_34878,N_33218,N_32082);
and U34879 (N_34879,N_32535,N_33329);
nor U34880 (N_34880,N_33685,N_32174);
nor U34881 (N_34881,N_33852,N_33293);
nand U34882 (N_34882,N_32303,N_33497);
nand U34883 (N_34883,N_32321,N_32801);
or U34884 (N_34884,N_33302,N_33698);
or U34885 (N_34885,N_33102,N_32999);
or U34886 (N_34886,N_33129,N_32831);
or U34887 (N_34887,N_32949,N_32913);
and U34888 (N_34888,N_32104,N_33942);
nand U34889 (N_34889,N_33826,N_32741);
nand U34890 (N_34890,N_33498,N_33231);
nor U34891 (N_34891,N_32757,N_33285);
or U34892 (N_34892,N_32433,N_33798);
or U34893 (N_34893,N_32006,N_33883);
nor U34894 (N_34894,N_33976,N_32417);
and U34895 (N_34895,N_32218,N_32497);
nand U34896 (N_34896,N_32415,N_33676);
xnor U34897 (N_34897,N_33158,N_33220);
and U34898 (N_34898,N_33232,N_33154);
nor U34899 (N_34899,N_32370,N_32056);
nor U34900 (N_34900,N_33869,N_32275);
nor U34901 (N_34901,N_33478,N_33416);
or U34902 (N_34902,N_33849,N_32183);
and U34903 (N_34903,N_32823,N_32595);
or U34904 (N_34904,N_32570,N_32426);
xnor U34905 (N_34905,N_32965,N_33125);
xnor U34906 (N_34906,N_32272,N_33391);
and U34907 (N_34907,N_32888,N_33363);
or U34908 (N_34908,N_32970,N_32352);
nand U34909 (N_34909,N_33943,N_32364);
or U34910 (N_34910,N_33745,N_32033);
or U34911 (N_34911,N_32410,N_33620);
nand U34912 (N_34912,N_32985,N_32902);
nand U34913 (N_34913,N_32374,N_32086);
xnor U34914 (N_34914,N_32726,N_33908);
or U34915 (N_34915,N_33116,N_33935);
nor U34916 (N_34916,N_32403,N_32116);
and U34917 (N_34917,N_32821,N_32197);
nand U34918 (N_34918,N_33142,N_33916);
and U34919 (N_34919,N_33570,N_33320);
xor U34920 (N_34920,N_32151,N_33260);
nor U34921 (N_34921,N_33075,N_33964);
and U34922 (N_34922,N_33893,N_33058);
nand U34923 (N_34923,N_33331,N_33611);
nand U34924 (N_34924,N_32692,N_33616);
and U34925 (N_34925,N_32951,N_32457);
xnor U34926 (N_34926,N_32558,N_32362);
nand U34927 (N_34927,N_33701,N_32637);
nand U34928 (N_34928,N_33316,N_33337);
xnor U34929 (N_34929,N_33348,N_33001);
or U34930 (N_34930,N_32681,N_32325);
nand U34931 (N_34931,N_32267,N_33703);
xnor U34932 (N_34932,N_32136,N_32820);
xor U34933 (N_34933,N_33958,N_33528);
nand U34934 (N_34934,N_32234,N_32011);
nand U34935 (N_34935,N_32123,N_33371);
nor U34936 (N_34936,N_33835,N_32180);
and U34937 (N_34937,N_32596,N_33377);
nand U34938 (N_34938,N_32012,N_33504);
or U34939 (N_34939,N_32026,N_32724);
xnor U34940 (N_34940,N_33262,N_32007);
or U34941 (N_34941,N_32318,N_33666);
nand U34942 (N_34942,N_32465,N_33506);
xnor U34943 (N_34943,N_32727,N_33931);
nor U34944 (N_34944,N_33324,N_33679);
nor U34945 (N_34945,N_33339,N_33577);
nor U34946 (N_34946,N_33981,N_32176);
nor U34947 (N_34947,N_32509,N_32583);
xnor U34948 (N_34948,N_32490,N_32266);
or U34949 (N_34949,N_32529,N_32332);
or U34950 (N_34950,N_32357,N_33461);
xnor U34951 (N_34951,N_33299,N_33532);
nand U34952 (N_34952,N_33723,N_32502);
or U34953 (N_34953,N_32242,N_33811);
or U34954 (N_34954,N_32671,N_32568);
nand U34955 (N_34955,N_32745,N_33051);
nand U34956 (N_34956,N_32419,N_33695);
and U34957 (N_34957,N_33373,N_32534);
and U34958 (N_34958,N_33004,N_32020);
or U34959 (N_34959,N_32612,N_32462);
xor U34960 (N_34960,N_32669,N_32428);
or U34961 (N_34961,N_33904,N_33929);
nand U34962 (N_34962,N_32919,N_32722);
and U34963 (N_34963,N_33525,N_33814);
or U34964 (N_34964,N_32201,N_33238);
xor U34965 (N_34965,N_33563,N_32881);
nand U34966 (N_34966,N_33306,N_32038);
nand U34967 (N_34967,N_32393,N_32469);
nor U34968 (N_34968,N_33624,N_33126);
and U34969 (N_34969,N_32904,N_32131);
xnor U34970 (N_34970,N_33903,N_33581);
or U34971 (N_34971,N_33780,N_33727);
nand U34972 (N_34972,N_32187,N_32564);
xor U34973 (N_34973,N_33214,N_33846);
xor U34974 (N_34974,N_33657,N_33601);
xor U34975 (N_34975,N_32302,N_32817);
xnor U34976 (N_34976,N_32049,N_32334);
and U34977 (N_34977,N_32566,N_33526);
xnor U34978 (N_34978,N_33017,N_33579);
xor U34979 (N_34979,N_32358,N_32846);
or U34980 (N_34980,N_32756,N_32576);
nor U34981 (N_34981,N_32728,N_33967);
nand U34982 (N_34982,N_33405,N_32769);
and U34983 (N_34983,N_32327,N_33031);
or U34984 (N_34984,N_32708,N_32989);
nand U34985 (N_34985,N_33615,N_33341);
nand U34986 (N_34986,N_33303,N_32189);
and U34987 (N_34987,N_32315,N_32909);
nand U34988 (N_34988,N_33699,N_32155);
and U34989 (N_34989,N_33789,N_33839);
nor U34990 (N_34990,N_32290,N_33453);
xor U34991 (N_34991,N_33456,N_32533);
and U34992 (N_34992,N_32027,N_32765);
nor U34993 (N_34993,N_33662,N_33920);
xnor U34994 (N_34994,N_32552,N_33538);
xnor U34995 (N_34995,N_33599,N_32384);
and U34996 (N_34996,N_33649,N_33149);
nand U34997 (N_34997,N_32440,N_32206);
nand U34998 (N_34998,N_32160,N_32876);
and U34999 (N_34999,N_32882,N_32016);
nor U35000 (N_35000,N_33508,N_32554);
and U35001 (N_35001,N_32970,N_32896);
xor U35002 (N_35002,N_32724,N_33502);
xnor U35003 (N_35003,N_32299,N_32719);
nor U35004 (N_35004,N_32329,N_33442);
or U35005 (N_35005,N_33870,N_33632);
and U35006 (N_35006,N_33725,N_33195);
and U35007 (N_35007,N_32891,N_32912);
or U35008 (N_35008,N_33000,N_33755);
and U35009 (N_35009,N_32562,N_33057);
nor U35010 (N_35010,N_32476,N_32495);
or U35011 (N_35011,N_33011,N_32856);
xor U35012 (N_35012,N_33815,N_32731);
or U35013 (N_35013,N_32186,N_33105);
nor U35014 (N_35014,N_32561,N_32318);
or U35015 (N_35015,N_33840,N_33900);
xor U35016 (N_35016,N_33518,N_33485);
xnor U35017 (N_35017,N_33595,N_32319);
xnor U35018 (N_35018,N_33987,N_33204);
xnor U35019 (N_35019,N_33246,N_33188);
xor U35020 (N_35020,N_33361,N_32774);
and U35021 (N_35021,N_33188,N_32779);
xor U35022 (N_35022,N_32135,N_32377);
and U35023 (N_35023,N_32976,N_32198);
xnor U35024 (N_35024,N_33667,N_32983);
nor U35025 (N_35025,N_33689,N_32594);
nand U35026 (N_35026,N_32916,N_33221);
and U35027 (N_35027,N_33135,N_32079);
nand U35028 (N_35028,N_32152,N_32918);
nor U35029 (N_35029,N_32133,N_33441);
and U35030 (N_35030,N_33961,N_32693);
or U35031 (N_35031,N_32488,N_33822);
or U35032 (N_35032,N_33731,N_33977);
or U35033 (N_35033,N_32212,N_32740);
or U35034 (N_35034,N_33480,N_32182);
nand U35035 (N_35035,N_33613,N_33553);
and U35036 (N_35036,N_33991,N_32578);
or U35037 (N_35037,N_33068,N_32196);
xor U35038 (N_35038,N_32513,N_33078);
nand U35039 (N_35039,N_32455,N_32444);
and U35040 (N_35040,N_32681,N_33339);
xor U35041 (N_35041,N_32492,N_32439);
nor U35042 (N_35042,N_33964,N_33843);
and U35043 (N_35043,N_32969,N_32927);
nand U35044 (N_35044,N_32659,N_33037);
or U35045 (N_35045,N_33800,N_32798);
and U35046 (N_35046,N_33227,N_33265);
or U35047 (N_35047,N_32813,N_32887);
or U35048 (N_35048,N_33428,N_32638);
nor U35049 (N_35049,N_33113,N_32331);
nand U35050 (N_35050,N_32570,N_32291);
or U35051 (N_35051,N_32347,N_33124);
nor U35052 (N_35052,N_33209,N_33533);
nor U35053 (N_35053,N_33261,N_33477);
or U35054 (N_35054,N_33509,N_32373);
and U35055 (N_35055,N_33757,N_32329);
nor U35056 (N_35056,N_32528,N_32753);
and U35057 (N_35057,N_33087,N_33581);
xnor U35058 (N_35058,N_32338,N_33438);
or U35059 (N_35059,N_32884,N_32100);
or U35060 (N_35060,N_33911,N_32344);
nand U35061 (N_35061,N_33388,N_33111);
or U35062 (N_35062,N_32090,N_32071);
nor U35063 (N_35063,N_32704,N_32925);
and U35064 (N_35064,N_32577,N_33045);
or U35065 (N_35065,N_32728,N_32986);
xnor U35066 (N_35066,N_33182,N_33046);
and U35067 (N_35067,N_33312,N_32694);
and U35068 (N_35068,N_32786,N_33092);
nand U35069 (N_35069,N_32042,N_32806);
nand U35070 (N_35070,N_33970,N_33154);
and U35071 (N_35071,N_32623,N_33682);
or U35072 (N_35072,N_33710,N_32183);
nor U35073 (N_35073,N_33846,N_33407);
or U35074 (N_35074,N_33694,N_32109);
nor U35075 (N_35075,N_33269,N_33772);
nor U35076 (N_35076,N_33905,N_32611);
or U35077 (N_35077,N_33659,N_33317);
or U35078 (N_35078,N_32181,N_33354);
xor U35079 (N_35079,N_33028,N_33200);
xor U35080 (N_35080,N_32257,N_32187);
xor U35081 (N_35081,N_32131,N_33106);
nand U35082 (N_35082,N_33657,N_33398);
and U35083 (N_35083,N_32625,N_32557);
and U35084 (N_35084,N_33788,N_33449);
or U35085 (N_35085,N_33727,N_33618);
xnor U35086 (N_35086,N_33978,N_32313);
nand U35087 (N_35087,N_33841,N_32705);
nor U35088 (N_35088,N_32396,N_32492);
or U35089 (N_35089,N_32819,N_32728);
or U35090 (N_35090,N_32798,N_33296);
and U35091 (N_35091,N_33155,N_33362);
or U35092 (N_35092,N_33431,N_33684);
nor U35093 (N_35093,N_32188,N_33130);
xnor U35094 (N_35094,N_32058,N_32353);
nor U35095 (N_35095,N_32340,N_32712);
or U35096 (N_35096,N_33959,N_32536);
or U35097 (N_35097,N_32987,N_33699);
xor U35098 (N_35098,N_33240,N_33438);
nand U35099 (N_35099,N_32108,N_33258);
nand U35100 (N_35100,N_33991,N_33920);
nand U35101 (N_35101,N_32141,N_32325);
and U35102 (N_35102,N_32688,N_33513);
nor U35103 (N_35103,N_32664,N_32370);
or U35104 (N_35104,N_33937,N_33460);
and U35105 (N_35105,N_33966,N_33394);
nand U35106 (N_35106,N_33195,N_32223);
and U35107 (N_35107,N_33905,N_32139);
nor U35108 (N_35108,N_33969,N_32643);
nor U35109 (N_35109,N_32908,N_33676);
xnor U35110 (N_35110,N_32496,N_33859);
or U35111 (N_35111,N_32107,N_32008);
or U35112 (N_35112,N_33672,N_32787);
nand U35113 (N_35113,N_33833,N_32642);
xor U35114 (N_35114,N_32809,N_33484);
xnor U35115 (N_35115,N_33304,N_32315);
or U35116 (N_35116,N_32831,N_32599);
and U35117 (N_35117,N_33394,N_32452);
and U35118 (N_35118,N_33923,N_32177);
or U35119 (N_35119,N_32305,N_32324);
nand U35120 (N_35120,N_32810,N_33920);
nor U35121 (N_35121,N_32116,N_32737);
nand U35122 (N_35122,N_32487,N_33126);
and U35123 (N_35123,N_33068,N_33240);
xor U35124 (N_35124,N_33236,N_33721);
and U35125 (N_35125,N_32540,N_33557);
nor U35126 (N_35126,N_32250,N_32956);
or U35127 (N_35127,N_32047,N_32130);
nor U35128 (N_35128,N_33333,N_33936);
and U35129 (N_35129,N_32427,N_33532);
and U35130 (N_35130,N_33903,N_33409);
nand U35131 (N_35131,N_33532,N_32462);
xnor U35132 (N_35132,N_33594,N_32111);
nor U35133 (N_35133,N_33345,N_32216);
xnor U35134 (N_35134,N_33321,N_33498);
and U35135 (N_35135,N_33943,N_33159);
and U35136 (N_35136,N_33792,N_32196);
nor U35137 (N_35137,N_33336,N_33584);
nand U35138 (N_35138,N_33441,N_33723);
nand U35139 (N_35139,N_33664,N_32296);
xor U35140 (N_35140,N_32410,N_32882);
and U35141 (N_35141,N_33646,N_32554);
xor U35142 (N_35142,N_33419,N_33588);
nand U35143 (N_35143,N_32052,N_33541);
xor U35144 (N_35144,N_32322,N_32165);
xor U35145 (N_35145,N_32911,N_32204);
and U35146 (N_35146,N_32191,N_33887);
nand U35147 (N_35147,N_32410,N_33132);
and U35148 (N_35148,N_32325,N_33604);
and U35149 (N_35149,N_32712,N_33119);
or U35150 (N_35150,N_32024,N_32917);
nor U35151 (N_35151,N_32582,N_32409);
xnor U35152 (N_35152,N_32877,N_33470);
nor U35153 (N_35153,N_33847,N_32269);
nand U35154 (N_35154,N_32664,N_32042);
xor U35155 (N_35155,N_32272,N_33839);
nor U35156 (N_35156,N_33990,N_33775);
nor U35157 (N_35157,N_33546,N_32363);
and U35158 (N_35158,N_33599,N_33305);
and U35159 (N_35159,N_32678,N_32248);
or U35160 (N_35160,N_32652,N_33434);
nor U35161 (N_35161,N_32542,N_32570);
nand U35162 (N_35162,N_33560,N_32705);
and U35163 (N_35163,N_33936,N_32614);
or U35164 (N_35164,N_33528,N_32607);
xor U35165 (N_35165,N_33677,N_32367);
xnor U35166 (N_35166,N_33325,N_32127);
xor U35167 (N_35167,N_33061,N_32264);
nand U35168 (N_35168,N_33933,N_32381);
nand U35169 (N_35169,N_32913,N_33946);
nand U35170 (N_35170,N_32218,N_33151);
or U35171 (N_35171,N_32706,N_32624);
nand U35172 (N_35172,N_32222,N_32552);
nand U35173 (N_35173,N_33397,N_33246);
nor U35174 (N_35174,N_32648,N_33808);
and U35175 (N_35175,N_33731,N_33139);
xor U35176 (N_35176,N_32486,N_33950);
nand U35177 (N_35177,N_32357,N_33834);
xor U35178 (N_35178,N_33562,N_32815);
xor U35179 (N_35179,N_33441,N_32306);
and U35180 (N_35180,N_33265,N_33323);
nor U35181 (N_35181,N_32768,N_32941);
or U35182 (N_35182,N_33955,N_33752);
nand U35183 (N_35183,N_33305,N_32143);
and U35184 (N_35184,N_33421,N_33769);
nand U35185 (N_35185,N_33382,N_33052);
xor U35186 (N_35186,N_32526,N_33658);
or U35187 (N_35187,N_32402,N_32843);
nor U35188 (N_35188,N_33889,N_32007);
and U35189 (N_35189,N_33156,N_33561);
nor U35190 (N_35190,N_32418,N_32479);
and U35191 (N_35191,N_33703,N_32901);
or U35192 (N_35192,N_32402,N_32863);
and U35193 (N_35193,N_33527,N_32232);
and U35194 (N_35194,N_32052,N_32514);
xnor U35195 (N_35195,N_33930,N_33055);
xor U35196 (N_35196,N_32317,N_32336);
and U35197 (N_35197,N_32185,N_32761);
or U35198 (N_35198,N_32424,N_33685);
nor U35199 (N_35199,N_33374,N_32288);
xnor U35200 (N_35200,N_32991,N_33907);
and U35201 (N_35201,N_32399,N_33633);
and U35202 (N_35202,N_32707,N_32219);
or U35203 (N_35203,N_33180,N_33322);
nand U35204 (N_35204,N_32253,N_32512);
and U35205 (N_35205,N_32431,N_33457);
and U35206 (N_35206,N_33657,N_32185);
and U35207 (N_35207,N_32842,N_33873);
nand U35208 (N_35208,N_33293,N_33562);
nand U35209 (N_35209,N_32882,N_32961);
nor U35210 (N_35210,N_33595,N_33974);
nand U35211 (N_35211,N_33601,N_32449);
or U35212 (N_35212,N_32314,N_32476);
and U35213 (N_35213,N_33516,N_33145);
xor U35214 (N_35214,N_32842,N_32526);
nor U35215 (N_35215,N_33023,N_33164);
nor U35216 (N_35216,N_33323,N_33674);
xnor U35217 (N_35217,N_32537,N_33829);
or U35218 (N_35218,N_33003,N_33796);
nand U35219 (N_35219,N_32900,N_32919);
or U35220 (N_35220,N_32085,N_32801);
nor U35221 (N_35221,N_32474,N_33621);
or U35222 (N_35222,N_33304,N_32637);
or U35223 (N_35223,N_33324,N_32226);
or U35224 (N_35224,N_33023,N_33265);
or U35225 (N_35225,N_32217,N_33660);
and U35226 (N_35226,N_32835,N_32277);
or U35227 (N_35227,N_33455,N_33898);
xnor U35228 (N_35228,N_32489,N_33845);
nand U35229 (N_35229,N_33667,N_33797);
and U35230 (N_35230,N_33158,N_33785);
and U35231 (N_35231,N_32320,N_32336);
and U35232 (N_35232,N_33766,N_32459);
nor U35233 (N_35233,N_33885,N_33621);
nand U35234 (N_35234,N_32858,N_32117);
and U35235 (N_35235,N_33784,N_32664);
nand U35236 (N_35236,N_32472,N_33775);
nor U35237 (N_35237,N_32818,N_33427);
or U35238 (N_35238,N_32231,N_33545);
and U35239 (N_35239,N_32119,N_32429);
nor U35240 (N_35240,N_33159,N_33702);
and U35241 (N_35241,N_32783,N_33298);
nor U35242 (N_35242,N_33436,N_33001);
or U35243 (N_35243,N_33862,N_32261);
nand U35244 (N_35244,N_32680,N_32610);
nor U35245 (N_35245,N_33379,N_33429);
xor U35246 (N_35246,N_33820,N_33453);
xor U35247 (N_35247,N_33372,N_33498);
nor U35248 (N_35248,N_33670,N_32823);
and U35249 (N_35249,N_32697,N_33255);
and U35250 (N_35250,N_33221,N_33197);
nand U35251 (N_35251,N_33931,N_33104);
xor U35252 (N_35252,N_32529,N_32565);
nand U35253 (N_35253,N_33099,N_33742);
and U35254 (N_35254,N_33958,N_32322);
nor U35255 (N_35255,N_32623,N_32292);
or U35256 (N_35256,N_32104,N_32666);
nor U35257 (N_35257,N_32984,N_33822);
nand U35258 (N_35258,N_32662,N_33494);
nor U35259 (N_35259,N_33400,N_33510);
xor U35260 (N_35260,N_32315,N_33306);
or U35261 (N_35261,N_32997,N_33613);
xnor U35262 (N_35262,N_33604,N_33762);
and U35263 (N_35263,N_32942,N_33451);
nor U35264 (N_35264,N_32748,N_33957);
nor U35265 (N_35265,N_32753,N_32100);
or U35266 (N_35266,N_32393,N_33093);
or U35267 (N_35267,N_33340,N_33355);
and U35268 (N_35268,N_33701,N_32588);
nand U35269 (N_35269,N_33704,N_33822);
nor U35270 (N_35270,N_32751,N_32120);
or U35271 (N_35271,N_33202,N_32965);
xor U35272 (N_35272,N_33107,N_32409);
and U35273 (N_35273,N_32026,N_33161);
and U35274 (N_35274,N_32085,N_33217);
xor U35275 (N_35275,N_32741,N_33267);
nor U35276 (N_35276,N_32568,N_33272);
or U35277 (N_35277,N_33310,N_33210);
nand U35278 (N_35278,N_32168,N_32933);
or U35279 (N_35279,N_32071,N_33969);
xnor U35280 (N_35280,N_32284,N_32296);
or U35281 (N_35281,N_33487,N_33714);
nor U35282 (N_35282,N_33122,N_33239);
xor U35283 (N_35283,N_33684,N_33589);
nand U35284 (N_35284,N_32689,N_32258);
xnor U35285 (N_35285,N_32541,N_32241);
and U35286 (N_35286,N_33567,N_32679);
nor U35287 (N_35287,N_33852,N_32819);
nand U35288 (N_35288,N_32039,N_33174);
nand U35289 (N_35289,N_33519,N_32774);
nor U35290 (N_35290,N_32340,N_33567);
and U35291 (N_35291,N_32367,N_32373);
nor U35292 (N_35292,N_32467,N_32656);
or U35293 (N_35293,N_32022,N_33300);
nor U35294 (N_35294,N_33575,N_32000);
nand U35295 (N_35295,N_33239,N_32632);
and U35296 (N_35296,N_32871,N_33867);
and U35297 (N_35297,N_32036,N_33081);
nand U35298 (N_35298,N_33851,N_32991);
nand U35299 (N_35299,N_32937,N_33498);
xor U35300 (N_35300,N_32797,N_33472);
nand U35301 (N_35301,N_33711,N_33518);
nor U35302 (N_35302,N_33845,N_33083);
xor U35303 (N_35303,N_33526,N_33254);
and U35304 (N_35304,N_33060,N_32230);
nor U35305 (N_35305,N_32206,N_33137);
and U35306 (N_35306,N_33685,N_32186);
xor U35307 (N_35307,N_32706,N_32941);
or U35308 (N_35308,N_33170,N_32162);
and U35309 (N_35309,N_32507,N_32006);
nor U35310 (N_35310,N_33069,N_32192);
xor U35311 (N_35311,N_32366,N_33953);
xnor U35312 (N_35312,N_32902,N_32833);
or U35313 (N_35313,N_33527,N_33775);
and U35314 (N_35314,N_33183,N_33416);
nor U35315 (N_35315,N_33714,N_32361);
and U35316 (N_35316,N_33321,N_32546);
nor U35317 (N_35317,N_32141,N_32419);
or U35318 (N_35318,N_32815,N_32230);
nand U35319 (N_35319,N_33205,N_33972);
nor U35320 (N_35320,N_32749,N_32952);
nor U35321 (N_35321,N_33717,N_32307);
xnor U35322 (N_35322,N_33847,N_33915);
nor U35323 (N_35323,N_32721,N_32479);
and U35324 (N_35324,N_33760,N_33149);
or U35325 (N_35325,N_33562,N_33721);
nor U35326 (N_35326,N_32465,N_32670);
and U35327 (N_35327,N_32043,N_33506);
xor U35328 (N_35328,N_33128,N_32025);
nor U35329 (N_35329,N_33588,N_33015);
nor U35330 (N_35330,N_32621,N_32683);
nand U35331 (N_35331,N_32712,N_33863);
nand U35332 (N_35332,N_32398,N_33017);
xor U35333 (N_35333,N_33417,N_32220);
or U35334 (N_35334,N_32256,N_32603);
nor U35335 (N_35335,N_33323,N_33277);
and U35336 (N_35336,N_32559,N_32614);
xor U35337 (N_35337,N_32379,N_33806);
xor U35338 (N_35338,N_33349,N_33406);
and U35339 (N_35339,N_32992,N_32106);
xor U35340 (N_35340,N_32794,N_33258);
nor U35341 (N_35341,N_32603,N_33096);
xor U35342 (N_35342,N_33133,N_33853);
and U35343 (N_35343,N_32271,N_33132);
and U35344 (N_35344,N_33189,N_33483);
and U35345 (N_35345,N_33662,N_32736);
nor U35346 (N_35346,N_33280,N_33598);
and U35347 (N_35347,N_32521,N_32365);
nand U35348 (N_35348,N_33427,N_33127);
nand U35349 (N_35349,N_32067,N_33642);
nand U35350 (N_35350,N_33381,N_32491);
or U35351 (N_35351,N_33251,N_32274);
and U35352 (N_35352,N_33031,N_33306);
nor U35353 (N_35353,N_32949,N_32903);
and U35354 (N_35354,N_32369,N_33861);
and U35355 (N_35355,N_32722,N_33634);
nor U35356 (N_35356,N_33130,N_33926);
and U35357 (N_35357,N_33581,N_32803);
nor U35358 (N_35358,N_33514,N_32495);
and U35359 (N_35359,N_33504,N_32668);
and U35360 (N_35360,N_32696,N_32610);
xnor U35361 (N_35361,N_33427,N_32536);
or U35362 (N_35362,N_33876,N_32184);
xor U35363 (N_35363,N_33886,N_33239);
nand U35364 (N_35364,N_32820,N_33227);
nor U35365 (N_35365,N_33341,N_33151);
xor U35366 (N_35366,N_32549,N_33900);
nor U35367 (N_35367,N_33595,N_33039);
or U35368 (N_35368,N_33766,N_33938);
nand U35369 (N_35369,N_32485,N_33178);
xor U35370 (N_35370,N_32746,N_32693);
or U35371 (N_35371,N_32423,N_33469);
xor U35372 (N_35372,N_32671,N_33050);
or U35373 (N_35373,N_33422,N_33598);
nor U35374 (N_35374,N_33493,N_32706);
xor U35375 (N_35375,N_32061,N_32621);
xor U35376 (N_35376,N_32464,N_32434);
and U35377 (N_35377,N_33716,N_33614);
xnor U35378 (N_35378,N_33258,N_33090);
nor U35379 (N_35379,N_33247,N_33304);
nand U35380 (N_35380,N_33856,N_33982);
nor U35381 (N_35381,N_32769,N_32056);
or U35382 (N_35382,N_33528,N_33687);
nand U35383 (N_35383,N_33417,N_33349);
xor U35384 (N_35384,N_33866,N_33871);
nor U35385 (N_35385,N_32689,N_33941);
and U35386 (N_35386,N_33921,N_33001);
xnor U35387 (N_35387,N_33001,N_33452);
nor U35388 (N_35388,N_33202,N_33377);
nor U35389 (N_35389,N_33963,N_33775);
nand U35390 (N_35390,N_32425,N_32221);
and U35391 (N_35391,N_32229,N_33638);
or U35392 (N_35392,N_33978,N_32553);
nor U35393 (N_35393,N_32695,N_33758);
and U35394 (N_35394,N_33128,N_32952);
or U35395 (N_35395,N_33173,N_32232);
xnor U35396 (N_35396,N_32249,N_33194);
nor U35397 (N_35397,N_32190,N_32981);
or U35398 (N_35398,N_33347,N_33490);
xor U35399 (N_35399,N_32257,N_33398);
and U35400 (N_35400,N_32301,N_33093);
nand U35401 (N_35401,N_33596,N_33410);
nand U35402 (N_35402,N_33797,N_32675);
or U35403 (N_35403,N_32342,N_33274);
nor U35404 (N_35404,N_33810,N_32993);
xnor U35405 (N_35405,N_32156,N_33849);
xnor U35406 (N_35406,N_33882,N_32115);
xor U35407 (N_35407,N_33957,N_32278);
and U35408 (N_35408,N_33963,N_33822);
nor U35409 (N_35409,N_33563,N_33147);
xnor U35410 (N_35410,N_32694,N_32640);
and U35411 (N_35411,N_33995,N_32993);
or U35412 (N_35412,N_32366,N_32893);
nand U35413 (N_35413,N_33687,N_32747);
nand U35414 (N_35414,N_33133,N_33036);
xor U35415 (N_35415,N_33411,N_33182);
nor U35416 (N_35416,N_32939,N_32211);
nand U35417 (N_35417,N_32709,N_33062);
xor U35418 (N_35418,N_32797,N_33886);
nand U35419 (N_35419,N_33736,N_33414);
and U35420 (N_35420,N_32794,N_33430);
nand U35421 (N_35421,N_32572,N_32425);
and U35422 (N_35422,N_32360,N_32380);
and U35423 (N_35423,N_32451,N_33582);
and U35424 (N_35424,N_32181,N_32016);
nor U35425 (N_35425,N_32284,N_33759);
xnor U35426 (N_35426,N_32736,N_33334);
nand U35427 (N_35427,N_33782,N_33806);
nor U35428 (N_35428,N_32974,N_32618);
or U35429 (N_35429,N_33189,N_32179);
and U35430 (N_35430,N_33805,N_32992);
or U35431 (N_35431,N_33130,N_33610);
nand U35432 (N_35432,N_33116,N_33314);
nor U35433 (N_35433,N_32177,N_32166);
and U35434 (N_35434,N_32867,N_33607);
nor U35435 (N_35435,N_33902,N_32522);
xor U35436 (N_35436,N_32227,N_33210);
nor U35437 (N_35437,N_33694,N_33579);
nand U35438 (N_35438,N_33071,N_32602);
xnor U35439 (N_35439,N_33779,N_33535);
nand U35440 (N_35440,N_33271,N_32378);
or U35441 (N_35441,N_33113,N_32325);
nor U35442 (N_35442,N_32637,N_33394);
or U35443 (N_35443,N_32509,N_33004);
and U35444 (N_35444,N_32577,N_33778);
xnor U35445 (N_35445,N_32973,N_33621);
nor U35446 (N_35446,N_33530,N_33646);
nor U35447 (N_35447,N_32537,N_32187);
or U35448 (N_35448,N_32801,N_32809);
nor U35449 (N_35449,N_32655,N_33868);
nand U35450 (N_35450,N_32030,N_32552);
nor U35451 (N_35451,N_32901,N_32171);
nand U35452 (N_35452,N_32258,N_32088);
nor U35453 (N_35453,N_32313,N_32616);
xor U35454 (N_35454,N_33145,N_32388);
nor U35455 (N_35455,N_33063,N_33564);
xor U35456 (N_35456,N_33108,N_32865);
or U35457 (N_35457,N_33139,N_33185);
and U35458 (N_35458,N_33919,N_33715);
or U35459 (N_35459,N_33982,N_32757);
xor U35460 (N_35460,N_32356,N_32528);
xnor U35461 (N_35461,N_33139,N_32339);
and U35462 (N_35462,N_33932,N_33910);
nand U35463 (N_35463,N_32162,N_32661);
nand U35464 (N_35464,N_33299,N_32093);
or U35465 (N_35465,N_32651,N_33570);
and U35466 (N_35466,N_33140,N_32287);
xnor U35467 (N_35467,N_32306,N_33204);
nor U35468 (N_35468,N_33168,N_32971);
nand U35469 (N_35469,N_32935,N_33705);
xnor U35470 (N_35470,N_32568,N_32332);
xnor U35471 (N_35471,N_33422,N_33339);
or U35472 (N_35472,N_33893,N_33100);
and U35473 (N_35473,N_33469,N_32987);
or U35474 (N_35474,N_33110,N_33735);
xnor U35475 (N_35475,N_32126,N_33409);
nor U35476 (N_35476,N_33377,N_32969);
or U35477 (N_35477,N_33968,N_33188);
xnor U35478 (N_35478,N_32204,N_33041);
xnor U35479 (N_35479,N_33036,N_33418);
nand U35480 (N_35480,N_32001,N_32274);
nor U35481 (N_35481,N_32833,N_32835);
nand U35482 (N_35482,N_32695,N_32315);
nor U35483 (N_35483,N_32161,N_32609);
and U35484 (N_35484,N_32492,N_33454);
xor U35485 (N_35485,N_33228,N_32176);
nand U35486 (N_35486,N_32455,N_32057);
xor U35487 (N_35487,N_32235,N_33948);
or U35488 (N_35488,N_33348,N_33152);
and U35489 (N_35489,N_33803,N_33761);
nand U35490 (N_35490,N_33195,N_33201);
and U35491 (N_35491,N_33460,N_33481);
or U35492 (N_35492,N_32276,N_32985);
nand U35493 (N_35493,N_32401,N_33264);
nand U35494 (N_35494,N_33698,N_32928);
and U35495 (N_35495,N_32251,N_33417);
nand U35496 (N_35496,N_33252,N_32918);
xnor U35497 (N_35497,N_32386,N_33127);
nor U35498 (N_35498,N_33115,N_33522);
and U35499 (N_35499,N_32639,N_33111);
and U35500 (N_35500,N_32050,N_33157);
xnor U35501 (N_35501,N_33223,N_33198);
xor U35502 (N_35502,N_32507,N_32697);
nor U35503 (N_35503,N_33906,N_32936);
or U35504 (N_35504,N_32971,N_33248);
or U35505 (N_35505,N_33175,N_33267);
and U35506 (N_35506,N_32514,N_32499);
or U35507 (N_35507,N_33260,N_33791);
nand U35508 (N_35508,N_33243,N_33497);
xor U35509 (N_35509,N_33880,N_33445);
and U35510 (N_35510,N_33838,N_33932);
xor U35511 (N_35511,N_33315,N_33669);
xor U35512 (N_35512,N_33756,N_32926);
or U35513 (N_35513,N_33059,N_32221);
xor U35514 (N_35514,N_32062,N_32583);
nand U35515 (N_35515,N_32096,N_32186);
xnor U35516 (N_35516,N_32986,N_32023);
or U35517 (N_35517,N_32857,N_32213);
nor U35518 (N_35518,N_33822,N_33862);
xor U35519 (N_35519,N_32251,N_32353);
and U35520 (N_35520,N_33005,N_32758);
and U35521 (N_35521,N_32767,N_32788);
and U35522 (N_35522,N_33916,N_32491);
xor U35523 (N_35523,N_32317,N_32329);
nand U35524 (N_35524,N_32237,N_33076);
and U35525 (N_35525,N_32429,N_32698);
or U35526 (N_35526,N_33555,N_32484);
or U35527 (N_35527,N_32514,N_32310);
nor U35528 (N_35528,N_33834,N_33544);
and U35529 (N_35529,N_33052,N_33027);
xor U35530 (N_35530,N_32887,N_33600);
and U35531 (N_35531,N_33176,N_32795);
and U35532 (N_35532,N_33227,N_33942);
or U35533 (N_35533,N_32597,N_32967);
and U35534 (N_35534,N_33630,N_32960);
nand U35535 (N_35535,N_33482,N_33460);
nor U35536 (N_35536,N_33694,N_32554);
nand U35537 (N_35537,N_32557,N_32237);
nor U35538 (N_35538,N_32159,N_32173);
and U35539 (N_35539,N_33346,N_32265);
or U35540 (N_35540,N_33959,N_32643);
nor U35541 (N_35541,N_32323,N_32087);
or U35542 (N_35542,N_32254,N_33609);
nor U35543 (N_35543,N_33097,N_33244);
nor U35544 (N_35544,N_32180,N_33559);
and U35545 (N_35545,N_32440,N_32823);
or U35546 (N_35546,N_33537,N_33904);
or U35547 (N_35547,N_33485,N_33534);
nand U35548 (N_35548,N_33329,N_33878);
and U35549 (N_35549,N_33969,N_32658);
xnor U35550 (N_35550,N_33640,N_33369);
nand U35551 (N_35551,N_33675,N_33055);
nor U35552 (N_35552,N_33307,N_33906);
nand U35553 (N_35553,N_32298,N_33339);
xnor U35554 (N_35554,N_32960,N_32917);
or U35555 (N_35555,N_33879,N_33004);
nand U35556 (N_35556,N_32929,N_32455);
nor U35557 (N_35557,N_33011,N_32455);
xor U35558 (N_35558,N_33746,N_32537);
nand U35559 (N_35559,N_32215,N_32235);
xor U35560 (N_35560,N_32018,N_32716);
and U35561 (N_35561,N_32967,N_33098);
or U35562 (N_35562,N_32034,N_32300);
nand U35563 (N_35563,N_33813,N_32836);
and U35564 (N_35564,N_33599,N_33375);
or U35565 (N_35565,N_32161,N_33030);
or U35566 (N_35566,N_33081,N_33773);
nor U35567 (N_35567,N_32691,N_33433);
and U35568 (N_35568,N_33980,N_33408);
nor U35569 (N_35569,N_33211,N_33059);
xnor U35570 (N_35570,N_33679,N_32741);
nand U35571 (N_35571,N_33423,N_32660);
nor U35572 (N_35572,N_33473,N_33302);
nand U35573 (N_35573,N_33749,N_32630);
nand U35574 (N_35574,N_33350,N_32338);
nor U35575 (N_35575,N_33740,N_33285);
nand U35576 (N_35576,N_33628,N_32214);
and U35577 (N_35577,N_33753,N_32365);
and U35578 (N_35578,N_33061,N_32834);
xor U35579 (N_35579,N_32854,N_33363);
nand U35580 (N_35580,N_33774,N_33694);
nand U35581 (N_35581,N_33054,N_33503);
nor U35582 (N_35582,N_33312,N_32797);
nand U35583 (N_35583,N_33732,N_32447);
and U35584 (N_35584,N_32734,N_32073);
nand U35585 (N_35585,N_33063,N_32024);
and U35586 (N_35586,N_33581,N_32550);
nor U35587 (N_35587,N_32761,N_32377);
xnor U35588 (N_35588,N_32876,N_32408);
and U35589 (N_35589,N_33560,N_32869);
and U35590 (N_35590,N_32574,N_33523);
nor U35591 (N_35591,N_32778,N_32002);
or U35592 (N_35592,N_33216,N_32274);
and U35593 (N_35593,N_33784,N_33118);
nor U35594 (N_35594,N_32763,N_32123);
and U35595 (N_35595,N_32789,N_33221);
or U35596 (N_35596,N_32820,N_33123);
nand U35597 (N_35597,N_33768,N_33182);
or U35598 (N_35598,N_32362,N_32726);
nand U35599 (N_35599,N_32111,N_33077);
or U35600 (N_35600,N_32163,N_32865);
or U35601 (N_35601,N_32223,N_33844);
nor U35602 (N_35602,N_32714,N_33047);
nor U35603 (N_35603,N_32250,N_33290);
xnor U35604 (N_35604,N_32104,N_33853);
and U35605 (N_35605,N_33937,N_32996);
xor U35606 (N_35606,N_32049,N_32630);
and U35607 (N_35607,N_32492,N_32648);
and U35608 (N_35608,N_32388,N_33776);
xnor U35609 (N_35609,N_33715,N_33885);
nor U35610 (N_35610,N_32501,N_33616);
xor U35611 (N_35611,N_32833,N_33771);
or U35612 (N_35612,N_33616,N_32173);
nor U35613 (N_35613,N_33740,N_33402);
nor U35614 (N_35614,N_32093,N_33059);
xor U35615 (N_35615,N_32147,N_32252);
nor U35616 (N_35616,N_32670,N_32247);
or U35617 (N_35617,N_33718,N_33904);
nand U35618 (N_35618,N_33128,N_32847);
nor U35619 (N_35619,N_32498,N_33896);
or U35620 (N_35620,N_33682,N_32081);
or U35621 (N_35621,N_33972,N_32581);
or U35622 (N_35622,N_32172,N_32148);
or U35623 (N_35623,N_32131,N_33492);
and U35624 (N_35624,N_32773,N_32333);
nand U35625 (N_35625,N_33890,N_33829);
nor U35626 (N_35626,N_32068,N_32786);
nor U35627 (N_35627,N_33344,N_32024);
and U35628 (N_35628,N_33058,N_33411);
and U35629 (N_35629,N_33023,N_33573);
and U35630 (N_35630,N_33546,N_33104);
nor U35631 (N_35631,N_33814,N_32226);
or U35632 (N_35632,N_33818,N_33932);
xnor U35633 (N_35633,N_33173,N_33354);
or U35634 (N_35634,N_33279,N_33098);
nor U35635 (N_35635,N_33361,N_32224);
nor U35636 (N_35636,N_32190,N_33809);
and U35637 (N_35637,N_32052,N_32793);
nand U35638 (N_35638,N_32496,N_32558);
or U35639 (N_35639,N_33205,N_32857);
xnor U35640 (N_35640,N_32229,N_32996);
or U35641 (N_35641,N_32100,N_32434);
or U35642 (N_35642,N_32603,N_32992);
or U35643 (N_35643,N_33901,N_32105);
or U35644 (N_35644,N_33935,N_33334);
nand U35645 (N_35645,N_33431,N_33686);
nor U35646 (N_35646,N_33484,N_32531);
and U35647 (N_35647,N_33307,N_33135);
nor U35648 (N_35648,N_33832,N_33865);
xor U35649 (N_35649,N_32294,N_32803);
or U35650 (N_35650,N_32756,N_33209);
nand U35651 (N_35651,N_33649,N_33575);
and U35652 (N_35652,N_32728,N_33484);
xor U35653 (N_35653,N_32106,N_33501);
nand U35654 (N_35654,N_33183,N_32920);
nor U35655 (N_35655,N_32462,N_32807);
nand U35656 (N_35656,N_32440,N_33822);
xnor U35657 (N_35657,N_32153,N_33696);
xor U35658 (N_35658,N_33170,N_32733);
nand U35659 (N_35659,N_33717,N_33631);
or U35660 (N_35660,N_33672,N_32311);
nor U35661 (N_35661,N_32565,N_33075);
xor U35662 (N_35662,N_32925,N_32536);
and U35663 (N_35663,N_33906,N_33900);
nor U35664 (N_35664,N_33966,N_33941);
nor U35665 (N_35665,N_32730,N_32419);
or U35666 (N_35666,N_32561,N_33432);
xnor U35667 (N_35667,N_32682,N_33932);
nand U35668 (N_35668,N_32227,N_33672);
nand U35669 (N_35669,N_32121,N_33718);
or U35670 (N_35670,N_32469,N_32787);
xor U35671 (N_35671,N_32993,N_33594);
and U35672 (N_35672,N_33656,N_32978);
and U35673 (N_35673,N_32774,N_33298);
or U35674 (N_35674,N_33654,N_32350);
and U35675 (N_35675,N_33223,N_33638);
xnor U35676 (N_35676,N_32716,N_33468);
and U35677 (N_35677,N_33430,N_32910);
or U35678 (N_35678,N_32773,N_32569);
xor U35679 (N_35679,N_32902,N_33255);
nor U35680 (N_35680,N_33531,N_33063);
nor U35681 (N_35681,N_32306,N_33525);
nor U35682 (N_35682,N_33396,N_33344);
or U35683 (N_35683,N_32432,N_33376);
nor U35684 (N_35684,N_32295,N_32415);
or U35685 (N_35685,N_33381,N_32985);
or U35686 (N_35686,N_32298,N_33436);
nand U35687 (N_35687,N_33073,N_33727);
and U35688 (N_35688,N_32516,N_33476);
and U35689 (N_35689,N_33981,N_32212);
and U35690 (N_35690,N_33858,N_33945);
xnor U35691 (N_35691,N_32888,N_32006);
or U35692 (N_35692,N_33000,N_33571);
nand U35693 (N_35693,N_32608,N_32827);
xnor U35694 (N_35694,N_33430,N_33956);
nand U35695 (N_35695,N_32629,N_32702);
or U35696 (N_35696,N_33287,N_33436);
and U35697 (N_35697,N_33734,N_33633);
xor U35698 (N_35698,N_33426,N_33336);
nand U35699 (N_35699,N_33732,N_33077);
or U35700 (N_35700,N_32245,N_32832);
and U35701 (N_35701,N_32499,N_33981);
and U35702 (N_35702,N_32835,N_33767);
nand U35703 (N_35703,N_33519,N_33781);
xor U35704 (N_35704,N_32395,N_32807);
or U35705 (N_35705,N_32190,N_33867);
xnor U35706 (N_35706,N_32778,N_32201);
or U35707 (N_35707,N_32270,N_32048);
nor U35708 (N_35708,N_33469,N_33959);
nand U35709 (N_35709,N_33194,N_33154);
nand U35710 (N_35710,N_33439,N_32678);
and U35711 (N_35711,N_33466,N_33087);
xnor U35712 (N_35712,N_33754,N_32344);
xnor U35713 (N_35713,N_33404,N_33128);
nor U35714 (N_35714,N_32024,N_33426);
nand U35715 (N_35715,N_32706,N_32028);
nor U35716 (N_35716,N_32477,N_33921);
xor U35717 (N_35717,N_32703,N_33318);
nor U35718 (N_35718,N_33867,N_33602);
or U35719 (N_35719,N_33893,N_33759);
nand U35720 (N_35720,N_32581,N_33356);
nand U35721 (N_35721,N_33382,N_33267);
nor U35722 (N_35722,N_32436,N_33137);
and U35723 (N_35723,N_33682,N_32660);
or U35724 (N_35724,N_32900,N_32314);
nand U35725 (N_35725,N_33511,N_33431);
or U35726 (N_35726,N_32989,N_33002);
nor U35727 (N_35727,N_33192,N_32256);
or U35728 (N_35728,N_33961,N_33272);
or U35729 (N_35729,N_32138,N_33800);
or U35730 (N_35730,N_32882,N_33537);
nand U35731 (N_35731,N_32657,N_33016);
and U35732 (N_35732,N_32766,N_32607);
nand U35733 (N_35733,N_33224,N_32840);
nor U35734 (N_35734,N_33155,N_32813);
nor U35735 (N_35735,N_33529,N_32872);
xnor U35736 (N_35736,N_33587,N_33048);
xnor U35737 (N_35737,N_33371,N_33974);
and U35738 (N_35738,N_33567,N_33170);
and U35739 (N_35739,N_33148,N_33643);
and U35740 (N_35740,N_32189,N_32418);
or U35741 (N_35741,N_32870,N_33026);
nor U35742 (N_35742,N_33987,N_32335);
xor U35743 (N_35743,N_33004,N_33041);
or U35744 (N_35744,N_33720,N_32141);
xor U35745 (N_35745,N_32839,N_33921);
xor U35746 (N_35746,N_32752,N_32071);
or U35747 (N_35747,N_32909,N_33708);
nor U35748 (N_35748,N_33031,N_33565);
and U35749 (N_35749,N_32217,N_32078);
and U35750 (N_35750,N_32906,N_33344);
and U35751 (N_35751,N_32751,N_33580);
nand U35752 (N_35752,N_32258,N_32227);
xnor U35753 (N_35753,N_33158,N_33197);
nor U35754 (N_35754,N_32319,N_32209);
nand U35755 (N_35755,N_33738,N_33175);
and U35756 (N_35756,N_33564,N_33566);
nand U35757 (N_35757,N_33972,N_32346);
or U35758 (N_35758,N_32342,N_33347);
and U35759 (N_35759,N_32515,N_32314);
and U35760 (N_35760,N_33738,N_32882);
xnor U35761 (N_35761,N_32701,N_32270);
nand U35762 (N_35762,N_32430,N_32174);
and U35763 (N_35763,N_33858,N_32903);
nand U35764 (N_35764,N_33646,N_33871);
nor U35765 (N_35765,N_32292,N_32473);
nor U35766 (N_35766,N_33698,N_33589);
nor U35767 (N_35767,N_33203,N_32915);
and U35768 (N_35768,N_33380,N_33745);
or U35769 (N_35769,N_32713,N_33913);
nand U35770 (N_35770,N_32097,N_32876);
xnor U35771 (N_35771,N_32046,N_33381);
and U35772 (N_35772,N_33847,N_32487);
nand U35773 (N_35773,N_33395,N_32014);
xor U35774 (N_35774,N_33519,N_33010);
and U35775 (N_35775,N_32224,N_33993);
nand U35776 (N_35776,N_33939,N_32257);
nor U35777 (N_35777,N_33324,N_32591);
nor U35778 (N_35778,N_32939,N_32212);
nand U35779 (N_35779,N_33926,N_32982);
and U35780 (N_35780,N_32527,N_33679);
nor U35781 (N_35781,N_32118,N_32236);
or U35782 (N_35782,N_33723,N_33199);
nor U35783 (N_35783,N_32084,N_32276);
or U35784 (N_35784,N_33382,N_32102);
and U35785 (N_35785,N_32425,N_32091);
nor U35786 (N_35786,N_32100,N_33360);
nand U35787 (N_35787,N_33729,N_33304);
xnor U35788 (N_35788,N_33584,N_32316);
xor U35789 (N_35789,N_32545,N_32985);
or U35790 (N_35790,N_32598,N_32574);
nand U35791 (N_35791,N_32165,N_32840);
and U35792 (N_35792,N_33660,N_32654);
nand U35793 (N_35793,N_32085,N_32542);
xor U35794 (N_35794,N_33871,N_33960);
xnor U35795 (N_35795,N_33099,N_33326);
nor U35796 (N_35796,N_33777,N_32206);
and U35797 (N_35797,N_32779,N_33189);
xnor U35798 (N_35798,N_32637,N_33534);
or U35799 (N_35799,N_32357,N_32649);
xor U35800 (N_35800,N_33350,N_32065);
or U35801 (N_35801,N_33237,N_32884);
or U35802 (N_35802,N_33755,N_32378);
xor U35803 (N_35803,N_32681,N_33542);
xnor U35804 (N_35804,N_32667,N_33252);
or U35805 (N_35805,N_33638,N_32778);
and U35806 (N_35806,N_33591,N_32228);
and U35807 (N_35807,N_32548,N_33644);
nor U35808 (N_35808,N_32551,N_32225);
and U35809 (N_35809,N_32243,N_33770);
or U35810 (N_35810,N_33795,N_33889);
xnor U35811 (N_35811,N_33524,N_33203);
nand U35812 (N_35812,N_33814,N_32666);
or U35813 (N_35813,N_33902,N_32427);
or U35814 (N_35814,N_33129,N_32432);
xor U35815 (N_35815,N_32577,N_32726);
and U35816 (N_35816,N_33302,N_33931);
and U35817 (N_35817,N_33018,N_32497);
nand U35818 (N_35818,N_32503,N_32913);
or U35819 (N_35819,N_33502,N_32480);
nor U35820 (N_35820,N_33060,N_32046);
nor U35821 (N_35821,N_32369,N_32364);
and U35822 (N_35822,N_32201,N_32591);
or U35823 (N_35823,N_33785,N_33053);
nand U35824 (N_35824,N_33727,N_32050);
and U35825 (N_35825,N_32891,N_32917);
and U35826 (N_35826,N_33628,N_32758);
nor U35827 (N_35827,N_33945,N_33357);
or U35828 (N_35828,N_32563,N_32872);
and U35829 (N_35829,N_32489,N_32422);
and U35830 (N_35830,N_33108,N_33152);
nand U35831 (N_35831,N_32162,N_32742);
nand U35832 (N_35832,N_32849,N_32031);
nand U35833 (N_35833,N_33868,N_32153);
and U35834 (N_35834,N_33717,N_33883);
nor U35835 (N_35835,N_32781,N_33604);
and U35836 (N_35836,N_33026,N_33167);
or U35837 (N_35837,N_33291,N_33159);
nor U35838 (N_35838,N_32738,N_32984);
or U35839 (N_35839,N_32402,N_32882);
nand U35840 (N_35840,N_32546,N_33481);
or U35841 (N_35841,N_32012,N_32714);
nand U35842 (N_35842,N_32705,N_33021);
nor U35843 (N_35843,N_32890,N_32165);
nand U35844 (N_35844,N_33840,N_33107);
nor U35845 (N_35845,N_33505,N_33441);
and U35846 (N_35846,N_32402,N_32436);
or U35847 (N_35847,N_33983,N_32197);
nor U35848 (N_35848,N_32784,N_32044);
and U35849 (N_35849,N_32720,N_32125);
nor U35850 (N_35850,N_33160,N_33294);
and U35851 (N_35851,N_33819,N_33918);
nor U35852 (N_35852,N_32183,N_33698);
xnor U35853 (N_35853,N_32433,N_33236);
and U35854 (N_35854,N_32152,N_33756);
or U35855 (N_35855,N_32246,N_33593);
nor U35856 (N_35856,N_32303,N_32515);
nor U35857 (N_35857,N_32557,N_32390);
and U35858 (N_35858,N_32702,N_32757);
nand U35859 (N_35859,N_32583,N_33929);
xor U35860 (N_35860,N_33896,N_32535);
nand U35861 (N_35861,N_33364,N_33256);
nor U35862 (N_35862,N_32202,N_33604);
xor U35863 (N_35863,N_32437,N_33589);
nand U35864 (N_35864,N_33238,N_32028);
xnor U35865 (N_35865,N_32783,N_33500);
xnor U35866 (N_35866,N_33373,N_32945);
xor U35867 (N_35867,N_33015,N_33281);
or U35868 (N_35868,N_32397,N_32177);
nor U35869 (N_35869,N_32054,N_32071);
and U35870 (N_35870,N_32522,N_33946);
and U35871 (N_35871,N_33351,N_33216);
nor U35872 (N_35872,N_32175,N_32309);
nand U35873 (N_35873,N_33880,N_32297);
or U35874 (N_35874,N_32970,N_32938);
nand U35875 (N_35875,N_32647,N_32106);
xnor U35876 (N_35876,N_33309,N_32860);
and U35877 (N_35877,N_32784,N_33136);
or U35878 (N_35878,N_32038,N_33708);
or U35879 (N_35879,N_33704,N_33652);
and U35880 (N_35880,N_33546,N_33851);
xnor U35881 (N_35881,N_33237,N_32487);
xnor U35882 (N_35882,N_33445,N_33342);
nand U35883 (N_35883,N_32504,N_32302);
xor U35884 (N_35884,N_33795,N_33814);
or U35885 (N_35885,N_33252,N_32610);
or U35886 (N_35886,N_32567,N_32614);
or U35887 (N_35887,N_33644,N_32478);
or U35888 (N_35888,N_32443,N_33486);
and U35889 (N_35889,N_33751,N_32561);
or U35890 (N_35890,N_33547,N_33316);
and U35891 (N_35891,N_32752,N_33694);
or U35892 (N_35892,N_33993,N_33974);
xor U35893 (N_35893,N_32037,N_33885);
or U35894 (N_35894,N_32993,N_32575);
nor U35895 (N_35895,N_33573,N_32565);
xnor U35896 (N_35896,N_32060,N_32903);
nor U35897 (N_35897,N_32112,N_33972);
or U35898 (N_35898,N_32322,N_32640);
and U35899 (N_35899,N_32580,N_33385);
and U35900 (N_35900,N_32538,N_32915);
xnor U35901 (N_35901,N_32770,N_33653);
xor U35902 (N_35902,N_33336,N_32787);
or U35903 (N_35903,N_32001,N_32582);
nor U35904 (N_35904,N_33670,N_33337);
nand U35905 (N_35905,N_32256,N_32719);
and U35906 (N_35906,N_33189,N_33527);
xor U35907 (N_35907,N_33837,N_33078);
and U35908 (N_35908,N_33069,N_33864);
or U35909 (N_35909,N_32084,N_33130);
nand U35910 (N_35910,N_32122,N_32956);
xnor U35911 (N_35911,N_33341,N_32679);
and U35912 (N_35912,N_33633,N_32123);
xor U35913 (N_35913,N_32751,N_33734);
or U35914 (N_35914,N_33309,N_33558);
nor U35915 (N_35915,N_32715,N_33138);
nand U35916 (N_35916,N_33265,N_32097);
nand U35917 (N_35917,N_32511,N_33128);
nand U35918 (N_35918,N_33442,N_32630);
and U35919 (N_35919,N_32352,N_33261);
nor U35920 (N_35920,N_32095,N_33652);
and U35921 (N_35921,N_32637,N_33214);
nor U35922 (N_35922,N_32326,N_32314);
nor U35923 (N_35923,N_32990,N_33129);
nand U35924 (N_35924,N_32446,N_32611);
xnor U35925 (N_35925,N_33803,N_33450);
and U35926 (N_35926,N_33498,N_32393);
and U35927 (N_35927,N_33949,N_32133);
xor U35928 (N_35928,N_33835,N_32816);
or U35929 (N_35929,N_32088,N_33675);
nand U35930 (N_35930,N_33852,N_33667);
nor U35931 (N_35931,N_32894,N_32386);
nand U35932 (N_35932,N_33663,N_32139);
and U35933 (N_35933,N_33786,N_33904);
xor U35934 (N_35934,N_33224,N_33751);
nor U35935 (N_35935,N_32032,N_33164);
xor U35936 (N_35936,N_32936,N_33646);
xnor U35937 (N_35937,N_32112,N_32592);
nor U35938 (N_35938,N_33232,N_33273);
or U35939 (N_35939,N_33477,N_32120);
nor U35940 (N_35940,N_32529,N_32373);
and U35941 (N_35941,N_33625,N_33222);
xor U35942 (N_35942,N_33166,N_33999);
xor U35943 (N_35943,N_33131,N_32477);
and U35944 (N_35944,N_33448,N_32398);
nor U35945 (N_35945,N_33292,N_33516);
nor U35946 (N_35946,N_33463,N_33752);
or U35947 (N_35947,N_32563,N_33164);
and U35948 (N_35948,N_33282,N_32309);
and U35949 (N_35949,N_32045,N_32661);
xnor U35950 (N_35950,N_32499,N_32646);
xor U35951 (N_35951,N_33887,N_32689);
xor U35952 (N_35952,N_32044,N_32279);
and U35953 (N_35953,N_33759,N_33192);
or U35954 (N_35954,N_32011,N_33621);
nor U35955 (N_35955,N_32913,N_32453);
or U35956 (N_35956,N_33242,N_32726);
or U35957 (N_35957,N_33360,N_33754);
xnor U35958 (N_35958,N_32099,N_33031);
nand U35959 (N_35959,N_33106,N_32463);
nor U35960 (N_35960,N_32857,N_33339);
nand U35961 (N_35961,N_33893,N_32887);
nor U35962 (N_35962,N_33759,N_32185);
nor U35963 (N_35963,N_32350,N_32483);
or U35964 (N_35964,N_33525,N_33508);
nand U35965 (N_35965,N_32733,N_33438);
xor U35966 (N_35966,N_32636,N_33129);
or U35967 (N_35967,N_32157,N_33271);
xnor U35968 (N_35968,N_33133,N_32317);
nand U35969 (N_35969,N_32953,N_32222);
and U35970 (N_35970,N_33349,N_33590);
nor U35971 (N_35971,N_32685,N_33467);
or U35972 (N_35972,N_33219,N_33762);
and U35973 (N_35973,N_33975,N_32361);
xor U35974 (N_35974,N_33047,N_33785);
xor U35975 (N_35975,N_33801,N_32537);
nor U35976 (N_35976,N_33174,N_32543);
or U35977 (N_35977,N_33010,N_33074);
or U35978 (N_35978,N_33959,N_32373);
xnor U35979 (N_35979,N_32484,N_33484);
nand U35980 (N_35980,N_32908,N_33749);
or U35981 (N_35981,N_32473,N_33587);
xor U35982 (N_35982,N_33369,N_32022);
nand U35983 (N_35983,N_33600,N_32223);
or U35984 (N_35984,N_32588,N_32059);
and U35985 (N_35985,N_33266,N_33340);
and U35986 (N_35986,N_32601,N_33094);
nand U35987 (N_35987,N_32384,N_32738);
nand U35988 (N_35988,N_32498,N_33597);
or U35989 (N_35989,N_33418,N_32917);
or U35990 (N_35990,N_32446,N_33526);
nor U35991 (N_35991,N_33304,N_33558);
nor U35992 (N_35992,N_32265,N_32753);
nor U35993 (N_35993,N_33875,N_33653);
nor U35994 (N_35994,N_32374,N_33852);
xor U35995 (N_35995,N_33182,N_33063);
xor U35996 (N_35996,N_32165,N_33563);
and U35997 (N_35997,N_32351,N_32772);
nand U35998 (N_35998,N_33997,N_32356);
nand U35999 (N_35999,N_33027,N_33392);
and U36000 (N_36000,N_34506,N_34349);
nor U36001 (N_36001,N_34295,N_34819);
nor U36002 (N_36002,N_35806,N_35557);
and U36003 (N_36003,N_34475,N_34781);
and U36004 (N_36004,N_34529,N_34438);
nand U36005 (N_36005,N_34510,N_34820);
or U36006 (N_36006,N_34296,N_34593);
or U36007 (N_36007,N_35258,N_34472);
nand U36008 (N_36008,N_35254,N_35326);
nor U36009 (N_36009,N_34653,N_34788);
xor U36010 (N_36010,N_34067,N_35956);
or U36011 (N_36011,N_34218,N_34103);
xor U36012 (N_36012,N_35588,N_35859);
and U36013 (N_36013,N_35300,N_34659);
nor U36014 (N_36014,N_34646,N_35202);
xor U36015 (N_36015,N_35069,N_35522);
or U36016 (N_36016,N_35028,N_34992);
and U36017 (N_36017,N_34715,N_34531);
xor U36018 (N_36018,N_35175,N_34070);
xor U36019 (N_36019,N_35286,N_34004);
nand U36020 (N_36020,N_35215,N_35890);
xnor U36021 (N_36021,N_35887,N_34880);
and U36022 (N_36022,N_34031,N_34937);
or U36023 (N_36023,N_35501,N_34487);
or U36024 (N_36024,N_35066,N_34876);
and U36025 (N_36025,N_34246,N_34851);
xnor U36026 (N_36026,N_35304,N_34971);
and U36027 (N_36027,N_35660,N_35907);
xnor U36028 (N_36028,N_35461,N_34194);
and U36029 (N_36029,N_35610,N_34912);
nor U36030 (N_36030,N_34754,N_35064);
xor U36031 (N_36031,N_35969,N_34838);
or U36032 (N_36032,N_34058,N_35166);
or U36033 (N_36033,N_35950,N_35414);
or U36034 (N_36034,N_35460,N_34907);
xnor U36035 (N_36035,N_34027,N_35044);
nand U36036 (N_36036,N_35306,N_34842);
xor U36037 (N_36037,N_34150,N_35569);
xnor U36038 (N_36038,N_35477,N_34508);
and U36039 (N_36039,N_35566,N_35087);
xnor U36040 (N_36040,N_34342,N_34165);
nand U36041 (N_36041,N_35640,N_34595);
and U36042 (N_36042,N_35912,N_34669);
nand U36043 (N_36043,N_34474,N_34827);
or U36044 (N_36044,N_34071,N_35365);
nor U36045 (N_36045,N_35129,N_34704);
nor U36046 (N_36046,N_34227,N_34883);
xor U36047 (N_36047,N_34877,N_35279);
and U36048 (N_36048,N_35251,N_34947);
and U36049 (N_36049,N_34046,N_35035);
and U36050 (N_36050,N_34463,N_35307);
nand U36051 (N_36051,N_35713,N_34364);
xor U36052 (N_36052,N_34893,N_34234);
or U36053 (N_36053,N_35140,N_35707);
nand U36054 (N_36054,N_35464,N_35818);
xor U36055 (N_36055,N_35631,N_35019);
and U36056 (N_36056,N_35778,N_35421);
xnor U36057 (N_36057,N_34513,N_34914);
nand U36058 (N_36058,N_35364,N_35292);
nor U36059 (N_36059,N_35256,N_35895);
nand U36060 (N_36060,N_34901,N_35076);
nor U36061 (N_36061,N_34760,N_35669);
and U36062 (N_36062,N_35596,N_34505);
and U36063 (N_36063,N_35194,N_34677);
xnor U36064 (N_36064,N_34161,N_35149);
nand U36065 (N_36065,N_34414,N_35313);
nand U36066 (N_36066,N_34716,N_35172);
or U36067 (N_36067,N_34634,N_35081);
nor U36068 (N_36068,N_34128,N_34750);
and U36069 (N_36069,N_35828,N_34658);
nor U36070 (N_36070,N_34941,N_34039);
and U36071 (N_36071,N_35975,N_35978);
xor U36072 (N_36072,N_34624,N_35622);
and U36073 (N_36073,N_34331,N_35330);
nor U36074 (N_36074,N_34675,N_34256);
nand U36075 (N_36075,N_34483,N_35368);
nor U36076 (N_36076,N_35687,N_35100);
or U36077 (N_36077,N_35635,N_35556);
and U36078 (N_36078,N_34584,N_34963);
xnor U36079 (N_36079,N_35674,N_34322);
or U36080 (N_36080,N_34352,N_35787);
nand U36081 (N_36081,N_35985,N_34378);
or U36082 (N_36082,N_34823,N_35104);
xnor U36083 (N_36083,N_35416,N_34733);
nor U36084 (N_36084,N_35271,N_34579);
or U36085 (N_36085,N_35219,N_35079);
and U36086 (N_36086,N_34988,N_34664);
and U36087 (N_36087,N_34787,N_35428);
nand U36088 (N_36088,N_34740,N_35725);
or U36089 (N_36089,N_34840,N_35942);
or U36090 (N_36090,N_34396,N_34588);
xor U36091 (N_36091,N_34292,N_35268);
nor U36092 (N_36092,N_35263,N_34010);
nand U36093 (N_36093,N_35020,N_34351);
xor U36094 (N_36094,N_34251,N_35362);
nand U36095 (N_36095,N_35591,N_34905);
and U36096 (N_36096,N_35633,N_34144);
or U36097 (N_36097,N_35496,N_34320);
and U36098 (N_36098,N_35112,N_34069);
nand U36099 (N_36099,N_34359,N_35745);
or U36100 (N_36100,N_35191,N_35555);
xor U36101 (N_36101,N_34940,N_34345);
or U36102 (N_36102,N_35683,N_35170);
nand U36103 (N_36103,N_35957,N_35996);
nor U36104 (N_36104,N_35425,N_35356);
nand U36105 (N_36105,N_34999,N_35351);
nor U36106 (N_36106,N_35614,N_34553);
nand U36107 (N_36107,N_35879,N_34237);
and U36108 (N_36108,N_34863,N_35335);
nand U36109 (N_36109,N_35916,N_35546);
xor U36110 (N_36110,N_34477,N_35308);
and U36111 (N_36111,N_34835,N_34499);
and U36112 (N_36112,N_34620,N_34722);
and U36113 (N_36113,N_35214,N_34942);
and U36114 (N_36114,N_35483,N_35002);
and U36115 (N_36115,N_35370,N_35992);
xnor U36116 (N_36116,N_35734,N_34460);
xnor U36117 (N_36117,N_34416,N_35667);
or U36118 (N_36118,N_35411,N_35708);
nand U36119 (N_36119,N_34393,N_35201);
xor U36120 (N_36120,N_34622,N_35444);
xor U36121 (N_36121,N_35060,N_35539);
nand U36122 (N_36122,N_34362,N_35726);
or U36123 (N_36123,N_35661,N_35662);
nand U36124 (N_36124,N_35590,N_35114);
nor U36125 (N_36125,N_35026,N_34795);
or U36126 (N_36126,N_34891,N_34156);
and U36127 (N_36127,N_34337,N_35116);
and U36128 (N_36128,N_35280,N_34271);
or U36129 (N_36129,N_35663,N_34696);
and U36130 (N_36130,N_35796,N_34129);
xnor U36131 (N_36131,N_35767,N_34864);
nand U36132 (N_36132,N_35310,N_34343);
xnor U36133 (N_36133,N_35835,N_35217);
or U36134 (N_36134,N_34741,N_35653);
nand U36135 (N_36135,N_34803,N_35491);
or U36136 (N_36136,N_34132,N_35827);
nor U36137 (N_36137,N_34488,N_34806);
nor U36138 (N_36138,N_34169,N_35743);
and U36139 (N_36139,N_35868,N_34661);
nor U36140 (N_36140,N_35873,N_34037);
nor U36141 (N_36141,N_34258,N_34617);
xor U36142 (N_36142,N_34307,N_35914);
or U36143 (N_36143,N_34384,N_35502);
nand U36144 (N_36144,N_34968,N_34466);
nand U36145 (N_36145,N_35513,N_35717);
nand U36146 (N_36146,N_34059,N_34752);
nand U36147 (N_36147,N_35180,N_35489);
nand U36148 (N_36148,N_34417,N_35456);
nand U36149 (N_36149,N_34871,N_35131);
xor U36150 (N_36150,N_34253,N_34524);
xor U36151 (N_36151,N_35185,N_34955);
or U36152 (N_36152,N_35010,N_35520);
or U36153 (N_36153,N_35469,N_35070);
or U36154 (N_36154,N_34205,N_34728);
nand U36155 (N_36155,N_35511,N_34420);
xor U36156 (N_36156,N_34509,N_34674);
nand U36157 (N_36157,N_35145,N_35541);
and U36158 (N_36158,N_35382,N_35647);
nor U36159 (N_36159,N_35626,N_35312);
nand U36160 (N_36160,N_35877,N_35809);
or U36161 (N_36161,N_35565,N_35223);
or U36162 (N_36162,N_35999,N_35212);
or U36163 (N_36163,N_35007,N_34742);
nor U36164 (N_36164,N_35107,N_34494);
nand U36165 (N_36165,N_35686,N_35597);
nand U36166 (N_36166,N_35936,N_35244);
nand U36167 (N_36167,N_34166,N_34973);
xnor U36168 (N_36168,N_34764,N_35903);
xnor U36169 (N_36169,N_35001,N_35623);
or U36170 (N_36170,N_34002,N_35467);
and U36171 (N_36171,N_35295,N_34327);
and U36172 (N_36172,N_34257,N_34152);
or U36173 (N_36173,N_35923,N_35492);
or U36174 (N_36174,N_34338,N_34422);
nor U36175 (N_36175,N_34418,N_35536);
and U36176 (N_36176,N_35573,N_35142);
and U36177 (N_36177,N_35053,N_34934);
nand U36178 (N_36178,N_34596,N_35773);
and U36179 (N_36179,N_34878,N_34365);
nand U36180 (N_36180,N_35840,N_35023);
nand U36181 (N_36181,N_34044,N_34757);
and U36182 (N_36182,N_35420,N_34288);
or U36183 (N_36183,N_34172,N_35606);
and U36184 (N_36184,N_34175,N_35514);
or U36185 (N_36185,N_34177,N_34633);
and U36186 (N_36186,N_34998,N_35729);
or U36187 (N_36187,N_35866,N_34151);
xor U36188 (N_36188,N_34939,N_34134);
and U36189 (N_36189,N_35415,N_35457);
and U36190 (N_36190,N_34770,N_34323);
nand U36191 (N_36191,N_34329,N_34511);
nor U36192 (N_36192,N_35432,N_35147);
or U36193 (N_36193,N_34647,N_35911);
nor U36194 (N_36194,N_34133,N_34708);
nand U36195 (N_36195,N_35602,N_35341);
nand U36196 (N_36196,N_35438,N_34316);
and U36197 (N_36197,N_34125,N_34926);
or U36198 (N_36198,N_34832,N_35904);
and U36199 (N_36199,N_34945,N_34665);
and U36200 (N_36200,N_35384,N_34147);
nor U36201 (N_36201,N_35752,N_35406);
xor U36202 (N_36202,N_34294,N_35710);
or U36203 (N_36203,N_34346,N_35052);
or U36204 (N_36204,N_35284,N_34068);
xnor U36205 (N_36205,N_35481,N_34373);
or U36206 (N_36206,N_34461,N_34273);
nand U36207 (N_36207,N_35527,N_34627);
nand U36208 (N_36208,N_34171,N_35898);
nand U36209 (N_36209,N_34552,N_35908);
or U36210 (N_36210,N_34935,N_35848);
xnor U36211 (N_36211,N_34626,N_34569);
nand U36212 (N_36212,N_35419,N_35771);
xnor U36213 (N_36213,N_35274,N_35727);
nand U36214 (N_36214,N_35466,N_34279);
xor U36215 (N_36215,N_35858,N_34435);
xnor U36216 (N_36216,N_34102,N_35151);
or U36217 (N_36217,N_34649,N_35232);
nand U36218 (N_36218,N_34215,N_34314);
nor U36219 (N_36219,N_35870,N_34501);
and U36220 (N_36220,N_34679,N_35600);
nor U36221 (N_36221,N_35652,N_34145);
nor U36222 (N_36222,N_35990,N_34225);
nand U36223 (N_36223,N_35878,N_34113);
nor U36224 (N_36224,N_35148,N_35399);
or U36225 (N_36225,N_34607,N_35862);
xor U36226 (N_36226,N_34604,N_34922);
or U36227 (N_36227,N_35495,N_35762);
and U36228 (N_36228,N_35377,N_34654);
and U36229 (N_36229,N_34810,N_35188);
or U36230 (N_36230,N_35518,N_34812);
xor U36231 (N_36231,N_34481,N_35508);
nor U36232 (N_36232,N_34680,N_35046);
nand U36233 (N_36233,N_34034,N_34382);
nand U36234 (N_36234,N_35599,N_35476);
or U36235 (N_36235,N_35413,N_34784);
nand U36236 (N_36236,N_35789,N_34693);
nand U36237 (N_36237,N_35658,N_35298);
nand U36238 (N_36238,N_34448,N_35974);
or U36239 (N_36239,N_35494,N_34407);
or U36240 (N_36240,N_34413,N_34909);
xnor U36241 (N_36241,N_34022,N_34594);
nor U36242 (N_36242,N_35621,N_35523);
or U36243 (N_36243,N_35031,N_34745);
and U36244 (N_36244,N_34135,N_35794);
or U36245 (N_36245,N_35774,N_35287);
xnor U36246 (N_36246,N_35473,N_35009);
nor U36247 (N_36247,N_34987,N_34038);
and U36248 (N_36248,N_35181,N_34243);
nand U36249 (N_36249,N_34564,N_35487);
or U36250 (N_36250,N_34771,N_34798);
nand U36251 (N_36251,N_34211,N_35689);
nor U36252 (N_36252,N_34141,N_34280);
or U36253 (N_36253,N_35283,N_35792);
or U36254 (N_36254,N_35917,N_34437);
xnor U36255 (N_36255,N_34858,N_35960);
and U36256 (N_36256,N_35799,N_34920);
and U36257 (N_36257,N_35500,N_34906);
and U36258 (N_36258,N_35865,N_34097);
nor U36259 (N_36259,N_35884,N_35861);
xnor U36260 (N_36260,N_35121,N_34259);
nor U36261 (N_36261,N_34032,N_35594);
and U36262 (N_36262,N_35735,N_35378);
nand U36263 (N_36263,N_34539,N_34252);
xor U36264 (N_36264,N_34550,N_35932);
nand U36265 (N_36265,N_35073,N_35839);
or U36266 (N_36266,N_34328,N_34186);
xor U36267 (N_36267,N_35775,N_34179);
or U36268 (N_36268,N_35182,N_34790);
nor U36269 (N_36269,N_34377,N_35324);
and U36270 (N_36270,N_35519,N_35299);
nand U36271 (N_36271,N_34140,N_35478);
or U36272 (N_36272,N_34495,N_35748);
nor U36273 (N_36273,N_35925,N_35234);
and U36274 (N_36274,N_35401,N_35246);
and U36275 (N_36275,N_34719,N_34092);
or U36276 (N_36276,N_35243,N_34219);
nand U36277 (N_36277,N_35127,N_35437);
nor U36278 (N_36278,N_35951,N_34240);
nand U36279 (N_36279,N_35819,N_35721);
xor U36280 (N_36280,N_35552,N_35252);
xor U36281 (N_36281,N_34572,N_34800);
nand U36282 (N_36282,N_34138,N_34326);
nor U36283 (N_36283,N_35442,N_35650);
and U36284 (N_36284,N_35515,N_34869);
or U36285 (N_36285,N_34489,N_35327);
and U36286 (N_36286,N_34542,N_35450);
xor U36287 (N_36287,N_34779,N_35386);
or U36288 (N_36288,N_35165,N_35770);
xnor U36289 (N_36289,N_35963,N_35245);
nor U36290 (N_36290,N_35190,N_35247);
or U36291 (N_36291,N_35269,N_34119);
xnor U36292 (N_36292,N_35682,N_34597);
or U36293 (N_36293,N_34458,N_35688);
or U36294 (N_36294,N_35747,N_34376);
xnor U36295 (N_36295,N_34107,N_34615);
nor U36296 (N_36296,N_34578,N_34056);
and U36297 (N_36297,N_34678,N_34452);
and U36298 (N_36298,N_35183,N_35436);
and U36299 (N_36299,N_34546,N_34302);
or U36300 (N_36300,N_34713,N_34821);
xnor U36301 (N_36301,N_35732,N_35032);
xnor U36302 (N_36302,N_34099,N_35940);
or U36303 (N_36303,N_34555,N_34471);
nor U36304 (N_36304,N_34585,N_35323);
or U36305 (N_36305,N_35915,N_34155);
and U36306 (N_36306,N_35349,N_35115);
or U36307 (N_36307,N_34303,N_34986);
nor U36308 (N_36308,N_34230,N_35654);
nor U36309 (N_36309,N_35159,N_34723);
and U36310 (N_36310,N_34241,N_35352);
or U36311 (N_36311,N_35920,N_34967);
and U36312 (N_36312,N_34662,N_34686);
and U36313 (N_36313,N_34599,N_35355);
xnor U36314 (N_36314,N_34563,N_34982);
xor U36315 (N_36315,N_34720,N_34143);
nor U36316 (N_36316,N_35062,N_35933);
and U36317 (N_36317,N_34231,N_34330);
nor U36318 (N_36318,N_35435,N_34498);
and U36319 (N_36319,N_35959,N_35237);
or U36320 (N_36320,N_34195,N_35656);
xor U36321 (N_36321,N_35037,N_35119);
nand U36322 (N_36322,N_34024,N_35968);
or U36323 (N_36323,N_34568,N_35322);
or U36324 (N_36324,N_34429,N_34379);
nand U36325 (N_36325,N_35550,N_34535);
nand U36326 (N_36326,N_35665,N_35132);
or U36327 (N_36327,N_35843,N_35703);
xnor U36328 (N_36328,N_35091,N_35314);
or U36329 (N_36329,N_34042,N_34347);
and U36330 (N_36330,N_35547,N_34250);
xnor U36331 (N_36331,N_34262,N_35337);
nand U36332 (N_36332,N_35637,N_35369);
or U36333 (N_36333,N_35278,N_35856);
nand U36334 (N_36334,N_34093,N_34671);
xor U36335 (N_36335,N_34110,N_35768);
nor U36336 (N_36336,N_34206,N_34473);
nor U36337 (N_36337,N_35516,N_34375);
or U36338 (N_36338,N_35333,N_34198);
nor U36339 (N_36339,N_35443,N_34029);
nand U36340 (N_36340,N_34682,N_35901);
nand U36341 (N_36341,N_35883,N_35067);
nor U36342 (N_36342,N_35608,N_34792);
and U36343 (N_36343,N_35231,N_35967);
nand U36344 (N_36344,N_34312,N_34888);
nand U36345 (N_36345,N_35178,N_34399);
xor U36346 (N_36346,N_35266,N_35293);
or U36347 (N_36347,N_35184,N_34885);
nand U36348 (N_36348,N_34687,N_35022);
nand U36349 (N_36349,N_34370,N_35636);
and U36350 (N_36350,N_35952,N_35240);
nand U36351 (N_36351,N_34469,N_34805);
and U36352 (N_36352,N_34777,N_34845);
and U36353 (N_36353,N_34561,N_34534);
nand U36354 (N_36354,N_35117,N_35719);
xnor U36355 (N_36355,N_34213,N_34462);
and U36356 (N_36356,N_34242,N_35836);
xor U36357 (N_36357,N_34274,N_35851);
nor U36358 (N_36358,N_35576,N_35504);
and U36359 (N_36359,N_35711,N_35277);
xnor U36360 (N_36360,N_35302,N_34860);
and U36361 (N_36361,N_35801,N_34158);
nand U36362 (N_36362,N_35854,N_34758);
xnor U36363 (N_36363,N_34439,N_35685);
and U36364 (N_36364,N_35612,N_34707);
xnor U36365 (N_36365,N_34176,N_34870);
and U36366 (N_36366,N_35692,N_35065);
or U36367 (N_36367,N_35823,N_34814);
nand U36368 (N_36368,N_34759,N_35678);
and U36369 (N_36369,N_34642,N_34703);
or U36370 (N_36370,N_35003,N_34033);
or U36371 (N_36371,N_35134,N_34459);
or U36372 (N_36372,N_34287,N_34403);
or U36373 (N_36373,N_34008,N_35946);
nand U36374 (N_36374,N_35634,N_34636);
or U36375 (N_36375,N_35200,N_35982);
and U36376 (N_36376,N_35529,N_35888);
xnor U36377 (N_36377,N_35937,N_35397);
xnor U36378 (N_36378,N_34455,N_34515);
nand U36379 (N_36379,N_34577,N_35193);
or U36380 (N_36380,N_35677,N_34358);
and U36381 (N_36381,N_35058,N_34170);
nand U36382 (N_36382,N_35615,N_35482);
and U36383 (N_36383,N_35408,N_35611);
xor U36384 (N_36384,N_34829,N_34167);
xor U36385 (N_36385,N_35000,N_34924);
xor U36386 (N_36386,N_35392,N_34282);
or U36387 (N_36387,N_35761,N_35168);
nor U36388 (N_36388,N_35468,N_35821);
and U36389 (N_36389,N_35276,N_34791);
and U36390 (N_36390,N_34392,N_35681);
xor U36391 (N_36391,N_35849,N_35048);
and U36392 (N_36392,N_34854,N_34265);
nand U36393 (N_36393,N_35831,N_34104);
xnor U36394 (N_36394,N_34690,N_34921);
nor U36395 (N_36395,N_35820,N_35617);
nand U36396 (N_36396,N_35357,N_34804);
xor U36397 (N_36397,N_34434,N_34023);
xnor U36398 (N_36398,N_35570,N_34019);
and U36399 (N_36399,N_35099,N_34065);
nand U36400 (N_36400,N_34964,N_35451);
xor U36401 (N_36401,N_35571,N_34533);
or U36402 (N_36402,N_34268,N_34174);
xor U36403 (N_36403,N_35241,N_35296);
xor U36404 (N_36404,N_34073,N_35361);
nand U36405 (N_36405,N_34224,N_34736);
and U36406 (N_36406,N_35924,N_34576);
xor U36407 (N_36407,N_35403,N_35702);
or U36408 (N_36408,N_35824,N_34238);
and U36409 (N_36409,N_34575,N_35447);
or U36410 (N_36410,N_34521,N_35564);
nand U36411 (N_36411,N_34356,N_35675);
and U36412 (N_36412,N_34762,N_35077);
xor U36413 (N_36413,N_35998,N_35319);
or U36414 (N_36414,N_35128,N_34305);
or U36415 (N_36415,N_34444,N_35479);
nor U36416 (N_36416,N_35781,N_34726);
and U36417 (N_36417,N_35659,N_35387);
nor U36418 (N_36418,N_34867,N_34796);
and U36419 (N_36419,N_34491,N_35753);
nand U36420 (N_36420,N_34184,N_34782);
and U36421 (N_36421,N_34080,N_34486);
and U36422 (N_36422,N_35812,N_34310);
xnor U36423 (N_36423,N_35524,N_34290);
nor U36424 (N_36424,N_35086,N_34833);
xor U36425 (N_36425,N_35459,N_34043);
and U36426 (N_36426,N_35676,N_35122);
nand U36427 (N_36427,N_34443,N_34691);
xor U36428 (N_36428,N_35379,N_35926);
or U36429 (N_36429,N_35376,N_34514);
and U36430 (N_36430,N_35755,N_35016);
and U36431 (N_36431,N_35363,N_34015);
or U36432 (N_36432,N_35949,N_34427);
nand U36433 (N_36433,N_34666,N_34185);
or U36434 (N_36434,N_34711,N_34372);
xnor U36435 (N_36435,N_34793,N_35939);
or U36436 (N_36436,N_35930,N_34297);
xnor U36437 (N_36437,N_34390,N_34397);
and U36438 (N_36438,N_34517,N_35371);
xnor U36439 (N_36439,N_35641,N_35698);
nand U36440 (N_36440,N_34203,N_34724);
xnor U36441 (N_36441,N_35345,N_35561);
and U36442 (N_36442,N_35472,N_35701);
and U36443 (N_36443,N_34126,N_34299);
nand U36444 (N_36444,N_34101,N_34204);
nor U36445 (N_36445,N_35881,N_35716);
or U36446 (N_36446,N_34217,N_35746);
xor U36447 (N_36447,N_35106,N_35381);
xnor U36448 (N_36448,N_35173,N_35720);
xor U36449 (N_36449,N_34276,N_34978);
or U36450 (N_36450,N_34651,N_34807);
and U36451 (N_36451,N_35563,N_35021);
or U36452 (N_36452,N_35706,N_35577);
xor U36453 (N_36453,N_35754,N_35805);
xnor U36454 (N_36454,N_34739,N_35807);
or U36455 (N_36455,N_35410,N_35118);
and U36456 (N_36456,N_34340,N_35815);
and U36457 (N_36457,N_34025,N_34698);
xnor U36458 (N_36458,N_35648,N_35164);
xnor U36459 (N_36459,N_35374,N_35448);
nand U36460 (N_36460,N_34729,N_34368);
xnor U36461 (N_36461,N_34245,N_34743);
or U36462 (N_36462,N_35108,N_34084);
xnor U36463 (N_36463,N_34083,N_34537);
nand U36464 (N_36464,N_34269,N_35742);
nand U36465 (N_36465,N_34528,N_34400);
nor U36466 (N_36466,N_34612,N_35560);
or U36467 (N_36467,N_34774,N_34028);
nand U36468 (N_36468,N_34222,N_35033);
or U36469 (N_36469,N_35979,N_35506);
and U36470 (N_36470,N_35668,N_35691);
nand U36471 (N_36471,N_35125,N_34898);
nand U36472 (N_36472,N_34731,N_35434);
xnor U36473 (N_36473,N_34892,N_34974);
nand U36474 (N_36474,N_35723,N_35919);
and U36475 (N_36475,N_34775,N_34480);
nor U36476 (N_36476,N_35136,N_34753);
or U36477 (N_36477,N_34248,N_35350);
xor U36478 (N_36478,N_35417,N_34301);
and U36479 (N_36479,N_35315,N_35446);
and U36480 (N_36480,N_34394,N_34075);
or U36481 (N_36481,N_35061,N_34193);
nand U36482 (N_36482,N_35343,N_35607);
or U36483 (N_36483,N_35704,N_34717);
or U36484 (N_36484,N_35143,N_35589);
nor U36485 (N_36485,N_34096,N_35535);
nor U36486 (N_36486,N_35584,N_35680);
nor U36487 (N_36487,N_35490,N_35671);
nand U36488 (N_36488,N_35738,N_35900);
or U36489 (N_36489,N_34468,N_34380);
xnor U36490 (N_36490,N_35265,N_34718);
or U36491 (N_36491,N_35737,N_35788);
xor U36492 (N_36492,N_35196,N_34904);
nand U36493 (N_36493,N_35260,N_34862);
nor U36494 (N_36494,N_35339,N_35983);
nor U36495 (N_36495,N_35540,N_34446);
and U36496 (N_36496,N_34751,N_35453);
xor U36497 (N_36497,N_35705,N_35210);
nor U36498 (N_36498,N_34882,N_34601);
xnor U36499 (N_36499,N_34670,N_34079);
nor U36500 (N_36500,N_34115,N_34614);
or U36501 (N_36501,N_35036,N_34591);
nand U36502 (N_36502,N_35038,N_34146);
nand U36503 (N_36503,N_34350,N_34383);
xnor U36504 (N_36504,N_35559,N_34632);
nand U36505 (N_36505,N_34336,N_34843);
or U36506 (N_36506,N_35216,N_34688);
nor U36507 (N_36507,N_35630,N_35015);
xnor U36508 (N_36508,N_34783,N_34062);
nor U36509 (N_36509,N_34284,N_34057);
nand U36510 (N_36510,N_34913,N_35358);
and U36511 (N_36511,N_34405,N_35301);
nand U36512 (N_36512,N_35207,N_35709);
or U36513 (N_36513,N_35288,N_34220);
nand U36514 (N_36514,N_34853,N_35222);
xor U36515 (N_36515,N_34465,N_34908);
or U36516 (N_36516,N_34975,N_34197);
or U36517 (N_36517,N_34061,N_34628);
xnor U36518 (N_36518,N_34005,N_35981);
xnor U36519 (N_36519,N_35543,N_34625);
xor U36520 (N_36520,N_34081,N_35236);
xnor U36521 (N_36521,N_35281,N_35714);
or U36522 (N_36522,N_35034,N_34497);
and U36523 (N_36523,N_35613,N_34324);
nand U36524 (N_36524,N_34540,N_35290);
nor U36525 (N_36525,N_34267,N_34401);
xnor U36526 (N_36526,N_35156,N_35558);
and U36527 (N_36527,N_34500,N_34229);
nor U36528 (N_36528,N_35538,N_35297);
or U36529 (N_36529,N_35578,N_34985);
xnor U36530 (N_36530,N_34266,N_35405);
xor U36531 (N_36531,N_35463,N_35220);
or U36532 (N_36532,N_35736,N_35174);
and U36533 (N_36533,N_34836,N_35808);
xnor U36534 (N_36534,N_35645,N_34849);
nand U36535 (N_36535,N_35897,N_34091);
and U36536 (N_36536,N_34903,N_34421);
or U36537 (N_36537,N_35096,N_35012);
and U36538 (N_36538,N_35601,N_35534);
xnor U36539 (N_36539,N_34077,N_35609);
xnor U36540 (N_36540,N_35587,N_35206);
xnor U36541 (N_36541,N_34589,N_35488);
nor U36542 (N_36542,N_35690,N_34730);
nand U36543 (N_36543,N_35008,N_34482);
or U36544 (N_36544,N_34308,N_34911);
or U36545 (N_36545,N_34001,N_35779);
and U36546 (N_36546,N_34532,N_34549);
nand U36547 (N_36547,N_34012,N_34127);
xnor U36548 (N_36548,N_35605,N_35465);
or U36549 (N_36549,N_35089,N_34746);
nand U36550 (N_36550,N_35162,N_35830);
and U36551 (N_36551,N_34464,N_34333);
nor U36552 (N_36552,N_34051,N_34074);
nor U36553 (N_36553,N_35110,N_35892);
nor U36554 (N_36554,N_34164,N_35651);
or U36555 (N_36555,N_35389,N_34582);
xnor U36556 (N_36556,N_34656,N_34249);
or U36557 (N_36557,N_34890,N_35018);
and U36558 (N_36558,N_35718,N_35454);
nand U36559 (N_36559,N_34335,N_35209);
xnor U36560 (N_36560,N_35935,N_34943);
nor U36561 (N_36561,N_34496,N_34932);
nor U36562 (N_36562,N_34811,N_35869);
nand U36563 (N_36563,N_34440,N_34613);
and U36564 (N_36564,N_35876,N_34424);
xor U36565 (N_36565,N_34641,N_34319);
nor U36566 (N_36566,N_34162,N_35740);
xor U36567 (N_36567,N_34606,N_34078);
and U36568 (N_36568,N_34558,N_35505);
nand U36569 (N_36569,N_35109,N_34652);
xnor U36570 (N_36570,N_35430,N_34063);
nand U36571 (N_36571,N_34602,N_35730);
or U36572 (N_36572,N_35509,N_34306);
nand U36573 (N_36573,N_34961,N_34749);
nand U36574 (N_36574,N_34727,N_35291);
xnor U36575 (N_36575,N_35199,N_35152);
or U36576 (N_36576,N_35530,N_35804);
and U36577 (N_36577,N_35006,N_34936);
xor U36578 (N_36578,N_35537,N_34154);
nor U36579 (N_36579,N_34300,N_34629);
nor U36580 (N_36580,N_35567,N_35239);
nand U36581 (N_36581,N_34334,N_35955);
nand U36582 (N_36582,N_35431,N_34386);
or U36583 (N_36583,N_35013,N_34223);
xnor U36584 (N_36584,N_34712,N_34839);
xnor U36585 (N_36585,N_35989,N_34566);
nor U36586 (N_36586,N_35294,N_34233);
or U36587 (N_36587,N_34928,N_34744);
xnor U36588 (N_36588,N_35728,N_35455);
xor U36589 (N_36589,N_34738,N_34442);
xor U36590 (N_36590,N_34244,N_34014);
nand U36591 (N_36591,N_34859,N_35857);
or U36592 (N_36592,N_35953,N_34173);
nor U36593 (N_36593,N_34600,N_35449);
and U36594 (N_36594,N_34214,N_34423);
or U36595 (N_36595,N_35874,N_35249);
nand U36596 (N_36596,N_35684,N_35972);
nand U36597 (N_36597,N_35984,N_34426);
nand U36598 (N_36598,N_35139,N_34683);
and U36599 (N_36599,N_35072,N_34178);
nand U36600 (N_36600,N_35041,N_35643);
or U36601 (N_36601,N_34105,N_34090);
nand U36602 (N_36602,N_34697,N_35030);
nor U36603 (N_36603,N_34705,N_34021);
nor U36604 (N_36604,N_35604,N_34192);
and U36605 (N_36605,N_34949,N_35427);
and U36606 (N_36606,N_35625,N_34106);
nor U36607 (N_36607,N_35047,N_34554);
xor U36608 (N_36608,N_34122,N_34902);
or U36609 (N_36609,N_35526,N_35439);
and U36610 (N_36610,N_34398,N_35722);
xor U36611 (N_36611,N_35551,N_35964);
nand U36612 (N_36612,N_35944,N_34117);
and U36613 (N_36613,N_34428,N_34959);
nand U36614 (N_36614,N_34447,N_35696);
and U36615 (N_36615,N_34457,N_34492);
nor U36616 (N_36616,N_35750,N_34003);
xor U36617 (N_36617,N_34485,N_34763);
and U36618 (N_36618,N_34756,N_34610);
nor U36619 (N_36619,N_34076,N_34966);
nand U36620 (N_36620,N_34954,N_35791);
xnor U36621 (N_36621,N_35344,N_35120);
xnor U36622 (N_36622,N_34830,N_34374);
nand U36623 (N_36623,N_35407,N_35679);
xor U36624 (N_36624,N_35238,N_35424);
and U36625 (N_36625,N_35385,N_34341);
nor U36626 (N_36626,N_34086,N_35966);
or U36627 (N_36627,N_35712,N_35875);
and U36628 (N_36628,N_35179,N_34694);
and U36629 (N_36629,N_34484,N_35375);
nor U36630 (N_36630,N_35157,N_35189);
xnor U36631 (N_36631,N_34361,N_35948);
xor U36632 (N_36632,N_34035,N_34157);
or U36633 (N_36633,N_34953,N_35993);
or U36634 (N_36634,N_35646,N_35976);
and U36635 (N_36635,N_34958,N_34837);
nand U36636 (N_36636,N_34163,N_35627);
nand U36637 (N_36637,N_35548,N_35257);
xor U36638 (N_36638,N_34984,N_35198);
xor U36639 (N_36639,N_34590,N_34875);
xor U36640 (N_36640,N_34780,N_34737);
and U36641 (N_36641,N_34049,N_34923);
nor U36642 (N_36642,N_35011,N_34586);
and U36643 (N_36643,N_35583,N_35545);
nand U36644 (N_36644,N_35380,N_34765);
and U36645 (N_36645,N_34571,N_35798);
nor U36646 (N_36646,N_34668,N_35739);
nor U36647 (N_36647,N_34523,N_34794);
xor U36648 (N_36648,N_34799,N_35262);
nor U36649 (N_36649,N_34120,N_35057);
nand U36650 (N_36650,N_35941,N_35285);
or U36651 (N_36651,N_34692,N_34285);
nor U36652 (N_36652,N_35340,N_34917);
nor U36653 (N_36653,N_35338,N_34006);
nand U36654 (N_36654,N_34502,N_35097);
and U36655 (N_36655,N_35586,N_34567);
and U36656 (N_36656,N_34277,N_34983);
nand U36657 (N_36657,N_34121,N_34388);
nor U36658 (N_36658,N_34387,N_34815);
xnor U36659 (N_36659,N_35927,N_34470);
nand U36660 (N_36660,N_35383,N_35498);
nand U36661 (N_36661,N_35485,N_35130);
nand U36662 (N_36662,N_35867,N_35225);
xor U36663 (N_36663,N_34445,N_35757);
nand U36664 (N_36664,N_35480,N_35549);
nor U36665 (N_36665,N_34137,N_34275);
or U36666 (N_36666,N_35517,N_34366);
nor U36667 (N_36667,N_34478,N_34676);
xor U36668 (N_36668,N_35029,N_35850);
nor U36669 (N_36669,N_34339,N_35163);
nor U36670 (N_36670,N_35810,N_34456);
nor U36671 (N_36671,N_35970,N_35354);
and U36672 (N_36672,N_34834,N_35205);
or U36673 (N_36673,N_34706,N_35847);
nand U36674 (N_36674,N_35832,N_34619);
and U36675 (N_36675,N_34200,N_34865);
nand U36676 (N_36676,N_34395,N_35056);
nor U36677 (N_36677,N_34111,N_35749);
xor U36678 (N_36678,N_35331,N_35083);
xor U36679 (N_36679,N_34545,N_34520);
nor U36680 (N_36680,N_34994,N_34822);
nor U36681 (N_36681,N_34072,N_35724);
xnor U36682 (N_36682,N_35844,N_35103);
nor U36683 (N_36683,N_35947,N_34541);
nand U36684 (N_36684,N_34415,N_34060);
or U36685 (N_36685,N_35697,N_35782);
nor U36686 (N_36686,N_34512,N_35267);
or U36687 (N_36687,N_35412,N_34100);
nor U36688 (N_36688,N_34897,N_34562);
nor U36689 (N_36689,N_35880,N_35657);
xor U36690 (N_36690,N_35404,N_34289);
or U36691 (N_36691,N_35342,N_34235);
xnor U36692 (N_36692,N_34570,N_34872);
xnor U36693 (N_36693,N_35005,N_34965);
nand U36694 (N_36694,N_34354,N_34709);
nor U36695 (N_36695,N_34467,N_34247);
nor U36696 (N_36696,N_34357,N_35528);
or U36697 (N_36697,N_34451,N_34650);
and U36698 (N_36698,N_35863,N_34332);
and U36699 (N_36699,N_35309,N_35766);
xor U36700 (N_36700,N_35049,N_35853);
nor U36701 (N_36701,N_35226,N_35575);
and U36702 (N_36702,N_35248,N_34976);
and U36703 (N_36703,N_34052,N_34371);
nand U36704 (N_36704,N_34124,N_35088);
nor U36705 (N_36705,N_35320,N_34409);
nor U36706 (N_36706,N_35426,N_35670);
or U36707 (N_36707,N_34644,N_34990);
or U36708 (N_36708,N_34580,N_35039);
and U36709 (N_36709,N_35082,N_35014);
nor U36710 (N_36710,N_35388,N_35790);
or U36711 (N_36711,N_35141,N_34261);
or U36712 (N_36712,N_35272,N_34592);
or U36713 (N_36713,N_35797,N_35693);
nand U36714 (N_36714,N_35554,N_34824);
and U36715 (N_36715,N_35632,N_34281);
xnor U36716 (N_36716,N_34522,N_35177);
nand U36717 (N_36717,N_34808,N_34321);
or U36718 (N_36718,N_34209,N_35255);
nor U36719 (N_36719,N_34311,N_34479);
nand U36720 (N_36720,N_35332,N_34672);
nor U36721 (N_36721,N_34681,N_34408);
nor U36722 (N_36722,N_35084,N_34916);
and U36723 (N_36723,N_35593,N_35017);
nand U36724 (N_36724,N_34476,N_34977);
nand U36725 (N_36725,N_35872,N_34996);
or U36726 (N_36726,N_34710,N_35213);
xor U36727 (N_36727,N_35655,N_34436);
and U36728 (N_36728,N_35176,N_35988);
or U36729 (N_36729,N_34773,N_35580);
or U36730 (N_36730,N_34972,N_34797);
nor U36731 (N_36731,N_35433,N_34236);
and U36732 (N_36732,N_35160,N_35101);
or U36733 (N_36733,N_34673,N_34264);
or U36734 (N_36734,N_35074,N_35846);
xnor U36735 (N_36735,N_34896,N_35329);
nand U36736 (N_36736,N_35359,N_35235);
nor U36737 (N_36737,N_34637,N_34449);
xnor U36738 (N_36738,N_35510,N_35154);
or U36739 (N_36739,N_35167,N_34685);
xor U36740 (N_36740,N_34786,N_34118);
nor U36741 (N_36741,N_34816,N_34689);
xnor U36742 (N_36742,N_34293,N_34817);
nor U36743 (N_36743,N_35093,N_34938);
and U36744 (N_36744,N_35211,N_35921);
nor U36745 (N_36745,N_35758,N_35553);
nand U36746 (N_36746,N_35772,N_35574);
or U36747 (N_36747,N_34565,N_34657);
or U36748 (N_36748,N_34648,N_34263);
nor U36749 (N_36749,N_34385,N_35751);
xnor U36750 (N_36750,N_35224,N_35973);
xor U36751 (N_36751,N_34768,N_34210);
and U36752 (N_36752,N_35885,N_34254);
or U36753 (N_36753,N_35962,N_35860);
nand U36754 (N_36754,N_34139,N_34556);
nand U36755 (N_36755,N_35864,N_35644);
nor U36756 (N_36756,N_34066,N_35579);
or U36757 (N_36757,N_34410,N_35228);
nand U36758 (N_36758,N_35144,N_35051);
nand U36759 (N_36759,N_35731,N_34755);
nor U36760 (N_36760,N_35639,N_35891);
xor U36761 (N_36761,N_35282,N_34732);
xor U36762 (N_36762,N_34813,N_35043);
xnor U36763 (N_36763,N_34899,N_35229);
nand U36764 (N_36764,N_34270,N_35913);
and U36765 (N_36765,N_34884,N_35394);
xnor U36766 (N_36766,N_34818,N_35793);
or U36767 (N_36767,N_35155,N_34412);
and U36768 (N_36768,N_34411,N_35841);
and U36769 (N_36769,N_35786,N_35264);
nor U36770 (N_36770,N_35780,N_35253);
xor U36771 (N_36771,N_34000,N_34583);
or U36772 (N_36772,N_35195,N_34894);
and U36773 (N_36773,N_34702,N_34639);
nand U36774 (N_36774,N_35186,N_35261);
and U36775 (N_36775,N_34149,N_35592);
or U36776 (N_36776,N_35521,N_34979);
xnor U36777 (N_36777,N_35045,N_35318);
and U36778 (N_36778,N_35400,N_35095);
or U36779 (N_36779,N_34761,N_35497);
and U36780 (N_36780,N_34188,N_34183);
nor U36781 (N_36781,N_34587,N_34663);
or U36782 (N_36782,N_35833,N_35699);
or U36783 (N_36783,N_34844,N_35486);
nand U36784 (N_36784,N_35525,N_34048);
or U36785 (N_36785,N_34608,N_35133);
nor U36786 (N_36786,N_34232,N_34970);
nor U36787 (N_36787,N_34087,N_35227);
xor U36788 (N_36788,N_35954,N_35664);
nand U36789 (N_36789,N_34355,N_35889);
or U36790 (N_36790,N_34433,N_34918);
nor U36791 (N_36791,N_34291,N_35042);
or U36792 (N_36792,N_35871,N_34946);
xnor U36793 (N_36793,N_34547,N_34950);
xor U36794 (N_36794,N_34026,N_34283);
and U36795 (N_36795,N_34725,N_34381);
xnor U36796 (N_36796,N_35906,N_35094);
and U36797 (N_36797,N_34852,N_34573);
and U36798 (N_36798,N_35233,N_35259);
and U36799 (N_36799,N_35816,N_34182);
nand U36800 (N_36800,N_35931,N_34603);
and U36801 (N_36801,N_34189,N_34956);
nand U36802 (N_36802,N_35102,N_34766);
and U36803 (N_36803,N_35242,N_34700);
or U36804 (N_36804,N_34868,N_35756);
or U36805 (N_36805,N_34286,N_35393);
nor U36806 (N_36806,N_34112,N_34450);
nor U36807 (N_36807,N_35137,N_34551);
nor U36808 (N_36808,N_35852,N_34013);
nor U36809 (N_36809,N_35054,N_35899);
nor U36810 (N_36810,N_34778,N_34895);
nor U36811 (N_36811,N_34116,N_35055);
nand U36812 (N_36812,N_35273,N_35071);
xnor U36813 (N_36813,N_34298,N_35111);
or U36814 (N_36814,N_34402,N_35347);
nand U36815 (N_36815,N_35171,N_34313);
and U36816 (N_36816,N_34317,N_34925);
or U36817 (N_36817,N_35402,N_35997);
nand U36818 (N_36818,N_34425,N_34047);
xor U36819 (N_36819,N_34009,N_34856);
nor U36820 (N_36820,N_35040,N_34207);
or U36821 (N_36821,N_34148,N_35321);
and U36822 (N_36822,N_35694,N_34007);
nor U36823 (N_36823,N_35744,N_34353);
and U36824 (N_36824,N_35784,N_34933);
nor U36825 (N_36825,N_35080,N_35367);
nor U36826 (N_36826,N_34881,N_35126);
xnor U36827 (N_36827,N_34948,N_34507);
or U36828 (N_36828,N_34088,N_34640);
and U36829 (N_36829,N_35568,N_34050);
or U36830 (N_36830,N_34850,N_34855);
or U36831 (N_36831,N_35581,N_34559);
and U36832 (N_36832,N_35741,N_35918);
or U36833 (N_36833,N_34929,N_34041);
nand U36834 (N_36834,N_34887,N_35763);
and U36835 (N_36835,N_35471,N_34981);
nand U36836 (N_36836,N_35624,N_35063);
or U36837 (N_36837,N_35991,N_35759);
and U36838 (N_36838,N_35390,N_35348);
nand U36839 (N_36839,N_35507,N_34931);
and U36840 (N_36840,N_35275,N_35123);
or U36841 (N_36841,N_35218,N_34369);
nand U36842 (N_36842,N_34159,N_35618);
nor U36843 (N_36843,N_34082,N_34598);
nor U36844 (N_36844,N_35938,N_34526);
nor U36845 (N_36845,N_35896,N_34304);
and U36846 (N_36846,N_35795,N_35813);
nand U36847 (N_36847,N_34574,N_35025);
nand U36848 (N_36848,N_35462,N_34825);
or U36849 (N_36849,N_35429,N_34089);
xor U36850 (N_36850,N_34504,N_34618);
and U36851 (N_36851,N_35986,N_34997);
nand U36852 (N_36852,N_34201,N_34538);
and U36853 (N_36853,N_34454,N_35532);
xor U36854 (N_36854,N_34910,N_35595);
xor U36855 (N_36855,N_35672,N_35642);
xor U36856 (N_36856,N_34018,N_35398);
xnor U36857 (N_36857,N_35811,N_35585);
or U36858 (N_36858,N_35373,N_34831);
and U36859 (N_36859,N_35250,N_34993);
nand U36860 (N_36860,N_35153,N_34776);
nor U36861 (N_36861,N_34879,N_34040);
nor U36862 (N_36862,N_34847,N_35499);
and U36863 (N_36863,N_34490,N_34196);
nor U36864 (N_36864,N_35475,N_34181);
or U36865 (N_36865,N_35582,N_34969);
xor U36866 (N_36866,N_35270,N_35837);
xnor U36867 (N_36867,N_34623,N_35158);
xor U36868 (N_36868,N_34951,N_34202);
nor U36869 (N_36869,N_34216,N_34927);
nand U36870 (N_36870,N_34094,N_34536);
xor U36871 (N_36871,N_34389,N_35328);
nand U36872 (N_36872,N_34153,N_34525);
or U36873 (N_36873,N_34191,N_34180);
and U36874 (N_36874,N_35075,N_34208);
xnor U36875 (N_36875,N_35777,N_35336);
nor U36876 (N_36876,N_34826,N_34095);
nand U36877 (N_36877,N_35146,N_34432);
or U36878 (N_36878,N_35638,N_35396);
or U36879 (N_36879,N_35203,N_34857);
nor U36880 (N_36880,N_34212,N_35544);
or U36881 (N_36881,N_35395,N_35418);
and U36882 (N_36882,N_35882,N_34036);
or U36883 (N_36883,N_34085,N_34142);
xor U36884 (N_36884,N_34503,N_35620);
xnor U36885 (N_36885,N_34874,N_35817);
xor U36886 (N_36886,N_35204,N_35715);
or U36887 (N_36887,N_35221,N_34714);
nor U36888 (N_36888,N_34991,N_35169);
xnor U36889 (N_36889,N_35649,N_34020);
nand U36890 (N_36890,N_34846,N_35945);
nor U36891 (N_36891,N_35629,N_34919);
or U36892 (N_36892,N_35325,N_34699);
nor U36893 (N_36893,N_34609,N_35783);
or U36894 (N_36894,N_35829,N_35493);
or U36895 (N_36895,N_35838,N_35289);
nor U36896 (N_36896,N_34054,N_35943);
nor U36897 (N_36897,N_35922,N_35800);
and U36898 (N_36898,N_34631,N_34168);
nand U36899 (N_36899,N_35700,N_35971);
xnor U36900 (N_36900,N_34360,N_35977);
nand U36901 (N_36901,N_35098,N_34900);
nand U36902 (N_36902,N_34123,N_34789);
nand U36903 (N_36903,N_35995,N_34391);
nor U36904 (N_36904,N_35562,N_34030);
and U36905 (N_36905,N_35902,N_35090);
xnor U36906 (N_36906,N_35187,N_34543);
and U36907 (N_36907,N_35422,N_35105);
nand U36908 (N_36908,N_34557,N_35910);
nand U36909 (N_36909,N_35334,N_34785);
and U36910 (N_36910,N_34309,N_34944);
nor U36911 (N_36911,N_35484,N_35826);
nand U36912 (N_36912,N_34995,N_34581);
xnor U36913 (N_36913,N_34767,N_34419);
or U36914 (N_36914,N_35894,N_35024);
xnor U36915 (N_36915,N_34011,N_34930);
and U36916 (N_36916,N_34548,N_35027);
nor U36917 (N_36917,N_34493,N_34406);
xnor U36918 (N_36918,N_34348,N_34114);
xnor U36919 (N_36919,N_35842,N_34131);
nor U36920 (N_36920,N_34430,N_35845);
nor U36921 (N_36921,N_34516,N_34630);
or U36922 (N_36922,N_35317,N_34660);
nand U36923 (N_36923,N_34221,N_35572);
nand U36924 (N_36924,N_35980,N_35834);
nor U36925 (N_36925,N_35470,N_35208);
xnor U36926 (N_36926,N_34404,N_34643);
and U36927 (N_36927,N_34228,N_34016);
or U36928 (N_36928,N_34621,N_34199);
nand U36929 (N_36929,N_34053,N_34136);
xnor U36930 (N_36930,N_34873,N_35078);
and U36931 (N_36931,N_34667,N_34915);
and U36932 (N_36932,N_35150,N_34721);
or U36933 (N_36933,N_34453,N_34747);
and U36934 (N_36934,N_34989,N_34017);
nand U36935 (N_36935,N_34769,N_35987);
or U36936 (N_36936,N_35113,N_34748);
and U36937 (N_36937,N_35628,N_35353);
xor U36938 (N_36938,N_35050,N_35958);
and U36939 (N_36939,N_34441,N_35138);
or U36940 (N_36940,N_34801,N_34638);
or U36941 (N_36941,N_35372,N_34734);
nand U36942 (N_36942,N_35825,N_35474);
or U36943 (N_36943,N_34560,N_35161);
nor U36944 (N_36944,N_35802,N_35909);
and U36945 (N_36945,N_34160,N_34848);
and U36946 (N_36946,N_35458,N_35068);
nand U36947 (N_36947,N_35760,N_34735);
xor U36948 (N_36948,N_34109,N_34611);
nor U36949 (N_36949,N_34344,N_34645);
and U36950 (N_36950,N_35765,N_35961);
nand U36951 (N_36951,N_34325,N_34272);
nor U36952 (N_36952,N_35619,N_35440);
and U36953 (N_36953,N_35542,N_35135);
xnor U36954 (N_36954,N_34315,N_35822);
xnor U36955 (N_36955,N_34957,N_35603);
xor U36956 (N_36956,N_35305,N_34045);
xnor U36957 (N_36957,N_34544,N_34886);
nor U36958 (N_36958,N_35905,N_35531);
xnor U36959 (N_36959,N_35441,N_34828);
and U36960 (N_36960,N_35666,N_35503);
nand U36961 (N_36961,N_35673,N_35192);
and U36962 (N_36962,N_35769,N_35965);
nor U36963 (N_36963,N_35886,N_34802);
nand U36964 (N_36964,N_34055,N_35445);
xor U36965 (N_36965,N_35928,N_35803);
and U36966 (N_36966,N_35085,N_34363);
xnor U36967 (N_36967,N_34519,N_34684);
nand U36968 (N_36968,N_34260,N_35391);
xnor U36969 (N_36969,N_35814,N_34064);
xnor U36970 (N_36970,N_34655,N_34226);
and U36971 (N_36971,N_35855,N_34527);
and U36972 (N_36972,N_34367,N_34701);
nand U36973 (N_36973,N_34605,N_35197);
xnor U36974 (N_36974,N_35004,N_34278);
and U36975 (N_36975,N_34861,N_34530);
nand U36976 (N_36976,N_34098,N_34952);
nand U36977 (N_36977,N_34809,N_35366);
nand U36978 (N_36978,N_35360,N_34960);
xor U36979 (N_36979,N_35346,N_35092);
nand U36980 (N_36980,N_34187,N_35934);
and U36981 (N_36981,N_34889,N_35785);
and U36982 (N_36982,N_34635,N_34962);
nand U36983 (N_36983,N_35695,N_35230);
xnor U36984 (N_36984,N_34190,N_35929);
and U36985 (N_36985,N_35598,N_34239);
nand U36986 (N_36986,N_35423,N_34318);
and U36987 (N_36987,N_35124,N_35311);
nor U36988 (N_36988,N_34255,N_35409);
nand U36989 (N_36989,N_35059,N_35893);
xnor U36990 (N_36990,N_35776,N_34616);
nor U36991 (N_36991,N_34108,N_34841);
nand U36992 (N_36992,N_35616,N_35316);
nor U36993 (N_36993,N_34695,N_34130);
and U36994 (N_36994,N_34772,N_35452);
nor U36995 (N_36995,N_34431,N_34980);
xnor U36996 (N_36996,N_35303,N_35994);
or U36997 (N_36997,N_35512,N_35733);
or U36998 (N_36998,N_35533,N_34866);
or U36999 (N_36999,N_35764,N_34518);
xnor U37000 (N_37000,N_35899,N_34155);
nand U37001 (N_37001,N_35582,N_34654);
xor U37002 (N_37002,N_35302,N_34264);
nand U37003 (N_37003,N_35302,N_34622);
xor U37004 (N_37004,N_34290,N_34276);
and U37005 (N_37005,N_35623,N_35455);
nand U37006 (N_37006,N_34084,N_34501);
nand U37007 (N_37007,N_34777,N_35904);
and U37008 (N_37008,N_34990,N_35403);
or U37009 (N_37009,N_34682,N_34367);
and U37010 (N_37010,N_34019,N_35825);
nand U37011 (N_37011,N_34037,N_35798);
nand U37012 (N_37012,N_34057,N_35512);
nor U37013 (N_37013,N_35444,N_34441);
or U37014 (N_37014,N_34408,N_34671);
and U37015 (N_37015,N_35549,N_34290);
xor U37016 (N_37016,N_34273,N_35767);
and U37017 (N_37017,N_34942,N_34798);
nor U37018 (N_37018,N_34374,N_34920);
or U37019 (N_37019,N_34523,N_35118);
nor U37020 (N_37020,N_34646,N_35617);
nor U37021 (N_37021,N_34085,N_35355);
xor U37022 (N_37022,N_35778,N_34576);
xor U37023 (N_37023,N_35700,N_35332);
and U37024 (N_37024,N_35859,N_35560);
nor U37025 (N_37025,N_35434,N_34285);
xnor U37026 (N_37026,N_34555,N_34047);
or U37027 (N_37027,N_35761,N_34849);
or U37028 (N_37028,N_34735,N_35097);
xnor U37029 (N_37029,N_34807,N_34957);
and U37030 (N_37030,N_35715,N_34071);
or U37031 (N_37031,N_35256,N_34371);
or U37032 (N_37032,N_34714,N_35107);
or U37033 (N_37033,N_34189,N_34330);
nor U37034 (N_37034,N_34358,N_35514);
xor U37035 (N_37035,N_34193,N_35983);
or U37036 (N_37036,N_34788,N_35427);
nand U37037 (N_37037,N_35637,N_35450);
nand U37038 (N_37038,N_34105,N_34366);
nand U37039 (N_37039,N_34720,N_34911);
or U37040 (N_37040,N_35388,N_34952);
and U37041 (N_37041,N_35418,N_34050);
nand U37042 (N_37042,N_34545,N_35036);
xnor U37043 (N_37043,N_34855,N_34268);
xnor U37044 (N_37044,N_34686,N_34941);
xor U37045 (N_37045,N_34631,N_34767);
nor U37046 (N_37046,N_35890,N_35268);
nand U37047 (N_37047,N_34873,N_34413);
or U37048 (N_37048,N_35204,N_34426);
or U37049 (N_37049,N_34354,N_35079);
xor U37050 (N_37050,N_34973,N_35965);
or U37051 (N_37051,N_34360,N_35732);
nor U37052 (N_37052,N_34013,N_35862);
and U37053 (N_37053,N_35099,N_35084);
and U37054 (N_37054,N_34364,N_35143);
or U37055 (N_37055,N_34902,N_34909);
and U37056 (N_37056,N_34398,N_34240);
and U37057 (N_37057,N_34562,N_34641);
nand U37058 (N_37058,N_35850,N_34481);
xor U37059 (N_37059,N_34597,N_34114);
nand U37060 (N_37060,N_34020,N_35191);
nand U37061 (N_37061,N_34221,N_34399);
or U37062 (N_37062,N_34819,N_34440);
and U37063 (N_37063,N_35333,N_35119);
xor U37064 (N_37064,N_34955,N_35911);
and U37065 (N_37065,N_34254,N_34125);
nand U37066 (N_37066,N_35623,N_35149);
nand U37067 (N_37067,N_34814,N_35192);
and U37068 (N_37068,N_34929,N_34571);
and U37069 (N_37069,N_34442,N_34167);
nor U37070 (N_37070,N_35562,N_35565);
nand U37071 (N_37071,N_34010,N_35276);
nand U37072 (N_37072,N_34436,N_34724);
xnor U37073 (N_37073,N_35238,N_34418);
nand U37074 (N_37074,N_34595,N_35500);
nand U37075 (N_37075,N_34969,N_35860);
and U37076 (N_37076,N_35727,N_35122);
nor U37077 (N_37077,N_34699,N_34096);
and U37078 (N_37078,N_34302,N_34742);
nand U37079 (N_37079,N_35534,N_34128);
and U37080 (N_37080,N_35312,N_35259);
nor U37081 (N_37081,N_35164,N_34681);
or U37082 (N_37082,N_34490,N_35411);
and U37083 (N_37083,N_35004,N_34384);
nand U37084 (N_37084,N_34414,N_35696);
xnor U37085 (N_37085,N_34478,N_35619);
xnor U37086 (N_37086,N_35260,N_34356);
nand U37087 (N_37087,N_35905,N_34006);
nand U37088 (N_37088,N_34305,N_35302);
nand U37089 (N_37089,N_34573,N_34808);
nand U37090 (N_37090,N_34647,N_35227);
nand U37091 (N_37091,N_35998,N_35167);
and U37092 (N_37092,N_34051,N_35144);
nand U37093 (N_37093,N_34101,N_34929);
nor U37094 (N_37094,N_35055,N_34147);
nand U37095 (N_37095,N_34997,N_34009);
xnor U37096 (N_37096,N_35197,N_34262);
nand U37097 (N_37097,N_34737,N_34216);
or U37098 (N_37098,N_34014,N_34460);
or U37099 (N_37099,N_34645,N_34471);
nand U37100 (N_37100,N_35360,N_34410);
nor U37101 (N_37101,N_34476,N_34353);
or U37102 (N_37102,N_35372,N_35713);
or U37103 (N_37103,N_35147,N_34160);
and U37104 (N_37104,N_34842,N_34680);
xnor U37105 (N_37105,N_35774,N_35745);
nor U37106 (N_37106,N_35734,N_35156);
nand U37107 (N_37107,N_34581,N_35285);
nand U37108 (N_37108,N_35830,N_35401);
or U37109 (N_37109,N_35164,N_35230);
or U37110 (N_37110,N_34614,N_35227);
or U37111 (N_37111,N_34267,N_34520);
and U37112 (N_37112,N_34781,N_35841);
or U37113 (N_37113,N_35454,N_34031);
xnor U37114 (N_37114,N_35350,N_34579);
or U37115 (N_37115,N_34347,N_35857);
nand U37116 (N_37116,N_35263,N_34203);
xor U37117 (N_37117,N_34829,N_34120);
nand U37118 (N_37118,N_34384,N_35671);
nand U37119 (N_37119,N_35171,N_34885);
nor U37120 (N_37120,N_34035,N_34815);
or U37121 (N_37121,N_34178,N_35286);
xnor U37122 (N_37122,N_34490,N_35378);
or U37123 (N_37123,N_35388,N_34721);
or U37124 (N_37124,N_34520,N_35844);
or U37125 (N_37125,N_34527,N_34954);
or U37126 (N_37126,N_34326,N_35168);
and U37127 (N_37127,N_35303,N_34082);
xor U37128 (N_37128,N_34405,N_34728);
xnor U37129 (N_37129,N_35947,N_34680);
nand U37130 (N_37130,N_34036,N_35901);
xnor U37131 (N_37131,N_35968,N_34846);
nor U37132 (N_37132,N_35141,N_35273);
nor U37133 (N_37133,N_35757,N_35807);
nand U37134 (N_37134,N_34091,N_34236);
nor U37135 (N_37135,N_35375,N_34554);
xor U37136 (N_37136,N_34955,N_34685);
nor U37137 (N_37137,N_35749,N_34869);
xnor U37138 (N_37138,N_35818,N_34330);
and U37139 (N_37139,N_35368,N_34830);
nor U37140 (N_37140,N_34285,N_34859);
nand U37141 (N_37141,N_35593,N_34713);
or U37142 (N_37142,N_34703,N_35829);
nor U37143 (N_37143,N_35299,N_34891);
nand U37144 (N_37144,N_35133,N_34880);
or U37145 (N_37145,N_35236,N_34303);
nand U37146 (N_37146,N_34683,N_34741);
nand U37147 (N_37147,N_35006,N_34748);
nand U37148 (N_37148,N_35581,N_35311);
or U37149 (N_37149,N_35663,N_35482);
nor U37150 (N_37150,N_34422,N_34710);
nor U37151 (N_37151,N_35323,N_34303);
and U37152 (N_37152,N_34778,N_34354);
nor U37153 (N_37153,N_34282,N_34243);
xor U37154 (N_37154,N_35050,N_35341);
and U37155 (N_37155,N_35604,N_34734);
xor U37156 (N_37156,N_35647,N_34815);
nand U37157 (N_37157,N_35212,N_35779);
and U37158 (N_37158,N_35226,N_34442);
xor U37159 (N_37159,N_35823,N_34073);
nand U37160 (N_37160,N_34062,N_35879);
and U37161 (N_37161,N_35645,N_34457);
xnor U37162 (N_37162,N_35125,N_35399);
or U37163 (N_37163,N_34559,N_35684);
and U37164 (N_37164,N_34466,N_34123);
or U37165 (N_37165,N_34050,N_34743);
nand U37166 (N_37166,N_34322,N_34099);
nor U37167 (N_37167,N_34711,N_35470);
and U37168 (N_37168,N_35529,N_34532);
xnor U37169 (N_37169,N_34176,N_34536);
nand U37170 (N_37170,N_34681,N_34686);
xor U37171 (N_37171,N_35601,N_35936);
xor U37172 (N_37172,N_35487,N_35573);
nand U37173 (N_37173,N_34122,N_34483);
xor U37174 (N_37174,N_35919,N_34523);
nand U37175 (N_37175,N_35421,N_34850);
nor U37176 (N_37176,N_35544,N_35299);
nor U37177 (N_37177,N_35943,N_34635);
and U37178 (N_37178,N_34661,N_34105);
xnor U37179 (N_37179,N_34601,N_35983);
nor U37180 (N_37180,N_35397,N_34873);
xnor U37181 (N_37181,N_34901,N_35050);
nand U37182 (N_37182,N_34231,N_34052);
xor U37183 (N_37183,N_35031,N_35040);
and U37184 (N_37184,N_34995,N_34364);
nand U37185 (N_37185,N_35233,N_34246);
xnor U37186 (N_37186,N_34581,N_34436);
or U37187 (N_37187,N_35453,N_34590);
nor U37188 (N_37188,N_35380,N_34836);
nor U37189 (N_37189,N_34073,N_34896);
or U37190 (N_37190,N_35949,N_35215);
xor U37191 (N_37191,N_34687,N_35942);
and U37192 (N_37192,N_35655,N_35282);
xor U37193 (N_37193,N_35160,N_34684);
or U37194 (N_37194,N_35245,N_34912);
nand U37195 (N_37195,N_34674,N_35786);
and U37196 (N_37196,N_34401,N_35083);
nand U37197 (N_37197,N_34334,N_35614);
and U37198 (N_37198,N_35431,N_34141);
and U37199 (N_37199,N_34906,N_34133);
and U37200 (N_37200,N_35735,N_35590);
nor U37201 (N_37201,N_34590,N_35467);
nand U37202 (N_37202,N_35186,N_34019);
xor U37203 (N_37203,N_34655,N_34085);
xor U37204 (N_37204,N_34225,N_35765);
or U37205 (N_37205,N_34182,N_35337);
or U37206 (N_37206,N_34407,N_34954);
or U37207 (N_37207,N_35832,N_34523);
xor U37208 (N_37208,N_34396,N_35760);
nor U37209 (N_37209,N_35243,N_34360);
nand U37210 (N_37210,N_34807,N_34929);
xnor U37211 (N_37211,N_35226,N_34315);
nand U37212 (N_37212,N_34955,N_35535);
xor U37213 (N_37213,N_34155,N_34233);
and U37214 (N_37214,N_35307,N_34197);
xnor U37215 (N_37215,N_34645,N_34742);
nor U37216 (N_37216,N_34249,N_34362);
and U37217 (N_37217,N_34541,N_34214);
nor U37218 (N_37218,N_34549,N_34983);
or U37219 (N_37219,N_34122,N_34164);
nand U37220 (N_37220,N_35221,N_34482);
nor U37221 (N_37221,N_34413,N_35446);
or U37222 (N_37222,N_35160,N_34779);
nor U37223 (N_37223,N_34100,N_35247);
nor U37224 (N_37224,N_34549,N_35341);
nand U37225 (N_37225,N_34207,N_35312);
and U37226 (N_37226,N_34821,N_34274);
nand U37227 (N_37227,N_34010,N_35329);
or U37228 (N_37228,N_35008,N_35801);
or U37229 (N_37229,N_34362,N_34810);
xnor U37230 (N_37230,N_34097,N_35712);
and U37231 (N_37231,N_34081,N_34572);
and U37232 (N_37232,N_35191,N_35872);
or U37233 (N_37233,N_35744,N_34283);
nand U37234 (N_37234,N_34665,N_35408);
or U37235 (N_37235,N_34353,N_35627);
and U37236 (N_37236,N_34650,N_34248);
and U37237 (N_37237,N_34169,N_35700);
nand U37238 (N_37238,N_35084,N_35331);
nand U37239 (N_37239,N_34556,N_35324);
and U37240 (N_37240,N_34688,N_34348);
xor U37241 (N_37241,N_35571,N_34889);
and U37242 (N_37242,N_35920,N_34598);
nand U37243 (N_37243,N_35342,N_35087);
xnor U37244 (N_37244,N_34027,N_35028);
or U37245 (N_37245,N_34171,N_35878);
and U37246 (N_37246,N_34944,N_35033);
nand U37247 (N_37247,N_34233,N_34851);
nor U37248 (N_37248,N_35143,N_35286);
and U37249 (N_37249,N_34855,N_34204);
xnor U37250 (N_37250,N_35994,N_34022);
nor U37251 (N_37251,N_35040,N_34999);
and U37252 (N_37252,N_35730,N_35460);
and U37253 (N_37253,N_35046,N_35281);
xor U37254 (N_37254,N_35745,N_35043);
nor U37255 (N_37255,N_34580,N_34124);
nor U37256 (N_37256,N_35988,N_34048);
nand U37257 (N_37257,N_35110,N_35459);
nand U37258 (N_37258,N_34607,N_35412);
nand U37259 (N_37259,N_35588,N_34484);
xor U37260 (N_37260,N_35458,N_34665);
nor U37261 (N_37261,N_34021,N_34969);
xor U37262 (N_37262,N_34140,N_34907);
nand U37263 (N_37263,N_34741,N_35305);
nor U37264 (N_37264,N_34497,N_35392);
nand U37265 (N_37265,N_35403,N_35561);
nor U37266 (N_37266,N_35605,N_34182);
or U37267 (N_37267,N_35484,N_35899);
or U37268 (N_37268,N_34192,N_35945);
nand U37269 (N_37269,N_35946,N_35953);
or U37270 (N_37270,N_35900,N_35204);
nor U37271 (N_37271,N_35283,N_34496);
and U37272 (N_37272,N_34793,N_35214);
and U37273 (N_37273,N_35238,N_35472);
or U37274 (N_37274,N_34846,N_35255);
and U37275 (N_37275,N_34513,N_34640);
or U37276 (N_37276,N_34719,N_35287);
nand U37277 (N_37277,N_35211,N_35273);
nand U37278 (N_37278,N_34902,N_35556);
and U37279 (N_37279,N_35046,N_34894);
or U37280 (N_37280,N_35945,N_34286);
and U37281 (N_37281,N_35684,N_35203);
and U37282 (N_37282,N_35167,N_35434);
xor U37283 (N_37283,N_35740,N_34133);
nand U37284 (N_37284,N_34824,N_34068);
nor U37285 (N_37285,N_34200,N_34453);
nand U37286 (N_37286,N_35946,N_35357);
nor U37287 (N_37287,N_34905,N_35458);
nor U37288 (N_37288,N_35829,N_34846);
nand U37289 (N_37289,N_34378,N_35495);
nand U37290 (N_37290,N_34243,N_35476);
nor U37291 (N_37291,N_34458,N_35940);
xnor U37292 (N_37292,N_34589,N_35123);
and U37293 (N_37293,N_34662,N_35369);
nand U37294 (N_37294,N_35170,N_35705);
nor U37295 (N_37295,N_35304,N_34924);
xnor U37296 (N_37296,N_34614,N_35779);
xor U37297 (N_37297,N_34270,N_35577);
nand U37298 (N_37298,N_35308,N_35649);
and U37299 (N_37299,N_35336,N_34799);
and U37300 (N_37300,N_34271,N_34184);
nor U37301 (N_37301,N_34693,N_34215);
nor U37302 (N_37302,N_35092,N_35538);
or U37303 (N_37303,N_35214,N_35696);
and U37304 (N_37304,N_34569,N_34042);
and U37305 (N_37305,N_34333,N_35843);
xnor U37306 (N_37306,N_35959,N_34969);
nand U37307 (N_37307,N_35487,N_35533);
nor U37308 (N_37308,N_35993,N_35246);
xnor U37309 (N_37309,N_34983,N_35149);
and U37310 (N_37310,N_35391,N_34191);
xnor U37311 (N_37311,N_34966,N_35288);
or U37312 (N_37312,N_35753,N_35151);
xnor U37313 (N_37313,N_35108,N_34824);
nand U37314 (N_37314,N_34811,N_35076);
xor U37315 (N_37315,N_34809,N_35722);
or U37316 (N_37316,N_35142,N_35548);
xor U37317 (N_37317,N_34348,N_34029);
xnor U37318 (N_37318,N_34237,N_34681);
and U37319 (N_37319,N_34421,N_34895);
and U37320 (N_37320,N_35365,N_35064);
or U37321 (N_37321,N_35613,N_35389);
and U37322 (N_37322,N_35168,N_35651);
nor U37323 (N_37323,N_34111,N_34096);
nor U37324 (N_37324,N_34948,N_34873);
and U37325 (N_37325,N_34867,N_35625);
or U37326 (N_37326,N_34955,N_35728);
xnor U37327 (N_37327,N_35875,N_34974);
or U37328 (N_37328,N_34405,N_34439);
xor U37329 (N_37329,N_34120,N_34050);
and U37330 (N_37330,N_34348,N_35096);
nand U37331 (N_37331,N_35927,N_34098);
or U37332 (N_37332,N_34103,N_34807);
nor U37333 (N_37333,N_34489,N_34824);
nor U37334 (N_37334,N_34576,N_35356);
nand U37335 (N_37335,N_34403,N_35828);
xnor U37336 (N_37336,N_34916,N_34719);
or U37337 (N_37337,N_35831,N_34681);
or U37338 (N_37338,N_35963,N_34676);
nand U37339 (N_37339,N_34384,N_34081);
or U37340 (N_37340,N_35374,N_34170);
nor U37341 (N_37341,N_35753,N_35568);
nor U37342 (N_37342,N_34925,N_34649);
and U37343 (N_37343,N_35641,N_35719);
nand U37344 (N_37344,N_34819,N_34983);
nand U37345 (N_37345,N_35903,N_34901);
xnor U37346 (N_37346,N_34073,N_35623);
and U37347 (N_37347,N_34853,N_34836);
or U37348 (N_37348,N_35448,N_34426);
nor U37349 (N_37349,N_34486,N_34703);
and U37350 (N_37350,N_35190,N_34353);
nor U37351 (N_37351,N_34937,N_35826);
nand U37352 (N_37352,N_35915,N_35242);
nor U37353 (N_37353,N_35581,N_34906);
nor U37354 (N_37354,N_34758,N_34624);
nand U37355 (N_37355,N_35656,N_34669);
nand U37356 (N_37356,N_34513,N_35666);
and U37357 (N_37357,N_35831,N_35127);
or U37358 (N_37358,N_34656,N_34462);
nand U37359 (N_37359,N_35759,N_35695);
nor U37360 (N_37360,N_35656,N_34870);
and U37361 (N_37361,N_35348,N_34409);
nand U37362 (N_37362,N_34489,N_35990);
nor U37363 (N_37363,N_34280,N_34379);
and U37364 (N_37364,N_34839,N_34870);
xor U37365 (N_37365,N_34899,N_35946);
or U37366 (N_37366,N_35479,N_35396);
nand U37367 (N_37367,N_35458,N_34856);
nor U37368 (N_37368,N_34775,N_35052);
and U37369 (N_37369,N_35647,N_34603);
nand U37370 (N_37370,N_35920,N_35353);
and U37371 (N_37371,N_35578,N_35523);
and U37372 (N_37372,N_34121,N_35546);
nor U37373 (N_37373,N_34940,N_35217);
and U37374 (N_37374,N_34630,N_35744);
nor U37375 (N_37375,N_35928,N_34735);
nand U37376 (N_37376,N_34295,N_34846);
and U37377 (N_37377,N_34557,N_35225);
and U37378 (N_37378,N_35842,N_35582);
xnor U37379 (N_37379,N_35485,N_35758);
or U37380 (N_37380,N_35875,N_35733);
xnor U37381 (N_37381,N_34044,N_34057);
xor U37382 (N_37382,N_34111,N_35183);
and U37383 (N_37383,N_35705,N_34195);
nand U37384 (N_37384,N_34759,N_35580);
and U37385 (N_37385,N_34980,N_34884);
or U37386 (N_37386,N_35172,N_35934);
or U37387 (N_37387,N_34621,N_34245);
nor U37388 (N_37388,N_35774,N_35967);
nand U37389 (N_37389,N_35692,N_35894);
xor U37390 (N_37390,N_34116,N_35957);
xnor U37391 (N_37391,N_34102,N_34068);
xor U37392 (N_37392,N_34341,N_35125);
and U37393 (N_37393,N_35893,N_35621);
or U37394 (N_37394,N_34161,N_34737);
xor U37395 (N_37395,N_35422,N_34583);
or U37396 (N_37396,N_34237,N_34061);
and U37397 (N_37397,N_35342,N_35371);
nand U37398 (N_37398,N_34350,N_34007);
and U37399 (N_37399,N_35903,N_35661);
or U37400 (N_37400,N_35441,N_35269);
xnor U37401 (N_37401,N_35521,N_35095);
and U37402 (N_37402,N_34956,N_34987);
or U37403 (N_37403,N_35218,N_34215);
or U37404 (N_37404,N_34843,N_34157);
nand U37405 (N_37405,N_35422,N_34299);
nand U37406 (N_37406,N_34343,N_34235);
and U37407 (N_37407,N_34536,N_34877);
or U37408 (N_37408,N_34716,N_35540);
nand U37409 (N_37409,N_34247,N_34905);
xnor U37410 (N_37410,N_34549,N_34439);
and U37411 (N_37411,N_34331,N_35685);
xor U37412 (N_37412,N_34411,N_34890);
or U37413 (N_37413,N_34591,N_34888);
nand U37414 (N_37414,N_35007,N_34799);
nand U37415 (N_37415,N_35625,N_35905);
nand U37416 (N_37416,N_35532,N_34690);
and U37417 (N_37417,N_34806,N_34430);
nand U37418 (N_37418,N_34344,N_35797);
xnor U37419 (N_37419,N_35305,N_35050);
nor U37420 (N_37420,N_34996,N_35492);
nor U37421 (N_37421,N_35644,N_34666);
and U37422 (N_37422,N_35568,N_35280);
and U37423 (N_37423,N_34453,N_35151);
nand U37424 (N_37424,N_34371,N_34227);
xor U37425 (N_37425,N_34545,N_35378);
or U37426 (N_37426,N_35697,N_34934);
xor U37427 (N_37427,N_35925,N_34109);
nor U37428 (N_37428,N_34566,N_34623);
xor U37429 (N_37429,N_35385,N_34627);
xor U37430 (N_37430,N_34076,N_35237);
nand U37431 (N_37431,N_35510,N_34041);
or U37432 (N_37432,N_35019,N_35322);
or U37433 (N_37433,N_34735,N_34841);
and U37434 (N_37434,N_34638,N_35887);
xnor U37435 (N_37435,N_34019,N_35758);
xor U37436 (N_37436,N_34042,N_35705);
nand U37437 (N_37437,N_34549,N_34528);
nor U37438 (N_37438,N_35017,N_35258);
xor U37439 (N_37439,N_35299,N_34797);
nand U37440 (N_37440,N_35120,N_34080);
xnor U37441 (N_37441,N_34768,N_35661);
nor U37442 (N_37442,N_34736,N_34578);
or U37443 (N_37443,N_35382,N_35387);
xnor U37444 (N_37444,N_35721,N_35669);
xnor U37445 (N_37445,N_34385,N_35758);
nor U37446 (N_37446,N_34246,N_34544);
xnor U37447 (N_37447,N_35962,N_35660);
xor U37448 (N_37448,N_35233,N_35729);
and U37449 (N_37449,N_35273,N_35054);
nand U37450 (N_37450,N_34091,N_35116);
and U37451 (N_37451,N_34486,N_35000);
nand U37452 (N_37452,N_34951,N_34745);
and U37453 (N_37453,N_34563,N_34231);
and U37454 (N_37454,N_35727,N_35671);
xor U37455 (N_37455,N_34443,N_34676);
xor U37456 (N_37456,N_35570,N_34042);
and U37457 (N_37457,N_34445,N_34297);
and U37458 (N_37458,N_34431,N_35654);
nand U37459 (N_37459,N_35263,N_34772);
nor U37460 (N_37460,N_35814,N_34815);
or U37461 (N_37461,N_35179,N_35270);
nand U37462 (N_37462,N_35968,N_34054);
and U37463 (N_37463,N_35487,N_35645);
or U37464 (N_37464,N_34429,N_34325);
nor U37465 (N_37465,N_34838,N_34602);
xnor U37466 (N_37466,N_34534,N_35373);
and U37467 (N_37467,N_35805,N_34450);
xnor U37468 (N_37468,N_34199,N_35963);
and U37469 (N_37469,N_35244,N_35280);
and U37470 (N_37470,N_35068,N_35354);
and U37471 (N_37471,N_34071,N_34313);
and U37472 (N_37472,N_35822,N_35992);
nand U37473 (N_37473,N_35009,N_35147);
xor U37474 (N_37474,N_34027,N_35361);
nor U37475 (N_37475,N_35711,N_35816);
or U37476 (N_37476,N_34510,N_34328);
nand U37477 (N_37477,N_35235,N_34926);
xnor U37478 (N_37478,N_35624,N_34444);
and U37479 (N_37479,N_35491,N_35051);
or U37480 (N_37480,N_34850,N_34575);
or U37481 (N_37481,N_34615,N_35943);
or U37482 (N_37482,N_35079,N_35481);
nand U37483 (N_37483,N_35012,N_35840);
nor U37484 (N_37484,N_34030,N_34932);
or U37485 (N_37485,N_34903,N_35582);
xor U37486 (N_37486,N_34252,N_34584);
or U37487 (N_37487,N_35497,N_34249);
xor U37488 (N_37488,N_35356,N_34676);
nor U37489 (N_37489,N_34050,N_34430);
and U37490 (N_37490,N_35697,N_35203);
or U37491 (N_37491,N_35087,N_35260);
or U37492 (N_37492,N_35320,N_34882);
and U37493 (N_37493,N_35526,N_35853);
xor U37494 (N_37494,N_35773,N_34752);
nor U37495 (N_37495,N_35725,N_34671);
nand U37496 (N_37496,N_35699,N_34547);
xor U37497 (N_37497,N_35405,N_35971);
and U37498 (N_37498,N_35525,N_35578);
nor U37499 (N_37499,N_35135,N_35942);
and U37500 (N_37500,N_35904,N_35631);
or U37501 (N_37501,N_34732,N_35443);
nand U37502 (N_37502,N_34176,N_34338);
xnor U37503 (N_37503,N_34947,N_34925);
xnor U37504 (N_37504,N_34929,N_34038);
or U37505 (N_37505,N_35948,N_34390);
nand U37506 (N_37506,N_34529,N_35549);
and U37507 (N_37507,N_34111,N_35882);
nor U37508 (N_37508,N_34996,N_34541);
nand U37509 (N_37509,N_34439,N_34690);
xnor U37510 (N_37510,N_34960,N_35033);
and U37511 (N_37511,N_34191,N_34834);
or U37512 (N_37512,N_34581,N_34260);
or U37513 (N_37513,N_35291,N_35510);
xnor U37514 (N_37514,N_34284,N_34326);
nor U37515 (N_37515,N_35564,N_35859);
nor U37516 (N_37516,N_34070,N_35878);
nand U37517 (N_37517,N_34338,N_34636);
xor U37518 (N_37518,N_35462,N_34487);
xor U37519 (N_37519,N_35141,N_34014);
xnor U37520 (N_37520,N_34958,N_34694);
or U37521 (N_37521,N_34699,N_34973);
nand U37522 (N_37522,N_34287,N_35130);
xor U37523 (N_37523,N_35506,N_34867);
nand U37524 (N_37524,N_35693,N_34025);
nor U37525 (N_37525,N_35176,N_34824);
nor U37526 (N_37526,N_35349,N_34693);
nand U37527 (N_37527,N_34234,N_35586);
or U37528 (N_37528,N_35771,N_34072);
nor U37529 (N_37529,N_35679,N_34212);
or U37530 (N_37530,N_34727,N_34040);
or U37531 (N_37531,N_35004,N_34068);
and U37532 (N_37532,N_35546,N_35647);
nor U37533 (N_37533,N_35855,N_34445);
or U37534 (N_37534,N_35843,N_35135);
and U37535 (N_37535,N_35936,N_34565);
or U37536 (N_37536,N_34711,N_34623);
nor U37537 (N_37537,N_34555,N_35163);
or U37538 (N_37538,N_35816,N_35969);
nand U37539 (N_37539,N_34250,N_34354);
xor U37540 (N_37540,N_35229,N_34520);
nand U37541 (N_37541,N_34490,N_35676);
xnor U37542 (N_37542,N_35087,N_35915);
nor U37543 (N_37543,N_35030,N_34442);
nand U37544 (N_37544,N_35524,N_34538);
nand U37545 (N_37545,N_34169,N_34031);
nand U37546 (N_37546,N_34339,N_34296);
nand U37547 (N_37547,N_34922,N_35439);
nand U37548 (N_37548,N_35092,N_35412);
and U37549 (N_37549,N_34499,N_34245);
and U37550 (N_37550,N_34598,N_34828);
xor U37551 (N_37551,N_34895,N_34296);
or U37552 (N_37552,N_34578,N_35716);
and U37553 (N_37553,N_35115,N_35553);
nor U37554 (N_37554,N_35308,N_35583);
and U37555 (N_37555,N_35620,N_35408);
or U37556 (N_37556,N_34525,N_34848);
nand U37557 (N_37557,N_35287,N_35317);
nand U37558 (N_37558,N_34257,N_34767);
and U37559 (N_37559,N_35369,N_35624);
nor U37560 (N_37560,N_35377,N_35380);
xor U37561 (N_37561,N_34025,N_34992);
nand U37562 (N_37562,N_34454,N_35150);
and U37563 (N_37563,N_34694,N_35680);
and U37564 (N_37564,N_34675,N_35360);
nand U37565 (N_37565,N_34642,N_34102);
and U37566 (N_37566,N_34412,N_34297);
nor U37567 (N_37567,N_34310,N_35375);
nand U37568 (N_37568,N_35745,N_35520);
nand U37569 (N_37569,N_34469,N_34462);
nand U37570 (N_37570,N_34743,N_35080);
xnor U37571 (N_37571,N_34483,N_35359);
nand U37572 (N_37572,N_35701,N_34315);
xor U37573 (N_37573,N_34883,N_34221);
xnor U37574 (N_37574,N_34164,N_35038);
xor U37575 (N_37575,N_35031,N_35901);
or U37576 (N_37576,N_34321,N_35651);
nand U37577 (N_37577,N_35645,N_35510);
nand U37578 (N_37578,N_34235,N_34531);
and U37579 (N_37579,N_35563,N_35202);
or U37580 (N_37580,N_34735,N_34239);
or U37581 (N_37581,N_34482,N_35362);
xnor U37582 (N_37582,N_35352,N_35455);
or U37583 (N_37583,N_35595,N_34923);
xor U37584 (N_37584,N_35793,N_35741);
nand U37585 (N_37585,N_35000,N_35871);
or U37586 (N_37586,N_35297,N_35217);
nand U37587 (N_37587,N_34691,N_34871);
nand U37588 (N_37588,N_34008,N_35850);
or U37589 (N_37589,N_34784,N_34520);
xnor U37590 (N_37590,N_34036,N_34657);
or U37591 (N_37591,N_34742,N_34438);
xor U37592 (N_37592,N_34909,N_34181);
nor U37593 (N_37593,N_35083,N_34100);
or U37594 (N_37594,N_35455,N_34345);
xor U37595 (N_37595,N_34931,N_34491);
and U37596 (N_37596,N_34038,N_35467);
xor U37597 (N_37597,N_34470,N_35538);
and U37598 (N_37598,N_35942,N_34038);
or U37599 (N_37599,N_34400,N_34885);
xor U37600 (N_37600,N_34859,N_35073);
or U37601 (N_37601,N_34321,N_34821);
and U37602 (N_37602,N_35570,N_34648);
and U37603 (N_37603,N_34213,N_35835);
nor U37604 (N_37604,N_35401,N_35158);
and U37605 (N_37605,N_35170,N_35338);
and U37606 (N_37606,N_34433,N_34564);
nand U37607 (N_37607,N_35578,N_34500);
and U37608 (N_37608,N_35861,N_35784);
and U37609 (N_37609,N_35967,N_34647);
nor U37610 (N_37610,N_35488,N_35260);
xor U37611 (N_37611,N_34515,N_34256);
nand U37612 (N_37612,N_35527,N_35840);
and U37613 (N_37613,N_34832,N_35248);
xor U37614 (N_37614,N_34923,N_35473);
or U37615 (N_37615,N_35535,N_35387);
or U37616 (N_37616,N_35040,N_34288);
nand U37617 (N_37617,N_35564,N_35634);
and U37618 (N_37618,N_34697,N_34757);
nand U37619 (N_37619,N_35435,N_34102);
nor U37620 (N_37620,N_34712,N_35706);
or U37621 (N_37621,N_35464,N_35026);
or U37622 (N_37622,N_34874,N_34392);
nand U37623 (N_37623,N_35459,N_35719);
or U37624 (N_37624,N_34009,N_35462);
nor U37625 (N_37625,N_35640,N_35714);
xor U37626 (N_37626,N_34903,N_34399);
nand U37627 (N_37627,N_35734,N_34317);
and U37628 (N_37628,N_34654,N_34156);
nor U37629 (N_37629,N_35307,N_34206);
nor U37630 (N_37630,N_35692,N_34433);
or U37631 (N_37631,N_35114,N_34942);
nand U37632 (N_37632,N_35622,N_34578);
nand U37633 (N_37633,N_34491,N_34470);
nand U37634 (N_37634,N_35616,N_34061);
xor U37635 (N_37635,N_35027,N_35333);
nand U37636 (N_37636,N_35421,N_35893);
nand U37637 (N_37637,N_34353,N_35114);
nand U37638 (N_37638,N_35039,N_35224);
or U37639 (N_37639,N_34738,N_35463);
nand U37640 (N_37640,N_35160,N_34711);
or U37641 (N_37641,N_35064,N_34241);
nand U37642 (N_37642,N_35143,N_35497);
or U37643 (N_37643,N_34834,N_34779);
xnor U37644 (N_37644,N_34109,N_35899);
or U37645 (N_37645,N_34822,N_34070);
and U37646 (N_37646,N_35975,N_35571);
nor U37647 (N_37647,N_34628,N_34448);
nand U37648 (N_37648,N_34616,N_34974);
nand U37649 (N_37649,N_35059,N_34270);
nand U37650 (N_37650,N_34993,N_35264);
or U37651 (N_37651,N_34435,N_35952);
or U37652 (N_37652,N_35421,N_34104);
nor U37653 (N_37653,N_34257,N_35449);
and U37654 (N_37654,N_34677,N_34663);
xor U37655 (N_37655,N_34235,N_35376);
or U37656 (N_37656,N_34315,N_35536);
xor U37657 (N_37657,N_34379,N_35173);
and U37658 (N_37658,N_34945,N_35676);
and U37659 (N_37659,N_35611,N_34681);
xor U37660 (N_37660,N_35614,N_34104);
and U37661 (N_37661,N_34712,N_35054);
or U37662 (N_37662,N_35512,N_35126);
xnor U37663 (N_37663,N_35712,N_34309);
xnor U37664 (N_37664,N_35162,N_34451);
nor U37665 (N_37665,N_35403,N_34854);
nor U37666 (N_37666,N_35672,N_34024);
xor U37667 (N_37667,N_35948,N_34720);
nor U37668 (N_37668,N_34116,N_35527);
xor U37669 (N_37669,N_35447,N_35759);
nor U37670 (N_37670,N_34454,N_35299);
and U37671 (N_37671,N_35450,N_35596);
xnor U37672 (N_37672,N_34622,N_35324);
xor U37673 (N_37673,N_34346,N_35601);
xor U37674 (N_37674,N_34668,N_35091);
nor U37675 (N_37675,N_35750,N_34008);
nor U37676 (N_37676,N_35358,N_34872);
or U37677 (N_37677,N_34682,N_34958);
nand U37678 (N_37678,N_34717,N_35744);
or U37679 (N_37679,N_34696,N_34602);
nand U37680 (N_37680,N_35709,N_34466);
nor U37681 (N_37681,N_34433,N_35318);
nand U37682 (N_37682,N_35250,N_34088);
xnor U37683 (N_37683,N_34339,N_35889);
nor U37684 (N_37684,N_34947,N_34015);
and U37685 (N_37685,N_34676,N_34646);
or U37686 (N_37686,N_35223,N_35439);
nor U37687 (N_37687,N_34678,N_35778);
nor U37688 (N_37688,N_34625,N_34260);
xor U37689 (N_37689,N_34654,N_34961);
xor U37690 (N_37690,N_35174,N_35255);
and U37691 (N_37691,N_35154,N_34398);
nor U37692 (N_37692,N_35701,N_34606);
xor U37693 (N_37693,N_34202,N_35984);
and U37694 (N_37694,N_35192,N_35306);
nand U37695 (N_37695,N_34969,N_34108);
xor U37696 (N_37696,N_35372,N_35152);
or U37697 (N_37697,N_34707,N_34801);
nor U37698 (N_37698,N_35511,N_34436);
and U37699 (N_37699,N_34121,N_35494);
or U37700 (N_37700,N_34717,N_35847);
and U37701 (N_37701,N_35177,N_34523);
xor U37702 (N_37702,N_35555,N_34562);
and U37703 (N_37703,N_34687,N_34347);
nor U37704 (N_37704,N_34511,N_35655);
nand U37705 (N_37705,N_35067,N_35733);
and U37706 (N_37706,N_35160,N_35036);
xor U37707 (N_37707,N_34118,N_35070);
nor U37708 (N_37708,N_35570,N_34787);
nand U37709 (N_37709,N_34942,N_35089);
and U37710 (N_37710,N_34314,N_34781);
xnor U37711 (N_37711,N_34853,N_35207);
and U37712 (N_37712,N_35902,N_34134);
or U37713 (N_37713,N_34529,N_35005);
xnor U37714 (N_37714,N_35525,N_34635);
xnor U37715 (N_37715,N_34836,N_34774);
nand U37716 (N_37716,N_35115,N_35058);
xnor U37717 (N_37717,N_34446,N_35072);
nand U37718 (N_37718,N_34666,N_34007);
nor U37719 (N_37719,N_34283,N_34730);
nand U37720 (N_37720,N_34757,N_34566);
nand U37721 (N_37721,N_35809,N_34015);
xor U37722 (N_37722,N_35212,N_35122);
nand U37723 (N_37723,N_35656,N_35140);
xor U37724 (N_37724,N_34680,N_35556);
nor U37725 (N_37725,N_34685,N_35471);
nand U37726 (N_37726,N_35506,N_34404);
xnor U37727 (N_37727,N_34817,N_34837);
or U37728 (N_37728,N_34972,N_34286);
nor U37729 (N_37729,N_34340,N_35035);
xor U37730 (N_37730,N_35141,N_34499);
and U37731 (N_37731,N_34552,N_34236);
xor U37732 (N_37732,N_34465,N_35793);
nor U37733 (N_37733,N_34859,N_34864);
nand U37734 (N_37734,N_34236,N_35774);
nand U37735 (N_37735,N_34329,N_34809);
or U37736 (N_37736,N_35284,N_35366);
or U37737 (N_37737,N_34871,N_35882);
and U37738 (N_37738,N_34117,N_34144);
and U37739 (N_37739,N_34233,N_35921);
and U37740 (N_37740,N_34849,N_35515);
or U37741 (N_37741,N_35570,N_35992);
nand U37742 (N_37742,N_35745,N_34815);
nand U37743 (N_37743,N_35963,N_35659);
or U37744 (N_37744,N_35115,N_34374);
nor U37745 (N_37745,N_34485,N_35761);
xor U37746 (N_37746,N_34625,N_35454);
xnor U37747 (N_37747,N_34889,N_34685);
nor U37748 (N_37748,N_35165,N_35248);
xnor U37749 (N_37749,N_34666,N_35529);
or U37750 (N_37750,N_34510,N_34142);
or U37751 (N_37751,N_34275,N_35155);
xnor U37752 (N_37752,N_34052,N_35088);
xor U37753 (N_37753,N_34421,N_34740);
nand U37754 (N_37754,N_35109,N_34471);
xor U37755 (N_37755,N_35634,N_34303);
and U37756 (N_37756,N_34127,N_34383);
and U37757 (N_37757,N_34083,N_34257);
nand U37758 (N_37758,N_34350,N_35430);
xnor U37759 (N_37759,N_35825,N_35186);
nand U37760 (N_37760,N_35640,N_35341);
nand U37761 (N_37761,N_35494,N_34463);
nor U37762 (N_37762,N_34552,N_34348);
and U37763 (N_37763,N_35361,N_35721);
or U37764 (N_37764,N_35071,N_34042);
nand U37765 (N_37765,N_34111,N_35912);
nand U37766 (N_37766,N_34015,N_34806);
and U37767 (N_37767,N_34777,N_34610);
nand U37768 (N_37768,N_35719,N_34098);
xor U37769 (N_37769,N_35378,N_35080);
xnor U37770 (N_37770,N_34991,N_35584);
nor U37771 (N_37771,N_35999,N_34207);
or U37772 (N_37772,N_34467,N_35929);
xnor U37773 (N_37773,N_34149,N_34769);
nor U37774 (N_37774,N_34270,N_34034);
xor U37775 (N_37775,N_35342,N_35887);
xnor U37776 (N_37776,N_35782,N_34895);
xnor U37777 (N_37777,N_35232,N_34617);
and U37778 (N_37778,N_35558,N_35689);
nor U37779 (N_37779,N_34467,N_35490);
nor U37780 (N_37780,N_34647,N_34057);
and U37781 (N_37781,N_34890,N_35646);
xor U37782 (N_37782,N_34117,N_35719);
nor U37783 (N_37783,N_35135,N_35603);
nand U37784 (N_37784,N_35002,N_34889);
or U37785 (N_37785,N_35945,N_34652);
and U37786 (N_37786,N_35653,N_34547);
nor U37787 (N_37787,N_35106,N_34024);
xnor U37788 (N_37788,N_34525,N_34901);
or U37789 (N_37789,N_34957,N_35696);
or U37790 (N_37790,N_34241,N_34350);
nand U37791 (N_37791,N_34590,N_34313);
xor U37792 (N_37792,N_35409,N_35260);
nor U37793 (N_37793,N_35678,N_35588);
xnor U37794 (N_37794,N_34748,N_34401);
and U37795 (N_37795,N_34900,N_35691);
nand U37796 (N_37796,N_35718,N_35281);
xor U37797 (N_37797,N_35258,N_34742);
nand U37798 (N_37798,N_34388,N_35889);
and U37799 (N_37799,N_35678,N_35255);
xor U37800 (N_37800,N_35628,N_34093);
nor U37801 (N_37801,N_34942,N_34268);
and U37802 (N_37802,N_34708,N_34061);
nand U37803 (N_37803,N_35305,N_34945);
or U37804 (N_37804,N_34936,N_35703);
xor U37805 (N_37805,N_34451,N_34358);
and U37806 (N_37806,N_34113,N_35082);
nor U37807 (N_37807,N_34496,N_35236);
nor U37808 (N_37808,N_34471,N_34507);
and U37809 (N_37809,N_34043,N_35020);
xor U37810 (N_37810,N_34868,N_34257);
nand U37811 (N_37811,N_35014,N_34478);
nor U37812 (N_37812,N_35508,N_35820);
nor U37813 (N_37813,N_34493,N_35025);
nand U37814 (N_37814,N_34405,N_35851);
or U37815 (N_37815,N_35108,N_35282);
nand U37816 (N_37816,N_35212,N_35224);
and U37817 (N_37817,N_34420,N_34948);
or U37818 (N_37818,N_34610,N_34649);
or U37819 (N_37819,N_35188,N_35608);
nor U37820 (N_37820,N_34849,N_34192);
or U37821 (N_37821,N_35342,N_35422);
xor U37822 (N_37822,N_35277,N_35691);
nand U37823 (N_37823,N_34839,N_35821);
xnor U37824 (N_37824,N_34319,N_35565);
nor U37825 (N_37825,N_35527,N_35566);
nor U37826 (N_37826,N_34565,N_35652);
nand U37827 (N_37827,N_34259,N_34101);
xnor U37828 (N_37828,N_35542,N_35265);
and U37829 (N_37829,N_34878,N_34101);
or U37830 (N_37830,N_35355,N_35261);
or U37831 (N_37831,N_35579,N_34884);
xor U37832 (N_37832,N_34021,N_35110);
nor U37833 (N_37833,N_35605,N_35856);
and U37834 (N_37834,N_34914,N_35740);
xnor U37835 (N_37835,N_34888,N_34984);
and U37836 (N_37836,N_35762,N_35891);
nor U37837 (N_37837,N_35964,N_34127);
xnor U37838 (N_37838,N_35011,N_34161);
or U37839 (N_37839,N_34212,N_34789);
or U37840 (N_37840,N_35680,N_34573);
nand U37841 (N_37841,N_34464,N_35795);
or U37842 (N_37842,N_35729,N_34467);
nor U37843 (N_37843,N_35366,N_35397);
or U37844 (N_37844,N_34106,N_35871);
nand U37845 (N_37845,N_34397,N_35060);
xnor U37846 (N_37846,N_34226,N_34949);
nand U37847 (N_37847,N_35903,N_34364);
nor U37848 (N_37848,N_34716,N_35673);
and U37849 (N_37849,N_34769,N_35169);
nand U37850 (N_37850,N_34622,N_34037);
xor U37851 (N_37851,N_34789,N_34043);
or U37852 (N_37852,N_35936,N_34378);
xor U37853 (N_37853,N_34669,N_35381);
nand U37854 (N_37854,N_34445,N_35636);
or U37855 (N_37855,N_34764,N_35704);
nand U37856 (N_37856,N_35235,N_34917);
xnor U37857 (N_37857,N_35239,N_35255);
nand U37858 (N_37858,N_35902,N_35533);
xnor U37859 (N_37859,N_35008,N_34132);
or U37860 (N_37860,N_35955,N_34743);
nand U37861 (N_37861,N_34004,N_34604);
nor U37862 (N_37862,N_35158,N_35787);
xor U37863 (N_37863,N_35131,N_34765);
nand U37864 (N_37864,N_35997,N_35571);
nand U37865 (N_37865,N_34921,N_34963);
and U37866 (N_37866,N_34477,N_34715);
nor U37867 (N_37867,N_35341,N_34345);
or U37868 (N_37868,N_34119,N_34791);
xor U37869 (N_37869,N_34868,N_34387);
nand U37870 (N_37870,N_34909,N_34666);
nor U37871 (N_37871,N_35979,N_34400);
and U37872 (N_37872,N_35444,N_34349);
and U37873 (N_37873,N_34906,N_35795);
nor U37874 (N_37874,N_34352,N_34238);
nand U37875 (N_37875,N_35970,N_34739);
nor U37876 (N_37876,N_34346,N_35659);
or U37877 (N_37877,N_34708,N_34243);
or U37878 (N_37878,N_35803,N_34681);
nor U37879 (N_37879,N_34419,N_35707);
nand U37880 (N_37880,N_35042,N_34749);
xor U37881 (N_37881,N_34547,N_34540);
xor U37882 (N_37882,N_35641,N_34137);
nand U37883 (N_37883,N_35072,N_35774);
nor U37884 (N_37884,N_35627,N_35283);
and U37885 (N_37885,N_34646,N_34595);
xor U37886 (N_37886,N_34708,N_34908);
nand U37887 (N_37887,N_34906,N_34160);
xor U37888 (N_37888,N_34733,N_34374);
or U37889 (N_37889,N_35056,N_35349);
xnor U37890 (N_37890,N_35744,N_34774);
xor U37891 (N_37891,N_35202,N_35664);
nor U37892 (N_37892,N_34972,N_34479);
and U37893 (N_37893,N_34543,N_34443);
or U37894 (N_37894,N_35492,N_34107);
nand U37895 (N_37895,N_34052,N_34617);
nor U37896 (N_37896,N_35623,N_35866);
and U37897 (N_37897,N_34202,N_35871);
and U37898 (N_37898,N_34507,N_35829);
nor U37899 (N_37899,N_34791,N_34847);
xnor U37900 (N_37900,N_34481,N_34159);
xnor U37901 (N_37901,N_34184,N_35547);
nand U37902 (N_37902,N_35916,N_34646);
xor U37903 (N_37903,N_35671,N_34843);
xor U37904 (N_37904,N_35004,N_35873);
nand U37905 (N_37905,N_35252,N_34510);
xor U37906 (N_37906,N_35957,N_35562);
nand U37907 (N_37907,N_34699,N_35819);
nor U37908 (N_37908,N_34673,N_34560);
and U37909 (N_37909,N_35573,N_34081);
nor U37910 (N_37910,N_35636,N_34123);
nor U37911 (N_37911,N_35623,N_34954);
and U37912 (N_37912,N_35727,N_35665);
nand U37913 (N_37913,N_34168,N_35274);
and U37914 (N_37914,N_34197,N_34473);
nor U37915 (N_37915,N_34342,N_34969);
and U37916 (N_37916,N_35409,N_34824);
nand U37917 (N_37917,N_35305,N_34788);
xor U37918 (N_37918,N_35663,N_35793);
or U37919 (N_37919,N_34713,N_35300);
nor U37920 (N_37920,N_34342,N_34914);
nand U37921 (N_37921,N_34522,N_34107);
and U37922 (N_37922,N_35392,N_35255);
and U37923 (N_37923,N_34930,N_35217);
nand U37924 (N_37924,N_35956,N_34149);
or U37925 (N_37925,N_34874,N_35690);
nand U37926 (N_37926,N_35251,N_35736);
or U37927 (N_37927,N_35887,N_35680);
xor U37928 (N_37928,N_35880,N_34891);
nand U37929 (N_37929,N_34541,N_34385);
or U37930 (N_37930,N_35646,N_35575);
nor U37931 (N_37931,N_35923,N_35307);
nand U37932 (N_37932,N_34111,N_35730);
and U37933 (N_37933,N_35555,N_34646);
nor U37934 (N_37934,N_34430,N_35434);
nor U37935 (N_37935,N_34622,N_34864);
and U37936 (N_37936,N_35473,N_35916);
or U37937 (N_37937,N_34689,N_35174);
or U37938 (N_37938,N_34987,N_35896);
xor U37939 (N_37939,N_35048,N_34613);
nand U37940 (N_37940,N_34329,N_35230);
or U37941 (N_37941,N_35900,N_35733);
or U37942 (N_37942,N_35886,N_35111);
and U37943 (N_37943,N_34645,N_34473);
or U37944 (N_37944,N_34542,N_35201);
xor U37945 (N_37945,N_34505,N_34259);
xor U37946 (N_37946,N_35443,N_35805);
and U37947 (N_37947,N_34245,N_35788);
nor U37948 (N_37948,N_34364,N_35455);
nand U37949 (N_37949,N_35631,N_34186);
nor U37950 (N_37950,N_34581,N_34885);
nand U37951 (N_37951,N_35988,N_35440);
nor U37952 (N_37952,N_34114,N_34333);
nand U37953 (N_37953,N_35756,N_35726);
and U37954 (N_37954,N_34484,N_34154);
nand U37955 (N_37955,N_34077,N_35003);
nor U37956 (N_37956,N_35900,N_34562);
xnor U37957 (N_37957,N_34595,N_34693);
xnor U37958 (N_37958,N_35194,N_35509);
nor U37959 (N_37959,N_35847,N_34959);
and U37960 (N_37960,N_35119,N_35687);
nor U37961 (N_37961,N_34331,N_34307);
or U37962 (N_37962,N_35765,N_35133);
xnor U37963 (N_37963,N_35209,N_35570);
nor U37964 (N_37964,N_34529,N_34487);
or U37965 (N_37965,N_35889,N_35953);
nor U37966 (N_37966,N_35412,N_34600);
xnor U37967 (N_37967,N_34011,N_34288);
xnor U37968 (N_37968,N_35935,N_34406);
nor U37969 (N_37969,N_35030,N_35597);
nand U37970 (N_37970,N_35903,N_35634);
xnor U37971 (N_37971,N_35430,N_35139);
and U37972 (N_37972,N_34134,N_35210);
or U37973 (N_37973,N_34503,N_35531);
nor U37974 (N_37974,N_34101,N_34320);
nor U37975 (N_37975,N_34431,N_34767);
xnor U37976 (N_37976,N_34851,N_35622);
nand U37977 (N_37977,N_35120,N_34546);
nor U37978 (N_37978,N_34690,N_34815);
or U37979 (N_37979,N_34310,N_34715);
nor U37980 (N_37980,N_35677,N_35544);
nor U37981 (N_37981,N_34638,N_34270);
xnor U37982 (N_37982,N_34860,N_34733);
and U37983 (N_37983,N_35186,N_35030);
or U37984 (N_37984,N_35173,N_35168);
nand U37985 (N_37985,N_35290,N_35355);
and U37986 (N_37986,N_35403,N_34653);
or U37987 (N_37987,N_35981,N_34308);
or U37988 (N_37988,N_35848,N_34851);
and U37989 (N_37989,N_34109,N_34658);
or U37990 (N_37990,N_35806,N_34411);
nor U37991 (N_37991,N_35588,N_34433);
xnor U37992 (N_37992,N_35412,N_35349);
nor U37993 (N_37993,N_35432,N_35422);
xnor U37994 (N_37994,N_34145,N_34389);
or U37995 (N_37995,N_34753,N_34493);
nand U37996 (N_37996,N_35151,N_34766);
nor U37997 (N_37997,N_35626,N_34781);
and U37998 (N_37998,N_35954,N_34989);
or U37999 (N_37999,N_34706,N_34687);
nand U38000 (N_38000,N_36856,N_37656);
nor U38001 (N_38001,N_37475,N_37830);
xor U38002 (N_38002,N_37291,N_37378);
xnor U38003 (N_38003,N_37328,N_37855);
or U38004 (N_38004,N_36608,N_36842);
nor U38005 (N_38005,N_37095,N_36754);
nand U38006 (N_38006,N_36772,N_37148);
nand U38007 (N_38007,N_36675,N_36759);
nand U38008 (N_38008,N_37607,N_37247);
or U38009 (N_38009,N_37957,N_36936);
and U38010 (N_38010,N_36686,N_37817);
nor U38011 (N_38011,N_36069,N_37814);
and U38012 (N_38012,N_36108,N_37015);
or U38013 (N_38013,N_37780,N_36888);
xor U38014 (N_38014,N_36433,N_37728);
nand U38015 (N_38015,N_36828,N_37142);
and U38016 (N_38016,N_37982,N_37449);
or U38017 (N_38017,N_36177,N_37308);
nor U38018 (N_38018,N_36139,N_36379);
nor U38019 (N_38019,N_36629,N_37287);
and U38020 (N_38020,N_37663,N_36212);
nor U38021 (N_38021,N_36081,N_36438);
nor U38022 (N_38022,N_37258,N_37877);
and U38023 (N_38023,N_37377,N_36193);
nand U38024 (N_38024,N_37571,N_37596);
nand U38025 (N_38025,N_37051,N_37742);
and U38026 (N_38026,N_36573,N_36718);
nor U38027 (N_38027,N_36033,N_37803);
nor U38028 (N_38028,N_37366,N_36971);
and U38029 (N_38029,N_37821,N_36488);
xnor U38030 (N_38030,N_36037,N_37100);
or U38031 (N_38031,N_37954,N_36482);
nor U38032 (N_38032,N_37623,N_37457);
nor U38033 (N_38033,N_37909,N_37207);
or U38034 (N_38034,N_37845,N_36701);
xor U38035 (N_38035,N_37364,N_36190);
nand U38036 (N_38036,N_37360,N_37680);
xnor U38037 (N_38037,N_36343,N_37948);
nor U38038 (N_38038,N_37002,N_36959);
and U38039 (N_38039,N_37867,N_36363);
xor U38040 (N_38040,N_37195,N_36765);
or U38041 (N_38041,N_36246,N_36924);
xnor U38042 (N_38042,N_36451,N_36874);
nor U38043 (N_38043,N_36172,N_36219);
nor U38044 (N_38044,N_37779,N_36792);
nand U38045 (N_38045,N_37442,N_36783);
nand U38046 (N_38046,N_36990,N_37521);
or U38047 (N_38047,N_37276,N_36589);
and U38048 (N_38048,N_36627,N_36158);
nand U38049 (N_38049,N_37905,N_37427);
nor U38050 (N_38050,N_36764,N_37423);
and U38051 (N_38051,N_37911,N_37304);
or U38052 (N_38052,N_36838,N_37847);
and U38053 (N_38053,N_36272,N_36602);
or U38054 (N_38054,N_36742,N_36041);
or U38055 (N_38055,N_37242,N_36603);
xnor U38056 (N_38056,N_36642,N_36392);
xnor U38057 (N_38057,N_36975,N_37203);
and U38058 (N_38058,N_36598,N_37184);
nand U38059 (N_38059,N_37239,N_37603);
or U38060 (N_38060,N_37702,N_37332);
xnor U38061 (N_38061,N_37835,N_36773);
nor U38062 (N_38062,N_37856,N_36699);
nand U38063 (N_38063,N_36502,N_37923);
nor U38064 (N_38064,N_37143,N_36835);
nand U38065 (N_38065,N_37894,N_37172);
nand U38066 (N_38066,N_36152,N_36795);
nand U38067 (N_38067,N_36031,N_36143);
or U38068 (N_38068,N_37716,N_36105);
xor U38069 (N_38069,N_37083,N_36605);
and U38070 (N_38070,N_36386,N_37641);
nor U38071 (N_38071,N_36974,N_37336);
nand U38072 (N_38072,N_37975,N_36336);
and U38073 (N_38073,N_37474,N_37430);
and U38074 (N_38074,N_36584,N_37984);
nand U38075 (N_38075,N_37620,N_36113);
nand U38076 (N_38076,N_36122,N_36825);
nor U38077 (N_38077,N_37575,N_37587);
or U38078 (N_38078,N_36456,N_36442);
nand U38079 (N_38079,N_37168,N_37634);
xnor U38080 (N_38080,N_36922,N_36324);
and U38081 (N_38081,N_36993,N_36397);
or U38082 (N_38082,N_36030,N_37557);
xnor U38083 (N_38083,N_37135,N_36860);
xor U38084 (N_38084,N_36072,N_37260);
nor U38085 (N_38085,N_36820,N_36934);
nand U38086 (N_38086,N_37648,N_37114);
or U38087 (N_38087,N_36986,N_36720);
xor U38088 (N_38088,N_36221,N_36463);
nand U38089 (N_38089,N_37486,N_36455);
xor U38090 (N_38090,N_37055,N_37507);
nor U38091 (N_38091,N_36512,N_37349);
or U38092 (N_38092,N_36005,N_36716);
nand U38093 (N_38093,N_37979,N_37798);
nand U38094 (N_38094,N_37514,N_37050);
nand U38095 (N_38095,N_37773,N_36136);
or U38096 (N_38096,N_36557,N_37029);
or U38097 (N_38097,N_37109,N_37740);
nor U38098 (N_38098,N_36413,N_37660);
or U38099 (N_38099,N_36595,N_36779);
xor U38100 (N_38100,N_36123,N_37286);
xor U38101 (N_38101,N_36286,N_37469);
or U38102 (N_38102,N_37755,N_37551);
xor U38103 (N_38103,N_37283,N_37515);
nor U38104 (N_38104,N_37123,N_36138);
nor U38105 (N_38105,N_36307,N_36026);
and U38106 (N_38106,N_36093,N_36426);
nor U38107 (N_38107,N_37574,N_37056);
xor U38108 (N_38108,N_36529,N_36914);
and U38109 (N_38109,N_37189,N_36903);
and U38110 (N_38110,N_37542,N_37768);
or U38111 (N_38111,N_36878,N_36359);
nor U38112 (N_38112,N_37299,N_36427);
nand U38113 (N_38113,N_37137,N_37080);
and U38114 (N_38114,N_37043,N_37344);
nand U38115 (N_38115,N_36954,N_36962);
nor U38116 (N_38116,N_37625,N_37130);
or U38117 (N_38117,N_36991,N_37653);
nor U38118 (N_38118,N_36237,N_36090);
and U38119 (N_38119,N_36254,N_37916);
nor U38120 (N_38120,N_36917,N_37888);
nand U38121 (N_38121,N_37651,N_37464);
nor U38122 (N_38122,N_37085,N_36273);
xor U38123 (N_38123,N_37000,N_36200);
and U38124 (N_38124,N_37750,N_37690);
nand U38125 (N_38125,N_37782,N_36241);
nand U38126 (N_38126,N_37284,N_36331);
xor U38127 (N_38127,N_36395,N_37731);
nor U38128 (N_38128,N_36910,N_37506);
and U38129 (N_38129,N_36207,N_37554);
or U38130 (N_38130,N_36269,N_36592);
xor U38131 (N_38131,N_36414,N_37805);
or U38132 (N_38132,N_37776,N_36188);
and U38133 (N_38133,N_37853,N_36145);
and U38134 (N_38134,N_37637,N_37693);
xnor U38135 (N_38135,N_37222,N_37811);
nand U38136 (N_38136,N_36966,N_36201);
and U38137 (N_38137,N_37508,N_36416);
and U38138 (N_38138,N_36635,N_37035);
xor U38139 (N_38139,N_36407,N_37527);
nand U38140 (N_38140,N_36942,N_36466);
xor U38141 (N_38141,N_36788,N_37403);
nor U38142 (N_38142,N_37259,N_36024);
nor U38143 (N_38143,N_37616,N_37072);
or U38144 (N_38144,N_36186,N_36721);
and U38145 (N_38145,N_36362,N_36586);
xnor U38146 (N_38146,N_37495,N_37945);
nand U38147 (N_38147,N_37633,N_36869);
xnor U38148 (N_38148,N_37891,N_37529);
and U38149 (N_38149,N_36332,N_37558);
nor U38150 (N_38150,N_36761,N_36400);
xnor U38151 (N_38151,N_37268,N_37823);
or U38152 (N_38152,N_36728,N_37384);
or U38153 (N_38153,N_37180,N_36978);
nor U38154 (N_38154,N_36164,N_36571);
or U38155 (N_38155,N_37510,N_36384);
nor U38156 (N_38156,N_36429,N_36634);
xor U38157 (N_38157,N_36168,N_37272);
nor U38158 (N_38158,N_37339,N_36319);
nand U38159 (N_38159,N_36054,N_36238);
and U38160 (N_38160,N_36316,N_36387);
and U38161 (N_38161,N_36118,N_36926);
nand U38162 (N_38162,N_36098,N_36325);
xor U38163 (N_38163,N_36743,N_37233);
and U38164 (N_38164,N_36726,N_37482);
or U38165 (N_38165,N_37468,N_37411);
nand U38166 (N_38166,N_37194,N_36626);
or U38167 (N_38167,N_36089,N_36639);
or U38168 (N_38168,N_37580,N_37578);
xnor U38169 (N_38169,N_37864,N_36335);
or U38170 (N_38170,N_36941,N_36625);
xor U38171 (N_38171,N_36281,N_37090);
or U38172 (N_38172,N_37160,N_36255);
nor U38173 (N_38173,N_36579,N_37504);
or U38174 (N_38174,N_37273,N_37030);
or U38175 (N_38175,N_36045,N_36277);
nor U38176 (N_38176,N_37297,N_36330);
and U38177 (N_38177,N_37285,N_36722);
nand U38178 (N_38178,N_36566,N_37213);
xnor U38179 (N_38179,N_36001,N_37517);
xor U38180 (N_38180,N_36769,N_36983);
xor U38181 (N_38181,N_37157,N_36127);
nand U38182 (N_38182,N_36205,N_37372);
nor U38183 (N_38183,N_36929,N_37900);
or U38184 (N_38184,N_37324,N_37409);
nor U38185 (N_38185,N_36094,N_37009);
or U38186 (N_38186,N_37450,N_37813);
xnor U38187 (N_38187,N_36102,N_37115);
nor U38188 (N_38188,N_36656,N_37199);
nor U38189 (N_38189,N_37963,N_36252);
nand U38190 (N_38190,N_37765,N_36161);
nand U38191 (N_38191,N_37104,N_36620);
nor U38192 (N_38192,N_36554,N_37686);
nand U38193 (N_38193,N_36836,N_37590);
nor U38194 (N_38194,N_36467,N_36454);
nor U38195 (N_38195,N_37522,N_36802);
xnor U38196 (N_38196,N_37334,N_36863);
and U38197 (N_38197,N_37685,N_36636);
and U38198 (N_38198,N_36551,N_37576);
and U38199 (N_38199,N_37758,N_36474);
xor U38200 (N_38200,N_36961,N_37518);
or U38201 (N_38201,N_36412,N_36070);
nand U38202 (N_38202,N_37918,N_36774);
or U38203 (N_38203,N_36622,N_37669);
xnor U38204 (N_38204,N_37434,N_36778);
nor U38205 (N_38205,N_37860,N_37008);
xnor U38206 (N_38206,N_37628,N_37069);
and U38207 (N_38207,N_37235,N_36537);
nand U38208 (N_38208,N_36445,N_37593);
or U38209 (N_38209,N_36198,N_36854);
xnor U38210 (N_38210,N_36327,N_36453);
nor U38211 (N_38211,N_36898,N_36260);
xor U38212 (N_38212,N_37210,N_36766);
nor U38213 (N_38213,N_37244,N_36021);
nand U38214 (N_38214,N_36091,N_37246);
xnor U38215 (N_38215,N_36646,N_36691);
nand U38216 (N_38216,N_37155,N_36022);
or U38217 (N_38217,N_37599,N_36748);
or U38218 (N_38218,N_36768,N_36837);
nand U38219 (N_38219,N_37441,N_37020);
xnor U38220 (N_38220,N_37812,N_36298);
nand U38221 (N_38221,N_37145,N_36394);
and U38222 (N_38222,N_37126,N_36956);
and U38223 (N_38223,N_36399,N_36514);
nor U38224 (N_38224,N_37484,N_37255);
nand U38225 (N_38225,N_37226,N_37451);
or U38226 (N_38226,N_36358,N_36333);
xnor U38227 (N_38227,N_36457,N_37939);
nand U38228 (N_38228,N_36807,N_37256);
or U38229 (N_38229,N_36628,N_36723);
nor U38230 (N_38230,N_37022,N_36476);
or U38231 (N_38231,N_37121,N_37969);
and U38232 (N_38232,N_37602,N_36692);
and U38233 (N_38233,N_36717,N_37117);
nor U38234 (N_38234,N_36497,N_37579);
and U38235 (N_38235,N_37186,N_36321);
xnor U38236 (N_38236,N_36234,N_37941);
nor U38237 (N_38237,N_36988,N_37828);
and U38238 (N_38238,N_36524,N_36657);
and U38239 (N_38239,N_36816,N_36496);
or U38240 (N_38240,N_36509,N_36310);
or U38241 (N_38241,N_37519,N_37146);
nor U38242 (N_38242,N_37262,N_36060);
xnor U38243 (N_38243,N_37307,N_36674);
xnor U38244 (N_38244,N_37858,N_37133);
and U38245 (N_38245,N_36431,N_37343);
nand U38246 (N_38246,N_37293,N_37443);
or U38247 (N_38247,N_36346,N_37566);
or U38248 (N_38248,N_37044,N_37591);
xnor U38249 (N_38249,N_36727,N_37532);
nor U38250 (N_38250,N_36075,N_37116);
or U38251 (N_38251,N_36248,N_37924);
or U38252 (N_38252,N_36032,N_37190);
nand U38253 (N_38253,N_36367,N_37490);
nor U38254 (N_38254,N_36977,N_37151);
nor U38255 (N_38255,N_36505,N_36369);
xor U38256 (N_38256,N_37747,N_36055);
nor U38257 (N_38257,N_36227,N_37325);
nand U38258 (N_38258,N_36087,N_36339);
nand U38259 (N_38259,N_37219,N_37980);
xnor U38260 (N_38260,N_37715,N_36401);
and U38261 (N_38261,N_36284,N_37730);
nand U38262 (N_38262,N_36420,N_36040);
nor U38263 (N_38263,N_37707,N_36443);
nor U38264 (N_38264,N_36419,N_36360);
or U38265 (N_38265,N_36980,N_37296);
and U38266 (N_38266,N_36334,N_37368);
nor U38267 (N_38267,N_37487,N_36553);
xor U38268 (N_38268,N_36705,N_36853);
nand U38269 (N_38269,N_37573,N_37752);
xor U38270 (N_38270,N_36713,N_37488);
nor U38271 (N_38271,N_37241,N_36673);
and U38272 (N_38272,N_37706,N_37799);
and U38273 (N_38273,N_36489,N_36029);
nand U38274 (N_38274,N_36121,N_36857);
and U38275 (N_38275,N_36963,N_36377);
or U38276 (N_38276,N_37800,N_36209);
or U38277 (N_38277,N_37668,N_36866);
or U38278 (N_38278,N_36671,N_37559);
xnor U38279 (N_38279,N_37319,N_36141);
and U38280 (N_38280,N_37406,N_36353);
and U38281 (N_38281,N_37027,N_36739);
xnor U38282 (N_38282,N_37895,N_36985);
or U38283 (N_38283,N_36880,N_37705);
or U38284 (N_38284,N_37738,N_36299);
nand U38285 (N_38285,N_36504,N_37141);
and U38286 (N_38286,N_36654,N_37717);
nand U38287 (N_38287,N_36789,N_36588);
and U38288 (N_38288,N_37049,N_36871);
nand U38289 (N_38289,N_36908,N_37250);
nor U38290 (N_38290,N_37661,N_36550);
nand U38291 (N_38291,N_37436,N_36043);
nor U38292 (N_38292,N_36314,N_36770);
nor U38293 (N_38293,N_36689,N_37187);
nor U38294 (N_38294,N_37962,N_37215);
or U38295 (N_38295,N_36696,N_36340);
nand U38296 (N_38296,N_36065,N_36902);
or U38297 (N_38297,N_37562,N_37251);
or U38298 (N_38298,N_36933,N_37321);
nand U38299 (N_38299,N_37694,N_37746);
or U38300 (N_38300,N_36895,N_37288);
xnor U38301 (N_38301,N_37087,N_37333);
nor U38302 (N_38302,N_36681,N_37066);
nand U38303 (N_38303,N_37081,N_37108);
nand U38304 (N_38304,N_36879,N_37756);
nand U38305 (N_38305,N_37868,N_36852);
nor U38306 (N_38306,N_37162,N_36428);
and U38307 (N_38307,N_37810,N_36710);
or U38308 (N_38308,N_36296,N_37363);
nand U38309 (N_38309,N_36841,N_37606);
nor U38310 (N_38310,N_36591,N_36736);
xnor U38311 (N_38311,N_36694,N_36301);
and U38312 (N_38312,N_36561,N_37809);
nor U38313 (N_38313,N_36932,N_37408);
nor U38314 (N_38314,N_37645,N_37549);
xor U38315 (N_38315,N_37405,N_37615);
or U38316 (N_38316,N_36452,N_37445);
nor U38317 (N_38317,N_37401,N_37785);
or U38318 (N_38318,N_37604,N_36848);
or U38319 (N_38319,N_36892,N_36655);
xor U38320 (N_38320,N_36746,N_36305);
and U38321 (N_38321,N_37552,N_37470);
xnor U38322 (N_38322,N_37791,N_37940);
or U38323 (N_38323,N_37511,N_36703);
nor U38324 (N_38324,N_36434,N_37624);
nand U38325 (N_38325,N_36011,N_36672);
and U38326 (N_38326,N_36485,N_36599);
or U38327 (N_38327,N_36160,N_36601);
xor U38328 (N_38328,N_37600,N_37388);
xor U38329 (N_38329,N_36994,N_37136);
and U38330 (N_38330,N_37166,N_37974);
nand U38331 (N_38331,N_37410,N_37889);
nor U38332 (N_38332,N_36149,N_36751);
nor U38333 (N_38333,N_36490,N_37666);
xnor U38334 (N_38334,N_37238,N_37499);
or U38335 (N_38335,N_37833,N_37429);
xnor U38336 (N_38336,N_37958,N_37509);
and U38337 (N_38337,N_36230,N_36028);
nand U38338 (N_38338,N_36583,N_37440);
nor U38339 (N_38339,N_37582,N_37539);
nand U38340 (N_38340,N_37097,N_36465);
and U38341 (N_38341,N_36424,N_37149);
or U38342 (N_38342,N_36432,N_37424);
nor U38343 (N_38343,N_37840,N_37067);
nand U38344 (N_38344,N_37311,N_36540);
nor U38345 (N_38345,N_37901,N_37844);
or U38346 (N_38346,N_36618,N_37959);
xnor U38347 (N_38347,N_37640,N_36249);
and U38348 (N_38348,N_37672,N_36955);
nand U38349 (N_38349,N_36015,N_36745);
nor U38350 (N_38350,N_36725,N_37883);
or U38351 (N_38351,N_36818,N_37169);
or U38352 (N_38352,N_37881,N_37524);
nor U38353 (N_38353,N_37419,N_37245);
nor U38354 (N_38354,N_37535,N_36006);
nand U38355 (N_38355,N_36192,N_37647);
xnor U38356 (N_38356,N_36698,N_37998);
nor U38357 (N_38357,N_36515,N_36663);
nand U38358 (N_38358,N_37842,N_37387);
or U38359 (N_38359,N_37389,N_36337);
nor U38360 (N_38360,N_36132,N_36704);
xnor U38361 (N_38361,N_36763,N_36992);
and U38362 (N_38362,N_37614,N_36365);
nor U38363 (N_38363,N_36831,N_37556);
nor U38364 (N_38364,N_36025,N_36714);
xnor U38365 (N_38365,N_36501,N_37721);
or U38366 (N_38366,N_37362,N_37064);
nor U38367 (N_38367,N_37546,N_36947);
nor U38368 (N_38368,N_37896,N_37699);
xor U38369 (N_38369,N_36827,N_36750);
nand U38370 (N_38370,N_36350,N_37113);
nand U38371 (N_38371,N_37253,N_36265);
nor U38372 (N_38372,N_36128,N_37063);
or U38373 (N_38373,N_37357,N_37091);
xnor U38374 (N_38374,N_37985,N_37692);
xor U38375 (N_38375,N_36076,N_37956);
nor U38376 (N_38376,N_37161,N_36056);
and U38377 (N_38377,N_37502,N_37052);
or U38378 (N_38378,N_36410,N_36872);
nor U38379 (N_38379,N_36843,N_36661);
nor U38380 (N_38380,N_36938,N_37264);
nor U38381 (N_38381,N_36526,N_37897);
xnor U38382 (N_38382,N_36907,N_37903);
xor U38383 (N_38383,N_37735,N_37743);
nand U38384 (N_38384,N_37447,N_37536);
nor U38385 (N_38385,N_36315,N_37836);
xnor U38386 (N_38386,N_37492,N_37681);
nor U38387 (N_38387,N_37684,N_36111);
xor U38388 (N_38388,N_37310,N_37089);
or U38389 (N_38389,N_37820,N_36737);
and U38390 (N_38390,N_36832,N_36295);
and U38391 (N_38391,N_37209,N_37071);
and U38392 (N_38392,N_36930,N_36999);
nor U38393 (N_38393,N_36533,N_37435);
xor U38394 (N_38394,N_37316,N_36215);
nor U38395 (N_38395,N_37088,N_37218);
xnor U38396 (N_38396,N_37892,N_36349);
and U38397 (N_38397,N_36050,N_37649);
and U38398 (N_38398,N_37178,N_36719);
xnor U38399 (N_38399,N_37134,N_37876);
and U38400 (N_38400,N_36899,N_36664);
nand U38401 (N_38401,N_37598,N_37402);
and U38402 (N_38402,N_37760,N_36063);
nand U38403 (N_38403,N_36347,N_37677);
xnor U38404 (N_38404,N_37884,N_36053);
nor U38405 (N_38405,N_36288,N_37555);
and U38406 (N_38406,N_36906,N_36855);
or U38407 (N_38407,N_36189,N_36256);
or U38408 (N_38408,N_37277,N_36797);
nor U38409 (N_38409,N_36126,N_36080);
nand U38410 (N_38410,N_36821,N_36066);
nand U38411 (N_38411,N_36357,N_37550);
nor U38412 (N_38412,N_37306,N_36450);
nand U38413 (N_38413,N_37950,N_36095);
and U38414 (N_38414,N_37105,N_36968);
nand U38415 (N_38415,N_36381,N_37483);
nor U38416 (N_38416,N_36049,N_36912);
and U38417 (N_38417,N_36306,N_36944);
nand U38418 (N_38418,N_36261,N_36199);
nand U38419 (N_38419,N_36312,N_37323);
xnor U38420 (N_38420,N_36730,N_37586);
nor U38421 (N_38421,N_36817,N_36590);
nand U38422 (N_38422,N_37202,N_36799);
xor U38423 (N_38423,N_36103,N_36612);
or U38424 (N_38424,N_36470,N_36928);
and U38425 (N_38425,N_36157,N_36208);
nand U38426 (N_38426,N_37300,N_37024);
and U38427 (N_38427,N_37214,N_37947);
nand U38428 (N_38428,N_36970,N_37869);
xnor U38429 (N_38429,N_36709,N_37709);
or U38430 (N_38430,N_37094,N_37619);
xor U38431 (N_38431,N_36004,N_36733);
or U38432 (N_38432,N_36931,N_37459);
or U38433 (N_38433,N_37118,N_36178);
and U38434 (N_38434,N_36293,N_37978);
or U38435 (N_38435,N_36425,N_37739);
or U38436 (N_38436,N_37762,N_37320);
nand U38437 (N_38437,N_36829,N_36014);
nor U38438 (N_38438,N_36421,N_36224);
nand U38439 (N_38439,N_37568,N_37972);
xor U38440 (N_38440,N_36345,N_37041);
nor U38441 (N_38441,N_36146,N_37843);
nand U38442 (N_38442,N_37046,N_36020);
or U38443 (N_38443,N_37997,N_37103);
nand U38444 (N_38444,N_36997,N_36275);
and U38445 (N_38445,N_37386,N_37417);
or U38446 (N_38446,N_36685,N_36225);
and U38447 (N_38447,N_37912,N_37786);
xnor U38448 (N_38448,N_36798,N_36137);
or U38449 (N_38449,N_37970,N_37374);
xor U38450 (N_38450,N_36495,N_36616);
or U38451 (N_38451,N_37444,N_36973);
nor U38452 (N_38452,N_36744,N_37414);
and U38453 (N_38453,N_37356,N_37534);
nand U38454 (N_38454,N_37062,N_36251);
or U38455 (N_38455,N_37512,N_37953);
xnor U38456 (N_38456,N_36749,N_37494);
and U38457 (N_38457,N_36404,N_36389);
nor U38458 (N_38458,N_37862,N_37794);
nand U38459 (N_38459,N_37461,N_37951);
and U38460 (N_38460,N_37585,N_37352);
or U38461 (N_38461,N_36376,N_37872);
xnor U38462 (N_38462,N_36417,N_36244);
xnor U38463 (N_38463,N_36567,N_36184);
nor U38464 (N_38464,N_36088,N_37899);
or U38465 (N_38465,N_36562,N_37026);
nor U38466 (N_38466,N_36348,N_36245);
xnor U38467 (N_38467,N_37824,N_36558);
nor U38468 (N_38468,N_36061,N_36545);
xor U38469 (N_38469,N_36464,N_36271);
or U38470 (N_38470,N_37068,N_37584);
xnor U38471 (N_38471,N_37965,N_37560);
or U38472 (N_38472,N_37928,N_37446);
nor U38473 (N_38473,N_36896,N_36609);
nand U38474 (N_38474,N_36753,N_37926);
xor U38475 (N_38475,N_36845,N_36734);
nor U38476 (N_38476,N_36995,N_37154);
or U38477 (N_38477,N_36623,N_37211);
nor U38478 (N_38478,N_37432,N_36805);
nand U38479 (N_38479,N_36796,N_37175);
nand U38480 (N_38480,N_36163,N_37463);
xnor U38481 (N_38481,N_36173,N_37439);
and U38482 (N_38482,N_36731,N_36239);
nor U38483 (N_38483,N_37875,N_37770);
nand U38484 (N_38484,N_37825,N_37561);
xor U38485 (N_38485,N_37375,N_37932);
or U38486 (N_38486,N_37347,N_37057);
and U38487 (N_38487,N_37946,N_36338);
or U38488 (N_38488,N_37526,N_36461);
or U38489 (N_38489,N_37193,N_36707);
nand U38490 (N_38490,N_36697,N_36581);
xor U38491 (N_38491,N_36624,N_36702);
and U38492 (N_38492,N_37943,N_36864);
and U38493 (N_38493,N_37757,N_36242);
and U38494 (N_38494,N_37305,N_37221);
xor U38495 (N_38495,N_37132,N_36106);
xor U38496 (N_38496,N_37831,N_37093);
xnor U38497 (N_38497,N_36677,N_36940);
nor U38498 (N_38498,N_37348,N_36278);
nor U38499 (N_38499,N_37373,N_36822);
nand U38500 (N_38500,N_37048,N_37480);
or U38501 (N_38501,N_37110,N_37601);
xnor U38502 (N_38502,N_37744,N_37385);
nand U38503 (N_38503,N_36647,N_37720);
nor U38504 (N_38504,N_36965,N_37632);
and U38505 (N_38505,N_37496,N_37290);
nand U38506 (N_38506,N_37167,N_36660);
nor U38507 (N_38507,N_36150,N_37395);
nor U38508 (N_38508,N_37302,N_37719);
nand U38509 (N_38509,N_37431,N_36073);
and U38510 (N_38510,N_36180,N_36834);
nand U38511 (N_38511,N_36130,N_37503);
nand U38512 (N_38512,N_37010,N_37034);
or U38513 (N_38513,N_37201,N_37538);
nand U38514 (N_38514,N_36447,N_36481);
or U38515 (N_38515,N_37196,N_37882);
or U38516 (N_38516,N_37745,N_36285);
xnor U38517 (N_38517,N_36536,N_36574);
nor U38518 (N_38518,N_37129,N_36506);
nand U38519 (N_38519,N_36289,N_36738);
and U38520 (N_38520,N_37124,N_37379);
nor U38521 (N_38521,N_36806,N_36191);
nor U38522 (N_38522,N_37917,N_37675);
and U38523 (N_38523,N_36510,N_37077);
and U38524 (N_38524,N_36148,N_37500);
or U38525 (N_38525,N_36297,N_36396);
and U38526 (N_38526,N_36361,N_37177);
and U38527 (N_38527,N_36987,N_36840);
or U38528 (N_38528,N_37331,N_37631);
xnor U38529 (N_38529,N_36576,N_37231);
and U38530 (N_38530,N_36522,N_37569);
xor U38531 (N_38531,N_36368,N_36259);
nor U38532 (N_38532,N_36920,N_37778);
or U38533 (N_38533,N_36957,N_36523);
nand U38534 (N_38534,N_37695,N_36943);
nand U38535 (N_38535,N_37122,N_37983);
and U38536 (N_38536,N_37465,N_36166);
and U38537 (N_38537,N_36036,N_36606);
nor U38538 (N_38538,N_37878,N_36676);
nor U38539 (N_38539,N_36051,N_37764);
or U38540 (N_38540,N_36439,N_36290);
xor U38541 (N_38541,N_36174,N_37254);
or U38542 (N_38542,N_36679,N_37322);
nand U38543 (N_38543,N_36531,N_36116);
and U38544 (N_38544,N_36876,N_37942);
and U38545 (N_38545,N_36587,N_36409);
or U38546 (N_38546,N_37315,N_37934);
and U38547 (N_38547,N_37777,N_37748);
or U38548 (N_38548,N_36861,N_36964);
and U38549 (N_38549,N_36600,N_36378);
or U38550 (N_38550,N_37863,N_36155);
and U38551 (N_38551,N_36596,N_36939);
xnor U38552 (N_38552,N_37082,N_36218);
or U38553 (N_38553,N_36905,N_37275);
nand U38554 (N_38554,N_37006,N_36303);
nor U38555 (N_38555,N_37525,N_37854);
nand U38556 (N_38556,N_36862,N_37120);
nand U38557 (N_38557,N_36263,N_36617);
and U38558 (N_38558,N_36027,N_36700);
nor U38559 (N_38559,N_36989,N_37257);
and U38560 (N_38560,N_37084,N_36187);
and U38561 (N_38561,N_37544,N_36729);
xnor U38562 (N_38562,N_37040,N_37153);
or U38563 (N_38563,N_36354,N_36867);
or U38564 (N_38564,N_37564,N_36074);
or U38565 (N_38565,N_37548,N_36142);
xor U38566 (N_38566,N_37070,N_37643);
nor U38567 (N_38567,N_36494,N_36649);
and U38568 (N_38568,N_36067,N_37528);
xor U38569 (N_38569,N_37737,N_36276);
or U38570 (N_38570,N_36117,N_36478);
and U38571 (N_38571,N_37437,N_36326);
nand U38572 (N_38572,N_37837,N_37960);
xor U38573 (N_38573,N_37294,N_37350);
nor U38574 (N_38574,N_37271,N_37170);
nand U38575 (N_38575,N_36658,N_36909);
and U38576 (N_38576,N_36253,N_37880);
or U38577 (N_38577,N_37466,N_37381);
or U38578 (N_38578,N_36125,N_36740);
and U38579 (N_38579,N_36133,N_37493);
nor U38580 (N_38580,N_37994,N_37609);
xor U38581 (N_38581,N_37674,N_37354);
xnor U38582 (N_38582,N_37053,N_36621);
and U38583 (N_38583,N_36715,N_37295);
xor U38584 (N_38584,N_36527,N_37237);
xor U38585 (N_38585,N_37991,N_37023);
xnor U38586 (N_38586,N_37657,N_37838);
or U38587 (N_38587,N_36473,N_37138);
or U38588 (N_38588,N_37234,N_36508);
or U38589 (N_38589,N_37804,N_37981);
or U38590 (N_38590,N_37795,N_36950);
nand U38591 (N_38591,N_36270,N_36632);
nand U38592 (N_38592,N_36607,N_37563);
or U38593 (N_38593,N_36039,N_36544);
nor U38594 (N_38594,N_37472,N_37664);
or U38595 (N_38595,N_36197,N_37317);
nor U38596 (N_38596,N_36372,N_36758);
and U38597 (N_38597,N_36388,N_37313);
and U38598 (N_38598,N_37433,N_37626);
nor U38599 (N_38599,N_36107,N_37212);
nand U38600 (N_38600,N_36171,N_37783);
and U38601 (N_38601,N_36328,N_37583);
or U38602 (N_38602,N_37065,N_37061);
nor U38603 (N_38603,N_36684,N_36952);
or U38604 (N_38604,N_36294,N_37806);
nor U38605 (N_38605,N_36555,N_36801);
and U38606 (N_38606,N_36516,N_37228);
or U38607 (N_38607,N_37567,N_36493);
xnor U38608 (N_38608,N_37987,N_36223);
xnor U38609 (N_38609,N_37312,N_37318);
nor U38610 (N_38610,N_37176,N_36958);
and U38611 (N_38611,N_37874,N_36194);
nand U38612 (N_38612,N_36695,N_36366);
xnor U38613 (N_38613,N_37491,N_37204);
nor U38614 (N_38614,N_37734,N_36134);
xor U38615 (N_38615,N_36534,N_37540);
and U38616 (N_38616,N_37976,N_37298);
xnor U38617 (N_38617,N_37772,N_37086);
nor U38618 (N_38618,N_37781,N_37904);
or U38619 (N_38619,N_37890,N_37413);
nand U38620 (N_38620,N_37769,N_36058);
xor U38621 (N_38621,N_37042,N_37140);
nand U38622 (N_38622,N_37025,N_37826);
nor U38623 (N_38623,N_36786,N_36868);
and U38624 (N_38624,N_36889,N_36232);
nor U38625 (N_38625,N_37964,N_37125);
nand U38626 (N_38626,N_37111,N_37278);
nor U38627 (N_38627,N_37197,N_36147);
xnor U38628 (N_38628,N_37390,N_36984);
xnor U38629 (N_38629,N_37485,N_36809);
xnor U38630 (N_38630,N_36911,N_36231);
nor U38631 (N_38631,N_37229,N_37144);
or U38632 (N_38632,N_36034,N_36546);
and U38633 (N_38633,N_37473,N_37404);
or U38634 (N_38634,N_37047,N_36687);
or U38635 (N_38635,N_36195,N_37673);
nand U38636 (N_38636,N_37396,N_37400);
xnor U38637 (N_38637,N_37870,N_37037);
nand U38638 (N_38638,N_36267,N_37269);
xnor U38639 (N_38639,N_36131,N_37289);
nand U38640 (N_38640,N_36097,N_36391);
xnor U38641 (N_38641,N_36901,N_37280);
xor U38642 (N_38642,N_36448,N_37767);
xor U38643 (N_38643,N_37131,N_37497);
or U38644 (N_38644,N_36548,N_37642);
and U38645 (N_38645,N_36375,N_36945);
nand U38646 (N_38646,N_36780,N_36279);
xor U38647 (N_38647,N_37252,N_36541);
xnor U38648 (N_38648,N_36499,N_36904);
nor U38649 (N_38649,N_36057,N_36921);
nand U38650 (N_38650,N_36803,N_37179);
nor U38651 (N_38651,N_36078,N_37696);
and U38652 (N_38652,N_36491,N_37908);
nor U38653 (N_38653,N_37003,N_37188);
or U38654 (N_38654,N_37613,N_36385);
nand U38655 (N_38655,N_36615,N_36948);
xor U38656 (N_38656,N_36398,N_37452);
or U38657 (N_38657,N_36329,N_36532);
and U38658 (N_38658,N_36308,N_36865);
and U38659 (N_38659,N_36222,N_37028);
nor U38660 (N_38660,N_37652,N_36528);
xor U38661 (N_38661,N_37266,N_37793);
nor U38662 (N_38662,N_36519,N_36217);
or U38663 (N_38663,N_36309,N_37938);
nand U38664 (N_38664,N_37516,N_37292);
xor U38665 (N_38665,N_36850,N_37351);
nor U38666 (N_38666,N_36323,N_36678);
xnor U38667 (N_38667,N_36793,N_36582);
xnor U38668 (N_38668,N_36165,N_37107);
and U38669 (N_38669,N_36300,N_37700);
nand U38670 (N_38670,N_36167,N_37949);
nand U38671 (N_38671,N_37171,N_37438);
or U38672 (N_38672,N_36240,N_37914);
or U38673 (N_38673,N_36785,N_37887);
and U38674 (N_38674,N_36220,N_37687);
and U38675 (N_38675,N_36471,N_36355);
nor U38676 (N_38676,N_36408,N_36637);
xnor U38677 (N_38677,N_36787,N_37263);
nor U38678 (N_38678,N_36500,N_37852);
nand U38679 (N_38679,N_36170,N_37834);
nor U38680 (N_38680,N_36894,N_37724);
or U38681 (N_38681,N_36538,N_37416);
nand U38682 (N_38682,N_36479,N_36498);
nor U38683 (N_38683,N_37007,N_37425);
nor U38684 (N_38684,N_37930,N_37629);
nand U38685 (N_38685,N_36469,N_36951);
nand U38686 (N_38686,N_37697,N_37224);
nor U38687 (N_38687,N_36211,N_36569);
xor U38688 (N_38688,N_36374,N_36100);
xnor U38689 (N_38689,N_36341,N_37230);
nand U38690 (N_38690,N_37627,N_37365);
and U38691 (N_38691,N_36844,N_37032);
or U38692 (N_38692,N_36870,N_36086);
xnor U38693 (N_38693,N_37165,N_36046);
nand U38694 (N_38694,N_36884,N_37096);
nor U38695 (N_38695,N_37610,N_37337);
xnor U38696 (N_38696,N_37654,N_36342);
xnor U38697 (N_38697,N_36570,N_37547);
and U38698 (N_38698,N_36492,N_37012);
or U38699 (N_38699,N_36112,N_36613);
nor U38700 (N_38700,N_37973,N_37857);
and U38701 (N_38701,N_37581,N_36507);
xnor U38702 (N_38702,N_37751,N_36549);
and U38703 (N_38703,N_36668,N_37995);
xnor U38704 (N_38704,N_36830,N_37541);
nand U38705 (N_38705,N_37232,N_37454);
nand U38706 (N_38706,N_36437,N_37102);
and U38707 (N_38707,N_36585,N_36370);
xnor U38708 (N_38708,N_37992,N_36882);
xnor U38709 (N_38709,N_37345,N_36652);
or U38710 (N_38710,N_36210,N_36115);
nand U38711 (N_38711,N_36846,N_37058);
xnor U38712 (N_38712,N_37802,N_37955);
xnor U38713 (N_38713,N_37977,N_37163);
xnor U38714 (N_38714,N_36513,N_37019);
or U38715 (N_38715,N_37726,N_36009);
xnor U38716 (N_38716,N_37281,N_36176);
nand U38717 (N_38717,N_36972,N_37759);
xnor U38718 (N_38718,N_36214,N_37989);
and U38719 (N_38719,N_36851,N_37014);
nor U38720 (N_38720,N_37471,N_37075);
nand U38721 (N_38721,N_36651,N_36946);
xor U38722 (N_38722,N_37458,N_36169);
nor U38723 (N_38723,N_36756,N_36580);
and U38724 (N_38724,N_36712,N_37426);
nand U38725 (N_38725,N_37045,N_36762);
nor U38726 (N_38726,N_36311,N_36960);
nand U38727 (N_38727,N_36918,N_37993);
or U38728 (N_38728,N_37303,N_37192);
nand U38729 (N_38729,N_37832,N_36919);
nor U38730 (N_38730,N_36520,N_36274);
or U38731 (N_38731,N_37099,N_37489);
xor U38732 (N_38732,N_37152,N_37248);
nand U38733 (N_38733,N_36403,N_36564);
nand U38734 (N_38734,N_36120,N_37033);
nor U38735 (N_38735,N_37873,N_36282);
nor U38736 (N_38736,N_37966,N_37523);
or U38737 (N_38737,N_37279,N_36643);
and U38738 (N_38738,N_37208,N_37016);
xor U38739 (N_38739,N_37412,N_37787);
and U38740 (N_38740,N_36008,N_36648);
nand U38741 (N_38741,N_36487,N_36925);
or U38742 (N_38742,N_36824,N_37592);
xnor U38743 (N_38743,N_36542,N_37005);
or U38744 (N_38744,N_36814,N_36760);
xor U38745 (N_38745,N_36291,N_36815);
nand U38746 (N_38746,N_37861,N_37462);
and U38747 (N_38747,N_37150,N_36129);
xor U38748 (N_38748,N_36665,N_37944);
or U38749 (N_38749,N_36976,N_36826);
xnor U38750 (N_38750,N_37198,N_37236);
and U38751 (N_38751,N_37646,N_36156);
and U38752 (N_38752,N_37682,N_37846);
and U38753 (N_38753,N_36042,N_37383);
xnor U38754 (N_38754,N_37788,N_37565);
nor U38755 (N_38755,N_37689,N_37183);
nand U38756 (N_38756,N_36423,N_36402);
nor U38757 (N_38757,N_36644,N_37421);
and U38758 (N_38758,N_36371,N_37608);
nand U38759 (N_38759,N_37839,N_36153);
nand U38760 (N_38760,N_36873,N_37013);
nor U38761 (N_38761,N_36486,N_37644);
and U38762 (N_38762,N_37418,N_37467);
xor U38763 (N_38763,N_37327,N_36044);
and U38764 (N_38764,N_37505,N_36085);
or U38765 (N_38765,N_36823,N_37849);
xnor U38766 (N_38766,N_36560,N_37358);
and U38767 (N_38767,N_37340,N_37807);
nand U38768 (N_38768,N_36079,N_37927);
nor U38769 (N_38769,N_37611,N_37101);
and U38770 (N_38770,N_37698,N_37808);
and U38771 (N_38771,N_37448,N_37936);
and U38772 (N_38772,N_36236,N_36669);
and U38773 (N_38773,N_37147,N_36283);
nor U38774 (N_38774,N_37671,N_37370);
nand U38775 (N_38775,N_37530,N_36518);
xor U38776 (N_38776,N_36099,N_37031);
xor U38777 (N_38777,N_37498,N_37701);
nor U38778 (N_38778,N_37815,N_36182);
nor U38779 (N_38779,N_37754,N_37217);
nand U38780 (N_38780,N_37971,N_37572);
nand U38781 (N_38781,N_37827,N_36257);
and U38782 (N_38782,N_37915,N_37796);
or U38783 (N_38783,N_36666,N_36578);
or U38784 (N_38784,N_37618,N_36318);
nor U38785 (N_38785,N_37801,N_36547);
or U38786 (N_38786,N_36650,N_36477);
or U38787 (N_38787,N_36781,N_37722);
and U38788 (N_38788,N_36183,N_36052);
or U38789 (N_38789,N_36619,N_36317);
xor U38790 (N_38790,N_37220,N_37341);
nand U38791 (N_38791,N_36411,N_37249);
or U38792 (N_38792,N_37392,N_37329);
xnor U38793 (N_38793,N_37453,N_36446);
and U38794 (N_38794,N_37545,N_37382);
or U38795 (N_38795,N_36287,N_37173);
or U38796 (N_38796,N_37309,N_36135);
nand U38797 (N_38797,N_37011,N_37240);
and U38798 (N_38798,N_36953,N_36877);
nor U38799 (N_38799,N_37703,N_36247);
nand U38800 (N_38800,N_36483,N_36268);
or U38801 (N_38801,N_37605,N_36196);
nor U38802 (N_38802,N_36811,N_36572);
nor U38803 (N_38803,N_36693,N_36304);
or U38804 (N_38804,N_36682,N_36144);
and U38805 (N_38805,N_36264,N_36262);
nor U38806 (N_38806,N_37741,N_37346);
nand U38807 (N_38807,N_36556,N_37919);
nor U38808 (N_38808,N_37723,N_36104);
nand U38809 (N_38809,N_36804,N_37021);
and U38810 (N_38810,N_37369,N_37397);
nor U38811 (N_38811,N_37159,N_37659);
nand U38812 (N_38812,N_37399,N_37079);
xnor U38813 (N_38813,N_37655,N_36351);
or U38814 (N_38814,N_36708,N_37865);
nor U38815 (N_38815,N_37185,N_36662);
and U38816 (N_38816,N_37371,N_37898);
nor U38817 (N_38817,N_37879,N_37921);
or U38818 (N_38818,N_36202,N_37906);
nand U38819 (N_38819,N_36048,N_37713);
nor U38820 (N_38820,N_37907,N_36982);
or U38821 (N_38821,N_37910,N_37330);
xnor U38822 (N_38822,N_36390,N_36010);
xnor U38823 (N_38823,N_37004,N_36382);
xnor U38824 (N_38824,N_37216,N_36435);
xnor U38825 (N_38825,N_37933,N_37790);
nor U38826 (N_38826,N_37073,N_37597);
nor U38827 (N_38827,N_37479,N_36688);
xor U38828 (N_38828,N_37570,N_36002);
nand U38829 (N_38829,N_37763,N_37380);
or U38830 (N_38830,N_37859,N_36969);
and U38831 (N_38831,N_36593,N_37886);
xnor U38832 (N_38832,N_36352,N_37017);
and U38833 (N_38833,N_36441,N_37543);
and U38834 (N_38834,N_36575,N_37267);
xor U38835 (N_38835,N_36813,N_37456);
xnor U38836 (N_38836,N_36344,N_36068);
or U38837 (N_38837,N_36559,N_36140);
and U38838 (N_38838,N_37261,N_36228);
and U38839 (N_38839,N_36110,N_36849);
xnor U38840 (N_38840,N_36364,N_37986);
and U38841 (N_38841,N_36383,N_36280);
xor U38842 (N_38842,N_36777,N_36013);
or U38843 (N_38843,N_37501,N_37714);
nand U38844 (N_38844,N_36886,N_36440);
and U38845 (N_38845,N_36109,N_36181);
xor U38846 (N_38846,N_37710,N_37513);
or U38847 (N_38847,N_37935,N_36071);
or U38848 (N_38848,N_37182,N_36393);
xnor U38849 (N_38849,N_37520,N_36468);
and U38850 (N_38850,N_36083,N_37191);
xor U38851 (N_38851,N_36858,N_37156);
nor U38852 (N_38852,N_36062,N_36082);
xnor U38853 (N_38853,N_37174,N_36233);
nand U38854 (N_38854,N_37996,N_36243);
xor U38855 (N_38855,N_37635,N_36449);
and U38856 (N_38856,N_37393,N_36923);
nand U38857 (N_38857,N_36690,N_37074);
nor U38858 (N_38858,N_37662,N_37227);
xor U38859 (N_38859,N_37622,N_37533);
xnor U38860 (N_38860,N_36356,N_37732);
nor U38861 (N_38861,N_36373,N_36462);
nor U38862 (N_38862,N_37128,N_37422);
and U38863 (N_38863,N_37481,N_36935);
nand U38864 (N_38864,N_36302,N_37774);
or U38865 (N_38865,N_37537,N_37929);
and U38866 (N_38866,N_37531,N_37766);
nor U38867 (N_38867,N_37181,N_37999);
and U38868 (N_38868,N_36430,N_37617);
nand U38869 (N_38869,N_36521,N_36900);
or U38870 (N_38870,N_36000,N_36484);
nor U38871 (N_38871,N_36735,N_37098);
and U38872 (N_38872,N_36018,N_36003);
and U38873 (N_38873,N_36175,N_37394);
nor U38874 (N_38874,N_36151,N_37729);
or U38875 (N_38875,N_36405,N_37711);
and U38876 (N_38876,N_37206,N_37455);
or U38877 (N_38877,N_37988,N_37428);
or U38878 (N_38878,N_37595,N_37797);
or U38879 (N_38879,N_37718,N_36313);
nor U38880 (N_38880,N_37001,N_37391);
or U38881 (N_38881,N_36752,N_36023);
nor U38882 (N_38882,N_36154,N_36258);
and U38883 (N_38883,N_36767,N_36213);
and U38884 (N_38884,N_36927,N_36119);
nand U38885 (N_38885,N_36981,N_36683);
nor U38886 (N_38886,N_37018,N_36530);
nand U38887 (N_38887,N_37127,N_36064);
and U38888 (N_38888,N_37139,N_36667);
or U38889 (N_38889,N_36883,N_36979);
xnor U38890 (N_38890,N_36755,N_37478);
xnor U38891 (N_38891,N_37038,N_36577);
nor U38892 (N_38892,N_37076,N_37733);
nand U38893 (N_38893,N_37059,N_37420);
nand U38894 (N_38894,N_37670,N_36503);
nand U38895 (N_38895,N_36406,N_37314);
and U38896 (N_38896,N_36597,N_36511);
nor U38897 (N_38897,N_37789,N_36633);
and U38898 (N_38898,N_36800,N_37636);
xor U38899 (N_38899,N_37106,N_36897);
or U38900 (N_38900,N_37819,N_37223);
and U38901 (N_38901,N_37822,N_36019);
nand U38902 (N_38902,N_37078,N_36659);
or U38903 (N_38903,N_37850,N_36784);
or U38904 (N_38904,N_36881,N_37200);
xor U38905 (N_38905,N_37588,N_36937);
xnor U38906 (N_38906,N_36645,N_37342);
nor U38907 (N_38907,N_36819,N_36114);
xor U38908 (N_38908,N_36077,N_36790);
nor U38909 (N_38909,N_36859,N_36012);
xor U38910 (N_38910,N_36610,N_37338);
xnor U38911 (N_38911,N_37205,N_36771);
and U38912 (N_38912,N_36179,N_37359);
nor U38913 (N_38913,N_36380,N_37968);
and U38914 (N_38914,N_36724,N_37829);
or U38915 (N_38915,N_37679,N_36444);
nor U38916 (N_38916,N_36638,N_37112);
nor U38917 (N_38917,N_37784,N_36747);
and U38918 (N_38918,N_37967,N_36235);
and U38919 (N_38919,N_36711,N_36847);
xnor U38920 (N_38920,N_36016,N_36459);
nor U38921 (N_38921,N_37937,N_36436);
nand U38922 (N_38922,N_36885,N_36732);
nand U38923 (N_38923,N_36292,N_36611);
and U38924 (N_38924,N_36084,N_36565);
nand U38925 (N_38925,N_36680,N_36967);
nand U38926 (N_38926,N_37725,N_36568);
or U38927 (N_38927,N_37164,N_36833);
and U38928 (N_38928,N_36543,N_37816);
nor U38929 (N_38929,N_37398,N_36206);
and U38930 (N_38930,N_36017,N_37119);
or U38931 (N_38931,N_36458,N_37931);
and U38932 (N_38932,N_37727,N_36916);
nor U38933 (N_38933,N_37712,N_36092);
or U38934 (N_38934,N_36162,N_36839);
nor U38935 (N_38935,N_36320,N_36875);
nor U38936 (N_38936,N_36035,N_36890);
nor U38937 (N_38937,N_36266,N_36949);
or U38938 (N_38938,N_36535,N_37630);
nor U38939 (N_38939,N_37792,N_36706);
nor U38940 (N_38940,N_37704,N_36322);
or U38941 (N_38941,N_37577,N_37650);
and U38942 (N_38942,N_37335,N_36810);
nor U38943 (N_38943,N_37665,N_36124);
or U38944 (N_38944,N_37039,N_37367);
xnor U38945 (N_38945,N_37761,N_37952);
nor U38946 (N_38946,N_37658,N_36203);
and U38947 (N_38947,N_36159,N_36913);
nand U38948 (N_38948,N_37691,N_37054);
xnor U38949 (N_38949,N_36775,N_36204);
xor U38950 (N_38950,N_37848,N_37708);
nor U38951 (N_38951,N_37301,N_37460);
nor U38952 (N_38952,N_36670,N_36998);
nor U38953 (N_38953,N_37688,N_36893);
or U38954 (N_38954,N_37667,N_37476);
and U38955 (N_38955,N_36996,N_36517);
xor U38956 (N_38956,N_36757,N_37621);
nand U38957 (N_38957,N_36038,N_37265);
nor U38958 (N_38958,N_36418,N_37818);
xnor U38959 (N_38959,N_37353,N_37589);
nor U38960 (N_38960,N_36641,N_37355);
nor U38961 (N_38961,N_36552,N_36741);
and U38962 (N_38962,N_36096,N_37922);
nor U38963 (N_38963,N_37841,N_36250);
nor U38964 (N_38964,N_36794,N_37594);
and U38965 (N_38965,N_36539,N_37866);
or U38966 (N_38966,N_36640,N_37683);
xnor U38967 (N_38967,N_36229,N_36047);
or U38968 (N_38968,N_37638,N_37326);
and U38969 (N_38969,N_37376,N_37361);
nor U38970 (N_38970,N_37678,N_36216);
or U38971 (N_38971,N_36782,N_37225);
nand U38972 (N_38972,N_37885,N_36460);
xnor U38973 (N_38973,N_36812,N_37639);
and U38974 (N_38974,N_37851,N_36475);
and U38975 (N_38975,N_37920,N_37913);
nor U38976 (N_38976,N_37060,N_36563);
nor U38977 (N_38977,N_36808,N_36101);
nand U38978 (N_38978,N_37415,N_37676);
and U38979 (N_38979,N_37771,N_36887);
nand U38980 (N_38980,N_37961,N_37990);
nand U38981 (N_38981,N_36185,N_37753);
xor U38982 (N_38982,N_37749,N_36614);
or U38983 (N_38983,N_36059,N_36415);
nand U38984 (N_38984,N_37736,N_36653);
nand U38985 (N_38985,N_36472,N_37902);
and U38986 (N_38986,N_36915,N_36891);
and U38987 (N_38987,N_36594,N_37893);
xor U38988 (N_38988,N_37925,N_37270);
xor U38989 (N_38989,N_36791,N_37036);
nor U38990 (N_38990,N_37553,N_37477);
or U38991 (N_38991,N_36631,N_36604);
xnor U38992 (N_38992,N_37871,N_37092);
or U38993 (N_38993,N_36226,N_36630);
and U38994 (N_38994,N_36422,N_36007);
and U38995 (N_38995,N_37775,N_36525);
nand U38996 (N_38996,N_37407,N_37243);
xor U38997 (N_38997,N_37274,N_36776);
nand U38998 (N_38998,N_37282,N_36480);
nor U38999 (N_38999,N_37158,N_37612);
nor U39000 (N_39000,N_37439,N_37201);
nor U39001 (N_39001,N_37546,N_37566);
or U39002 (N_39002,N_37925,N_36102);
xnor U39003 (N_39003,N_36377,N_37234);
xnor U39004 (N_39004,N_37407,N_37178);
nor U39005 (N_39005,N_36359,N_36397);
nand U39006 (N_39006,N_36649,N_37342);
nand U39007 (N_39007,N_37934,N_36473);
and U39008 (N_39008,N_36325,N_36488);
and U39009 (N_39009,N_37978,N_37452);
xnor U39010 (N_39010,N_37294,N_36695);
xnor U39011 (N_39011,N_37849,N_37730);
and U39012 (N_39012,N_36014,N_37601);
nand U39013 (N_39013,N_37368,N_37125);
and U39014 (N_39014,N_36255,N_36662);
nand U39015 (N_39015,N_37993,N_36650);
xor U39016 (N_39016,N_37702,N_37290);
and U39017 (N_39017,N_36616,N_36114);
xnor U39018 (N_39018,N_37071,N_37258);
xor U39019 (N_39019,N_37478,N_37138);
xnor U39020 (N_39020,N_37029,N_37351);
or U39021 (N_39021,N_36905,N_37983);
and U39022 (N_39022,N_36081,N_37755);
nor U39023 (N_39023,N_36374,N_36329);
nor U39024 (N_39024,N_37170,N_37228);
nand U39025 (N_39025,N_36466,N_36014);
and U39026 (N_39026,N_36175,N_36969);
nor U39027 (N_39027,N_36684,N_37675);
and U39028 (N_39028,N_37626,N_37228);
or U39029 (N_39029,N_36269,N_36865);
xor U39030 (N_39030,N_37020,N_37297);
xnor U39031 (N_39031,N_36549,N_36597);
nand U39032 (N_39032,N_37511,N_37157);
nand U39033 (N_39033,N_36614,N_36516);
or U39034 (N_39034,N_36059,N_37147);
nand U39035 (N_39035,N_36363,N_36653);
nand U39036 (N_39036,N_37659,N_36213);
xnor U39037 (N_39037,N_37791,N_37327);
and U39038 (N_39038,N_37857,N_36273);
and U39039 (N_39039,N_36775,N_36422);
or U39040 (N_39040,N_36774,N_36872);
or U39041 (N_39041,N_36040,N_36599);
and U39042 (N_39042,N_36848,N_36930);
and U39043 (N_39043,N_37756,N_37559);
or U39044 (N_39044,N_36648,N_37644);
and U39045 (N_39045,N_36035,N_37258);
nor U39046 (N_39046,N_36631,N_36230);
and U39047 (N_39047,N_36653,N_36519);
nand U39048 (N_39048,N_36981,N_37522);
or U39049 (N_39049,N_37781,N_36931);
nand U39050 (N_39050,N_36551,N_37855);
and U39051 (N_39051,N_37771,N_36924);
nand U39052 (N_39052,N_37030,N_36589);
nor U39053 (N_39053,N_36592,N_37561);
and U39054 (N_39054,N_36682,N_36945);
nand U39055 (N_39055,N_37358,N_37715);
nand U39056 (N_39056,N_36935,N_37240);
or U39057 (N_39057,N_36972,N_36271);
nand U39058 (N_39058,N_36493,N_37992);
nand U39059 (N_39059,N_37992,N_37033);
or U39060 (N_39060,N_36752,N_37889);
xnor U39061 (N_39061,N_36154,N_37282);
nand U39062 (N_39062,N_36904,N_37604);
nand U39063 (N_39063,N_37327,N_36207);
xor U39064 (N_39064,N_37594,N_37089);
and U39065 (N_39065,N_36924,N_36098);
nand U39066 (N_39066,N_36411,N_36913);
or U39067 (N_39067,N_36751,N_37427);
and U39068 (N_39068,N_37200,N_37506);
nand U39069 (N_39069,N_36906,N_36228);
xor U39070 (N_39070,N_36791,N_37976);
and U39071 (N_39071,N_37837,N_36686);
or U39072 (N_39072,N_36442,N_36700);
or U39073 (N_39073,N_37989,N_37099);
nand U39074 (N_39074,N_36304,N_36247);
nor U39075 (N_39075,N_36343,N_37680);
and U39076 (N_39076,N_36205,N_36324);
or U39077 (N_39077,N_37990,N_37056);
or U39078 (N_39078,N_37299,N_37820);
nand U39079 (N_39079,N_37226,N_36536);
nor U39080 (N_39080,N_37524,N_37615);
nor U39081 (N_39081,N_36325,N_36789);
nor U39082 (N_39082,N_37701,N_37195);
nor U39083 (N_39083,N_37644,N_36884);
or U39084 (N_39084,N_36707,N_37645);
nor U39085 (N_39085,N_37003,N_36364);
nor U39086 (N_39086,N_36401,N_37860);
or U39087 (N_39087,N_37281,N_37554);
and U39088 (N_39088,N_36004,N_36229);
nor U39089 (N_39089,N_37595,N_36268);
nor U39090 (N_39090,N_36923,N_36272);
nand U39091 (N_39091,N_37190,N_36650);
or U39092 (N_39092,N_37747,N_37208);
and U39093 (N_39093,N_37471,N_36020);
and U39094 (N_39094,N_37409,N_37674);
nand U39095 (N_39095,N_37421,N_37648);
or U39096 (N_39096,N_37605,N_37697);
nand U39097 (N_39097,N_36473,N_36274);
and U39098 (N_39098,N_37837,N_37948);
and U39099 (N_39099,N_37580,N_37844);
xor U39100 (N_39100,N_37322,N_37948);
xor U39101 (N_39101,N_36731,N_36065);
nor U39102 (N_39102,N_37794,N_37550);
or U39103 (N_39103,N_37928,N_36850);
xor U39104 (N_39104,N_37119,N_37100);
and U39105 (N_39105,N_36247,N_36136);
nand U39106 (N_39106,N_36458,N_37892);
nor U39107 (N_39107,N_37179,N_36407);
nor U39108 (N_39108,N_36372,N_36883);
and U39109 (N_39109,N_37789,N_37256);
nand U39110 (N_39110,N_37053,N_36036);
xor U39111 (N_39111,N_37243,N_37052);
nand U39112 (N_39112,N_37360,N_37351);
and U39113 (N_39113,N_37321,N_36159);
xnor U39114 (N_39114,N_36413,N_37690);
nor U39115 (N_39115,N_36399,N_36056);
xor U39116 (N_39116,N_36687,N_36091);
and U39117 (N_39117,N_36121,N_37654);
or U39118 (N_39118,N_37766,N_36291);
nand U39119 (N_39119,N_37343,N_37066);
or U39120 (N_39120,N_37168,N_37480);
and U39121 (N_39121,N_37980,N_36270);
xnor U39122 (N_39122,N_37405,N_36762);
nor U39123 (N_39123,N_36078,N_36270);
and U39124 (N_39124,N_36055,N_36022);
nand U39125 (N_39125,N_37124,N_37653);
nand U39126 (N_39126,N_36953,N_36003);
nor U39127 (N_39127,N_37325,N_36750);
or U39128 (N_39128,N_36395,N_36311);
nand U39129 (N_39129,N_36499,N_36752);
and U39130 (N_39130,N_36006,N_37595);
nor U39131 (N_39131,N_36788,N_37622);
nor U39132 (N_39132,N_36011,N_37216);
nor U39133 (N_39133,N_37032,N_37905);
nor U39134 (N_39134,N_36373,N_37677);
xnor U39135 (N_39135,N_37591,N_37368);
nor U39136 (N_39136,N_37263,N_36635);
xor U39137 (N_39137,N_36333,N_37186);
nand U39138 (N_39138,N_36067,N_36743);
xor U39139 (N_39139,N_37113,N_37593);
xor U39140 (N_39140,N_37511,N_37979);
xnor U39141 (N_39141,N_37870,N_37130);
nand U39142 (N_39142,N_36256,N_36744);
xnor U39143 (N_39143,N_37581,N_37726);
and U39144 (N_39144,N_36021,N_36441);
xnor U39145 (N_39145,N_36654,N_37921);
xnor U39146 (N_39146,N_37043,N_36313);
nand U39147 (N_39147,N_36370,N_37956);
and U39148 (N_39148,N_37721,N_36076);
xnor U39149 (N_39149,N_36195,N_36374);
and U39150 (N_39150,N_36393,N_37517);
nor U39151 (N_39151,N_36596,N_37987);
nand U39152 (N_39152,N_36980,N_36774);
nor U39153 (N_39153,N_37771,N_37616);
xor U39154 (N_39154,N_36423,N_36462);
nand U39155 (N_39155,N_36981,N_36799);
and U39156 (N_39156,N_36008,N_37262);
xnor U39157 (N_39157,N_37819,N_36423);
and U39158 (N_39158,N_37968,N_37066);
and U39159 (N_39159,N_37987,N_36973);
and U39160 (N_39160,N_37490,N_37237);
xnor U39161 (N_39161,N_37762,N_36082);
or U39162 (N_39162,N_36905,N_37800);
nand U39163 (N_39163,N_36070,N_36199);
nor U39164 (N_39164,N_36991,N_37284);
nand U39165 (N_39165,N_36422,N_36783);
nor U39166 (N_39166,N_36470,N_37829);
nand U39167 (N_39167,N_36719,N_37798);
nor U39168 (N_39168,N_36539,N_37605);
nand U39169 (N_39169,N_37452,N_37244);
nand U39170 (N_39170,N_37321,N_37082);
and U39171 (N_39171,N_36659,N_36148);
nor U39172 (N_39172,N_36538,N_36124);
xor U39173 (N_39173,N_36457,N_37227);
xnor U39174 (N_39174,N_37654,N_37419);
nor U39175 (N_39175,N_36349,N_36172);
or U39176 (N_39176,N_36757,N_37468);
xnor U39177 (N_39177,N_37245,N_36136);
nand U39178 (N_39178,N_36851,N_36317);
nor U39179 (N_39179,N_36868,N_37885);
nand U39180 (N_39180,N_36231,N_36864);
nor U39181 (N_39181,N_37714,N_37907);
xor U39182 (N_39182,N_36113,N_36740);
xnor U39183 (N_39183,N_37420,N_36322);
and U39184 (N_39184,N_37281,N_36836);
nand U39185 (N_39185,N_37460,N_37752);
or U39186 (N_39186,N_36389,N_36678);
nor U39187 (N_39187,N_37693,N_36274);
xor U39188 (N_39188,N_37661,N_36584);
or U39189 (N_39189,N_36263,N_36450);
nand U39190 (N_39190,N_37926,N_36990);
nand U39191 (N_39191,N_36484,N_37041);
and U39192 (N_39192,N_37819,N_37211);
and U39193 (N_39193,N_37502,N_37559);
or U39194 (N_39194,N_36176,N_37433);
nand U39195 (N_39195,N_36243,N_37642);
xnor U39196 (N_39196,N_36873,N_36521);
or U39197 (N_39197,N_36579,N_37658);
nand U39198 (N_39198,N_36290,N_37445);
nor U39199 (N_39199,N_36815,N_37890);
and U39200 (N_39200,N_37940,N_36849);
or U39201 (N_39201,N_36377,N_36149);
nor U39202 (N_39202,N_36922,N_37840);
nand U39203 (N_39203,N_37473,N_36453);
nor U39204 (N_39204,N_37361,N_37136);
and U39205 (N_39205,N_37197,N_36983);
nand U39206 (N_39206,N_36005,N_37217);
or U39207 (N_39207,N_36582,N_37096);
xnor U39208 (N_39208,N_36352,N_37889);
and U39209 (N_39209,N_37499,N_36048);
and U39210 (N_39210,N_37997,N_37100);
and U39211 (N_39211,N_37225,N_36801);
nand U39212 (N_39212,N_37505,N_37470);
or U39213 (N_39213,N_37897,N_37208);
nor U39214 (N_39214,N_37434,N_37584);
and U39215 (N_39215,N_36297,N_36739);
nor U39216 (N_39216,N_37256,N_37058);
or U39217 (N_39217,N_36527,N_36275);
and U39218 (N_39218,N_36013,N_37068);
nor U39219 (N_39219,N_36609,N_36300);
and U39220 (N_39220,N_37944,N_37966);
or U39221 (N_39221,N_36584,N_36786);
or U39222 (N_39222,N_37704,N_37771);
xor U39223 (N_39223,N_36734,N_37253);
nor U39224 (N_39224,N_36308,N_36734);
nand U39225 (N_39225,N_37001,N_37506);
xor U39226 (N_39226,N_36105,N_37326);
nand U39227 (N_39227,N_37316,N_36723);
xor U39228 (N_39228,N_37657,N_37006);
nand U39229 (N_39229,N_36295,N_37093);
nor U39230 (N_39230,N_36632,N_37381);
xor U39231 (N_39231,N_36120,N_36338);
and U39232 (N_39232,N_37147,N_37290);
nor U39233 (N_39233,N_37686,N_36124);
xnor U39234 (N_39234,N_36718,N_36211);
or U39235 (N_39235,N_36043,N_37772);
nor U39236 (N_39236,N_37217,N_36384);
and U39237 (N_39237,N_37561,N_37632);
nand U39238 (N_39238,N_36347,N_37741);
xnor U39239 (N_39239,N_37402,N_36721);
nand U39240 (N_39240,N_36467,N_37880);
and U39241 (N_39241,N_36323,N_37250);
or U39242 (N_39242,N_36597,N_37673);
and U39243 (N_39243,N_36351,N_37917);
or U39244 (N_39244,N_37554,N_36407);
nor U39245 (N_39245,N_37574,N_37306);
and U39246 (N_39246,N_37168,N_36646);
nor U39247 (N_39247,N_36373,N_37623);
nand U39248 (N_39248,N_36476,N_36036);
or U39249 (N_39249,N_37251,N_36308);
and U39250 (N_39250,N_36592,N_37903);
nand U39251 (N_39251,N_36755,N_36872);
nand U39252 (N_39252,N_36277,N_36152);
nor U39253 (N_39253,N_36548,N_36088);
nand U39254 (N_39254,N_36370,N_36060);
and U39255 (N_39255,N_36878,N_36512);
and U39256 (N_39256,N_37411,N_37426);
and U39257 (N_39257,N_37274,N_36504);
and U39258 (N_39258,N_36495,N_36818);
nand U39259 (N_39259,N_36476,N_36969);
nand U39260 (N_39260,N_36329,N_37177);
and U39261 (N_39261,N_36543,N_36535);
xor U39262 (N_39262,N_37499,N_36404);
and U39263 (N_39263,N_37441,N_37469);
nor U39264 (N_39264,N_37065,N_37640);
nand U39265 (N_39265,N_36856,N_37070);
nor U39266 (N_39266,N_37044,N_36224);
nand U39267 (N_39267,N_37808,N_37653);
and U39268 (N_39268,N_37975,N_36453);
and U39269 (N_39269,N_36019,N_36961);
and U39270 (N_39270,N_36266,N_37786);
nand U39271 (N_39271,N_37323,N_37566);
nor U39272 (N_39272,N_36860,N_37714);
xnor U39273 (N_39273,N_36494,N_36098);
nor U39274 (N_39274,N_36866,N_36167);
or U39275 (N_39275,N_37582,N_36057);
nor U39276 (N_39276,N_37997,N_36210);
or U39277 (N_39277,N_37122,N_37678);
nor U39278 (N_39278,N_37561,N_37526);
or U39279 (N_39279,N_37248,N_36909);
and U39280 (N_39280,N_37800,N_36706);
nand U39281 (N_39281,N_37569,N_37842);
or U39282 (N_39282,N_37769,N_37579);
nand U39283 (N_39283,N_37894,N_36670);
xnor U39284 (N_39284,N_36192,N_37872);
xor U39285 (N_39285,N_36758,N_37379);
nand U39286 (N_39286,N_36988,N_36253);
xor U39287 (N_39287,N_37422,N_37876);
xor U39288 (N_39288,N_36887,N_37647);
or U39289 (N_39289,N_37128,N_36629);
and U39290 (N_39290,N_36780,N_37527);
nor U39291 (N_39291,N_37919,N_36650);
xnor U39292 (N_39292,N_36240,N_37220);
and U39293 (N_39293,N_36827,N_37197);
nand U39294 (N_39294,N_36699,N_36299);
and U39295 (N_39295,N_37699,N_36979);
xor U39296 (N_39296,N_36239,N_36177);
xor U39297 (N_39297,N_36896,N_37292);
and U39298 (N_39298,N_37301,N_37033);
and U39299 (N_39299,N_36346,N_36393);
xnor U39300 (N_39300,N_36243,N_36574);
or U39301 (N_39301,N_36910,N_37324);
nand U39302 (N_39302,N_36082,N_37826);
or U39303 (N_39303,N_36715,N_37974);
xor U39304 (N_39304,N_36817,N_37200);
nor U39305 (N_39305,N_37682,N_37716);
or U39306 (N_39306,N_37599,N_36243);
and U39307 (N_39307,N_37199,N_36072);
or U39308 (N_39308,N_37566,N_36009);
or U39309 (N_39309,N_36145,N_37026);
nand U39310 (N_39310,N_37251,N_36028);
nor U39311 (N_39311,N_37769,N_37524);
nand U39312 (N_39312,N_37307,N_37078);
nor U39313 (N_39313,N_37104,N_36545);
xor U39314 (N_39314,N_37354,N_36592);
nand U39315 (N_39315,N_36683,N_36611);
nor U39316 (N_39316,N_36600,N_37796);
or U39317 (N_39317,N_36636,N_37612);
xnor U39318 (N_39318,N_36973,N_36261);
nor U39319 (N_39319,N_36329,N_36411);
and U39320 (N_39320,N_37597,N_37676);
nor U39321 (N_39321,N_36948,N_37884);
or U39322 (N_39322,N_37089,N_37618);
or U39323 (N_39323,N_36074,N_37763);
xnor U39324 (N_39324,N_36626,N_36324);
nand U39325 (N_39325,N_37710,N_37988);
or U39326 (N_39326,N_37264,N_36167);
xor U39327 (N_39327,N_37132,N_36304);
and U39328 (N_39328,N_37458,N_37779);
xnor U39329 (N_39329,N_37075,N_36485);
nand U39330 (N_39330,N_36008,N_36354);
and U39331 (N_39331,N_36244,N_36897);
xor U39332 (N_39332,N_36273,N_37395);
and U39333 (N_39333,N_37158,N_37271);
or U39334 (N_39334,N_36483,N_36879);
nor U39335 (N_39335,N_37982,N_37008);
xnor U39336 (N_39336,N_37692,N_37605);
nand U39337 (N_39337,N_36201,N_36912);
nand U39338 (N_39338,N_37133,N_37615);
or U39339 (N_39339,N_36494,N_36804);
nor U39340 (N_39340,N_36295,N_37821);
nand U39341 (N_39341,N_36890,N_36983);
nand U39342 (N_39342,N_37268,N_37273);
nand U39343 (N_39343,N_36134,N_36966);
nand U39344 (N_39344,N_37612,N_36134);
and U39345 (N_39345,N_37455,N_36942);
xnor U39346 (N_39346,N_37072,N_36565);
nand U39347 (N_39347,N_36581,N_36474);
xor U39348 (N_39348,N_36635,N_37500);
and U39349 (N_39349,N_37958,N_36693);
xnor U39350 (N_39350,N_36835,N_37693);
or U39351 (N_39351,N_36019,N_37975);
and U39352 (N_39352,N_37967,N_36339);
nand U39353 (N_39353,N_36754,N_37799);
nor U39354 (N_39354,N_36325,N_36465);
nand U39355 (N_39355,N_37990,N_37443);
nor U39356 (N_39356,N_36811,N_37198);
xor U39357 (N_39357,N_37071,N_37260);
and U39358 (N_39358,N_36517,N_37520);
and U39359 (N_39359,N_37689,N_37027);
or U39360 (N_39360,N_37671,N_37394);
nand U39361 (N_39361,N_37856,N_37316);
xor U39362 (N_39362,N_37978,N_37624);
and U39363 (N_39363,N_37276,N_37782);
and U39364 (N_39364,N_37820,N_37535);
xnor U39365 (N_39365,N_37795,N_36378);
nor U39366 (N_39366,N_36557,N_36429);
or U39367 (N_39367,N_36884,N_36120);
or U39368 (N_39368,N_37731,N_36457);
xnor U39369 (N_39369,N_37511,N_37480);
and U39370 (N_39370,N_36949,N_37119);
nor U39371 (N_39371,N_36928,N_36252);
and U39372 (N_39372,N_36462,N_37627);
or U39373 (N_39373,N_37265,N_37309);
or U39374 (N_39374,N_37315,N_36731);
or U39375 (N_39375,N_37679,N_37885);
and U39376 (N_39376,N_36273,N_36568);
nor U39377 (N_39377,N_37604,N_37522);
or U39378 (N_39378,N_37374,N_36435);
nor U39379 (N_39379,N_37246,N_37176);
nor U39380 (N_39380,N_37480,N_36023);
nand U39381 (N_39381,N_37783,N_37291);
xnor U39382 (N_39382,N_37028,N_37854);
nand U39383 (N_39383,N_36698,N_36699);
nor U39384 (N_39384,N_36402,N_37838);
or U39385 (N_39385,N_36950,N_36791);
or U39386 (N_39386,N_37349,N_37042);
or U39387 (N_39387,N_37105,N_36485);
and U39388 (N_39388,N_37267,N_36925);
nor U39389 (N_39389,N_36257,N_37646);
or U39390 (N_39390,N_37314,N_37673);
or U39391 (N_39391,N_36379,N_37792);
or U39392 (N_39392,N_37969,N_36800);
nor U39393 (N_39393,N_36298,N_36852);
nor U39394 (N_39394,N_36005,N_36640);
or U39395 (N_39395,N_37397,N_37606);
nand U39396 (N_39396,N_36842,N_37907);
nor U39397 (N_39397,N_36354,N_36716);
nor U39398 (N_39398,N_37844,N_37053);
nand U39399 (N_39399,N_37248,N_37943);
nand U39400 (N_39400,N_37983,N_37592);
xor U39401 (N_39401,N_37461,N_36893);
nor U39402 (N_39402,N_36387,N_36784);
xor U39403 (N_39403,N_36527,N_36516);
or U39404 (N_39404,N_36314,N_37496);
and U39405 (N_39405,N_37195,N_37260);
or U39406 (N_39406,N_36483,N_37881);
nor U39407 (N_39407,N_36842,N_37838);
nand U39408 (N_39408,N_36253,N_36517);
nor U39409 (N_39409,N_36806,N_36906);
and U39410 (N_39410,N_36194,N_37489);
nor U39411 (N_39411,N_36735,N_37773);
nor U39412 (N_39412,N_37891,N_36210);
nor U39413 (N_39413,N_36735,N_37500);
xnor U39414 (N_39414,N_36704,N_36847);
and U39415 (N_39415,N_37761,N_37812);
and U39416 (N_39416,N_36101,N_36886);
or U39417 (N_39417,N_36789,N_37051);
or U39418 (N_39418,N_36359,N_36611);
nor U39419 (N_39419,N_36895,N_36384);
or U39420 (N_39420,N_36565,N_37446);
or U39421 (N_39421,N_36633,N_36763);
nor U39422 (N_39422,N_37175,N_37524);
xnor U39423 (N_39423,N_37009,N_37234);
nor U39424 (N_39424,N_37872,N_36712);
nand U39425 (N_39425,N_37441,N_36409);
nor U39426 (N_39426,N_37497,N_37409);
and U39427 (N_39427,N_36792,N_37842);
and U39428 (N_39428,N_37724,N_36057);
nand U39429 (N_39429,N_37602,N_36332);
nor U39430 (N_39430,N_37025,N_37474);
xor U39431 (N_39431,N_37242,N_36697);
nor U39432 (N_39432,N_37943,N_36983);
or U39433 (N_39433,N_37197,N_36664);
nand U39434 (N_39434,N_36282,N_37032);
or U39435 (N_39435,N_37450,N_37183);
xor U39436 (N_39436,N_37093,N_36874);
nor U39437 (N_39437,N_37176,N_36584);
or U39438 (N_39438,N_37347,N_36703);
xnor U39439 (N_39439,N_37231,N_36839);
nand U39440 (N_39440,N_36265,N_37390);
nand U39441 (N_39441,N_37721,N_36704);
and U39442 (N_39442,N_37355,N_37709);
nand U39443 (N_39443,N_36959,N_36183);
xor U39444 (N_39444,N_36939,N_37527);
or U39445 (N_39445,N_36025,N_36893);
xnor U39446 (N_39446,N_37163,N_37244);
xnor U39447 (N_39447,N_36703,N_36055);
and U39448 (N_39448,N_36806,N_37225);
and U39449 (N_39449,N_37460,N_36192);
or U39450 (N_39450,N_37111,N_36290);
nor U39451 (N_39451,N_36170,N_37853);
nor U39452 (N_39452,N_37813,N_36219);
nand U39453 (N_39453,N_36031,N_36569);
and U39454 (N_39454,N_36510,N_37413);
xnor U39455 (N_39455,N_37143,N_36748);
and U39456 (N_39456,N_37082,N_36105);
nor U39457 (N_39457,N_36911,N_37692);
and U39458 (N_39458,N_37814,N_36984);
or U39459 (N_39459,N_36514,N_36822);
and U39460 (N_39460,N_37389,N_36474);
or U39461 (N_39461,N_37296,N_36903);
or U39462 (N_39462,N_37306,N_36998);
nor U39463 (N_39463,N_36896,N_36151);
or U39464 (N_39464,N_37315,N_37943);
nor U39465 (N_39465,N_36906,N_37508);
or U39466 (N_39466,N_37176,N_37711);
nor U39467 (N_39467,N_37285,N_37564);
xnor U39468 (N_39468,N_37242,N_36407);
or U39469 (N_39469,N_36568,N_37444);
and U39470 (N_39470,N_37098,N_36053);
nand U39471 (N_39471,N_36956,N_36729);
and U39472 (N_39472,N_37157,N_37420);
nand U39473 (N_39473,N_36448,N_36269);
and U39474 (N_39474,N_37116,N_36953);
and U39475 (N_39475,N_36579,N_37853);
or U39476 (N_39476,N_37032,N_36840);
nand U39477 (N_39477,N_37224,N_37401);
xor U39478 (N_39478,N_36335,N_36440);
xnor U39479 (N_39479,N_37905,N_37172);
or U39480 (N_39480,N_36595,N_36777);
and U39481 (N_39481,N_36540,N_36477);
or U39482 (N_39482,N_36315,N_36650);
or U39483 (N_39483,N_37224,N_36594);
xnor U39484 (N_39484,N_36707,N_37223);
or U39485 (N_39485,N_37594,N_37543);
or U39486 (N_39486,N_36097,N_36260);
or U39487 (N_39487,N_36231,N_36783);
nand U39488 (N_39488,N_36983,N_36688);
nand U39489 (N_39489,N_36283,N_36866);
or U39490 (N_39490,N_36482,N_37114);
or U39491 (N_39491,N_37353,N_37516);
and U39492 (N_39492,N_36660,N_37061);
nor U39493 (N_39493,N_37221,N_37471);
nand U39494 (N_39494,N_36497,N_36623);
nand U39495 (N_39495,N_37083,N_36894);
or U39496 (N_39496,N_37714,N_37140);
nand U39497 (N_39497,N_36952,N_36985);
nand U39498 (N_39498,N_37977,N_36267);
or U39499 (N_39499,N_36907,N_37006);
or U39500 (N_39500,N_37345,N_36530);
nor U39501 (N_39501,N_37990,N_36516);
or U39502 (N_39502,N_37048,N_36137);
xor U39503 (N_39503,N_36689,N_37239);
nor U39504 (N_39504,N_37783,N_37755);
xnor U39505 (N_39505,N_37170,N_37549);
xnor U39506 (N_39506,N_37342,N_37321);
and U39507 (N_39507,N_37034,N_37264);
nor U39508 (N_39508,N_37883,N_37841);
and U39509 (N_39509,N_37588,N_36575);
xnor U39510 (N_39510,N_37720,N_36671);
and U39511 (N_39511,N_37723,N_37430);
and U39512 (N_39512,N_37546,N_37603);
or U39513 (N_39513,N_37981,N_36311);
xor U39514 (N_39514,N_36284,N_36411);
or U39515 (N_39515,N_37273,N_36423);
xnor U39516 (N_39516,N_36518,N_36531);
and U39517 (N_39517,N_37957,N_37552);
xor U39518 (N_39518,N_36796,N_36687);
nor U39519 (N_39519,N_37818,N_36336);
and U39520 (N_39520,N_36447,N_37875);
nand U39521 (N_39521,N_37127,N_36929);
xnor U39522 (N_39522,N_36605,N_37208);
nor U39523 (N_39523,N_36337,N_36637);
and U39524 (N_39524,N_36036,N_36621);
xnor U39525 (N_39525,N_37260,N_37111);
nor U39526 (N_39526,N_36431,N_37133);
xnor U39527 (N_39527,N_37270,N_37940);
nor U39528 (N_39528,N_36048,N_36779);
nand U39529 (N_39529,N_36727,N_36719);
xnor U39530 (N_39530,N_37112,N_37589);
xnor U39531 (N_39531,N_36022,N_37823);
nand U39532 (N_39532,N_37548,N_36947);
or U39533 (N_39533,N_37904,N_36770);
nor U39534 (N_39534,N_37479,N_36742);
or U39535 (N_39535,N_37482,N_37893);
and U39536 (N_39536,N_36921,N_36062);
or U39537 (N_39537,N_37868,N_36373);
and U39538 (N_39538,N_36566,N_36930);
nor U39539 (N_39539,N_37245,N_37692);
and U39540 (N_39540,N_36788,N_37052);
xor U39541 (N_39541,N_37200,N_36707);
nor U39542 (N_39542,N_37438,N_37127);
or U39543 (N_39543,N_36961,N_37695);
and U39544 (N_39544,N_36863,N_37035);
nand U39545 (N_39545,N_36783,N_37625);
nand U39546 (N_39546,N_36493,N_36789);
nand U39547 (N_39547,N_37244,N_36663);
xor U39548 (N_39548,N_36418,N_37875);
nand U39549 (N_39549,N_36291,N_37584);
or U39550 (N_39550,N_36439,N_36167);
nand U39551 (N_39551,N_36661,N_36718);
and U39552 (N_39552,N_36169,N_36377);
nand U39553 (N_39553,N_36456,N_37724);
nand U39554 (N_39554,N_37153,N_36553);
nand U39555 (N_39555,N_37597,N_37388);
or U39556 (N_39556,N_37510,N_37715);
and U39557 (N_39557,N_37031,N_36573);
or U39558 (N_39558,N_36082,N_37468);
and U39559 (N_39559,N_36132,N_37222);
nor U39560 (N_39560,N_36020,N_36749);
xnor U39561 (N_39561,N_37094,N_36377);
or U39562 (N_39562,N_36920,N_37466);
or U39563 (N_39563,N_36449,N_36372);
and U39564 (N_39564,N_36885,N_36214);
xnor U39565 (N_39565,N_37619,N_36358);
xnor U39566 (N_39566,N_36810,N_37363);
or U39567 (N_39567,N_37138,N_36816);
and U39568 (N_39568,N_36258,N_37363);
nor U39569 (N_39569,N_36021,N_36750);
and U39570 (N_39570,N_36960,N_36012);
nor U39571 (N_39571,N_37092,N_36429);
xor U39572 (N_39572,N_37498,N_36359);
xor U39573 (N_39573,N_36941,N_36345);
or U39574 (N_39574,N_36733,N_36728);
nand U39575 (N_39575,N_37017,N_37503);
nor U39576 (N_39576,N_36714,N_37086);
xor U39577 (N_39577,N_36940,N_37279);
or U39578 (N_39578,N_36113,N_37953);
and U39579 (N_39579,N_37959,N_36314);
xor U39580 (N_39580,N_37440,N_36890);
or U39581 (N_39581,N_36524,N_36334);
nor U39582 (N_39582,N_37077,N_36095);
xnor U39583 (N_39583,N_37921,N_37857);
and U39584 (N_39584,N_37756,N_36997);
xnor U39585 (N_39585,N_37434,N_36538);
nand U39586 (N_39586,N_36405,N_36867);
nand U39587 (N_39587,N_37239,N_36273);
and U39588 (N_39588,N_36441,N_37372);
nor U39589 (N_39589,N_37837,N_36165);
nand U39590 (N_39590,N_37901,N_37507);
nor U39591 (N_39591,N_37661,N_37119);
nand U39592 (N_39592,N_37049,N_36731);
or U39593 (N_39593,N_36944,N_36142);
nor U39594 (N_39594,N_36754,N_36124);
or U39595 (N_39595,N_36070,N_37607);
nor U39596 (N_39596,N_36011,N_36859);
and U39597 (N_39597,N_37210,N_37928);
nor U39598 (N_39598,N_36889,N_37763);
nor U39599 (N_39599,N_37156,N_36390);
nand U39600 (N_39600,N_36439,N_36450);
and U39601 (N_39601,N_36205,N_36303);
and U39602 (N_39602,N_36400,N_36814);
or U39603 (N_39603,N_37854,N_36326);
nor U39604 (N_39604,N_36787,N_37809);
and U39605 (N_39605,N_36103,N_37904);
nor U39606 (N_39606,N_37502,N_36559);
xor U39607 (N_39607,N_37228,N_36573);
xnor U39608 (N_39608,N_36244,N_37337);
xor U39609 (N_39609,N_37310,N_37364);
xnor U39610 (N_39610,N_36533,N_36506);
and U39611 (N_39611,N_37892,N_37911);
nor U39612 (N_39612,N_37746,N_36719);
or U39613 (N_39613,N_36640,N_37373);
nand U39614 (N_39614,N_37303,N_36422);
or U39615 (N_39615,N_36037,N_36938);
or U39616 (N_39616,N_36332,N_37229);
and U39617 (N_39617,N_36842,N_37830);
xor U39618 (N_39618,N_37837,N_36519);
and U39619 (N_39619,N_36682,N_37163);
xor U39620 (N_39620,N_36292,N_37985);
and U39621 (N_39621,N_37962,N_36922);
or U39622 (N_39622,N_36552,N_36513);
and U39623 (N_39623,N_37338,N_37821);
xor U39624 (N_39624,N_36774,N_37631);
xnor U39625 (N_39625,N_37777,N_37988);
nand U39626 (N_39626,N_36097,N_36282);
xor U39627 (N_39627,N_36724,N_36954);
xnor U39628 (N_39628,N_36835,N_36271);
and U39629 (N_39629,N_37075,N_37772);
xor U39630 (N_39630,N_37337,N_37775);
xnor U39631 (N_39631,N_37331,N_36888);
and U39632 (N_39632,N_36354,N_37224);
nor U39633 (N_39633,N_37983,N_37674);
nor U39634 (N_39634,N_37095,N_36652);
xor U39635 (N_39635,N_36243,N_36669);
and U39636 (N_39636,N_37689,N_37324);
or U39637 (N_39637,N_36348,N_36975);
xor U39638 (N_39638,N_36647,N_37429);
or U39639 (N_39639,N_36821,N_36896);
and U39640 (N_39640,N_37485,N_36153);
and U39641 (N_39641,N_37484,N_37281);
and U39642 (N_39642,N_37848,N_37853);
nand U39643 (N_39643,N_36610,N_36586);
nor U39644 (N_39644,N_37895,N_36671);
or U39645 (N_39645,N_37974,N_37463);
and U39646 (N_39646,N_36894,N_37054);
xnor U39647 (N_39647,N_36762,N_36834);
xnor U39648 (N_39648,N_37549,N_37364);
xor U39649 (N_39649,N_36073,N_37357);
nor U39650 (N_39650,N_36202,N_36293);
or U39651 (N_39651,N_36730,N_37061);
nor U39652 (N_39652,N_37045,N_36564);
xnor U39653 (N_39653,N_37049,N_37650);
and U39654 (N_39654,N_36342,N_37929);
and U39655 (N_39655,N_37702,N_36397);
or U39656 (N_39656,N_36538,N_36626);
xnor U39657 (N_39657,N_36268,N_36972);
or U39658 (N_39658,N_36526,N_36408);
or U39659 (N_39659,N_37182,N_36320);
xor U39660 (N_39660,N_37282,N_37005);
nor U39661 (N_39661,N_37169,N_36293);
or U39662 (N_39662,N_36398,N_37008);
nor U39663 (N_39663,N_37654,N_36624);
or U39664 (N_39664,N_37458,N_37845);
nor U39665 (N_39665,N_36802,N_36839);
and U39666 (N_39666,N_37595,N_36855);
nor U39667 (N_39667,N_36801,N_37773);
nand U39668 (N_39668,N_36114,N_37104);
and U39669 (N_39669,N_36022,N_36574);
nor U39670 (N_39670,N_37817,N_36647);
nand U39671 (N_39671,N_36463,N_37887);
nor U39672 (N_39672,N_36454,N_36413);
nand U39673 (N_39673,N_36766,N_37883);
nand U39674 (N_39674,N_36067,N_36339);
nand U39675 (N_39675,N_37364,N_37884);
nand U39676 (N_39676,N_37911,N_37806);
nand U39677 (N_39677,N_36237,N_36774);
xor U39678 (N_39678,N_36829,N_36240);
xor U39679 (N_39679,N_36616,N_37735);
nand U39680 (N_39680,N_36038,N_37167);
xor U39681 (N_39681,N_36513,N_37224);
nand U39682 (N_39682,N_37744,N_37677);
or U39683 (N_39683,N_36521,N_36749);
nor U39684 (N_39684,N_36122,N_36653);
nor U39685 (N_39685,N_36495,N_36461);
nor U39686 (N_39686,N_36109,N_37245);
nor U39687 (N_39687,N_36934,N_37076);
nor U39688 (N_39688,N_37185,N_37367);
xor U39689 (N_39689,N_37539,N_37203);
and U39690 (N_39690,N_37898,N_36213);
or U39691 (N_39691,N_37465,N_37885);
nand U39692 (N_39692,N_37324,N_37773);
nor U39693 (N_39693,N_37348,N_36652);
or U39694 (N_39694,N_37083,N_37026);
nand U39695 (N_39695,N_37400,N_36074);
nand U39696 (N_39696,N_36510,N_37578);
nand U39697 (N_39697,N_36644,N_37804);
nor U39698 (N_39698,N_37555,N_37464);
nor U39699 (N_39699,N_36392,N_36287);
and U39700 (N_39700,N_37747,N_37409);
nand U39701 (N_39701,N_36380,N_37067);
nor U39702 (N_39702,N_36549,N_37933);
nor U39703 (N_39703,N_37182,N_36603);
or U39704 (N_39704,N_36747,N_37709);
nor U39705 (N_39705,N_36540,N_37049);
or U39706 (N_39706,N_37628,N_37234);
or U39707 (N_39707,N_36404,N_36648);
xor U39708 (N_39708,N_37274,N_36046);
nand U39709 (N_39709,N_37431,N_37094);
or U39710 (N_39710,N_36771,N_37712);
xor U39711 (N_39711,N_37997,N_36445);
and U39712 (N_39712,N_36891,N_37960);
or U39713 (N_39713,N_36104,N_37764);
and U39714 (N_39714,N_37654,N_36765);
nor U39715 (N_39715,N_36700,N_37702);
nor U39716 (N_39716,N_36651,N_36181);
nand U39717 (N_39717,N_36385,N_36207);
or U39718 (N_39718,N_37442,N_37184);
nand U39719 (N_39719,N_36180,N_36963);
xnor U39720 (N_39720,N_37471,N_36128);
nor U39721 (N_39721,N_36474,N_37404);
xor U39722 (N_39722,N_37641,N_36962);
nor U39723 (N_39723,N_36783,N_36367);
nor U39724 (N_39724,N_37413,N_36786);
and U39725 (N_39725,N_37606,N_37417);
nor U39726 (N_39726,N_36208,N_37608);
and U39727 (N_39727,N_36866,N_36649);
and U39728 (N_39728,N_36029,N_36398);
or U39729 (N_39729,N_37989,N_36670);
xnor U39730 (N_39730,N_37821,N_37835);
nand U39731 (N_39731,N_37769,N_37200);
or U39732 (N_39732,N_37500,N_36311);
and U39733 (N_39733,N_37887,N_36195);
xor U39734 (N_39734,N_37514,N_36597);
or U39735 (N_39735,N_37607,N_37331);
and U39736 (N_39736,N_37959,N_36900);
nor U39737 (N_39737,N_37538,N_37894);
xor U39738 (N_39738,N_37082,N_37307);
nand U39739 (N_39739,N_36598,N_36947);
nand U39740 (N_39740,N_36326,N_36174);
xor U39741 (N_39741,N_37056,N_37791);
or U39742 (N_39742,N_37214,N_36332);
nand U39743 (N_39743,N_36163,N_36996);
nand U39744 (N_39744,N_37067,N_37178);
nand U39745 (N_39745,N_36305,N_36643);
xor U39746 (N_39746,N_37453,N_36629);
and U39747 (N_39747,N_37233,N_37893);
or U39748 (N_39748,N_36019,N_36772);
or U39749 (N_39749,N_36245,N_37451);
nor U39750 (N_39750,N_36952,N_36546);
nand U39751 (N_39751,N_36741,N_36270);
xor U39752 (N_39752,N_36192,N_36609);
or U39753 (N_39753,N_36002,N_37066);
xor U39754 (N_39754,N_36747,N_36407);
and U39755 (N_39755,N_37023,N_37891);
and U39756 (N_39756,N_37151,N_36946);
or U39757 (N_39757,N_37654,N_37595);
xor U39758 (N_39758,N_37829,N_36818);
nor U39759 (N_39759,N_36795,N_36068);
and U39760 (N_39760,N_36346,N_37189);
nand U39761 (N_39761,N_37883,N_36829);
or U39762 (N_39762,N_36889,N_37446);
nor U39763 (N_39763,N_36951,N_36054);
or U39764 (N_39764,N_36383,N_36865);
and U39765 (N_39765,N_37634,N_37423);
nand U39766 (N_39766,N_36552,N_36200);
xor U39767 (N_39767,N_37987,N_36907);
nor U39768 (N_39768,N_36317,N_36725);
and U39769 (N_39769,N_36832,N_36786);
and U39770 (N_39770,N_36155,N_37892);
and U39771 (N_39771,N_36027,N_37011);
nand U39772 (N_39772,N_36346,N_36296);
xor U39773 (N_39773,N_36818,N_36469);
nand U39774 (N_39774,N_37094,N_36364);
and U39775 (N_39775,N_36821,N_36978);
and U39776 (N_39776,N_36622,N_37959);
or U39777 (N_39777,N_36063,N_37244);
or U39778 (N_39778,N_36119,N_37340);
or U39779 (N_39779,N_37178,N_37245);
or U39780 (N_39780,N_37778,N_37757);
xor U39781 (N_39781,N_37523,N_36694);
or U39782 (N_39782,N_37077,N_37466);
and U39783 (N_39783,N_36742,N_36519);
nor U39784 (N_39784,N_37862,N_36360);
nor U39785 (N_39785,N_36107,N_37224);
nand U39786 (N_39786,N_36969,N_36666);
nand U39787 (N_39787,N_36785,N_36082);
nor U39788 (N_39788,N_36936,N_37622);
nor U39789 (N_39789,N_36403,N_36419);
nor U39790 (N_39790,N_37853,N_37525);
or U39791 (N_39791,N_37559,N_37146);
and U39792 (N_39792,N_37181,N_37238);
or U39793 (N_39793,N_37928,N_37477);
xor U39794 (N_39794,N_36531,N_36812);
and U39795 (N_39795,N_36337,N_37469);
nand U39796 (N_39796,N_37109,N_37235);
and U39797 (N_39797,N_36772,N_37085);
and U39798 (N_39798,N_37455,N_37659);
nor U39799 (N_39799,N_37874,N_36039);
xnor U39800 (N_39800,N_36489,N_37651);
nand U39801 (N_39801,N_37544,N_37278);
and U39802 (N_39802,N_37302,N_36836);
nand U39803 (N_39803,N_36987,N_36737);
and U39804 (N_39804,N_37211,N_37288);
or U39805 (N_39805,N_36254,N_36520);
or U39806 (N_39806,N_36713,N_36703);
xor U39807 (N_39807,N_36843,N_36950);
and U39808 (N_39808,N_36571,N_37708);
nand U39809 (N_39809,N_37421,N_36827);
nand U39810 (N_39810,N_36692,N_36756);
or U39811 (N_39811,N_36991,N_36103);
xnor U39812 (N_39812,N_37729,N_36824);
or U39813 (N_39813,N_36317,N_36332);
nand U39814 (N_39814,N_37010,N_36996);
nand U39815 (N_39815,N_37642,N_37878);
nor U39816 (N_39816,N_36213,N_37658);
and U39817 (N_39817,N_37592,N_37314);
or U39818 (N_39818,N_37060,N_37822);
nor U39819 (N_39819,N_36911,N_36355);
and U39820 (N_39820,N_36773,N_37132);
xor U39821 (N_39821,N_37332,N_37613);
nand U39822 (N_39822,N_37036,N_36964);
or U39823 (N_39823,N_37283,N_36373);
nor U39824 (N_39824,N_37511,N_36129);
and U39825 (N_39825,N_36358,N_36794);
and U39826 (N_39826,N_37014,N_37359);
nor U39827 (N_39827,N_36706,N_36326);
xnor U39828 (N_39828,N_37756,N_37717);
or U39829 (N_39829,N_36877,N_37417);
nand U39830 (N_39830,N_36544,N_36342);
and U39831 (N_39831,N_37061,N_37244);
and U39832 (N_39832,N_37228,N_36441);
xor U39833 (N_39833,N_37497,N_37731);
nor U39834 (N_39834,N_37177,N_36927);
and U39835 (N_39835,N_37486,N_37719);
and U39836 (N_39836,N_37686,N_37040);
nor U39837 (N_39837,N_37138,N_37505);
or U39838 (N_39838,N_37712,N_37482);
nor U39839 (N_39839,N_36302,N_36388);
nor U39840 (N_39840,N_36778,N_37496);
or U39841 (N_39841,N_36040,N_37848);
and U39842 (N_39842,N_36275,N_37665);
and U39843 (N_39843,N_36060,N_36687);
nand U39844 (N_39844,N_36784,N_37692);
xor U39845 (N_39845,N_37412,N_36292);
xnor U39846 (N_39846,N_36414,N_36687);
and U39847 (N_39847,N_37500,N_37269);
nor U39848 (N_39848,N_37838,N_37550);
and U39849 (N_39849,N_36321,N_37275);
nand U39850 (N_39850,N_37572,N_36306);
nor U39851 (N_39851,N_37680,N_36217);
or U39852 (N_39852,N_36369,N_37632);
or U39853 (N_39853,N_37117,N_36434);
and U39854 (N_39854,N_36467,N_36395);
xnor U39855 (N_39855,N_37055,N_36369);
nor U39856 (N_39856,N_37638,N_37902);
or U39857 (N_39857,N_36514,N_36602);
nand U39858 (N_39858,N_36119,N_37932);
nor U39859 (N_39859,N_37355,N_36265);
nor U39860 (N_39860,N_37786,N_37976);
nand U39861 (N_39861,N_37613,N_36337);
nand U39862 (N_39862,N_37399,N_37777);
or U39863 (N_39863,N_36825,N_37564);
or U39864 (N_39864,N_37838,N_36693);
or U39865 (N_39865,N_37308,N_36515);
xor U39866 (N_39866,N_36795,N_36297);
xnor U39867 (N_39867,N_36485,N_36549);
nor U39868 (N_39868,N_36594,N_36900);
or U39869 (N_39869,N_36604,N_37634);
and U39870 (N_39870,N_37575,N_37050);
or U39871 (N_39871,N_36981,N_36742);
xnor U39872 (N_39872,N_37887,N_37692);
nand U39873 (N_39873,N_36854,N_37547);
and U39874 (N_39874,N_37500,N_37955);
xor U39875 (N_39875,N_37084,N_36023);
and U39876 (N_39876,N_36406,N_36984);
and U39877 (N_39877,N_37864,N_36005);
nand U39878 (N_39878,N_37163,N_37986);
and U39879 (N_39879,N_36409,N_37934);
nand U39880 (N_39880,N_37980,N_36218);
and U39881 (N_39881,N_36625,N_37219);
or U39882 (N_39882,N_36360,N_37259);
nand U39883 (N_39883,N_36673,N_36768);
or U39884 (N_39884,N_36718,N_37197);
nand U39885 (N_39885,N_37936,N_37489);
nor U39886 (N_39886,N_36027,N_36516);
or U39887 (N_39887,N_37728,N_37740);
nor U39888 (N_39888,N_37130,N_36951);
or U39889 (N_39889,N_36776,N_37255);
nor U39890 (N_39890,N_36604,N_36079);
nand U39891 (N_39891,N_37805,N_36701);
xor U39892 (N_39892,N_36534,N_36967);
xor U39893 (N_39893,N_37370,N_36496);
xnor U39894 (N_39894,N_36478,N_36485);
or U39895 (N_39895,N_37037,N_36471);
nor U39896 (N_39896,N_36982,N_36219);
xor U39897 (N_39897,N_36454,N_37896);
nor U39898 (N_39898,N_37527,N_37377);
nor U39899 (N_39899,N_36929,N_36891);
nor U39900 (N_39900,N_36013,N_36126);
nor U39901 (N_39901,N_36251,N_37701);
and U39902 (N_39902,N_36715,N_36697);
and U39903 (N_39903,N_36896,N_36842);
and U39904 (N_39904,N_36429,N_36664);
or U39905 (N_39905,N_36109,N_37040);
nand U39906 (N_39906,N_36778,N_37269);
or U39907 (N_39907,N_37757,N_37500);
and U39908 (N_39908,N_36063,N_36819);
nand U39909 (N_39909,N_36486,N_36227);
xnor U39910 (N_39910,N_37216,N_37343);
and U39911 (N_39911,N_36668,N_37119);
xnor U39912 (N_39912,N_36226,N_36886);
nor U39913 (N_39913,N_37701,N_37809);
nand U39914 (N_39914,N_37751,N_37401);
nor U39915 (N_39915,N_37857,N_37001);
nand U39916 (N_39916,N_36561,N_37560);
nand U39917 (N_39917,N_37299,N_36511);
and U39918 (N_39918,N_37222,N_36325);
nand U39919 (N_39919,N_36158,N_36715);
nor U39920 (N_39920,N_36197,N_37028);
xor U39921 (N_39921,N_37893,N_37333);
and U39922 (N_39922,N_37119,N_36503);
nor U39923 (N_39923,N_37684,N_36099);
nand U39924 (N_39924,N_37527,N_37602);
or U39925 (N_39925,N_36607,N_36650);
xor U39926 (N_39926,N_37321,N_36190);
and U39927 (N_39927,N_36589,N_37381);
and U39928 (N_39928,N_36131,N_37411);
nor U39929 (N_39929,N_36877,N_36323);
nand U39930 (N_39930,N_36852,N_36739);
xor U39931 (N_39931,N_36982,N_37564);
and U39932 (N_39932,N_36670,N_36770);
nand U39933 (N_39933,N_37686,N_37278);
or U39934 (N_39934,N_37417,N_36915);
or U39935 (N_39935,N_36545,N_37244);
nor U39936 (N_39936,N_36172,N_37533);
and U39937 (N_39937,N_36875,N_36618);
or U39938 (N_39938,N_37602,N_37181);
or U39939 (N_39939,N_36683,N_37293);
nor U39940 (N_39940,N_37042,N_36816);
nand U39941 (N_39941,N_37537,N_36608);
nor U39942 (N_39942,N_37992,N_36945);
or U39943 (N_39943,N_37563,N_37854);
or U39944 (N_39944,N_36821,N_36812);
nand U39945 (N_39945,N_37304,N_36645);
or U39946 (N_39946,N_37780,N_36843);
nand U39947 (N_39947,N_37824,N_37735);
nand U39948 (N_39948,N_37484,N_36945);
xor U39949 (N_39949,N_36685,N_36655);
or U39950 (N_39950,N_36124,N_36283);
and U39951 (N_39951,N_37294,N_36034);
and U39952 (N_39952,N_36129,N_36158);
nand U39953 (N_39953,N_37245,N_37765);
and U39954 (N_39954,N_36619,N_36414);
or U39955 (N_39955,N_36171,N_37155);
nand U39956 (N_39956,N_37357,N_36627);
nor U39957 (N_39957,N_37190,N_37462);
and U39958 (N_39958,N_36209,N_37481);
nand U39959 (N_39959,N_37538,N_37576);
nor U39960 (N_39960,N_36905,N_37648);
nand U39961 (N_39961,N_36594,N_37025);
nor U39962 (N_39962,N_37385,N_36131);
and U39963 (N_39963,N_37709,N_37146);
xnor U39964 (N_39964,N_36121,N_37780);
xor U39965 (N_39965,N_36613,N_37162);
and U39966 (N_39966,N_36324,N_36628);
and U39967 (N_39967,N_37304,N_37163);
and U39968 (N_39968,N_36585,N_36276);
nand U39969 (N_39969,N_36680,N_37674);
nand U39970 (N_39970,N_37864,N_36964);
xor U39971 (N_39971,N_37654,N_37529);
or U39972 (N_39972,N_37955,N_36854);
and U39973 (N_39973,N_36847,N_36680);
or U39974 (N_39974,N_37078,N_37821);
nor U39975 (N_39975,N_37038,N_36789);
xor U39976 (N_39976,N_36555,N_36986);
nand U39977 (N_39977,N_36795,N_36532);
or U39978 (N_39978,N_37730,N_36180);
and U39979 (N_39979,N_36173,N_37850);
or U39980 (N_39980,N_36162,N_36670);
xnor U39981 (N_39981,N_37664,N_36350);
nand U39982 (N_39982,N_37410,N_37395);
nand U39983 (N_39983,N_36488,N_36153);
or U39984 (N_39984,N_36991,N_37359);
xnor U39985 (N_39985,N_36876,N_36906);
nand U39986 (N_39986,N_36203,N_36814);
nor U39987 (N_39987,N_36035,N_36554);
nand U39988 (N_39988,N_37724,N_37506);
xnor U39989 (N_39989,N_37908,N_37454);
or U39990 (N_39990,N_36389,N_37640);
nor U39991 (N_39991,N_37693,N_36092);
and U39992 (N_39992,N_36047,N_36370);
or U39993 (N_39993,N_36857,N_36074);
or U39994 (N_39994,N_36332,N_37401);
or U39995 (N_39995,N_36996,N_36475);
nor U39996 (N_39996,N_37114,N_37581);
nor U39997 (N_39997,N_37573,N_37245);
nor U39998 (N_39998,N_36960,N_36302);
and U39999 (N_39999,N_36146,N_37498);
and U40000 (N_40000,N_39176,N_38083);
nor U40001 (N_40001,N_39153,N_39717);
nor U40002 (N_40002,N_39072,N_38265);
and U40003 (N_40003,N_39621,N_39952);
xor U40004 (N_40004,N_38211,N_39350);
or U40005 (N_40005,N_38797,N_38806);
nor U40006 (N_40006,N_38516,N_38964);
nand U40007 (N_40007,N_38236,N_38412);
and U40008 (N_40008,N_38608,N_38930);
and U40009 (N_40009,N_38268,N_39385);
nor U40010 (N_40010,N_38543,N_39925);
nand U40011 (N_40011,N_39310,N_39093);
and U40012 (N_40012,N_39727,N_39288);
nand U40013 (N_40013,N_38775,N_38400);
and U40014 (N_40014,N_39500,N_39149);
and U40015 (N_40015,N_38899,N_39331);
nand U40016 (N_40016,N_39316,N_38135);
or U40017 (N_40017,N_39516,N_38942);
or U40018 (N_40018,N_38283,N_38985);
and U40019 (N_40019,N_38905,N_39212);
nor U40020 (N_40020,N_38491,N_38151);
and U40021 (N_40021,N_39896,N_39029);
and U40022 (N_40022,N_39195,N_38718);
xnor U40023 (N_40023,N_38218,N_38909);
xor U40024 (N_40024,N_38673,N_38632);
nor U40025 (N_40025,N_39325,N_38851);
nand U40026 (N_40026,N_38091,N_38109);
or U40027 (N_40027,N_38809,N_39617);
or U40028 (N_40028,N_39349,N_39730);
nand U40029 (N_40029,N_38731,N_39731);
and U40030 (N_40030,N_38856,N_39902);
xnor U40031 (N_40031,N_39642,N_38871);
or U40032 (N_40032,N_38936,N_38393);
and U40033 (N_40033,N_38790,N_38857);
and U40034 (N_40034,N_38814,N_39892);
xnor U40035 (N_40035,N_39619,N_39081);
nor U40036 (N_40036,N_39131,N_38363);
or U40037 (N_40037,N_39336,N_38604);
and U40038 (N_40038,N_39311,N_38453);
nand U40039 (N_40039,N_38888,N_39495);
nor U40040 (N_40040,N_38063,N_39564);
and U40041 (N_40041,N_38503,N_38147);
xor U40042 (N_40042,N_39358,N_38891);
xor U40043 (N_40043,N_38597,N_38407);
nor U40044 (N_40044,N_39102,N_39686);
and U40045 (N_40045,N_39339,N_38685);
and U40046 (N_40046,N_39109,N_38892);
or U40047 (N_40047,N_39620,N_38782);
nand U40048 (N_40048,N_38486,N_38337);
and U40049 (N_40049,N_39048,N_38781);
nor U40050 (N_40050,N_38348,N_39887);
nand U40051 (N_40051,N_39772,N_38327);
nor U40052 (N_40052,N_39735,N_39696);
or U40053 (N_40053,N_38522,N_39571);
and U40054 (N_40054,N_39026,N_39613);
and U40055 (N_40055,N_38767,N_39874);
nor U40056 (N_40056,N_39913,N_39127);
nand U40057 (N_40057,N_39742,N_38499);
nand U40058 (N_40058,N_39200,N_39476);
xor U40059 (N_40059,N_38049,N_38196);
nor U40060 (N_40060,N_38875,N_38678);
or U40061 (N_40061,N_38575,N_39684);
or U40062 (N_40062,N_38528,N_38020);
or U40063 (N_40063,N_38434,N_38170);
xnor U40064 (N_40064,N_39830,N_39858);
or U40065 (N_40065,N_38935,N_38601);
nand U40066 (N_40066,N_39294,N_38569);
or U40067 (N_40067,N_38445,N_39474);
nand U40068 (N_40068,N_39003,N_39544);
nand U40069 (N_40069,N_38086,N_38341);
or U40070 (N_40070,N_39572,N_39144);
xnor U40071 (N_40071,N_39369,N_39503);
and U40072 (N_40072,N_39025,N_38640);
xnor U40073 (N_40073,N_39086,N_39443);
nor U40074 (N_40074,N_38457,N_38563);
and U40075 (N_40075,N_38869,N_38527);
or U40076 (N_40076,N_39893,N_39122);
nor U40077 (N_40077,N_39205,N_39707);
xor U40078 (N_40078,N_39427,N_39412);
or U40079 (N_40079,N_38843,N_39929);
nor U40080 (N_40080,N_39984,N_38367);
and U40081 (N_40081,N_38037,N_39537);
nor U40082 (N_40082,N_38354,N_39335);
nand U40083 (N_40083,N_38150,N_38773);
nor U40084 (N_40084,N_38810,N_39805);
and U40085 (N_40085,N_38255,N_38550);
and U40086 (N_40086,N_39843,N_39279);
nand U40087 (N_40087,N_38183,N_38258);
xor U40088 (N_40088,N_38276,N_39302);
xnor U40089 (N_40089,N_39654,N_39021);
or U40090 (N_40090,N_38284,N_39956);
nand U40091 (N_40091,N_39275,N_38431);
xnor U40092 (N_40092,N_39317,N_39511);
and U40093 (N_40093,N_39290,N_39567);
and U40094 (N_40094,N_38047,N_39228);
nor U40095 (N_40095,N_39258,N_38429);
nor U40096 (N_40096,N_39065,N_38315);
nor U40097 (N_40097,N_38920,N_38073);
nor U40098 (N_40098,N_39607,N_39608);
xor U40099 (N_40099,N_39099,N_39560);
and U40100 (N_40100,N_39752,N_39273);
xor U40101 (N_40101,N_39857,N_38243);
nor U40102 (N_40102,N_39491,N_38906);
xor U40103 (N_40103,N_38842,N_39870);
nand U40104 (N_40104,N_39804,N_39246);
nand U40105 (N_40105,N_38730,N_38154);
and U40106 (N_40106,N_38970,N_39594);
nand U40107 (N_40107,N_39761,N_39950);
xor U40108 (N_40108,N_38532,N_39970);
and U40109 (N_40109,N_39169,N_39538);
nand U40110 (N_40110,N_38002,N_39070);
nor U40111 (N_40111,N_38743,N_39994);
nor U40112 (N_40112,N_38387,N_38981);
or U40113 (N_40113,N_38143,N_39862);
nand U40114 (N_40114,N_39019,N_39531);
or U40115 (N_40115,N_39418,N_38697);
nand U40116 (N_40116,N_38441,N_39423);
nand U40117 (N_40117,N_39390,N_39561);
nand U40118 (N_40118,N_39298,N_38646);
nand U40119 (N_40119,N_38165,N_39927);
nand U40120 (N_40120,N_38749,N_39126);
xnor U40121 (N_40121,N_39392,N_39507);
and U40122 (N_40122,N_39043,N_38370);
nand U40123 (N_40123,N_38616,N_39055);
or U40124 (N_40124,N_38353,N_39827);
nand U40125 (N_40125,N_39340,N_38314);
or U40126 (N_40126,N_38475,N_39911);
or U40127 (N_40127,N_38826,N_38325);
or U40128 (N_40128,N_38253,N_39801);
nor U40129 (N_40129,N_39393,N_38539);
nor U40130 (N_40130,N_38022,N_39701);
or U40131 (N_40131,N_38798,N_39875);
nor U40132 (N_40132,N_38128,N_39067);
and U40133 (N_40133,N_39628,N_39915);
and U40134 (N_40134,N_39869,N_38096);
xnor U40135 (N_40135,N_39433,N_38986);
xnor U40136 (N_40136,N_39087,N_38162);
xnor U40137 (N_40137,N_39809,N_38644);
nand U40138 (N_40138,N_38684,N_39330);
and U40139 (N_40139,N_38228,N_38657);
xor U40140 (N_40140,N_38947,N_39213);
nor U40141 (N_40141,N_39464,N_38090);
or U40142 (N_40142,N_39227,N_39168);
or U40143 (N_40143,N_38694,N_39630);
and U40144 (N_40144,N_39973,N_39615);
nand U40145 (N_40145,N_39196,N_39557);
and U40146 (N_40146,N_38229,N_38862);
and U40147 (N_40147,N_38870,N_38378);
and U40148 (N_40148,N_38804,N_39563);
nand U40149 (N_40149,N_39876,N_38141);
xor U40150 (N_40150,N_38541,N_38591);
nor U40151 (N_40151,N_38028,N_39400);
nand U40152 (N_40152,N_38304,N_39850);
nor U40153 (N_40153,N_38799,N_39525);
xor U40154 (N_40154,N_39224,N_38662);
nor U40155 (N_40155,N_38536,N_39420);
or U40156 (N_40156,N_38368,N_38753);
and U40157 (N_40157,N_38984,N_39979);
nand U40158 (N_40158,N_39705,N_39983);
or U40159 (N_40159,N_38661,N_39849);
nand U40160 (N_40160,N_39441,N_39825);
nor U40161 (N_40161,N_39199,N_38706);
nor U40162 (N_40162,N_39481,N_38023);
nor U40163 (N_40163,N_39091,N_38670);
and U40164 (N_40164,N_39475,N_38254);
nor U40165 (N_40165,N_39105,N_38783);
xor U40166 (N_40166,N_39562,N_39004);
or U40167 (N_40167,N_38776,N_39776);
nor U40168 (N_40168,N_39382,N_39765);
nand U40169 (N_40169,N_38588,N_39023);
or U40170 (N_40170,N_39535,N_39609);
nand U40171 (N_40171,N_38745,N_38562);
xnor U40172 (N_40172,N_39906,N_38709);
and U40173 (N_40173,N_38958,N_39863);
xor U40174 (N_40174,N_38950,N_38358);
nand U40175 (N_40175,N_39177,N_39885);
nand U40176 (N_40176,N_38902,N_39883);
nand U40177 (N_40177,N_39838,N_38117);
or U40178 (N_40178,N_39920,N_39380);
and U40179 (N_40179,N_39257,N_38722);
nand U40180 (N_40180,N_38852,N_38940);
nand U40181 (N_40181,N_39991,N_38894);
nand U40182 (N_40182,N_38224,N_38778);
xor U40183 (N_40183,N_39136,N_39729);
or U40184 (N_40184,N_39499,N_39512);
nor U40185 (N_40185,N_38373,N_39243);
nand U40186 (N_40186,N_39990,N_39467);
nand U40187 (N_40187,N_38605,N_39156);
and U40188 (N_40188,N_38800,N_39817);
nor U40189 (N_40189,N_38040,N_38113);
or U40190 (N_40190,N_39494,N_39775);
xnor U40191 (N_40191,N_39834,N_39178);
or U40192 (N_40192,N_38351,N_39027);
xor U40193 (N_40193,N_38329,N_38688);
nor U40194 (N_40194,N_39379,N_39450);
and U40195 (N_40195,N_39219,N_38227);
or U40196 (N_40196,N_39389,N_38655);
or U40197 (N_40197,N_39673,N_39753);
or U40198 (N_40198,N_38295,N_38967);
and U40199 (N_40199,N_39051,N_38298);
and U40200 (N_40200,N_38712,N_39364);
or U40201 (N_40201,N_39030,N_39388);
or U40202 (N_40202,N_39370,N_38222);
xnor U40203 (N_40203,N_39147,N_39683);
nor U40204 (N_40204,N_38250,N_38787);
nand U40205 (N_40205,N_38683,N_39362);
and U40206 (N_40206,N_38951,N_39092);
nand U40207 (N_40207,N_38647,N_39437);
nor U40208 (N_40208,N_38450,N_39103);
and U40209 (N_40209,N_39704,N_39645);
or U40210 (N_40210,N_38285,N_39581);
and U40211 (N_40211,N_38133,N_39044);
nor U40212 (N_40212,N_38038,N_39189);
xnor U40213 (N_40213,N_38883,N_39163);
xor U40214 (N_40214,N_39540,N_39632);
or U40215 (N_40215,N_39300,N_39376);
xnor U40216 (N_40216,N_38840,N_38786);
nand U40217 (N_40217,N_38677,N_38500);
nand U40218 (N_40218,N_38651,N_38312);
and U40219 (N_40219,N_38244,N_38910);
and U40220 (N_40220,N_39890,N_38669);
xor U40221 (N_40221,N_39234,N_39745);
or U40222 (N_40222,N_38596,N_39315);
xnor U40223 (N_40223,N_38956,N_39725);
or U40224 (N_40224,N_39924,N_38231);
xor U40225 (N_40225,N_39101,N_38580);
nand U40226 (N_40226,N_39658,N_38829);
xnor U40227 (N_40227,N_38844,N_38997);
nor U40228 (N_40228,N_39904,N_39134);
or U40229 (N_40229,N_39647,N_39605);
and U40230 (N_40230,N_38469,N_39050);
or U40231 (N_40231,N_38217,N_39554);
or U40232 (N_40232,N_39971,N_38146);
xor U40233 (N_40233,N_38079,N_39650);
nand U40234 (N_40234,N_38357,N_39969);
or U40235 (N_40235,N_38025,N_38733);
or U40236 (N_40236,N_39305,N_39665);
nand U40237 (N_40237,N_39945,N_39789);
xnor U40238 (N_40238,N_38957,N_39785);
nand U40239 (N_40239,N_38705,N_38919);
or U40240 (N_40240,N_39712,N_39342);
or U40241 (N_40241,N_38080,N_38366);
and U40242 (N_40242,N_39792,N_39465);
and U40243 (N_40243,N_39098,N_39239);
nand U40244 (N_40244,N_39853,N_38582);
xnor U40245 (N_40245,N_39711,N_38839);
xnor U40246 (N_40246,N_38896,N_39552);
nand U40247 (N_40247,N_38832,N_39457);
nor U40248 (N_40248,N_39011,N_39680);
nor U40249 (N_40249,N_39308,N_38521);
xor U40250 (N_40250,N_38638,N_39341);
xnor U40251 (N_40251,N_39541,N_38269);
and U40252 (N_40252,N_39409,N_39659);
and U40253 (N_40253,N_38451,N_39872);
nand U40254 (N_40254,N_38242,N_38506);
and U40255 (N_40255,N_39010,N_39723);
or U40256 (N_40256,N_38009,N_39784);
or U40257 (N_40257,N_38430,N_38511);
nor U40258 (N_40258,N_39528,N_38111);
nor U40259 (N_40259,N_38791,N_39151);
nor U40260 (N_40260,N_38264,N_38708);
xor U40261 (N_40261,N_38728,N_39414);
or U40262 (N_40262,N_39555,N_39269);
nor U40263 (N_40263,N_38310,N_38579);
and U40264 (N_40264,N_38794,N_39881);
nand U40265 (N_40265,N_38741,N_39656);
nand U40266 (N_40266,N_39842,N_39117);
xnor U40267 (N_40267,N_39822,N_39488);
nand U40268 (N_40268,N_38496,N_39319);
xor U40269 (N_40269,N_39271,N_38637);
nand U40270 (N_40270,N_38130,N_38779);
and U40271 (N_40271,N_38623,N_39988);
and U40272 (N_40272,N_38505,N_38937);
nand U40273 (N_40273,N_39054,N_38927);
nor U40274 (N_40274,N_38051,N_38618);
and U40275 (N_40275,N_38477,N_39530);
and U40276 (N_40276,N_38234,N_39301);
or U40277 (N_40277,N_39919,N_38710);
nand U40278 (N_40278,N_39773,N_39754);
or U40279 (N_40279,N_38725,N_39936);
nor U40280 (N_40280,N_39415,N_38012);
or U40281 (N_40281,N_39997,N_39068);
or U40282 (N_40282,N_38538,N_38995);
and U40283 (N_40283,N_39867,N_39695);
nand U40284 (N_40284,N_38874,N_38483);
nand U40285 (N_40285,N_39550,N_39798);
and U40286 (N_40286,N_39677,N_39962);
and U40287 (N_40287,N_39959,N_38901);
and U40288 (N_40288,N_38139,N_38629);
xnor U40289 (N_40289,N_38816,N_39624);
and U40290 (N_40290,N_38006,N_39599);
xnor U40291 (N_40291,N_38793,N_38723);
nor U40292 (N_40292,N_39847,N_39836);
nand U40293 (N_40293,N_39931,N_39185);
and U40294 (N_40294,N_38311,N_39618);
nand U40295 (N_40295,N_39631,N_38692);
xnor U40296 (N_40296,N_38121,N_39737);
xor U40297 (N_40297,N_38026,N_38593);
xnor U40298 (N_40298,N_38200,N_38365);
nor U40299 (N_40299,N_39174,N_39006);
xnor U40300 (N_40300,N_38897,N_38059);
and U40301 (N_40301,N_39209,N_39247);
xor U40302 (N_40302,N_38460,N_38561);
or U40303 (N_40303,N_39606,N_38176);
and U40304 (N_40304,N_39261,N_38360);
or U40305 (N_40305,N_38858,N_38645);
and U40306 (N_40306,N_38201,N_38900);
nand U40307 (N_40307,N_39118,N_38567);
and U40308 (N_40308,N_39734,N_39974);
nor U40309 (N_40309,N_38966,N_39018);
xnor U40310 (N_40310,N_38755,N_39164);
or U40311 (N_40311,N_39405,N_39688);
nand U40312 (N_40312,N_38145,N_38933);
nor U40313 (N_40313,N_38520,N_39732);
or U40314 (N_40314,N_38017,N_39855);
and U40315 (N_40315,N_39460,N_38458);
xor U40316 (N_40316,N_39816,N_38112);
xor U40317 (N_40317,N_39953,N_39452);
nor U40318 (N_40318,N_38713,N_39715);
or U40319 (N_40319,N_39254,N_38886);
or U40320 (N_40320,N_39496,N_38598);
or U40321 (N_40321,N_38214,N_39877);
nor U40322 (N_40322,N_39413,N_38526);
nor U40323 (N_40323,N_39739,N_39192);
and U40324 (N_40324,N_39839,N_38204);
xnor U40325 (N_40325,N_39778,N_38385);
and U40326 (N_40326,N_38383,N_39113);
and U40327 (N_40327,N_38621,N_39949);
nor U40328 (N_40328,N_38485,N_38418);
nor U40329 (N_40329,N_38476,N_38402);
and U40330 (N_40330,N_38884,N_38277);
nand U40331 (N_40331,N_39461,N_39106);
xnor U40332 (N_40332,N_39095,N_39646);
xor U40333 (N_40333,N_39946,N_38292);
nor U40334 (N_40334,N_38737,N_39791);
nand U40335 (N_40335,N_39878,N_39932);
xnor U40336 (N_40336,N_39756,N_38168);
nand U40337 (N_40337,N_39262,N_38473);
nor U40338 (N_40338,N_38568,N_39795);
xor U40339 (N_40339,N_39399,N_39546);
and U40340 (N_40340,N_39755,N_38992);
xor U40341 (N_40341,N_38414,N_39374);
nor U40342 (N_40342,N_38554,N_39277);
and U40343 (N_40343,N_39080,N_39985);
and U40344 (N_40344,N_39241,N_38974);
nor U40345 (N_40345,N_38849,N_39972);
or U40346 (N_40346,N_38946,N_38488);
nor U40347 (N_40347,N_38278,N_39000);
xor U40348 (N_40348,N_39611,N_39485);
and U40349 (N_40349,N_39318,N_38388);
xnor U40350 (N_40350,N_39322,N_38043);
nand U40351 (N_40351,N_39668,N_39282);
nand U40352 (N_40352,N_39748,N_38297);
and U40353 (N_40353,N_39509,N_39671);
nand U40354 (N_40354,N_38847,N_39865);
or U40355 (N_40355,N_39996,N_39142);
nand U40356 (N_40356,N_39639,N_39966);
or U40357 (N_40357,N_39057,N_38939);
and U40358 (N_40358,N_39909,N_39718);
nand U40359 (N_40359,N_38690,N_38889);
or U40360 (N_40360,N_38260,N_39375);
nand U40361 (N_40361,N_38399,N_38693);
nor U40362 (N_40362,N_39998,N_38462);
and U40363 (N_40363,N_38738,N_39439);
nor U40364 (N_40364,N_39139,N_39137);
xnor U40365 (N_40365,N_38194,N_38479);
nor U40366 (N_40366,N_39764,N_39455);
and U40367 (N_40367,N_38758,N_39907);
nor U40368 (N_40368,N_39272,N_39861);
xnor U40369 (N_40369,N_39542,N_39899);
nand U40370 (N_40370,N_39833,N_38795);
nor U40371 (N_40371,N_38225,N_38286);
or U40372 (N_40372,N_38846,N_39150);
and U40373 (N_40373,N_38424,N_39558);
xnor U40374 (N_40374,N_39252,N_39202);
xnor U40375 (N_40375,N_39210,N_39506);
or U40376 (N_40376,N_38926,N_38355);
xor U40377 (N_40377,N_38053,N_38911);
or U40378 (N_40378,N_39333,N_39832);
and U40379 (N_40379,N_38665,N_39135);
and U40380 (N_40380,N_39186,N_39267);
nor U40381 (N_40381,N_38160,N_39750);
nor U40382 (N_40382,N_39284,N_39759);
and U40383 (N_40383,N_38811,N_38792);
nor U40384 (N_40384,N_38863,N_39944);
nor U40385 (N_40385,N_38099,N_39416);
nand U40386 (N_40386,N_38386,N_39041);
and U40387 (N_40387,N_39037,N_38817);
and U40388 (N_40388,N_39851,N_38291);
or U40389 (N_40389,N_39394,N_38282);
xnor U40390 (N_40390,N_39536,N_39141);
nand U40391 (N_40391,N_39038,N_39864);
nor U40392 (N_40392,N_39720,N_39638);
and U40393 (N_40393,N_39407,N_38834);
or U40394 (N_40394,N_39600,N_38700);
nand U40395 (N_40395,N_38841,N_38195);
xnor U40396 (N_40396,N_39976,N_38784);
nor U40397 (N_40397,N_38108,N_39928);
nor U40398 (N_40398,N_39280,N_39593);
nor U40399 (N_40399,N_39088,N_38308);
xnor U40400 (N_40400,N_39360,N_38021);
nand U40401 (N_40401,N_38078,N_39125);
xor U40402 (N_40402,N_38409,N_39447);
and U40403 (N_40403,N_39303,N_38603);
and U40404 (N_40404,N_39373,N_38129);
and U40405 (N_40405,N_38633,N_39253);
xnor U40406 (N_40406,N_38490,N_38118);
nor U40407 (N_40407,N_39844,N_38232);
or U40408 (N_40408,N_39498,N_39480);
nor U40409 (N_40409,N_39066,N_39097);
and U40410 (N_40410,N_38115,N_38008);
xnor U40411 (N_40411,N_39326,N_39435);
nor U40412 (N_40412,N_38924,N_38125);
or U40413 (N_40413,N_39487,N_38456);
xnor U40414 (N_40414,N_39104,N_38379);
and U40415 (N_40415,N_38679,N_39534);
xnor U40416 (N_40416,N_39579,N_38531);
and U40417 (N_40417,N_38313,N_38853);
xor U40418 (N_40418,N_39110,N_38333);
nand U40419 (N_40419,N_39762,N_38267);
or U40420 (N_40420,N_39289,N_38318);
or U40421 (N_40421,N_39217,N_38237);
xor U40422 (N_40422,N_38084,N_39046);
or U40423 (N_40423,N_38868,N_38835);
nor U40424 (N_40424,N_39513,N_38761);
xor U40425 (N_40425,N_39458,N_38239);
and U40426 (N_40426,N_38766,N_39459);
nand U40427 (N_40427,N_39591,N_39578);
and U40428 (N_40428,N_38288,N_39989);
nand U40429 (N_40429,N_39504,N_38004);
nand U40430 (N_40430,N_39672,N_39493);
nor U40431 (N_40431,N_38624,N_39527);
xor U40432 (N_40432,N_39760,N_39281);
nand U40433 (N_40433,N_39157,N_39930);
or U40434 (N_40434,N_39521,N_39022);
nand U40435 (N_40435,N_39245,N_39079);
nor U40436 (N_40436,N_39446,N_39840);
and U40437 (N_40437,N_38923,N_38192);
xnor U40438 (N_40438,N_38559,N_38600);
and U40439 (N_40439,N_38752,N_38262);
and U40440 (N_40440,N_38821,N_39559);
nor U40441 (N_40441,N_39229,N_38498);
nor U40442 (N_40442,N_38345,N_39669);
nor U40443 (N_40443,N_39580,N_38501);
and U40444 (N_40444,N_39306,N_38836);
and U40445 (N_40445,N_39017,N_39859);
nor U40446 (N_40446,N_38331,N_38606);
xor U40447 (N_40447,N_38953,N_39069);
or U40448 (N_40448,N_38819,N_39889);
or U40449 (N_40449,N_38155,N_38595);
nand U40450 (N_40450,N_38893,N_39894);
xnor U40451 (N_40451,N_39955,N_39678);
nand U40452 (N_40452,N_38564,N_38861);
and U40453 (N_40453,N_39112,N_38962);
and U40454 (N_40454,N_38674,N_38560);
or U40455 (N_40455,N_39032,N_39751);
and U40456 (N_40456,N_39436,N_39967);
and U40457 (N_40457,N_38305,N_38320);
and U40458 (N_40458,N_38454,N_39225);
and U40459 (N_40459,N_38885,N_39598);
nand U40460 (N_40460,N_39033,N_38959);
xor U40461 (N_40461,N_39575,N_39508);
and U40462 (N_40462,N_39700,N_39741);
nand U40463 (N_40463,N_39343,N_38076);
nand U40464 (N_40464,N_39582,N_38398);
nor U40465 (N_40465,N_39898,N_38654);
and U40466 (N_40466,N_38374,N_38044);
and U40467 (N_40467,N_39597,N_38290);
and U40468 (N_40468,N_39515,N_39133);
xnor U40469 (N_40469,N_39526,N_38198);
xor U40470 (N_40470,N_39589,N_38184);
and U40471 (N_40471,N_38463,N_39396);
nand U40472 (N_40472,N_38850,N_38701);
nand U40473 (N_40473,N_39052,N_38153);
nand U40474 (N_40474,N_38586,N_38736);
xor U40475 (N_40475,N_38326,N_39363);
xor U40476 (N_40476,N_38158,N_39815);
nor U40477 (N_40477,N_38517,N_38216);
and U40478 (N_40478,N_39674,N_38416);
and U40479 (N_40479,N_39943,N_39009);
and U40480 (N_40480,N_39492,N_39693);
nand U40481 (N_40481,N_39781,N_38042);
nand U40482 (N_40482,N_38512,N_38879);
nor U40483 (N_40483,N_38495,N_39757);
xnor U40484 (N_40484,N_39726,N_38510);
nor U40485 (N_40485,N_39666,N_38046);
xor U40486 (N_40486,N_39657,N_38789);
and U40487 (N_40487,N_38573,N_38003);
and U40488 (N_40488,N_39198,N_39001);
and U40489 (N_40489,N_38210,N_38576);
nor U40490 (N_40490,N_39180,N_38551);
and U40491 (N_40491,N_39634,N_38391);
and U40492 (N_40492,N_39384,N_39662);
and U40493 (N_40493,N_39082,N_39811);
nor U40494 (N_40494,N_38540,N_39297);
xnor U40495 (N_40495,N_39162,N_38831);
xnor U40496 (N_40496,N_39128,N_39138);
nor U40497 (N_40497,N_39719,N_39215);
and U40498 (N_40498,N_38069,N_39190);
and U40499 (N_40499,N_39519,N_39166);
xor U40500 (N_40500,N_38359,N_39992);
nand U40501 (N_40501,N_38306,N_39181);
nand U40502 (N_40502,N_39299,N_38085);
nor U40503 (N_40503,N_38173,N_38468);
and U40504 (N_40504,N_39221,N_39738);
nand U40505 (N_40505,N_38018,N_39551);
and U40506 (N_40506,N_38663,N_39111);
or U40507 (N_40507,N_39445,N_38093);
nand U40508 (N_40508,N_38747,N_38307);
and U40509 (N_40509,N_39556,N_39545);
or U40510 (N_40510,N_38720,N_39637);
nand U40511 (N_40511,N_38954,N_38751);
nand U40512 (N_40512,N_38916,N_39244);
or U40513 (N_40513,N_39401,N_38482);
xnor U40514 (N_40514,N_38928,N_38087);
nor U40515 (N_40515,N_39083,N_38838);
xnor U40516 (N_40516,N_39584,N_39073);
nand U40517 (N_40517,N_39251,N_38759);
xnor U40518 (N_40518,N_38714,N_39249);
nand U40519 (N_40519,N_39810,N_38171);
and U40520 (N_40520,N_39482,N_39236);
xnor U40521 (N_40521,N_38455,N_38686);
nor U40522 (N_40522,N_38872,N_39986);
nor U40523 (N_40523,N_38484,N_38478);
and U40524 (N_40524,N_39648,N_38050);
or U40525 (N_40525,N_39747,N_38818);
and U40526 (N_40526,N_38261,N_38103);
nand U40527 (N_40527,N_39649,N_39365);
nor U40528 (N_40528,N_39942,N_39235);
nor U40529 (N_40529,N_38240,N_39813);
nor U40530 (N_40530,N_38566,N_38915);
nor U40531 (N_40531,N_38502,N_38880);
or U40532 (N_40532,N_39263,N_39886);
nand U40533 (N_40533,N_38072,N_38732);
nand U40534 (N_40534,N_38611,N_39100);
or U40535 (N_40535,N_39947,N_39434);
xnor U40536 (N_40536,N_38696,N_39059);
and U40537 (N_40537,N_38159,N_39155);
xnor U40538 (N_40538,N_38124,N_38279);
or U40539 (N_40539,N_39324,N_39577);
and U40540 (N_40540,N_39586,N_39987);
and U40541 (N_40541,N_39337,N_39404);
or U40542 (N_40542,N_38036,N_39084);
nor U40543 (N_40543,N_39218,N_38656);
nor U40544 (N_40544,N_39918,N_38584);
or U40545 (N_40545,N_39570,N_38763);
nor U40546 (N_40546,N_38599,N_39047);
xnor U40547 (N_40547,N_39689,N_39793);
or U40548 (N_40548,N_39078,N_38263);
xnor U40549 (N_40549,N_39312,N_39880);
nor U40550 (N_40550,N_39682,N_38614);
xnor U40551 (N_40551,N_38980,N_39171);
and U40552 (N_40552,N_39814,N_38167);
or U40553 (N_40553,N_39916,N_38381);
nand U40554 (N_40554,N_38054,N_39161);
or U40555 (N_40555,N_38515,N_39266);
xor U40556 (N_40556,N_39502,N_38122);
or U40557 (N_40557,N_38045,N_38065);
and U40558 (N_40558,N_38098,N_39831);
xnor U40559 (N_40559,N_39472,N_39345);
nor U40560 (N_40560,N_39510,N_39015);
xnor U40561 (N_40561,N_39045,N_38185);
nor U40562 (N_40562,N_38815,N_39116);
and U40563 (N_40563,N_39016,N_39633);
nand U40564 (N_40564,N_39014,N_38489);
nand U40565 (N_40565,N_38726,N_38976);
xnor U40566 (N_40566,N_38617,N_39408);
and U40567 (N_40567,N_38119,N_38592);
xor U40568 (N_40568,N_38396,N_39933);
nand U40569 (N_40569,N_39170,N_39685);
or U40570 (N_40570,N_38395,N_39444);
xnor U40571 (N_40571,N_38549,N_38371);
or U40572 (N_40572,N_38756,N_38492);
nand U40573 (N_40573,N_38610,N_38780);
xor U40574 (N_40574,N_38627,N_38620);
and U40575 (N_40575,N_38770,N_38824);
xnor U40576 (N_40576,N_39361,N_38887);
nand U40577 (N_40577,N_38349,N_39470);
and U40578 (N_40578,N_39895,N_38000);
and U40579 (N_40579,N_38104,N_39856);
nand U40580 (N_40580,N_39203,N_39381);
nand U40581 (N_40581,N_38771,N_38796);
nor U40582 (N_40582,N_38281,N_39291);
nor U40583 (N_40583,N_39692,N_39623);
nand U40584 (N_40584,N_39207,N_38188);
xor U40585 (N_40585,N_38163,N_39714);
and U40586 (N_40586,N_38294,N_39961);
xor U40587 (N_40587,N_38626,N_39703);
xnor U40588 (N_40588,N_39490,N_39265);
and U40589 (N_40589,N_38724,N_39152);
nand U40590 (N_40590,N_38914,N_39808);
and U40591 (N_40591,N_38029,N_38634);
xor U40592 (N_40592,N_38533,N_38177);
xnor U40593 (N_40593,N_38570,N_39238);
and U40594 (N_40594,N_38854,N_38989);
xnor U40595 (N_40595,N_38208,N_38922);
nor U40596 (N_40596,N_38397,N_39264);
and U40597 (N_40597,N_38077,N_38405);
nor U40598 (N_40598,N_39806,N_38180);
and U40599 (N_40599,N_39891,N_39583);
and U40600 (N_40600,N_38270,N_38581);
nand U40601 (N_40601,N_39823,N_38015);
or U40602 (N_40602,N_39901,N_38729);
xor U40603 (N_40603,N_38825,N_38619);
and U40604 (N_40604,N_38768,N_39590);
nand U40605 (N_40605,N_39285,N_38472);
nand U40606 (N_40606,N_38319,N_38859);
and U40607 (N_40607,N_39965,N_39543);
and U40608 (N_40608,N_38334,N_39819);
nor U40609 (N_40609,N_39391,N_39794);
nor U40610 (N_40610,N_38082,N_38344);
xnor U40611 (N_40611,N_39518,N_39644);
nor U40612 (N_40612,N_38206,N_39140);
and U40613 (N_40613,N_38668,N_39442);
and U40614 (N_40614,N_39471,N_39402);
xor U40615 (N_40615,N_38999,N_39501);
and U40616 (N_40616,N_39232,N_39453);
xnor U40617 (N_40617,N_38943,N_38426);
nand U40618 (N_40618,N_38362,N_38175);
xor U40619 (N_40619,N_38556,N_39077);
and U40620 (N_40620,N_38864,N_39270);
and U40621 (N_40621,N_39351,N_38565);
or U40622 (N_40622,N_39154,N_38833);
nand U40623 (N_40623,N_39905,N_38812);
and U40624 (N_40624,N_39287,N_38010);
nand U40625 (N_40625,N_38116,N_39222);
or U40626 (N_40626,N_38259,N_39841);
nand U40627 (N_40627,N_38494,N_39604);
nor U40628 (N_40628,N_38097,N_39432);
nand U40629 (N_40629,N_39681,N_38765);
xor U40630 (N_40630,N_38289,N_38977);
xnor U40631 (N_40631,N_39121,N_38001);
and U40632 (N_40632,N_38808,N_38338);
nand U40633 (N_40633,N_38436,N_38978);
nand U40634 (N_40634,N_39060,N_38241);
nand U40635 (N_40635,N_38574,N_38474);
and U40636 (N_40636,N_38174,N_38390);
xnor U40637 (N_40637,N_38552,N_39763);
or U40638 (N_40638,N_38056,N_39074);
xnor U40639 (N_40639,N_39368,N_38332);
xnor U40640 (N_40640,N_38235,N_38181);
xor U40641 (N_40641,N_39426,N_38055);
nor U40642 (N_40642,N_39592,N_38190);
xor U40643 (N_40643,N_38132,N_39596);
xnor U40644 (N_40644,N_38433,N_38470);
or U40645 (N_40645,N_38209,N_39477);
xor U40646 (N_40646,N_38404,N_39226);
or U40647 (N_40647,N_39058,N_38979);
nor U40648 (N_40648,N_39332,N_39233);
nand U40649 (N_40649,N_38350,N_38578);
xor U40650 (N_40650,N_38982,N_39430);
nand U40651 (N_40651,N_38993,N_38058);
and U40652 (N_40652,N_39746,N_38867);
nand U40653 (N_40653,N_38347,N_38882);
or U40654 (N_40654,N_39352,N_38123);
nand U40655 (N_40655,N_39835,N_39803);
and U40656 (N_40656,N_38944,N_38423);
nand U40657 (N_40657,N_38207,N_38607);
or U40658 (N_40658,N_38376,N_39664);
nand U40659 (N_40659,N_39173,N_38878);
or U40660 (N_40660,N_39002,N_39698);
or U40661 (N_40661,N_39914,N_39796);
nand U40662 (N_40662,N_39119,N_39020);
or U40663 (N_40663,N_38750,N_39826);
nand U40664 (N_40664,N_39912,N_39917);
or U40665 (N_40665,N_38965,N_39663);
and U40666 (N_40666,N_39328,N_38921);
and U40667 (N_40667,N_38542,N_38774);
or U40668 (N_40668,N_39585,N_38589);
nand U40669 (N_40669,N_39403,N_38949);
xor U40670 (N_40670,N_38033,N_39356);
nand U40671 (N_40671,N_39636,N_38070);
or U40672 (N_40672,N_39197,N_38092);
nand U40673 (N_40673,N_38427,N_38827);
xor U40674 (N_40674,N_38913,N_39852);
xor U40675 (N_40675,N_39158,N_38546);
xor U40676 (N_40676,N_39124,N_39206);
nand U40677 (N_40677,N_39900,N_38807);
nor U40678 (N_40678,N_38583,N_39039);
nor U40679 (N_40679,N_39184,N_38302);
xor U40680 (N_40680,N_39935,N_39089);
and U40681 (N_40681,N_39655,N_39548);
nand U40682 (N_40682,N_38039,N_38523);
xnor U40683 (N_40683,N_38524,N_39787);
nand U40684 (N_40684,N_39007,N_39661);
xnor U40685 (N_40685,N_38609,N_39980);
nand U40686 (N_40686,N_39296,N_39231);
or U40687 (N_40687,N_39652,N_38466);
xnor U40688 (N_40688,N_39367,N_38716);
xor U40689 (N_40689,N_39937,N_38403);
nand U40690 (N_40690,N_39024,N_38643);
nor U40691 (N_40691,N_39802,N_39941);
and U40692 (N_40692,N_39214,N_38230);
xnor U40693 (N_40693,N_38342,N_39334);
nand U40694 (N_40694,N_39208,N_39995);
and U40695 (N_40695,N_38219,N_39295);
nor U40696 (N_40696,N_38945,N_39828);
nor U40697 (N_40697,N_39602,N_38642);
nor U40698 (N_40698,N_39651,N_39062);
and U40699 (N_40699,N_39660,N_39837);
xor U40700 (N_40700,N_38248,N_39372);
xor U40701 (N_40701,N_39107,N_38557);
nor U40702 (N_40702,N_38748,N_38246);
nor U40703 (N_40703,N_38131,N_39130);
nor U40704 (N_40704,N_38805,N_38178);
nand U40705 (N_40705,N_38757,N_39722);
nand U40706 (N_40706,N_39820,N_39627);
xor U40707 (N_40707,N_38449,N_38555);
nand U40708 (N_40708,N_38998,N_39766);
nand U40709 (N_40709,N_38249,N_39694);
and U40710 (N_40710,N_39194,N_39071);
and U40711 (N_40711,N_38157,N_38446);
nand U40712 (N_40712,N_39524,N_39565);
nand U40713 (N_40713,N_39610,N_39424);
and U40714 (N_40714,N_38437,N_39250);
nand U40715 (N_40715,N_39309,N_38587);
and U40716 (N_40716,N_39774,N_38164);
nor U40717 (N_40717,N_39860,N_38890);
nor U40718 (N_40718,N_39397,N_38727);
and U40719 (N_40719,N_39629,N_39129);
and U40720 (N_40720,N_39635,N_38813);
and U40721 (N_40721,N_38675,N_39462);
xnor U40722 (N_40722,N_38461,N_39146);
or U40723 (N_40723,N_38513,N_38064);
nor U40724 (N_40724,N_38100,N_39473);
or U40725 (N_40725,N_38411,N_38650);
nor U40726 (N_40726,N_38410,N_39123);
xnor U40727 (N_40727,N_38881,N_38487);
nand U40728 (N_40728,N_38442,N_38548);
and U40729 (N_40729,N_39159,N_38081);
or U40730 (N_40730,N_39934,N_38687);
xnor U40731 (N_40731,N_39641,N_38508);
or U40732 (N_40732,N_39523,N_39148);
nand U40733 (N_40733,N_38186,N_38658);
and U40734 (N_40734,N_38339,N_38535);
nor U40735 (N_40735,N_38537,N_39640);
nand U40736 (N_40736,N_39709,N_38088);
nand U40737 (N_40737,N_39256,N_39145);
xnor U40738 (N_40738,N_39643,N_38971);
or U40739 (N_40739,N_38335,N_38120);
and U40740 (N_40740,N_38742,N_39539);
nor U40741 (N_40741,N_38068,N_38299);
nor U40742 (N_40742,N_38764,N_38691);
and U40743 (N_40743,N_39276,N_38220);
nor U40744 (N_40744,N_38585,N_38744);
and U40745 (N_40745,N_38788,N_38649);
or U40746 (N_40746,N_39160,N_38212);
and U40747 (N_40747,N_38252,N_38994);
nand U40748 (N_40748,N_38682,N_38534);
nor U40749 (N_40749,N_38389,N_38075);
nand U40750 (N_40750,N_38011,N_38032);
nand U40751 (N_40751,N_39268,N_38380);
nor U40752 (N_40752,N_39483,N_39569);
xnor U40753 (N_40753,N_38273,N_39165);
xnor U40754 (N_40754,N_38497,N_38664);
nor U40755 (N_40755,N_38074,N_38558);
or U40756 (N_40756,N_38848,N_38238);
and U40757 (N_40757,N_39978,N_39964);
nor U40758 (N_40758,N_39829,N_39573);
or U40759 (N_40759,N_38707,N_39786);
nor U40760 (N_40760,N_38659,N_38760);
nand U40761 (N_40761,N_38680,N_38464);
or U40762 (N_40762,N_39255,N_39724);
nor U40763 (N_40763,N_38066,N_38612);
and U40764 (N_40764,N_39451,N_38622);
nand U40765 (N_40765,N_39697,N_38547);
nor U40766 (N_40766,N_38191,N_39223);
and U40767 (N_40767,N_38904,N_39468);
xnor U40768 (N_40768,N_38903,N_38027);
and U40769 (N_40769,N_38590,N_38772);
and U40770 (N_40770,N_38452,N_39191);
xor U40771 (N_40771,N_39846,N_38802);
nor U40772 (N_40772,N_38777,N_39449);
nor U40773 (N_40773,N_38907,N_39260);
nor U40774 (N_40774,N_39304,N_38179);
xor U40775 (N_40775,N_39175,N_38005);
or U40776 (N_40776,N_38828,N_39522);
and U40777 (N_40777,N_39463,N_39975);
or U40778 (N_40778,N_38671,N_38233);
nand U40779 (N_40779,N_38602,N_38504);
or U40780 (N_40780,N_39691,N_38149);
and U40781 (N_40781,N_39329,N_38114);
xor U40782 (N_40782,N_38530,N_39879);
xor U40783 (N_40783,N_38465,N_38625);
nor U40784 (N_40784,N_38444,N_38193);
nand U40785 (N_40785,N_39484,N_38182);
nand U40786 (N_40786,N_38960,N_38137);
and U40787 (N_40787,N_39728,N_38256);
nand U40788 (N_40788,N_38932,N_38356);
and U40789 (N_40789,N_38955,N_38421);
nor U40790 (N_40790,N_38754,N_39993);
xnor U40791 (N_40791,N_39348,N_38330);
nor U40792 (N_40792,N_38301,N_38991);
nor U40793 (N_40793,N_38837,N_39240);
or U40794 (N_40794,N_39085,N_38983);
nor U40795 (N_40795,N_38101,N_38106);
and U40796 (N_40796,N_39771,N_38975);
or U40797 (N_40797,N_39283,N_39797);
nor U40798 (N_40798,N_39957,N_38830);
nor U40799 (N_40799,N_39999,N_39094);
xor U40800 (N_40800,N_38107,N_39120);
nand U40801 (N_40801,N_38702,N_38635);
and U40802 (N_40802,N_39888,N_38202);
xor U40803 (N_40803,N_39670,N_38721);
and U40804 (N_40804,N_38031,N_39568);
or U40805 (N_40805,N_38672,N_39035);
nand U40806 (N_40806,N_38425,N_39293);
nand U40807 (N_40807,N_38507,N_38615);
or U40808 (N_40808,N_38447,N_39601);
xor U40809 (N_40809,N_39061,N_39005);
or U40810 (N_40810,N_38140,N_39603);
xnor U40811 (N_40811,N_38364,N_39736);
xnor U40812 (N_40812,N_39977,N_38681);
nor U40813 (N_40813,N_39076,N_38877);
xor U40814 (N_40814,N_39353,N_39923);
or U40815 (N_40815,N_39882,N_38060);
and U40816 (N_40816,N_38309,N_38912);
nor U40817 (N_40817,N_38413,N_39800);
xor U40818 (N_40818,N_39323,N_39667);
and U40819 (N_40819,N_38822,N_38873);
and U40820 (N_40820,N_39866,N_38019);
xnor U40821 (N_40821,N_38667,N_39201);
and U40822 (N_40822,N_39788,N_38415);
or U40823 (N_40823,N_39417,N_39008);
xnor U40824 (N_40824,N_38245,N_38422);
xnor U40825 (N_40825,N_39172,N_39721);
and U40826 (N_40826,N_38406,N_38459);
nor U40827 (N_40827,N_39777,N_39479);
and U40828 (N_40828,N_38963,N_38346);
nor U40829 (N_40829,N_39702,N_38917);
or U40830 (N_40830,N_38417,N_38271);
nor U40831 (N_40831,N_38938,N_39675);
and U40832 (N_40832,N_38336,N_38408);
nand U40833 (N_40833,N_39307,N_39910);
or U40834 (N_40834,N_38929,N_38525);
nand U40835 (N_40835,N_39922,N_38866);
or U40836 (N_40836,N_39958,N_38996);
xnor U40837 (N_40837,N_39749,N_38639);
or U40838 (N_40838,N_38372,N_38518);
or U40839 (N_40839,N_39096,N_38666);
nand U40840 (N_40840,N_39075,N_38052);
and U40841 (N_40841,N_39049,N_39371);
and U40842 (N_40842,N_38509,N_39779);
nor U40843 (N_40843,N_39314,N_39780);
and U40844 (N_40844,N_38013,N_38553);
and U40845 (N_40845,N_39626,N_39622);
xnor U40846 (N_40846,N_38734,N_38034);
or U40847 (N_40847,N_39981,N_38303);
nand U40848 (N_40848,N_39347,N_38095);
nor U40849 (N_40849,N_39422,N_38544);
nor U40850 (N_40850,N_38007,N_38719);
nand U40851 (N_40851,N_38471,N_38152);
nand U40852 (N_40852,N_39056,N_38438);
and U40853 (N_40853,N_39425,N_38375);
or U40854 (N_40854,N_39440,N_38247);
nand U40855 (N_40855,N_38698,N_39824);
nor U40856 (N_40856,N_38223,N_39744);
nand U40857 (N_40857,N_39115,N_39963);
xnor U40858 (N_40858,N_38660,N_38280);
or U40859 (N_40859,N_38740,N_39486);
and U40860 (N_40860,N_39574,N_38030);
and U40861 (N_40861,N_39395,N_38860);
and U40862 (N_40862,N_39366,N_39954);
nor U40863 (N_40863,N_39466,N_39587);
nor U40864 (N_40864,N_38205,N_38845);
or U40865 (N_40865,N_38699,N_39320);
nand U40866 (N_40866,N_38251,N_39982);
xor U40867 (N_40867,N_38918,N_38948);
nor U40868 (N_40868,N_39469,N_39679);
nor U40869 (N_40869,N_38952,N_38689);
and U40870 (N_40870,N_38287,N_38169);
or U40871 (N_40871,N_39897,N_38641);
nor U40872 (N_40872,N_39706,N_39871);
nand U40873 (N_40873,N_39216,N_38908);
nand U40874 (N_40874,N_39758,N_38648);
or U40875 (N_40875,N_39429,N_39505);
and U40876 (N_40876,N_38769,N_39938);
and U40877 (N_40877,N_39716,N_39114);
or U40878 (N_40878,N_39532,N_39713);
nand U40879 (N_40879,N_39687,N_39438);
xnor U40880 (N_40880,N_38317,N_39383);
and U40881 (N_40881,N_38762,N_38988);
nor U40882 (N_40882,N_38394,N_38529);
and U40883 (N_40883,N_38545,N_38343);
nor U40884 (N_40884,N_39031,N_39188);
xnor U40885 (N_40885,N_38316,N_39848);
nor U40886 (N_40886,N_38990,N_39355);
xnor U40887 (N_40887,N_38048,N_38016);
or U40888 (N_40888,N_38746,N_39398);
xor U40889 (N_40889,N_38435,N_38865);
nand U40890 (N_40890,N_38820,N_38296);
or U40891 (N_40891,N_38275,N_38631);
nand U40892 (N_40892,N_39286,N_38105);
and U40893 (N_40893,N_39421,N_38197);
nor U40894 (N_40894,N_39182,N_39653);
xor U40895 (N_40895,N_39812,N_39743);
xnor U40896 (N_40896,N_39378,N_38653);
or U40897 (N_40897,N_38035,N_38266);
or U40898 (N_40898,N_38419,N_38089);
or U40899 (N_40899,N_39845,N_39710);
or U40900 (N_40900,N_38715,N_39951);
xnor U40901 (N_40901,N_39921,N_38189);
nand U40902 (N_40902,N_39616,N_39132);
xnor U40903 (N_40903,N_38711,N_39873);
or U40904 (N_40904,N_38274,N_39799);
nor U40905 (N_40905,N_38024,N_38968);
nand U40906 (N_40906,N_39790,N_39028);
and U40907 (N_40907,N_39514,N_39338);
nand U40908 (N_40908,N_38428,N_38801);
or U40909 (N_40909,N_38328,N_39357);
nor U40910 (N_40910,N_38514,N_39884);
and U40911 (N_40911,N_39588,N_39386);
nand U40912 (N_40912,N_38324,N_38493);
or U40913 (N_40913,N_38961,N_38057);
xor U40914 (N_40914,N_39040,N_39053);
nor U40915 (N_40915,N_39211,N_38138);
or U40916 (N_40916,N_39676,N_38895);
nand U40917 (N_40917,N_39576,N_39948);
xnor U40918 (N_40918,N_39768,N_38392);
or U40919 (N_40919,N_39529,N_38931);
nand U40920 (N_40920,N_38628,N_38695);
or U40921 (N_40921,N_39242,N_38519);
and U40922 (N_40922,N_39237,N_39595);
nor U40923 (N_40923,N_39167,N_38352);
and U40924 (N_40924,N_38676,N_39090);
and U40925 (N_40925,N_39354,N_38094);
xnor U40926 (N_40926,N_38972,N_39960);
nor U40927 (N_40927,N_38439,N_38717);
nor U40928 (N_40928,N_38221,N_38577);
nand U40929 (N_40929,N_39143,N_39410);
or U40930 (N_40930,N_38203,N_38361);
or U40931 (N_40931,N_39733,N_39411);
and U40932 (N_40932,N_38199,N_39278);
and U40933 (N_40933,N_38443,N_38401);
nand U40934 (N_40934,N_38384,N_38127);
or U40935 (N_40935,N_39818,N_39478);
nor U40936 (N_40936,N_38300,N_38321);
or U40937 (N_40937,N_38785,N_38340);
nand U40938 (N_40938,N_38144,N_39553);
nor U40939 (N_40939,N_38630,N_39968);
or U40940 (N_40940,N_38855,N_39313);
nand U40941 (N_40941,N_38369,N_38172);
and U40942 (N_40942,N_38652,N_38420);
or U40943 (N_40943,N_39821,N_38636);
and U40944 (N_40944,N_39740,N_39770);
nand U40945 (N_40945,N_38062,N_39940);
and U40946 (N_40946,N_39903,N_38156);
xor U40947 (N_40947,N_38110,N_39042);
and U40948 (N_40948,N_39034,N_38148);
and U40949 (N_40949,N_39108,N_39520);
nor U40950 (N_40950,N_39614,N_39359);
xor U40951 (N_40951,N_39036,N_39783);
xor U40952 (N_40952,N_38973,N_39782);
or U40953 (N_40953,N_39387,N_38014);
nor U40954 (N_40954,N_38467,N_38613);
xor U40955 (N_40955,N_39346,N_39327);
nand U40956 (N_40956,N_39377,N_38594);
or U40957 (N_40957,N_38925,N_39344);
or U40958 (N_40958,N_38876,N_39183);
and U40959 (N_40959,N_38823,N_38481);
nor U40960 (N_40960,N_39431,N_38061);
xor U40961 (N_40961,N_38432,N_38572);
or U40962 (N_40962,N_38323,N_38071);
and U40963 (N_40963,N_38448,N_39064);
or U40964 (N_40964,N_38136,N_39259);
xor U40965 (N_40965,N_38126,N_39274);
nand U40966 (N_40966,N_39187,N_39767);
and U40967 (N_40967,N_39769,N_38161);
xnor U40968 (N_40968,N_39456,N_38142);
xor U40969 (N_40969,N_39406,N_39230);
or U40970 (N_40970,N_39419,N_38803);
nor U40971 (N_40971,N_38272,N_38969);
xor U40972 (N_40972,N_39612,N_39708);
nand U40973 (N_40973,N_39063,N_39248);
nand U40974 (N_40974,N_38293,N_39533);
nand U40975 (N_40975,N_39625,N_38941);
xnor U40976 (N_40976,N_38322,N_39549);
and U40977 (N_40977,N_39939,N_39854);
xnor U40978 (N_40978,N_38226,N_38166);
nor U40979 (N_40979,N_38213,N_38987);
and U40980 (N_40980,N_39807,N_38440);
or U40981 (N_40981,N_39517,N_39566);
or U40982 (N_40982,N_39454,N_38480);
or U40983 (N_40983,N_39489,N_39204);
xnor U40984 (N_40984,N_39193,N_38934);
nor U40985 (N_40985,N_38187,N_39292);
nand U40986 (N_40986,N_38571,N_38067);
nand U40987 (N_40987,N_39497,N_39448);
and U40988 (N_40988,N_39013,N_39547);
nor U40989 (N_40989,N_38257,N_38215);
and U40990 (N_40990,N_39908,N_39220);
and U40991 (N_40991,N_38041,N_39690);
and U40992 (N_40992,N_38377,N_39699);
nand U40993 (N_40993,N_39012,N_39179);
or U40994 (N_40994,N_38898,N_39926);
nor U40995 (N_40995,N_38382,N_39428);
nor U40996 (N_40996,N_38735,N_38704);
nand U40997 (N_40997,N_38134,N_38703);
nand U40998 (N_40998,N_39868,N_38739);
or U40999 (N_40999,N_39321,N_38102);
nor U41000 (N_41000,N_39593,N_38300);
nor U41001 (N_41001,N_39303,N_39287);
nor U41002 (N_41002,N_38169,N_39167);
and U41003 (N_41003,N_39789,N_38569);
and U41004 (N_41004,N_39531,N_39955);
and U41005 (N_41005,N_38297,N_39407);
xor U41006 (N_41006,N_39947,N_38234);
nor U41007 (N_41007,N_38393,N_38139);
nand U41008 (N_41008,N_38737,N_39311);
or U41009 (N_41009,N_38969,N_38717);
nand U41010 (N_41010,N_39480,N_38872);
and U41011 (N_41011,N_39780,N_38128);
nand U41012 (N_41012,N_39223,N_38935);
and U41013 (N_41013,N_39629,N_38781);
nand U41014 (N_41014,N_39938,N_38696);
nand U41015 (N_41015,N_38419,N_39370);
xor U41016 (N_41016,N_39652,N_38176);
xor U41017 (N_41017,N_39260,N_38570);
or U41018 (N_41018,N_38696,N_38660);
or U41019 (N_41019,N_39144,N_38436);
and U41020 (N_41020,N_38694,N_39382);
or U41021 (N_41021,N_38450,N_39362);
nand U41022 (N_41022,N_39333,N_39102);
and U41023 (N_41023,N_38577,N_39925);
nand U41024 (N_41024,N_39193,N_39680);
nor U41025 (N_41025,N_39114,N_38809);
and U41026 (N_41026,N_38333,N_39646);
nand U41027 (N_41027,N_39540,N_38921);
and U41028 (N_41028,N_39841,N_38062);
xnor U41029 (N_41029,N_39882,N_39121);
xor U41030 (N_41030,N_39448,N_39943);
and U41031 (N_41031,N_39765,N_38926);
xnor U41032 (N_41032,N_38165,N_39066);
and U41033 (N_41033,N_39558,N_39043);
nor U41034 (N_41034,N_39486,N_39351);
nand U41035 (N_41035,N_39475,N_39913);
and U41036 (N_41036,N_38331,N_39913);
nand U41037 (N_41037,N_39602,N_38211);
and U41038 (N_41038,N_39940,N_39823);
or U41039 (N_41039,N_39881,N_39893);
nand U41040 (N_41040,N_39295,N_38393);
or U41041 (N_41041,N_39843,N_39074);
nor U41042 (N_41042,N_39918,N_39008);
or U41043 (N_41043,N_38082,N_38463);
and U41044 (N_41044,N_38496,N_39391);
nand U41045 (N_41045,N_38819,N_38637);
xor U41046 (N_41046,N_38492,N_39652);
nor U41047 (N_41047,N_39961,N_38521);
or U41048 (N_41048,N_38456,N_38881);
and U41049 (N_41049,N_38042,N_39392);
nand U41050 (N_41050,N_39292,N_38721);
nor U41051 (N_41051,N_38103,N_39643);
nor U41052 (N_41052,N_39261,N_39206);
and U41053 (N_41053,N_38358,N_38686);
or U41054 (N_41054,N_38959,N_38975);
xor U41055 (N_41055,N_39997,N_39492);
nor U41056 (N_41056,N_39465,N_39933);
and U41057 (N_41057,N_39892,N_39434);
nor U41058 (N_41058,N_39328,N_38161);
xnor U41059 (N_41059,N_39149,N_38330);
or U41060 (N_41060,N_38562,N_39692);
and U41061 (N_41061,N_38210,N_38964);
nor U41062 (N_41062,N_38256,N_38466);
and U41063 (N_41063,N_38645,N_38931);
xor U41064 (N_41064,N_39335,N_38092);
or U41065 (N_41065,N_39342,N_39173);
xnor U41066 (N_41066,N_39954,N_38195);
nor U41067 (N_41067,N_39793,N_38923);
xnor U41068 (N_41068,N_38318,N_38306);
and U41069 (N_41069,N_39750,N_38692);
or U41070 (N_41070,N_38468,N_38664);
or U41071 (N_41071,N_39747,N_38872);
xor U41072 (N_41072,N_38623,N_39733);
nand U41073 (N_41073,N_38055,N_39061);
xor U41074 (N_41074,N_39816,N_38093);
and U41075 (N_41075,N_39292,N_39619);
nand U41076 (N_41076,N_38595,N_39269);
nor U41077 (N_41077,N_38854,N_38693);
nor U41078 (N_41078,N_38986,N_39558);
nor U41079 (N_41079,N_38437,N_39047);
and U41080 (N_41080,N_38965,N_38802);
and U41081 (N_41081,N_38767,N_39762);
xor U41082 (N_41082,N_38178,N_39245);
xnor U41083 (N_41083,N_39596,N_39145);
nor U41084 (N_41084,N_39541,N_39942);
or U41085 (N_41085,N_39534,N_38595);
nand U41086 (N_41086,N_39946,N_39031);
nor U41087 (N_41087,N_38361,N_38519);
and U41088 (N_41088,N_39770,N_38840);
and U41089 (N_41089,N_38918,N_38389);
and U41090 (N_41090,N_39740,N_38639);
and U41091 (N_41091,N_39070,N_38110);
or U41092 (N_41092,N_39002,N_38839);
xor U41093 (N_41093,N_39734,N_39318);
and U41094 (N_41094,N_39394,N_39178);
or U41095 (N_41095,N_38475,N_38547);
nor U41096 (N_41096,N_38707,N_39897);
or U41097 (N_41097,N_38987,N_39490);
or U41098 (N_41098,N_38141,N_39015);
nand U41099 (N_41099,N_39216,N_39155);
or U41100 (N_41100,N_38885,N_38233);
nand U41101 (N_41101,N_38546,N_39031);
or U41102 (N_41102,N_39877,N_39846);
xnor U41103 (N_41103,N_38479,N_38636);
or U41104 (N_41104,N_39814,N_38568);
or U41105 (N_41105,N_39377,N_38397);
nand U41106 (N_41106,N_39877,N_39823);
nand U41107 (N_41107,N_38773,N_39154);
nor U41108 (N_41108,N_39662,N_38125);
and U41109 (N_41109,N_38567,N_38729);
nand U41110 (N_41110,N_39151,N_39767);
nand U41111 (N_41111,N_38199,N_38432);
xnor U41112 (N_41112,N_38812,N_38947);
xor U41113 (N_41113,N_38022,N_38336);
nor U41114 (N_41114,N_38335,N_38490);
xnor U41115 (N_41115,N_39949,N_39858);
xor U41116 (N_41116,N_39488,N_38298);
xnor U41117 (N_41117,N_38509,N_39586);
or U41118 (N_41118,N_38922,N_39354);
or U41119 (N_41119,N_39169,N_39014);
xnor U41120 (N_41120,N_39054,N_38241);
or U41121 (N_41121,N_38655,N_39259);
nand U41122 (N_41122,N_38628,N_38694);
nor U41123 (N_41123,N_38062,N_39792);
or U41124 (N_41124,N_39305,N_39548);
nor U41125 (N_41125,N_38669,N_39257);
or U41126 (N_41126,N_39552,N_38298);
nor U41127 (N_41127,N_39757,N_38738);
nand U41128 (N_41128,N_38905,N_38024);
xnor U41129 (N_41129,N_39115,N_38970);
and U41130 (N_41130,N_38298,N_38605);
nor U41131 (N_41131,N_39373,N_38685);
and U41132 (N_41132,N_39616,N_39344);
nand U41133 (N_41133,N_39686,N_39159);
and U41134 (N_41134,N_38792,N_38463);
nor U41135 (N_41135,N_38881,N_39688);
and U41136 (N_41136,N_38289,N_38645);
and U41137 (N_41137,N_39280,N_39182);
and U41138 (N_41138,N_39529,N_39151);
nand U41139 (N_41139,N_38076,N_39025);
and U41140 (N_41140,N_39742,N_39331);
nand U41141 (N_41141,N_39860,N_38748);
nor U41142 (N_41142,N_39353,N_39618);
or U41143 (N_41143,N_39450,N_39429);
nor U41144 (N_41144,N_38731,N_38026);
or U41145 (N_41145,N_39639,N_39485);
or U41146 (N_41146,N_38744,N_38010);
and U41147 (N_41147,N_38913,N_39513);
xor U41148 (N_41148,N_39089,N_38870);
nand U41149 (N_41149,N_38840,N_38792);
or U41150 (N_41150,N_38017,N_39809);
or U41151 (N_41151,N_38119,N_38322);
nand U41152 (N_41152,N_38558,N_39084);
or U41153 (N_41153,N_38916,N_38949);
xnor U41154 (N_41154,N_38691,N_38037);
xor U41155 (N_41155,N_38295,N_38692);
or U41156 (N_41156,N_38987,N_39859);
or U41157 (N_41157,N_38624,N_38021);
and U41158 (N_41158,N_38572,N_38609);
nand U41159 (N_41159,N_38561,N_38470);
or U41160 (N_41160,N_38701,N_38085);
and U41161 (N_41161,N_38051,N_39638);
or U41162 (N_41162,N_38087,N_39922);
and U41163 (N_41163,N_38950,N_39127);
nand U41164 (N_41164,N_39703,N_38288);
nor U41165 (N_41165,N_38757,N_38331);
or U41166 (N_41166,N_39161,N_39426);
nand U41167 (N_41167,N_39399,N_38180);
xor U41168 (N_41168,N_38646,N_39944);
xor U41169 (N_41169,N_38869,N_38269);
xor U41170 (N_41170,N_38584,N_39453);
nor U41171 (N_41171,N_38029,N_39302);
and U41172 (N_41172,N_39397,N_39048);
nor U41173 (N_41173,N_38306,N_38847);
nor U41174 (N_41174,N_38235,N_38625);
and U41175 (N_41175,N_39219,N_38731);
nor U41176 (N_41176,N_38499,N_39469);
or U41177 (N_41177,N_38866,N_39827);
or U41178 (N_41178,N_38207,N_38029);
and U41179 (N_41179,N_39259,N_39030);
and U41180 (N_41180,N_39742,N_38933);
nor U41181 (N_41181,N_38325,N_38181);
nor U41182 (N_41182,N_39053,N_38336);
xor U41183 (N_41183,N_39609,N_39975);
xor U41184 (N_41184,N_39240,N_38667);
and U41185 (N_41185,N_38842,N_38224);
xnor U41186 (N_41186,N_39631,N_39442);
and U41187 (N_41187,N_38172,N_39187);
nor U41188 (N_41188,N_39396,N_39724);
and U41189 (N_41189,N_39897,N_38774);
and U41190 (N_41190,N_38463,N_38326);
and U41191 (N_41191,N_39045,N_39965);
xor U41192 (N_41192,N_38054,N_38175);
nor U41193 (N_41193,N_39305,N_39851);
nor U41194 (N_41194,N_38377,N_39145);
or U41195 (N_41195,N_39072,N_38835);
xor U41196 (N_41196,N_39460,N_38244);
and U41197 (N_41197,N_39456,N_38358);
and U41198 (N_41198,N_39929,N_39110);
or U41199 (N_41199,N_38378,N_38535);
nor U41200 (N_41200,N_38772,N_38293);
nand U41201 (N_41201,N_38045,N_39278);
xnor U41202 (N_41202,N_39085,N_39271);
nand U41203 (N_41203,N_39234,N_38952);
nand U41204 (N_41204,N_38739,N_39642);
and U41205 (N_41205,N_39437,N_39677);
and U41206 (N_41206,N_38453,N_38686);
and U41207 (N_41207,N_38045,N_39171);
nand U41208 (N_41208,N_38461,N_39093);
and U41209 (N_41209,N_39543,N_39226);
nand U41210 (N_41210,N_39070,N_38349);
nand U41211 (N_41211,N_39301,N_39068);
nor U41212 (N_41212,N_39270,N_38863);
nor U41213 (N_41213,N_39982,N_39552);
or U41214 (N_41214,N_38791,N_38770);
nand U41215 (N_41215,N_38444,N_39294);
nor U41216 (N_41216,N_39979,N_39345);
nand U41217 (N_41217,N_39854,N_39315);
and U41218 (N_41218,N_38468,N_38226);
nand U41219 (N_41219,N_39513,N_38920);
or U41220 (N_41220,N_38157,N_39005);
nand U41221 (N_41221,N_38702,N_39661);
or U41222 (N_41222,N_38007,N_39149);
and U41223 (N_41223,N_39461,N_39261);
xnor U41224 (N_41224,N_38423,N_38253);
nand U41225 (N_41225,N_39150,N_39249);
or U41226 (N_41226,N_39930,N_39781);
xor U41227 (N_41227,N_38354,N_38526);
and U41228 (N_41228,N_38092,N_39314);
xor U41229 (N_41229,N_38874,N_39130);
and U41230 (N_41230,N_39521,N_39556);
nand U41231 (N_41231,N_38287,N_39130);
xnor U41232 (N_41232,N_39819,N_38238);
xor U41233 (N_41233,N_39859,N_38132);
xor U41234 (N_41234,N_38025,N_39333);
nand U41235 (N_41235,N_38901,N_39350);
nand U41236 (N_41236,N_39351,N_38011);
and U41237 (N_41237,N_38125,N_38001);
nand U41238 (N_41238,N_39269,N_39928);
and U41239 (N_41239,N_39943,N_39378);
or U41240 (N_41240,N_39530,N_38216);
nor U41241 (N_41241,N_38095,N_39124);
or U41242 (N_41242,N_38627,N_39640);
xor U41243 (N_41243,N_39892,N_38484);
or U41244 (N_41244,N_39304,N_38143);
nor U41245 (N_41245,N_38486,N_39678);
nor U41246 (N_41246,N_38489,N_38901);
nand U41247 (N_41247,N_39157,N_38257);
nor U41248 (N_41248,N_38433,N_39394);
xor U41249 (N_41249,N_38427,N_38594);
nand U41250 (N_41250,N_39062,N_39032);
and U41251 (N_41251,N_39368,N_39517);
xnor U41252 (N_41252,N_39749,N_39917);
xnor U41253 (N_41253,N_39829,N_38029);
nor U41254 (N_41254,N_38333,N_39096);
and U41255 (N_41255,N_39834,N_38568);
nand U41256 (N_41256,N_39602,N_38160);
nand U41257 (N_41257,N_39450,N_39146);
nor U41258 (N_41258,N_38601,N_38186);
nand U41259 (N_41259,N_39261,N_38318);
and U41260 (N_41260,N_38363,N_39679);
and U41261 (N_41261,N_39818,N_39286);
and U41262 (N_41262,N_38421,N_38718);
nand U41263 (N_41263,N_38694,N_39786);
nand U41264 (N_41264,N_38016,N_38042);
nand U41265 (N_41265,N_39446,N_38962);
nor U41266 (N_41266,N_38630,N_38361);
nor U41267 (N_41267,N_39650,N_39163);
nor U41268 (N_41268,N_38603,N_38687);
nand U41269 (N_41269,N_38386,N_38224);
xor U41270 (N_41270,N_38250,N_38154);
or U41271 (N_41271,N_39229,N_39722);
nor U41272 (N_41272,N_38474,N_39830);
or U41273 (N_41273,N_39207,N_38733);
xnor U41274 (N_41274,N_38999,N_38521);
nand U41275 (N_41275,N_38645,N_38669);
and U41276 (N_41276,N_39106,N_38701);
xor U41277 (N_41277,N_39294,N_38185);
xnor U41278 (N_41278,N_39417,N_39372);
xor U41279 (N_41279,N_38314,N_38922);
or U41280 (N_41280,N_38569,N_38254);
nor U41281 (N_41281,N_39307,N_39020);
or U41282 (N_41282,N_39179,N_39430);
or U41283 (N_41283,N_38636,N_39652);
xor U41284 (N_41284,N_39561,N_39636);
xor U41285 (N_41285,N_39803,N_39300);
or U41286 (N_41286,N_38704,N_38829);
and U41287 (N_41287,N_38409,N_39637);
xor U41288 (N_41288,N_39778,N_39578);
nand U41289 (N_41289,N_39293,N_38301);
nor U41290 (N_41290,N_38271,N_39214);
xnor U41291 (N_41291,N_39609,N_38901);
xnor U41292 (N_41292,N_39469,N_39123);
or U41293 (N_41293,N_39066,N_39382);
nor U41294 (N_41294,N_39049,N_38214);
xor U41295 (N_41295,N_38985,N_39022);
or U41296 (N_41296,N_39815,N_38733);
nand U41297 (N_41297,N_38132,N_38111);
nor U41298 (N_41298,N_39220,N_38825);
or U41299 (N_41299,N_38528,N_38228);
xor U41300 (N_41300,N_38176,N_38397);
and U41301 (N_41301,N_39769,N_39704);
and U41302 (N_41302,N_38811,N_39273);
nand U41303 (N_41303,N_38925,N_38621);
or U41304 (N_41304,N_38850,N_39574);
nand U41305 (N_41305,N_38018,N_39149);
xnor U41306 (N_41306,N_39938,N_39707);
xor U41307 (N_41307,N_39532,N_38063);
nor U41308 (N_41308,N_39177,N_39024);
and U41309 (N_41309,N_38438,N_39785);
nor U41310 (N_41310,N_39997,N_38933);
nor U41311 (N_41311,N_39450,N_38925);
nor U41312 (N_41312,N_38870,N_38249);
and U41313 (N_41313,N_39326,N_38729);
nor U41314 (N_41314,N_38528,N_38272);
xor U41315 (N_41315,N_38070,N_38445);
and U41316 (N_41316,N_39910,N_38551);
and U41317 (N_41317,N_39321,N_39230);
nand U41318 (N_41318,N_39030,N_38156);
or U41319 (N_41319,N_38462,N_38254);
xor U41320 (N_41320,N_38142,N_39429);
xor U41321 (N_41321,N_39297,N_38437);
nor U41322 (N_41322,N_38564,N_38488);
nor U41323 (N_41323,N_39822,N_39352);
nand U41324 (N_41324,N_39586,N_39537);
and U41325 (N_41325,N_39845,N_38690);
xor U41326 (N_41326,N_39361,N_38332);
or U41327 (N_41327,N_39777,N_38007);
nor U41328 (N_41328,N_38025,N_38703);
and U41329 (N_41329,N_39230,N_38356);
nand U41330 (N_41330,N_38193,N_39119);
xor U41331 (N_41331,N_38917,N_39655);
nor U41332 (N_41332,N_38943,N_39466);
and U41333 (N_41333,N_38013,N_39008);
nand U41334 (N_41334,N_38812,N_39398);
or U41335 (N_41335,N_39132,N_39021);
nand U41336 (N_41336,N_39911,N_38009);
nand U41337 (N_41337,N_38374,N_39880);
xor U41338 (N_41338,N_39697,N_39073);
nor U41339 (N_41339,N_38158,N_38181);
xnor U41340 (N_41340,N_39083,N_39202);
and U41341 (N_41341,N_39964,N_38052);
xor U41342 (N_41342,N_39001,N_39212);
nand U41343 (N_41343,N_39064,N_39645);
xor U41344 (N_41344,N_39657,N_38183);
or U41345 (N_41345,N_39045,N_38771);
nor U41346 (N_41346,N_39469,N_38328);
or U41347 (N_41347,N_38512,N_38747);
nand U41348 (N_41348,N_38749,N_38911);
nor U41349 (N_41349,N_39266,N_39951);
or U41350 (N_41350,N_38082,N_38637);
xor U41351 (N_41351,N_39376,N_39746);
and U41352 (N_41352,N_38114,N_38179);
and U41353 (N_41353,N_39764,N_38955);
nand U41354 (N_41354,N_39678,N_38504);
xor U41355 (N_41355,N_39159,N_38183);
xnor U41356 (N_41356,N_38267,N_39917);
or U41357 (N_41357,N_39135,N_39912);
and U41358 (N_41358,N_39723,N_38863);
xor U41359 (N_41359,N_39669,N_39450);
and U41360 (N_41360,N_38155,N_38406);
or U41361 (N_41361,N_39956,N_38428);
or U41362 (N_41362,N_39344,N_38000);
xnor U41363 (N_41363,N_38755,N_38261);
nand U41364 (N_41364,N_39348,N_38210);
nor U41365 (N_41365,N_39617,N_38866);
nand U41366 (N_41366,N_39987,N_39429);
and U41367 (N_41367,N_38554,N_39440);
nand U41368 (N_41368,N_38772,N_39808);
and U41369 (N_41369,N_39460,N_38654);
nor U41370 (N_41370,N_38008,N_39056);
nand U41371 (N_41371,N_38840,N_39812);
nor U41372 (N_41372,N_38331,N_38232);
or U41373 (N_41373,N_39844,N_38505);
nor U41374 (N_41374,N_38975,N_39066);
xnor U41375 (N_41375,N_39952,N_38375);
nand U41376 (N_41376,N_38910,N_38948);
and U41377 (N_41377,N_38489,N_39628);
and U41378 (N_41378,N_38644,N_39546);
or U41379 (N_41379,N_39898,N_38147);
or U41380 (N_41380,N_39591,N_39423);
xor U41381 (N_41381,N_39563,N_38435);
or U41382 (N_41382,N_38639,N_39028);
and U41383 (N_41383,N_39439,N_38791);
xor U41384 (N_41384,N_38847,N_38211);
xor U41385 (N_41385,N_38763,N_38861);
nor U41386 (N_41386,N_39130,N_39306);
and U41387 (N_41387,N_38636,N_39428);
nand U41388 (N_41388,N_39641,N_39719);
nor U41389 (N_41389,N_38906,N_38211);
nand U41390 (N_41390,N_39246,N_39649);
and U41391 (N_41391,N_38681,N_38920);
xor U41392 (N_41392,N_38425,N_39545);
nand U41393 (N_41393,N_38587,N_38736);
xnor U41394 (N_41394,N_39221,N_39536);
xor U41395 (N_41395,N_39066,N_38671);
nor U41396 (N_41396,N_38876,N_39856);
xor U41397 (N_41397,N_39039,N_38434);
nor U41398 (N_41398,N_38063,N_39899);
xnor U41399 (N_41399,N_38324,N_39879);
xnor U41400 (N_41400,N_38285,N_39393);
xnor U41401 (N_41401,N_38133,N_38497);
nor U41402 (N_41402,N_39685,N_38745);
nor U41403 (N_41403,N_38693,N_38518);
xor U41404 (N_41404,N_38886,N_39539);
nand U41405 (N_41405,N_38045,N_38905);
nand U41406 (N_41406,N_38075,N_39223);
or U41407 (N_41407,N_38997,N_38211);
and U41408 (N_41408,N_39667,N_39295);
nor U41409 (N_41409,N_39773,N_38589);
or U41410 (N_41410,N_38936,N_39668);
or U41411 (N_41411,N_38324,N_39951);
nand U41412 (N_41412,N_38099,N_39317);
or U41413 (N_41413,N_39526,N_38517);
xor U41414 (N_41414,N_38544,N_38555);
or U41415 (N_41415,N_39065,N_39808);
nor U41416 (N_41416,N_39006,N_38405);
nor U41417 (N_41417,N_38861,N_38490);
nand U41418 (N_41418,N_39021,N_38560);
or U41419 (N_41419,N_39340,N_38367);
and U41420 (N_41420,N_39530,N_39988);
and U41421 (N_41421,N_38410,N_39114);
and U41422 (N_41422,N_39469,N_38187);
and U41423 (N_41423,N_38878,N_38000);
nand U41424 (N_41424,N_38045,N_39142);
nor U41425 (N_41425,N_39058,N_39414);
xor U41426 (N_41426,N_38563,N_39644);
or U41427 (N_41427,N_38424,N_38329);
xnor U41428 (N_41428,N_38055,N_39422);
nand U41429 (N_41429,N_39545,N_39865);
or U41430 (N_41430,N_39165,N_39212);
nor U41431 (N_41431,N_39062,N_39473);
nand U41432 (N_41432,N_38094,N_38750);
nor U41433 (N_41433,N_38686,N_39972);
xnor U41434 (N_41434,N_39696,N_38675);
and U41435 (N_41435,N_38667,N_38894);
xor U41436 (N_41436,N_38624,N_38584);
or U41437 (N_41437,N_39185,N_38920);
nand U41438 (N_41438,N_39482,N_39914);
and U41439 (N_41439,N_38709,N_39042);
nor U41440 (N_41440,N_38310,N_38294);
and U41441 (N_41441,N_38006,N_38421);
nor U41442 (N_41442,N_39547,N_38350);
xor U41443 (N_41443,N_38337,N_38324);
nand U41444 (N_41444,N_39671,N_38785);
nor U41445 (N_41445,N_39384,N_38836);
or U41446 (N_41446,N_38571,N_39296);
or U41447 (N_41447,N_39934,N_39115);
and U41448 (N_41448,N_38162,N_39770);
xor U41449 (N_41449,N_39618,N_38571);
or U41450 (N_41450,N_39611,N_38348);
or U41451 (N_41451,N_38932,N_39127);
or U41452 (N_41452,N_38271,N_38602);
and U41453 (N_41453,N_38816,N_39472);
xor U41454 (N_41454,N_38859,N_38989);
and U41455 (N_41455,N_39041,N_39124);
or U41456 (N_41456,N_38638,N_39344);
nand U41457 (N_41457,N_38833,N_39424);
nor U41458 (N_41458,N_39599,N_39659);
nor U41459 (N_41459,N_38513,N_39918);
and U41460 (N_41460,N_38529,N_39308);
or U41461 (N_41461,N_39274,N_38837);
nand U41462 (N_41462,N_39590,N_39519);
nor U41463 (N_41463,N_39681,N_38972);
and U41464 (N_41464,N_38899,N_38531);
and U41465 (N_41465,N_38052,N_39042);
nand U41466 (N_41466,N_39333,N_38020);
and U41467 (N_41467,N_38854,N_39321);
nand U41468 (N_41468,N_39334,N_39804);
nand U41469 (N_41469,N_38063,N_39385);
or U41470 (N_41470,N_39350,N_38638);
nor U41471 (N_41471,N_38575,N_38782);
xnor U41472 (N_41472,N_39406,N_39134);
and U41473 (N_41473,N_38042,N_38272);
nor U41474 (N_41474,N_38525,N_39205);
and U41475 (N_41475,N_38976,N_39821);
nand U41476 (N_41476,N_39948,N_38497);
nor U41477 (N_41477,N_38960,N_39280);
nand U41478 (N_41478,N_38270,N_38372);
nor U41479 (N_41479,N_39229,N_39264);
nor U41480 (N_41480,N_38172,N_39595);
xor U41481 (N_41481,N_38020,N_39234);
or U41482 (N_41482,N_39102,N_39104);
or U41483 (N_41483,N_38035,N_39297);
xor U41484 (N_41484,N_38947,N_39523);
nor U41485 (N_41485,N_39707,N_38540);
xnor U41486 (N_41486,N_39793,N_38474);
or U41487 (N_41487,N_38602,N_38514);
and U41488 (N_41488,N_38308,N_38508);
and U41489 (N_41489,N_39238,N_38400);
and U41490 (N_41490,N_39938,N_39287);
xnor U41491 (N_41491,N_39608,N_38446);
and U41492 (N_41492,N_39385,N_39683);
or U41493 (N_41493,N_38955,N_38477);
and U41494 (N_41494,N_38032,N_39558);
nand U41495 (N_41495,N_39319,N_39615);
nor U41496 (N_41496,N_39734,N_39241);
nor U41497 (N_41497,N_38321,N_38172);
or U41498 (N_41498,N_38421,N_39612);
nor U41499 (N_41499,N_39026,N_39288);
nand U41500 (N_41500,N_38044,N_38173);
xor U41501 (N_41501,N_38041,N_39823);
nand U41502 (N_41502,N_39743,N_39008);
or U41503 (N_41503,N_39745,N_39626);
and U41504 (N_41504,N_38445,N_38576);
xor U41505 (N_41505,N_38518,N_39043);
nand U41506 (N_41506,N_39539,N_38601);
xnor U41507 (N_41507,N_39996,N_38129);
or U41508 (N_41508,N_38302,N_38212);
and U41509 (N_41509,N_38517,N_39321);
nor U41510 (N_41510,N_39150,N_38283);
or U41511 (N_41511,N_38670,N_39256);
or U41512 (N_41512,N_39763,N_39417);
or U41513 (N_41513,N_39588,N_39335);
nand U41514 (N_41514,N_39584,N_38062);
nor U41515 (N_41515,N_38519,N_38049);
nor U41516 (N_41516,N_38629,N_38235);
nor U41517 (N_41517,N_39390,N_38992);
nor U41518 (N_41518,N_39274,N_39559);
xor U41519 (N_41519,N_39499,N_39444);
or U41520 (N_41520,N_39226,N_38329);
or U41521 (N_41521,N_39651,N_38624);
xor U41522 (N_41522,N_39482,N_38453);
nor U41523 (N_41523,N_38737,N_38408);
or U41524 (N_41524,N_38519,N_39506);
or U41525 (N_41525,N_39961,N_39393);
nor U41526 (N_41526,N_38947,N_39629);
or U41527 (N_41527,N_38750,N_38242);
xor U41528 (N_41528,N_39632,N_38881);
and U41529 (N_41529,N_39839,N_38248);
nor U41530 (N_41530,N_38532,N_39053);
nor U41531 (N_41531,N_39515,N_39030);
or U41532 (N_41532,N_39347,N_39979);
xnor U41533 (N_41533,N_39917,N_39548);
xor U41534 (N_41534,N_39000,N_39703);
nand U41535 (N_41535,N_38451,N_39154);
nand U41536 (N_41536,N_39770,N_38777);
xnor U41537 (N_41537,N_39047,N_38891);
or U41538 (N_41538,N_38020,N_38643);
nor U41539 (N_41539,N_38939,N_39681);
nor U41540 (N_41540,N_39643,N_39016);
or U41541 (N_41541,N_38633,N_38256);
nand U41542 (N_41542,N_38189,N_38446);
xnor U41543 (N_41543,N_39630,N_38003);
xor U41544 (N_41544,N_38010,N_38004);
nor U41545 (N_41545,N_39175,N_38160);
nand U41546 (N_41546,N_39810,N_39553);
and U41547 (N_41547,N_39753,N_39437);
and U41548 (N_41548,N_38027,N_39623);
and U41549 (N_41549,N_38720,N_38000);
or U41550 (N_41550,N_38126,N_38355);
nand U41551 (N_41551,N_39613,N_38214);
or U41552 (N_41552,N_39376,N_39543);
and U41553 (N_41553,N_39901,N_39903);
and U41554 (N_41554,N_38243,N_38087);
nor U41555 (N_41555,N_39642,N_38383);
nand U41556 (N_41556,N_39477,N_39841);
and U41557 (N_41557,N_39118,N_39792);
nand U41558 (N_41558,N_38256,N_39862);
nor U41559 (N_41559,N_39951,N_39492);
xor U41560 (N_41560,N_38203,N_38916);
nand U41561 (N_41561,N_39601,N_39711);
and U41562 (N_41562,N_39134,N_38288);
nor U41563 (N_41563,N_38126,N_39728);
nor U41564 (N_41564,N_38138,N_38214);
nand U41565 (N_41565,N_38938,N_38424);
and U41566 (N_41566,N_39565,N_39183);
and U41567 (N_41567,N_38123,N_39011);
or U41568 (N_41568,N_38530,N_38842);
or U41569 (N_41569,N_38469,N_38993);
and U41570 (N_41570,N_38638,N_38415);
and U41571 (N_41571,N_39473,N_38491);
and U41572 (N_41572,N_39332,N_38514);
nand U41573 (N_41573,N_38133,N_38143);
xor U41574 (N_41574,N_38903,N_39282);
xnor U41575 (N_41575,N_38032,N_39944);
xor U41576 (N_41576,N_39771,N_38942);
nand U41577 (N_41577,N_38978,N_39689);
and U41578 (N_41578,N_38031,N_39727);
and U41579 (N_41579,N_39187,N_38781);
xor U41580 (N_41580,N_39255,N_38141);
nor U41581 (N_41581,N_39882,N_38457);
xor U41582 (N_41582,N_39973,N_38311);
and U41583 (N_41583,N_38559,N_39623);
or U41584 (N_41584,N_39438,N_38131);
xnor U41585 (N_41585,N_39305,N_38383);
or U41586 (N_41586,N_38065,N_39187);
and U41587 (N_41587,N_39635,N_39095);
xor U41588 (N_41588,N_38098,N_39706);
or U41589 (N_41589,N_39861,N_38883);
xnor U41590 (N_41590,N_39117,N_39331);
and U41591 (N_41591,N_39278,N_39632);
nor U41592 (N_41592,N_38789,N_38754);
or U41593 (N_41593,N_38095,N_39520);
or U41594 (N_41594,N_38730,N_39191);
and U41595 (N_41595,N_39878,N_38228);
nor U41596 (N_41596,N_39253,N_39545);
nor U41597 (N_41597,N_38630,N_39368);
xor U41598 (N_41598,N_39304,N_39440);
nand U41599 (N_41599,N_39890,N_38205);
nor U41600 (N_41600,N_38521,N_38435);
nor U41601 (N_41601,N_39816,N_38917);
xnor U41602 (N_41602,N_38871,N_39056);
nor U41603 (N_41603,N_39930,N_38903);
xnor U41604 (N_41604,N_39476,N_38734);
xor U41605 (N_41605,N_38384,N_38196);
nand U41606 (N_41606,N_38621,N_38731);
nand U41607 (N_41607,N_39339,N_38149);
and U41608 (N_41608,N_38208,N_38938);
and U41609 (N_41609,N_39661,N_39610);
xnor U41610 (N_41610,N_39491,N_38155);
nor U41611 (N_41611,N_38346,N_38863);
xor U41612 (N_41612,N_38018,N_39022);
nor U41613 (N_41613,N_38050,N_39195);
xnor U41614 (N_41614,N_38013,N_39405);
xnor U41615 (N_41615,N_38634,N_39800);
nor U41616 (N_41616,N_38958,N_39538);
xnor U41617 (N_41617,N_39830,N_39208);
and U41618 (N_41618,N_38933,N_39013);
nand U41619 (N_41619,N_38170,N_38786);
nand U41620 (N_41620,N_38951,N_38607);
and U41621 (N_41621,N_38888,N_39946);
or U41622 (N_41622,N_38646,N_38250);
and U41623 (N_41623,N_39864,N_38755);
and U41624 (N_41624,N_38133,N_39685);
nor U41625 (N_41625,N_38644,N_39353);
nor U41626 (N_41626,N_38496,N_38220);
nand U41627 (N_41627,N_38790,N_39972);
or U41628 (N_41628,N_38121,N_38735);
nand U41629 (N_41629,N_39084,N_39641);
and U41630 (N_41630,N_39709,N_38697);
nand U41631 (N_41631,N_39221,N_39238);
xor U41632 (N_41632,N_39888,N_38057);
nand U41633 (N_41633,N_39170,N_39949);
and U41634 (N_41634,N_38238,N_39499);
and U41635 (N_41635,N_39813,N_38441);
nand U41636 (N_41636,N_38128,N_38252);
and U41637 (N_41637,N_38200,N_38364);
xor U41638 (N_41638,N_38721,N_38694);
nor U41639 (N_41639,N_38488,N_38998);
or U41640 (N_41640,N_38966,N_39083);
xor U41641 (N_41641,N_39463,N_38083);
nand U41642 (N_41642,N_38539,N_39452);
nand U41643 (N_41643,N_39126,N_38866);
nor U41644 (N_41644,N_38896,N_39250);
xnor U41645 (N_41645,N_38038,N_39150);
xor U41646 (N_41646,N_38448,N_38128);
or U41647 (N_41647,N_39880,N_39416);
or U41648 (N_41648,N_39877,N_39967);
xor U41649 (N_41649,N_38799,N_39729);
or U41650 (N_41650,N_39345,N_38268);
and U41651 (N_41651,N_38772,N_39106);
nor U41652 (N_41652,N_39875,N_39145);
nor U41653 (N_41653,N_38485,N_39234);
xnor U41654 (N_41654,N_38319,N_39187);
xnor U41655 (N_41655,N_38687,N_38012);
nand U41656 (N_41656,N_39969,N_38823);
nor U41657 (N_41657,N_38494,N_39148);
xor U41658 (N_41658,N_39426,N_39747);
nor U41659 (N_41659,N_39472,N_39758);
or U41660 (N_41660,N_38724,N_39060);
nor U41661 (N_41661,N_38265,N_38750);
nand U41662 (N_41662,N_39014,N_39344);
or U41663 (N_41663,N_38746,N_39373);
or U41664 (N_41664,N_38681,N_38555);
or U41665 (N_41665,N_38763,N_39229);
and U41666 (N_41666,N_38812,N_39628);
and U41667 (N_41667,N_39354,N_39229);
nor U41668 (N_41668,N_39339,N_38362);
xor U41669 (N_41669,N_38559,N_38850);
nand U41670 (N_41670,N_38422,N_38110);
xnor U41671 (N_41671,N_39853,N_38250);
and U41672 (N_41672,N_38029,N_38154);
nand U41673 (N_41673,N_38462,N_38147);
and U41674 (N_41674,N_38675,N_38706);
or U41675 (N_41675,N_38835,N_39381);
nor U41676 (N_41676,N_38192,N_38852);
and U41677 (N_41677,N_39283,N_38007);
nand U41678 (N_41678,N_39994,N_39159);
and U41679 (N_41679,N_39191,N_38532);
and U41680 (N_41680,N_39762,N_38823);
xnor U41681 (N_41681,N_39442,N_38619);
nand U41682 (N_41682,N_38370,N_39954);
and U41683 (N_41683,N_38422,N_38977);
or U41684 (N_41684,N_38305,N_39824);
nor U41685 (N_41685,N_39595,N_38447);
or U41686 (N_41686,N_39909,N_39260);
or U41687 (N_41687,N_39318,N_39276);
and U41688 (N_41688,N_39587,N_38307);
or U41689 (N_41689,N_39069,N_38346);
nand U41690 (N_41690,N_39153,N_38487);
or U41691 (N_41691,N_39755,N_38503);
or U41692 (N_41692,N_39233,N_38089);
or U41693 (N_41693,N_38531,N_38333);
nor U41694 (N_41694,N_38869,N_39715);
nor U41695 (N_41695,N_38870,N_39947);
nor U41696 (N_41696,N_39116,N_39132);
xnor U41697 (N_41697,N_39494,N_39738);
nand U41698 (N_41698,N_38047,N_38656);
and U41699 (N_41699,N_38168,N_38006);
nor U41700 (N_41700,N_38418,N_39013);
or U41701 (N_41701,N_39889,N_39906);
nor U41702 (N_41702,N_38712,N_38893);
nor U41703 (N_41703,N_38472,N_38159);
xor U41704 (N_41704,N_38784,N_39965);
nor U41705 (N_41705,N_38603,N_38487);
and U41706 (N_41706,N_38655,N_39668);
xnor U41707 (N_41707,N_39502,N_38702);
and U41708 (N_41708,N_38589,N_38658);
xor U41709 (N_41709,N_39076,N_39260);
nand U41710 (N_41710,N_38483,N_38071);
or U41711 (N_41711,N_38414,N_38339);
xnor U41712 (N_41712,N_38754,N_39066);
nor U41713 (N_41713,N_38121,N_39820);
nor U41714 (N_41714,N_39512,N_39484);
nor U41715 (N_41715,N_39479,N_38134);
and U41716 (N_41716,N_39364,N_38480);
xnor U41717 (N_41717,N_39566,N_38019);
xor U41718 (N_41718,N_39309,N_39576);
and U41719 (N_41719,N_39671,N_38880);
nand U41720 (N_41720,N_38957,N_38240);
or U41721 (N_41721,N_38758,N_39942);
and U41722 (N_41722,N_38710,N_39389);
nor U41723 (N_41723,N_39761,N_39594);
nor U41724 (N_41724,N_39510,N_39783);
and U41725 (N_41725,N_38351,N_38480);
nor U41726 (N_41726,N_38719,N_38888);
and U41727 (N_41727,N_39299,N_39029);
nor U41728 (N_41728,N_39783,N_39009);
nor U41729 (N_41729,N_39176,N_39333);
or U41730 (N_41730,N_39461,N_39091);
and U41731 (N_41731,N_38603,N_39512);
and U41732 (N_41732,N_39802,N_38000);
nor U41733 (N_41733,N_38251,N_38232);
nor U41734 (N_41734,N_39670,N_39649);
nand U41735 (N_41735,N_39699,N_38907);
nand U41736 (N_41736,N_38266,N_38913);
and U41737 (N_41737,N_39396,N_39457);
or U41738 (N_41738,N_39289,N_38580);
and U41739 (N_41739,N_39893,N_39486);
or U41740 (N_41740,N_39248,N_39659);
xnor U41741 (N_41741,N_39457,N_39077);
xnor U41742 (N_41742,N_39014,N_39613);
or U41743 (N_41743,N_38328,N_38652);
xnor U41744 (N_41744,N_39368,N_38884);
and U41745 (N_41745,N_39061,N_39499);
xor U41746 (N_41746,N_39764,N_38763);
xor U41747 (N_41747,N_39385,N_38881);
nor U41748 (N_41748,N_39140,N_38216);
and U41749 (N_41749,N_39943,N_39581);
or U41750 (N_41750,N_39750,N_39211);
nor U41751 (N_41751,N_38163,N_39438);
nand U41752 (N_41752,N_38183,N_38355);
nand U41753 (N_41753,N_38692,N_39364);
xnor U41754 (N_41754,N_38136,N_38164);
xor U41755 (N_41755,N_39547,N_39373);
or U41756 (N_41756,N_39420,N_38204);
nand U41757 (N_41757,N_39430,N_39733);
nor U41758 (N_41758,N_38353,N_39918);
xnor U41759 (N_41759,N_38294,N_39162);
or U41760 (N_41760,N_39684,N_39867);
xor U41761 (N_41761,N_38687,N_38589);
nand U41762 (N_41762,N_39788,N_39294);
and U41763 (N_41763,N_38436,N_38775);
xnor U41764 (N_41764,N_39173,N_38351);
xnor U41765 (N_41765,N_39781,N_39822);
or U41766 (N_41766,N_38003,N_38063);
nor U41767 (N_41767,N_39480,N_39444);
xnor U41768 (N_41768,N_39543,N_38659);
nor U41769 (N_41769,N_39500,N_38037);
nand U41770 (N_41770,N_38617,N_38940);
and U41771 (N_41771,N_39151,N_39032);
or U41772 (N_41772,N_39604,N_38052);
xor U41773 (N_41773,N_38013,N_38089);
or U41774 (N_41774,N_38547,N_38502);
nor U41775 (N_41775,N_38024,N_38974);
or U41776 (N_41776,N_39868,N_38616);
xor U41777 (N_41777,N_38793,N_39458);
and U41778 (N_41778,N_38608,N_38461);
nand U41779 (N_41779,N_38675,N_38561);
xor U41780 (N_41780,N_38688,N_39580);
nor U41781 (N_41781,N_38484,N_39975);
nor U41782 (N_41782,N_38053,N_39446);
nand U41783 (N_41783,N_39949,N_38272);
and U41784 (N_41784,N_38473,N_39213);
nand U41785 (N_41785,N_38006,N_38468);
nor U41786 (N_41786,N_39052,N_39768);
nor U41787 (N_41787,N_39299,N_39104);
xor U41788 (N_41788,N_38843,N_38069);
xor U41789 (N_41789,N_38164,N_39342);
nand U41790 (N_41790,N_39128,N_39359);
xor U41791 (N_41791,N_39050,N_38022);
xor U41792 (N_41792,N_38207,N_38310);
xor U41793 (N_41793,N_39209,N_38809);
or U41794 (N_41794,N_38026,N_38472);
nor U41795 (N_41795,N_38757,N_38683);
nand U41796 (N_41796,N_38406,N_38488);
nand U41797 (N_41797,N_38685,N_39535);
and U41798 (N_41798,N_38695,N_38774);
nand U41799 (N_41799,N_39646,N_39887);
nand U41800 (N_41800,N_39131,N_38539);
nor U41801 (N_41801,N_38357,N_38166);
xnor U41802 (N_41802,N_39099,N_38703);
xor U41803 (N_41803,N_39495,N_38791);
nor U41804 (N_41804,N_39719,N_39595);
and U41805 (N_41805,N_38654,N_38650);
and U41806 (N_41806,N_38673,N_38551);
xnor U41807 (N_41807,N_38057,N_39249);
xor U41808 (N_41808,N_38659,N_39935);
nor U41809 (N_41809,N_39921,N_38617);
or U41810 (N_41810,N_38217,N_39472);
nand U41811 (N_41811,N_39385,N_39248);
xor U41812 (N_41812,N_38999,N_38033);
xnor U41813 (N_41813,N_38950,N_38599);
nor U41814 (N_41814,N_39442,N_38079);
xnor U41815 (N_41815,N_38453,N_38488);
or U41816 (N_41816,N_38813,N_39170);
nor U41817 (N_41817,N_39585,N_39922);
or U41818 (N_41818,N_39437,N_38527);
xnor U41819 (N_41819,N_39920,N_38117);
or U41820 (N_41820,N_39865,N_39754);
or U41821 (N_41821,N_38723,N_38597);
xor U41822 (N_41822,N_39540,N_38500);
nor U41823 (N_41823,N_38416,N_38235);
or U41824 (N_41824,N_39537,N_38110);
nor U41825 (N_41825,N_38771,N_38300);
nor U41826 (N_41826,N_39418,N_38119);
and U41827 (N_41827,N_38445,N_38899);
or U41828 (N_41828,N_39572,N_38572);
xor U41829 (N_41829,N_39845,N_38886);
nor U41830 (N_41830,N_39622,N_39989);
nand U41831 (N_41831,N_38557,N_39592);
nor U41832 (N_41832,N_39511,N_39573);
or U41833 (N_41833,N_39371,N_39825);
nand U41834 (N_41834,N_38547,N_38232);
nor U41835 (N_41835,N_39576,N_38375);
or U41836 (N_41836,N_39255,N_39570);
or U41837 (N_41837,N_39434,N_38975);
nand U41838 (N_41838,N_39936,N_39630);
or U41839 (N_41839,N_39754,N_39473);
or U41840 (N_41840,N_38824,N_38391);
nand U41841 (N_41841,N_39297,N_38352);
or U41842 (N_41842,N_38117,N_38354);
and U41843 (N_41843,N_39540,N_39210);
nand U41844 (N_41844,N_38361,N_39722);
xnor U41845 (N_41845,N_39457,N_39035);
nand U41846 (N_41846,N_39297,N_39723);
and U41847 (N_41847,N_38608,N_38394);
or U41848 (N_41848,N_38767,N_38251);
or U41849 (N_41849,N_38446,N_39008);
xor U41850 (N_41850,N_38879,N_39668);
or U41851 (N_41851,N_39728,N_39348);
nand U41852 (N_41852,N_38241,N_39890);
or U41853 (N_41853,N_39840,N_39715);
nand U41854 (N_41854,N_38603,N_38277);
xor U41855 (N_41855,N_38785,N_39996);
and U41856 (N_41856,N_39562,N_39294);
xor U41857 (N_41857,N_38680,N_39921);
or U41858 (N_41858,N_38174,N_39952);
and U41859 (N_41859,N_38662,N_38968);
xnor U41860 (N_41860,N_38528,N_38375);
nand U41861 (N_41861,N_38880,N_38770);
and U41862 (N_41862,N_38505,N_38056);
or U41863 (N_41863,N_38098,N_38958);
xnor U41864 (N_41864,N_38204,N_39372);
xnor U41865 (N_41865,N_38314,N_38172);
xor U41866 (N_41866,N_39634,N_38952);
nor U41867 (N_41867,N_39700,N_39197);
nand U41868 (N_41868,N_39002,N_38795);
and U41869 (N_41869,N_39518,N_39167);
and U41870 (N_41870,N_39510,N_38590);
and U41871 (N_41871,N_39596,N_38726);
or U41872 (N_41872,N_39032,N_38134);
xnor U41873 (N_41873,N_38984,N_38890);
xnor U41874 (N_41874,N_38146,N_38762);
xnor U41875 (N_41875,N_38522,N_39321);
nor U41876 (N_41876,N_38758,N_38990);
xnor U41877 (N_41877,N_39711,N_38313);
or U41878 (N_41878,N_38475,N_38343);
nand U41879 (N_41879,N_38113,N_39426);
xor U41880 (N_41880,N_39979,N_38782);
xnor U41881 (N_41881,N_38662,N_38522);
and U41882 (N_41882,N_39892,N_38426);
nor U41883 (N_41883,N_38418,N_39751);
nor U41884 (N_41884,N_38836,N_38625);
xnor U41885 (N_41885,N_38168,N_39191);
nand U41886 (N_41886,N_38820,N_39341);
and U41887 (N_41887,N_38457,N_39239);
or U41888 (N_41888,N_39348,N_38755);
and U41889 (N_41889,N_38904,N_39709);
and U41890 (N_41890,N_39842,N_39612);
nor U41891 (N_41891,N_38968,N_38677);
and U41892 (N_41892,N_38720,N_38347);
or U41893 (N_41893,N_39716,N_39788);
nand U41894 (N_41894,N_38873,N_39925);
nor U41895 (N_41895,N_38258,N_38444);
xor U41896 (N_41896,N_38300,N_39282);
nand U41897 (N_41897,N_38204,N_38326);
and U41898 (N_41898,N_38459,N_39594);
nor U41899 (N_41899,N_39089,N_39486);
and U41900 (N_41900,N_39435,N_39279);
nand U41901 (N_41901,N_38827,N_38287);
and U41902 (N_41902,N_38782,N_39228);
xnor U41903 (N_41903,N_38470,N_39747);
xor U41904 (N_41904,N_38431,N_38808);
or U41905 (N_41905,N_38158,N_38288);
nor U41906 (N_41906,N_39725,N_38350);
nor U41907 (N_41907,N_38000,N_38437);
nor U41908 (N_41908,N_38463,N_38368);
or U41909 (N_41909,N_38088,N_38103);
and U41910 (N_41910,N_39053,N_38819);
and U41911 (N_41911,N_38641,N_38317);
nand U41912 (N_41912,N_39569,N_38171);
nand U41913 (N_41913,N_39000,N_38539);
nand U41914 (N_41914,N_39076,N_39645);
and U41915 (N_41915,N_38987,N_38353);
and U41916 (N_41916,N_38724,N_39655);
or U41917 (N_41917,N_39592,N_38706);
and U41918 (N_41918,N_38334,N_39341);
nand U41919 (N_41919,N_39681,N_39981);
xor U41920 (N_41920,N_38757,N_38220);
xor U41921 (N_41921,N_38191,N_38753);
or U41922 (N_41922,N_38830,N_39312);
nor U41923 (N_41923,N_39419,N_38691);
nor U41924 (N_41924,N_39579,N_39105);
xor U41925 (N_41925,N_38152,N_39434);
and U41926 (N_41926,N_39342,N_38562);
or U41927 (N_41927,N_38798,N_39498);
and U41928 (N_41928,N_38257,N_38907);
nand U41929 (N_41929,N_38005,N_38885);
or U41930 (N_41930,N_39534,N_39586);
nand U41931 (N_41931,N_39347,N_39864);
nor U41932 (N_41932,N_38740,N_39258);
or U41933 (N_41933,N_39710,N_39304);
nor U41934 (N_41934,N_39311,N_39915);
and U41935 (N_41935,N_39399,N_39723);
nor U41936 (N_41936,N_39034,N_38655);
nand U41937 (N_41937,N_38655,N_39176);
nand U41938 (N_41938,N_38913,N_39947);
xnor U41939 (N_41939,N_39055,N_38047);
nand U41940 (N_41940,N_38812,N_38382);
xor U41941 (N_41941,N_38259,N_38640);
nand U41942 (N_41942,N_38135,N_39482);
and U41943 (N_41943,N_38328,N_39128);
nand U41944 (N_41944,N_38869,N_38883);
nor U41945 (N_41945,N_38021,N_39160);
nand U41946 (N_41946,N_39623,N_39668);
or U41947 (N_41947,N_38527,N_39297);
xnor U41948 (N_41948,N_39360,N_38056);
nand U41949 (N_41949,N_39919,N_39370);
or U41950 (N_41950,N_39818,N_39839);
xor U41951 (N_41951,N_39252,N_38888);
and U41952 (N_41952,N_39568,N_38098);
and U41953 (N_41953,N_38771,N_39499);
xnor U41954 (N_41954,N_39422,N_38456);
nand U41955 (N_41955,N_39639,N_38172);
and U41956 (N_41956,N_38533,N_38518);
or U41957 (N_41957,N_38160,N_38078);
nor U41958 (N_41958,N_38019,N_39129);
xnor U41959 (N_41959,N_39347,N_38403);
nand U41960 (N_41960,N_38687,N_38948);
nand U41961 (N_41961,N_38860,N_39705);
nand U41962 (N_41962,N_38466,N_39801);
nor U41963 (N_41963,N_38183,N_38086);
nor U41964 (N_41964,N_39359,N_38300);
nor U41965 (N_41965,N_38561,N_38625);
nand U41966 (N_41966,N_38147,N_38326);
or U41967 (N_41967,N_38040,N_38796);
and U41968 (N_41968,N_38639,N_39577);
nand U41969 (N_41969,N_38492,N_39843);
xnor U41970 (N_41970,N_38625,N_39145);
nor U41971 (N_41971,N_39771,N_38654);
nor U41972 (N_41972,N_39344,N_38125);
or U41973 (N_41973,N_39461,N_38043);
and U41974 (N_41974,N_38791,N_38000);
nand U41975 (N_41975,N_39983,N_39312);
or U41976 (N_41976,N_38772,N_39195);
and U41977 (N_41977,N_39578,N_39832);
and U41978 (N_41978,N_38200,N_39433);
xnor U41979 (N_41979,N_38574,N_39274);
or U41980 (N_41980,N_39013,N_38468);
xnor U41981 (N_41981,N_39998,N_38231);
nor U41982 (N_41982,N_38765,N_39552);
or U41983 (N_41983,N_39163,N_38648);
nor U41984 (N_41984,N_38986,N_39975);
nand U41985 (N_41985,N_39819,N_38368);
and U41986 (N_41986,N_38338,N_39494);
and U41987 (N_41987,N_38541,N_38174);
xor U41988 (N_41988,N_38463,N_39604);
nand U41989 (N_41989,N_38913,N_38641);
xnor U41990 (N_41990,N_38894,N_38765);
and U41991 (N_41991,N_38809,N_38931);
nand U41992 (N_41992,N_39102,N_39542);
nor U41993 (N_41993,N_38248,N_38960);
xnor U41994 (N_41994,N_39441,N_38504);
nand U41995 (N_41995,N_39908,N_38037);
nand U41996 (N_41996,N_39619,N_39072);
nor U41997 (N_41997,N_38597,N_39785);
or U41998 (N_41998,N_39191,N_39641);
nor U41999 (N_41999,N_38829,N_39382);
xor U42000 (N_42000,N_41069,N_40950);
and U42001 (N_42001,N_41167,N_41921);
or U42002 (N_42002,N_40425,N_41857);
nor U42003 (N_42003,N_41257,N_40590);
nand U42004 (N_42004,N_41404,N_40356);
xor U42005 (N_42005,N_40757,N_41516);
and U42006 (N_42006,N_40948,N_40061);
or U42007 (N_42007,N_40611,N_41077);
nand U42008 (N_42008,N_41452,N_41053);
or U42009 (N_42009,N_41523,N_40522);
and U42010 (N_42010,N_41218,N_40753);
nor U42011 (N_42011,N_40949,N_41133);
nand U42012 (N_42012,N_40612,N_41242);
xnor U42013 (N_42013,N_40306,N_41393);
or U42014 (N_42014,N_41935,N_40199);
xor U42015 (N_42015,N_41056,N_41586);
xnor U42016 (N_42016,N_41677,N_40070);
and U42017 (N_42017,N_40558,N_40194);
and U42018 (N_42018,N_41325,N_40797);
and U42019 (N_42019,N_41214,N_40803);
nand U42020 (N_42020,N_41634,N_40768);
or U42021 (N_42021,N_41927,N_40835);
and U42022 (N_42022,N_41878,N_41776);
xor U42023 (N_42023,N_40890,N_41459);
nor U42024 (N_42024,N_40637,N_40386);
and U42025 (N_42025,N_41993,N_40037);
and U42026 (N_42026,N_41071,N_40318);
and U42027 (N_42027,N_40747,N_40717);
nor U42028 (N_42028,N_41276,N_41864);
nand U42029 (N_42029,N_41912,N_40490);
or U42030 (N_42030,N_40456,N_40363);
nand U42031 (N_42031,N_41846,N_40682);
xor U42032 (N_42032,N_40785,N_40352);
nand U42033 (N_42033,N_41684,N_41746);
or U42034 (N_42034,N_40654,N_41751);
xor U42035 (N_42035,N_41322,N_41389);
or U42036 (N_42036,N_41345,N_41201);
xor U42037 (N_42037,N_41984,N_41615);
nand U42038 (N_42038,N_41052,N_41565);
and U42039 (N_42039,N_40715,N_41964);
nor U42040 (N_42040,N_41161,N_41850);
nor U42041 (N_42041,N_40414,N_40703);
nor U42042 (N_42042,N_40938,N_41600);
xnor U42043 (N_42043,N_40610,N_40931);
or U42044 (N_42044,N_41807,N_40775);
nor U42045 (N_42045,N_40173,N_41683);
nand U42046 (N_42046,N_40354,N_40680);
xor U42047 (N_42047,N_40521,N_41844);
or U42048 (N_42048,N_41206,N_41624);
nor U42049 (N_42049,N_40200,N_40546);
and U42050 (N_42050,N_40706,N_40377);
xor U42051 (N_42051,N_41465,N_41224);
or U42052 (N_42052,N_41032,N_41008);
or U42053 (N_42053,N_40591,N_40259);
or U42054 (N_42054,N_40211,N_41955);
nor U42055 (N_42055,N_40164,N_40373);
or U42056 (N_42056,N_41756,N_41068);
xnor U42057 (N_42057,N_41670,N_40067);
nor U42058 (N_42058,N_40023,N_40412);
xnor U42059 (N_42059,N_40174,N_40622);
and U42060 (N_42060,N_40537,N_40817);
or U42061 (N_42061,N_40805,N_41779);
nand U42062 (N_42062,N_41996,N_41190);
xor U42063 (N_42063,N_41660,N_41637);
nor U42064 (N_42064,N_41287,N_41527);
xnor U42065 (N_42065,N_40069,N_41035);
or U42066 (N_42066,N_40481,N_40374);
and U42067 (N_42067,N_41438,N_41079);
nor U42068 (N_42068,N_40427,N_40663);
or U42069 (N_42069,N_41832,N_40629);
nor U42070 (N_42070,N_41617,N_41140);
and U42071 (N_42071,N_41488,N_41903);
xnor U42072 (N_42072,N_41687,N_41557);
and U42073 (N_42073,N_41040,N_41361);
nand U42074 (N_42074,N_40660,N_40782);
nand U42075 (N_42075,N_40662,N_40336);
nor U42076 (N_42076,N_40976,N_41753);
nor U42077 (N_42077,N_40979,N_41093);
nand U42078 (N_42078,N_41948,N_40764);
xnor U42079 (N_42079,N_41471,N_40201);
nor U42080 (N_42080,N_41428,N_40968);
nand U42081 (N_42081,N_40900,N_40721);
and U42082 (N_42082,N_40407,N_41820);
or U42083 (N_42083,N_41936,N_41399);
nor U42084 (N_42084,N_41142,N_41463);
nor U42085 (N_42085,N_41232,N_41095);
nor U42086 (N_42086,N_40655,N_41942);
or U42087 (N_42087,N_41741,N_40276);
nand U42088 (N_42088,N_41171,N_40464);
or U42089 (N_42089,N_41479,N_41961);
xnor U42090 (N_42090,N_41674,N_41450);
nor U42091 (N_42091,N_41063,N_40846);
xor U42092 (N_42092,N_40402,N_40207);
xnor U42093 (N_42093,N_41039,N_41494);
nand U42094 (N_42094,N_40419,N_41327);
nor U42095 (N_42095,N_41227,N_41701);
nand U42096 (N_42096,N_41410,N_41642);
nor U42097 (N_42097,N_41806,N_41983);
nand U42098 (N_42098,N_40760,N_41496);
nand U42099 (N_42099,N_40585,N_41693);
and U42100 (N_42100,N_41107,N_40428);
and U42101 (N_42101,N_41239,N_41332);
and U42102 (N_42102,N_40874,N_41635);
nor U42103 (N_42103,N_40268,N_40294);
nand U42104 (N_42104,N_40727,N_41922);
nor U42105 (N_42105,N_41729,N_41286);
xnor U42106 (N_42106,N_40209,N_41669);
or U42107 (N_42107,N_40270,N_41202);
or U42108 (N_42108,N_41413,N_40997);
nand U42109 (N_42109,N_40615,N_41688);
and U42110 (N_42110,N_41639,N_41765);
xnor U42111 (N_42111,N_40163,N_40618);
and U42112 (N_42112,N_41915,N_40810);
xor U42113 (N_42113,N_40617,N_41667);
and U42114 (N_42114,N_41290,N_41217);
nand U42115 (N_42115,N_40093,N_40406);
nor U42116 (N_42116,N_40080,N_40573);
xor U42117 (N_42117,N_40112,N_40978);
and U42118 (N_42118,N_40244,N_40853);
nor U42119 (N_42119,N_41969,N_41241);
nor U42120 (N_42120,N_40914,N_41229);
and U42121 (N_42121,N_40015,N_41192);
nor U42122 (N_42122,N_40994,N_41976);
nor U42123 (N_42123,N_41231,N_41708);
or U42124 (N_42124,N_41436,N_40873);
nand U42125 (N_42125,N_41368,N_41260);
nor U42126 (N_42126,N_40170,N_41582);
nor U42127 (N_42127,N_40883,N_40324);
nor U42128 (N_42128,N_40310,N_41676);
and U42129 (N_42129,N_41177,N_41132);
xor U42130 (N_42130,N_41947,N_40179);
and U42131 (N_42131,N_40471,N_40254);
nand U42132 (N_42132,N_41011,N_41681);
nand U42133 (N_42133,N_40519,N_40542);
nand U42134 (N_42134,N_40752,N_41308);
xnor U42135 (N_42135,N_41261,N_41986);
nor U42136 (N_42136,N_40601,N_41205);
xor U42137 (N_42137,N_40770,N_41973);
xor U42138 (N_42138,N_41834,N_41431);
nor U42139 (N_42139,N_40053,N_41380);
xor U42140 (N_42140,N_41900,N_41946);
or U42141 (N_42141,N_41330,N_41117);
or U42142 (N_42142,N_41147,N_40413);
xor U42143 (N_42143,N_40694,N_41106);
xor U42144 (N_42144,N_41129,N_40332);
or U42145 (N_42145,N_41065,N_40541);
nand U42146 (N_42146,N_40579,N_41162);
and U42147 (N_42147,N_40424,N_41491);
nand U42148 (N_42148,N_40527,N_40913);
nor U42149 (N_42149,N_41890,N_41520);
and U42150 (N_42150,N_40957,N_40535);
nor U42151 (N_42151,N_40256,N_40713);
nor U42152 (N_42152,N_40295,N_41285);
nor U42153 (N_42153,N_40232,N_40832);
xnor U42154 (N_42154,N_41933,N_40676);
nand U42155 (N_42155,N_41118,N_41838);
nor U42156 (N_42156,N_41930,N_40441);
xnor U42157 (N_42157,N_40800,N_41994);
and U42158 (N_42158,N_41583,N_41213);
or U42159 (N_42159,N_40987,N_40172);
xor U42160 (N_42160,N_41180,N_40333);
xnor U42161 (N_42161,N_40644,N_41033);
nand U42162 (N_42162,N_40799,N_41732);
xor U42163 (N_42163,N_40111,N_40879);
xnor U42164 (N_42164,N_40885,N_40133);
xor U42165 (N_42165,N_40952,N_41607);
or U42166 (N_42166,N_40423,N_40139);
nor U42167 (N_42167,N_40841,N_41679);
xnor U42168 (N_42168,N_41775,N_40507);
or U42169 (N_42169,N_41090,N_40935);
or U42170 (N_42170,N_41186,N_41443);
or U42171 (N_42171,N_41909,N_40765);
and U42172 (N_42172,N_41415,N_40998);
xnor U42173 (N_42173,N_41626,N_41610);
nor U42174 (N_42174,N_41121,N_40132);
nand U42175 (N_42175,N_41547,N_41312);
or U42176 (N_42176,N_41892,N_41164);
xor U42177 (N_42177,N_40831,N_40493);
or U42178 (N_42178,N_41665,N_40548);
or U42179 (N_42179,N_41247,N_40038);
or U42180 (N_42180,N_41889,N_40146);
and U42181 (N_42181,N_40524,N_41458);
xnor U42182 (N_42182,N_40346,N_40967);
nor U42183 (N_42183,N_40578,N_40759);
nor U42184 (N_42184,N_40897,N_41737);
nand U42185 (N_42185,N_41784,N_41370);
or U42186 (N_42186,N_41387,N_40287);
nand U42187 (N_42187,N_40556,N_41847);
or U42188 (N_42188,N_40911,N_40247);
nor U42189 (N_42189,N_41707,N_41868);
or U42190 (N_42190,N_40126,N_41066);
nand U42191 (N_42191,N_41883,N_40042);
xnor U42192 (N_42192,N_40300,N_41103);
and U42193 (N_42193,N_41621,N_41255);
nand U42194 (N_42194,N_41636,N_40708);
nand U42195 (N_42195,N_40545,N_40495);
xor U42196 (N_42196,N_41704,N_41975);
nor U42197 (N_42197,N_41021,N_40145);
xor U42198 (N_42198,N_41828,N_41897);
and U42199 (N_42199,N_40589,N_41644);
nand U42200 (N_42200,N_41997,N_41489);
and U42201 (N_42201,N_41159,N_41024);
or U42202 (N_42202,N_41685,N_41219);
nor U42203 (N_42203,N_40864,N_40410);
nand U42204 (N_42204,N_40855,N_40964);
nand U42205 (N_42205,N_41706,N_41244);
or U42206 (N_42206,N_41781,N_41796);
or U42207 (N_42207,N_41061,N_40730);
nand U42208 (N_42208,N_40555,N_40494);
and U42209 (N_42209,N_41764,N_40550);
and U42210 (N_42210,N_40060,N_41613);
or U42211 (N_42211,N_40129,N_41154);
and U42212 (N_42212,N_40085,N_40466);
or U42213 (N_42213,N_40435,N_41277);
and U42214 (N_42214,N_40695,N_40587);
nand U42215 (N_42215,N_41991,N_41861);
xor U42216 (N_42216,N_40588,N_41966);
or U42217 (N_42217,N_40261,N_40095);
or U42218 (N_42218,N_40681,N_40762);
or U42219 (N_42219,N_40448,N_40279);
or U42220 (N_42220,N_41910,N_41357);
nand U42221 (N_42221,N_41603,N_40055);
xnor U42222 (N_42222,N_40195,N_40833);
and U42223 (N_42223,N_40923,N_41697);
and U42224 (N_42224,N_40784,N_40652);
and U42225 (N_42225,N_41441,N_41541);
nor U42226 (N_42226,N_40280,N_40297);
xnor U42227 (N_42227,N_41735,N_40736);
nand U42228 (N_42228,N_41067,N_41618);
and U42229 (N_42229,N_41495,N_40812);
nor U42230 (N_42230,N_41843,N_41376);
xor U42231 (N_42231,N_40278,N_41267);
xor U42232 (N_42232,N_41989,N_41896);
or U42233 (N_42233,N_40315,N_40263);
or U42234 (N_42234,N_40778,N_41367);
and U42235 (N_42235,N_41348,N_40749);
nor U42236 (N_42236,N_40175,N_41388);
and U42237 (N_42237,N_40193,N_40005);
or U42238 (N_42238,N_40742,N_40344);
or U42239 (N_42239,N_40600,N_41058);
xor U42240 (N_42240,N_41266,N_40806);
and U42241 (N_42241,N_41733,N_40272);
nor U42242 (N_42242,N_41478,N_41533);
nor U42243 (N_42243,N_41875,N_40404);
nand U42244 (N_42244,N_41315,N_41694);
nand U42245 (N_42245,N_41015,N_40417);
xor U42246 (N_42246,N_40131,N_41654);
xnor U42247 (N_42247,N_40202,N_41082);
nand U42248 (N_42248,N_40288,N_40996);
nand U42249 (N_42249,N_41451,N_40469);
nand U42250 (N_42250,N_40583,N_40616);
or U42251 (N_42251,N_40106,N_41251);
or U42252 (N_42252,N_40071,N_40699);
nor U42253 (N_42253,N_40366,N_41867);
nor U42254 (N_42254,N_41633,N_41175);
nor U42255 (N_42255,N_40851,N_40636);
nand U42256 (N_42256,N_41770,N_41731);
xor U42257 (N_42257,N_41931,N_41439);
xnor U42258 (N_42258,N_41866,N_40926);
and U42259 (N_42259,N_41371,N_41340);
xor U42260 (N_42260,N_41466,N_40933);
and U42261 (N_42261,N_40839,N_41762);
xnor U42262 (N_42262,N_40523,N_40274);
xor U42263 (N_42263,N_40500,N_40385);
or U42264 (N_42264,N_41881,N_40237);
or U42265 (N_42265,N_41675,N_40758);
xnor U42266 (N_42266,N_40050,N_40031);
nor U42267 (N_42267,N_41259,N_40461);
nand U42268 (N_42268,N_41150,N_41884);
nand U42269 (N_42269,N_40698,N_40837);
nand U42270 (N_42270,N_40847,N_40322);
nand U42271 (N_42271,N_40025,N_41373);
or U42272 (N_42272,N_40326,N_40943);
or U42273 (N_42273,N_41409,N_40271);
or U42274 (N_42274,N_40491,N_40656);
and U42275 (N_42275,N_41941,N_41502);
and U42276 (N_42276,N_40484,N_41222);
or U42277 (N_42277,N_41906,N_40642);
nor U42278 (N_42278,N_40186,N_41477);
nor U42279 (N_42279,N_41456,N_40342);
and U42280 (N_42280,N_41097,N_41759);
nand U42281 (N_42281,N_41629,N_41321);
nand U42282 (N_42282,N_40375,N_41929);
nor U42283 (N_42283,N_41385,N_40230);
and U42284 (N_42284,N_41017,N_41280);
nor U42285 (N_42285,N_40744,N_40361);
nand U42286 (N_42286,N_41026,N_41510);
nor U42287 (N_42287,N_40970,N_40290);
xor U42288 (N_42288,N_41377,N_41084);
or U42289 (N_42289,N_40769,N_40668);
and U42290 (N_42290,N_40125,N_40819);
or U42291 (N_42291,N_40974,N_41482);
and U42292 (N_42292,N_41009,N_40684);
and U42293 (N_42293,N_40169,N_40450);
nand U42294 (N_42294,N_40360,N_41543);
nor U42295 (N_42295,N_40956,N_40307);
nand U42296 (N_42296,N_40395,N_40657);
nand U42297 (N_42297,N_40989,N_40786);
and U42298 (N_42298,N_41006,N_40192);
xor U42299 (N_42299,N_40604,N_41437);
and U42300 (N_42300,N_40845,N_41880);
nand U42301 (N_42301,N_40626,N_40510);
and U42302 (N_42302,N_40219,N_40825);
or U42303 (N_42303,N_41156,N_41396);
nor U42304 (N_42304,N_40433,N_40856);
nand U42305 (N_42305,N_40137,N_40766);
nand U42306 (N_42306,N_40852,N_41604);
nand U42307 (N_42307,N_40403,N_41390);
or U42308 (N_42308,N_40737,N_40705);
xnor U42309 (N_42309,N_40205,N_41418);
nand U42310 (N_42310,N_40795,N_40303);
nand U42311 (N_42311,N_41158,N_40909);
xor U42312 (N_42312,N_40334,N_41183);
nor U42313 (N_42313,N_40569,N_40993);
nand U42314 (N_42314,N_41663,N_41209);
nand U42315 (N_42315,N_41666,N_41027);
and U42316 (N_42316,N_41101,N_40678);
nand U42317 (N_42317,N_41073,N_40458);
nor U42318 (N_42318,N_40824,N_40418);
xor U42319 (N_42319,N_40214,N_40865);
or U42320 (N_42320,N_41453,N_41328);
nor U42321 (N_42321,N_41475,N_41905);
nand U42322 (N_42322,N_41601,N_41934);
or U42323 (N_42323,N_40777,N_41965);
and U42324 (N_42324,N_40317,N_40718);
or U42325 (N_42325,N_41137,N_41135);
nand U42326 (N_42326,N_40249,N_41360);
nor U42327 (N_42327,N_40960,N_40975);
xor U42328 (N_42328,N_41394,N_40000);
and U42329 (N_42329,N_41372,N_41263);
or U42330 (N_42330,N_40862,N_41078);
or U42331 (N_42331,N_41144,N_41054);
xnor U42332 (N_42332,N_40581,N_40104);
xor U42333 (N_42333,N_40432,N_41856);
and U42334 (N_42334,N_41913,N_40866);
xnor U42335 (N_42335,N_41578,N_40741);
and U42336 (N_42336,N_41959,N_40014);
nor U42337 (N_42337,N_40343,N_40614);
and U42338 (N_42338,N_41157,N_40798);
and U42339 (N_42339,N_40246,N_41822);
and U42340 (N_42340,N_40697,N_41303);
and U42341 (N_42341,N_41873,N_40154);
or U42342 (N_42342,N_41800,N_41787);
xnor U42343 (N_42343,N_40099,N_41457);
or U42344 (N_42344,N_40599,N_40683);
nor U42345 (N_42345,N_41254,N_40962);
nor U42346 (N_42346,N_41661,N_41352);
nand U42347 (N_42347,N_41808,N_41987);
xnor U42348 (N_42348,N_40506,N_40181);
xnor U42349 (N_42349,N_41166,N_41146);
and U42350 (N_42350,N_40893,N_41795);
and U42351 (N_42351,N_41819,N_40226);
xor U42352 (N_42352,N_41374,N_40144);
nand U42353 (N_42353,N_41230,N_40714);
nand U42354 (N_42354,N_41019,N_41734);
or U42355 (N_42355,N_41165,N_41627);
nor U42356 (N_42356,N_41712,N_41128);
or U42357 (N_42357,N_41356,N_41754);
nand U42358 (N_42358,N_41087,N_40582);
nand U42359 (N_42359,N_41840,N_40575);
and U42360 (N_42360,N_40946,N_40150);
and U42361 (N_42361,N_41163,N_40574);
and U42362 (N_42362,N_41126,N_40942);
nor U42363 (N_42363,N_41358,N_41282);
and U42364 (N_42364,N_40529,N_41778);
nor U42365 (N_42365,N_41608,N_41649);
and U42366 (N_42366,N_41782,N_40189);
or U42367 (N_42367,N_41853,N_41074);
or U42368 (N_42368,N_41235,N_41777);
or U42369 (N_42369,N_41518,N_41785);
nand U42370 (N_42370,N_41937,N_41023);
xnor U42371 (N_42371,N_41234,N_41531);
nor U42372 (N_42372,N_41306,N_40539);
nand U42373 (N_42373,N_41049,N_40944);
nor U42374 (N_42374,N_40880,N_41329);
nand U42375 (N_42375,N_41817,N_41728);
xor U42376 (N_42376,N_40750,N_40048);
and U42377 (N_42377,N_41748,N_40628);
and U42378 (N_42378,N_41297,N_41561);
nand U42379 (N_42379,N_40870,N_41029);
and U42380 (N_42380,N_40298,N_40498);
nor U42381 (N_42381,N_40525,N_40468);
or U42382 (N_42382,N_41152,N_40844);
nor U42383 (N_42383,N_41110,N_41891);
nor U42384 (N_42384,N_40400,N_40659);
nand U42385 (N_42385,N_41485,N_40543);
nor U42386 (N_42386,N_40783,N_40266);
or U42387 (N_42387,N_40850,N_41919);
or U42388 (N_42388,N_40508,N_40399);
xnor U42389 (N_42389,N_40330,N_41597);
and U42390 (N_42390,N_41378,N_40664);
and U42391 (N_42391,N_41236,N_41355);
or U42392 (N_42392,N_40028,N_41739);
nor U42393 (N_42393,N_41115,N_40653);
or U42394 (N_42394,N_41928,N_41824);
and U42395 (N_42395,N_40379,N_40961);
and U42396 (N_42396,N_40827,N_40225);
or U42397 (N_42397,N_41226,N_40396);
and U42398 (N_42398,N_41750,N_41326);
nand U42399 (N_42399,N_41199,N_40667);
and U42400 (N_42400,N_40632,N_41588);
nand U42401 (N_42401,N_41412,N_40073);
xor U42402 (N_42402,N_41203,N_40475);
or U42403 (N_42403,N_41480,N_40184);
nand U42404 (N_42404,N_41574,N_40118);
and U42405 (N_42405,N_40138,N_41408);
nor U42406 (N_42406,N_40459,N_41407);
xnor U42407 (N_42407,N_40089,N_41270);
nand U42408 (N_42408,N_40701,N_41823);
nor U42409 (N_42409,N_40002,N_40216);
xor U42410 (N_42410,N_41577,N_41493);
nand U42411 (N_42411,N_41514,N_40155);
nor U42412 (N_42412,N_41316,N_40408);
and U42413 (N_42413,N_40711,N_41148);
xor U42414 (N_42414,N_40592,N_40840);
xor U42415 (N_42415,N_41894,N_40560);
xnor U42416 (N_42416,N_40492,N_40380);
or U42417 (N_42417,N_40003,N_40905);
nand U42418 (N_42418,N_40834,N_40745);
and U42419 (N_42419,N_40958,N_41172);
nand U42420 (N_42420,N_40212,N_41978);
or U42421 (N_42421,N_40439,N_41403);
xnor U42422 (N_42422,N_40820,N_40647);
xnor U42423 (N_42423,N_41826,N_41513);
nand U42424 (N_42424,N_41419,N_40082);
xnor U42425 (N_42425,N_41564,N_41014);
xor U42426 (N_42426,N_41791,N_40917);
nor U42427 (N_42427,N_41473,N_40415);
or U42428 (N_42428,N_41522,N_41013);
nand U42429 (N_42429,N_40901,N_41500);
xor U42430 (N_42430,N_40140,N_41050);
and U42431 (N_42431,N_40327,N_40382);
and U42432 (N_42432,N_40661,N_41532);
nand U42433 (N_42433,N_40160,N_41446);
xor U42434 (N_42434,N_40335,N_41651);
xnor U42435 (N_42435,N_40098,N_41744);
xor U42436 (N_42436,N_40672,N_40731);
xnor U42437 (N_42437,N_40563,N_41141);
nor U42438 (N_42438,N_40135,N_40635);
or U42439 (N_42439,N_40503,N_40971);
and U42440 (N_42440,N_40057,N_41302);
nor U42441 (N_42441,N_41099,N_41818);
nor U42442 (N_42442,N_41250,N_40097);
nor U42443 (N_42443,N_40729,N_40319);
or U42444 (N_42444,N_41766,N_40984);
or U42445 (N_42445,N_41363,N_40358);
nor U42446 (N_42446,N_41127,N_41151);
or U42447 (N_42447,N_40690,N_41570);
xor U42448 (N_42448,N_41365,N_41758);
or U42449 (N_42449,N_41469,N_40995);
xnor U42450 (N_42450,N_41193,N_41515);
nor U42451 (N_42451,N_41908,N_41421);
and U42452 (N_42452,N_41558,N_41974);
or U42453 (N_42453,N_40191,N_41562);
xnor U42454 (N_42454,N_41657,N_41225);
and U42455 (N_42455,N_41022,N_40876);
nor U42456 (N_42456,N_41804,N_40309);
nor U42457 (N_42457,N_40609,N_40362);
nand U42458 (N_42458,N_40159,N_41401);
xor U42459 (N_42459,N_40781,N_41695);
and U42460 (N_42460,N_41342,N_40046);
nand U42461 (N_42461,N_40811,N_40584);
xor U42462 (N_42462,N_40252,N_40505);
nor U42463 (N_42463,N_40738,N_41503);
nand U42464 (N_42464,N_40117,N_40122);
nor U42465 (N_42465,N_40381,N_40848);
xnor U42466 (N_42466,N_40292,N_40536);
nor U42467 (N_42467,N_40058,N_41549);
and U42468 (N_42468,N_40677,N_40571);
and U42469 (N_42469,N_41007,N_41105);
nand U42470 (N_42470,N_40687,N_41333);
or U42471 (N_42471,N_40483,N_40026);
xor U42472 (N_42472,N_41470,N_41000);
or U42473 (N_42473,N_41104,N_40836);
and U42474 (N_42474,N_41977,N_41004);
or U42475 (N_42475,N_41349,N_40564);
or U42476 (N_42476,N_40512,N_41420);
or U42477 (N_42477,N_40001,N_41671);
xor U42478 (N_42478,N_40357,N_41999);
nor U42479 (N_42479,N_41318,N_41249);
nor U42480 (N_42480,N_41181,N_41080);
and U42481 (N_42481,N_40992,N_41723);
nor U42482 (N_42482,N_41952,N_41094);
nor U42483 (N_42483,N_40710,N_41539);
and U42484 (N_42484,N_40919,N_40894);
and U42485 (N_42485,N_40017,N_41346);
xor U42486 (N_42486,N_41170,N_40951);
nor U42487 (N_42487,N_40902,N_40052);
or U42488 (N_42488,N_40646,N_40177);
or U42489 (N_42489,N_40241,N_40047);
nor U42490 (N_42490,N_40480,N_41064);
nand U42491 (N_42491,N_40253,N_41273);
nor U42492 (N_42492,N_41526,N_40022);
xnor U42493 (N_42493,N_40349,N_41112);
nand U42494 (N_42494,N_41831,N_41085);
nand U42495 (N_42495,N_40056,N_41720);
nand U42496 (N_42496,N_41536,N_41591);
nand U42497 (N_42497,N_41611,N_41051);
xnor U42498 (N_42498,N_40688,N_40488);
and U42499 (N_42499,N_41851,N_40032);
nand U42500 (N_42500,N_40224,N_40457);
nor U42501 (N_42501,N_41113,N_41300);
nand U42502 (N_42502,N_40816,N_40389);
nor U42503 (N_42503,N_40113,N_41528);
nand U42504 (N_42504,N_40595,N_41963);
nand U42505 (N_42505,N_41645,N_40586);
xnor U42506 (N_42506,N_40544,N_41567);
nor U42507 (N_42507,N_41837,N_41246);
nand U42508 (N_42508,N_40829,N_41044);
nor U42509 (N_42509,N_40185,N_41210);
and U42510 (N_42510,N_40675,N_40359);
and U42511 (N_42511,N_41534,N_41812);
nand U42512 (N_42512,N_41815,N_41461);
xnor U42513 (N_42513,N_40221,N_41805);
nand U42514 (N_42514,N_41031,N_41709);
or U42515 (N_42515,N_40473,N_41003);
nor U42516 (N_42516,N_40557,N_40740);
or U42517 (N_42517,N_40814,N_41131);
and U42518 (N_42518,N_41590,N_41108);
and U42519 (N_42519,N_41673,N_41338);
or U42520 (N_42520,N_40904,N_41870);
or U42521 (N_42521,N_40096,N_41572);
nor U42522 (N_42522,N_41484,N_40891);
nor U42523 (N_42523,N_40559,N_40040);
and U42524 (N_42524,N_40692,N_41958);
or U42525 (N_42525,N_40161,N_40449);
nor U42526 (N_42526,N_40603,N_41237);
and U42527 (N_42527,N_41350,N_40281);
xnor U42528 (N_42528,N_41659,N_41658);
nor U42529 (N_42529,N_40387,N_41030);
xnor U42530 (N_42530,N_40972,N_41717);
or U42531 (N_42531,N_41631,N_40369);
or U42532 (N_42532,N_41816,N_41985);
or U42533 (N_42533,N_40818,N_40455);
xor U42534 (N_42534,N_40102,N_41620);
xor U42535 (N_42535,N_40265,N_40763);
nor U42536 (N_42536,N_41416,N_41323);
or U42537 (N_42537,N_40101,N_41914);
and U42538 (N_42538,N_40474,N_41417);
xnor U42539 (N_42539,N_40045,N_41797);
nand U42540 (N_42540,N_40233,N_41788);
or U42541 (N_42541,N_41519,N_40054);
nor U42542 (N_42542,N_40210,N_41716);
nand U42543 (N_42543,N_40064,N_40947);
or U42544 (N_42544,N_41895,N_41295);
xnor U42545 (N_42545,N_41619,N_40308);
xor U42546 (N_42546,N_41271,N_41499);
nand U42547 (N_42547,N_41814,N_41967);
nand U42548 (N_42548,N_41335,N_41957);
and U42549 (N_42549,N_40420,N_41092);
or U42550 (N_42550,N_40815,N_41845);
and U42551 (N_42551,N_40320,N_41801);
nor U42552 (N_42552,N_41045,N_41691);
xor U42553 (N_42553,N_41467,N_40092);
or U42554 (N_42554,N_40884,N_41992);
or U42555 (N_42555,N_41311,N_40255);
xnor U42556 (N_42556,N_41072,N_40051);
nor U42557 (N_42557,N_40932,N_41972);
nand U42558 (N_42558,N_40963,N_40822);
and U42559 (N_42559,N_40044,N_41768);
nor U42560 (N_42560,N_40134,N_40401);
xor U42561 (N_42561,N_40316,N_41869);
nor U42562 (N_42562,N_41507,N_40702);
nor U42563 (N_42563,N_41509,N_41444);
nor U42564 (N_42564,N_40789,N_41043);
and U42565 (N_42565,N_40291,N_40700);
xor U42566 (N_42566,N_40454,N_40966);
xnor U42567 (N_42567,N_41556,N_40321);
and U42568 (N_42568,N_40328,N_41490);
nor U42569 (N_42569,N_40090,N_41454);
nor U42570 (N_42570,N_40842,N_40639);
xor U42571 (N_42571,N_40036,N_41429);
and U42572 (N_42572,N_41689,N_40465);
xnor U42573 (N_42573,N_40877,N_40638);
nand U42574 (N_42574,N_41130,N_40075);
and U42575 (N_42575,N_40345,N_40183);
and U42576 (N_42576,N_40062,N_41641);
nand U42577 (N_42577,N_40367,N_41529);
xnor U42578 (N_42578,N_41088,N_41191);
nor U42579 (N_42579,N_40509,N_41245);
nor U42580 (N_42580,N_40983,N_40733);
xnor U42581 (N_42581,N_40477,N_41757);
and U42582 (N_42582,N_41395,N_40857);
xnor U42583 (N_42583,N_40912,N_40472);
or U42584 (N_42584,N_41690,N_41476);
nand U42585 (N_42585,N_40934,N_40302);
xnor U42586 (N_42586,N_40598,N_40826);
or U42587 (N_42587,N_41028,N_41120);
nor U42588 (N_42588,N_40086,N_40120);
and U42589 (N_42589,N_41176,N_41882);
xor U42590 (N_42590,N_41354,N_41672);
xor U42591 (N_42591,N_41979,N_40442);
nor U42592 (N_42592,N_40776,N_40236);
nand U42593 (N_42593,N_40889,N_41783);
or U42594 (N_42594,N_40444,N_41647);
and U42595 (N_42595,N_41319,N_41736);
and U42596 (N_42596,N_41576,N_41625);
nand U42597 (N_42597,N_40860,N_40669);
xnor U42598 (N_42598,N_41272,N_41652);
nor U42599 (N_42599,N_41719,N_41143);
nand U42600 (N_42600,N_40059,N_40872);
xor U42601 (N_42601,N_40517,N_41086);
nor U42602 (N_42602,N_41511,N_40035);
and U42603 (N_42603,N_40147,N_41362);
xor U42604 (N_42604,N_40376,N_40903);
nor U42605 (N_42605,N_41208,N_40447);
nand U42606 (N_42606,N_41696,N_40124);
or U42607 (N_42607,N_41501,N_41859);
nor U42608 (N_42608,N_40220,N_41648);
xnor U42609 (N_42609,N_41483,N_41037);
or U42610 (N_42610,N_40323,N_40734);
nand U42611 (N_42611,N_41460,N_41833);
xor U42612 (N_42612,N_40787,N_41102);
xor U42613 (N_42613,N_41046,N_41070);
or U42614 (N_42614,N_41664,N_41305);
nor U42615 (N_42615,N_41424,N_41761);
nand U42616 (N_42616,N_40674,N_40446);
and U42617 (N_42617,N_40213,N_41569);
nand U42618 (N_42618,N_41299,N_41885);
or U42619 (N_42619,N_40565,N_40533);
xnor U42620 (N_42620,N_41727,N_41005);
nor U42621 (N_42621,N_41016,N_41449);
nor U42622 (N_42622,N_40105,N_41081);
and U42623 (N_42623,N_41292,N_41863);
nand U42624 (N_42624,N_41508,N_41911);
nand U42625 (N_42625,N_41988,N_40801);
nand U42626 (N_42626,N_41705,N_40553);
and U42627 (N_42627,N_41149,N_40016);
nand U42628 (N_42628,N_40547,N_41339);
or U42629 (N_42629,N_41012,N_40928);
nor U42630 (N_42630,N_41060,N_40426);
or U42631 (N_42631,N_40940,N_41252);
nand U42632 (N_42632,N_41274,N_41568);
and U42633 (N_42633,N_40620,N_40453);
nand U42634 (N_42634,N_40716,N_40130);
or U42635 (N_42635,N_40723,N_40892);
and U42636 (N_42636,N_41196,N_40227);
and U42637 (N_42637,N_40019,N_40792);
and U42638 (N_42638,N_40937,N_40467);
xor U42639 (N_42639,N_40083,N_40651);
nand U42640 (N_42640,N_41430,N_40722);
xor U42641 (N_42641,N_40514,N_40421);
or U42642 (N_42642,N_41842,N_41153);
and U42643 (N_42643,N_41512,N_40613);
nor U42644 (N_42644,N_40597,N_40114);
nor U42645 (N_42645,N_41923,N_40091);
nor U42646 (N_42646,N_40910,N_40416);
nand U42647 (N_42647,N_40924,N_40772);
or U42648 (N_42648,N_41980,N_41083);
and U42649 (N_42649,N_41742,N_40925);
and U42650 (N_42650,N_40761,N_40081);
and U42651 (N_42651,N_41293,N_41123);
nand U42652 (N_42652,N_41920,N_40094);
nor U42653 (N_42653,N_41075,N_41331);
nor U42654 (N_42654,N_41713,N_41700);
or U42655 (N_42655,N_40438,N_41609);
or U42656 (N_42656,N_40338,N_41835);
nand U42657 (N_42657,N_40930,N_40121);
and U42658 (N_42658,N_41901,N_41573);
and U42659 (N_42659,N_40078,N_40049);
xnor U42660 (N_42660,N_40486,N_41763);
and U42661 (N_42661,N_41369,N_41848);
nor U42662 (N_42662,N_40607,N_41337);
nor U42663 (N_42663,N_40347,N_41655);
nor U42664 (N_42664,N_40838,N_41160);
and U42665 (N_42665,N_40869,N_40709);
xnor U42666 (N_42666,N_41802,N_41793);
nor U42667 (N_42667,N_40187,N_41760);
xnor U42668 (N_42668,N_41215,N_41893);
nand U42669 (N_42669,N_41579,N_41552);
or U42670 (N_42670,N_40364,N_41907);
or U42671 (N_42671,N_40411,N_40182);
xnor U42672 (N_42672,N_41076,N_41904);
or U42673 (N_42673,N_41100,N_41268);
nand U42674 (N_42674,N_40854,N_40828);
xnor U42675 (N_42675,N_40712,N_41811);
nor U42676 (N_42676,N_41774,N_40128);
nor U42677 (N_42677,N_41048,N_40888);
nand U42678 (N_42678,N_41411,N_40074);
or U42679 (N_42679,N_40299,N_41686);
or U42680 (N_42680,N_41710,N_40431);
and U42681 (N_42681,N_41580,N_41598);
nor U42682 (N_42682,N_40732,N_41351);
and U42683 (N_42683,N_40679,N_41269);
and U42684 (N_42684,N_41020,N_41595);
and U42685 (N_42685,N_41279,N_41364);
nand U42686 (N_42686,N_41938,N_41968);
or U42687 (N_42687,N_40532,N_41145);
and U42688 (N_42688,N_40243,N_40029);
and U42689 (N_42689,N_40264,N_41402);
nor U42690 (N_42690,N_40470,N_41738);
or U42691 (N_42691,N_40719,N_40568);
nor U42692 (N_42692,N_41125,N_41699);
and U42693 (N_42693,N_41038,N_40823);
xnor U42694 (N_42694,N_40378,N_41771);
xnor U42695 (N_42695,N_40821,N_40277);
or U42696 (N_42696,N_41262,N_40394);
nand U42697 (N_42697,N_40240,N_41602);
or U42698 (N_42698,N_40813,N_41898);
or U42699 (N_42699,N_40217,N_40939);
xor U42700 (N_42700,N_40251,N_41950);
or U42701 (N_42701,N_41301,N_40371);
and U42702 (N_42702,N_41646,N_40631);
xor U42703 (N_42703,N_40076,N_40430);
nand U42704 (N_42704,N_40955,N_40570);
and U42705 (N_42705,N_40107,N_40282);
and U42706 (N_42706,N_40286,N_41310);
or U42707 (N_42707,N_40437,N_40649);
nor U42708 (N_42708,N_41468,N_40878);
nor U42709 (N_42709,N_41207,N_41139);
nand U42710 (N_42710,N_41943,N_40393);
nand U42711 (N_42711,N_40728,N_41492);
and U42712 (N_42712,N_41284,N_41546);
or U42713 (N_42713,N_41545,N_41010);
and U42714 (N_42714,N_40685,N_41433);
nor U42715 (N_42715,N_40171,N_40965);
or U42716 (N_42716,N_40314,N_40671);
nand U42717 (N_42717,N_41256,N_40020);
nand U42718 (N_42718,N_40666,N_41275);
nor U42719 (N_42719,N_40008,N_40153);
nand U42720 (N_42720,N_40397,N_41178);
nor U42721 (N_42721,N_41109,N_40779);
or U42722 (N_42722,N_41442,N_41813);
nand U42723 (N_42723,N_41982,N_40907);
or U42724 (N_42724,N_40296,N_41698);
and U42725 (N_42725,N_41098,N_41810);
nand U42726 (N_42726,N_41487,N_40391);
nand U42727 (N_42727,N_40250,N_41786);
or U42728 (N_42728,N_41384,N_40858);
xor U42729 (N_42729,N_41628,N_41852);
and U42730 (N_42730,N_40501,N_40068);
or U42731 (N_42731,N_41382,N_41560);
and U42732 (N_42732,N_41530,N_40203);
nor U42733 (N_42733,N_40165,N_40895);
nand U42734 (N_42734,N_41584,N_41702);
nor U42735 (N_42735,N_41971,N_40531);
nand U42736 (N_42736,N_40518,N_40788);
and U42737 (N_42737,N_40198,N_40260);
nand U42738 (N_42738,N_41397,N_40222);
nand U42739 (N_42739,N_40790,N_41119);
nand U42740 (N_42740,N_40868,N_41854);
nor U42741 (N_42741,N_41096,N_41767);
nor U42742 (N_42742,N_41497,N_41551);
xor U42743 (N_42743,N_41535,N_41612);
nand U42744 (N_42744,N_40511,N_40499);
or U42745 (N_42745,N_40353,N_41223);
xnor U42746 (N_42746,N_41990,N_41902);
and U42747 (N_42747,N_40941,N_41692);
xor U42748 (N_42748,N_41939,N_40881);
and U42749 (N_42749,N_40549,N_41916);
and U42750 (N_42750,N_41538,N_41212);
xnor U42751 (N_42751,N_40033,N_41721);
or U42752 (N_42752,N_40830,N_40136);
nand U42753 (N_42753,N_40643,N_41258);
or U42754 (N_42754,N_41353,N_40304);
and U42755 (N_42755,N_41198,N_40988);
xnor U42756 (N_42756,N_41876,N_40009);
nor U42757 (N_42757,N_41593,N_41550);
nand U42758 (N_42758,N_40673,N_40562);
or U42759 (N_42759,N_40665,N_41114);
nor U42760 (N_42760,N_41638,N_40027);
and U42761 (N_42761,N_40650,N_40331);
nor U42762 (N_42762,N_41383,N_40151);
and U42763 (N_42763,N_41724,N_40370);
or U42764 (N_42764,N_40982,N_40043);
or U42765 (N_42765,N_40640,N_40239);
xnor U42766 (N_42766,N_41122,N_40365);
nor U42767 (N_42767,N_41780,N_41940);
nand U42768 (N_42768,N_41294,N_40110);
and U42769 (N_42769,N_40325,N_41111);
nand U42770 (N_42770,N_40482,N_40502);
and U42771 (N_42771,N_41858,N_40348);
xnor U42772 (N_42772,N_41445,N_40624);
or U42773 (N_42773,N_41216,N_41836);
nor U42774 (N_42774,N_40720,N_41962);
nand U42775 (N_42775,N_41711,N_40340);
nor U42776 (N_42776,N_40630,N_41917);
and U42777 (N_42777,N_40223,N_40796);
or U42778 (N_42778,N_41656,N_41240);
nand U42779 (N_42779,N_40746,N_40258);
and U42780 (N_42780,N_41745,N_41304);
and U42781 (N_42781,N_41291,N_41877);
xnor U42782 (N_42782,N_41317,N_41945);
nor U42783 (N_42783,N_40981,N_41924);
nor U42784 (N_42784,N_40538,N_41566);
or U42785 (N_42785,N_41435,N_41392);
and U42786 (N_42786,N_41918,N_40141);
nand U42787 (N_42787,N_41228,N_40339);
nand U42788 (N_42788,N_41422,N_41622);
or U42789 (N_42789,N_40959,N_41521);
xnor U42790 (N_42790,N_40526,N_40504);
or U42791 (N_42791,N_41951,N_41243);
nand U42792 (N_42792,N_40476,N_41798);
nand U42793 (N_42793,N_41440,N_41587);
or U42794 (N_42794,N_41124,N_41872);
or U42795 (N_42795,N_41195,N_40691);
nor U42796 (N_42796,N_40072,N_40497);
xnor U42797 (N_42797,N_41002,N_41347);
or U42798 (N_42798,N_40351,N_40530);
nand U42799 (N_42799,N_40242,N_40686);
nand U42800 (N_42800,N_40301,N_41464);
or U42801 (N_42801,N_40337,N_40561);
and U42802 (N_42802,N_40528,N_40704);
and U42803 (N_42803,N_40100,N_40990);
and U42804 (N_42804,N_41265,N_41187);
nand U42805 (N_42805,N_40409,N_41498);
nor U42806 (N_42806,N_40929,N_41041);
nor U42807 (N_42807,N_41899,N_41359);
and U42808 (N_42808,N_40269,N_40915);
nor U42809 (N_42809,N_40696,N_41668);
and U42810 (N_42810,N_41718,N_41324);
or U42811 (N_42811,N_41554,N_40875);
xor U42812 (N_42812,N_40487,N_41730);
nor U42813 (N_42813,N_40229,N_40084);
nand U42814 (N_42814,N_40257,N_40496);
nand U42815 (N_42815,N_40899,N_40843);
nor U42816 (N_42816,N_41581,N_40780);
xor U42817 (N_42817,N_41888,N_41289);
nor U42818 (N_42818,N_41606,N_41472);
nor U42819 (N_42819,N_40024,N_41585);
and U42820 (N_42820,N_40576,N_41283);
and U42821 (N_42821,N_41517,N_40283);
nor U42822 (N_42822,N_40953,N_40754);
nand U42823 (N_42823,N_41662,N_40980);
nand U42824 (N_42824,N_40513,N_40887);
or U42825 (N_42825,N_41887,N_40516);
nor U42826 (N_42826,N_40802,N_40807);
and U42827 (N_42827,N_40079,N_40350);
and U42828 (N_42828,N_40372,N_41336);
and U42829 (N_42829,N_40977,N_41253);
or U42830 (N_42830,N_41343,N_40771);
or U42831 (N_42831,N_40262,N_40142);
nor U42832 (N_42832,N_41414,N_40341);
nand U42833 (N_42833,N_40554,N_41616);
or U42834 (N_42834,N_41211,N_41925);
xor U42835 (N_42835,N_40013,N_40594);
nand U42836 (N_42836,N_40390,N_40012);
xnor U42837 (N_42837,N_41185,N_41926);
xor U42838 (N_42838,N_41309,N_41134);
or U42839 (N_42839,N_40918,N_41307);
nor U42840 (N_42840,N_41204,N_41571);
and U42841 (N_42841,N_40030,N_41432);
nand U42842 (N_42842,N_40368,N_40273);
and U42843 (N_42843,N_40443,N_40006);
xnor U42844 (N_42844,N_40572,N_40927);
nor U42845 (N_42845,N_41427,N_41400);
xnor U42846 (N_42846,N_41643,N_41375);
nand U42847 (N_42847,N_41825,N_40969);
nor U42848 (N_42848,N_40794,N_41599);
nand U42849 (N_42849,N_40999,N_41555);
xnor U42850 (N_42850,N_40645,N_40007);
or U42851 (N_42851,N_40479,N_41506);
nor U42852 (N_42852,N_40921,N_41423);
xor U42853 (N_42853,N_40388,N_40178);
xor U42854 (N_42854,N_40234,N_41743);
nor U42855 (N_42855,N_41790,N_40735);
nand U42856 (N_42856,N_40384,N_41447);
nand U42857 (N_42857,N_40641,N_41189);
and U42858 (N_42858,N_40755,N_41653);
or U42859 (N_42859,N_40284,N_40920);
xor U42860 (N_42860,N_41703,N_41789);
or U42861 (N_42861,N_40148,N_40004);
or U42862 (N_42862,N_41179,N_40218);
nand U42863 (N_42863,N_41341,N_41953);
or U42864 (N_42864,N_40991,N_40774);
nand U42865 (N_42865,N_41794,N_40973);
nand U42866 (N_42866,N_40355,N_40011);
or U42867 (N_42867,N_41288,N_41055);
xnor U42868 (N_42868,N_40460,N_41630);
or U42869 (N_42869,N_40228,N_40577);
or U42870 (N_42870,N_41879,N_40063);
xor U42871 (N_42871,N_40551,N_40285);
and U42872 (N_42872,N_41042,N_41047);
xor U42873 (N_42873,N_40648,N_40398);
or U42874 (N_42874,N_40275,N_40289);
or U42875 (N_42875,N_41998,N_41773);
nor U42876 (N_42876,N_41849,N_41220);
nor U42877 (N_42877,N_40127,N_41116);
nor U42878 (N_42878,N_40552,N_40267);
nand U42879 (N_42879,N_41281,N_41886);
nand U42880 (N_42880,N_40445,N_40808);
nand U42881 (N_42881,N_41650,N_40039);
xor U42882 (N_42882,N_41314,N_40077);
nand U42883 (N_42883,N_41238,N_40634);
xor U42884 (N_42884,N_40606,N_41474);
and U42885 (N_42885,N_41184,N_41821);
nand U42886 (N_42886,N_41386,N_41932);
xnor U42887 (N_42887,N_40658,N_41248);
xor U42888 (N_42888,N_41725,N_41174);
nor U42889 (N_42889,N_41320,N_41960);
or U42890 (N_42890,N_40724,N_40670);
nor U42891 (N_42891,N_40065,N_41715);
and U42892 (N_42892,N_41448,N_40434);
and U42893 (N_42893,N_41434,N_40440);
and U42894 (N_42894,N_40190,N_41596);
nand U42895 (N_42895,N_40793,N_40429);
and U42896 (N_42896,N_41803,N_40849);
nand U42897 (N_42897,N_40149,N_41504);
xnor U42898 (N_42898,N_41264,N_41455);
or U42899 (N_42899,N_40896,N_40103);
or U42900 (N_42900,N_40313,N_40608);
nand U42901 (N_42901,N_41486,N_41169);
nand U42902 (N_42902,N_41034,N_41747);
xnor U42903 (N_42903,N_41188,N_40886);
and U42904 (N_42904,N_41623,N_40152);
nor U42905 (N_42905,N_41168,N_41525);
or U42906 (N_42906,N_41194,N_40088);
or U42907 (N_42907,N_40176,N_40034);
nor U42908 (N_42908,N_41334,N_41138);
nand U42909 (N_42909,N_40238,N_40605);
xnor U42910 (N_42910,N_40436,N_41632);
xnor U42911 (N_42911,N_40751,N_40451);
nand U42912 (N_42912,N_41605,N_40707);
nand U42913 (N_42913,N_40621,N_41772);
nand U42914 (N_42914,N_41036,N_41956);
nor U42915 (N_42915,N_40908,N_40021);
nor U42916 (N_42916,N_40123,N_40898);
or U42917 (N_42917,N_41995,N_41233);
or U42918 (N_42918,N_40739,N_40293);
and U42919 (N_42919,N_41830,N_40804);
or U42920 (N_42920,N_40515,N_41155);
xor U42921 (N_42921,N_40208,N_41970);
nor U42922 (N_42922,N_40383,N_40867);
nor U42923 (N_42923,N_40168,N_41799);
and U42924 (N_42924,N_41057,N_40143);
or U42925 (N_42925,N_41379,N_40197);
xor U42926 (N_42926,N_40619,N_40534);
and U42927 (N_42927,N_40906,N_41862);
nand U42928 (N_42928,N_40462,N_41366);
and U42929 (N_42929,N_40602,N_41594);
nor U42930 (N_42930,N_41524,N_41406);
and U42931 (N_42931,N_41874,N_41182);
xnor U42932 (N_42932,N_41553,N_41059);
nor U42933 (N_42933,N_41462,N_40954);
xor U42934 (N_42934,N_40116,N_41398);
xor U42935 (N_42935,N_41752,N_41592);
xor U42936 (N_42936,N_41865,N_40248);
nor U42937 (N_42937,N_40452,N_40627);
nand U42938 (N_42938,N_40871,N_40693);
nor U42939 (N_42939,N_41792,N_40188);
and U42940 (N_42940,N_41769,N_41197);
xnor U42941 (N_42941,N_40305,N_41871);
or U42942 (N_42942,N_41001,N_41313);
xor U42943 (N_42943,N_41381,N_40593);
and U42944 (N_42944,N_40235,N_40567);
xor U42945 (N_42945,N_40215,N_40196);
xor U42946 (N_42946,N_41405,N_41855);
or U42947 (N_42947,N_40119,N_41575);
nor U42948 (N_42948,N_40859,N_41589);
nor U42949 (N_42949,N_41173,N_41954);
and U42950 (N_42950,N_40623,N_41425);
xnor U42951 (N_42951,N_41544,N_40109);
or U42952 (N_42952,N_40726,N_40773);
and U42953 (N_42953,N_41841,N_40463);
nand U42954 (N_42954,N_40756,N_40882);
nand U42955 (N_42955,N_40157,N_40580);
nor U42956 (N_42956,N_40936,N_41682);
and U42957 (N_42957,N_40156,N_40162);
and U42958 (N_42958,N_41827,N_40861);
nor U42959 (N_42959,N_41563,N_41391);
and U42960 (N_42960,N_41018,N_41829);
or U42961 (N_42961,N_40743,N_41726);
nor U42962 (N_42962,N_41542,N_41614);
xor U42963 (N_42963,N_41221,N_40809);
or U42964 (N_42964,N_41740,N_40945);
nor U42965 (N_42965,N_40010,N_41949);
xnor U42966 (N_42966,N_41505,N_41749);
xor U42967 (N_42967,N_40922,N_41714);
nand U42968 (N_42968,N_40916,N_40245);
nor U42969 (N_42969,N_40158,N_41025);
or U42970 (N_42970,N_40311,N_41481);
nand U42971 (N_42971,N_41678,N_41089);
nor U42972 (N_42972,N_40478,N_41640);
nand U42973 (N_42973,N_40725,N_41981);
xnor U42974 (N_42974,N_41344,N_41200);
or U42975 (N_42975,N_40180,N_41944);
nor U42976 (N_42976,N_40489,N_40633);
nand U42977 (N_42977,N_41136,N_41809);
or U42978 (N_42978,N_40566,N_40204);
nor U42979 (N_42979,N_40986,N_41860);
or U42980 (N_42980,N_40863,N_40791);
nand U42981 (N_42981,N_40166,N_40405);
nor U42982 (N_42982,N_41540,N_40108);
nand U42983 (N_42983,N_40748,N_41548);
nand U42984 (N_42984,N_41298,N_41755);
nand U42985 (N_42985,N_40985,N_40422);
nor U42986 (N_42986,N_40485,N_40041);
xor U42987 (N_42987,N_40520,N_40596);
and U42988 (N_42988,N_40767,N_41722);
nand U42989 (N_42989,N_40625,N_40312);
or U42990 (N_42990,N_40018,N_40231);
and U42991 (N_42991,N_40329,N_41426);
nor U42992 (N_42992,N_40167,N_40540);
or U42993 (N_42993,N_41062,N_41091);
and U42994 (N_42994,N_41559,N_41680);
nand U42995 (N_42995,N_40206,N_40689);
nor U42996 (N_42996,N_40115,N_40392);
and U42997 (N_42997,N_40087,N_41278);
or U42998 (N_42998,N_41296,N_41839);
xor U42999 (N_42999,N_41537,N_40066);
nand U43000 (N_43000,N_40896,N_41929);
or U43001 (N_43001,N_41281,N_41671);
xnor U43002 (N_43002,N_41244,N_41486);
or U43003 (N_43003,N_40832,N_41175);
nand U43004 (N_43004,N_41236,N_41192);
xor U43005 (N_43005,N_41606,N_41840);
xor U43006 (N_43006,N_40401,N_40332);
or U43007 (N_43007,N_41442,N_41383);
nor U43008 (N_43008,N_40455,N_41906);
nor U43009 (N_43009,N_41198,N_40357);
xor U43010 (N_43010,N_41259,N_40417);
xor U43011 (N_43011,N_41039,N_41790);
and U43012 (N_43012,N_41350,N_40669);
or U43013 (N_43013,N_41702,N_40304);
xnor U43014 (N_43014,N_40472,N_41307);
and U43015 (N_43015,N_40687,N_40545);
nor U43016 (N_43016,N_40122,N_40192);
or U43017 (N_43017,N_41094,N_41037);
and U43018 (N_43018,N_41071,N_40775);
xnor U43019 (N_43019,N_40258,N_41814);
xor U43020 (N_43020,N_40347,N_40061);
nor U43021 (N_43021,N_41966,N_41184);
or U43022 (N_43022,N_40188,N_41198);
or U43023 (N_43023,N_40841,N_41619);
and U43024 (N_43024,N_41021,N_40355);
or U43025 (N_43025,N_40207,N_41583);
nor U43026 (N_43026,N_41842,N_41570);
nor U43027 (N_43027,N_41167,N_41058);
or U43028 (N_43028,N_41281,N_41646);
or U43029 (N_43029,N_41241,N_41682);
or U43030 (N_43030,N_41456,N_40231);
nor U43031 (N_43031,N_40267,N_40501);
nand U43032 (N_43032,N_40474,N_40214);
or U43033 (N_43033,N_41993,N_40069);
nor U43034 (N_43034,N_41994,N_40165);
and U43035 (N_43035,N_40977,N_40939);
and U43036 (N_43036,N_40451,N_41369);
or U43037 (N_43037,N_41996,N_40610);
nor U43038 (N_43038,N_41324,N_40684);
nand U43039 (N_43039,N_40457,N_40298);
nand U43040 (N_43040,N_40124,N_41567);
xnor U43041 (N_43041,N_40397,N_40699);
and U43042 (N_43042,N_40173,N_41384);
nor U43043 (N_43043,N_40203,N_40398);
nor U43044 (N_43044,N_40835,N_40268);
or U43045 (N_43045,N_40321,N_40309);
nand U43046 (N_43046,N_40315,N_40523);
xnor U43047 (N_43047,N_40054,N_40352);
and U43048 (N_43048,N_41407,N_41235);
or U43049 (N_43049,N_41101,N_40726);
and U43050 (N_43050,N_40961,N_41844);
xor U43051 (N_43051,N_40211,N_40370);
or U43052 (N_43052,N_41000,N_41529);
and U43053 (N_43053,N_40763,N_41240);
nand U43054 (N_43054,N_41509,N_41700);
and U43055 (N_43055,N_40991,N_40036);
xor U43056 (N_43056,N_40829,N_40508);
xnor U43057 (N_43057,N_40698,N_41185);
or U43058 (N_43058,N_40871,N_41213);
nand U43059 (N_43059,N_41295,N_40081);
or U43060 (N_43060,N_40181,N_41382);
and U43061 (N_43061,N_40014,N_41809);
and U43062 (N_43062,N_41604,N_40769);
xnor U43063 (N_43063,N_41966,N_41475);
nor U43064 (N_43064,N_41714,N_40720);
and U43065 (N_43065,N_40817,N_40298);
xor U43066 (N_43066,N_40900,N_41903);
nor U43067 (N_43067,N_41751,N_40824);
or U43068 (N_43068,N_40052,N_41684);
xnor U43069 (N_43069,N_40918,N_41925);
nand U43070 (N_43070,N_40557,N_41568);
xor U43071 (N_43071,N_41757,N_41079);
or U43072 (N_43072,N_41818,N_41812);
nand U43073 (N_43073,N_40335,N_40935);
xnor U43074 (N_43074,N_40904,N_41357);
or U43075 (N_43075,N_40287,N_41333);
or U43076 (N_43076,N_41356,N_41600);
or U43077 (N_43077,N_40139,N_40048);
or U43078 (N_43078,N_40891,N_40487);
and U43079 (N_43079,N_41740,N_41696);
xnor U43080 (N_43080,N_40621,N_40061);
xnor U43081 (N_43081,N_40887,N_40831);
nor U43082 (N_43082,N_41745,N_41343);
xor U43083 (N_43083,N_41275,N_41839);
nor U43084 (N_43084,N_40304,N_40839);
or U43085 (N_43085,N_41021,N_40416);
xor U43086 (N_43086,N_41191,N_41629);
nor U43087 (N_43087,N_41727,N_40235);
nand U43088 (N_43088,N_41605,N_40175);
nand U43089 (N_43089,N_40276,N_41707);
nand U43090 (N_43090,N_41796,N_41414);
xnor U43091 (N_43091,N_40507,N_40408);
xor U43092 (N_43092,N_40933,N_40144);
or U43093 (N_43093,N_41849,N_40011);
nor U43094 (N_43094,N_40031,N_41789);
nand U43095 (N_43095,N_40748,N_40000);
nor U43096 (N_43096,N_41831,N_40954);
nor U43097 (N_43097,N_40940,N_41686);
or U43098 (N_43098,N_41747,N_41428);
nor U43099 (N_43099,N_40238,N_41213);
and U43100 (N_43100,N_40930,N_40664);
nand U43101 (N_43101,N_40249,N_41736);
nor U43102 (N_43102,N_41590,N_40123);
or U43103 (N_43103,N_41548,N_40772);
nand U43104 (N_43104,N_40134,N_40876);
and U43105 (N_43105,N_41097,N_41654);
nor U43106 (N_43106,N_40589,N_40411);
nand U43107 (N_43107,N_40565,N_40973);
xor U43108 (N_43108,N_41052,N_40109);
nor U43109 (N_43109,N_40548,N_40366);
and U43110 (N_43110,N_41616,N_41537);
nor U43111 (N_43111,N_40466,N_41542);
and U43112 (N_43112,N_41622,N_41569);
and U43113 (N_43113,N_40040,N_41826);
and U43114 (N_43114,N_41808,N_40982);
nand U43115 (N_43115,N_41361,N_41002);
xor U43116 (N_43116,N_41114,N_40973);
nor U43117 (N_43117,N_40080,N_41871);
or U43118 (N_43118,N_40815,N_41520);
or U43119 (N_43119,N_40368,N_41553);
and U43120 (N_43120,N_41804,N_41793);
nor U43121 (N_43121,N_40545,N_41537);
xnor U43122 (N_43122,N_40499,N_40096);
and U43123 (N_43123,N_41918,N_40330);
or U43124 (N_43124,N_40010,N_41162);
or U43125 (N_43125,N_41144,N_41951);
nor U43126 (N_43126,N_40412,N_41882);
or U43127 (N_43127,N_40534,N_41048);
or U43128 (N_43128,N_40802,N_40108);
and U43129 (N_43129,N_41186,N_40277);
nand U43130 (N_43130,N_41656,N_40649);
nand U43131 (N_43131,N_41522,N_41816);
and U43132 (N_43132,N_40164,N_41281);
and U43133 (N_43133,N_41018,N_41355);
and U43134 (N_43134,N_40674,N_41811);
nand U43135 (N_43135,N_41174,N_40002);
or U43136 (N_43136,N_40768,N_41361);
or U43137 (N_43137,N_41170,N_41502);
or U43138 (N_43138,N_40462,N_41387);
or U43139 (N_43139,N_41287,N_40605);
or U43140 (N_43140,N_40955,N_41964);
and U43141 (N_43141,N_41220,N_41940);
nor U43142 (N_43142,N_41938,N_40655);
and U43143 (N_43143,N_41328,N_41127);
nand U43144 (N_43144,N_41002,N_40445);
and U43145 (N_43145,N_41065,N_40888);
nand U43146 (N_43146,N_40208,N_40051);
nand U43147 (N_43147,N_40497,N_41637);
xnor U43148 (N_43148,N_41733,N_41667);
and U43149 (N_43149,N_40021,N_40990);
xor U43150 (N_43150,N_40469,N_41103);
and U43151 (N_43151,N_41465,N_40010);
nand U43152 (N_43152,N_40825,N_40210);
and U43153 (N_43153,N_41430,N_41535);
xor U43154 (N_43154,N_41465,N_40024);
and U43155 (N_43155,N_40629,N_40635);
xor U43156 (N_43156,N_41197,N_40263);
or U43157 (N_43157,N_40037,N_40096);
or U43158 (N_43158,N_40493,N_41464);
xnor U43159 (N_43159,N_41239,N_41480);
nand U43160 (N_43160,N_41364,N_40750);
nand U43161 (N_43161,N_41388,N_41065);
xor U43162 (N_43162,N_40073,N_40584);
nand U43163 (N_43163,N_40332,N_41584);
nor U43164 (N_43164,N_41161,N_41829);
nand U43165 (N_43165,N_40187,N_40976);
xnor U43166 (N_43166,N_41757,N_40491);
nor U43167 (N_43167,N_41635,N_40896);
or U43168 (N_43168,N_41643,N_40572);
xor U43169 (N_43169,N_40117,N_41578);
and U43170 (N_43170,N_40508,N_40236);
xor U43171 (N_43171,N_41512,N_40416);
nand U43172 (N_43172,N_40463,N_40586);
nand U43173 (N_43173,N_40110,N_41481);
nand U43174 (N_43174,N_40622,N_41297);
or U43175 (N_43175,N_40194,N_40178);
nand U43176 (N_43176,N_41912,N_41059);
nand U43177 (N_43177,N_40226,N_40396);
xor U43178 (N_43178,N_40163,N_40463);
xnor U43179 (N_43179,N_41446,N_41861);
nor U43180 (N_43180,N_41913,N_41483);
or U43181 (N_43181,N_40397,N_40212);
nor U43182 (N_43182,N_41659,N_41308);
xnor U43183 (N_43183,N_41726,N_41606);
and U43184 (N_43184,N_40705,N_41640);
xnor U43185 (N_43185,N_41792,N_41499);
nor U43186 (N_43186,N_40927,N_41788);
nand U43187 (N_43187,N_40882,N_41648);
nor U43188 (N_43188,N_40153,N_40097);
and U43189 (N_43189,N_40755,N_40657);
and U43190 (N_43190,N_40532,N_40871);
xor U43191 (N_43191,N_40618,N_41391);
nor U43192 (N_43192,N_40499,N_40358);
or U43193 (N_43193,N_41292,N_40577);
xnor U43194 (N_43194,N_40761,N_41227);
or U43195 (N_43195,N_41514,N_40480);
xnor U43196 (N_43196,N_41236,N_40913);
and U43197 (N_43197,N_40817,N_41469);
nor U43198 (N_43198,N_41838,N_41340);
nand U43199 (N_43199,N_40363,N_41105);
nor U43200 (N_43200,N_40859,N_40909);
nor U43201 (N_43201,N_40234,N_40043);
xnor U43202 (N_43202,N_41059,N_40296);
xnor U43203 (N_43203,N_41506,N_41784);
xnor U43204 (N_43204,N_40918,N_40008);
nor U43205 (N_43205,N_40158,N_40026);
and U43206 (N_43206,N_40239,N_41697);
nor U43207 (N_43207,N_41650,N_40688);
xor U43208 (N_43208,N_41892,N_41967);
nand U43209 (N_43209,N_40913,N_41906);
xor U43210 (N_43210,N_40746,N_41261);
and U43211 (N_43211,N_41843,N_40752);
nor U43212 (N_43212,N_41395,N_41287);
or U43213 (N_43213,N_40680,N_40727);
nor U43214 (N_43214,N_40477,N_41204);
nor U43215 (N_43215,N_41029,N_40533);
and U43216 (N_43216,N_41923,N_41758);
and U43217 (N_43217,N_40214,N_41084);
and U43218 (N_43218,N_40814,N_40017);
nand U43219 (N_43219,N_41491,N_41142);
nor U43220 (N_43220,N_40388,N_40242);
xnor U43221 (N_43221,N_41472,N_41217);
and U43222 (N_43222,N_41295,N_40608);
or U43223 (N_43223,N_41683,N_41789);
nor U43224 (N_43224,N_40944,N_41927);
xnor U43225 (N_43225,N_41369,N_41950);
nor U43226 (N_43226,N_41235,N_41318);
and U43227 (N_43227,N_40941,N_41580);
or U43228 (N_43228,N_41027,N_40908);
nand U43229 (N_43229,N_40965,N_41367);
nor U43230 (N_43230,N_40158,N_40910);
nand U43231 (N_43231,N_41623,N_41796);
or U43232 (N_43232,N_41259,N_40580);
nor U43233 (N_43233,N_41277,N_40367);
or U43234 (N_43234,N_40698,N_41772);
and U43235 (N_43235,N_41583,N_40996);
nor U43236 (N_43236,N_41961,N_40297);
nand U43237 (N_43237,N_40276,N_41052);
xnor U43238 (N_43238,N_41786,N_41886);
and U43239 (N_43239,N_40735,N_40075);
xor U43240 (N_43240,N_40612,N_40481);
xor U43241 (N_43241,N_41381,N_40373);
or U43242 (N_43242,N_40215,N_41391);
nor U43243 (N_43243,N_41318,N_41760);
or U43244 (N_43244,N_40912,N_40935);
or U43245 (N_43245,N_40910,N_40692);
nor U43246 (N_43246,N_41033,N_40932);
xor U43247 (N_43247,N_40485,N_41480);
nand U43248 (N_43248,N_40663,N_41237);
and U43249 (N_43249,N_41427,N_40170);
nand U43250 (N_43250,N_41725,N_41866);
nor U43251 (N_43251,N_40968,N_40204);
and U43252 (N_43252,N_40343,N_40516);
or U43253 (N_43253,N_40658,N_40842);
nor U43254 (N_43254,N_41385,N_40767);
nand U43255 (N_43255,N_41696,N_41678);
or U43256 (N_43256,N_40246,N_41221);
and U43257 (N_43257,N_41974,N_40833);
and U43258 (N_43258,N_41896,N_41774);
xor U43259 (N_43259,N_41235,N_41642);
xnor U43260 (N_43260,N_40731,N_41576);
xnor U43261 (N_43261,N_40539,N_40917);
nor U43262 (N_43262,N_41110,N_40934);
xor U43263 (N_43263,N_40421,N_41983);
nand U43264 (N_43264,N_41504,N_41383);
and U43265 (N_43265,N_40547,N_41492);
or U43266 (N_43266,N_40137,N_40663);
or U43267 (N_43267,N_40286,N_40926);
nor U43268 (N_43268,N_40021,N_40244);
nor U43269 (N_43269,N_41076,N_41390);
and U43270 (N_43270,N_41903,N_40608);
nand U43271 (N_43271,N_40065,N_41429);
xnor U43272 (N_43272,N_41338,N_40355);
or U43273 (N_43273,N_41803,N_40904);
and U43274 (N_43274,N_41378,N_40409);
nand U43275 (N_43275,N_41863,N_41416);
xnor U43276 (N_43276,N_41494,N_41810);
nand U43277 (N_43277,N_40246,N_41536);
and U43278 (N_43278,N_40177,N_40541);
and U43279 (N_43279,N_40096,N_40131);
xor U43280 (N_43280,N_40936,N_40186);
and U43281 (N_43281,N_40353,N_41374);
nand U43282 (N_43282,N_41395,N_41612);
xnor U43283 (N_43283,N_40905,N_40221);
nand U43284 (N_43284,N_40362,N_40382);
or U43285 (N_43285,N_40006,N_40345);
xor U43286 (N_43286,N_41415,N_41910);
xnor U43287 (N_43287,N_40016,N_41382);
xor U43288 (N_43288,N_41226,N_40634);
xnor U43289 (N_43289,N_40390,N_41449);
nor U43290 (N_43290,N_41873,N_41676);
xnor U43291 (N_43291,N_41315,N_40900);
nor U43292 (N_43292,N_41884,N_40442);
nor U43293 (N_43293,N_41156,N_41434);
xor U43294 (N_43294,N_41320,N_41697);
nand U43295 (N_43295,N_40572,N_40722);
or U43296 (N_43296,N_41565,N_40201);
nor U43297 (N_43297,N_40164,N_40362);
or U43298 (N_43298,N_40533,N_40613);
and U43299 (N_43299,N_41251,N_40068);
nand U43300 (N_43300,N_40743,N_40803);
nand U43301 (N_43301,N_40607,N_41952);
and U43302 (N_43302,N_40086,N_40448);
nand U43303 (N_43303,N_40985,N_40490);
nand U43304 (N_43304,N_40677,N_40129);
nand U43305 (N_43305,N_41075,N_41593);
nor U43306 (N_43306,N_41924,N_40752);
and U43307 (N_43307,N_40481,N_40949);
nand U43308 (N_43308,N_40930,N_41022);
nor U43309 (N_43309,N_41477,N_41487);
nor U43310 (N_43310,N_41912,N_40012);
nor U43311 (N_43311,N_40684,N_40304);
nand U43312 (N_43312,N_40959,N_41686);
xor U43313 (N_43313,N_40005,N_41606);
xnor U43314 (N_43314,N_40169,N_41590);
or U43315 (N_43315,N_41505,N_41846);
nand U43316 (N_43316,N_40160,N_40455);
xnor U43317 (N_43317,N_40236,N_40790);
xor U43318 (N_43318,N_41298,N_40661);
and U43319 (N_43319,N_40384,N_40264);
nand U43320 (N_43320,N_41993,N_40591);
and U43321 (N_43321,N_40263,N_41279);
and U43322 (N_43322,N_40400,N_40799);
and U43323 (N_43323,N_41916,N_40601);
or U43324 (N_43324,N_41495,N_41485);
or U43325 (N_43325,N_40435,N_40930);
and U43326 (N_43326,N_40624,N_41530);
or U43327 (N_43327,N_40685,N_40781);
and U43328 (N_43328,N_40425,N_40177);
xor U43329 (N_43329,N_41151,N_41395);
and U43330 (N_43330,N_41059,N_40959);
nand U43331 (N_43331,N_40117,N_40041);
xnor U43332 (N_43332,N_40562,N_40897);
or U43333 (N_43333,N_41322,N_41238);
or U43334 (N_43334,N_41803,N_40932);
and U43335 (N_43335,N_41350,N_40505);
nor U43336 (N_43336,N_41612,N_40989);
nor U43337 (N_43337,N_41251,N_41348);
nor U43338 (N_43338,N_41977,N_41725);
and U43339 (N_43339,N_41735,N_41171);
nand U43340 (N_43340,N_41227,N_41872);
nand U43341 (N_43341,N_40061,N_41615);
or U43342 (N_43342,N_40043,N_41583);
nand U43343 (N_43343,N_41324,N_41034);
nor U43344 (N_43344,N_41440,N_40395);
nor U43345 (N_43345,N_40225,N_40891);
nand U43346 (N_43346,N_41446,N_41224);
and U43347 (N_43347,N_41206,N_41952);
and U43348 (N_43348,N_41063,N_41928);
and U43349 (N_43349,N_41244,N_41549);
or U43350 (N_43350,N_41939,N_40526);
or U43351 (N_43351,N_40338,N_41130);
nand U43352 (N_43352,N_40526,N_40894);
or U43353 (N_43353,N_40405,N_41458);
nor U43354 (N_43354,N_41969,N_40232);
xor U43355 (N_43355,N_40671,N_40705);
nand U43356 (N_43356,N_41943,N_41078);
nand U43357 (N_43357,N_40632,N_40440);
nand U43358 (N_43358,N_40093,N_41353);
nor U43359 (N_43359,N_40811,N_40206);
or U43360 (N_43360,N_40009,N_40624);
nor U43361 (N_43361,N_40051,N_41924);
or U43362 (N_43362,N_40654,N_41871);
nor U43363 (N_43363,N_40090,N_41522);
nand U43364 (N_43364,N_40352,N_40350);
and U43365 (N_43365,N_40649,N_41338);
and U43366 (N_43366,N_40521,N_41342);
nor U43367 (N_43367,N_40428,N_40280);
and U43368 (N_43368,N_41932,N_40291);
or U43369 (N_43369,N_41520,N_41971);
xnor U43370 (N_43370,N_40276,N_40507);
nand U43371 (N_43371,N_41073,N_40634);
nand U43372 (N_43372,N_41753,N_41650);
and U43373 (N_43373,N_40896,N_41022);
and U43374 (N_43374,N_41345,N_40830);
nand U43375 (N_43375,N_41204,N_40602);
or U43376 (N_43376,N_41174,N_40504);
xnor U43377 (N_43377,N_40572,N_41768);
xor U43378 (N_43378,N_40166,N_41610);
xor U43379 (N_43379,N_41833,N_41686);
or U43380 (N_43380,N_40472,N_40794);
and U43381 (N_43381,N_41811,N_41850);
or U43382 (N_43382,N_40602,N_41679);
xor U43383 (N_43383,N_40220,N_41766);
nor U43384 (N_43384,N_40469,N_41011);
or U43385 (N_43385,N_40493,N_40770);
and U43386 (N_43386,N_40655,N_40344);
nor U43387 (N_43387,N_40701,N_40568);
or U43388 (N_43388,N_41822,N_41884);
and U43389 (N_43389,N_41571,N_41510);
or U43390 (N_43390,N_40337,N_40214);
or U43391 (N_43391,N_40581,N_41416);
nor U43392 (N_43392,N_40150,N_41916);
nor U43393 (N_43393,N_40137,N_41473);
xor U43394 (N_43394,N_40604,N_40974);
nor U43395 (N_43395,N_41541,N_40883);
and U43396 (N_43396,N_40737,N_41249);
or U43397 (N_43397,N_41229,N_40031);
xor U43398 (N_43398,N_40263,N_40183);
xor U43399 (N_43399,N_41171,N_41384);
xor U43400 (N_43400,N_41932,N_40203);
and U43401 (N_43401,N_40875,N_40368);
or U43402 (N_43402,N_40410,N_41434);
xor U43403 (N_43403,N_40928,N_41718);
or U43404 (N_43404,N_41167,N_41006);
nand U43405 (N_43405,N_40042,N_40888);
and U43406 (N_43406,N_40904,N_41358);
nand U43407 (N_43407,N_40749,N_41547);
or U43408 (N_43408,N_40788,N_40177);
xnor U43409 (N_43409,N_40392,N_41005);
or U43410 (N_43410,N_40363,N_40094);
nand U43411 (N_43411,N_41694,N_41565);
xnor U43412 (N_43412,N_41966,N_41295);
nand U43413 (N_43413,N_40722,N_41988);
or U43414 (N_43414,N_40867,N_41587);
nand U43415 (N_43415,N_40194,N_41909);
and U43416 (N_43416,N_41881,N_41267);
nand U43417 (N_43417,N_41289,N_41342);
nand U43418 (N_43418,N_41008,N_41065);
or U43419 (N_43419,N_40938,N_41575);
and U43420 (N_43420,N_41513,N_40683);
nand U43421 (N_43421,N_41759,N_40765);
or U43422 (N_43422,N_40684,N_40806);
nand U43423 (N_43423,N_40764,N_40484);
or U43424 (N_43424,N_40353,N_41356);
nand U43425 (N_43425,N_41059,N_41154);
and U43426 (N_43426,N_41472,N_40762);
or U43427 (N_43427,N_40306,N_40683);
xnor U43428 (N_43428,N_40089,N_40070);
or U43429 (N_43429,N_41759,N_41424);
or U43430 (N_43430,N_41614,N_41604);
nor U43431 (N_43431,N_40401,N_40639);
and U43432 (N_43432,N_41051,N_40152);
nor U43433 (N_43433,N_41766,N_41466);
xnor U43434 (N_43434,N_41491,N_41821);
and U43435 (N_43435,N_41688,N_40195);
or U43436 (N_43436,N_41562,N_40599);
and U43437 (N_43437,N_40291,N_41459);
nor U43438 (N_43438,N_41520,N_40172);
xor U43439 (N_43439,N_40103,N_40638);
nand U43440 (N_43440,N_41653,N_40025);
nor U43441 (N_43441,N_41175,N_41711);
and U43442 (N_43442,N_40648,N_40252);
and U43443 (N_43443,N_41431,N_41415);
or U43444 (N_43444,N_41646,N_40020);
xnor U43445 (N_43445,N_41118,N_40188);
and U43446 (N_43446,N_41013,N_41396);
xnor U43447 (N_43447,N_40558,N_41036);
and U43448 (N_43448,N_40694,N_41023);
and U43449 (N_43449,N_40468,N_40543);
nand U43450 (N_43450,N_41340,N_41242);
xnor U43451 (N_43451,N_41069,N_41661);
and U43452 (N_43452,N_40757,N_40880);
and U43453 (N_43453,N_40326,N_41329);
nand U43454 (N_43454,N_41326,N_40421);
nor U43455 (N_43455,N_41958,N_40264);
nor U43456 (N_43456,N_40442,N_41835);
xor U43457 (N_43457,N_41190,N_41358);
xnor U43458 (N_43458,N_40501,N_40948);
xnor U43459 (N_43459,N_41905,N_41647);
nand U43460 (N_43460,N_40319,N_40876);
and U43461 (N_43461,N_40877,N_40899);
nand U43462 (N_43462,N_40569,N_41817);
and U43463 (N_43463,N_40485,N_41118);
and U43464 (N_43464,N_41791,N_41587);
nor U43465 (N_43465,N_40846,N_40329);
nand U43466 (N_43466,N_41950,N_40216);
nor U43467 (N_43467,N_41492,N_40821);
and U43468 (N_43468,N_41220,N_41890);
nand U43469 (N_43469,N_40834,N_41627);
nand U43470 (N_43470,N_41228,N_40229);
xor U43471 (N_43471,N_41437,N_40785);
and U43472 (N_43472,N_41056,N_40155);
or U43473 (N_43473,N_40067,N_40234);
nand U43474 (N_43474,N_40673,N_41578);
or U43475 (N_43475,N_41102,N_40043);
or U43476 (N_43476,N_40496,N_40323);
and U43477 (N_43477,N_41786,N_41870);
nor U43478 (N_43478,N_41043,N_40390);
xnor U43479 (N_43479,N_40781,N_40998);
xor U43480 (N_43480,N_41144,N_40604);
and U43481 (N_43481,N_41368,N_40465);
nand U43482 (N_43482,N_40249,N_41799);
or U43483 (N_43483,N_41597,N_40335);
and U43484 (N_43484,N_40394,N_40348);
nor U43485 (N_43485,N_41622,N_41611);
or U43486 (N_43486,N_40882,N_41452);
and U43487 (N_43487,N_40252,N_41406);
nor U43488 (N_43488,N_40645,N_40146);
xor U43489 (N_43489,N_40116,N_40062);
nor U43490 (N_43490,N_40383,N_40599);
and U43491 (N_43491,N_40638,N_41334);
or U43492 (N_43492,N_41445,N_40258);
xor U43493 (N_43493,N_40818,N_40978);
and U43494 (N_43494,N_40408,N_41119);
xor U43495 (N_43495,N_40226,N_40273);
and U43496 (N_43496,N_40838,N_41618);
nor U43497 (N_43497,N_41150,N_40837);
nand U43498 (N_43498,N_41445,N_40044);
nand U43499 (N_43499,N_41891,N_40108);
nor U43500 (N_43500,N_41532,N_41024);
xnor U43501 (N_43501,N_41318,N_40742);
or U43502 (N_43502,N_40948,N_40131);
xor U43503 (N_43503,N_40853,N_41298);
nand U43504 (N_43504,N_41340,N_40915);
xor U43505 (N_43505,N_41899,N_40698);
nand U43506 (N_43506,N_41139,N_40799);
and U43507 (N_43507,N_40978,N_41916);
nand U43508 (N_43508,N_40215,N_41331);
xnor U43509 (N_43509,N_41419,N_41271);
xnor U43510 (N_43510,N_40270,N_41528);
and U43511 (N_43511,N_40836,N_40934);
nand U43512 (N_43512,N_41208,N_41994);
and U43513 (N_43513,N_41264,N_40208);
or U43514 (N_43514,N_41232,N_40818);
nand U43515 (N_43515,N_40969,N_40971);
and U43516 (N_43516,N_41111,N_40190);
xor U43517 (N_43517,N_41628,N_41728);
nor U43518 (N_43518,N_41026,N_41025);
xor U43519 (N_43519,N_41637,N_40788);
and U43520 (N_43520,N_40485,N_40856);
and U43521 (N_43521,N_41673,N_41230);
nor U43522 (N_43522,N_40868,N_41171);
nor U43523 (N_43523,N_41789,N_41688);
nor U43524 (N_43524,N_41662,N_40161);
or U43525 (N_43525,N_41957,N_41921);
xnor U43526 (N_43526,N_41871,N_41386);
and U43527 (N_43527,N_40939,N_40794);
and U43528 (N_43528,N_40360,N_41325);
and U43529 (N_43529,N_40879,N_41433);
and U43530 (N_43530,N_41254,N_40327);
nor U43531 (N_43531,N_40587,N_40463);
xor U43532 (N_43532,N_41713,N_40544);
or U43533 (N_43533,N_41844,N_40100);
and U43534 (N_43534,N_40466,N_40444);
and U43535 (N_43535,N_41444,N_41730);
and U43536 (N_43536,N_41900,N_41239);
nand U43537 (N_43537,N_41558,N_40468);
nor U43538 (N_43538,N_40966,N_41832);
nand U43539 (N_43539,N_40853,N_41079);
or U43540 (N_43540,N_40423,N_41329);
xor U43541 (N_43541,N_40964,N_41069);
nor U43542 (N_43542,N_41661,N_41681);
or U43543 (N_43543,N_40298,N_41829);
or U43544 (N_43544,N_40015,N_40126);
nor U43545 (N_43545,N_41919,N_41637);
and U43546 (N_43546,N_40265,N_41745);
xnor U43547 (N_43547,N_41842,N_40831);
nor U43548 (N_43548,N_40333,N_41493);
xor U43549 (N_43549,N_40121,N_41292);
xor U43550 (N_43550,N_41242,N_41045);
or U43551 (N_43551,N_41294,N_41026);
xnor U43552 (N_43552,N_41282,N_41741);
or U43553 (N_43553,N_40265,N_40845);
and U43554 (N_43554,N_40379,N_41512);
or U43555 (N_43555,N_40519,N_40365);
nand U43556 (N_43556,N_41070,N_40169);
or U43557 (N_43557,N_41854,N_40993);
xnor U43558 (N_43558,N_41007,N_40103);
nor U43559 (N_43559,N_40854,N_41158);
and U43560 (N_43560,N_40865,N_40966);
and U43561 (N_43561,N_40329,N_41259);
or U43562 (N_43562,N_41062,N_41184);
nand U43563 (N_43563,N_40453,N_41821);
xor U43564 (N_43564,N_40530,N_41672);
nand U43565 (N_43565,N_40205,N_41020);
nand U43566 (N_43566,N_40142,N_40558);
nand U43567 (N_43567,N_41389,N_41224);
nor U43568 (N_43568,N_40997,N_41845);
or U43569 (N_43569,N_41482,N_40302);
xnor U43570 (N_43570,N_41409,N_41085);
or U43571 (N_43571,N_41245,N_40790);
or U43572 (N_43572,N_41745,N_40873);
or U43573 (N_43573,N_40201,N_40533);
and U43574 (N_43574,N_40407,N_41833);
xor U43575 (N_43575,N_40582,N_40587);
nor U43576 (N_43576,N_41559,N_40321);
xnor U43577 (N_43577,N_40825,N_40052);
or U43578 (N_43578,N_41409,N_40168);
or U43579 (N_43579,N_41138,N_41408);
xor U43580 (N_43580,N_41610,N_41239);
nor U43581 (N_43581,N_40263,N_40127);
nor U43582 (N_43582,N_41811,N_40177);
and U43583 (N_43583,N_40641,N_40424);
nand U43584 (N_43584,N_41473,N_41048);
xor U43585 (N_43585,N_40286,N_41572);
and U43586 (N_43586,N_40141,N_40401);
xor U43587 (N_43587,N_40779,N_41912);
and U43588 (N_43588,N_40688,N_41326);
nor U43589 (N_43589,N_41244,N_41001);
nand U43590 (N_43590,N_40806,N_40836);
xor U43591 (N_43591,N_41712,N_40385);
nand U43592 (N_43592,N_40484,N_40870);
nand U43593 (N_43593,N_40375,N_40120);
or U43594 (N_43594,N_41940,N_40974);
nand U43595 (N_43595,N_41143,N_41603);
nor U43596 (N_43596,N_41146,N_41021);
or U43597 (N_43597,N_40285,N_41616);
nor U43598 (N_43598,N_41365,N_40948);
xor U43599 (N_43599,N_40485,N_41731);
nor U43600 (N_43600,N_40548,N_41747);
or U43601 (N_43601,N_40993,N_41771);
nand U43602 (N_43602,N_41464,N_40213);
nor U43603 (N_43603,N_40132,N_40336);
or U43604 (N_43604,N_40084,N_40444);
and U43605 (N_43605,N_41487,N_41538);
or U43606 (N_43606,N_40324,N_41369);
nand U43607 (N_43607,N_40859,N_41452);
nand U43608 (N_43608,N_41487,N_41307);
nand U43609 (N_43609,N_40424,N_41987);
nor U43610 (N_43610,N_40280,N_41851);
xnor U43611 (N_43611,N_40072,N_40027);
nand U43612 (N_43612,N_41572,N_40930);
xnor U43613 (N_43613,N_40953,N_41589);
xnor U43614 (N_43614,N_40307,N_40038);
and U43615 (N_43615,N_40999,N_40978);
xor U43616 (N_43616,N_41653,N_40204);
and U43617 (N_43617,N_41621,N_41637);
nor U43618 (N_43618,N_41429,N_40821);
and U43619 (N_43619,N_41395,N_40824);
nand U43620 (N_43620,N_40761,N_41999);
and U43621 (N_43621,N_40820,N_40176);
xor U43622 (N_43622,N_40567,N_41520);
and U43623 (N_43623,N_40373,N_40622);
nand U43624 (N_43624,N_41451,N_41903);
xnor U43625 (N_43625,N_40269,N_41262);
or U43626 (N_43626,N_40666,N_40566);
or U43627 (N_43627,N_40721,N_40005);
nor U43628 (N_43628,N_41234,N_41635);
and U43629 (N_43629,N_41449,N_40328);
nand U43630 (N_43630,N_41429,N_41355);
and U43631 (N_43631,N_40371,N_40134);
or U43632 (N_43632,N_40498,N_41233);
and U43633 (N_43633,N_40001,N_41268);
nor U43634 (N_43634,N_41616,N_41356);
nor U43635 (N_43635,N_41752,N_40722);
or U43636 (N_43636,N_40858,N_40311);
xnor U43637 (N_43637,N_40501,N_41499);
nand U43638 (N_43638,N_41070,N_40859);
or U43639 (N_43639,N_40179,N_40140);
or U43640 (N_43640,N_41939,N_41235);
or U43641 (N_43641,N_41512,N_41596);
nand U43642 (N_43642,N_40353,N_40534);
nand U43643 (N_43643,N_40544,N_41937);
nor U43644 (N_43644,N_41726,N_40559);
or U43645 (N_43645,N_41773,N_40484);
xor U43646 (N_43646,N_40908,N_41825);
nor U43647 (N_43647,N_40507,N_41748);
and U43648 (N_43648,N_40498,N_40959);
or U43649 (N_43649,N_40546,N_41210);
nor U43650 (N_43650,N_41087,N_41353);
and U43651 (N_43651,N_40310,N_40017);
nand U43652 (N_43652,N_41642,N_40729);
xnor U43653 (N_43653,N_41017,N_41914);
nor U43654 (N_43654,N_40599,N_40921);
nor U43655 (N_43655,N_40869,N_40525);
nand U43656 (N_43656,N_41972,N_40961);
or U43657 (N_43657,N_40900,N_41714);
and U43658 (N_43658,N_40380,N_40665);
and U43659 (N_43659,N_40399,N_40007);
or U43660 (N_43660,N_41973,N_41732);
and U43661 (N_43661,N_40294,N_40045);
xor U43662 (N_43662,N_41826,N_40245);
nor U43663 (N_43663,N_40130,N_41898);
nor U43664 (N_43664,N_41348,N_40654);
nand U43665 (N_43665,N_40176,N_41674);
and U43666 (N_43666,N_40446,N_40055);
nor U43667 (N_43667,N_41566,N_40670);
or U43668 (N_43668,N_41588,N_40499);
nor U43669 (N_43669,N_41394,N_40571);
nand U43670 (N_43670,N_40873,N_41934);
and U43671 (N_43671,N_41553,N_41987);
nor U43672 (N_43672,N_40677,N_41441);
and U43673 (N_43673,N_41832,N_40294);
nor U43674 (N_43674,N_41011,N_41619);
xnor U43675 (N_43675,N_40967,N_41858);
nand U43676 (N_43676,N_41433,N_40098);
xnor U43677 (N_43677,N_40889,N_41078);
xor U43678 (N_43678,N_41463,N_41231);
nor U43679 (N_43679,N_41370,N_41433);
and U43680 (N_43680,N_40126,N_40345);
nor U43681 (N_43681,N_40611,N_40895);
and U43682 (N_43682,N_41994,N_41902);
or U43683 (N_43683,N_41483,N_40549);
xor U43684 (N_43684,N_40480,N_41399);
or U43685 (N_43685,N_40080,N_40188);
nor U43686 (N_43686,N_40591,N_40668);
and U43687 (N_43687,N_40031,N_41952);
and U43688 (N_43688,N_41111,N_41951);
xor U43689 (N_43689,N_40105,N_40968);
nor U43690 (N_43690,N_40714,N_40751);
xnor U43691 (N_43691,N_40937,N_40218);
xnor U43692 (N_43692,N_40454,N_40202);
nor U43693 (N_43693,N_41843,N_41925);
and U43694 (N_43694,N_41660,N_41381);
or U43695 (N_43695,N_41974,N_40764);
xor U43696 (N_43696,N_40901,N_40025);
and U43697 (N_43697,N_41477,N_41250);
xor U43698 (N_43698,N_41815,N_41190);
xnor U43699 (N_43699,N_40448,N_40506);
nor U43700 (N_43700,N_41015,N_41872);
nor U43701 (N_43701,N_40736,N_40382);
and U43702 (N_43702,N_40420,N_40387);
and U43703 (N_43703,N_41791,N_40195);
nor U43704 (N_43704,N_40600,N_40548);
xnor U43705 (N_43705,N_40274,N_41842);
nor U43706 (N_43706,N_40525,N_41828);
nor U43707 (N_43707,N_41752,N_40621);
xnor U43708 (N_43708,N_41326,N_40138);
xor U43709 (N_43709,N_40610,N_40912);
xor U43710 (N_43710,N_40161,N_40603);
xor U43711 (N_43711,N_40752,N_41356);
nand U43712 (N_43712,N_40870,N_40982);
nor U43713 (N_43713,N_40084,N_41751);
or U43714 (N_43714,N_41603,N_41068);
nand U43715 (N_43715,N_40509,N_41238);
or U43716 (N_43716,N_41447,N_41763);
and U43717 (N_43717,N_40107,N_41933);
or U43718 (N_43718,N_40106,N_40407);
or U43719 (N_43719,N_41180,N_41857);
xor U43720 (N_43720,N_41327,N_40661);
nand U43721 (N_43721,N_41924,N_40034);
and U43722 (N_43722,N_40317,N_41580);
and U43723 (N_43723,N_41576,N_41274);
xor U43724 (N_43724,N_41124,N_40540);
or U43725 (N_43725,N_41990,N_41481);
nand U43726 (N_43726,N_41942,N_40804);
xnor U43727 (N_43727,N_40936,N_41964);
and U43728 (N_43728,N_40417,N_40138);
nor U43729 (N_43729,N_41789,N_40670);
xor U43730 (N_43730,N_40801,N_40313);
and U43731 (N_43731,N_41708,N_41995);
nor U43732 (N_43732,N_40490,N_41452);
or U43733 (N_43733,N_40681,N_40354);
or U43734 (N_43734,N_40774,N_40293);
and U43735 (N_43735,N_41126,N_40143);
nor U43736 (N_43736,N_40021,N_41431);
xnor U43737 (N_43737,N_40001,N_40418);
and U43738 (N_43738,N_40004,N_40619);
nand U43739 (N_43739,N_41481,N_41321);
or U43740 (N_43740,N_40270,N_40621);
and U43741 (N_43741,N_41131,N_41591);
xor U43742 (N_43742,N_40500,N_41724);
and U43743 (N_43743,N_40969,N_40133);
or U43744 (N_43744,N_41787,N_41066);
nor U43745 (N_43745,N_40065,N_41556);
or U43746 (N_43746,N_41838,N_40216);
and U43747 (N_43747,N_41168,N_40344);
and U43748 (N_43748,N_41733,N_40485);
xor U43749 (N_43749,N_40726,N_41448);
nor U43750 (N_43750,N_41970,N_41571);
or U43751 (N_43751,N_41191,N_40539);
xnor U43752 (N_43752,N_41571,N_41665);
or U43753 (N_43753,N_40382,N_41965);
and U43754 (N_43754,N_41633,N_40281);
or U43755 (N_43755,N_41713,N_41669);
xnor U43756 (N_43756,N_41758,N_41232);
or U43757 (N_43757,N_41758,N_41180);
and U43758 (N_43758,N_41598,N_40461);
nand U43759 (N_43759,N_40096,N_41172);
xor U43760 (N_43760,N_41173,N_40765);
or U43761 (N_43761,N_41816,N_40300);
nor U43762 (N_43762,N_40743,N_40691);
and U43763 (N_43763,N_41608,N_41738);
nor U43764 (N_43764,N_41650,N_41992);
nor U43765 (N_43765,N_41671,N_41576);
nor U43766 (N_43766,N_40186,N_40469);
nor U43767 (N_43767,N_41848,N_40863);
and U43768 (N_43768,N_40921,N_40496);
or U43769 (N_43769,N_41982,N_41996);
xnor U43770 (N_43770,N_40600,N_41059);
xor U43771 (N_43771,N_40854,N_40071);
xor U43772 (N_43772,N_40805,N_41878);
nand U43773 (N_43773,N_40445,N_40865);
and U43774 (N_43774,N_40817,N_41545);
nor U43775 (N_43775,N_41097,N_40996);
or U43776 (N_43776,N_40651,N_41436);
xnor U43777 (N_43777,N_40620,N_40121);
or U43778 (N_43778,N_41638,N_41653);
xor U43779 (N_43779,N_41642,N_40011);
nand U43780 (N_43780,N_41320,N_41297);
and U43781 (N_43781,N_40961,N_40812);
xnor U43782 (N_43782,N_41391,N_41723);
nor U43783 (N_43783,N_40915,N_40225);
and U43784 (N_43784,N_41156,N_41418);
and U43785 (N_43785,N_41654,N_40302);
and U43786 (N_43786,N_41395,N_40059);
nor U43787 (N_43787,N_40725,N_40427);
nand U43788 (N_43788,N_41797,N_41544);
nand U43789 (N_43789,N_41563,N_40194);
and U43790 (N_43790,N_41298,N_41599);
nand U43791 (N_43791,N_40590,N_40057);
and U43792 (N_43792,N_40947,N_41278);
xor U43793 (N_43793,N_40991,N_40587);
nor U43794 (N_43794,N_41906,N_40662);
nand U43795 (N_43795,N_40572,N_41616);
and U43796 (N_43796,N_41208,N_41126);
nand U43797 (N_43797,N_41341,N_40656);
and U43798 (N_43798,N_41675,N_41770);
and U43799 (N_43799,N_41967,N_41545);
or U43800 (N_43800,N_40057,N_41536);
or U43801 (N_43801,N_40645,N_41724);
xor U43802 (N_43802,N_40876,N_41953);
or U43803 (N_43803,N_41151,N_40860);
nor U43804 (N_43804,N_41286,N_40064);
and U43805 (N_43805,N_40607,N_41402);
and U43806 (N_43806,N_40499,N_40032);
nor U43807 (N_43807,N_41175,N_40248);
nor U43808 (N_43808,N_41822,N_40439);
nand U43809 (N_43809,N_40236,N_41384);
nand U43810 (N_43810,N_40370,N_41584);
and U43811 (N_43811,N_40814,N_40347);
nand U43812 (N_43812,N_40601,N_41891);
nand U43813 (N_43813,N_40689,N_40358);
nand U43814 (N_43814,N_40217,N_41149);
xnor U43815 (N_43815,N_41116,N_41622);
nor U43816 (N_43816,N_41392,N_41754);
nor U43817 (N_43817,N_40414,N_41884);
xor U43818 (N_43818,N_40144,N_40563);
xor U43819 (N_43819,N_40504,N_41474);
and U43820 (N_43820,N_41746,N_40715);
nand U43821 (N_43821,N_41917,N_40489);
xor U43822 (N_43822,N_41026,N_41411);
and U43823 (N_43823,N_41493,N_40424);
and U43824 (N_43824,N_40861,N_40109);
nand U43825 (N_43825,N_41059,N_40672);
nor U43826 (N_43826,N_40962,N_41834);
nand U43827 (N_43827,N_40140,N_40402);
and U43828 (N_43828,N_41487,N_41016);
nor U43829 (N_43829,N_40614,N_40712);
or U43830 (N_43830,N_41038,N_40729);
or U43831 (N_43831,N_40852,N_41681);
nor U43832 (N_43832,N_40016,N_41066);
nor U43833 (N_43833,N_40915,N_40440);
and U43834 (N_43834,N_40560,N_40503);
nor U43835 (N_43835,N_41292,N_40920);
nand U43836 (N_43836,N_40837,N_40579);
nand U43837 (N_43837,N_41556,N_41543);
or U43838 (N_43838,N_40552,N_41345);
and U43839 (N_43839,N_41400,N_40537);
nor U43840 (N_43840,N_41004,N_40857);
nor U43841 (N_43841,N_41354,N_41637);
xnor U43842 (N_43842,N_40173,N_41397);
xnor U43843 (N_43843,N_41339,N_40710);
xnor U43844 (N_43844,N_40436,N_40502);
xor U43845 (N_43845,N_41298,N_40257);
nand U43846 (N_43846,N_40929,N_41824);
xor U43847 (N_43847,N_41891,N_40525);
xnor U43848 (N_43848,N_40907,N_41406);
nand U43849 (N_43849,N_41614,N_40389);
and U43850 (N_43850,N_41883,N_40254);
nor U43851 (N_43851,N_40139,N_40734);
nand U43852 (N_43852,N_41983,N_41447);
or U43853 (N_43853,N_41927,N_41884);
nor U43854 (N_43854,N_41686,N_40310);
xnor U43855 (N_43855,N_40869,N_41352);
and U43856 (N_43856,N_40146,N_41452);
and U43857 (N_43857,N_40605,N_40339);
xnor U43858 (N_43858,N_40521,N_40737);
and U43859 (N_43859,N_41342,N_40945);
or U43860 (N_43860,N_40028,N_41293);
and U43861 (N_43861,N_41639,N_40735);
or U43862 (N_43862,N_40541,N_41901);
xor U43863 (N_43863,N_41491,N_40674);
nand U43864 (N_43864,N_41092,N_40884);
or U43865 (N_43865,N_40256,N_40600);
or U43866 (N_43866,N_41805,N_40849);
or U43867 (N_43867,N_40954,N_41183);
or U43868 (N_43868,N_40006,N_40670);
nor U43869 (N_43869,N_41936,N_41395);
xor U43870 (N_43870,N_40181,N_41208);
xor U43871 (N_43871,N_40077,N_41287);
or U43872 (N_43872,N_40714,N_40627);
or U43873 (N_43873,N_40504,N_40814);
xnor U43874 (N_43874,N_41280,N_41797);
xor U43875 (N_43875,N_40006,N_40867);
nand U43876 (N_43876,N_41564,N_40899);
xor U43877 (N_43877,N_41226,N_40588);
nand U43878 (N_43878,N_41804,N_40096);
nor U43879 (N_43879,N_40117,N_40003);
nand U43880 (N_43880,N_41709,N_40790);
nor U43881 (N_43881,N_41039,N_41956);
and U43882 (N_43882,N_41703,N_40832);
or U43883 (N_43883,N_40477,N_41389);
nor U43884 (N_43884,N_41475,N_41247);
nor U43885 (N_43885,N_41309,N_40935);
and U43886 (N_43886,N_41072,N_41687);
nor U43887 (N_43887,N_40481,N_41052);
nor U43888 (N_43888,N_41671,N_40034);
or U43889 (N_43889,N_40962,N_40989);
nor U43890 (N_43890,N_40462,N_40821);
xor U43891 (N_43891,N_41991,N_41406);
and U43892 (N_43892,N_40986,N_40264);
xor U43893 (N_43893,N_40801,N_41680);
or U43894 (N_43894,N_41079,N_41781);
or U43895 (N_43895,N_40828,N_40058);
xor U43896 (N_43896,N_40008,N_40311);
nor U43897 (N_43897,N_40529,N_40823);
and U43898 (N_43898,N_41893,N_40676);
or U43899 (N_43899,N_40669,N_40029);
and U43900 (N_43900,N_41771,N_40411);
or U43901 (N_43901,N_40477,N_40048);
and U43902 (N_43902,N_41673,N_40102);
xnor U43903 (N_43903,N_40688,N_40432);
and U43904 (N_43904,N_40263,N_40094);
xor U43905 (N_43905,N_41934,N_41424);
nor U43906 (N_43906,N_41758,N_40880);
or U43907 (N_43907,N_41449,N_40109);
xor U43908 (N_43908,N_40320,N_41386);
xor U43909 (N_43909,N_41600,N_41545);
xor U43910 (N_43910,N_41934,N_40821);
xnor U43911 (N_43911,N_40491,N_41721);
or U43912 (N_43912,N_41112,N_41488);
xnor U43913 (N_43913,N_41293,N_41960);
xor U43914 (N_43914,N_41070,N_41832);
nor U43915 (N_43915,N_40776,N_41936);
xor U43916 (N_43916,N_41083,N_40381);
and U43917 (N_43917,N_41171,N_40273);
and U43918 (N_43918,N_41661,N_40397);
and U43919 (N_43919,N_41527,N_41963);
and U43920 (N_43920,N_40816,N_41302);
and U43921 (N_43921,N_41634,N_41586);
xor U43922 (N_43922,N_41193,N_40640);
or U43923 (N_43923,N_41207,N_40161);
and U43924 (N_43924,N_41542,N_41722);
xnor U43925 (N_43925,N_40060,N_41638);
nor U43926 (N_43926,N_40947,N_40540);
or U43927 (N_43927,N_41767,N_41509);
nor U43928 (N_43928,N_41259,N_41036);
nand U43929 (N_43929,N_40677,N_40108);
nand U43930 (N_43930,N_40087,N_41010);
and U43931 (N_43931,N_41281,N_40743);
nand U43932 (N_43932,N_41329,N_40277);
xnor U43933 (N_43933,N_41115,N_40081);
nand U43934 (N_43934,N_41378,N_41578);
nand U43935 (N_43935,N_40054,N_40194);
xor U43936 (N_43936,N_40485,N_41385);
xnor U43937 (N_43937,N_40363,N_41379);
or U43938 (N_43938,N_41354,N_41963);
and U43939 (N_43939,N_40540,N_41518);
and U43940 (N_43940,N_41688,N_41399);
or U43941 (N_43941,N_40439,N_40885);
and U43942 (N_43942,N_40802,N_41669);
nor U43943 (N_43943,N_40858,N_41142);
xor U43944 (N_43944,N_40590,N_40187);
xnor U43945 (N_43945,N_40835,N_41740);
nand U43946 (N_43946,N_40967,N_41350);
xor U43947 (N_43947,N_41144,N_40160);
and U43948 (N_43948,N_41193,N_41276);
nor U43949 (N_43949,N_41474,N_40072);
or U43950 (N_43950,N_40255,N_40007);
nand U43951 (N_43951,N_41267,N_41730);
nor U43952 (N_43952,N_41974,N_41749);
and U43953 (N_43953,N_40510,N_40135);
and U43954 (N_43954,N_40615,N_41819);
or U43955 (N_43955,N_41338,N_40039);
and U43956 (N_43956,N_41737,N_40523);
or U43957 (N_43957,N_41804,N_41100);
xnor U43958 (N_43958,N_41777,N_41046);
and U43959 (N_43959,N_40742,N_40533);
nor U43960 (N_43960,N_41686,N_41500);
or U43961 (N_43961,N_41279,N_41618);
nand U43962 (N_43962,N_41506,N_40296);
xor U43963 (N_43963,N_40579,N_40278);
or U43964 (N_43964,N_41104,N_40589);
and U43965 (N_43965,N_40784,N_41336);
nor U43966 (N_43966,N_40777,N_41513);
nand U43967 (N_43967,N_40493,N_40916);
xnor U43968 (N_43968,N_41459,N_41801);
nor U43969 (N_43969,N_41017,N_40484);
or U43970 (N_43970,N_41857,N_40188);
or U43971 (N_43971,N_40894,N_40354);
or U43972 (N_43972,N_41172,N_40293);
nor U43973 (N_43973,N_40805,N_40505);
nor U43974 (N_43974,N_41579,N_40587);
nor U43975 (N_43975,N_40773,N_40077);
nor U43976 (N_43976,N_40861,N_41099);
nor U43977 (N_43977,N_41789,N_41182);
nor U43978 (N_43978,N_41167,N_41498);
and U43979 (N_43979,N_40530,N_40766);
nand U43980 (N_43980,N_41374,N_41607);
nand U43981 (N_43981,N_41580,N_40957);
or U43982 (N_43982,N_41856,N_40669);
nand U43983 (N_43983,N_40010,N_40902);
nand U43984 (N_43984,N_41216,N_41113);
xnor U43985 (N_43985,N_41120,N_41634);
xor U43986 (N_43986,N_40080,N_40874);
nand U43987 (N_43987,N_41953,N_41754);
xor U43988 (N_43988,N_40301,N_41408);
nor U43989 (N_43989,N_41707,N_40470);
and U43990 (N_43990,N_40264,N_41570);
xor U43991 (N_43991,N_40756,N_40138);
xor U43992 (N_43992,N_41879,N_40271);
nor U43993 (N_43993,N_41828,N_40723);
or U43994 (N_43994,N_41571,N_40948);
or U43995 (N_43995,N_40664,N_41112);
nor U43996 (N_43996,N_41629,N_40582);
and U43997 (N_43997,N_40283,N_41748);
nor U43998 (N_43998,N_41525,N_41436);
xnor U43999 (N_43999,N_41768,N_40193);
or U44000 (N_44000,N_42552,N_42930);
nor U44001 (N_44001,N_42408,N_42216);
and U44002 (N_44002,N_43293,N_43432);
and U44003 (N_44003,N_43831,N_42296);
or U44004 (N_44004,N_42993,N_42271);
and U44005 (N_44005,N_42331,N_42272);
or U44006 (N_44006,N_43077,N_42302);
and U44007 (N_44007,N_43693,N_43544);
xor U44008 (N_44008,N_42460,N_42193);
nor U44009 (N_44009,N_43346,N_43316);
nand U44010 (N_44010,N_42488,N_43951);
xnor U44011 (N_44011,N_42896,N_43015);
and U44012 (N_44012,N_43967,N_42194);
or U44013 (N_44013,N_42637,N_42045);
nand U44014 (N_44014,N_42595,N_43333);
or U44015 (N_44015,N_42487,N_43404);
or U44016 (N_44016,N_42075,N_42107);
nand U44017 (N_44017,N_43428,N_42779);
xor U44018 (N_44018,N_42529,N_43340);
nand U44019 (N_44019,N_43061,N_43002);
xnor U44020 (N_44020,N_42725,N_43983);
nand U44021 (N_44021,N_42961,N_43562);
xnor U44022 (N_44022,N_43781,N_43561);
nor U44023 (N_44023,N_42139,N_42617);
nand U44024 (N_44024,N_43052,N_43175);
and U44025 (N_44025,N_42692,N_42517);
nand U44026 (N_44026,N_43248,N_43878);
or U44027 (N_44027,N_42413,N_43185);
xnor U44028 (N_44028,N_42079,N_42124);
nor U44029 (N_44029,N_43296,N_43301);
nand U44030 (N_44030,N_43977,N_42866);
and U44031 (N_44031,N_42613,N_42132);
nand U44032 (N_44032,N_43552,N_42220);
xnor U44033 (N_44033,N_42979,N_42941);
nand U44034 (N_44034,N_43522,N_42059);
xnor U44035 (N_44035,N_42570,N_43226);
nor U44036 (N_44036,N_43940,N_42039);
xnor U44037 (N_44037,N_42023,N_43383);
or U44038 (N_44038,N_42818,N_42334);
nand U44039 (N_44039,N_42395,N_43076);
nand U44040 (N_44040,N_43926,N_42061);
or U44041 (N_44041,N_42910,N_42957);
or U44042 (N_44042,N_43919,N_43496);
nor U44043 (N_44043,N_42058,N_42428);
or U44044 (N_44044,N_43412,N_42577);
or U44045 (N_44045,N_43516,N_42750);
and U44046 (N_44046,N_42335,N_43583);
nand U44047 (N_44047,N_42849,N_43348);
nor U44048 (N_44048,N_42421,N_43643);
nand U44049 (N_44049,N_43551,N_42375);
or U44050 (N_44050,N_43176,N_42490);
nor U44051 (N_44051,N_42110,N_43987);
and U44052 (N_44052,N_42618,N_43311);
and U44053 (N_44053,N_42855,N_42596);
nand U44054 (N_44054,N_43267,N_43514);
nand U44055 (N_44055,N_43427,N_42018);
nor U44056 (N_44056,N_42664,N_42677);
and U44057 (N_44057,N_42576,N_42820);
nor U44058 (N_44058,N_43986,N_43691);
nor U44059 (N_44059,N_43549,N_43250);
and U44060 (N_44060,N_42532,N_43897);
xnor U44061 (N_44061,N_43354,N_42877);
nand U44062 (N_44062,N_43230,N_43109);
nor U44063 (N_44063,N_43107,N_43893);
nand U44064 (N_44064,N_43793,N_43374);
nand U44065 (N_44065,N_43202,N_43669);
and U44066 (N_44066,N_43445,N_43692);
xnor U44067 (N_44067,N_42603,N_42537);
or U44068 (N_44068,N_42102,N_43082);
xor U44069 (N_44069,N_42417,N_43547);
or U44070 (N_44070,N_43658,N_43007);
nor U44071 (N_44071,N_42129,N_42682);
or U44072 (N_44072,N_43278,N_42323);
nor U44073 (N_44073,N_42287,N_43063);
nor U44074 (N_44074,N_43336,N_42906);
nand U44075 (N_44075,N_42815,N_42550);
nor U44076 (N_44076,N_42269,N_43116);
nand U44077 (N_44077,N_42890,N_43845);
xor U44078 (N_44078,N_42086,N_42869);
nand U44079 (N_44079,N_43212,N_43511);
and U44080 (N_44080,N_42624,N_43168);
xor U44081 (N_44081,N_42245,N_42306);
nor U44082 (N_44082,N_42733,N_42469);
nor U44083 (N_44083,N_43913,N_42142);
and U44084 (N_44084,N_42827,N_42717);
and U44085 (N_44085,N_43459,N_43513);
xnor U44086 (N_44086,N_43523,N_42859);
nor U44087 (N_44087,N_42505,N_42420);
nor U44088 (N_44088,N_42044,N_42557);
and U44089 (N_44089,N_43736,N_43995);
and U44090 (N_44090,N_43727,N_43553);
xor U44091 (N_44091,N_43679,N_43075);
or U44092 (N_44092,N_43169,N_42825);
or U44093 (N_44093,N_43671,N_43517);
xor U44094 (N_44094,N_43215,N_42527);
and U44095 (N_44095,N_42609,N_43638);
or U44096 (N_44096,N_42212,N_42981);
xnor U44097 (N_44097,N_43803,N_42011);
and U44098 (N_44098,N_42431,N_42034);
nand U44099 (N_44099,N_42486,N_43442);
nor U44100 (N_44100,N_42600,N_42708);
and U44101 (N_44101,N_42085,N_42580);
nor U44102 (N_44102,N_43053,N_43330);
xnor U44103 (N_44103,N_42461,N_42400);
xnor U44104 (N_44104,N_42837,N_42791);
nand U44105 (N_44105,N_42073,N_43028);
nand U44106 (N_44106,N_43471,N_42797);
nand U44107 (N_44107,N_43395,N_43603);
and U44108 (N_44108,N_42250,N_42703);
xor U44109 (N_44109,N_43120,N_42761);
nand U44110 (N_44110,N_43121,N_43635);
and U44111 (N_44111,N_43319,N_42242);
nand U44112 (N_44112,N_42756,N_42858);
and U44113 (N_44113,N_42160,N_43399);
nand U44114 (N_44114,N_42736,N_43582);
xnor U44115 (N_44115,N_42622,N_43214);
and U44116 (N_44116,N_43453,N_42716);
nor U44117 (N_44117,N_43304,N_42391);
nor U44118 (N_44118,N_42556,N_43473);
or U44119 (N_44119,N_43580,N_43096);
nor U44120 (N_44120,N_42084,N_42484);
xnor U44121 (N_44121,N_42027,N_43824);
nand U44122 (N_44122,N_43850,N_42824);
nand U44123 (N_44123,N_42265,N_43836);
and U44124 (N_44124,N_43686,N_42214);
nand U44125 (N_44125,N_43978,N_43078);
and U44126 (N_44126,N_42281,N_43555);
nand U44127 (N_44127,N_43481,N_42351);
or U44128 (N_44128,N_43159,N_42493);
xor U44129 (N_44129,N_43999,N_42597);
or U44130 (N_44130,N_42987,N_43402);
xor U44131 (N_44131,N_43435,N_43125);
nand U44132 (N_44132,N_42076,N_43280);
xor U44133 (N_44133,N_43859,N_42501);
and U44134 (N_44134,N_43773,N_42237);
or U44135 (N_44135,N_43541,N_42623);
nand U44136 (N_44136,N_42332,N_43943);
xor U44137 (N_44137,N_43767,N_42711);
and U44138 (N_44138,N_43675,N_43771);
and U44139 (N_44139,N_42933,N_43676);
or U44140 (N_44140,N_42659,N_43678);
nand U44141 (N_44141,N_42713,N_43759);
nand U44142 (N_44142,N_42872,N_42819);
or U44143 (N_44143,N_43191,N_42355);
and U44144 (N_44144,N_43567,N_43928);
nor U44145 (N_44145,N_43416,N_43937);
nand U44146 (N_44146,N_43801,N_43006);
and U44147 (N_44147,N_43495,N_43022);
and U44148 (N_44148,N_43408,N_43653);
nand U44149 (N_44149,N_43622,N_42346);
and U44150 (N_44150,N_43989,N_43313);
nand U44151 (N_44151,N_42328,N_43810);
nand U44152 (N_44152,N_42317,N_43600);
nand U44153 (N_44153,N_43840,N_43018);
and U44154 (N_44154,N_43560,N_43003);
and U44155 (N_44155,N_43477,N_43729);
xnor U44156 (N_44156,N_42738,N_43392);
and U44157 (N_44157,N_43982,N_42678);
and U44158 (N_44158,N_43659,N_43642);
nor U44159 (N_44159,N_43529,N_42052);
or U44160 (N_44160,N_43208,N_42513);
and U44161 (N_44161,N_43414,N_42902);
or U44162 (N_44162,N_43703,N_43135);
and U44163 (N_44163,N_43013,N_42908);
xnor U44164 (N_44164,N_43540,N_42412);
nand U44165 (N_44165,N_42706,N_42764);
xnor U44166 (N_44166,N_42316,N_42919);
nand U44167 (N_44167,N_43749,N_43229);
and U44168 (N_44168,N_43266,N_43757);
or U44169 (N_44169,N_42667,N_42546);
xor U44170 (N_44170,N_43525,N_42345);
nor U44171 (N_44171,N_42369,N_42122);
nand U44172 (N_44172,N_43420,N_42240);
or U44173 (N_44173,N_42186,N_42985);
nand U44174 (N_44174,N_42514,N_42439);
and U44175 (N_44175,N_43466,N_42012);
nand U44176 (N_44176,N_42868,N_43242);
nand U44177 (N_44177,N_42816,N_42275);
nand U44178 (N_44178,N_43032,N_43908);
and U44179 (N_44179,N_42581,N_43133);
and U44180 (N_44180,N_42781,N_42473);
nand U44181 (N_44181,N_42239,N_42326);
nand U44182 (N_44182,N_42367,N_42917);
nand U44183 (N_44183,N_43934,N_42862);
xor U44184 (N_44184,N_43772,N_43775);
nand U44185 (N_44185,N_42422,N_42679);
or U44186 (N_44186,N_42203,N_43487);
nor U44187 (N_44187,N_43876,N_42798);
nor U44188 (N_44188,N_43961,N_42019);
and U44189 (N_44189,N_42728,N_42904);
nand U44190 (N_44190,N_43699,N_43581);
nor U44191 (N_44191,N_42774,N_42080);
and U44192 (N_44192,N_42313,N_43426);
and U44193 (N_44193,N_43371,N_43456);
or U44194 (N_44194,N_43375,N_42632);
nand U44195 (N_44195,N_42699,N_43865);
and U44196 (N_44196,N_43539,N_42991);
nand U44197 (N_44197,N_43646,N_42766);
and U44198 (N_44198,N_43656,N_43050);
or U44199 (N_44199,N_42481,N_42153);
nand U44200 (N_44200,N_42686,N_42893);
nand U44201 (N_44201,N_42530,N_42088);
and U44202 (N_44202,N_43964,N_42157);
or U44203 (N_44203,N_42494,N_42838);
nor U44204 (N_44204,N_43216,N_42378);
or U44205 (N_44205,N_42518,N_43283);
or U44206 (N_44206,N_42739,N_43722);
xnor U44207 (N_44207,N_42680,N_43388);
nor U44208 (N_44208,N_43751,N_42229);
or U44209 (N_44209,N_43180,N_43249);
or U44210 (N_44210,N_43049,N_43657);
nand U44211 (N_44211,N_43343,N_42318);
and U44212 (N_44212,N_42753,N_42333);
nor U44213 (N_44213,N_43766,N_43927);
or U44214 (N_44214,N_43485,N_43174);
nor U44215 (N_44215,N_42396,N_43713);
nor U44216 (N_44216,N_42655,N_42185);
xor U44217 (N_44217,N_43518,N_42471);
nor U44218 (N_44218,N_43558,N_43826);
nand U44219 (N_44219,N_42029,N_42244);
or U44220 (N_44220,N_42626,N_42545);
or U44221 (N_44221,N_42829,N_42971);
xor U44222 (N_44222,N_42995,N_42760);
or U44223 (N_44223,N_43704,N_43093);
xnor U44224 (N_44224,N_43938,N_42972);
and U44225 (N_44225,N_43536,N_42120);
nand U44226 (N_44226,N_42293,N_42565);
nor U44227 (N_44227,N_43430,N_43697);
or U44228 (N_44228,N_43717,N_42863);
nor U44229 (N_44229,N_43813,N_42236);
nor U44230 (N_44230,N_43595,N_43469);
nor U44231 (N_44231,N_43633,N_43302);
nand U44232 (N_44232,N_43177,N_42144);
and U44233 (N_44233,N_43470,N_43623);
and U44234 (N_44234,N_42543,N_42599);
nor U44235 (N_44235,N_43101,N_43117);
and U44236 (N_44236,N_43111,N_43353);
xnor U44237 (N_44237,N_43639,N_42322);
xor U44238 (N_44238,N_43058,N_42989);
or U44239 (N_44239,N_42476,N_43906);
or U44240 (N_44240,N_42681,N_43739);
nor U44241 (N_44241,N_43778,N_43941);
nand U44242 (N_44242,N_43322,N_42652);
nand U44243 (N_44243,N_42458,N_43498);
or U44244 (N_44244,N_42198,N_42453);
nor U44245 (N_44245,N_42286,N_43370);
nand U44246 (N_44246,N_43054,N_42572);
xor U44247 (N_44247,N_42382,N_42536);
xnor U44248 (N_44248,N_43834,N_43099);
nand U44249 (N_44249,N_43359,N_43955);
and U44250 (N_44250,N_42913,N_42035);
nor U44251 (N_44251,N_42867,N_42722);
nor U44252 (N_44252,N_43438,N_43042);
nor U44253 (N_44253,N_42665,N_43745);
xnor U44254 (N_44254,N_42593,N_42589);
and U44255 (N_44255,N_43956,N_43310);
or U44256 (N_44256,N_43463,N_43288);
xnor U44257 (N_44257,N_42020,N_42647);
xnor U44258 (N_44258,N_42575,N_43086);
and U44259 (N_44259,N_42372,N_43379);
nand U44260 (N_44260,N_42749,N_43196);
or U44261 (N_44261,N_42554,N_42591);
nand U44262 (N_44262,N_43533,N_43575);
nor U44263 (N_44263,N_42001,N_43387);
nor U44264 (N_44264,N_43060,N_42926);
nor U44265 (N_44265,N_42586,N_42055);
or U44266 (N_44266,N_43880,N_43452);
nor U44267 (N_44267,N_42446,N_43644);
or U44268 (N_44268,N_43357,N_43305);
and U44269 (N_44269,N_43920,N_43637);
nor U44270 (N_44270,N_42467,N_43724);
and U44271 (N_44271,N_43391,N_42964);
nor U44272 (N_44272,N_42279,N_42569);
and U44273 (N_44273,N_42925,N_42907);
xnor U44274 (N_44274,N_43415,N_42520);
xnor U44275 (N_44275,N_42892,N_42177);
xor U44276 (N_44276,N_42164,N_42504);
and U44277 (N_44277,N_43172,N_43730);
or U44278 (N_44278,N_43578,N_43979);
nand U44279 (N_44279,N_43589,N_42005);
and U44280 (N_44280,N_43335,N_42109);
and U44281 (N_44281,N_42525,N_43079);
and U44282 (N_44282,N_42232,N_42050);
nand U44283 (N_44283,N_42297,N_43349);
and U44284 (N_44284,N_42474,N_42089);
and U44285 (N_44285,N_42365,N_43474);
or U44286 (N_44286,N_43634,N_42419);
and U44287 (N_44287,N_43882,N_43268);
xnor U44288 (N_44288,N_43431,N_43000);
and U44289 (N_44289,N_43742,N_43220);
or U44290 (N_44290,N_43548,N_42672);
nand U44291 (N_44291,N_42721,N_43044);
and U44292 (N_44292,N_43209,N_43894);
nor U44293 (N_44293,N_43672,N_43256);
nor U44294 (N_44294,N_43532,N_43531);
nand U44295 (N_44295,N_42793,N_43667);
xor U44296 (N_44296,N_42879,N_42782);
xor U44297 (N_44297,N_42495,N_42411);
nor U44298 (N_44298,N_42406,N_43504);
and U44299 (N_44299,N_42191,N_43696);
or U44300 (N_44300,N_43141,N_42909);
nand U44301 (N_44301,N_42887,N_43508);
and U44302 (N_44302,N_43774,N_42688);
nand U44303 (N_44303,N_43382,N_42388);
or U44304 (N_44304,N_43240,N_43695);
nand U44305 (N_44305,N_42507,N_42112);
xnor U44306 (N_44306,N_43262,N_43568);
or U44307 (N_44307,N_42920,N_43809);
and U44308 (N_44308,N_43936,N_43102);
and U44309 (N_44309,N_43963,N_42834);
nor U44310 (N_44310,N_42573,N_43275);
xor U44311 (N_44311,N_43534,N_42741);
xor U44312 (N_44312,N_43158,N_43451);
nor U44313 (N_44313,N_43613,N_43652);
nand U44314 (N_44314,N_43503,N_42154);
xnor U44315 (N_44315,N_42414,N_43907);
xnor U44316 (N_44316,N_43486,N_42805);
and U44317 (N_44317,N_43569,N_43537);
xor U44318 (N_44318,N_42685,N_43641);
xor U44319 (N_44319,N_42409,N_42723);
or U44320 (N_44320,N_42189,N_42389);
nand U44321 (N_44321,N_43588,N_42929);
nand U44322 (N_44322,N_43949,N_43796);
nand U44323 (N_44323,N_43139,N_42559);
xor U44324 (N_44324,N_42178,N_42730);
or U44325 (N_44325,N_43380,N_43478);
nand U44326 (N_44326,N_43087,N_42095);
nor U44327 (N_44327,N_42455,N_43621);
and U44328 (N_44328,N_42702,N_43615);
or U44329 (N_44329,N_42321,N_43129);
nand U44330 (N_44330,N_43853,N_43297);
nor U44331 (N_44331,N_43750,N_42888);
nor U44332 (N_44332,N_43405,N_43318);
nand U44333 (N_44333,N_43663,N_42071);
nor U44334 (N_44334,N_43723,N_43687);
and U44335 (N_44335,N_43614,N_43519);
nand U44336 (N_44336,N_42982,N_42967);
and U44337 (N_44337,N_42523,N_42642);
or U44338 (N_44338,N_42151,N_43609);
nor U44339 (N_44339,N_43841,N_42511);
nor U44340 (N_44340,N_42640,N_43606);
nor U44341 (N_44341,N_43546,N_43838);
nor U44342 (N_44342,N_43792,N_43800);
xor U44343 (N_44343,N_42763,N_43417);
nor U44344 (N_44344,N_42258,N_43846);
and U44345 (N_44345,N_42225,N_42249);
or U44346 (N_44346,N_43762,N_43423);
or U44347 (N_44347,N_42168,N_42839);
nor U44348 (N_44348,N_43797,N_42912);
and U44349 (N_44349,N_43236,N_43163);
or U44350 (N_44350,N_42209,N_43458);
xnor U44351 (N_44351,N_42590,N_43795);
nand U44352 (N_44352,N_42115,N_42370);
or U44353 (N_44353,N_42082,N_42470);
and U44354 (N_44354,N_43239,N_43476);
nor U44355 (N_44355,N_42983,N_43231);
nand U44356 (N_44356,N_43871,N_42502);
xnor U44357 (N_44357,N_42263,N_42024);
xor U44358 (N_44358,N_43872,N_43818);
or U44359 (N_44359,N_42025,N_43976);
nor U44360 (N_44360,N_43827,N_42277);
and U44361 (N_44361,N_42111,N_43953);
and U44362 (N_44362,N_43026,N_43443);
and U44363 (N_44363,N_42003,N_43024);
xnor U44364 (N_44364,N_43655,N_42794);
nor U44365 (N_44365,N_43368,N_42385);
xor U44366 (N_44366,N_42459,N_43234);
nand U44367 (N_44367,N_43530,N_42905);
nor U44368 (N_44368,N_43170,N_43221);
xnor U44369 (N_44369,N_43317,N_42881);
and U44370 (N_44370,N_42398,N_43320);
or U44371 (N_44371,N_43932,N_43030);
or U44372 (N_44372,N_42171,N_42383);
nand U44373 (N_44373,N_42980,N_43909);
and U44374 (N_44374,N_43483,N_43807);
nor U44375 (N_44375,N_43741,N_43572);
or U44376 (N_44376,N_43673,N_43945);
or U44377 (N_44377,N_42648,N_42535);
nor U44378 (N_44378,N_43715,N_42731);
and U44379 (N_44379,N_42072,N_43410);
nor U44380 (N_44380,N_42284,N_43178);
and U44381 (N_44381,N_43903,N_42935);
nand U44382 (N_44382,N_43143,N_43034);
nor U44383 (N_44383,N_42689,N_42435);
nor U44384 (N_44384,N_42004,N_42835);
nor U44385 (N_44385,N_42063,N_42117);
nand U44386 (N_44386,N_43535,N_43011);
xnor U44387 (N_44387,N_43041,N_42740);
or U44388 (N_44388,N_43764,N_42758);
or U44389 (N_44389,N_43036,N_43915);
or U44390 (N_44390,N_43363,N_43988);
xnor U44391 (N_44391,N_43263,N_42942);
xor U44392 (N_44392,N_42687,N_42006);
xnor U44393 (N_44393,N_43334,N_43136);
and U44394 (N_44394,N_42578,N_42639);
nand U44395 (N_44395,N_43651,N_43365);
and U44396 (N_44396,N_42671,N_43883);
nor U44397 (N_44397,N_42347,N_43390);
or U44398 (N_44398,N_43429,N_42870);
xor U44399 (N_44399,N_43570,N_43985);
and U44400 (N_44400,N_42548,N_43005);
nand U44401 (N_44401,N_43587,N_42658);
or U44402 (N_44402,N_42970,N_42174);
xor U44403 (N_44403,N_42368,N_42694);
nor U44404 (N_44404,N_42895,N_43700);
nor U44405 (N_44405,N_43062,N_43607);
nor U44406 (N_44406,N_42998,N_42450);
nor U44407 (N_44407,N_42231,N_43092);
nand U44408 (N_44408,N_42551,N_43246);
and U44409 (N_44409,N_42836,N_42038);
xnor U44410 (N_44410,N_43489,N_43789);
xor U44411 (N_44411,N_43756,N_42744);
nand U44412 (N_44412,N_42362,N_42288);
nand U44413 (N_44413,N_43312,N_42742);
nand U44414 (N_44414,N_42108,N_42918);
and U44415 (N_44415,N_43065,N_43247);
nand U44416 (N_44416,N_42950,N_43484);
nand U44417 (N_44417,N_42588,N_42243);
or U44418 (N_44418,N_43142,N_43303);
nand U44419 (N_44419,N_43085,N_42503);
and U44420 (N_44420,N_42437,N_42841);
or U44421 (N_44421,N_42399,N_42434);
xnor U44422 (N_44422,N_43631,N_43059);
or U44423 (N_44423,N_43350,N_43261);
xor U44424 (N_44424,N_43206,N_42619);
xnor U44425 (N_44425,N_43981,N_42668);
nand U44426 (N_44426,N_43197,N_42036);
nor U44427 (N_44427,N_42564,N_43130);
or U44428 (N_44428,N_43866,N_42436);
and U44429 (N_44429,N_42715,N_43372);
xor U44430 (N_44430,N_43858,N_43817);
xor U44431 (N_44431,N_42047,N_42701);
nand U44432 (N_44432,N_42192,N_42945);
nand U44433 (N_44433,N_42438,N_42010);
nand U44434 (N_44434,N_43106,N_43021);
xnor U44435 (N_44435,N_43994,N_43144);
nor U44436 (N_44436,N_43596,N_43755);
and U44437 (N_44437,N_43625,N_43194);
and U44438 (N_44438,N_43798,N_42077);
nor U44439 (N_44439,N_43731,N_43110);
nand U44440 (N_44440,N_43480,N_43166);
or U44441 (N_44441,N_42187,N_42662);
nor U44442 (N_44442,N_42230,N_43344);
nand U44443 (N_44443,N_43381,N_43397);
or U44444 (N_44444,N_42051,N_43457);
and U44445 (N_44445,N_42130,N_42974);
xor U44446 (N_44446,N_43930,N_42848);
nor U44447 (N_44447,N_42291,N_42657);
nor U44448 (N_44448,N_43012,N_43439);
nand U44449 (N_44449,N_42427,N_43584);
and U44450 (N_44450,N_42601,N_42812);
and U44451 (N_44451,N_42894,N_42498);
nor U44452 (N_44452,N_43091,N_43345);
xnor U44453 (N_44453,N_43472,N_43726);
nand U44454 (N_44454,N_43754,N_42801);
nand U44455 (N_44455,N_43527,N_42393);
nor U44456 (N_44456,N_43455,N_43748);
and U44457 (N_44457,N_42202,N_43324);
and U44458 (N_44458,N_42500,N_42510);
nand U44459 (N_44459,N_43946,N_42298);
nor U44460 (N_44460,N_42629,N_43966);
and U44461 (N_44461,N_43661,N_42889);
and U44462 (N_44462,N_42135,N_43660);
nand U44463 (N_44463,N_42712,N_42831);
and U44464 (N_44464,N_42828,N_42947);
nor U44465 (N_44465,N_43124,N_43822);
nor U44466 (N_44466,N_43251,N_43709);
xnor U44467 (N_44467,N_42560,N_42976);
nand U44468 (N_44468,N_42311,N_43199);
or U44469 (N_44469,N_43400,N_43556);
nor U44470 (N_44470,N_42424,N_42022);
nand U44471 (N_44471,N_43097,N_43187);
xnor U44472 (N_44472,N_42644,N_42196);
nand U44473 (N_44473,N_42770,N_42349);
and U44474 (N_44474,N_43787,N_42963);
xor U44475 (N_44475,N_42506,N_43403);
or U44476 (N_44476,N_43608,N_43825);
nor U44477 (N_44477,N_42170,N_43497);
xor U44478 (N_44478,N_43892,N_42114);
and U44479 (N_44479,N_43554,N_42238);
nor U44480 (N_44480,N_43879,N_43815);
xnor U44481 (N_44481,N_43257,N_43645);
or U44482 (N_44482,N_43160,N_42579);
or U44483 (N_44483,N_42924,N_43662);
nor U44484 (N_44484,N_42773,N_42211);
nand U44485 (N_44485,N_43701,N_42292);
nor U44486 (N_44486,N_42410,N_42602);
and U44487 (N_44487,N_42954,N_42254);
xnor U44488 (N_44488,N_43171,N_43122);
nor U44489 (N_44489,N_42745,N_42339);
xor U44490 (N_44490,N_42883,N_42726);
nand U44491 (N_44491,N_42915,N_42582);
and U44492 (N_44492,N_42802,N_43629);
or U44493 (N_44493,N_42462,N_42337);
or U44494 (N_44494,N_42280,N_43138);
xor U44495 (N_44495,N_42856,N_42423);
or U44496 (N_44496,N_43342,N_42853);
and U44497 (N_44497,N_42295,N_43152);
nor U44498 (N_44498,N_42452,N_42053);
nand U44499 (N_44499,N_42207,N_42343);
or U44500 (N_44500,N_43465,N_42817);
nor U44501 (N_44501,N_42654,N_42986);
and U44502 (N_44502,N_42247,N_43794);
or U44503 (N_44503,N_43738,N_42137);
nand U44504 (N_44504,N_43201,N_42751);
xnor U44505 (N_44505,N_42121,N_43591);
nor U44506 (N_44506,N_42994,N_42900);
nand U44507 (N_44507,N_43464,N_43183);
nor U44508 (N_44508,N_42070,N_42253);
nor U44509 (N_44509,N_42847,N_42483);
nand U44510 (N_44510,N_42392,N_43274);
or U44511 (N_44511,N_42641,N_43942);
nand U44512 (N_44512,N_43808,N_43528);
and U44513 (N_44513,N_42145,N_42800);
nor U44514 (N_44514,N_42524,N_42934);
xor U44515 (N_44515,N_43828,N_42734);
nand U44516 (N_44516,N_43156,N_42821);
xnor U44517 (N_44517,N_43620,N_42627);
nor U44518 (N_44518,N_42743,N_42669);
or U44519 (N_44519,N_43361,N_42612);
and U44520 (N_44520,N_42808,N_43680);
or U44521 (N_44521,N_43326,N_42464);
nand U44522 (N_44522,N_43273,N_43874);
nor U44523 (N_44523,N_42394,N_43378);
nand U44524 (N_44524,N_42405,N_42608);
nor U44525 (N_44525,N_42903,N_42604);
or U44526 (N_44526,N_42468,N_43628);
and U44527 (N_44527,N_43586,N_43482);
or U44528 (N_44528,N_43744,N_42531);
or U44529 (N_44529,N_43098,N_43812);
and U44530 (N_44530,N_43066,N_42792);
nand U44531 (N_44531,N_43746,N_43108);
or U44532 (N_44532,N_42809,N_43524);
and U44533 (N_44533,N_43161,N_43965);
nor U44534 (N_44534,N_43500,N_43565);
nand U44535 (N_44535,N_43210,N_43115);
and U44536 (N_44536,N_42946,N_43924);
or U44537 (N_44537,N_42155,N_42377);
or U44538 (N_44538,N_43888,N_43592);
nor U44539 (N_44539,N_43799,N_43113);
or U44540 (N_44540,N_42309,N_43193);
nand U44541 (N_44541,N_43992,N_43259);
nand U44542 (N_44542,N_43475,N_42282);
nand U44543 (N_44543,N_43038,N_42465);
and U44544 (N_44544,N_42143,N_42729);
nand U44545 (N_44545,N_43167,N_43505);
nand U44546 (N_44546,N_42997,N_42965);
nand U44547 (N_44547,N_42148,N_42000);
and U44548 (N_44548,N_42813,N_42033);
or U44549 (N_44549,N_42966,N_42775);
and U44550 (N_44550,N_42666,N_42342);
and U44551 (N_44551,N_42276,N_43014);
nor U44552 (N_44552,N_42566,N_42940);
nor U44553 (N_44553,N_42851,N_42615);
and U44554 (N_44554,N_42320,N_43848);
and U44555 (N_44555,N_42732,N_42442);
nor U44556 (N_44556,N_43270,N_42538);
nor U44557 (N_44557,N_43881,N_42992);
or U44558 (N_44558,N_43490,N_43467);
or U44559 (N_44559,N_43362,N_43126);
or U44560 (N_44560,N_43681,N_43502);
xor U44561 (N_44561,N_42336,N_42528);
nor U44562 (N_44562,N_42097,N_43770);
or U44563 (N_44563,N_42718,N_43616);
and U44564 (N_44564,N_42056,N_42636);
xor U44565 (N_44565,N_42709,N_42166);
and U44566 (N_44566,N_42163,N_43244);
nor U44567 (N_44567,N_43281,N_43132);
and U44568 (N_44568,N_42106,N_42923);
and U44569 (N_44569,N_42016,N_42754);
or U44570 (N_44570,N_43890,N_42778);
or U44571 (N_44571,N_43619,N_42183);
nand U44572 (N_44572,N_43367,N_42134);
xnor U44573 (N_44573,N_42181,N_42273);
nor U44574 (N_44574,N_42563,N_43182);
nor U44575 (N_44575,N_43910,N_42584);
and U44576 (N_44576,N_42625,N_43181);
or U44577 (N_44577,N_42633,N_42182);
and U44578 (N_44578,N_43150,N_42670);
nand U44579 (N_44579,N_42042,N_43377);
nand U44580 (N_44580,N_43401,N_43806);
nand U44581 (N_44581,N_43690,N_43441);
nand U44582 (N_44582,N_43947,N_43260);
nor U44583 (N_44583,N_42131,N_42046);
xnor U44584 (N_44584,N_43088,N_42100);
xnor U44585 (N_44585,N_43409,N_42028);
and U44586 (N_44586,N_43839,N_42650);
or U44587 (N_44587,N_43237,N_43157);
or U44588 (N_44588,N_43852,N_42136);
xor U44589 (N_44589,N_42891,N_42840);
nor U44590 (N_44590,N_42960,N_42833);
nand U44591 (N_44591,N_43819,N_42826);
nand U44592 (N_44592,N_43788,N_42663);
nor U44593 (N_44593,N_43914,N_43040);
and U44594 (N_44594,N_42251,N_42401);
nand U44595 (N_44595,N_42990,N_42264);
nand U44596 (N_44596,N_42882,N_42113);
xnor U44597 (N_44597,N_42832,N_43939);
nor U44598 (N_44598,N_42845,N_43684);
nor U44599 (N_44599,N_42330,N_43479);
and U44600 (N_44600,N_43677,N_43286);
nor U44601 (N_44601,N_43957,N_42223);
xor U44602 (N_44602,N_43698,N_42661);
nand U44603 (N_44603,N_43993,N_43705);
nand U44604 (N_44604,N_42013,N_43067);
xnor U44605 (N_44605,N_42127,N_43188);
nand U44606 (N_44606,N_43422,N_43520);
and U44607 (N_44607,N_42790,N_43916);
or U44608 (N_44608,N_42842,N_42014);
and U44609 (N_44609,N_42541,N_43491);
nand U44610 (N_44610,N_43019,N_43720);
or U44611 (N_44611,N_42860,N_43868);
or U44612 (N_44612,N_42449,N_43462);
or U44613 (N_44613,N_42674,N_42364);
or U44614 (N_44614,N_42737,N_43605);
nor U44615 (N_44615,N_42371,N_43118);
and U44616 (N_44616,N_43833,N_42583);
nand U44617 (N_44617,N_43666,N_43786);
and U44618 (N_44618,N_43752,N_42324);
nor U44619 (N_44619,N_42886,N_43148);
or U44620 (N_44620,N_42938,N_42948);
nand U44621 (N_44621,N_42675,N_42429);
or U44622 (N_44622,N_43406,N_43290);
xor U44623 (N_44623,N_42735,N_43235);
nor U44624 (N_44624,N_43384,N_43074);
or U44625 (N_44625,N_42210,N_42268);
nor U44626 (N_44626,N_42844,N_43298);
and U44627 (N_44627,N_43721,N_43081);
xnor U44628 (N_44628,N_42252,N_42125);
nand U44629 (N_44629,N_43991,N_43933);
or U44630 (N_44630,N_42516,N_42386);
or U44631 (N_44631,N_42141,N_43725);
nand U44632 (N_44632,N_43104,N_43017);
xor U44633 (N_44633,N_42188,N_43119);
and U44634 (N_44634,N_42384,N_43090);
or U44635 (N_44635,N_42260,N_42200);
xnor U44636 (N_44636,N_42621,N_43935);
or U44637 (N_44637,N_43025,N_43071);
and U44638 (N_44638,N_43219,N_42305);
nor U44639 (N_44639,N_42542,N_43029);
or U44640 (N_44640,N_43867,N_42255);
xnor U44641 (N_44641,N_43105,N_43016);
and U44642 (N_44642,N_43538,N_43542);
or U44643 (N_44643,N_43421,N_43559);
nor U44644 (N_44644,N_42521,N_42943);
or U44645 (N_44645,N_42289,N_43418);
nor U44646 (N_44646,N_42156,N_43385);
and U44647 (N_44647,N_42147,N_43083);
nand U44648 (N_44648,N_43205,N_42041);
xnor U44649 (N_44649,N_42356,N_43925);
and U44650 (N_44650,N_43654,N_42508);
nand U44651 (N_44651,N_43694,N_43647);
and U44652 (N_44652,N_42772,N_42190);
and U44653 (N_44653,N_42246,N_43094);
or U44654 (N_44654,N_43306,N_42492);
nand U44655 (N_44655,N_43728,N_43223);
or U44656 (N_44656,N_43328,N_43747);
and U44657 (N_44657,N_43579,N_42354);
or U44658 (N_44658,N_42359,N_43023);
xor U44659 (N_44659,N_42746,N_42397);
nor U44660 (N_44660,N_42221,N_42594);
xnor U44661 (N_44661,N_42402,N_42126);
nand U44662 (N_44662,N_43972,N_42197);
xor U44663 (N_44663,N_42707,N_43970);
xor U44664 (N_44664,N_43389,N_43140);
xor U44665 (N_44665,N_43233,N_43198);
xnor U44666 (N_44666,N_43186,N_43901);
or U44667 (N_44667,N_42307,N_43207);
or U44668 (N_44668,N_43877,N_43931);
xnor U44669 (N_44669,N_43594,N_43740);
nand U44670 (N_44670,N_42257,N_43055);
and U44671 (N_44671,N_42592,N_42628);
and U44672 (N_44672,N_42958,N_43184);
nand U44673 (N_44673,N_43364,N_42683);
xor U44674 (N_44674,N_43332,N_42777);
xor U44675 (N_44675,N_43515,N_43394);
and U44676 (N_44676,N_42962,N_42823);
and U44677 (N_44677,N_43969,N_43047);
nor U44678 (N_44678,N_43447,N_42704);
nor U44679 (N_44679,N_43904,N_42944);
nand U44680 (N_44680,N_42485,N_42932);
nor U44681 (N_44681,N_43407,N_43149);
nand U44682 (N_44682,N_42463,N_42562);
nand U44683 (N_44683,N_42340,N_43702);
nor U44684 (N_44684,N_42123,N_43873);
or U44685 (N_44685,N_43064,N_42094);
xor U44686 (N_44686,N_43376,N_43763);
and U44687 (N_44687,N_43688,N_42444);
nand U44688 (N_44688,N_43351,N_42533);
nand U44689 (N_44689,N_42146,N_42939);
nor U44690 (N_44690,N_42092,N_42752);
xnor U44691 (N_44691,N_42205,N_43204);
or U44692 (N_44692,N_43618,N_43070);
nand U44693 (N_44693,N_43352,N_43980);
or U44694 (N_44694,N_43599,N_42327);
and U44695 (N_44695,N_42158,N_42172);
xor U44696 (N_44696,N_43039,N_42314);
nor U44697 (N_44697,N_42285,N_43905);
xnor U44698 (N_44698,N_43779,N_42771);
and U44699 (N_44699,N_42299,N_42899);
xnor U44700 (N_44700,N_43020,N_42489);
xor U44701 (N_44701,N_43411,N_43009);
nand U44702 (N_44702,N_43743,N_42068);
and U44703 (N_44703,N_43566,N_42204);
xnor U44704 (N_44704,N_42610,N_42472);
nand U44705 (N_44705,N_43413,N_43844);
and U44706 (N_44706,N_42755,N_42814);
nor U44707 (N_44707,N_42864,N_43832);
or U44708 (N_44708,N_43857,N_43791);
nand U44709 (N_44709,N_43632,N_43665);
and U44710 (N_44710,N_42066,N_42574);
nand U44711 (N_44711,N_43493,N_42030);
or U44712 (N_44712,N_42783,N_43521);
nand U44713 (N_44713,N_43294,N_42757);
and U44714 (N_44714,N_43341,N_43433);
or U44715 (N_44715,N_43734,N_43636);
nor U44716 (N_44716,N_43849,N_43805);
xnor U44717 (N_44717,N_43004,N_42953);
xor U44718 (N_44718,N_43863,N_42357);
nand U44719 (N_44719,N_42747,N_43162);
or U44720 (N_44720,N_43889,N_42169);
or U44721 (N_44721,N_43010,N_42228);
and U44722 (N_44722,N_43648,N_42700);
and U44723 (N_44723,N_43835,N_42922);
nand U44724 (N_44724,N_43624,N_43682);
and U44725 (N_44725,N_42048,N_42567);
and U44726 (N_44726,N_43785,N_43252);
nand U44727 (N_44727,N_43649,N_43610);
nand U44728 (N_44728,N_42161,N_42499);
nor U44729 (N_44729,N_43285,N_43271);
xnor U44730 (N_44730,N_43545,N_43543);
nor U44731 (N_44731,N_43861,N_42914);
nor U44732 (N_44732,N_42645,N_43155);
xor U44733 (N_44733,N_42235,N_43960);
and U44734 (N_44734,N_42457,N_43821);
nand U44735 (N_44735,N_43501,N_43954);
or U44736 (N_44736,N_42303,N_43975);
and U44737 (N_44737,N_42344,N_42009);
nand U44738 (N_44738,N_42150,N_42547);
or U44739 (N_44739,N_42233,N_42865);
xor U44740 (N_44740,N_42312,N_42660);
nand U44741 (N_44741,N_42380,N_43790);
nor U44742 (N_44742,N_43898,N_42358);
xnor U44743 (N_44743,N_43900,N_42379);
xor U44744 (N_44744,N_42116,N_42226);
or U44745 (N_44745,N_43308,N_42037);
xnor U44746 (N_44746,N_43507,N_42256);
xor U44747 (N_44747,N_42969,N_42241);
or U44748 (N_44748,N_42850,N_42638);
and U44749 (N_44749,N_42329,N_43814);
nor U44750 (N_44750,N_43674,N_42348);
or U44751 (N_44751,N_42634,N_42568);
nand U44752 (N_44752,N_43253,N_42955);
xor U44753 (N_44753,N_43597,N_42315);
or U44754 (N_44754,N_43847,N_42553);
and U44755 (N_44755,N_42690,N_43911);
nand U44756 (N_44756,N_43804,N_42065);
or U44757 (N_44757,N_43593,N_42616);
nor U44758 (N_44758,N_43027,N_42184);
nand U44759 (N_44759,N_42007,N_43923);
or U44760 (N_44760,N_42043,N_43855);
or U44761 (N_44761,N_42294,N_43902);
nand U44762 (N_44762,N_42876,N_42308);
nor U44763 (N_44763,N_42418,N_43444);
xnor U44764 (N_44764,N_43998,N_43689);
or U44765 (N_44765,N_43776,N_42884);
or U44766 (N_44766,N_43114,N_42806);
nand U44767 (N_44767,N_42387,N_42635);
and U44768 (N_44768,N_43617,N_42101);
and U44769 (N_44769,N_43147,N_43258);
xor U44770 (N_44770,N_42031,N_43037);
and U44771 (N_44771,N_42049,N_42319);
nor U44772 (N_44772,N_43284,N_42885);
nand U44773 (N_44773,N_43046,N_43035);
or U44774 (N_44774,N_42175,N_42693);
xnor U44775 (N_44775,N_42558,N_43753);
nor U44776 (N_44776,N_43891,N_42149);
or U44777 (N_44777,N_43112,N_42857);
nand U44778 (N_44778,N_43918,N_43424);
nand U44779 (N_44779,N_43222,N_42540);
nor U44780 (N_44780,N_43265,N_43571);
nor U44781 (N_44781,N_43287,N_43425);
and U44782 (N_44782,N_43436,N_42199);
xor U44783 (N_44783,N_43506,N_42653);
nor U44784 (N_44784,N_42878,N_43153);
nor U44785 (N_44785,N_43712,N_43710);
or U44786 (N_44786,N_42937,N_43760);
nor U44787 (N_44787,N_43626,N_43719);
and U44788 (N_44788,N_42614,N_43664);
and U44789 (N_44789,N_43811,N_42534);
nor U44790 (N_44790,N_42512,N_42787);
nand U44791 (N_44791,N_42788,N_43045);
nor U44792 (N_44792,N_43668,N_42795);
or U44793 (N_44793,N_42539,N_43494);
and U44794 (N_44794,N_43200,N_43173);
nor U44795 (N_44795,N_42720,N_42128);
nand U44796 (N_44796,N_43048,N_42780);
nor U44797 (N_44797,N_43830,N_42432);
xnor U44798 (N_44798,N_43232,N_43950);
or U44799 (N_44799,N_42219,N_42390);
xor U44800 (N_44800,N_42363,N_43073);
xnor U44801 (N_44801,N_42090,N_42482);
and U44802 (N_44802,N_42952,N_43103);
xor U44803 (N_44803,N_43095,N_42180);
nand U44804 (N_44804,N_42975,N_42496);
or U44805 (N_44805,N_43057,N_42973);
and U44806 (N_44806,N_43488,N_42765);
nor U44807 (N_44807,N_42040,N_43323);
xor U44808 (N_44808,N_42360,N_43043);
and U44809 (N_44809,N_42916,N_43131);
nor U44810 (N_44810,N_42448,N_43856);
nor U44811 (N_44811,N_42338,N_42874);
nor U44812 (N_44812,N_43292,N_42977);
and U44813 (N_44813,N_42843,N_42456);
and U44814 (N_44814,N_43782,N_42032);
nand U44815 (N_44815,N_42133,N_43990);
nand U44816 (N_44816,N_43860,N_43134);
nand U44817 (N_44817,N_42373,N_42227);
or U44818 (N_44818,N_42830,N_43761);
xnor U44819 (N_44819,N_42475,N_42098);
nand U44820 (N_44820,N_43944,N_42949);
and U44821 (N_44821,N_42786,N_43492);
and U44822 (N_44822,N_42407,N_42433);
or U44823 (N_44823,N_43369,N_43958);
nor U44824 (N_44824,N_42099,N_43711);
and U44825 (N_44825,N_43917,N_43509);
xnor U44826 (N_44826,N_43254,N_42021);
xnor U44827 (N_44827,N_43300,N_42561);
nand U44828 (N_44828,N_42999,N_43895);
and U44829 (N_44829,N_42159,N_42325);
nor U44830 (N_44830,N_42705,N_42799);
nand U44831 (N_44831,N_42875,N_43227);
xnor U44832 (N_44832,N_42673,N_42519);
xnor U44833 (N_44833,N_42769,N_42785);
nand U44834 (N_44834,N_43510,N_43769);
nand U44835 (N_44835,N_42789,N_43564);
xor U44836 (N_44836,N_43154,N_43164);
nand U44837 (N_44837,N_43217,N_42968);
nand U44838 (N_44838,N_42093,N_43449);
and U44839 (N_44839,N_43128,N_42440);
or U44840 (N_44840,N_43355,N_42491);
xor U44841 (N_44841,N_43899,N_42234);
or U44842 (N_44842,N_42374,N_42103);
nand U44843 (N_44843,N_43255,N_43737);
and U44844 (N_44844,N_42684,N_42768);
and U44845 (N_44845,N_42811,N_42698);
or U44846 (N_44846,N_43585,N_43434);
xor U44847 (N_44847,N_43008,N_43190);
or U44848 (N_44848,N_43264,N_42606);
and U44849 (N_44849,N_43948,N_42631);
nand U44850 (N_44850,N_42376,N_42695);
or U44851 (N_44851,N_43854,N_43331);
and U44852 (N_44852,N_42083,N_42526);
and U44853 (N_44853,N_43213,N_42861);
and U44854 (N_44854,N_42515,N_43896);
nand U44855 (N_44855,N_43358,N_42479);
xor U44856 (N_44856,N_43245,N_43768);
or U44857 (N_44857,N_42366,N_42697);
xor U44858 (N_44858,N_42555,N_43885);
and U44859 (N_44859,N_43707,N_43461);
xor U44860 (N_44860,N_43137,N_42300);
nor U44861 (N_44861,N_43386,N_42871);
xor U44862 (N_44862,N_43450,N_43360);
or U44863 (N_44863,N_42477,N_43783);
nor U44864 (N_44864,N_42008,N_42176);
and U44865 (N_44865,N_43192,N_42901);
xnor U44866 (N_44866,N_42605,N_43165);
nand U44867 (N_44867,N_43224,N_43780);
and U44868 (N_44868,N_42301,N_43068);
xor U44869 (N_44869,N_43837,N_43716);
and U44870 (N_44870,N_42361,N_43446);
nand U44871 (N_44871,N_42956,N_43460);
nor U44872 (N_44872,N_42852,N_42091);
nor U44873 (N_44873,N_42096,N_42017);
xor U44874 (N_44874,N_43929,N_42443);
nand U44875 (N_44875,N_42430,N_43080);
nand U44876 (N_44876,N_43218,N_42283);
and U44877 (N_44877,N_42165,N_42804);
or U44878 (N_44878,N_43203,N_42067);
nand U44879 (N_44879,N_42002,N_42224);
and U44880 (N_44880,N_43243,N_42776);
nand U44881 (N_44881,N_42873,N_43031);
xor U44882 (N_44882,N_43851,N_43314);
and U44883 (N_44883,N_43347,N_43886);
and U44884 (N_44884,N_43884,N_42381);
or U44885 (N_44885,N_42087,N_42206);
nand U44886 (N_44886,N_43339,N_42931);
nor U44887 (N_44887,N_42404,N_42140);
nand U44888 (N_44888,N_43611,N_43573);
xor U44889 (N_44889,N_42270,N_42259);
and U44890 (N_44890,N_42784,N_42762);
nand U44891 (N_44891,N_42951,N_42509);
nand U44892 (N_44892,N_42266,N_42119);
nor U44893 (N_44893,N_43454,N_42649);
xnor U44894 (N_44894,N_42643,N_43123);
xor U44895 (N_44895,N_42544,N_43842);
nor U44896 (N_44896,N_42152,N_43823);
nand U44897 (N_44897,N_43971,N_42105);
nor U44898 (N_44898,N_42898,N_42290);
xor U44899 (N_44899,N_43356,N_43225);
or U44900 (N_44900,N_42217,N_43685);
and U44901 (N_44901,N_42928,N_43448);
xor U44902 (N_44902,N_42646,N_42897);
xnor U44903 (N_44903,N_43550,N_42810);
and U44904 (N_44904,N_43777,N_43627);
or U44905 (N_44905,N_42403,N_43650);
nand U44906 (N_44906,N_42719,N_43338);
nand U44907 (N_44907,N_43974,N_42676);
xor U44908 (N_44908,N_42807,N_42267);
or U44909 (N_44909,N_43864,N_42167);
xnor U44910 (N_44910,N_42656,N_43829);
xnor U44911 (N_44911,N_43396,N_43952);
and U44912 (N_44912,N_43084,N_42927);
xnor U44913 (N_44913,N_43598,N_42138);
and U44914 (N_44914,N_43419,N_43269);
xor U44915 (N_44915,N_43373,N_42415);
xor U44916 (N_44916,N_43366,N_42984);
xnor U44917 (N_44917,N_43968,N_42611);
nand U44918 (N_44918,N_43001,N_42057);
xnor U44919 (N_44919,N_42480,N_42724);
nand U44920 (N_44920,N_42549,N_43870);
nand U44921 (N_44921,N_43512,N_43714);
xor U44922 (N_44922,N_42803,N_42710);
or U44923 (N_44923,N_43959,N_43802);
xor U44924 (N_44924,N_42478,N_43499);
nand U44925 (N_44925,N_42447,N_43151);
nor U44926 (N_44926,N_43309,N_43051);
and U44927 (N_44927,N_43279,N_42426);
and U44928 (N_44928,N_43393,N_42218);
xnor U44929 (N_44929,N_43321,N_42598);
nand U44930 (N_44930,N_42441,N_43706);
nand U44931 (N_44931,N_43732,N_43437);
and U44932 (N_44932,N_43289,N_42081);
nand U44933 (N_44933,N_42630,N_42522);
and U44934 (N_44934,N_43887,N_43557);
nor U44935 (N_44935,N_43277,N_43602);
and U44936 (N_44936,N_43276,N_43640);
nor U44937 (N_44937,N_42880,N_42262);
xor U44938 (N_44938,N_43127,N_42846);
nor U44939 (N_44939,N_42691,N_43912);
xnor U44940 (N_44940,N_42696,N_43526);
xor U44941 (N_44941,N_43325,N_42936);
nand U44942 (N_44942,N_42078,N_43089);
xnor U44943 (N_44943,N_42620,N_42607);
xor U44944 (N_44944,N_43145,N_43295);
or U44945 (N_44945,N_43146,N_43843);
nor U44946 (N_44946,N_43179,N_43282);
nand U44947 (N_44947,N_43307,N_43577);
nand U44948 (N_44948,N_42341,N_43962);
nor U44949 (N_44949,N_43398,N_42727);
or U44950 (N_44950,N_42201,N_43291);
or U44951 (N_44951,N_43272,N_42353);
or U44952 (N_44952,N_42585,N_42445);
and U44953 (N_44953,N_42222,N_43440);
and U44954 (N_44954,N_42026,N_43228);
or U44955 (N_44955,N_43984,N_42959);
and U44956 (N_44956,N_42069,N_42104);
and U44957 (N_44957,N_42304,N_42466);
and U44958 (N_44958,N_42350,N_43875);
nor U44959 (N_44959,N_42195,N_43576);
xor U44960 (N_44960,N_43996,N_43973);
and U44961 (N_44961,N_43056,N_42571);
nand U44962 (N_44962,N_42996,N_42451);
xnor U44963 (N_44963,N_42767,N_42054);
nand U44964 (N_44964,N_43718,N_42822);
or U44965 (N_44965,N_42988,N_42118);
xor U44966 (N_44966,N_42060,N_43683);
nor U44967 (N_44967,N_43241,N_42497);
xnor U44968 (N_44968,N_43735,N_42213);
and U44969 (N_44969,N_43327,N_43590);
nor U44970 (N_44970,N_43869,N_42015);
nor U44971 (N_44971,N_43069,N_43468);
and U44972 (N_44972,N_42064,N_42274);
nor U44973 (N_44973,N_43195,N_42854);
and U44974 (N_44974,N_43329,N_43072);
or U44975 (N_44975,N_42162,N_43820);
nor U44976 (N_44976,N_42978,N_42310);
and U44977 (N_44977,N_43563,N_42278);
nand U44978 (N_44978,N_42416,N_42748);
nor U44979 (N_44979,N_42248,N_42215);
or U44980 (N_44980,N_43604,N_43574);
and U44981 (N_44981,N_43601,N_43670);
nor U44982 (N_44982,N_43238,N_43612);
xor U44983 (N_44983,N_42651,N_43784);
xnor U44984 (N_44984,N_43211,N_43100);
or U44985 (N_44985,N_42759,N_42454);
and U44986 (N_44986,N_43708,N_42352);
xnor U44987 (N_44987,N_42911,N_42587);
xor U44988 (N_44988,N_43315,N_43299);
or U44989 (N_44989,N_43921,N_43997);
nand U44990 (N_44990,N_43189,N_42261);
and U44991 (N_44991,N_43337,N_43033);
nand U44992 (N_44992,N_42062,N_43816);
and U44993 (N_44993,N_42179,N_42208);
nand U44994 (N_44994,N_42173,N_43733);
or U44995 (N_44995,N_42921,N_42714);
and U44996 (N_44996,N_43862,N_42425);
nor U44997 (N_44997,N_42074,N_43765);
and U44998 (N_44998,N_43758,N_42796);
and U44999 (N_44999,N_43630,N_43922);
and U45000 (N_45000,N_43742,N_42280);
or U45001 (N_45001,N_43326,N_42330);
or U45002 (N_45002,N_42923,N_42887);
nor U45003 (N_45003,N_43519,N_42328);
or U45004 (N_45004,N_43555,N_42318);
nand U45005 (N_45005,N_42195,N_42738);
and U45006 (N_45006,N_43125,N_42875);
xnor U45007 (N_45007,N_43653,N_43119);
nor U45008 (N_45008,N_43858,N_43302);
or U45009 (N_45009,N_43797,N_43940);
nor U45010 (N_45010,N_43414,N_42849);
nor U45011 (N_45011,N_42963,N_43514);
xor U45012 (N_45012,N_42292,N_43569);
xnor U45013 (N_45013,N_43399,N_43318);
xnor U45014 (N_45014,N_42492,N_43908);
and U45015 (N_45015,N_42697,N_43226);
and U45016 (N_45016,N_43822,N_42994);
nor U45017 (N_45017,N_43802,N_42177);
xnor U45018 (N_45018,N_43517,N_42251);
nand U45019 (N_45019,N_42254,N_43177);
xnor U45020 (N_45020,N_42433,N_43977);
and U45021 (N_45021,N_43283,N_42964);
nor U45022 (N_45022,N_43481,N_43388);
nor U45023 (N_45023,N_42785,N_43405);
nand U45024 (N_45024,N_43476,N_43441);
and U45025 (N_45025,N_42615,N_43278);
or U45026 (N_45026,N_43268,N_42392);
nand U45027 (N_45027,N_43958,N_42178);
xor U45028 (N_45028,N_43886,N_43133);
nand U45029 (N_45029,N_43401,N_42525);
and U45030 (N_45030,N_43223,N_43377);
nand U45031 (N_45031,N_42058,N_42234);
nor U45032 (N_45032,N_43067,N_42711);
or U45033 (N_45033,N_42038,N_42346);
nand U45034 (N_45034,N_42628,N_42939);
nor U45035 (N_45035,N_43829,N_42870);
nor U45036 (N_45036,N_43975,N_43845);
and U45037 (N_45037,N_43724,N_43431);
xor U45038 (N_45038,N_42121,N_42309);
xor U45039 (N_45039,N_42124,N_43302);
nor U45040 (N_45040,N_42690,N_43880);
xnor U45041 (N_45041,N_43554,N_42855);
nor U45042 (N_45042,N_43694,N_43704);
and U45043 (N_45043,N_42150,N_43159);
nor U45044 (N_45044,N_42271,N_43702);
nor U45045 (N_45045,N_42848,N_42348);
nor U45046 (N_45046,N_42148,N_42473);
or U45047 (N_45047,N_43794,N_43388);
or U45048 (N_45048,N_43147,N_43256);
and U45049 (N_45049,N_42721,N_42712);
xnor U45050 (N_45050,N_43177,N_43821);
nor U45051 (N_45051,N_42739,N_42626);
xor U45052 (N_45052,N_43547,N_43861);
and U45053 (N_45053,N_43423,N_42661);
and U45054 (N_45054,N_43374,N_43216);
nor U45055 (N_45055,N_42027,N_42934);
xnor U45056 (N_45056,N_43228,N_43454);
or U45057 (N_45057,N_43670,N_42401);
xnor U45058 (N_45058,N_43431,N_43327);
or U45059 (N_45059,N_43904,N_42984);
nor U45060 (N_45060,N_42665,N_43801);
nand U45061 (N_45061,N_42764,N_42567);
nor U45062 (N_45062,N_43589,N_42932);
nor U45063 (N_45063,N_43159,N_43380);
or U45064 (N_45064,N_43452,N_42003);
nor U45065 (N_45065,N_42681,N_42660);
nand U45066 (N_45066,N_42078,N_42128);
and U45067 (N_45067,N_42088,N_43964);
or U45068 (N_45068,N_42663,N_43652);
or U45069 (N_45069,N_43324,N_43723);
nand U45070 (N_45070,N_42715,N_43414);
xnor U45071 (N_45071,N_43656,N_42285);
nand U45072 (N_45072,N_43824,N_42373);
and U45073 (N_45073,N_43270,N_43206);
nor U45074 (N_45074,N_42276,N_43820);
nand U45075 (N_45075,N_42962,N_42828);
nand U45076 (N_45076,N_42247,N_43211);
xnor U45077 (N_45077,N_43676,N_43132);
and U45078 (N_45078,N_42396,N_42534);
nor U45079 (N_45079,N_42714,N_42200);
nand U45080 (N_45080,N_42193,N_42074);
or U45081 (N_45081,N_43169,N_43720);
nand U45082 (N_45082,N_42382,N_42858);
or U45083 (N_45083,N_43719,N_42906);
xor U45084 (N_45084,N_42600,N_42172);
and U45085 (N_45085,N_43039,N_42540);
nor U45086 (N_45086,N_43074,N_42394);
nor U45087 (N_45087,N_43555,N_42728);
nor U45088 (N_45088,N_42784,N_43258);
or U45089 (N_45089,N_43813,N_43311);
and U45090 (N_45090,N_42302,N_43110);
and U45091 (N_45091,N_42305,N_43773);
and U45092 (N_45092,N_42686,N_43583);
or U45093 (N_45093,N_42963,N_42455);
nor U45094 (N_45094,N_42967,N_43133);
xnor U45095 (N_45095,N_42262,N_43376);
xor U45096 (N_45096,N_43765,N_43643);
or U45097 (N_45097,N_42915,N_43216);
nand U45098 (N_45098,N_42082,N_42522);
or U45099 (N_45099,N_43556,N_42920);
nor U45100 (N_45100,N_43848,N_42077);
nor U45101 (N_45101,N_43303,N_43173);
xor U45102 (N_45102,N_42814,N_43501);
nand U45103 (N_45103,N_43996,N_42939);
and U45104 (N_45104,N_42325,N_43543);
or U45105 (N_45105,N_43514,N_43542);
and U45106 (N_45106,N_43795,N_43641);
xnor U45107 (N_45107,N_42170,N_43164);
and U45108 (N_45108,N_42240,N_43908);
nand U45109 (N_45109,N_43316,N_43956);
nor U45110 (N_45110,N_42759,N_42568);
nand U45111 (N_45111,N_42854,N_42649);
nor U45112 (N_45112,N_42581,N_42075);
or U45113 (N_45113,N_43017,N_43675);
and U45114 (N_45114,N_42772,N_43030);
nor U45115 (N_45115,N_43695,N_42641);
and U45116 (N_45116,N_43274,N_42438);
or U45117 (N_45117,N_43333,N_42806);
nor U45118 (N_45118,N_43565,N_43733);
or U45119 (N_45119,N_42176,N_42215);
or U45120 (N_45120,N_42284,N_43104);
and U45121 (N_45121,N_42032,N_43646);
nand U45122 (N_45122,N_42787,N_42586);
or U45123 (N_45123,N_42867,N_43080);
and U45124 (N_45124,N_43846,N_43218);
xnor U45125 (N_45125,N_42415,N_42214);
and U45126 (N_45126,N_42539,N_43953);
nor U45127 (N_45127,N_42133,N_43589);
nand U45128 (N_45128,N_42819,N_42255);
nand U45129 (N_45129,N_43394,N_42144);
xnor U45130 (N_45130,N_42134,N_42933);
or U45131 (N_45131,N_42802,N_42388);
or U45132 (N_45132,N_42123,N_42301);
nand U45133 (N_45133,N_42603,N_42270);
xnor U45134 (N_45134,N_42722,N_42974);
nor U45135 (N_45135,N_43456,N_43732);
nand U45136 (N_45136,N_42209,N_43207);
and U45137 (N_45137,N_42180,N_42327);
nand U45138 (N_45138,N_42551,N_43627);
xnor U45139 (N_45139,N_42562,N_43200);
nand U45140 (N_45140,N_43627,N_43891);
nand U45141 (N_45141,N_43496,N_42272);
nor U45142 (N_45142,N_42410,N_42982);
or U45143 (N_45143,N_43086,N_42056);
nor U45144 (N_45144,N_42431,N_43498);
nand U45145 (N_45145,N_43144,N_42462);
and U45146 (N_45146,N_43119,N_42882);
nand U45147 (N_45147,N_42389,N_42854);
and U45148 (N_45148,N_43954,N_43009);
xnor U45149 (N_45149,N_42967,N_43842);
or U45150 (N_45150,N_43903,N_43706);
nor U45151 (N_45151,N_43431,N_42382);
or U45152 (N_45152,N_43533,N_43535);
or U45153 (N_45153,N_43366,N_43908);
nor U45154 (N_45154,N_43597,N_43919);
xnor U45155 (N_45155,N_43651,N_43793);
or U45156 (N_45156,N_42310,N_42184);
nor U45157 (N_45157,N_43532,N_43674);
nor U45158 (N_45158,N_43981,N_42711);
nand U45159 (N_45159,N_42175,N_42705);
nor U45160 (N_45160,N_42480,N_43799);
or U45161 (N_45161,N_43731,N_42383);
nor U45162 (N_45162,N_42233,N_43518);
nor U45163 (N_45163,N_42028,N_42855);
nand U45164 (N_45164,N_43570,N_43107);
or U45165 (N_45165,N_42863,N_42191);
xnor U45166 (N_45166,N_43073,N_43805);
or U45167 (N_45167,N_43618,N_43469);
or U45168 (N_45168,N_42019,N_42374);
nand U45169 (N_45169,N_43853,N_43864);
or U45170 (N_45170,N_42036,N_42950);
nor U45171 (N_45171,N_43689,N_42545);
xor U45172 (N_45172,N_43954,N_42833);
xnor U45173 (N_45173,N_43879,N_43774);
nand U45174 (N_45174,N_43550,N_43373);
nand U45175 (N_45175,N_42915,N_43403);
xor U45176 (N_45176,N_43601,N_43869);
and U45177 (N_45177,N_42621,N_42520);
xor U45178 (N_45178,N_43431,N_43282);
xor U45179 (N_45179,N_43676,N_43103);
or U45180 (N_45180,N_42265,N_43074);
or U45181 (N_45181,N_43599,N_43606);
and U45182 (N_45182,N_43253,N_43335);
or U45183 (N_45183,N_43680,N_42216);
or U45184 (N_45184,N_43789,N_42375);
and U45185 (N_45185,N_42654,N_43045);
or U45186 (N_45186,N_42982,N_42806);
nor U45187 (N_45187,N_42729,N_42519);
xnor U45188 (N_45188,N_43577,N_43315);
nand U45189 (N_45189,N_43630,N_43948);
xnor U45190 (N_45190,N_43554,N_42712);
or U45191 (N_45191,N_42174,N_42372);
xor U45192 (N_45192,N_43659,N_42729);
xnor U45193 (N_45193,N_42508,N_43821);
nor U45194 (N_45194,N_42105,N_42889);
xnor U45195 (N_45195,N_42228,N_43105);
nand U45196 (N_45196,N_43810,N_42510);
or U45197 (N_45197,N_43195,N_42419);
and U45198 (N_45198,N_43236,N_43959);
nor U45199 (N_45199,N_42656,N_42814);
nand U45200 (N_45200,N_42032,N_42584);
nor U45201 (N_45201,N_42835,N_43891);
nand U45202 (N_45202,N_42510,N_42310);
or U45203 (N_45203,N_42532,N_43143);
nand U45204 (N_45204,N_43862,N_42331);
and U45205 (N_45205,N_42993,N_43705);
nor U45206 (N_45206,N_43515,N_42768);
and U45207 (N_45207,N_43035,N_42821);
nand U45208 (N_45208,N_42533,N_42697);
nor U45209 (N_45209,N_43886,N_42825);
xnor U45210 (N_45210,N_42575,N_43076);
nand U45211 (N_45211,N_42331,N_42795);
or U45212 (N_45212,N_43601,N_42816);
or U45213 (N_45213,N_42022,N_42792);
and U45214 (N_45214,N_43174,N_43809);
nor U45215 (N_45215,N_42632,N_42394);
or U45216 (N_45216,N_43761,N_43689);
xnor U45217 (N_45217,N_42730,N_43757);
nand U45218 (N_45218,N_42191,N_43584);
and U45219 (N_45219,N_42411,N_42048);
or U45220 (N_45220,N_43000,N_42967);
nand U45221 (N_45221,N_43680,N_42888);
nor U45222 (N_45222,N_43108,N_42293);
and U45223 (N_45223,N_42653,N_43858);
and U45224 (N_45224,N_42189,N_42872);
nor U45225 (N_45225,N_43032,N_43160);
nor U45226 (N_45226,N_42986,N_43061);
nand U45227 (N_45227,N_43372,N_42847);
nand U45228 (N_45228,N_42897,N_43503);
nand U45229 (N_45229,N_43806,N_42816);
nor U45230 (N_45230,N_43224,N_43356);
nor U45231 (N_45231,N_42664,N_42832);
nor U45232 (N_45232,N_43736,N_42441);
or U45233 (N_45233,N_42813,N_42359);
or U45234 (N_45234,N_43174,N_43558);
nor U45235 (N_45235,N_42020,N_43841);
xnor U45236 (N_45236,N_43620,N_42136);
nor U45237 (N_45237,N_43559,N_42466);
nor U45238 (N_45238,N_43814,N_43433);
xnor U45239 (N_45239,N_42765,N_42145);
or U45240 (N_45240,N_42119,N_43526);
nor U45241 (N_45241,N_42481,N_42844);
or U45242 (N_45242,N_43029,N_43268);
and U45243 (N_45243,N_42974,N_42681);
xor U45244 (N_45244,N_42887,N_43556);
nand U45245 (N_45245,N_43400,N_43953);
and U45246 (N_45246,N_42362,N_42425);
and U45247 (N_45247,N_42233,N_43401);
nor U45248 (N_45248,N_43749,N_42529);
or U45249 (N_45249,N_43712,N_42179);
nor U45250 (N_45250,N_42089,N_42751);
xor U45251 (N_45251,N_43881,N_43741);
and U45252 (N_45252,N_43075,N_43671);
and U45253 (N_45253,N_42881,N_43772);
nand U45254 (N_45254,N_42386,N_43197);
nand U45255 (N_45255,N_43631,N_42463);
nand U45256 (N_45256,N_42266,N_43164);
or U45257 (N_45257,N_42104,N_43821);
xnor U45258 (N_45258,N_43894,N_42455);
or U45259 (N_45259,N_42105,N_43455);
and U45260 (N_45260,N_42499,N_42532);
and U45261 (N_45261,N_43226,N_43646);
or U45262 (N_45262,N_43597,N_43533);
and U45263 (N_45263,N_43888,N_43093);
nor U45264 (N_45264,N_42403,N_42533);
and U45265 (N_45265,N_43982,N_42638);
nor U45266 (N_45266,N_43968,N_43596);
nand U45267 (N_45267,N_42983,N_43287);
and U45268 (N_45268,N_43454,N_43233);
xnor U45269 (N_45269,N_42418,N_43983);
and U45270 (N_45270,N_43581,N_43642);
nor U45271 (N_45271,N_42537,N_42222);
nor U45272 (N_45272,N_42178,N_43436);
nand U45273 (N_45273,N_42470,N_43598);
nor U45274 (N_45274,N_42768,N_42135);
and U45275 (N_45275,N_43494,N_43862);
and U45276 (N_45276,N_42191,N_42632);
and U45277 (N_45277,N_42997,N_43501);
and U45278 (N_45278,N_42038,N_43731);
xor U45279 (N_45279,N_43982,N_43743);
or U45280 (N_45280,N_43073,N_43898);
xnor U45281 (N_45281,N_42021,N_42546);
or U45282 (N_45282,N_43444,N_42881);
or U45283 (N_45283,N_42898,N_42404);
xnor U45284 (N_45284,N_42838,N_42194);
and U45285 (N_45285,N_43033,N_43167);
or U45286 (N_45286,N_42929,N_42406);
and U45287 (N_45287,N_43198,N_43403);
nor U45288 (N_45288,N_43493,N_43454);
or U45289 (N_45289,N_43536,N_42505);
and U45290 (N_45290,N_43424,N_42821);
nor U45291 (N_45291,N_43416,N_43253);
or U45292 (N_45292,N_43734,N_43067);
or U45293 (N_45293,N_43922,N_43813);
nand U45294 (N_45294,N_43880,N_42516);
nor U45295 (N_45295,N_43863,N_43072);
nand U45296 (N_45296,N_42137,N_42524);
xor U45297 (N_45297,N_43375,N_42802);
nor U45298 (N_45298,N_43505,N_43586);
xnor U45299 (N_45299,N_43614,N_42323);
nor U45300 (N_45300,N_43525,N_43638);
and U45301 (N_45301,N_43681,N_43123);
nor U45302 (N_45302,N_42230,N_42519);
nand U45303 (N_45303,N_43324,N_42725);
and U45304 (N_45304,N_43413,N_42167);
or U45305 (N_45305,N_43396,N_42473);
nand U45306 (N_45306,N_43469,N_43413);
or U45307 (N_45307,N_42287,N_43203);
and U45308 (N_45308,N_42038,N_42288);
nand U45309 (N_45309,N_43531,N_43179);
xnor U45310 (N_45310,N_42933,N_43718);
xor U45311 (N_45311,N_43141,N_43077);
nor U45312 (N_45312,N_43972,N_43113);
nand U45313 (N_45313,N_42106,N_42859);
nand U45314 (N_45314,N_42266,N_42831);
xor U45315 (N_45315,N_43601,N_43442);
and U45316 (N_45316,N_43521,N_42027);
and U45317 (N_45317,N_42576,N_43106);
and U45318 (N_45318,N_43595,N_43641);
and U45319 (N_45319,N_43127,N_43710);
nand U45320 (N_45320,N_42104,N_43994);
xor U45321 (N_45321,N_43148,N_43675);
and U45322 (N_45322,N_43889,N_42024);
nand U45323 (N_45323,N_42340,N_43451);
nor U45324 (N_45324,N_43473,N_43878);
and U45325 (N_45325,N_43606,N_42754);
nor U45326 (N_45326,N_43716,N_42390);
nand U45327 (N_45327,N_43843,N_42483);
xnor U45328 (N_45328,N_43110,N_43670);
nor U45329 (N_45329,N_43196,N_42961);
or U45330 (N_45330,N_42735,N_43511);
or U45331 (N_45331,N_42029,N_43389);
nand U45332 (N_45332,N_43239,N_42231);
nor U45333 (N_45333,N_42290,N_43488);
xor U45334 (N_45334,N_43961,N_43741);
or U45335 (N_45335,N_42056,N_42696);
and U45336 (N_45336,N_42329,N_43234);
nor U45337 (N_45337,N_42206,N_43071);
or U45338 (N_45338,N_42459,N_42660);
nor U45339 (N_45339,N_43320,N_43481);
nand U45340 (N_45340,N_43036,N_43626);
or U45341 (N_45341,N_43626,N_43943);
and U45342 (N_45342,N_42848,N_43162);
or U45343 (N_45343,N_43489,N_43173);
nand U45344 (N_45344,N_43145,N_42747);
nand U45345 (N_45345,N_42091,N_43059);
nand U45346 (N_45346,N_42485,N_43239);
nor U45347 (N_45347,N_43364,N_42598);
or U45348 (N_45348,N_43840,N_42207);
xor U45349 (N_45349,N_42659,N_43059);
or U45350 (N_45350,N_43828,N_43424);
and U45351 (N_45351,N_42245,N_42764);
nor U45352 (N_45352,N_42477,N_42262);
nand U45353 (N_45353,N_43556,N_43809);
nand U45354 (N_45354,N_43302,N_42772);
or U45355 (N_45355,N_43748,N_42751);
nor U45356 (N_45356,N_43715,N_42742);
or U45357 (N_45357,N_43191,N_43667);
nand U45358 (N_45358,N_42932,N_43164);
nand U45359 (N_45359,N_43689,N_43115);
xnor U45360 (N_45360,N_42567,N_43474);
nor U45361 (N_45361,N_43901,N_43602);
xnor U45362 (N_45362,N_42471,N_43468);
or U45363 (N_45363,N_43801,N_43245);
xor U45364 (N_45364,N_43774,N_42530);
or U45365 (N_45365,N_43020,N_42631);
or U45366 (N_45366,N_43226,N_43607);
nand U45367 (N_45367,N_42493,N_43132);
xor U45368 (N_45368,N_42454,N_42516);
nand U45369 (N_45369,N_43338,N_43109);
nor U45370 (N_45370,N_42076,N_43102);
xor U45371 (N_45371,N_42495,N_42046);
and U45372 (N_45372,N_43339,N_43277);
nor U45373 (N_45373,N_43827,N_42834);
nor U45374 (N_45374,N_42312,N_42845);
and U45375 (N_45375,N_42050,N_42847);
and U45376 (N_45376,N_43548,N_43322);
xnor U45377 (N_45377,N_43755,N_42096);
nand U45378 (N_45378,N_43717,N_42004);
and U45379 (N_45379,N_42845,N_42038);
nand U45380 (N_45380,N_42621,N_43679);
nor U45381 (N_45381,N_42162,N_43979);
xor U45382 (N_45382,N_42043,N_43773);
or U45383 (N_45383,N_42899,N_42741);
nand U45384 (N_45384,N_43882,N_42569);
nand U45385 (N_45385,N_42751,N_42558);
or U45386 (N_45386,N_43930,N_43072);
xor U45387 (N_45387,N_42222,N_42271);
nor U45388 (N_45388,N_42320,N_42864);
nor U45389 (N_45389,N_42988,N_42283);
xor U45390 (N_45390,N_43686,N_43918);
nand U45391 (N_45391,N_42908,N_43677);
or U45392 (N_45392,N_43159,N_43756);
nand U45393 (N_45393,N_43143,N_42198);
nand U45394 (N_45394,N_42820,N_43070);
and U45395 (N_45395,N_43984,N_42299);
and U45396 (N_45396,N_43741,N_42487);
and U45397 (N_45397,N_43086,N_42371);
nor U45398 (N_45398,N_43694,N_43717);
and U45399 (N_45399,N_42459,N_43297);
nor U45400 (N_45400,N_42521,N_42776);
nand U45401 (N_45401,N_42691,N_42837);
xnor U45402 (N_45402,N_43926,N_42641);
and U45403 (N_45403,N_43207,N_42814);
xor U45404 (N_45404,N_42854,N_42613);
nor U45405 (N_45405,N_43281,N_42493);
xnor U45406 (N_45406,N_43245,N_42363);
xnor U45407 (N_45407,N_43094,N_42312);
or U45408 (N_45408,N_43688,N_42935);
and U45409 (N_45409,N_43683,N_42676);
xnor U45410 (N_45410,N_42889,N_43377);
nor U45411 (N_45411,N_43535,N_43642);
nand U45412 (N_45412,N_43942,N_42738);
xor U45413 (N_45413,N_43587,N_42746);
nand U45414 (N_45414,N_43816,N_43519);
xnor U45415 (N_45415,N_42280,N_43049);
nor U45416 (N_45416,N_42554,N_43234);
or U45417 (N_45417,N_42545,N_42676);
nand U45418 (N_45418,N_43475,N_42480);
nor U45419 (N_45419,N_42307,N_42174);
xor U45420 (N_45420,N_42946,N_43908);
nor U45421 (N_45421,N_42292,N_42842);
nand U45422 (N_45422,N_42061,N_42480);
and U45423 (N_45423,N_42590,N_43366);
nand U45424 (N_45424,N_43609,N_42779);
xor U45425 (N_45425,N_43395,N_43008);
and U45426 (N_45426,N_43995,N_43352);
xor U45427 (N_45427,N_43493,N_42440);
or U45428 (N_45428,N_42851,N_42689);
and U45429 (N_45429,N_43888,N_43865);
nand U45430 (N_45430,N_43513,N_42361);
nand U45431 (N_45431,N_43088,N_43794);
or U45432 (N_45432,N_42826,N_43101);
xor U45433 (N_45433,N_42575,N_42734);
or U45434 (N_45434,N_43902,N_42067);
nor U45435 (N_45435,N_43872,N_43873);
nand U45436 (N_45436,N_43728,N_43369);
and U45437 (N_45437,N_43345,N_43928);
and U45438 (N_45438,N_42027,N_43513);
nor U45439 (N_45439,N_43657,N_42502);
nand U45440 (N_45440,N_43338,N_43849);
xor U45441 (N_45441,N_43621,N_43245);
or U45442 (N_45442,N_43739,N_42034);
or U45443 (N_45443,N_43859,N_42627);
or U45444 (N_45444,N_43138,N_43592);
nor U45445 (N_45445,N_42956,N_43879);
nand U45446 (N_45446,N_42658,N_42527);
or U45447 (N_45447,N_43309,N_43181);
nand U45448 (N_45448,N_43053,N_43995);
and U45449 (N_45449,N_43477,N_42630);
nor U45450 (N_45450,N_43257,N_43643);
nor U45451 (N_45451,N_42603,N_43019);
and U45452 (N_45452,N_43994,N_43337);
nor U45453 (N_45453,N_42236,N_43095);
and U45454 (N_45454,N_42451,N_42419);
nand U45455 (N_45455,N_43232,N_42035);
and U45456 (N_45456,N_42050,N_43087);
nor U45457 (N_45457,N_43280,N_43034);
nand U45458 (N_45458,N_43456,N_43027);
and U45459 (N_45459,N_43401,N_42806);
or U45460 (N_45460,N_43080,N_43155);
nand U45461 (N_45461,N_43798,N_43808);
nor U45462 (N_45462,N_42143,N_42392);
nor U45463 (N_45463,N_42182,N_43196);
nor U45464 (N_45464,N_42906,N_42063);
nor U45465 (N_45465,N_43412,N_43404);
nor U45466 (N_45466,N_42930,N_42626);
nand U45467 (N_45467,N_42434,N_43319);
xnor U45468 (N_45468,N_43583,N_43413);
xor U45469 (N_45469,N_42283,N_43068);
or U45470 (N_45470,N_42934,N_42818);
or U45471 (N_45471,N_42702,N_42575);
and U45472 (N_45472,N_42737,N_42765);
and U45473 (N_45473,N_42280,N_43713);
nand U45474 (N_45474,N_43019,N_43844);
and U45475 (N_45475,N_42659,N_43293);
or U45476 (N_45476,N_43776,N_42937);
or U45477 (N_45477,N_43983,N_43991);
or U45478 (N_45478,N_43506,N_42888);
nor U45479 (N_45479,N_42974,N_42214);
xnor U45480 (N_45480,N_42874,N_42045);
nor U45481 (N_45481,N_42269,N_43863);
nand U45482 (N_45482,N_43216,N_43455);
nor U45483 (N_45483,N_43616,N_42777);
nor U45484 (N_45484,N_43343,N_42132);
nor U45485 (N_45485,N_42810,N_42223);
nand U45486 (N_45486,N_43669,N_42241);
and U45487 (N_45487,N_42792,N_42655);
or U45488 (N_45488,N_43156,N_43680);
and U45489 (N_45489,N_43897,N_43200);
and U45490 (N_45490,N_42092,N_42579);
and U45491 (N_45491,N_43609,N_42856);
nor U45492 (N_45492,N_42296,N_42247);
nor U45493 (N_45493,N_43909,N_43537);
or U45494 (N_45494,N_42038,N_42285);
nand U45495 (N_45495,N_42785,N_42315);
nor U45496 (N_45496,N_42091,N_42845);
and U45497 (N_45497,N_42004,N_43767);
xor U45498 (N_45498,N_42140,N_42619);
nand U45499 (N_45499,N_42888,N_42054);
nor U45500 (N_45500,N_42460,N_43818);
and U45501 (N_45501,N_42344,N_43958);
xor U45502 (N_45502,N_43741,N_42973);
or U45503 (N_45503,N_43271,N_43842);
nor U45504 (N_45504,N_42528,N_43062);
nor U45505 (N_45505,N_43211,N_42294);
nor U45506 (N_45506,N_43503,N_42761);
nor U45507 (N_45507,N_43863,N_43595);
nor U45508 (N_45508,N_42501,N_42698);
nand U45509 (N_45509,N_43836,N_42614);
nor U45510 (N_45510,N_43629,N_43730);
xor U45511 (N_45511,N_42431,N_43607);
xor U45512 (N_45512,N_43868,N_42048);
and U45513 (N_45513,N_43535,N_43221);
nor U45514 (N_45514,N_42839,N_43577);
nor U45515 (N_45515,N_42931,N_43292);
xor U45516 (N_45516,N_43007,N_43283);
nand U45517 (N_45517,N_43769,N_42195);
nor U45518 (N_45518,N_42662,N_42050);
nor U45519 (N_45519,N_42400,N_43896);
nor U45520 (N_45520,N_43219,N_43316);
nor U45521 (N_45521,N_43001,N_43203);
xor U45522 (N_45522,N_42090,N_43354);
nor U45523 (N_45523,N_43578,N_42137);
xnor U45524 (N_45524,N_43822,N_43231);
and U45525 (N_45525,N_43311,N_43757);
nand U45526 (N_45526,N_43514,N_43720);
xnor U45527 (N_45527,N_43347,N_42298);
or U45528 (N_45528,N_43489,N_42738);
nor U45529 (N_45529,N_43176,N_43819);
nor U45530 (N_45530,N_43166,N_42934);
xor U45531 (N_45531,N_43501,N_43935);
nand U45532 (N_45532,N_42735,N_43442);
and U45533 (N_45533,N_43193,N_43898);
nand U45534 (N_45534,N_43893,N_43685);
nand U45535 (N_45535,N_43234,N_43311);
or U45536 (N_45536,N_43122,N_43835);
or U45537 (N_45537,N_42515,N_43936);
nand U45538 (N_45538,N_42316,N_42100);
xor U45539 (N_45539,N_42784,N_42211);
and U45540 (N_45540,N_43393,N_42231);
xnor U45541 (N_45541,N_42135,N_42537);
or U45542 (N_45542,N_42924,N_43058);
xor U45543 (N_45543,N_43524,N_42470);
nand U45544 (N_45544,N_43572,N_43629);
or U45545 (N_45545,N_43287,N_42474);
xnor U45546 (N_45546,N_43776,N_42616);
or U45547 (N_45547,N_42658,N_42310);
or U45548 (N_45548,N_43246,N_42749);
or U45549 (N_45549,N_42484,N_42526);
nor U45550 (N_45550,N_43809,N_43156);
and U45551 (N_45551,N_42885,N_42412);
nor U45552 (N_45552,N_43086,N_43649);
xor U45553 (N_45553,N_43406,N_43572);
and U45554 (N_45554,N_43203,N_42899);
or U45555 (N_45555,N_43012,N_42209);
or U45556 (N_45556,N_42303,N_43959);
xor U45557 (N_45557,N_43669,N_43380);
xnor U45558 (N_45558,N_42995,N_43796);
or U45559 (N_45559,N_42066,N_43705);
and U45560 (N_45560,N_42719,N_42958);
xnor U45561 (N_45561,N_42991,N_43154);
nor U45562 (N_45562,N_43378,N_42306);
nand U45563 (N_45563,N_43971,N_42273);
or U45564 (N_45564,N_42961,N_43871);
xor U45565 (N_45565,N_42518,N_43824);
or U45566 (N_45566,N_42988,N_43340);
or U45567 (N_45567,N_43973,N_42693);
or U45568 (N_45568,N_42006,N_42015);
nand U45569 (N_45569,N_42133,N_42855);
or U45570 (N_45570,N_42918,N_42905);
nand U45571 (N_45571,N_42378,N_43979);
xnor U45572 (N_45572,N_43159,N_42106);
nor U45573 (N_45573,N_43417,N_43375);
nand U45574 (N_45574,N_42220,N_42630);
nor U45575 (N_45575,N_43631,N_43027);
or U45576 (N_45576,N_43250,N_42856);
or U45577 (N_45577,N_43171,N_42885);
or U45578 (N_45578,N_42526,N_42876);
xor U45579 (N_45579,N_43129,N_43305);
and U45580 (N_45580,N_42646,N_43977);
nor U45581 (N_45581,N_43179,N_43422);
nand U45582 (N_45582,N_42213,N_42547);
nand U45583 (N_45583,N_43822,N_42486);
and U45584 (N_45584,N_43928,N_43925);
nor U45585 (N_45585,N_42589,N_43889);
or U45586 (N_45586,N_43756,N_43314);
xnor U45587 (N_45587,N_42980,N_42077);
nand U45588 (N_45588,N_42690,N_42337);
xnor U45589 (N_45589,N_43134,N_42830);
and U45590 (N_45590,N_43732,N_43287);
or U45591 (N_45591,N_42763,N_43315);
nand U45592 (N_45592,N_42318,N_42715);
or U45593 (N_45593,N_42500,N_43297);
and U45594 (N_45594,N_43188,N_43944);
nand U45595 (N_45595,N_43525,N_42929);
xnor U45596 (N_45596,N_42169,N_42768);
and U45597 (N_45597,N_43343,N_42084);
nor U45598 (N_45598,N_42351,N_42993);
nor U45599 (N_45599,N_42166,N_42318);
xnor U45600 (N_45600,N_42485,N_42321);
or U45601 (N_45601,N_43896,N_43778);
and U45602 (N_45602,N_42829,N_43782);
nor U45603 (N_45603,N_42851,N_42761);
nand U45604 (N_45604,N_43219,N_42268);
xor U45605 (N_45605,N_42311,N_43170);
or U45606 (N_45606,N_42275,N_43121);
nand U45607 (N_45607,N_42983,N_42475);
or U45608 (N_45608,N_42587,N_43608);
nand U45609 (N_45609,N_42821,N_42555);
and U45610 (N_45610,N_42468,N_43996);
or U45611 (N_45611,N_43036,N_42578);
and U45612 (N_45612,N_42659,N_43519);
nor U45613 (N_45613,N_43802,N_43926);
or U45614 (N_45614,N_43993,N_43694);
or U45615 (N_45615,N_43923,N_42781);
and U45616 (N_45616,N_43166,N_42822);
nand U45617 (N_45617,N_42734,N_43026);
xnor U45618 (N_45618,N_43330,N_42621);
or U45619 (N_45619,N_42188,N_43872);
nand U45620 (N_45620,N_42652,N_43504);
nor U45621 (N_45621,N_43146,N_43537);
xnor U45622 (N_45622,N_42997,N_42689);
nor U45623 (N_45623,N_42239,N_42248);
nand U45624 (N_45624,N_42152,N_43753);
nand U45625 (N_45625,N_43980,N_42084);
nand U45626 (N_45626,N_42769,N_42800);
xor U45627 (N_45627,N_43670,N_42016);
nand U45628 (N_45628,N_43725,N_42400);
and U45629 (N_45629,N_42108,N_42174);
and U45630 (N_45630,N_42185,N_42418);
xnor U45631 (N_45631,N_43092,N_42084);
nor U45632 (N_45632,N_43085,N_42097);
xor U45633 (N_45633,N_42170,N_42193);
nor U45634 (N_45634,N_43169,N_42094);
nor U45635 (N_45635,N_42694,N_43973);
and U45636 (N_45636,N_42122,N_42319);
xor U45637 (N_45637,N_42194,N_42395);
xnor U45638 (N_45638,N_43517,N_42340);
xnor U45639 (N_45639,N_43784,N_42461);
nor U45640 (N_45640,N_42795,N_43933);
and U45641 (N_45641,N_43835,N_43953);
xor U45642 (N_45642,N_43674,N_43962);
and U45643 (N_45643,N_42450,N_42401);
nand U45644 (N_45644,N_43700,N_42470);
or U45645 (N_45645,N_42700,N_43305);
or U45646 (N_45646,N_42809,N_42004);
xor U45647 (N_45647,N_42724,N_42086);
xnor U45648 (N_45648,N_42741,N_43656);
nand U45649 (N_45649,N_43471,N_43201);
xnor U45650 (N_45650,N_42510,N_43333);
xnor U45651 (N_45651,N_43257,N_43246);
and U45652 (N_45652,N_42652,N_43827);
nor U45653 (N_45653,N_42218,N_43794);
nor U45654 (N_45654,N_42940,N_43244);
or U45655 (N_45655,N_42658,N_42900);
nand U45656 (N_45656,N_42334,N_43699);
and U45657 (N_45657,N_42065,N_42616);
nand U45658 (N_45658,N_43909,N_42817);
and U45659 (N_45659,N_42194,N_43449);
or U45660 (N_45660,N_42765,N_42490);
and U45661 (N_45661,N_42317,N_42572);
nand U45662 (N_45662,N_42962,N_43863);
nand U45663 (N_45663,N_43739,N_43625);
nand U45664 (N_45664,N_42996,N_42970);
and U45665 (N_45665,N_43533,N_43009);
nand U45666 (N_45666,N_43850,N_43848);
and U45667 (N_45667,N_43637,N_42268);
xnor U45668 (N_45668,N_42359,N_42198);
xnor U45669 (N_45669,N_43510,N_42382);
nand U45670 (N_45670,N_43467,N_42317);
and U45671 (N_45671,N_42697,N_42534);
xnor U45672 (N_45672,N_42432,N_43071);
or U45673 (N_45673,N_42887,N_43580);
xor U45674 (N_45674,N_43176,N_43957);
nand U45675 (N_45675,N_42530,N_43472);
nand U45676 (N_45676,N_43360,N_42540);
or U45677 (N_45677,N_43227,N_42004);
xnor U45678 (N_45678,N_43143,N_42184);
nor U45679 (N_45679,N_43048,N_43240);
and U45680 (N_45680,N_42495,N_43422);
nor U45681 (N_45681,N_42550,N_42099);
nand U45682 (N_45682,N_42683,N_42039);
xnor U45683 (N_45683,N_42153,N_43290);
and U45684 (N_45684,N_42834,N_42559);
nand U45685 (N_45685,N_43524,N_42311);
and U45686 (N_45686,N_43935,N_42786);
nor U45687 (N_45687,N_42125,N_42320);
nor U45688 (N_45688,N_43532,N_43597);
xor U45689 (N_45689,N_43335,N_43548);
nor U45690 (N_45690,N_43832,N_43935);
and U45691 (N_45691,N_42616,N_42124);
xnor U45692 (N_45692,N_43349,N_43210);
nor U45693 (N_45693,N_43790,N_43830);
nand U45694 (N_45694,N_43895,N_43453);
nand U45695 (N_45695,N_43279,N_43656);
and U45696 (N_45696,N_42762,N_43569);
and U45697 (N_45697,N_42003,N_43412);
nand U45698 (N_45698,N_42463,N_43284);
xnor U45699 (N_45699,N_42900,N_42547);
nand U45700 (N_45700,N_43505,N_42235);
xor U45701 (N_45701,N_42567,N_43245);
xnor U45702 (N_45702,N_42252,N_42232);
and U45703 (N_45703,N_43100,N_43036);
nand U45704 (N_45704,N_42886,N_43508);
xor U45705 (N_45705,N_43472,N_42372);
nand U45706 (N_45706,N_43983,N_43250);
nor U45707 (N_45707,N_42794,N_43144);
nor U45708 (N_45708,N_43752,N_43262);
nor U45709 (N_45709,N_42618,N_42801);
and U45710 (N_45710,N_43855,N_43242);
xor U45711 (N_45711,N_42980,N_43044);
xnor U45712 (N_45712,N_43546,N_43701);
nor U45713 (N_45713,N_43130,N_42459);
and U45714 (N_45714,N_42252,N_42350);
nor U45715 (N_45715,N_43665,N_42378);
or U45716 (N_45716,N_42743,N_43044);
xnor U45717 (N_45717,N_43443,N_43850);
xor U45718 (N_45718,N_43558,N_42115);
nor U45719 (N_45719,N_42823,N_42180);
xor U45720 (N_45720,N_42374,N_42929);
and U45721 (N_45721,N_42661,N_43632);
and U45722 (N_45722,N_43511,N_42571);
xor U45723 (N_45723,N_42532,N_43271);
or U45724 (N_45724,N_43584,N_43040);
or U45725 (N_45725,N_43820,N_42687);
nand U45726 (N_45726,N_43539,N_43887);
nand U45727 (N_45727,N_43329,N_42750);
xnor U45728 (N_45728,N_42729,N_42616);
nor U45729 (N_45729,N_43850,N_43300);
and U45730 (N_45730,N_43521,N_43359);
and U45731 (N_45731,N_42301,N_42543);
nor U45732 (N_45732,N_42693,N_42154);
or U45733 (N_45733,N_42309,N_42187);
and U45734 (N_45734,N_42251,N_42796);
nand U45735 (N_45735,N_42562,N_42372);
nor U45736 (N_45736,N_42112,N_43747);
nor U45737 (N_45737,N_42849,N_42419);
nand U45738 (N_45738,N_43346,N_42733);
or U45739 (N_45739,N_43118,N_43520);
nor U45740 (N_45740,N_42480,N_43233);
nor U45741 (N_45741,N_42384,N_43506);
and U45742 (N_45742,N_43383,N_43062);
nand U45743 (N_45743,N_42475,N_42347);
nand U45744 (N_45744,N_43507,N_43198);
nor U45745 (N_45745,N_42714,N_42187);
or U45746 (N_45746,N_42185,N_42001);
xor U45747 (N_45747,N_43050,N_43422);
and U45748 (N_45748,N_43328,N_42508);
or U45749 (N_45749,N_43769,N_43906);
xor U45750 (N_45750,N_42496,N_42656);
xnor U45751 (N_45751,N_43265,N_42884);
nand U45752 (N_45752,N_43880,N_43964);
nor U45753 (N_45753,N_42707,N_43411);
or U45754 (N_45754,N_42340,N_42255);
nand U45755 (N_45755,N_43071,N_43551);
and U45756 (N_45756,N_42212,N_42967);
nor U45757 (N_45757,N_43145,N_42631);
xor U45758 (N_45758,N_42034,N_43339);
nor U45759 (N_45759,N_43146,N_42148);
nor U45760 (N_45760,N_43499,N_43554);
and U45761 (N_45761,N_43434,N_43730);
xnor U45762 (N_45762,N_43595,N_42959);
nand U45763 (N_45763,N_43034,N_42607);
nand U45764 (N_45764,N_42410,N_42586);
nand U45765 (N_45765,N_42017,N_42344);
xor U45766 (N_45766,N_42759,N_42725);
or U45767 (N_45767,N_43767,N_42759);
and U45768 (N_45768,N_42850,N_42008);
xnor U45769 (N_45769,N_42021,N_43002);
or U45770 (N_45770,N_43959,N_42456);
nand U45771 (N_45771,N_42727,N_43478);
or U45772 (N_45772,N_43531,N_42880);
nand U45773 (N_45773,N_43087,N_42294);
or U45774 (N_45774,N_43095,N_42227);
xnor U45775 (N_45775,N_43184,N_43612);
or U45776 (N_45776,N_42185,N_43905);
or U45777 (N_45777,N_42257,N_42138);
nor U45778 (N_45778,N_43764,N_42005);
nor U45779 (N_45779,N_43981,N_43947);
nand U45780 (N_45780,N_42164,N_42689);
xor U45781 (N_45781,N_42893,N_43055);
nand U45782 (N_45782,N_43112,N_43877);
or U45783 (N_45783,N_43247,N_42903);
or U45784 (N_45784,N_43842,N_42448);
and U45785 (N_45785,N_43465,N_43673);
nor U45786 (N_45786,N_42665,N_43116);
and U45787 (N_45787,N_43838,N_43108);
xnor U45788 (N_45788,N_43044,N_42202);
and U45789 (N_45789,N_42986,N_43712);
nand U45790 (N_45790,N_43883,N_42002);
nand U45791 (N_45791,N_43208,N_43582);
nor U45792 (N_45792,N_43717,N_43821);
or U45793 (N_45793,N_43903,N_43060);
xor U45794 (N_45794,N_42395,N_42130);
or U45795 (N_45795,N_43151,N_43339);
nor U45796 (N_45796,N_42342,N_43931);
or U45797 (N_45797,N_42113,N_43808);
or U45798 (N_45798,N_42672,N_42696);
and U45799 (N_45799,N_42449,N_42573);
xnor U45800 (N_45800,N_42014,N_43718);
and U45801 (N_45801,N_43775,N_43962);
nor U45802 (N_45802,N_42317,N_43362);
or U45803 (N_45803,N_43409,N_42304);
or U45804 (N_45804,N_43958,N_42240);
xnor U45805 (N_45805,N_42498,N_43138);
nor U45806 (N_45806,N_43418,N_43133);
nor U45807 (N_45807,N_43878,N_43750);
and U45808 (N_45808,N_42053,N_42164);
nor U45809 (N_45809,N_42130,N_42111);
nor U45810 (N_45810,N_42569,N_42678);
nor U45811 (N_45811,N_43355,N_42788);
or U45812 (N_45812,N_42954,N_42679);
nor U45813 (N_45813,N_42559,N_43558);
and U45814 (N_45814,N_43292,N_43029);
nand U45815 (N_45815,N_43012,N_43797);
nor U45816 (N_45816,N_42881,N_43981);
xnor U45817 (N_45817,N_43740,N_43646);
nand U45818 (N_45818,N_43321,N_42832);
nand U45819 (N_45819,N_42898,N_43403);
nand U45820 (N_45820,N_42176,N_43175);
xnor U45821 (N_45821,N_43282,N_42310);
and U45822 (N_45822,N_42715,N_42007);
nand U45823 (N_45823,N_43362,N_43203);
xnor U45824 (N_45824,N_43010,N_42181);
nand U45825 (N_45825,N_42411,N_43811);
and U45826 (N_45826,N_42552,N_43186);
nor U45827 (N_45827,N_43435,N_42740);
xnor U45828 (N_45828,N_42606,N_43356);
nand U45829 (N_45829,N_42574,N_43983);
and U45830 (N_45830,N_43582,N_43385);
nand U45831 (N_45831,N_42602,N_42728);
xnor U45832 (N_45832,N_43790,N_42795);
nand U45833 (N_45833,N_43713,N_43758);
nand U45834 (N_45834,N_42492,N_42456);
and U45835 (N_45835,N_42281,N_43984);
nand U45836 (N_45836,N_43337,N_43562);
or U45837 (N_45837,N_42188,N_43559);
nand U45838 (N_45838,N_42247,N_43858);
nor U45839 (N_45839,N_43829,N_42786);
nand U45840 (N_45840,N_42379,N_42964);
or U45841 (N_45841,N_42162,N_43186);
nand U45842 (N_45842,N_42146,N_43476);
nand U45843 (N_45843,N_42766,N_43574);
nand U45844 (N_45844,N_42921,N_42656);
xnor U45845 (N_45845,N_43025,N_42216);
or U45846 (N_45846,N_42335,N_42160);
nor U45847 (N_45847,N_42428,N_43614);
nand U45848 (N_45848,N_42733,N_43474);
nand U45849 (N_45849,N_43557,N_42436);
nand U45850 (N_45850,N_42569,N_43540);
nand U45851 (N_45851,N_42627,N_43182);
or U45852 (N_45852,N_43231,N_42600);
or U45853 (N_45853,N_42467,N_43834);
nand U45854 (N_45854,N_43071,N_43413);
nor U45855 (N_45855,N_43941,N_42335);
and U45856 (N_45856,N_43835,N_43238);
nand U45857 (N_45857,N_42866,N_43057);
xnor U45858 (N_45858,N_42879,N_42869);
xor U45859 (N_45859,N_42340,N_43646);
xor U45860 (N_45860,N_43795,N_43015);
or U45861 (N_45861,N_43814,N_43981);
nor U45862 (N_45862,N_42441,N_42830);
nor U45863 (N_45863,N_42424,N_42963);
and U45864 (N_45864,N_42998,N_42295);
xor U45865 (N_45865,N_42630,N_43910);
xor U45866 (N_45866,N_42271,N_43268);
and U45867 (N_45867,N_43615,N_42918);
nor U45868 (N_45868,N_42313,N_42697);
xnor U45869 (N_45869,N_42113,N_42606);
xor U45870 (N_45870,N_42202,N_43106);
nor U45871 (N_45871,N_42860,N_43151);
or U45872 (N_45872,N_42035,N_42487);
nor U45873 (N_45873,N_43289,N_43246);
nor U45874 (N_45874,N_42923,N_42538);
nor U45875 (N_45875,N_42598,N_43729);
and U45876 (N_45876,N_43050,N_42245);
or U45877 (N_45877,N_42596,N_43380);
and U45878 (N_45878,N_43161,N_43641);
nand U45879 (N_45879,N_42646,N_43680);
nand U45880 (N_45880,N_42676,N_42965);
or U45881 (N_45881,N_43955,N_43841);
nor U45882 (N_45882,N_42034,N_43427);
and U45883 (N_45883,N_42826,N_43329);
xor U45884 (N_45884,N_43092,N_42386);
nand U45885 (N_45885,N_43950,N_43778);
and U45886 (N_45886,N_42273,N_42506);
nand U45887 (N_45887,N_43081,N_43768);
nor U45888 (N_45888,N_42521,N_42566);
and U45889 (N_45889,N_42426,N_43395);
or U45890 (N_45890,N_43354,N_43077);
nand U45891 (N_45891,N_43501,N_43163);
or U45892 (N_45892,N_42615,N_43178);
and U45893 (N_45893,N_43722,N_43236);
nor U45894 (N_45894,N_42139,N_42320);
nor U45895 (N_45895,N_42427,N_43467);
xnor U45896 (N_45896,N_42587,N_42716);
nand U45897 (N_45897,N_43716,N_43305);
nor U45898 (N_45898,N_43616,N_42265);
or U45899 (N_45899,N_43713,N_42881);
xor U45900 (N_45900,N_43164,N_42865);
nand U45901 (N_45901,N_42026,N_42932);
nand U45902 (N_45902,N_42644,N_42056);
xnor U45903 (N_45903,N_42510,N_43640);
and U45904 (N_45904,N_42843,N_43553);
nand U45905 (N_45905,N_42542,N_43883);
nand U45906 (N_45906,N_42669,N_42962);
nand U45907 (N_45907,N_42168,N_42299);
nor U45908 (N_45908,N_42692,N_43996);
and U45909 (N_45909,N_43347,N_43022);
xnor U45910 (N_45910,N_42718,N_43365);
nor U45911 (N_45911,N_42237,N_43503);
nor U45912 (N_45912,N_42205,N_42276);
and U45913 (N_45913,N_43742,N_43215);
xor U45914 (N_45914,N_42221,N_43574);
xnor U45915 (N_45915,N_42115,N_43398);
xor U45916 (N_45916,N_43061,N_42113);
and U45917 (N_45917,N_43928,N_43711);
nand U45918 (N_45918,N_43572,N_43840);
nand U45919 (N_45919,N_42880,N_42751);
nand U45920 (N_45920,N_42257,N_43422);
xor U45921 (N_45921,N_43342,N_42486);
xor U45922 (N_45922,N_42845,N_43172);
nor U45923 (N_45923,N_43262,N_42086);
and U45924 (N_45924,N_42223,N_43019);
or U45925 (N_45925,N_43408,N_43176);
nor U45926 (N_45926,N_42745,N_43729);
nand U45927 (N_45927,N_42946,N_42806);
and U45928 (N_45928,N_43966,N_43723);
nand U45929 (N_45929,N_43083,N_43708);
and U45930 (N_45930,N_42551,N_42412);
nand U45931 (N_45931,N_43955,N_42283);
nor U45932 (N_45932,N_42447,N_42617);
and U45933 (N_45933,N_43448,N_42329);
and U45934 (N_45934,N_43770,N_43822);
or U45935 (N_45935,N_42715,N_42435);
and U45936 (N_45936,N_42840,N_43664);
nor U45937 (N_45937,N_43216,N_42187);
xnor U45938 (N_45938,N_43523,N_42542);
xnor U45939 (N_45939,N_43003,N_43497);
and U45940 (N_45940,N_43574,N_42300);
xor U45941 (N_45941,N_43392,N_43827);
nand U45942 (N_45942,N_43121,N_43560);
or U45943 (N_45943,N_43281,N_42724);
nor U45944 (N_45944,N_42565,N_43880);
nand U45945 (N_45945,N_43472,N_42511);
nor U45946 (N_45946,N_43469,N_43490);
and U45947 (N_45947,N_43861,N_43944);
nor U45948 (N_45948,N_43368,N_42230);
and U45949 (N_45949,N_43741,N_43450);
and U45950 (N_45950,N_43179,N_42402);
and U45951 (N_45951,N_43045,N_43447);
nor U45952 (N_45952,N_42788,N_42182);
or U45953 (N_45953,N_43467,N_42304);
nor U45954 (N_45954,N_43636,N_43622);
nor U45955 (N_45955,N_43076,N_42251);
nor U45956 (N_45956,N_43733,N_42628);
nor U45957 (N_45957,N_42721,N_43306);
nor U45958 (N_45958,N_42378,N_42191);
nor U45959 (N_45959,N_42066,N_43317);
and U45960 (N_45960,N_43989,N_43003);
nand U45961 (N_45961,N_43238,N_42966);
nand U45962 (N_45962,N_43825,N_42479);
or U45963 (N_45963,N_43960,N_43645);
or U45964 (N_45964,N_43795,N_43554);
nor U45965 (N_45965,N_42323,N_42812);
nand U45966 (N_45966,N_42485,N_43745);
and U45967 (N_45967,N_43981,N_43111);
nand U45968 (N_45968,N_42617,N_42653);
xnor U45969 (N_45969,N_42715,N_42635);
and U45970 (N_45970,N_43873,N_42519);
xnor U45971 (N_45971,N_43952,N_42946);
xnor U45972 (N_45972,N_42657,N_42258);
and U45973 (N_45973,N_42955,N_42392);
nor U45974 (N_45974,N_43897,N_42175);
nor U45975 (N_45975,N_42669,N_43867);
nor U45976 (N_45976,N_43620,N_43269);
nand U45977 (N_45977,N_43412,N_42519);
xor U45978 (N_45978,N_42754,N_42677);
and U45979 (N_45979,N_43213,N_42841);
nand U45980 (N_45980,N_43418,N_43460);
nand U45981 (N_45981,N_43764,N_43185);
and U45982 (N_45982,N_43711,N_42342);
nand U45983 (N_45983,N_43840,N_42900);
xor U45984 (N_45984,N_43930,N_42636);
or U45985 (N_45985,N_43929,N_43777);
nor U45986 (N_45986,N_42037,N_42634);
or U45987 (N_45987,N_42190,N_42044);
xnor U45988 (N_45988,N_42282,N_43337);
and U45989 (N_45989,N_42680,N_42636);
nand U45990 (N_45990,N_42256,N_43104);
or U45991 (N_45991,N_43731,N_43432);
and U45992 (N_45992,N_42444,N_42113);
nand U45993 (N_45993,N_43926,N_43118);
and U45994 (N_45994,N_43524,N_43794);
xnor U45995 (N_45995,N_43523,N_42793);
or U45996 (N_45996,N_43680,N_43724);
or U45997 (N_45997,N_42367,N_43182);
xor U45998 (N_45998,N_42966,N_43408);
nor U45999 (N_45999,N_42548,N_43598);
and U46000 (N_46000,N_45047,N_45844);
nand U46001 (N_46001,N_45258,N_45354);
nand U46002 (N_46002,N_45292,N_45468);
or U46003 (N_46003,N_45841,N_45801);
and U46004 (N_46004,N_45981,N_44543);
nand U46005 (N_46005,N_45315,N_45752);
and U46006 (N_46006,N_45529,N_45026);
nand U46007 (N_46007,N_44456,N_44175);
or U46008 (N_46008,N_45359,N_45308);
or U46009 (N_46009,N_44332,N_44271);
xnor U46010 (N_46010,N_44832,N_44667);
nor U46011 (N_46011,N_45858,N_44459);
nand U46012 (N_46012,N_44468,N_44068);
or U46013 (N_46013,N_44009,N_45902);
or U46014 (N_46014,N_45362,N_45299);
nor U46015 (N_46015,N_45126,N_45073);
xor U46016 (N_46016,N_44631,N_45928);
nor U46017 (N_46017,N_45432,N_45069);
xor U46018 (N_46018,N_45297,N_44433);
xor U46019 (N_46019,N_45358,N_45211);
or U46020 (N_46020,N_44576,N_44732);
xor U46021 (N_46021,N_44041,N_44428);
nand U46022 (N_46022,N_44016,N_44539);
nand U46023 (N_46023,N_44161,N_44300);
xor U46024 (N_46024,N_45685,N_44876);
nor U46025 (N_46025,N_45578,N_44623);
and U46026 (N_46026,N_44387,N_45426);
nor U46027 (N_46027,N_44689,N_44244);
or U46028 (N_46028,N_44642,N_45754);
nor U46029 (N_46029,N_44839,N_44610);
xnor U46030 (N_46030,N_45042,N_45747);
and U46031 (N_46031,N_44299,N_44995);
or U46032 (N_46032,N_44211,N_45443);
and U46033 (N_46033,N_45093,N_45163);
nor U46034 (N_46034,N_45038,N_45753);
or U46035 (N_46035,N_44402,N_45409);
nor U46036 (N_46036,N_45104,N_45484);
or U46037 (N_46037,N_45786,N_45151);
nand U46038 (N_46038,N_45540,N_45001);
xor U46039 (N_46039,N_44403,N_45382);
xor U46040 (N_46040,N_45182,N_44824);
nand U46041 (N_46041,N_44940,N_44635);
or U46042 (N_46042,N_44954,N_45653);
xnor U46043 (N_46043,N_44682,N_45764);
nand U46044 (N_46044,N_44508,N_44024);
and U46045 (N_46045,N_44624,N_44880);
nand U46046 (N_46046,N_45373,N_44987);
nand U46047 (N_46047,N_45614,N_44854);
nand U46048 (N_46048,N_44809,N_45994);
or U46049 (N_46049,N_44498,N_44568);
or U46050 (N_46050,N_45993,N_44182);
nand U46051 (N_46051,N_45652,N_45569);
and U46052 (N_46052,N_44239,N_44149);
and U46053 (N_46053,N_44183,N_45879);
xor U46054 (N_46054,N_44220,N_44385);
nor U46055 (N_46055,N_44895,N_45076);
nor U46056 (N_46056,N_45474,N_45797);
nand U46057 (N_46057,N_45551,N_44168);
or U46058 (N_46058,N_44565,N_44618);
xor U46059 (N_46059,N_44958,N_44890);
and U46060 (N_46060,N_45880,N_45364);
nand U46061 (N_46061,N_45859,N_45554);
or U46062 (N_46062,N_45015,N_45709);
nand U46063 (N_46063,N_45556,N_44503);
nor U46064 (N_46064,N_45559,N_45194);
or U46065 (N_46065,N_45196,N_45787);
xnor U46066 (N_46066,N_45116,N_44362);
xnor U46067 (N_46067,N_44422,N_45264);
nand U46068 (N_46068,N_44959,N_45134);
and U46069 (N_46069,N_45146,N_44946);
and U46070 (N_46070,N_44546,N_44267);
nor U46071 (N_46071,N_44720,N_44556);
nor U46072 (N_46072,N_45465,N_44548);
xor U46073 (N_46073,N_44857,N_45102);
xnor U46074 (N_46074,N_45565,N_44308);
and U46075 (N_46075,N_44103,N_44943);
nand U46076 (N_46076,N_45077,N_44626);
and U46077 (N_46077,N_44098,N_45657);
xnor U46078 (N_46078,N_44821,N_45564);
and U46079 (N_46079,N_45087,N_45715);
or U46080 (N_46080,N_45118,N_44046);
nand U46081 (N_46081,N_45183,N_44006);
nand U46082 (N_46082,N_44401,N_44741);
or U46083 (N_46083,N_45371,N_44935);
nor U46084 (N_46084,N_45226,N_44998);
nand U46085 (N_46085,N_45998,N_45604);
nand U46086 (N_46086,N_44653,N_44996);
and U46087 (N_46087,N_44432,N_45227);
and U46088 (N_46088,N_45717,N_45539);
nand U46089 (N_46089,N_44721,N_45985);
and U46090 (N_46090,N_44101,N_45959);
or U46091 (N_46091,N_44847,N_44658);
xnor U46092 (N_46092,N_44279,N_45602);
nor U46093 (N_46093,N_44289,N_44569);
nand U46094 (N_46094,N_44043,N_44039);
or U46095 (N_46095,N_45473,N_45143);
nand U46096 (N_46096,N_44140,N_45745);
nor U46097 (N_46097,N_44862,N_44894);
and U46098 (N_46098,N_44188,N_45796);
nand U46099 (N_46099,N_45510,N_45321);
nand U46100 (N_46100,N_44481,N_44045);
nand U46101 (N_46101,N_44662,N_44216);
or U46102 (N_46102,N_45004,N_44540);
nand U46103 (N_46103,N_45271,N_44476);
or U46104 (N_46104,N_45930,N_44804);
xor U46105 (N_46105,N_45907,N_44636);
nor U46106 (N_46106,N_45722,N_45255);
or U46107 (N_46107,N_44609,N_45641);
and U46108 (N_46108,N_45275,N_45535);
nand U46109 (N_46109,N_44205,N_44352);
and U46110 (N_46110,N_44163,N_44517);
or U46111 (N_46111,N_44266,N_44097);
nor U46112 (N_46112,N_44315,N_44001);
nand U46113 (N_46113,N_44155,N_44739);
nor U46114 (N_46114,N_45585,N_44888);
or U46115 (N_46115,N_44057,N_44482);
xor U46116 (N_46116,N_44745,N_44709);
xnor U46117 (N_46117,N_45721,N_45220);
nand U46118 (N_46118,N_44458,N_44105);
and U46119 (N_46119,N_45009,N_44889);
and U46120 (N_46120,N_44747,N_45545);
nor U46121 (N_46121,N_45910,N_44474);
xor U46122 (N_46122,N_44694,N_45582);
nor U46123 (N_46123,N_44255,N_45957);
and U46124 (N_46124,N_44632,N_44554);
and U46125 (N_46125,N_44963,N_44107);
nand U46126 (N_46126,N_45562,N_45719);
nand U46127 (N_46127,N_45783,N_44817);
xor U46128 (N_46128,N_44335,N_45405);
nand U46129 (N_46129,N_45702,N_44297);
and U46130 (N_46130,N_45229,N_44965);
or U46131 (N_46131,N_45326,N_44537);
nor U46132 (N_46132,N_45988,N_45932);
xnor U46133 (N_46133,N_45978,N_44675);
or U46134 (N_46134,N_45363,N_45034);
nand U46135 (N_46135,N_44871,N_44264);
and U46136 (N_46136,N_45495,N_45472);
or U46137 (N_46137,N_45131,N_45915);
xor U46138 (N_46138,N_45421,N_45322);
and U46139 (N_46139,N_44766,N_44934);
and U46140 (N_46140,N_44851,N_44671);
xnor U46141 (N_46141,N_45566,N_45658);
and U46142 (N_46142,N_44699,N_44203);
xnor U46143 (N_46143,N_44840,N_44989);
nor U46144 (N_46144,N_45045,N_45272);
nor U46145 (N_46145,N_44716,N_44404);
xnor U46146 (N_46146,N_44598,N_45332);
xor U46147 (N_46147,N_45336,N_44521);
nand U46148 (N_46148,N_45889,N_45068);
or U46149 (N_46149,N_44274,N_45574);
or U46150 (N_46150,N_45014,N_45697);
xnor U46151 (N_46151,N_45725,N_44391);
or U46152 (N_46152,N_44177,N_44859);
and U46153 (N_46153,N_44852,N_45282);
nor U46154 (N_46154,N_45813,N_45804);
xor U46155 (N_46155,N_45238,N_45387);
or U46156 (N_46156,N_45631,N_44535);
nor U46157 (N_46157,N_44110,N_44595);
nor U46158 (N_46158,N_44324,N_44596);
nand U46159 (N_46159,N_44722,N_44286);
or U46160 (N_46160,N_44270,N_45052);
or U46161 (N_46161,N_44676,N_45445);
nor U46162 (N_46162,N_44683,N_45692);
and U46163 (N_46163,N_44415,N_44648);
xnor U46164 (N_46164,N_45485,N_44160);
and U46165 (N_46165,N_45157,N_45313);
nor U46166 (N_46166,N_45541,N_45711);
or U46167 (N_46167,N_45408,N_45412);
and U46168 (N_46168,N_45638,N_44487);
and U46169 (N_46169,N_44158,N_45707);
or U46170 (N_46170,N_45534,N_45145);
nor U46171 (N_46171,N_44520,N_44504);
xor U46172 (N_46172,N_44444,N_44059);
xnor U46173 (N_46173,N_45795,N_45329);
or U46174 (N_46174,N_45028,N_45235);
nor U46175 (N_46175,N_45378,N_44269);
nor U46176 (N_46176,N_45521,N_45938);
xnor U46177 (N_46177,N_44661,N_44639);
or U46178 (N_46178,N_44908,N_44135);
and U46179 (N_46179,N_45953,N_45865);
nand U46180 (N_46180,N_44905,N_44780);
xor U46181 (N_46181,N_45324,N_44020);
or U46182 (N_46182,N_45760,N_45411);
xnor U46183 (N_46183,N_44003,N_44820);
and U46184 (N_46184,N_44597,N_44374);
nand U46185 (N_46185,N_44086,N_44070);
or U46186 (N_46186,N_44583,N_45428);
xnor U46187 (N_46187,N_45463,N_44420);
nand U46188 (N_46188,N_45188,N_45289);
or U46189 (N_46189,N_44261,N_44969);
nand U46190 (N_46190,N_44350,N_45355);
nand U46191 (N_46191,N_44861,N_45856);
or U46192 (N_46192,N_45430,N_44029);
nand U46193 (N_46193,N_45413,N_44828);
nand U46194 (N_46194,N_44717,N_44680);
nor U46195 (N_46195,N_45814,N_44524);
or U46196 (N_46196,N_45690,N_44186);
or U46197 (N_46197,N_44710,N_44621);
or U46198 (N_46198,N_44475,N_45862);
and U46199 (N_46199,N_44552,N_45201);
nand U46200 (N_46200,N_44678,N_44083);
nand U46201 (N_46201,N_45788,N_44955);
nand U46202 (N_46202,N_45759,N_44838);
nor U46203 (N_46203,N_45970,N_45096);
nand U46204 (N_46204,N_45012,N_45972);
or U46205 (N_46205,N_45492,N_44967);
and U46206 (N_46206,N_45509,N_44230);
nand U46207 (N_46207,N_44341,N_45800);
or U46208 (N_46208,N_45245,N_45007);
or U46209 (N_46209,N_44296,N_44509);
nor U46210 (N_46210,N_44902,N_45132);
or U46211 (N_46211,N_44754,N_45518);
and U46212 (N_46212,N_45030,N_44536);
and U46213 (N_46213,N_45058,N_45346);
nor U46214 (N_46214,N_45156,N_45898);
and U46215 (N_46215,N_44263,N_45422);
nor U46216 (N_46216,N_45608,N_45025);
nor U46217 (N_46217,N_45647,N_45961);
or U46218 (N_46218,N_44947,N_45537);
xnor U46219 (N_46219,N_45650,N_45318);
or U46220 (N_46220,N_44223,N_44002);
nor U46221 (N_46221,N_44370,N_45820);
nand U46222 (N_46222,N_44375,N_44591);
or U46223 (N_46223,N_44439,N_44930);
nand U46224 (N_46224,N_44047,N_45388);
nor U46225 (N_46225,N_45607,N_44630);
nand U46226 (N_46226,N_44496,N_45525);
nor U46227 (N_46227,N_45123,N_44891);
and U46228 (N_46228,N_45195,N_45829);
xor U46229 (N_46229,N_45464,N_44976);
and U46230 (N_46230,N_44379,N_44152);
nor U46231 (N_46231,N_45304,N_45016);
or U46232 (N_46232,N_45241,N_44903);
xor U46233 (N_46233,N_45664,N_45746);
nand U46234 (N_46234,N_45875,N_44282);
nand U46235 (N_46235,N_45868,N_44157);
nand U46236 (N_46236,N_44765,N_45057);
nor U46237 (N_46237,N_44073,N_44629);
or U46238 (N_46238,N_44855,N_44613);
xor U46239 (N_46239,N_44421,N_44912);
nand U46240 (N_46240,N_44281,N_45114);
or U46241 (N_46241,N_44752,N_45017);
nor U46242 (N_46242,N_45097,N_45224);
and U46243 (N_46243,N_45153,N_44363);
nand U46244 (N_46244,N_44873,N_44457);
nand U46245 (N_46245,N_45834,N_44663);
xor U46246 (N_46246,N_44793,N_44132);
and U46247 (N_46247,N_45256,N_44376);
or U46248 (N_46248,N_45071,N_44910);
nor U46249 (N_46249,N_45150,N_44392);
nor U46250 (N_46250,N_44711,N_45279);
and U46251 (N_46251,N_44846,N_45298);
xnor U46252 (N_46252,N_44460,N_44849);
and U46253 (N_46253,N_45941,N_45105);
xor U46254 (N_46254,N_44084,N_45266);
or U46255 (N_46255,N_44557,N_44964);
xnor U46256 (N_46256,N_45849,N_45897);
or U46257 (N_46257,N_45637,N_45221);
or U46258 (N_46258,N_45673,N_45398);
nor U46259 (N_46259,N_44283,N_44225);
nand U46260 (N_46260,N_45723,N_45349);
xnor U46261 (N_46261,N_44810,N_45807);
and U46262 (N_46262,N_44397,N_45667);
or U46263 (N_46263,N_45901,N_44365);
xor U46264 (N_46264,N_45418,N_45878);
nand U46265 (N_46265,N_45293,N_44226);
and U46266 (N_46266,N_45505,N_45619);
or U46267 (N_46267,N_45812,N_44449);
nor U46268 (N_46268,N_45103,N_45606);
nand U46269 (N_46269,N_45850,N_44124);
nor U46270 (N_46270,N_45032,N_44147);
and U46271 (N_46271,N_45688,N_45665);
or U46272 (N_46272,N_44681,N_45617);
nor U46273 (N_46273,N_44982,N_44904);
xor U46274 (N_46274,N_45403,N_44842);
nand U46275 (N_46275,N_44767,N_44058);
nor U46276 (N_46276,N_45439,N_44306);
nand U46277 (N_46277,N_44406,N_44075);
nand U46278 (N_46278,N_44151,N_45946);
or U46279 (N_46279,N_45768,N_44394);
nor U46280 (N_46280,N_44833,N_44377);
or U46281 (N_46281,N_45916,N_45138);
nand U46282 (N_46282,N_44398,N_44495);
and U46283 (N_46283,N_45686,N_45496);
or U46284 (N_46284,N_45084,N_45823);
and U46285 (N_46285,N_45700,N_45782);
xor U46286 (N_46286,N_44823,N_45698);
and U46287 (N_46287,N_45228,N_44346);
nand U46288 (N_46288,N_45213,N_45693);
and U46289 (N_46289,N_44069,N_44695);
and U46290 (N_46290,N_44241,N_45461);
or U46291 (N_46291,N_44590,N_45240);
nand U46292 (N_46292,N_45035,N_45695);
xor U46293 (N_46293,N_45740,N_45533);
xor U46294 (N_46294,N_44913,N_44813);
xor U46295 (N_46295,N_44114,N_45863);
xnor U46296 (N_46296,N_45943,N_45416);
and U46297 (N_46297,N_44054,N_45530);
or U46298 (N_46298,N_44237,N_45402);
nand U46299 (N_46299,N_44528,N_44490);
nor U46300 (N_46300,N_44616,N_45733);
xor U46301 (N_46301,N_45599,N_45851);
or U46302 (N_46302,N_45549,N_45254);
nand U46303 (N_46303,N_44939,N_45467);
nor U46304 (N_46304,N_44096,N_45483);
nand U46305 (N_46305,N_45189,N_45864);
or U46306 (N_46306,N_44584,N_44419);
or U46307 (N_46307,N_45605,N_45470);
or U46308 (N_46308,N_44115,N_44423);
or U46309 (N_46309,N_44962,N_45501);
and U46310 (N_46310,N_45542,N_45062);
and U46311 (N_46311,N_44060,N_45049);
xor U46312 (N_46312,N_45805,N_45763);
or U46313 (N_46313,N_45347,N_44483);
and U46314 (N_46314,N_44911,N_44815);
nand U46315 (N_46315,N_44166,N_44215);
xor U46316 (N_46316,N_45497,N_44164);
xnor U46317 (N_46317,N_45632,N_45634);
nand U46318 (N_46318,N_45269,N_44492);
and U46319 (N_46319,N_45059,N_44123);
nor U46320 (N_46320,N_44417,N_44395);
nor U46321 (N_46321,N_44200,N_45724);
or U46322 (N_46322,N_44794,N_44893);
nor U46323 (N_46323,N_44570,N_44950);
or U46324 (N_46324,N_44856,N_44627);
nand U46325 (N_46325,N_44129,N_45645);
or U46326 (N_46326,N_45469,N_45531);
nor U46327 (N_46327,N_44864,N_44664);
nand U46328 (N_46328,N_45216,N_44679);
nand U46329 (N_46329,N_45417,N_45660);
xor U46330 (N_46330,N_44219,N_45333);
xnor U46331 (N_46331,N_45767,N_44272);
nor U46332 (N_46332,N_44858,N_44127);
nor U46333 (N_46333,N_45793,N_44870);
nor U46334 (N_46334,N_44325,N_44562);
nand U46335 (N_46335,N_44302,N_44887);
xor U46336 (N_46336,N_44513,N_44801);
nand U46337 (N_46337,N_44802,N_44280);
nand U46338 (N_46338,N_45450,N_45511);
nor U46339 (N_46339,N_44462,N_44102);
or U46340 (N_46340,N_45615,N_45338);
or U46341 (N_46341,N_44844,N_45583);
or U46342 (N_46342,N_45952,N_44235);
nand U46343 (N_46343,N_45039,N_44882);
nor U46344 (N_46344,N_45586,N_45479);
nand U46345 (N_46345,N_44011,N_45375);
or U46346 (N_46346,N_44900,N_45335);
xor U46347 (N_46347,N_44812,N_45595);
nand U46348 (N_46348,N_44555,N_45169);
and U46349 (N_46349,N_44589,N_44800);
nand U46350 (N_46350,N_45283,N_45185);
xnor U46351 (N_46351,N_44431,N_44309);
xor U46352 (N_46352,N_45506,N_44768);
nor U46353 (N_46353,N_45117,N_45395);
and U46354 (N_46354,N_44000,N_44080);
xor U46355 (N_46355,N_45276,N_45425);
and U46356 (N_46356,N_44799,N_44587);
nand U46357 (N_46357,N_45527,N_44953);
nor U46358 (N_46358,N_44606,N_44090);
or U46359 (N_46359,N_45410,N_45678);
nand U46360 (N_46360,N_45203,N_44727);
or U46361 (N_46361,N_45963,N_45517);
or U46362 (N_46362,N_45011,N_45438);
or U46363 (N_46363,N_44005,N_45260);
and U46364 (N_46364,N_44276,N_44008);
xor U46365 (N_46365,N_44469,N_44577);
xnor U46366 (N_46366,N_44477,N_45817);
nor U46367 (N_46367,N_45307,N_45265);
nor U46368 (N_46368,N_44787,N_44723);
or U46369 (N_46369,N_45681,N_44333);
and U46370 (N_46370,N_45177,N_44329);
or U46371 (N_46371,N_44696,N_45319);
or U46372 (N_46372,N_44668,N_44657);
xor U46373 (N_46373,N_44845,N_45066);
nand U46374 (N_46374,N_45231,N_44227);
xor U46375 (N_46375,N_45656,N_44336);
nor U46376 (N_46376,N_45682,N_44038);
and U46377 (N_46377,N_44049,N_45893);
nor U46378 (N_46378,N_44704,N_45215);
and U46379 (N_46379,N_45340,N_45712);
nor U46380 (N_46380,N_45987,N_44921);
xor U46381 (N_46381,N_45154,N_45852);
xor U46382 (N_46382,N_44410,N_45785);
xor U46383 (N_46383,N_44522,N_44441);
nor U46384 (N_46384,N_44874,N_45158);
xnor U46385 (N_46385,N_44733,N_45662);
nand U46386 (N_46386,N_44715,N_45091);
nor U46387 (N_46387,N_45268,N_45048);
or U46388 (N_46388,N_44085,N_44180);
xor U46389 (N_46389,N_44233,N_44703);
or U46390 (N_46390,N_45186,N_45065);
or U46391 (N_46391,N_44604,N_44748);
or U46392 (N_46392,N_45869,N_44051);
or U46393 (N_46393,N_45120,N_44373);
nor U46394 (N_46394,N_44178,N_45968);
and U46395 (N_46395,N_45573,N_45342);
nor U46396 (N_46396,N_44452,N_44938);
nor U46397 (N_46397,N_44907,N_45935);
xor U46398 (N_46398,N_45598,N_45923);
nand U46399 (N_46399,N_45728,N_44478);
nand U46400 (N_46400,N_44826,N_45022);
or U46401 (N_46401,N_44447,N_45086);
and U46402 (N_46402,N_44254,N_45927);
and U46403 (N_46403,N_45743,N_45137);
or U46404 (N_46404,N_44320,N_44759);
xor U46405 (N_46405,N_45210,N_44351);
and U46406 (N_46406,N_44659,N_44600);
nor U46407 (N_46407,N_44811,N_44510);
xnor U46408 (N_46408,N_44119,N_45589);
nand U46409 (N_46409,N_44927,N_44571);
nor U46410 (N_46410,N_44301,N_44654);
or U46411 (N_46411,N_44637,N_44991);
nand U46412 (N_46412,N_45273,N_45819);
nor U46413 (N_46413,N_44067,N_44055);
nor U46414 (N_46414,N_45029,N_44429);
nand U46415 (N_46415,N_45597,N_44424);
nor U46416 (N_46416,N_45872,N_44295);
nand U46417 (N_46417,N_44789,N_44615);
and U46418 (N_46418,N_45471,N_44651);
nor U46419 (N_46419,N_45085,N_45644);
nor U46420 (N_46420,N_44383,N_45280);
nor U46421 (N_46421,N_44378,N_45591);
nand U46422 (N_46422,N_45951,N_44952);
and U46423 (N_46423,N_45237,N_45334);
or U46424 (N_46424,N_44666,N_45181);
or U46425 (N_46425,N_44652,N_45677);
nand U46426 (N_46426,N_45167,N_45141);
and U46427 (N_46427,N_45899,N_45092);
or U46428 (N_46428,N_45033,N_44511);
xnor U46429 (N_46429,N_44848,N_44757);
nor U46430 (N_46430,N_44121,N_44078);
and U46431 (N_46431,N_45202,N_45661);
or U46432 (N_46432,N_44181,N_45601);
or U46433 (N_46433,N_45791,N_44674);
nor U46434 (N_46434,N_45730,N_45848);
or U46435 (N_46435,N_44172,N_45960);
and U46436 (N_46436,N_44082,N_44247);
or U46437 (N_46437,N_45078,N_45798);
nor U46438 (N_46438,N_44036,N_45672);
nor U46439 (N_46439,N_45088,N_45942);
xor U46440 (N_46440,N_45480,N_45436);
nand U46441 (N_46441,N_44142,N_45734);
xor U46442 (N_46442,N_45703,N_45262);
nand U46443 (N_46443,N_44619,N_45895);
nor U46444 (N_46444,N_44698,N_44560);
xor U46445 (N_46445,N_45995,N_45906);
and U46446 (N_46446,N_45802,N_44707);
or U46447 (N_46447,N_45931,N_45560);
nand U46448 (N_46448,N_44647,N_45587);
xor U46449 (N_46449,N_45152,N_45984);
nand U46450 (N_46450,N_44340,N_44310);
or U46451 (N_46451,N_45792,N_45288);
xor U46452 (N_46452,N_44617,N_45081);
or U46453 (N_46453,N_45552,N_44290);
nand U46454 (N_46454,N_44628,N_45727);
nor U46455 (N_46455,N_45374,N_45002);
and U46456 (N_46456,N_45133,N_44588);
and U46457 (N_46457,N_44742,N_45350);
or U46458 (N_46458,N_45516,N_45311);
and U46459 (N_46459,N_44026,N_44702);
or U46460 (N_46460,N_45553,N_44208);
and U46461 (N_46461,N_45179,N_45175);
nand U46462 (N_46462,N_44023,N_45918);
and U46463 (N_46463,N_45504,N_44240);
nand U46464 (N_46464,N_45381,N_45980);
nand U46465 (N_46465,N_45251,N_44738);
nand U46466 (N_46466,N_44542,N_45287);
nor U46467 (N_46467,N_44897,N_44022);
nor U46468 (N_46468,N_45629,N_45075);
and U46469 (N_46469,N_44735,N_45592);
nor U46470 (N_46470,N_45239,N_45735);
nand U46471 (N_46471,N_44926,N_44516);
or U46472 (N_46472,N_44917,N_45160);
xor U46473 (N_46473,N_45345,N_45544);
and U46474 (N_46474,N_44100,N_45072);
and U46475 (N_46475,N_44686,N_45861);
or U46476 (N_46476,N_44025,N_45018);
nor U46477 (N_46477,N_44829,N_45142);
nand U46478 (N_46478,N_44010,N_45394);
nand U46479 (N_46479,N_45285,N_45380);
xor U46480 (N_46480,N_44892,N_45976);
nand U46481 (N_46481,N_44620,N_45161);
nand U46482 (N_46482,N_44896,N_44430);
nor U46483 (N_46483,N_45838,N_44984);
nor U46484 (N_46484,N_45684,N_45296);
nor U46485 (N_46485,N_44836,N_44945);
nor U46486 (N_46486,N_44104,N_45003);
and U46487 (N_46487,N_44451,N_45036);
or U46488 (N_46488,N_44655,N_44328);
nand U46489 (N_46489,N_45316,N_45666);
xor U46490 (N_46490,N_44924,N_44763);
and U46491 (N_46491,N_45842,N_45128);
nand U46492 (N_46492,N_44956,N_45594);
and U46493 (N_46493,N_45714,N_45140);
and U46494 (N_46494,N_44331,N_44012);
xor U46495 (N_46495,N_45751,N_44563);
nor U46496 (N_46496,N_45546,N_44174);
xnor U46497 (N_46497,N_44355,N_45452);
or U46498 (N_46498,N_44941,N_45323);
nor U46499 (N_46499,N_44293,N_45777);
nor U46500 (N_46500,N_45781,N_45964);
or U46501 (N_46501,N_44827,N_44074);
nor U46502 (N_46502,N_44153,N_45263);
xnor U46503 (N_46503,N_45462,N_44983);
xor U46504 (N_46504,N_45286,N_45441);
nand U46505 (N_46505,N_44322,N_45356);
nand U46506 (N_46506,N_44256,N_44198);
nor U46507 (N_46507,N_44968,N_45873);
xor U46508 (N_46508,N_45309,N_44744);
and U46509 (N_46509,N_45164,N_44063);
nand U46510 (N_46510,N_45616,N_45190);
nand U46511 (N_46511,N_45784,N_45206);
and U46512 (N_46512,N_45500,N_45799);
nand U46513 (N_46513,N_45233,N_45242);
nor U46514 (N_46514,N_45668,N_44176);
xnor U46515 (N_46515,N_44236,N_45571);
or U46516 (N_46516,N_45491,N_44317);
and U46517 (N_46517,N_44712,N_45568);
nor U46518 (N_46518,N_44753,N_44273);
nand U46519 (N_46519,N_44027,N_45572);
nor U46520 (N_46520,N_44450,N_45343);
or U46521 (N_46521,N_44949,N_44017);
xnor U46522 (N_46522,N_45701,N_45639);
and U46523 (N_46523,N_45567,N_44512);
nor U46524 (N_46524,N_45121,N_45089);
nor U46525 (N_46525,N_45729,N_44217);
nor U46526 (N_46526,N_45996,N_44693);
or U46527 (N_46527,N_45070,N_45705);
nor U46528 (N_46528,N_45503,N_45596);
xor U46529 (N_46529,N_45648,N_44381);
xor U46530 (N_46530,N_44126,N_45147);
xnor U46531 (N_46531,N_45737,N_45352);
nand U46532 (N_46532,N_44438,N_44407);
nand U46533 (N_46533,N_44736,N_44971);
nor U46534 (N_46534,N_44783,N_45171);
nor U46535 (N_46535,N_45622,N_45748);
nand U46536 (N_46536,N_44865,N_45810);
and U46537 (N_46537,N_45522,N_45330);
or U46538 (N_46538,N_45561,N_45794);
nor U46539 (N_46539,N_44776,N_44948);
or U46540 (N_46540,N_44412,N_44788);
xnor U46541 (N_46541,N_45611,N_45958);
xor U46542 (N_46542,N_45174,N_44013);
nand U46543 (N_46543,N_45433,N_44734);
and U46544 (N_46544,N_44697,N_45769);
xor U46545 (N_46545,N_44194,N_45027);
xnor U46546 (N_46546,N_44665,N_44463);
nand U46547 (N_46547,N_45204,N_44872);
or U46548 (N_46548,N_44411,N_44034);
xor U46549 (N_46549,N_45144,N_45821);
and U46550 (N_46550,N_45310,N_45041);
xor U46551 (N_46551,N_44670,N_44507);
nor U46552 (N_46552,N_44353,N_44526);
nor U46553 (N_46553,N_44922,N_45259);
nand U46554 (N_46554,N_45172,N_44112);
and U46555 (N_46555,N_45843,N_44344);
and U46556 (N_46556,N_44224,N_45230);
nand U46557 (N_46557,N_45427,N_45905);
xor U46558 (N_46558,N_44396,N_44579);
nand U46559 (N_46559,N_44553,N_45979);
xor U46560 (N_46560,N_45835,N_45043);
nor U46561 (N_46561,N_45939,N_44530);
nand U46562 (N_46562,N_45627,N_44445);
and U46563 (N_46563,N_45393,N_45499);
xor U46564 (N_46564,N_45626,N_45888);
nand U46565 (N_46565,N_45139,N_44756);
xor U46566 (N_46566,N_44692,N_44544);
nand U46567 (N_46567,N_44973,N_45278);
xor U46568 (N_46568,N_44602,N_45543);
nor U46569 (N_46569,N_45588,N_45100);
xor U46570 (N_46570,N_44728,N_45713);
nor U46571 (N_46571,N_45000,N_45919);
nor U46572 (N_46572,N_45687,N_45882);
nor U46573 (N_46573,N_44506,N_44337);
nor U46574 (N_46574,N_45654,N_44660);
xnor U46575 (N_46575,N_44684,N_45399);
xnor U46576 (N_46576,N_44418,N_44349);
xnor U46577 (N_46577,N_45006,N_45366);
nor U46578 (N_46578,N_45921,N_45244);
nor U46579 (N_46579,N_45400,N_44981);
nand U46580 (N_46580,N_45295,N_44050);
or U46581 (N_46581,N_44361,N_44932);
xnor U46582 (N_46582,N_44366,N_45840);
xor U46583 (N_46583,N_44835,N_44467);
xor U46584 (N_46584,N_44388,N_45208);
xor U46585 (N_46585,N_44529,N_44312);
xor U46586 (N_46586,N_44518,N_45633);
nand U46587 (N_46587,N_45325,N_45129);
nor U46588 (N_46588,N_45415,N_44795);
nand U46589 (N_46589,N_44853,N_44822);
nor U46590 (N_46590,N_44586,N_45281);
xor U46591 (N_46591,N_45112,N_45824);
or U46592 (N_46592,N_45610,N_44505);
xnor U46593 (N_46593,N_45205,N_44750);
nand U46594 (N_46594,N_45680,N_45082);
xnor U46595 (N_46595,N_44298,N_44761);
and U46596 (N_46596,N_45977,N_45108);
nor U46597 (N_46597,N_44729,N_45876);
or U46598 (N_46598,N_45447,N_45524);
xnor U46599 (N_46599,N_44081,N_44758);
nand U46600 (N_46600,N_44923,N_44785);
xor U46601 (N_46601,N_45623,N_44204);
xor U46602 (N_46602,N_44534,N_45696);
xor U46603 (N_46603,N_44311,N_44782);
nor U46604 (N_46604,N_44144,N_45482);
and U46605 (N_46605,N_45060,N_44649);
and U46606 (N_46606,N_45947,N_45247);
and U46607 (N_46607,N_44440,N_45811);
xor U46608 (N_46608,N_44928,N_44755);
nand U46609 (N_46609,N_44426,N_44566);
xor U46610 (N_46610,N_44771,N_44162);
or U46611 (N_46611,N_45401,N_45671);
and U46612 (N_46612,N_45222,N_45351);
xnor U46613 (N_46613,N_44901,N_45718);
or U46614 (N_46614,N_45502,N_44106);
and U46615 (N_46615,N_45225,N_44705);
nand U46616 (N_46616,N_45435,N_44749);
and U46617 (N_46617,N_44677,N_44884);
nand U46618 (N_46618,N_44389,N_45762);
or U46619 (N_46619,N_44192,N_45742);
nor U46620 (N_46620,N_44318,N_45954);
xor U46621 (N_46621,N_44869,N_44130);
and U46622 (N_46622,N_44999,N_45446);
nor U46623 (N_46623,N_44564,N_45253);
nor U46624 (N_46624,N_44772,N_44561);
and U46625 (N_46625,N_44139,N_44154);
nand U46626 (N_46626,N_45903,N_45550);
and U46627 (N_46627,N_45050,N_44071);
xnor U46628 (N_46628,N_44357,N_44416);
nand U46629 (N_46629,N_44944,N_44866);
nor U46630 (N_46630,N_45476,N_45618);
and U46631 (N_46631,N_44169,N_45779);
and U46632 (N_46632,N_44867,N_44501);
or U46633 (N_46633,N_45771,N_45187);
and U46634 (N_46634,N_45386,N_44201);
nor U46635 (N_46635,N_45475,N_45494);
xnor U46636 (N_46636,N_45055,N_45317);
xnor U46637 (N_46637,N_44779,N_44714);
nor U46638 (N_46638,N_44493,N_44550);
nor U46639 (N_46639,N_44094,N_44726);
nor U46640 (N_46640,N_44622,N_45391);
or U46641 (N_46641,N_45625,N_45749);
xor U46642 (N_46642,N_45384,N_44035);
nand U46643 (N_46643,N_45414,N_45732);
nand U46644 (N_46644,N_44538,N_45372);
nor U46645 (N_46645,N_45867,N_44248);
nor U46646 (N_46646,N_44138,N_44136);
xnor U46647 (N_46647,N_45538,N_44148);
nor U46648 (N_46648,N_45106,N_44974);
or U46649 (N_46649,N_45054,N_45593);
xor U46650 (N_46650,N_45404,N_44197);
xor U46651 (N_46651,N_45037,N_45178);
and U46652 (N_46652,N_44380,N_44515);
or U46653 (N_46653,N_45095,N_44195);
nand U46654 (N_46654,N_45261,N_45881);
xor U46655 (N_46655,N_44258,N_45955);
and U46656 (N_46656,N_45738,N_44559);
and U46657 (N_46657,N_45920,N_44316);
nand U46658 (N_46658,N_45223,N_45917);
or U46659 (N_46659,N_44128,N_44189);
or U46660 (N_46660,N_44599,N_45830);
xor U46661 (N_46661,N_45064,N_44018);
nor U46662 (N_46662,N_44814,N_44980);
nand U46663 (N_46663,N_45726,N_45115);
or U46664 (N_46664,N_45236,N_44993);
nor U46665 (N_46665,N_44214,N_44488);
or U46666 (N_46666,N_44573,N_45936);
or U46667 (N_46667,N_45967,N_44724);
xor U46668 (N_46668,N_44775,N_44252);
or U46669 (N_46669,N_45890,N_44547);
xnor U46670 (N_46670,N_45997,N_44234);
xnor U46671 (N_46671,N_44218,N_45969);
and U46672 (N_46672,N_44089,N_44284);
or U46673 (N_46673,N_45284,N_44125);
or U46674 (N_46674,N_44358,N_45766);
xnor U46675 (N_46675,N_44713,N_44202);
or U46676 (N_46676,N_45109,N_44480);
nor U46677 (N_46677,N_44545,N_44500);
nor U46678 (N_46678,N_45558,N_45136);
and U46679 (N_46679,N_44919,N_44978);
and U46680 (N_46680,N_44687,N_44770);
or U46681 (N_46681,N_45406,N_44303);
nor U46682 (N_46682,N_45248,N_45294);
xnor U46683 (N_46683,N_44405,N_45217);
nor U46684 (N_46684,N_45192,N_44260);
nand U46685 (N_46685,N_45130,N_45111);
xnor U46686 (N_46686,N_45305,N_45520);
nand U46687 (N_46687,N_45214,N_44572);
xnor U46688 (N_46688,N_45808,N_44253);
or U46689 (N_46689,N_44243,N_45377);
xnor U46690 (N_46690,N_45514,N_45983);
nor U46691 (N_46691,N_44525,N_44485);
or U46692 (N_46692,N_44933,N_44193);
and U46693 (N_46693,N_45456,N_44957);
or U46694 (N_46694,N_45212,N_45512);
xnor U46695 (N_46695,N_44109,N_44133);
nand U46696 (N_46696,N_45871,N_44425);
nor U46697 (N_46697,N_44443,N_44931);
or U46698 (N_46698,N_45699,N_45563);
nand U46699 (N_46699,N_44486,N_45790);
and U46700 (N_46700,N_45973,N_44936);
and U46701 (N_46701,N_44951,N_44831);
nand U46702 (N_46702,N_44608,N_45389);
or U46703 (N_46703,N_44997,N_45392);
and U46704 (N_46704,N_44708,N_44778);
nand U46705 (N_46705,N_45945,N_44134);
and U46706 (N_46706,N_44614,N_45337);
and U46707 (N_46707,N_45803,N_44499);
xnor U46708 (N_46708,N_44131,N_44095);
or U46709 (N_46709,N_45098,N_45679);
nor U46710 (N_46710,N_44918,N_44899);
nor U46711 (N_46711,N_44268,N_45736);
or U46712 (N_46712,N_45925,N_44141);
nand U46713 (N_46713,N_45061,N_45368);
nand U46714 (N_46714,N_45451,N_45420);
xnor U46715 (N_46715,N_44287,N_44464);
nand U46716 (N_46716,N_44228,N_44818);
nand U46717 (N_46717,N_44929,N_44914);
and U46718 (N_46718,N_44338,N_44156);
and U46719 (N_46719,N_45816,N_45080);
and U46720 (N_46720,N_44808,N_44323);
and U46721 (N_46721,N_45755,N_44120);
and U46722 (N_46722,N_44850,N_44021);
nand U46723 (N_46723,N_44251,N_44093);
or U46724 (N_46724,N_45353,N_44731);
xnor U46725 (N_46725,N_44972,N_44145);
nand U46726 (N_46726,N_44209,N_44040);
or U46727 (N_46727,N_44033,N_44582);
xor U46728 (N_46728,N_45466,N_44327);
and U46729 (N_46729,N_45191,N_44718);
or U46730 (N_46730,N_44605,N_45860);
xnor U46731 (N_46731,N_44278,N_45312);
or U46732 (N_46732,N_45756,N_45886);
nand U46733 (N_46733,N_45434,N_45600);
nor U46734 (N_46734,N_44691,N_45040);
nand U46735 (N_46735,N_44446,N_45590);
xor U46736 (N_46736,N_44465,N_44643);
and U46737 (N_46737,N_44685,N_44603);
xnor U46738 (N_46738,N_45828,N_44196);
or U46739 (N_46739,N_45376,N_45458);
or U46740 (N_46740,N_44640,N_45706);
nor U46741 (N_46741,N_45933,N_45663);
nand U46742 (N_46742,N_45770,N_44916);
xor U46743 (N_46743,N_44436,N_45148);
nand U46744 (N_46744,N_45303,N_44232);
and U46745 (N_46745,N_45857,N_44399);
and U46746 (N_46746,N_45519,N_44004);
and U46747 (N_46747,N_45739,N_44805);
or U46748 (N_46748,N_45646,N_44898);
or U46749 (N_46749,N_44343,N_44612);
or U46750 (N_46750,N_44199,N_44032);
or U46751 (N_46751,N_45490,N_45489);
and U46752 (N_46752,N_45162,N_45455);
or U46753 (N_46753,N_45053,N_45971);
nor U46754 (N_46754,N_44334,N_44088);
xnor U46755 (N_46755,N_44920,N_44065);
and U46756 (N_46756,N_44113,N_44798);
nor U46757 (N_46757,N_44633,N_44014);
and U46758 (N_46758,N_45900,N_45581);
or U46759 (N_46759,N_44091,N_44356);
and U46760 (N_46760,N_44641,N_45635);
nor U46761 (N_46761,N_45498,N_45370);
nand U46762 (N_46762,N_44825,N_44245);
and U46763 (N_46763,N_44185,N_45159);
nand U46764 (N_46764,N_44259,N_45385);
and U46765 (N_46765,N_45710,N_44994);
nand U46766 (N_46766,N_44593,N_44786);
nor U46767 (N_46767,N_44191,N_45246);
and U46768 (N_46768,N_45676,N_44184);
nand U46769 (N_46769,N_45365,N_44435);
and U46770 (N_46770,N_45383,N_45827);
and U46771 (N_46771,N_45234,N_44672);
or U46772 (N_46772,N_45570,N_45990);
or U46773 (N_46773,N_45277,N_44167);
and U46774 (N_46774,N_44673,N_44764);
xor U46775 (N_46775,N_44807,N_45847);
nand U46776 (N_46776,N_45965,N_44171);
nand U46777 (N_46777,N_45328,N_44179);
nand U46778 (N_46778,N_44489,N_44531);
nor U46779 (N_46779,N_45986,N_45833);
nand U46780 (N_46780,N_45523,N_45119);
and U46781 (N_46781,N_44885,N_44937);
and U46782 (N_46782,N_44250,N_45674);
xor U46783 (N_46783,N_45507,N_45270);
nor U46784 (N_46784,N_44210,N_44368);
or U46785 (N_46785,N_44883,N_45584);
or U46786 (N_46786,N_45122,N_45008);
or U46787 (N_46787,N_44372,N_45962);
xor U46788 (N_46788,N_44288,N_44257);
or U46789 (N_46789,N_44030,N_45642);
xor U46790 (N_46790,N_45839,N_45621);
nand U46791 (N_46791,N_45005,N_45577);
xor U46792 (N_46792,N_44117,N_44644);
nand U46793 (N_46793,N_44567,N_45176);
nand U46794 (N_46794,N_45110,N_45170);
xnor U46795 (N_46795,N_44277,N_44961);
and U46796 (N_46796,N_45765,N_44986);
nor U46797 (N_46797,N_44330,N_44393);
nor U46798 (N_46798,N_45640,N_45643);
nand U46799 (N_46799,N_44108,N_45090);
xnor U46800 (N_46800,N_44915,N_45010);
nor U46801 (N_46801,N_45716,N_45854);
xor U46802 (N_46802,N_45896,N_44367);
or U46803 (N_46803,N_44792,N_44578);
and U46804 (N_46804,N_44345,N_44737);
or U46805 (N_46805,N_44427,N_45846);
or U46806 (N_46806,N_45826,N_44574);
xor U46807 (N_46807,N_45870,N_44796);
and U46808 (N_46808,N_45778,N_45892);
nor U46809 (N_46809,N_45348,N_45885);
nor U46810 (N_46810,N_44549,N_45515);
nor U46811 (N_46811,N_44137,N_44111);
nand U46812 (N_46812,N_44056,N_44719);
and U46813 (N_46813,N_44294,N_45776);
nand U46814 (N_46814,N_44830,N_44453);
xnor U46815 (N_46815,N_44066,N_44491);
nor U46816 (N_46816,N_45630,N_44238);
xnor U46817 (N_46817,N_45331,N_45548);
or U46818 (N_46818,N_44730,N_45825);
or U46819 (N_46819,N_44988,N_44502);
and U46820 (N_46820,N_45481,N_44292);
nand U46821 (N_46821,N_44307,N_45675);
or U46822 (N_46822,N_45950,N_45780);
and U46823 (N_46823,N_45866,N_45020);
and U46824 (N_46824,N_45099,N_45478);
nor U46825 (N_46825,N_45831,N_44650);
nor U46826 (N_46826,N_45135,N_45051);
xnor U46827 (N_46827,N_45757,N_45982);
nand U46828 (N_46828,N_45291,N_45855);
nand U46829 (N_46829,N_45419,N_44455);
or U46830 (N_46830,N_44669,N_44360);
or U46831 (N_46831,N_45891,N_44860);
or U46832 (N_46832,N_45199,N_44925);
nor U46833 (N_46833,N_45532,N_44448);
nand U46834 (N_46834,N_44688,N_44601);
nor U46835 (N_46835,N_44077,N_44314);
nor U46836 (N_46836,N_45290,N_44774);
xor U46837 (N_46837,N_44769,N_44146);
or U46838 (N_46838,N_44841,N_45576);
nand U46839 (N_46839,N_45024,N_45536);
xnor U46840 (N_46840,N_44053,N_45320);
nand U46841 (N_46841,N_44408,N_44992);
nor U46842 (N_46842,N_45689,N_45603);
nand U46843 (N_46843,N_44581,N_44881);
and U46844 (N_46844,N_45575,N_44863);
nor U46845 (N_46845,N_44028,N_44305);
nand U46846 (N_46846,N_44690,N_44472);
xor U46847 (N_46847,N_45056,N_45929);
nor U46848 (N_46848,N_45944,N_44347);
nand U46849 (N_46849,N_44580,N_45197);
and U46850 (N_46850,N_44514,N_45877);
nand U46851 (N_46851,N_45360,N_44611);
or U46852 (N_46852,N_45079,N_45218);
nand U46853 (N_46853,N_45314,N_45390);
or U46854 (N_46854,N_45429,N_44592);
nor U46855 (N_46855,N_45613,N_44414);
or U46856 (N_46856,N_44118,N_45442);
xor U46857 (N_46857,N_44242,N_44625);
xor U46858 (N_46858,N_45669,N_44190);
or U46859 (N_46859,N_45486,N_44523);
nand U46860 (N_46860,N_45708,N_45367);
nand U46861 (N_46861,N_44371,N_45651);
nand U46862 (N_46862,N_45620,N_44646);
xnor U46863 (N_46863,N_44837,N_44879);
nand U46864 (N_46864,N_44076,N_44048);
xor U46865 (N_46865,N_44222,N_44473);
nor U46866 (N_46866,N_45200,N_44409);
or U46867 (N_46867,N_44816,N_45926);
nand U46868 (N_46868,N_44634,N_45243);
nand U46869 (N_46869,N_45845,N_45019);
or U46870 (N_46870,N_44942,N_45125);
nor U46871 (N_46871,N_44313,N_44221);
or U46872 (N_46872,N_44843,N_45021);
nand U46873 (N_46873,N_44497,N_44834);
nand U46874 (N_46874,N_45547,N_45909);
or U46875 (N_46875,N_45636,N_44784);
nand U46876 (N_46876,N_45219,N_45252);
nand U46877 (N_46877,N_44173,N_45911);
and U46878 (N_46878,N_44743,N_45437);
or U46879 (N_46879,N_45992,N_45063);
and U46880 (N_46880,N_45720,N_45369);
or U46881 (N_46881,N_45339,N_45773);
xnor U46882 (N_46882,N_45913,N_44638);
nand U46883 (N_46883,N_45853,N_45956);
xnor U46884 (N_46884,N_44906,N_45460);
or U46885 (N_46885,N_45449,N_45249);
or U46886 (N_46886,N_44803,N_44558);
or U46887 (N_46887,N_45774,N_44479);
nand U46888 (N_46888,N_45274,N_45232);
xnor U46889 (N_46889,N_45628,N_44092);
or U46890 (N_46890,N_44212,N_45127);
xor U46891 (N_46891,N_44037,N_44087);
or U46892 (N_46892,N_45173,N_45612);
and U46893 (N_46893,N_45257,N_45966);
nand U46894 (N_46894,N_44400,N_45609);
and U46895 (N_46895,N_45444,N_45423);
xor U46896 (N_46896,N_45894,N_44231);
nor U46897 (N_46897,N_44868,N_45508);
and U46898 (N_46898,N_45887,N_44434);
and U46899 (N_46899,N_44527,N_45193);
nor U46900 (N_46900,N_45691,N_44979);
and U46901 (N_46901,N_44585,N_45327);
nor U46902 (N_46902,N_45198,N_45624);
and U46903 (N_46903,N_45761,N_44806);
xnor U46904 (N_46904,N_44015,N_44706);
or U46905 (N_46905,N_44072,N_45528);
nand U46906 (N_46906,N_45731,N_45883);
xnor U46907 (N_46907,N_44390,N_44275);
or U46908 (N_46908,N_44575,N_45083);
or U46909 (N_46909,N_44249,N_44533);
nand U46910 (N_46910,N_44773,N_44369);
xor U46911 (N_46911,N_44007,N_44985);
and U46912 (N_46912,N_44760,N_44791);
and U46913 (N_46913,N_44607,N_45013);
or U46914 (N_46914,N_45649,N_45836);
nand U46915 (N_46915,N_44326,N_45526);
nand U46916 (N_46916,N_45357,N_44645);
nor U46917 (N_46917,N_45046,N_44165);
nand U46918 (N_46918,N_45044,N_45694);
nor U46919 (N_46919,N_44019,N_44437);
nand U46920 (N_46920,N_44229,N_45991);
nand U46921 (N_46921,N_44116,N_45555);
xnor U46922 (N_46922,N_45579,N_44339);
or U46923 (N_46923,N_44384,N_45758);
nand U46924 (N_46924,N_44413,N_45165);
nand U46925 (N_46925,N_45975,N_45884);
nand U46926 (N_46926,N_45750,N_44061);
nor U46927 (N_46927,N_45300,N_45934);
or U46928 (N_46928,N_44990,N_45937);
nor U46929 (N_46929,N_44790,N_45124);
and U46930 (N_46930,N_44354,N_44960);
nand U46931 (N_46931,N_44143,N_45459);
or U46932 (N_46932,N_45301,N_45670);
nand U46933 (N_46933,N_45306,N_44725);
xnor U46934 (N_46934,N_45815,N_44454);
xor U46935 (N_46935,N_45023,N_45659);
nand U46936 (N_46936,N_44656,N_45922);
and U46937 (N_46937,N_45180,N_45457);
nor U46938 (N_46938,N_44762,N_44285);
and U46939 (N_46939,N_44207,N_45487);
nor U46940 (N_46940,N_45809,N_44304);
nand U46941 (N_46941,N_44150,N_44246);
nand U46942 (N_46942,N_45341,N_45914);
and U46943 (N_46943,N_44159,N_44265);
nor U46944 (N_46944,N_45741,N_45772);
or U46945 (N_46945,N_44966,N_44213);
nor U46946 (N_46946,N_45396,N_45440);
or U46947 (N_46947,N_45454,N_44291);
nor U46948 (N_46948,N_44977,N_45074);
xnor U46949 (N_46949,N_45775,N_45113);
xor U46950 (N_46950,N_44364,N_44122);
xor U46951 (N_46951,N_44170,N_45557);
or U46952 (N_46952,N_45267,N_45949);
nor U46953 (N_46953,N_44875,N_44359);
nand U46954 (N_46954,N_45067,N_44042);
nor U46955 (N_46955,N_45149,N_44909);
or U46956 (N_46956,N_44519,N_44442);
or U46957 (N_46957,N_44494,N_44466);
xnor U46958 (N_46958,N_45453,N_45904);
xor U46959 (N_46959,N_44819,N_45806);
or U46960 (N_46960,N_45209,N_45513);
xor U46961 (N_46961,N_45908,N_44342);
xnor U46962 (N_46962,N_45207,N_45999);
or U46963 (N_46963,N_45107,N_45302);
and U46964 (N_46964,N_45818,N_44319);
nand U46965 (N_46965,N_44262,N_44461);
and U46966 (N_46966,N_44062,N_45168);
xor U46967 (N_46967,N_44541,N_45431);
nor U46968 (N_46968,N_44064,N_45655);
nor U46969 (N_46969,N_45683,N_45822);
or U46970 (N_46970,N_45397,N_44484);
and U46971 (N_46971,N_44079,N_45912);
xor U46972 (N_46972,N_45744,N_44206);
and U46973 (N_46973,N_44700,N_44751);
and U46974 (N_46974,N_45924,N_45974);
nand U46975 (N_46975,N_44187,N_44740);
nand U46976 (N_46976,N_44551,N_44321);
nor U46977 (N_46977,N_45031,N_44382);
or U46978 (N_46978,N_44878,N_45407);
xnor U46979 (N_46979,N_45344,N_45477);
xor U46980 (N_46980,N_45184,N_44052);
nand U46981 (N_46981,N_44781,N_44975);
and U46982 (N_46982,N_44044,N_45837);
nor U46983 (N_46983,N_45101,N_44701);
and U46984 (N_46984,N_45832,N_44594);
nand U46985 (N_46985,N_45948,N_45424);
xor U46986 (N_46986,N_44746,N_45704);
nand U46987 (N_46987,N_44470,N_45488);
nand U46988 (N_46988,N_45250,N_44877);
nand U46989 (N_46989,N_45361,N_44970);
nand U46990 (N_46990,N_44777,N_45448);
or U46991 (N_46991,N_44886,N_45379);
and U46992 (N_46992,N_44099,N_44031);
or U46993 (N_46993,N_45493,N_45094);
xnor U46994 (N_46994,N_45874,N_44386);
xor U46995 (N_46995,N_45580,N_45989);
and U46996 (N_46996,N_44532,N_45789);
nand U46997 (N_46997,N_45940,N_44471);
xor U46998 (N_46998,N_44348,N_45166);
nand U46999 (N_46999,N_45155,N_44797);
nand U47000 (N_47000,N_45357,N_45663);
or U47001 (N_47001,N_44659,N_44451);
nand U47002 (N_47002,N_45068,N_44438);
and U47003 (N_47003,N_45584,N_44995);
and U47004 (N_47004,N_45668,N_44138);
xor U47005 (N_47005,N_45593,N_45760);
nor U47006 (N_47006,N_45615,N_44747);
xor U47007 (N_47007,N_44822,N_44555);
xor U47008 (N_47008,N_44795,N_44407);
or U47009 (N_47009,N_44370,N_45562);
and U47010 (N_47010,N_45806,N_45793);
nor U47011 (N_47011,N_45713,N_45897);
nor U47012 (N_47012,N_44904,N_45699);
nand U47013 (N_47013,N_45516,N_44040);
nor U47014 (N_47014,N_44942,N_44185);
nand U47015 (N_47015,N_45269,N_44131);
nand U47016 (N_47016,N_45444,N_45219);
nor U47017 (N_47017,N_45433,N_45590);
nand U47018 (N_47018,N_44409,N_45279);
nand U47019 (N_47019,N_44714,N_45320);
or U47020 (N_47020,N_45018,N_45242);
nand U47021 (N_47021,N_45364,N_45202);
or U47022 (N_47022,N_45079,N_44431);
or U47023 (N_47023,N_45214,N_44895);
xor U47024 (N_47024,N_44126,N_45405);
nor U47025 (N_47025,N_44744,N_45993);
nor U47026 (N_47026,N_44242,N_45488);
xor U47027 (N_47027,N_44587,N_44343);
nand U47028 (N_47028,N_45500,N_45120);
and U47029 (N_47029,N_45576,N_44755);
and U47030 (N_47030,N_44049,N_44837);
or U47031 (N_47031,N_45139,N_44014);
nand U47032 (N_47032,N_44318,N_44771);
or U47033 (N_47033,N_45425,N_44683);
nor U47034 (N_47034,N_45009,N_44746);
nand U47035 (N_47035,N_45288,N_45556);
xor U47036 (N_47036,N_44829,N_44921);
xor U47037 (N_47037,N_44895,N_44766);
nor U47038 (N_47038,N_44870,N_45981);
or U47039 (N_47039,N_44840,N_45727);
nand U47040 (N_47040,N_45021,N_44331);
nand U47041 (N_47041,N_44288,N_44095);
or U47042 (N_47042,N_45535,N_45208);
and U47043 (N_47043,N_45413,N_45753);
nand U47044 (N_47044,N_45767,N_44439);
nand U47045 (N_47045,N_44535,N_44777);
nand U47046 (N_47046,N_45260,N_45483);
xnor U47047 (N_47047,N_45100,N_44958);
nand U47048 (N_47048,N_44477,N_45829);
nand U47049 (N_47049,N_44652,N_45625);
nor U47050 (N_47050,N_44027,N_45679);
and U47051 (N_47051,N_45164,N_45112);
and U47052 (N_47052,N_44002,N_44989);
nand U47053 (N_47053,N_44968,N_44585);
nand U47054 (N_47054,N_44640,N_45750);
nor U47055 (N_47055,N_44854,N_45692);
or U47056 (N_47056,N_45644,N_45722);
nor U47057 (N_47057,N_45432,N_44404);
or U47058 (N_47058,N_45515,N_44572);
nor U47059 (N_47059,N_44681,N_45912);
and U47060 (N_47060,N_44285,N_45768);
nor U47061 (N_47061,N_44446,N_45253);
or U47062 (N_47062,N_44738,N_45763);
nor U47063 (N_47063,N_44868,N_44108);
nor U47064 (N_47064,N_45962,N_45576);
xor U47065 (N_47065,N_44794,N_45020);
nor U47066 (N_47066,N_45838,N_45767);
nand U47067 (N_47067,N_45598,N_44176);
nor U47068 (N_47068,N_44565,N_44236);
nand U47069 (N_47069,N_44899,N_44615);
nor U47070 (N_47070,N_45210,N_45021);
xor U47071 (N_47071,N_45249,N_45950);
nand U47072 (N_47072,N_45478,N_44376);
xnor U47073 (N_47073,N_44105,N_45677);
nand U47074 (N_47074,N_44256,N_44203);
nand U47075 (N_47075,N_45932,N_44834);
and U47076 (N_47076,N_44405,N_45388);
nor U47077 (N_47077,N_45607,N_45499);
nor U47078 (N_47078,N_44660,N_44186);
nor U47079 (N_47079,N_44695,N_45534);
and U47080 (N_47080,N_44236,N_45208);
or U47081 (N_47081,N_45862,N_44004);
or U47082 (N_47082,N_45771,N_45991);
nor U47083 (N_47083,N_44288,N_45205);
and U47084 (N_47084,N_44030,N_44529);
and U47085 (N_47085,N_45502,N_45405);
or U47086 (N_47086,N_45543,N_45718);
nor U47087 (N_47087,N_45161,N_45120);
or U47088 (N_47088,N_45747,N_44108);
xor U47089 (N_47089,N_44806,N_44610);
xnor U47090 (N_47090,N_44448,N_44524);
xnor U47091 (N_47091,N_45695,N_45397);
and U47092 (N_47092,N_44237,N_44499);
or U47093 (N_47093,N_44726,N_45146);
xnor U47094 (N_47094,N_45316,N_44752);
or U47095 (N_47095,N_45714,N_44590);
or U47096 (N_47096,N_45486,N_44619);
and U47097 (N_47097,N_45330,N_44334);
nand U47098 (N_47098,N_44687,N_45170);
and U47099 (N_47099,N_45285,N_44578);
nand U47100 (N_47100,N_44201,N_45641);
nor U47101 (N_47101,N_45340,N_45715);
or U47102 (N_47102,N_44809,N_45175);
or U47103 (N_47103,N_45767,N_45116);
nand U47104 (N_47104,N_44931,N_44625);
nor U47105 (N_47105,N_44000,N_45699);
nand U47106 (N_47106,N_44718,N_45270);
nor U47107 (N_47107,N_45246,N_45577);
or U47108 (N_47108,N_44954,N_45926);
and U47109 (N_47109,N_45079,N_44032);
nor U47110 (N_47110,N_44988,N_44802);
xor U47111 (N_47111,N_45086,N_45355);
xor U47112 (N_47112,N_44664,N_45378);
nor U47113 (N_47113,N_45936,N_45420);
xor U47114 (N_47114,N_45901,N_45532);
nand U47115 (N_47115,N_45081,N_44995);
nor U47116 (N_47116,N_45509,N_44842);
and U47117 (N_47117,N_44805,N_44534);
and U47118 (N_47118,N_45677,N_45974);
xnor U47119 (N_47119,N_45998,N_45011);
or U47120 (N_47120,N_44363,N_45332);
xor U47121 (N_47121,N_44309,N_44644);
nor U47122 (N_47122,N_45984,N_44528);
nor U47123 (N_47123,N_44740,N_45243);
nand U47124 (N_47124,N_44152,N_45582);
and U47125 (N_47125,N_44420,N_44213);
nor U47126 (N_47126,N_45775,N_45406);
or U47127 (N_47127,N_45388,N_44167);
and U47128 (N_47128,N_45811,N_44068);
or U47129 (N_47129,N_44888,N_44396);
xor U47130 (N_47130,N_44860,N_45869);
or U47131 (N_47131,N_45180,N_44415);
nand U47132 (N_47132,N_45940,N_45275);
nor U47133 (N_47133,N_45030,N_45666);
or U47134 (N_47134,N_44851,N_45252);
or U47135 (N_47135,N_44587,N_45991);
or U47136 (N_47136,N_45325,N_44891);
nand U47137 (N_47137,N_45220,N_44920);
or U47138 (N_47138,N_45978,N_44156);
or U47139 (N_47139,N_44113,N_45069);
nand U47140 (N_47140,N_45139,N_45081);
nand U47141 (N_47141,N_45115,N_45796);
xnor U47142 (N_47142,N_44268,N_45358);
nand U47143 (N_47143,N_45363,N_44985);
xor U47144 (N_47144,N_45494,N_45530);
or U47145 (N_47145,N_44298,N_44528);
nor U47146 (N_47146,N_45589,N_44158);
nand U47147 (N_47147,N_44664,N_45296);
nor U47148 (N_47148,N_44202,N_45683);
or U47149 (N_47149,N_45815,N_45490);
xnor U47150 (N_47150,N_45171,N_44875);
nand U47151 (N_47151,N_44889,N_45407);
nand U47152 (N_47152,N_44458,N_44273);
xor U47153 (N_47153,N_44101,N_44378);
or U47154 (N_47154,N_45933,N_45305);
xor U47155 (N_47155,N_45694,N_44211);
xnor U47156 (N_47156,N_44155,N_44899);
nand U47157 (N_47157,N_45012,N_45908);
nand U47158 (N_47158,N_44216,N_45657);
nand U47159 (N_47159,N_45358,N_44057);
and U47160 (N_47160,N_44644,N_45399);
and U47161 (N_47161,N_44915,N_44963);
or U47162 (N_47162,N_44208,N_44928);
xnor U47163 (N_47163,N_44645,N_45785);
xor U47164 (N_47164,N_44893,N_44776);
nand U47165 (N_47165,N_45649,N_45122);
or U47166 (N_47166,N_45973,N_44958);
and U47167 (N_47167,N_44154,N_45794);
nor U47168 (N_47168,N_45257,N_45968);
nor U47169 (N_47169,N_44115,N_45505);
nor U47170 (N_47170,N_44506,N_44009);
or U47171 (N_47171,N_45667,N_44413);
nor U47172 (N_47172,N_44890,N_44199);
nand U47173 (N_47173,N_45664,N_45001);
nand U47174 (N_47174,N_45131,N_44832);
and U47175 (N_47175,N_45385,N_44582);
nand U47176 (N_47176,N_45191,N_45814);
and U47177 (N_47177,N_45641,N_44348);
xor U47178 (N_47178,N_44113,N_44232);
and U47179 (N_47179,N_45671,N_45703);
and U47180 (N_47180,N_45012,N_45414);
and U47181 (N_47181,N_44269,N_44014);
or U47182 (N_47182,N_45021,N_45982);
and U47183 (N_47183,N_45797,N_44831);
and U47184 (N_47184,N_45092,N_44009);
and U47185 (N_47185,N_44812,N_44564);
and U47186 (N_47186,N_44874,N_45782);
xor U47187 (N_47187,N_45128,N_45582);
or U47188 (N_47188,N_45297,N_45703);
and U47189 (N_47189,N_45717,N_45996);
and U47190 (N_47190,N_44841,N_44311);
xor U47191 (N_47191,N_45962,N_45448);
and U47192 (N_47192,N_44565,N_45954);
or U47193 (N_47193,N_45080,N_44333);
and U47194 (N_47194,N_44691,N_45898);
xnor U47195 (N_47195,N_45809,N_45585);
nand U47196 (N_47196,N_44648,N_45721);
or U47197 (N_47197,N_45058,N_44023);
nor U47198 (N_47198,N_45154,N_45434);
nand U47199 (N_47199,N_44963,N_44601);
xnor U47200 (N_47200,N_45613,N_44074);
xor U47201 (N_47201,N_44917,N_45652);
and U47202 (N_47202,N_45368,N_45700);
xnor U47203 (N_47203,N_45421,N_45506);
and U47204 (N_47204,N_45129,N_44345);
and U47205 (N_47205,N_45576,N_44093);
nand U47206 (N_47206,N_45818,N_44396);
xor U47207 (N_47207,N_45429,N_44963);
and U47208 (N_47208,N_45262,N_44553);
nand U47209 (N_47209,N_45650,N_45480);
and U47210 (N_47210,N_45747,N_45514);
or U47211 (N_47211,N_45316,N_44671);
and U47212 (N_47212,N_44596,N_44004);
nor U47213 (N_47213,N_45597,N_45804);
or U47214 (N_47214,N_44334,N_45085);
xor U47215 (N_47215,N_44270,N_44908);
or U47216 (N_47216,N_44959,N_44113);
and U47217 (N_47217,N_45581,N_45915);
xnor U47218 (N_47218,N_45948,N_44475);
and U47219 (N_47219,N_45481,N_44557);
or U47220 (N_47220,N_45887,N_44844);
or U47221 (N_47221,N_45259,N_44240);
and U47222 (N_47222,N_45705,N_45163);
nor U47223 (N_47223,N_44060,N_44614);
nand U47224 (N_47224,N_45728,N_44565);
nor U47225 (N_47225,N_44919,N_44542);
nor U47226 (N_47226,N_44876,N_45043);
nand U47227 (N_47227,N_44788,N_44544);
nand U47228 (N_47228,N_45227,N_44716);
nand U47229 (N_47229,N_44606,N_44734);
nor U47230 (N_47230,N_45626,N_44791);
or U47231 (N_47231,N_44178,N_45633);
or U47232 (N_47232,N_45487,N_45978);
xnor U47233 (N_47233,N_45415,N_45186);
and U47234 (N_47234,N_44129,N_45780);
nand U47235 (N_47235,N_44499,N_44189);
nand U47236 (N_47236,N_44676,N_44337);
nand U47237 (N_47237,N_44819,N_45824);
or U47238 (N_47238,N_45309,N_45568);
nand U47239 (N_47239,N_44801,N_45064);
nor U47240 (N_47240,N_44406,N_44834);
and U47241 (N_47241,N_44970,N_45955);
xor U47242 (N_47242,N_45406,N_45261);
xnor U47243 (N_47243,N_44925,N_44871);
nor U47244 (N_47244,N_45720,N_45583);
xor U47245 (N_47245,N_45326,N_44398);
and U47246 (N_47246,N_45660,N_45143);
and U47247 (N_47247,N_45850,N_44328);
or U47248 (N_47248,N_45813,N_45845);
xnor U47249 (N_47249,N_44788,N_45812);
nand U47250 (N_47250,N_45663,N_44356);
or U47251 (N_47251,N_45486,N_44222);
nor U47252 (N_47252,N_45422,N_45359);
nand U47253 (N_47253,N_45464,N_44250);
nor U47254 (N_47254,N_44030,N_45661);
and U47255 (N_47255,N_44647,N_45134);
nand U47256 (N_47256,N_45086,N_44436);
xnor U47257 (N_47257,N_45835,N_44985);
xor U47258 (N_47258,N_44248,N_44471);
or U47259 (N_47259,N_45653,N_45683);
nand U47260 (N_47260,N_45626,N_45105);
or U47261 (N_47261,N_45746,N_45908);
and U47262 (N_47262,N_45268,N_44336);
or U47263 (N_47263,N_44545,N_45844);
and U47264 (N_47264,N_44977,N_44073);
or U47265 (N_47265,N_44628,N_45472);
xor U47266 (N_47266,N_44666,N_45211);
xor U47267 (N_47267,N_44174,N_44671);
nand U47268 (N_47268,N_45254,N_45735);
nor U47269 (N_47269,N_45984,N_44608);
nand U47270 (N_47270,N_45694,N_45512);
nand U47271 (N_47271,N_44177,N_44973);
and U47272 (N_47272,N_45805,N_45225);
and U47273 (N_47273,N_44933,N_45890);
nand U47274 (N_47274,N_45767,N_44520);
nor U47275 (N_47275,N_44060,N_44648);
nor U47276 (N_47276,N_45833,N_44487);
nand U47277 (N_47277,N_44203,N_45195);
xnor U47278 (N_47278,N_44406,N_44269);
nand U47279 (N_47279,N_45291,N_45521);
and U47280 (N_47280,N_44191,N_45827);
or U47281 (N_47281,N_45845,N_45396);
nor U47282 (N_47282,N_44296,N_45501);
nand U47283 (N_47283,N_45823,N_45990);
or U47284 (N_47284,N_44886,N_44226);
nor U47285 (N_47285,N_45514,N_44909);
or U47286 (N_47286,N_45144,N_45045);
nor U47287 (N_47287,N_45077,N_44550);
nor U47288 (N_47288,N_44090,N_45165);
xor U47289 (N_47289,N_44878,N_45085);
or U47290 (N_47290,N_45633,N_44675);
nand U47291 (N_47291,N_44813,N_44722);
or U47292 (N_47292,N_44842,N_45484);
nor U47293 (N_47293,N_45318,N_44515);
nand U47294 (N_47294,N_45598,N_45683);
or U47295 (N_47295,N_44670,N_44263);
nor U47296 (N_47296,N_44046,N_45344);
and U47297 (N_47297,N_45825,N_44273);
nor U47298 (N_47298,N_44550,N_44980);
nand U47299 (N_47299,N_44397,N_44072);
or U47300 (N_47300,N_45773,N_45384);
nand U47301 (N_47301,N_44134,N_44683);
xor U47302 (N_47302,N_45743,N_44146);
xnor U47303 (N_47303,N_44149,N_44959);
nand U47304 (N_47304,N_44948,N_44060);
nor U47305 (N_47305,N_45672,N_45911);
or U47306 (N_47306,N_44297,N_44838);
xnor U47307 (N_47307,N_44668,N_45433);
nand U47308 (N_47308,N_45831,N_44358);
and U47309 (N_47309,N_44887,N_44555);
or U47310 (N_47310,N_44910,N_45154);
nor U47311 (N_47311,N_45029,N_44164);
nor U47312 (N_47312,N_44268,N_45107);
and U47313 (N_47313,N_44219,N_45462);
and U47314 (N_47314,N_45011,N_44685);
nor U47315 (N_47315,N_45645,N_45820);
nor U47316 (N_47316,N_45239,N_44586);
or U47317 (N_47317,N_44537,N_45242);
nor U47318 (N_47318,N_45813,N_45581);
xnor U47319 (N_47319,N_45675,N_44143);
nand U47320 (N_47320,N_45755,N_44451);
nand U47321 (N_47321,N_45716,N_44109);
nor U47322 (N_47322,N_44064,N_44746);
nor U47323 (N_47323,N_45248,N_44659);
or U47324 (N_47324,N_44840,N_44360);
or U47325 (N_47325,N_44163,N_45128);
nor U47326 (N_47326,N_45149,N_45671);
and U47327 (N_47327,N_44305,N_44100);
nor U47328 (N_47328,N_44395,N_45055);
and U47329 (N_47329,N_44376,N_45421);
or U47330 (N_47330,N_45448,N_44099);
and U47331 (N_47331,N_45153,N_44235);
or U47332 (N_47332,N_45906,N_44976);
xnor U47333 (N_47333,N_45223,N_44994);
or U47334 (N_47334,N_45058,N_44218);
and U47335 (N_47335,N_45323,N_44744);
xor U47336 (N_47336,N_45359,N_44325);
nor U47337 (N_47337,N_44448,N_44282);
xor U47338 (N_47338,N_45500,N_44011);
or U47339 (N_47339,N_44762,N_44011);
nor U47340 (N_47340,N_45282,N_44694);
or U47341 (N_47341,N_44622,N_45557);
or U47342 (N_47342,N_44483,N_44248);
nand U47343 (N_47343,N_45553,N_45627);
or U47344 (N_47344,N_45084,N_45216);
or U47345 (N_47345,N_45262,N_44239);
nand U47346 (N_47346,N_45195,N_44779);
or U47347 (N_47347,N_44924,N_44075);
nand U47348 (N_47348,N_44344,N_44853);
and U47349 (N_47349,N_44591,N_44331);
nor U47350 (N_47350,N_44515,N_44797);
nand U47351 (N_47351,N_45177,N_45233);
or U47352 (N_47352,N_44733,N_45179);
and U47353 (N_47353,N_44147,N_45674);
and U47354 (N_47354,N_44548,N_44870);
nor U47355 (N_47355,N_45700,N_44717);
nand U47356 (N_47356,N_44678,N_44365);
nand U47357 (N_47357,N_45954,N_45527);
xnor U47358 (N_47358,N_45858,N_45398);
nand U47359 (N_47359,N_45284,N_44303);
xor U47360 (N_47360,N_44999,N_44793);
and U47361 (N_47361,N_45615,N_45255);
nor U47362 (N_47362,N_44010,N_44707);
nor U47363 (N_47363,N_44644,N_44896);
nand U47364 (N_47364,N_44455,N_44028);
nand U47365 (N_47365,N_45550,N_45378);
nand U47366 (N_47366,N_45746,N_44371);
and U47367 (N_47367,N_44806,N_45179);
nand U47368 (N_47368,N_44575,N_45987);
or U47369 (N_47369,N_44989,N_44373);
xor U47370 (N_47370,N_45812,N_44389);
xor U47371 (N_47371,N_44211,N_45759);
nor U47372 (N_47372,N_45893,N_45247);
or U47373 (N_47373,N_44608,N_45775);
nand U47374 (N_47374,N_45567,N_45165);
nor U47375 (N_47375,N_44388,N_45997);
xnor U47376 (N_47376,N_44871,N_45419);
nand U47377 (N_47377,N_45252,N_45561);
or U47378 (N_47378,N_44479,N_44334);
and U47379 (N_47379,N_44727,N_44341);
xnor U47380 (N_47380,N_44108,N_45511);
or U47381 (N_47381,N_44276,N_45047);
xnor U47382 (N_47382,N_44981,N_44498);
and U47383 (N_47383,N_44417,N_45992);
and U47384 (N_47384,N_44931,N_45761);
xnor U47385 (N_47385,N_44623,N_44063);
nand U47386 (N_47386,N_44516,N_45312);
or U47387 (N_47387,N_44554,N_45497);
and U47388 (N_47388,N_45198,N_44428);
nor U47389 (N_47389,N_44065,N_45410);
xor U47390 (N_47390,N_44177,N_45064);
xnor U47391 (N_47391,N_44859,N_45427);
nor U47392 (N_47392,N_44206,N_44036);
xor U47393 (N_47393,N_44869,N_45888);
nand U47394 (N_47394,N_44922,N_44491);
or U47395 (N_47395,N_45259,N_45084);
or U47396 (N_47396,N_45978,N_44245);
or U47397 (N_47397,N_45421,N_45848);
nor U47398 (N_47398,N_44801,N_44837);
xor U47399 (N_47399,N_45029,N_45059);
or U47400 (N_47400,N_45972,N_44599);
nor U47401 (N_47401,N_44268,N_44578);
nor U47402 (N_47402,N_44125,N_45853);
nor U47403 (N_47403,N_44381,N_44315);
nor U47404 (N_47404,N_44062,N_44316);
or U47405 (N_47405,N_45220,N_44506);
xnor U47406 (N_47406,N_45697,N_45652);
and U47407 (N_47407,N_44661,N_45770);
or U47408 (N_47408,N_44154,N_44877);
and U47409 (N_47409,N_45516,N_45939);
nor U47410 (N_47410,N_45785,N_44225);
and U47411 (N_47411,N_45109,N_45265);
or U47412 (N_47412,N_44193,N_44781);
nor U47413 (N_47413,N_44136,N_44924);
and U47414 (N_47414,N_45738,N_45876);
or U47415 (N_47415,N_44454,N_45336);
and U47416 (N_47416,N_45856,N_44290);
nand U47417 (N_47417,N_44390,N_44042);
nand U47418 (N_47418,N_45300,N_44849);
nand U47419 (N_47419,N_44765,N_45819);
nor U47420 (N_47420,N_45380,N_45493);
and U47421 (N_47421,N_45722,N_44249);
nor U47422 (N_47422,N_45689,N_45700);
nand U47423 (N_47423,N_45252,N_44555);
nand U47424 (N_47424,N_45806,N_45362);
xnor U47425 (N_47425,N_44232,N_45296);
nand U47426 (N_47426,N_45088,N_45249);
xnor U47427 (N_47427,N_45662,N_44083);
nor U47428 (N_47428,N_45212,N_45059);
and U47429 (N_47429,N_45394,N_44563);
xnor U47430 (N_47430,N_45096,N_45643);
and U47431 (N_47431,N_44376,N_44725);
nor U47432 (N_47432,N_44447,N_45567);
and U47433 (N_47433,N_45723,N_44786);
or U47434 (N_47434,N_45352,N_45560);
xnor U47435 (N_47435,N_45329,N_44006);
xor U47436 (N_47436,N_44510,N_44078);
xnor U47437 (N_47437,N_44896,N_44714);
xor U47438 (N_47438,N_45060,N_45499);
and U47439 (N_47439,N_44953,N_44386);
nand U47440 (N_47440,N_45520,N_45329);
nand U47441 (N_47441,N_44527,N_44565);
xnor U47442 (N_47442,N_44322,N_44055);
nor U47443 (N_47443,N_44837,N_44503);
xor U47444 (N_47444,N_44854,N_45955);
nand U47445 (N_47445,N_45406,N_44308);
or U47446 (N_47446,N_45808,N_45299);
or U47447 (N_47447,N_45872,N_45469);
xnor U47448 (N_47448,N_44951,N_45350);
nor U47449 (N_47449,N_44757,N_44546);
nand U47450 (N_47450,N_44269,N_45795);
and U47451 (N_47451,N_44700,N_44825);
nor U47452 (N_47452,N_45176,N_44769);
xor U47453 (N_47453,N_44401,N_45936);
or U47454 (N_47454,N_45874,N_45076);
and U47455 (N_47455,N_44919,N_44932);
xnor U47456 (N_47456,N_44229,N_45698);
nand U47457 (N_47457,N_45413,N_44829);
nor U47458 (N_47458,N_45051,N_44920);
nand U47459 (N_47459,N_45104,N_44845);
or U47460 (N_47460,N_45045,N_45219);
nand U47461 (N_47461,N_44534,N_44053);
xnor U47462 (N_47462,N_45230,N_44691);
nor U47463 (N_47463,N_44632,N_44284);
and U47464 (N_47464,N_44705,N_45579);
or U47465 (N_47465,N_44032,N_44061);
and U47466 (N_47466,N_44326,N_45056);
or U47467 (N_47467,N_45525,N_45203);
nor U47468 (N_47468,N_45515,N_45798);
or U47469 (N_47469,N_45019,N_45225);
or U47470 (N_47470,N_45003,N_44146);
xor U47471 (N_47471,N_45825,N_45570);
and U47472 (N_47472,N_45860,N_45845);
and U47473 (N_47473,N_44043,N_44545);
and U47474 (N_47474,N_44905,N_44131);
and U47475 (N_47475,N_44894,N_45657);
nand U47476 (N_47476,N_45347,N_45973);
nand U47477 (N_47477,N_45441,N_45036);
and U47478 (N_47478,N_44429,N_45409);
xor U47479 (N_47479,N_45577,N_45077);
or U47480 (N_47480,N_45290,N_44629);
xnor U47481 (N_47481,N_45652,N_44595);
nor U47482 (N_47482,N_44821,N_45754);
nor U47483 (N_47483,N_44327,N_45223);
and U47484 (N_47484,N_45464,N_45891);
and U47485 (N_47485,N_44572,N_44853);
or U47486 (N_47486,N_44193,N_44676);
nor U47487 (N_47487,N_45400,N_45306);
and U47488 (N_47488,N_45816,N_45497);
nor U47489 (N_47489,N_44874,N_44087);
or U47490 (N_47490,N_45347,N_44780);
nand U47491 (N_47491,N_45082,N_45509);
or U47492 (N_47492,N_44550,N_44336);
or U47493 (N_47493,N_45884,N_44932);
nand U47494 (N_47494,N_45326,N_45724);
and U47495 (N_47495,N_44432,N_44358);
and U47496 (N_47496,N_45780,N_45564);
xnor U47497 (N_47497,N_45605,N_44517);
nor U47498 (N_47498,N_45643,N_45037);
and U47499 (N_47499,N_44765,N_44633);
and U47500 (N_47500,N_45653,N_45687);
nand U47501 (N_47501,N_44837,N_45946);
xnor U47502 (N_47502,N_44122,N_45335);
nand U47503 (N_47503,N_45329,N_45855);
xor U47504 (N_47504,N_44295,N_44933);
nand U47505 (N_47505,N_45310,N_44490);
nand U47506 (N_47506,N_44042,N_45090);
and U47507 (N_47507,N_44875,N_44445);
nand U47508 (N_47508,N_45660,N_44283);
or U47509 (N_47509,N_44882,N_45759);
nor U47510 (N_47510,N_45636,N_44435);
or U47511 (N_47511,N_44365,N_44107);
or U47512 (N_47512,N_44427,N_44780);
and U47513 (N_47513,N_44608,N_45439);
or U47514 (N_47514,N_45633,N_45152);
and U47515 (N_47515,N_44278,N_45925);
or U47516 (N_47516,N_45997,N_44497);
nand U47517 (N_47517,N_45329,N_45653);
nor U47518 (N_47518,N_44521,N_45103);
xor U47519 (N_47519,N_45444,N_45096);
nand U47520 (N_47520,N_45730,N_45612);
and U47521 (N_47521,N_45545,N_45632);
nand U47522 (N_47522,N_45132,N_45610);
nand U47523 (N_47523,N_45481,N_44711);
nor U47524 (N_47524,N_44760,N_45021);
nand U47525 (N_47525,N_44354,N_44777);
or U47526 (N_47526,N_45107,N_44614);
nand U47527 (N_47527,N_45364,N_45183);
and U47528 (N_47528,N_44525,N_44007);
nor U47529 (N_47529,N_44044,N_45532);
nor U47530 (N_47530,N_45161,N_45167);
or U47531 (N_47531,N_45432,N_44722);
xor U47532 (N_47532,N_45708,N_44447);
xnor U47533 (N_47533,N_45573,N_44584);
nor U47534 (N_47534,N_45919,N_44060);
and U47535 (N_47535,N_45968,N_45090);
nor U47536 (N_47536,N_44331,N_44490);
and U47537 (N_47537,N_44262,N_44143);
nand U47538 (N_47538,N_44964,N_45891);
or U47539 (N_47539,N_44717,N_44229);
nand U47540 (N_47540,N_44052,N_44349);
or U47541 (N_47541,N_44309,N_44708);
nor U47542 (N_47542,N_44591,N_44145);
nor U47543 (N_47543,N_44749,N_45591);
or U47544 (N_47544,N_45813,N_44844);
nor U47545 (N_47545,N_45716,N_45125);
or U47546 (N_47546,N_44822,N_45812);
nor U47547 (N_47547,N_44454,N_45518);
nor U47548 (N_47548,N_44839,N_45999);
and U47549 (N_47549,N_45933,N_44153);
nand U47550 (N_47550,N_45176,N_45089);
and U47551 (N_47551,N_44607,N_45502);
or U47552 (N_47552,N_44250,N_44674);
nand U47553 (N_47553,N_44981,N_44302);
nand U47554 (N_47554,N_44100,N_45857);
xnor U47555 (N_47555,N_45571,N_45549);
xor U47556 (N_47556,N_44091,N_44271);
nand U47557 (N_47557,N_45992,N_44535);
nor U47558 (N_47558,N_45295,N_44207);
or U47559 (N_47559,N_44675,N_44657);
xor U47560 (N_47560,N_45473,N_45472);
or U47561 (N_47561,N_44254,N_45800);
nand U47562 (N_47562,N_45460,N_44984);
xor U47563 (N_47563,N_45741,N_44684);
and U47564 (N_47564,N_45816,N_44750);
nor U47565 (N_47565,N_44297,N_44093);
xor U47566 (N_47566,N_44046,N_44292);
nor U47567 (N_47567,N_44054,N_44436);
and U47568 (N_47568,N_44204,N_44366);
or U47569 (N_47569,N_44871,N_45027);
xor U47570 (N_47570,N_44711,N_45618);
or U47571 (N_47571,N_45478,N_44654);
nand U47572 (N_47572,N_44368,N_45303);
or U47573 (N_47573,N_44748,N_44661);
and U47574 (N_47574,N_44380,N_45962);
nand U47575 (N_47575,N_44415,N_45856);
or U47576 (N_47576,N_44081,N_45520);
nor U47577 (N_47577,N_44420,N_44750);
nand U47578 (N_47578,N_45923,N_44737);
or U47579 (N_47579,N_44565,N_45305);
nand U47580 (N_47580,N_44274,N_45225);
and U47581 (N_47581,N_45982,N_45954);
or U47582 (N_47582,N_44858,N_45266);
xnor U47583 (N_47583,N_44019,N_44696);
nand U47584 (N_47584,N_45262,N_45163);
and U47585 (N_47585,N_44252,N_45400);
nor U47586 (N_47586,N_44851,N_44122);
xor U47587 (N_47587,N_45645,N_45457);
nand U47588 (N_47588,N_44978,N_45411);
nand U47589 (N_47589,N_44128,N_45481);
nor U47590 (N_47590,N_44241,N_45175);
nor U47591 (N_47591,N_45647,N_44513);
nor U47592 (N_47592,N_45901,N_44290);
nor U47593 (N_47593,N_44698,N_44566);
and U47594 (N_47594,N_45819,N_45945);
or U47595 (N_47595,N_44322,N_44068);
xnor U47596 (N_47596,N_44170,N_44855);
nand U47597 (N_47597,N_44556,N_45974);
or U47598 (N_47598,N_44726,N_45748);
nand U47599 (N_47599,N_44084,N_45700);
and U47600 (N_47600,N_44844,N_45476);
and U47601 (N_47601,N_45618,N_45353);
nand U47602 (N_47602,N_44314,N_45356);
nor U47603 (N_47603,N_44664,N_44785);
or U47604 (N_47604,N_45957,N_45045);
and U47605 (N_47605,N_44223,N_44682);
or U47606 (N_47606,N_44021,N_45610);
nand U47607 (N_47607,N_44753,N_44167);
nand U47608 (N_47608,N_44798,N_45120);
and U47609 (N_47609,N_44418,N_45627);
nand U47610 (N_47610,N_45313,N_44776);
or U47611 (N_47611,N_45326,N_45270);
nor U47612 (N_47612,N_45344,N_45986);
xnor U47613 (N_47613,N_44431,N_44505);
nand U47614 (N_47614,N_44555,N_45999);
or U47615 (N_47615,N_44145,N_45005);
xor U47616 (N_47616,N_44543,N_44145);
xnor U47617 (N_47617,N_45886,N_45249);
nor U47618 (N_47618,N_45267,N_44818);
or U47619 (N_47619,N_45979,N_45620);
nand U47620 (N_47620,N_45260,N_44677);
and U47621 (N_47621,N_44970,N_45512);
nor U47622 (N_47622,N_45041,N_45778);
or U47623 (N_47623,N_44715,N_45428);
xor U47624 (N_47624,N_44187,N_44278);
xnor U47625 (N_47625,N_44549,N_45285);
nand U47626 (N_47626,N_44244,N_44169);
nand U47627 (N_47627,N_44465,N_45618);
or U47628 (N_47628,N_44022,N_45942);
and U47629 (N_47629,N_45171,N_45952);
or U47630 (N_47630,N_44755,N_45903);
or U47631 (N_47631,N_45123,N_44523);
and U47632 (N_47632,N_45838,N_45085);
xor U47633 (N_47633,N_45170,N_44000);
nor U47634 (N_47634,N_45430,N_44520);
and U47635 (N_47635,N_45694,N_44940);
and U47636 (N_47636,N_45247,N_44413);
nor U47637 (N_47637,N_45462,N_44337);
nor U47638 (N_47638,N_45088,N_45230);
or U47639 (N_47639,N_45411,N_45711);
xor U47640 (N_47640,N_45637,N_45262);
and U47641 (N_47641,N_45488,N_45567);
and U47642 (N_47642,N_45577,N_45562);
and U47643 (N_47643,N_44401,N_44395);
xnor U47644 (N_47644,N_45667,N_45048);
nand U47645 (N_47645,N_45162,N_45154);
and U47646 (N_47646,N_45295,N_45967);
or U47647 (N_47647,N_45895,N_45029);
nor U47648 (N_47648,N_45301,N_44324);
xor U47649 (N_47649,N_44940,N_44942);
nor U47650 (N_47650,N_45916,N_44619);
or U47651 (N_47651,N_44842,N_44477);
nand U47652 (N_47652,N_44641,N_44732);
and U47653 (N_47653,N_45792,N_45196);
xnor U47654 (N_47654,N_45477,N_44696);
and U47655 (N_47655,N_44030,N_45349);
and U47656 (N_47656,N_44974,N_45388);
nor U47657 (N_47657,N_44231,N_44253);
or U47658 (N_47658,N_45701,N_45616);
or U47659 (N_47659,N_44603,N_44364);
and U47660 (N_47660,N_44369,N_44457);
nor U47661 (N_47661,N_44223,N_45618);
and U47662 (N_47662,N_45592,N_44888);
and U47663 (N_47663,N_45742,N_45867);
nand U47664 (N_47664,N_45039,N_44102);
xor U47665 (N_47665,N_44583,N_44065);
xnor U47666 (N_47666,N_44854,N_45504);
nand U47667 (N_47667,N_44381,N_44961);
xor U47668 (N_47668,N_44947,N_44362);
and U47669 (N_47669,N_45040,N_45363);
nor U47670 (N_47670,N_44375,N_45657);
nand U47671 (N_47671,N_45828,N_44526);
or U47672 (N_47672,N_45901,N_45923);
or U47673 (N_47673,N_45958,N_45855);
and U47674 (N_47674,N_44926,N_44849);
xnor U47675 (N_47675,N_45833,N_44122);
xnor U47676 (N_47676,N_44317,N_45291);
and U47677 (N_47677,N_45031,N_44234);
nand U47678 (N_47678,N_44340,N_45660);
and U47679 (N_47679,N_45359,N_45313);
nand U47680 (N_47680,N_45280,N_45762);
nand U47681 (N_47681,N_44780,N_45932);
xnor U47682 (N_47682,N_44854,N_45651);
or U47683 (N_47683,N_44470,N_45223);
nor U47684 (N_47684,N_45330,N_45576);
nand U47685 (N_47685,N_44363,N_44901);
or U47686 (N_47686,N_45163,N_45582);
nand U47687 (N_47687,N_44021,N_44036);
or U47688 (N_47688,N_45207,N_44139);
and U47689 (N_47689,N_44458,N_44263);
nand U47690 (N_47690,N_44352,N_44251);
xor U47691 (N_47691,N_45208,N_44576);
xnor U47692 (N_47692,N_44718,N_45813);
xor U47693 (N_47693,N_45940,N_45480);
nand U47694 (N_47694,N_44537,N_44812);
nand U47695 (N_47695,N_44238,N_44013);
or U47696 (N_47696,N_44479,N_44102);
and U47697 (N_47697,N_44193,N_44568);
nor U47698 (N_47698,N_44367,N_45399);
and U47699 (N_47699,N_45889,N_45435);
xnor U47700 (N_47700,N_44812,N_44999);
nand U47701 (N_47701,N_44042,N_44037);
xor U47702 (N_47702,N_45881,N_44661);
nand U47703 (N_47703,N_44591,N_44311);
nor U47704 (N_47704,N_45980,N_45908);
and U47705 (N_47705,N_44962,N_44538);
or U47706 (N_47706,N_45983,N_44161);
xor U47707 (N_47707,N_45238,N_44598);
nand U47708 (N_47708,N_45307,N_45293);
or U47709 (N_47709,N_44806,N_44539);
or U47710 (N_47710,N_44527,N_45254);
nor U47711 (N_47711,N_45781,N_45589);
and U47712 (N_47712,N_44956,N_44108);
nand U47713 (N_47713,N_44746,N_45042);
or U47714 (N_47714,N_45669,N_45886);
and U47715 (N_47715,N_45077,N_44620);
and U47716 (N_47716,N_44597,N_45088);
and U47717 (N_47717,N_45287,N_44827);
or U47718 (N_47718,N_44814,N_44084);
nand U47719 (N_47719,N_45967,N_45869);
nand U47720 (N_47720,N_45811,N_44316);
nor U47721 (N_47721,N_44804,N_44531);
xnor U47722 (N_47722,N_44286,N_44629);
nand U47723 (N_47723,N_45897,N_45193);
or U47724 (N_47724,N_44691,N_44639);
xor U47725 (N_47725,N_45778,N_44908);
nand U47726 (N_47726,N_45685,N_45723);
nand U47727 (N_47727,N_44339,N_45632);
nand U47728 (N_47728,N_44879,N_45057);
nand U47729 (N_47729,N_44419,N_44583);
nor U47730 (N_47730,N_45301,N_44774);
and U47731 (N_47731,N_45864,N_44218);
xnor U47732 (N_47732,N_44295,N_44007);
xnor U47733 (N_47733,N_45135,N_44588);
xor U47734 (N_47734,N_45351,N_44117);
xor U47735 (N_47735,N_45539,N_45992);
nor U47736 (N_47736,N_45602,N_45589);
nor U47737 (N_47737,N_45083,N_44274);
and U47738 (N_47738,N_44736,N_45333);
nand U47739 (N_47739,N_44795,N_44854);
xnor U47740 (N_47740,N_44365,N_45036);
xnor U47741 (N_47741,N_44093,N_45535);
and U47742 (N_47742,N_45216,N_44755);
xor U47743 (N_47743,N_44034,N_44448);
or U47744 (N_47744,N_44244,N_44862);
and U47745 (N_47745,N_44787,N_44092);
or U47746 (N_47746,N_45520,N_44748);
nand U47747 (N_47747,N_45394,N_45354);
nand U47748 (N_47748,N_44667,N_44954);
nor U47749 (N_47749,N_45301,N_44781);
nor U47750 (N_47750,N_45844,N_45567);
nor U47751 (N_47751,N_45404,N_44845);
nand U47752 (N_47752,N_45553,N_44455);
and U47753 (N_47753,N_44603,N_44102);
or U47754 (N_47754,N_44537,N_45542);
nor U47755 (N_47755,N_45658,N_45119);
nor U47756 (N_47756,N_44273,N_44386);
xnor U47757 (N_47757,N_44754,N_45552);
and U47758 (N_47758,N_45547,N_44224);
and U47759 (N_47759,N_44067,N_44668);
and U47760 (N_47760,N_44059,N_45760);
and U47761 (N_47761,N_45746,N_45837);
and U47762 (N_47762,N_45331,N_44294);
and U47763 (N_47763,N_45305,N_45961);
xor U47764 (N_47764,N_44527,N_45379);
and U47765 (N_47765,N_45612,N_45903);
nand U47766 (N_47766,N_44411,N_44699);
nor U47767 (N_47767,N_45734,N_44437);
and U47768 (N_47768,N_45179,N_45690);
and U47769 (N_47769,N_44355,N_45284);
and U47770 (N_47770,N_44233,N_44677);
and U47771 (N_47771,N_45900,N_45165);
or U47772 (N_47772,N_45733,N_45028);
nor U47773 (N_47773,N_45762,N_45348);
and U47774 (N_47774,N_44651,N_44045);
nand U47775 (N_47775,N_45588,N_44356);
nor U47776 (N_47776,N_45330,N_44003);
nand U47777 (N_47777,N_44650,N_44647);
and U47778 (N_47778,N_44736,N_44903);
xor U47779 (N_47779,N_44679,N_44534);
nor U47780 (N_47780,N_45126,N_45380);
and U47781 (N_47781,N_44310,N_45113);
xnor U47782 (N_47782,N_45037,N_45940);
and U47783 (N_47783,N_45326,N_44557);
xnor U47784 (N_47784,N_45018,N_44738);
and U47785 (N_47785,N_44339,N_44480);
nand U47786 (N_47786,N_44747,N_44472);
and U47787 (N_47787,N_45209,N_44346);
nor U47788 (N_47788,N_45100,N_45667);
xor U47789 (N_47789,N_44433,N_45566);
xnor U47790 (N_47790,N_45607,N_45218);
nand U47791 (N_47791,N_45111,N_45278);
nand U47792 (N_47792,N_45923,N_44066);
xor U47793 (N_47793,N_45083,N_45231);
or U47794 (N_47794,N_45827,N_44494);
or U47795 (N_47795,N_44721,N_44149);
nand U47796 (N_47796,N_44635,N_45428);
nand U47797 (N_47797,N_44495,N_44503);
nand U47798 (N_47798,N_45319,N_44321);
or U47799 (N_47799,N_44505,N_44589);
xnor U47800 (N_47800,N_44498,N_45473);
or U47801 (N_47801,N_44941,N_45705);
or U47802 (N_47802,N_45437,N_44325);
or U47803 (N_47803,N_45481,N_44352);
nand U47804 (N_47804,N_44347,N_45701);
nor U47805 (N_47805,N_45791,N_44682);
and U47806 (N_47806,N_44804,N_44159);
nor U47807 (N_47807,N_45698,N_45627);
xor U47808 (N_47808,N_45882,N_45261);
or U47809 (N_47809,N_44765,N_44886);
xnor U47810 (N_47810,N_45350,N_44213);
xor U47811 (N_47811,N_44702,N_45074);
or U47812 (N_47812,N_45034,N_45928);
or U47813 (N_47813,N_44433,N_44809);
nand U47814 (N_47814,N_45029,N_44517);
or U47815 (N_47815,N_45317,N_44236);
nor U47816 (N_47816,N_45265,N_44303);
and U47817 (N_47817,N_45175,N_44956);
nor U47818 (N_47818,N_44545,N_44571);
xnor U47819 (N_47819,N_44543,N_44481);
and U47820 (N_47820,N_44940,N_44116);
nand U47821 (N_47821,N_45154,N_45264);
and U47822 (N_47822,N_45424,N_45527);
or U47823 (N_47823,N_45560,N_45890);
and U47824 (N_47824,N_45626,N_44946);
nand U47825 (N_47825,N_45655,N_45873);
and U47826 (N_47826,N_45745,N_44978);
nor U47827 (N_47827,N_44836,N_44711);
and U47828 (N_47828,N_45897,N_45719);
nand U47829 (N_47829,N_45095,N_45447);
and U47830 (N_47830,N_45369,N_44748);
nor U47831 (N_47831,N_44653,N_45877);
or U47832 (N_47832,N_45649,N_44762);
or U47833 (N_47833,N_44852,N_45347);
nand U47834 (N_47834,N_45119,N_45349);
and U47835 (N_47835,N_44301,N_44807);
and U47836 (N_47836,N_45940,N_45123);
or U47837 (N_47837,N_44092,N_44922);
and U47838 (N_47838,N_45496,N_44391);
xor U47839 (N_47839,N_45966,N_44883);
or U47840 (N_47840,N_45938,N_44319);
nand U47841 (N_47841,N_44579,N_44323);
nand U47842 (N_47842,N_45858,N_45507);
nor U47843 (N_47843,N_45819,N_45859);
and U47844 (N_47844,N_44212,N_44956);
xnor U47845 (N_47845,N_45804,N_44830);
nor U47846 (N_47846,N_45715,N_45607);
nand U47847 (N_47847,N_45772,N_44240);
or U47848 (N_47848,N_45796,N_45173);
nor U47849 (N_47849,N_44588,N_45266);
or U47850 (N_47850,N_44437,N_44911);
or U47851 (N_47851,N_44855,N_45247);
and U47852 (N_47852,N_44659,N_44932);
nor U47853 (N_47853,N_44001,N_45120);
and U47854 (N_47854,N_45676,N_44148);
or U47855 (N_47855,N_44666,N_44032);
or U47856 (N_47856,N_45089,N_45988);
nor U47857 (N_47857,N_44101,N_44632);
or U47858 (N_47858,N_44366,N_44851);
nand U47859 (N_47859,N_44778,N_45841);
or U47860 (N_47860,N_45444,N_44965);
xnor U47861 (N_47861,N_44733,N_45881);
nor U47862 (N_47862,N_45258,N_45055);
or U47863 (N_47863,N_45036,N_44040);
or U47864 (N_47864,N_45471,N_44499);
nand U47865 (N_47865,N_45870,N_45152);
xor U47866 (N_47866,N_45239,N_45834);
and U47867 (N_47867,N_45522,N_45422);
nand U47868 (N_47868,N_45814,N_45118);
and U47869 (N_47869,N_45958,N_45026);
xnor U47870 (N_47870,N_45848,N_44715);
and U47871 (N_47871,N_44334,N_45346);
xor U47872 (N_47872,N_44688,N_45666);
or U47873 (N_47873,N_45291,N_45380);
or U47874 (N_47874,N_44862,N_45172);
or U47875 (N_47875,N_45357,N_45304);
xor U47876 (N_47876,N_45532,N_44450);
nand U47877 (N_47877,N_45391,N_45898);
nand U47878 (N_47878,N_44609,N_44517);
nor U47879 (N_47879,N_44939,N_44422);
or U47880 (N_47880,N_44785,N_44377);
nor U47881 (N_47881,N_44389,N_45032);
nand U47882 (N_47882,N_44256,N_45121);
nor U47883 (N_47883,N_44907,N_44396);
nor U47884 (N_47884,N_44477,N_44408);
nand U47885 (N_47885,N_44293,N_44308);
nor U47886 (N_47886,N_45945,N_45158);
and U47887 (N_47887,N_44788,N_45434);
and U47888 (N_47888,N_44243,N_44862);
nor U47889 (N_47889,N_45319,N_45709);
and U47890 (N_47890,N_45781,N_45070);
xnor U47891 (N_47891,N_44195,N_45103);
nor U47892 (N_47892,N_45702,N_44004);
nand U47893 (N_47893,N_45555,N_45006);
nand U47894 (N_47894,N_45581,N_44067);
or U47895 (N_47895,N_44033,N_45166);
nand U47896 (N_47896,N_44806,N_44255);
nand U47897 (N_47897,N_44291,N_44255);
and U47898 (N_47898,N_44967,N_45302);
or U47899 (N_47899,N_44897,N_45267);
or U47900 (N_47900,N_45487,N_44922);
nor U47901 (N_47901,N_44875,N_44507);
and U47902 (N_47902,N_44539,N_45080);
or U47903 (N_47903,N_44585,N_45593);
nor U47904 (N_47904,N_45064,N_45387);
and U47905 (N_47905,N_44328,N_45395);
nor U47906 (N_47906,N_45908,N_45949);
xor U47907 (N_47907,N_45848,N_45370);
xor U47908 (N_47908,N_44172,N_44268);
or U47909 (N_47909,N_44245,N_45914);
nor U47910 (N_47910,N_45997,N_44806);
xnor U47911 (N_47911,N_45724,N_45813);
nor U47912 (N_47912,N_45301,N_45006);
nor U47913 (N_47913,N_44614,N_45959);
nand U47914 (N_47914,N_45032,N_45902);
nor U47915 (N_47915,N_45226,N_45229);
and U47916 (N_47916,N_45093,N_44391);
nor U47917 (N_47917,N_45031,N_45184);
nand U47918 (N_47918,N_44843,N_44938);
and U47919 (N_47919,N_44621,N_44383);
nand U47920 (N_47920,N_45596,N_45968);
nor U47921 (N_47921,N_45648,N_45391);
xnor U47922 (N_47922,N_44875,N_45191);
xor U47923 (N_47923,N_45710,N_44948);
and U47924 (N_47924,N_45655,N_45804);
nand U47925 (N_47925,N_45779,N_45976);
nand U47926 (N_47926,N_44751,N_44769);
nor U47927 (N_47927,N_45159,N_45915);
nor U47928 (N_47928,N_45334,N_44711);
or U47929 (N_47929,N_44830,N_45807);
xor U47930 (N_47930,N_45197,N_45434);
nor U47931 (N_47931,N_44981,N_45733);
xor U47932 (N_47932,N_44545,N_45660);
or U47933 (N_47933,N_45764,N_44725);
nor U47934 (N_47934,N_45820,N_44972);
nor U47935 (N_47935,N_45112,N_44391);
nor U47936 (N_47936,N_44753,N_45013);
or U47937 (N_47937,N_45891,N_44088);
and U47938 (N_47938,N_44248,N_44060);
or U47939 (N_47939,N_44337,N_44855);
and U47940 (N_47940,N_44519,N_44064);
nor U47941 (N_47941,N_44696,N_45430);
and U47942 (N_47942,N_44707,N_45238);
nand U47943 (N_47943,N_45433,N_44549);
nor U47944 (N_47944,N_45787,N_45599);
xnor U47945 (N_47945,N_44390,N_45629);
nor U47946 (N_47946,N_44377,N_44547);
or U47947 (N_47947,N_45644,N_45428);
and U47948 (N_47948,N_45687,N_44268);
or U47949 (N_47949,N_44389,N_45853);
or U47950 (N_47950,N_45303,N_44917);
xnor U47951 (N_47951,N_44856,N_44236);
nor U47952 (N_47952,N_44415,N_44418);
or U47953 (N_47953,N_44322,N_45485);
or U47954 (N_47954,N_45864,N_45842);
or U47955 (N_47955,N_44574,N_45839);
xnor U47956 (N_47956,N_45445,N_45391);
nor U47957 (N_47957,N_44503,N_44827);
xor U47958 (N_47958,N_45081,N_45521);
and U47959 (N_47959,N_44862,N_44326);
or U47960 (N_47960,N_45881,N_44966);
or U47961 (N_47961,N_44377,N_45387);
nor U47962 (N_47962,N_44589,N_45708);
nand U47963 (N_47963,N_45287,N_45506);
nand U47964 (N_47964,N_45502,N_45932);
xnor U47965 (N_47965,N_45027,N_44478);
nand U47966 (N_47966,N_45161,N_44637);
or U47967 (N_47967,N_45376,N_44057);
or U47968 (N_47968,N_44554,N_45057);
nor U47969 (N_47969,N_44878,N_45540);
nand U47970 (N_47970,N_45123,N_45036);
and U47971 (N_47971,N_45528,N_44903);
or U47972 (N_47972,N_44033,N_44352);
nand U47973 (N_47973,N_44245,N_44663);
nor U47974 (N_47974,N_45376,N_45289);
and U47975 (N_47975,N_45341,N_44550);
or U47976 (N_47976,N_45215,N_45575);
nand U47977 (N_47977,N_44008,N_44808);
or U47978 (N_47978,N_44506,N_44223);
nor U47979 (N_47979,N_44730,N_45583);
and U47980 (N_47980,N_45490,N_45743);
nor U47981 (N_47981,N_44351,N_44828);
and U47982 (N_47982,N_44148,N_44482);
or U47983 (N_47983,N_45435,N_45966);
or U47984 (N_47984,N_45609,N_45603);
xor U47985 (N_47985,N_44554,N_45409);
nor U47986 (N_47986,N_44745,N_44889);
and U47987 (N_47987,N_44747,N_45285);
xnor U47988 (N_47988,N_44909,N_45705);
xor U47989 (N_47989,N_44765,N_45736);
nand U47990 (N_47990,N_44212,N_45072);
nand U47991 (N_47991,N_44407,N_45128);
or U47992 (N_47992,N_45428,N_44594);
nand U47993 (N_47993,N_45931,N_45888);
xor U47994 (N_47994,N_44619,N_45018);
nor U47995 (N_47995,N_45935,N_44015);
or U47996 (N_47996,N_44386,N_44427);
nor U47997 (N_47997,N_45822,N_44394);
nor U47998 (N_47998,N_44192,N_45696);
or U47999 (N_47999,N_45871,N_45198);
nor U48000 (N_48000,N_47263,N_47182);
and U48001 (N_48001,N_46578,N_47489);
xnor U48002 (N_48002,N_47121,N_46826);
and U48003 (N_48003,N_46842,N_46856);
nor U48004 (N_48004,N_46443,N_47696);
nand U48005 (N_48005,N_46113,N_47599);
and U48006 (N_48006,N_47430,N_46374);
nor U48007 (N_48007,N_47268,N_47473);
and U48008 (N_48008,N_46684,N_46034);
or U48009 (N_48009,N_46143,N_46698);
and U48010 (N_48010,N_46899,N_47362);
or U48011 (N_48011,N_46975,N_46091);
nor U48012 (N_48012,N_46241,N_47654);
and U48013 (N_48013,N_47206,N_47485);
nor U48014 (N_48014,N_46930,N_46406);
nand U48015 (N_48015,N_46226,N_47822);
xnor U48016 (N_48016,N_46741,N_47701);
nor U48017 (N_48017,N_47666,N_46738);
and U48018 (N_48018,N_46915,N_47639);
xnor U48019 (N_48019,N_46840,N_46779);
and U48020 (N_48020,N_47275,N_46123);
and U48021 (N_48021,N_47222,N_46740);
nor U48022 (N_48022,N_47703,N_47921);
and U48023 (N_48023,N_46327,N_46714);
or U48024 (N_48024,N_46665,N_46978);
nand U48025 (N_48025,N_47176,N_46792);
nand U48026 (N_48026,N_46903,N_47071);
nand U48027 (N_48027,N_47949,N_46994);
xnor U48028 (N_48028,N_46950,N_47594);
and U48029 (N_48029,N_47997,N_47324);
xor U48030 (N_48030,N_47629,N_46094);
nor U48031 (N_48031,N_47285,N_47885);
nor U48032 (N_48032,N_47080,N_47815);
xnor U48033 (N_48033,N_47099,N_47742);
and U48034 (N_48034,N_47695,N_47297);
nand U48035 (N_48035,N_47502,N_46653);
nor U48036 (N_48036,N_46633,N_46832);
and U48037 (N_48037,N_46439,N_47951);
xnor U48038 (N_48038,N_47211,N_47950);
nor U48039 (N_48039,N_47294,N_47939);
xor U48040 (N_48040,N_47414,N_46254);
or U48041 (N_48041,N_46795,N_47563);
and U48042 (N_48042,N_47482,N_47513);
nand U48043 (N_48043,N_47245,N_46908);
nand U48044 (N_48044,N_46289,N_46202);
and U48045 (N_48045,N_47784,N_47795);
and U48046 (N_48046,N_47323,N_47011);
and U48047 (N_48047,N_47169,N_46763);
nand U48048 (N_48048,N_47787,N_46682);
or U48049 (N_48049,N_47461,N_46024);
and U48050 (N_48050,N_46223,N_47445);
or U48051 (N_48051,N_47491,N_47857);
xnor U48052 (N_48052,N_46862,N_47259);
nand U48053 (N_48053,N_47922,N_47349);
or U48054 (N_48054,N_46555,N_46829);
xor U48055 (N_48055,N_47284,N_47722);
nor U48056 (N_48056,N_47436,N_47013);
nor U48057 (N_48057,N_46947,N_47768);
xor U48058 (N_48058,N_46340,N_46520);
nand U48059 (N_48059,N_46552,N_46025);
nand U48060 (N_48060,N_46110,N_47904);
or U48061 (N_48061,N_47447,N_46086);
and U48062 (N_48062,N_47283,N_46918);
and U48063 (N_48063,N_47823,N_46464);
xor U48064 (N_48064,N_46373,N_47129);
xnor U48065 (N_48065,N_46619,N_47780);
xnor U48066 (N_48066,N_46215,N_47651);
and U48067 (N_48067,N_46463,N_46438);
and U48068 (N_48068,N_47912,N_47088);
and U48069 (N_48069,N_47170,N_46356);
and U48070 (N_48070,N_46193,N_47338);
xor U48071 (N_48071,N_47495,N_47753);
nor U48072 (N_48072,N_46958,N_46434);
or U48073 (N_48073,N_46906,N_47261);
and U48074 (N_48074,N_46135,N_47029);
and U48075 (N_48075,N_47942,N_47303);
nor U48076 (N_48076,N_47581,N_46368);
xor U48077 (N_48077,N_46594,N_47905);
nor U48078 (N_48078,N_47592,N_47167);
nor U48079 (N_48079,N_46852,N_47070);
xnor U48080 (N_48080,N_47794,N_46380);
xor U48081 (N_48081,N_46557,N_46784);
or U48082 (N_48082,N_46338,N_47640);
or U48083 (N_48083,N_46636,N_47340);
nor U48084 (N_48084,N_47091,N_46657);
or U48085 (N_48085,N_47327,N_47838);
nor U48086 (N_48086,N_46080,N_46582);
nor U48087 (N_48087,N_47896,N_47769);
xor U48088 (N_48088,N_47273,N_47940);
and U48089 (N_48089,N_47007,N_46554);
nand U48090 (N_48090,N_46956,N_46854);
nand U48091 (N_48091,N_46722,N_46651);
and U48092 (N_48092,N_46914,N_47184);
nand U48093 (N_48093,N_46361,N_46175);
or U48094 (N_48094,N_47936,N_47434);
or U48095 (N_48095,N_46359,N_47636);
nor U48096 (N_48096,N_47322,N_46833);
or U48097 (N_48097,N_47484,N_47943);
and U48098 (N_48098,N_46635,N_47153);
xor U48099 (N_48099,N_47188,N_47891);
nand U48100 (N_48100,N_46627,N_46272);
xor U48101 (N_48101,N_47510,N_46560);
nand U48102 (N_48102,N_46339,N_46543);
nand U48103 (N_48103,N_47288,N_46263);
xor U48104 (N_48104,N_46284,N_47138);
xnor U48105 (N_48105,N_47757,N_47791);
xor U48106 (N_48106,N_47927,N_46590);
nor U48107 (N_48107,N_47572,N_47957);
and U48108 (N_48108,N_47019,N_46810);
or U48109 (N_48109,N_47603,N_46706);
nand U48110 (N_48110,N_47133,N_47418);
nor U48111 (N_48111,N_47549,N_46404);
and U48112 (N_48112,N_47577,N_47365);
nor U48113 (N_48113,N_47413,N_47098);
nor U48114 (N_48114,N_47953,N_47149);
or U48115 (N_48115,N_46728,N_47755);
nor U48116 (N_48116,N_47821,N_47317);
nor U48117 (N_48117,N_46746,N_47713);
and U48118 (N_48118,N_47635,N_47670);
xnor U48119 (N_48119,N_47583,N_47628);
nand U48120 (N_48120,N_46939,N_47358);
nand U48121 (N_48121,N_47910,N_46184);
xnor U48122 (N_48122,N_47306,N_46343);
xnor U48123 (N_48123,N_47472,N_46358);
xnor U48124 (N_48124,N_47218,N_46020);
or U48125 (N_48125,N_46791,N_47889);
or U48126 (N_48126,N_47551,N_46616);
and U48127 (N_48127,N_46973,N_46109);
and U48128 (N_48128,N_46448,N_46285);
xor U48129 (N_48129,N_46321,N_47415);
or U48130 (N_48130,N_46496,N_47134);
and U48131 (N_48131,N_46154,N_46008);
xor U48132 (N_48132,N_46498,N_47870);
and U48133 (N_48133,N_46513,N_47638);
or U48134 (N_48134,N_46152,N_47747);
xnor U48135 (N_48135,N_46893,N_47678);
xor U48136 (N_48136,N_46046,N_46063);
nand U48137 (N_48137,N_46479,N_46467);
xor U48138 (N_48138,N_47089,N_47475);
xnor U48139 (N_48139,N_46730,N_47320);
or U48140 (N_48140,N_47952,N_47156);
nor U48141 (N_48141,N_47751,N_47689);
nor U48142 (N_48142,N_46157,N_46902);
nor U48143 (N_48143,N_46737,N_46435);
xor U48144 (N_48144,N_46172,N_46645);
nand U48145 (N_48145,N_47215,N_46153);
nor U48146 (N_48146,N_46476,N_47216);
nor U48147 (N_48147,N_47189,N_47137);
nor U48148 (N_48148,N_46989,N_47202);
or U48149 (N_48149,N_47253,N_46235);
nor U48150 (N_48150,N_46119,N_46752);
xor U48151 (N_48151,N_46692,N_47114);
nand U48152 (N_48152,N_46650,N_47803);
and U48153 (N_48153,N_47490,N_47839);
nand U48154 (N_48154,N_47084,N_46132);
or U48155 (N_48155,N_47076,N_46971);
and U48156 (N_48156,N_47251,N_46170);
or U48157 (N_48157,N_46988,N_47861);
nor U48158 (N_48158,N_46394,N_47824);
nor U48159 (N_48159,N_46882,N_47964);
and U48160 (N_48160,N_46984,N_46534);
or U48161 (N_48161,N_47179,N_47056);
nor U48162 (N_48162,N_46079,N_47183);
and U48163 (N_48163,N_47799,N_46201);
xnor U48164 (N_48164,N_47668,N_46995);
nand U48165 (N_48165,N_47985,N_47622);
and U48166 (N_48166,N_46585,N_47582);
xor U48167 (N_48167,N_46142,N_46458);
nor U48168 (N_48168,N_46589,N_47033);
and U48169 (N_48169,N_46867,N_46245);
nand U48170 (N_48170,N_47903,N_46058);
and U48171 (N_48171,N_47597,N_46219);
nand U48172 (N_48172,N_46487,N_47224);
and U48173 (N_48173,N_46983,N_47657);
nor U48174 (N_48174,N_46656,N_47230);
xnor U48175 (N_48175,N_46937,N_47858);
nand U48176 (N_48176,N_47965,N_47348);
xnor U48177 (N_48177,N_46828,N_47381);
nor U48178 (N_48178,N_47496,N_46910);
nor U48179 (N_48179,N_47938,N_47819);
nand U48180 (N_48180,N_47527,N_46033);
xnor U48181 (N_48181,N_47544,N_47093);
nand U48182 (N_48182,N_46583,N_46528);
nor U48183 (N_48183,N_47069,N_46690);
nor U48184 (N_48184,N_47522,N_47337);
xor U48185 (N_48185,N_46881,N_46688);
or U48186 (N_48186,N_46878,N_46281);
xnor U48187 (N_48187,N_47743,N_47166);
or U48188 (N_48188,N_46278,N_47034);
and U48189 (N_48189,N_46040,N_47372);
nand U48190 (N_48190,N_47781,N_47983);
xnor U48191 (N_48191,N_47924,N_46287);
or U48192 (N_48192,N_47431,N_46609);
or U48193 (N_48193,N_47669,N_46725);
nor U48194 (N_48194,N_46949,N_46797);
nand U48195 (N_48195,N_46953,N_46229);
xnor U48196 (N_48196,N_47173,N_46017);
nor U48197 (N_48197,N_46239,N_46734);
nor U48198 (N_48198,N_46409,N_47017);
nand U48199 (N_48199,N_46323,N_47319);
nand U48200 (N_48200,N_46250,N_47450);
or U48201 (N_48201,N_47947,N_46369);
or U48202 (N_48202,N_47658,N_46622);
and U48203 (N_48203,N_46019,N_46334);
or U48204 (N_48204,N_47433,N_46249);
nor U48205 (N_48205,N_47907,N_46127);
nor U48206 (N_48206,N_47444,N_47792);
nand U48207 (N_48207,N_47898,N_46385);
nor U48208 (N_48208,N_46853,N_46310);
nor U48209 (N_48209,N_46849,N_46408);
nand U48210 (N_48210,N_46824,N_47276);
nand U48211 (N_48211,N_47287,N_47305);
nand U48212 (N_48212,N_46586,N_46418);
xor U48213 (N_48213,N_47719,N_47290);
or U48214 (N_48214,N_46744,N_47617);
or U48215 (N_48215,N_46497,N_47602);
nand U48216 (N_48216,N_46642,N_46541);
and U48217 (N_48217,N_47046,N_47122);
nor U48218 (N_48218,N_47425,N_47830);
xor U48219 (N_48219,N_47750,N_46716);
or U48220 (N_48220,N_46236,N_46669);
or U48221 (N_48221,N_47835,N_46106);
nor U48222 (N_48222,N_46556,N_46037);
nor U48223 (N_48223,N_46141,N_47025);
nor U48224 (N_48224,N_46294,N_46612);
and U48225 (N_48225,N_46593,N_47200);
nand U48226 (N_48226,N_47960,N_47771);
and U48227 (N_48227,N_47441,N_47865);
nor U48228 (N_48228,N_46588,N_47726);
and U48229 (N_48229,N_47595,N_46739);
nand U48230 (N_48230,N_46005,N_46516);
or U48231 (N_48231,N_46233,N_47531);
nor U48232 (N_48232,N_46010,N_46449);
nand U48233 (N_48233,N_46494,N_46787);
xnor U48234 (N_48234,N_46545,N_47923);
and U48235 (N_48235,N_46927,N_47486);
xor U48236 (N_48236,N_47714,N_47351);
nand U48237 (N_48237,N_46894,N_46806);
nor U48238 (N_48238,N_47616,N_46117);
xor U48239 (N_48239,N_46446,N_46208);
or U48240 (N_48240,N_46630,N_47229);
nand U48241 (N_48241,N_47615,N_47452);
and U48242 (N_48242,N_47442,N_47191);
nand U48243 (N_48243,N_47682,N_46873);
nor U48244 (N_48244,N_47226,N_47257);
nor U48245 (N_48245,N_46944,N_46802);
nor U48246 (N_48246,N_46974,N_47102);
xor U48247 (N_48247,N_46089,N_46348);
or U48248 (N_48248,N_47042,N_47746);
or U48249 (N_48249,N_47552,N_47417);
nor U48250 (N_48250,N_46414,N_47342);
nand U48251 (N_48251,N_47556,N_46485);
nor U48252 (N_48252,N_46818,N_47095);
xor U48253 (N_48253,N_47567,N_47448);
nor U48254 (N_48254,N_46723,N_46081);
nand U48255 (N_48255,N_46194,N_46360);
nand U48256 (N_48256,N_46468,N_47868);
nor U48257 (N_48257,N_47971,N_46447);
xnor U48258 (N_48258,N_47432,N_47976);
nor U48259 (N_48259,N_47364,N_46453);
or U48260 (N_48260,N_46047,N_47832);
or U48261 (N_48261,N_46370,N_47107);
nand U48262 (N_48262,N_47346,N_46028);
nor U48263 (N_48263,N_47529,N_46053);
nor U48264 (N_48264,N_46531,N_47959);
xnor U48265 (N_48265,N_46951,N_46604);
nand U48266 (N_48266,N_46436,N_47511);
or U48267 (N_48267,N_46055,N_47270);
or U48268 (N_48268,N_46660,N_46632);
nor U48269 (N_48269,N_46337,N_46562);
or U48270 (N_48270,N_47464,N_47999);
nor U48271 (N_48271,N_46182,N_46847);
and U48272 (N_48272,N_47006,N_46301);
nor U48273 (N_48273,N_47203,N_46073);
nand U48274 (N_48274,N_47758,N_47248);
nand U48275 (N_48275,N_46704,N_47834);
nor U48276 (N_48276,N_47674,N_47506);
or U48277 (N_48277,N_47859,N_46721);
or U48278 (N_48278,N_46892,N_47962);
nor U48279 (N_48279,N_47756,N_47031);
xnor U48280 (N_48280,N_47789,N_46544);
nor U48281 (N_48281,N_47877,N_47647);
nand U48282 (N_48282,N_46372,N_46105);
nand U48283 (N_48283,N_46451,N_46965);
and U48284 (N_48284,N_46595,N_47866);
xor U48285 (N_48285,N_47687,N_47334);
xnor U48286 (N_48286,N_46793,N_46121);
nor U48287 (N_48287,N_46116,N_47902);
nand U48288 (N_48288,N_47238,N_46696);
nor U48289 (N_48289,N_47565,N_47528);
and U48290 (N_48290,N_46366,N_46014);
nand U48291 (N_48291,N_47776,N_46137);
nand U48292 (N_48292,N_47412,N_46298);
or U48293 (N_48293,N_46432,N_47851);
and U48294 (N_48294,N_46029,N_46232);
nor U48295 (N_48295,N_46648,N_46045);
nand U48296 (N_48296,N_47690,N_46176);
and U48297 (N_48297,N_47671,N_46820);
nand U48298 (N_48298,N_47398,N_46018);
and U48299 (N_48299,N_46535,N_47164);
xnor U48300 (N_48300,N_46518,N_47455);
xor U48301 (N_48301,N_47026,N_47731);
xor U48302 (N_48302,N_47061,N_47286);
nor U48303 (N_48303,N_47558,N_46068);
xor U48304 (N_48304,N_46478,N_46428);
nand U48305 (N_48305,N_46863,N_46398);
or U48306 (N_48306,N_47375,N_47384);
nor U48307 (N_48307,N_46615,N_46092);
or U48308 (N_48308,N_47483,N_46803);
nand U48309 (N_48309,N_47101,N_47220);
nand U48310 (N_48310,N_47086,N_46546);
or U48311 (N_48311,N_46678,N_46652);
and U48312 (N_48312,N_47734,N_47264);
or U48313 (N_48313,N_46084,N_46324);
or U48314 (N_48314,N_46526,N_46001);
nor U48315 (N_48315,N_46124,N_46277);
and U48316 (N_48316,N_47237,N_47729);
and U48317 (N_48317,N_47382,N_46602);
nor U48318 (N_48318,N_46512,N_47812);
or U48319 (N_48319,N_46259,N_46932);
and U48320 (N_48320,N_46568,N_46059);
or U48321 (N_48321,N_47335,N_47053);
and U48322 (N_48322,N_46715,N_46907);
and U48323 (N_48323,N_47570,N_46243);
or U48324 (N_48324,N_47730,N_47998);
nor U48325 (N_48325,N_47972,N_47623);
or U48326 (N_48326,N_47982,N_46773);
nand U48327 (N_48327,N_47610,N_46430);
nand U48328 (N_48328,N_46700,N_46357);
and U48329 (N_48329,N_47311,N_47621);
nand U48330 (N_48330,N_46411,N_46156);
and U48331 (N_48331,N_46805,N_47440);
nor U48332 (N_48332,N_47542,N_46794);
or U48333 (N_48333,N_46767,N_47419);
or U48334 (N_48334,N_46490,N_46611);
xnor U48335 (N_48335,N_47928,N_47360);
or U48336 (N_48336,N_46748,N_47443);
and U48337 (N_48337,N_46006,N_46049);
nand U48338 (N_48338,N_46759,N_47958);
and U48339 (N_48339,N_47207,N_46038);
or U48340 (N_48340,N_47562,N_46307);
and U48341 (N_48341,N_47967,N_47892);
nor U48342 (N_48342,N_46076,N_46713);
xor U48343 (N_48343,N_47359,N_46085);
or U48344 (N_48344,N_46836,N_46624);
xor U48345 (N_48345,N_46993,N_46605);
nand U48346 (N_48346,N_46811,N_47708);
and U48347 (N_48347,N_47589,N_47576);
nand U48348 (N_48348,N_47739,N_46169);
nand U48349 (N_48349,N_46222,N_46963);
nor U48350 (N_48350,N_46330,N_46050);
nor U48351 (N_48351,N_47136,N_46382);
nor U48352 (N_48352,N_46957,N_46150);
nand U48353 (N_48353,N_47837,N_47536);
nor U48354 (N_48354,N_46935,N_46484);
nor U48355 (N_48355,N_47347,N_47925);
or U48356 (N_48356,N_46561,N_47547);
nor U48357 (N_48357,N_46450,N_47426);
and U48358 (N_48358,N_47548,N_47901);
or U48359 (N_48359,N_47691,N_46911);
nor U48360 (N_48360,N_47427,N_47404);
xnor U48361 (N_48361,N_46683,N_47712);
and U48362 (N_48362,N_47204,N_46048);
nor U48363 (N_48363,N_46162,N_46776);
nand U48364 (N_48364,N_47140,N_46306);
or U48365 (N_48365,N_46371,N_46699);
nor U48366 (N_48366,N_47494,N_47937);
xnor U48367 (N_48367,N_47410,N_47908);
xor U48368 (N_48368,N_47702,N_46766);
nor U48369 (N_48369,N_46126,N_47884);
or U48370 (N_48370,N_46042,N_47018);
or U48371 (N_48371,N_46062,N_47596);
nor U48372 (N_48372,N_46618,N_47760);
xnor U48373 (N_48373,N_46098,N_46185);
or U48374 (N_48374,N_47266,N_47377);
and U48375 (N_48375,N_46032,N_47280);
xor U48376 (N_48376,N_47148,N_46712);
xnor U48377 (N_48377,N_47038,N_46822);
or U48378 (N_48378,N_46131,N_47874);
xor U48379 (N_48379,N_47763,N_46885);
and U48380 (N_48380,N_47460,N_46931);
and U48381 (N_48381,N_47895,N_46262);
or U48382 (N_48382,N_46689,N_47813);
xnor U48383 (N_48383,N_46318,N_47605);
nand U48384 (N_48384,N_46475,N_46256);
nand U48385 (N_48385,N_46355,N_47863);
or U48386 (N_48386,N_47208,N_46936);
or U48387 (N_48387,N_46663,N_47119);
nor U48388 (N_48388,N_47672,N_46674);
nor U48389 (N_48389,N_46720,N_47274);
nand U48390 (N_48390,N_46659,N_46489);
or U48391 (N_48391,N_46564,N_46013);
xor U48392 (N_48392,N_47537,N_47295);
xor U48393 (N_48393,N_46196,N_46655);
nand U48394 (N_48394,N_46078,N_46060);
nand U48395 (N_48395,N_46923,N_47788);
and U48396 (N_48396,N_47386,N_47574);
xor U48397 (N_48397,N_47130,N_47995);
or U48398 (N_48398,N_47391,N_47796);
nor U48399 (N_48399,N_46786,N_46328);
nand U48400 (N_48400,N_46871,N_46890);
nand U48401 (N_48401,N_47498,N_47254);
and U48402 (N_48402,N_47097,N_46331);
nor U48403 (N_48403,N_47161,N_46480);
or U48404 (N_48404,N_47112,N_47612);
or U48405 (N_48405,N_47064,N_47421);
nor U48406 (N_48406,N_46961,N_47804);
nand U48407 (N_48407,N_47676,N_46808);
nand U48408 (N_48408,N_47463,N_47326);
nor U48409 (N_48409,N_47242,N_46731);
nor U48410 (N_48410,N_46976,N_46444);
or U48411 (N_48411,N_47709,N_46870);
or U48412 (N_48412,N_46275,N_47989);
nor U48413 (N_48413,N_47591,N_47392);
and U48414 (N_48414,N_46015,N_46452);
or U48415 (N_48415,N_47036,N_46410);
or U48416 (N_48416,N_46225,N_46869);
xnor U48417 (N_48417,N_47683,N_47040);
or U48418 (N_48418,N_46095,N_46332);
nand U48419 (N_48419,N_47144,N_47109);
or U48420 (N_48420,N_46103,N_46921);
nor U48421 (N_48421,N_46115,N_46729);
and U48422 (N_48422,N_47973,N_46423);
nor U48423 (N_48423,N_47969,N_47648);
xor U48424 (N_48424,N_46523,N_46999);
or U48425 (N_48425,N_46403,N_46413);
or U48426 (N_48426,N_47492,N_46051);
xnor U48427 (N_48427,N_46326,N_47063);
xor U48428 (N_48428,N_47880,N_46350);
nor U48429 (N_48429,N_47198,N_46336);
xnor U48430 (N_48430,N_46897,N_47367);
nor U48431 (N_48431,N_47318,N_46772);
or U48432 (N_48432,N_47127,N_47199);
nor U48433 (N_48433,N_47401,N_47331);
nor U48434 (N_48434,N_47428,N_47843);
nand U48435 (N_48435,N_46732,N_47871);
and U48436 (N_48436,N_47728,N_47493);
or U48437 (N_48437,N_46997,N_46536);
or U48438 (N_48438,N_47438,N_46405);
xnor U48439 (N_48439,N_47785,N_46813);
and U48440 (N_48440,N_46992,N_46938);
nor U48441 (N_48441,N_46390,N_46011);
nand U48442 (N_48442,N_46522,N_47024);
nor U48443 (N_48443,N_46465,N_47631);
and U48444 (N_48444,N_47744,N_46192);
xnor U48445 (N_48445,N_46760,N_47194);
nor U48446 (N_48446,N_47515,N_47039);
xnor U48447 (N_48447,N_47001,N_46777);
nor U48448 (N_48448,N_47252,N_46621);
nor U48449 (N_48449,N_47062,N_46375);
and U48450 (N_48450,N_47963,N_47914);
nor U48451 (N_48451,N_47665,N_46253);
or U48452 (N_48452,N_47655,N_47197);
xnor U48453 (N_48453,N_46835,N_46641);
xor U48454 (N_48454,N_46133,N_47500);
nor U48455 (N_48455,N_46221,N_47000);
and U48456 (N_48456,N_46685,N_46981);
xor U48457 (N_48457,N_46389,N_47684);
nor U48458 (N_48458,N_47607,N_46668);
nor U48459 (N_48459,N_46664,N_47139);
xor U48460 (N_48460,N_47126,N_46661);
nand U48461 (N_48461,N_47175,N_47313);
and U48462 (N_48462,N_46527,N_46972);
and U48463 (N_48463,N_47059,N_47422);
or U48464 (N_48464,N_47291,N_46631);
and U48465 (N_48465,N_46378,N_46529);
nor U48466 (N_48466,N_47688,N_47241);
and U48467 (N_48467,N_47371,N_47424);
or U48468 (N_48468,N_47523,N_47541);
or U48469 (N_48469,N_47585,N_46164);
and U48470 (N_48470,N_47023,N_46821);
xor U48471 (N_48471,N_47979,N_47961);
nand U48472 (N_48472,N_47779,N_46841);
nor U48473 (N_48473,N_46858,N_46244);
and U48474 (N_48474,N_47519,N_46677);
or U48475 (N_48475,N_47256,N_47675);
or U48476 (N_48476,N_47474,N_46138);
nor U48477 (N_48477,N_46702,N_47573);
nor U48478 (N_48478,N_46474,N_46148);
and U48479 (N_48479,N_47399,N_47820);
nor U48480 (N_48480,N_47210,N_47356);
nor U48481 (N_48481,N_47948,N_46486);
nand U48482 (N_48482,N_46859,N_47705);
and U48483 (N_48483,N_47852,N_47790);
or U48484 (N_48484,N_47048,N_46139);
nand U48485 (N_48485,N_46422,N_46481);
nand U48486 (N_48486,N_47850,N_47535);
and U48487 (N_48487,N_46107,N_47190);
nand U48488 (N_48488,N_47125,N_46425);
xor U48489 (N_48489,N_46838,N_46851);
xor U48490 (N_48490,N_47488,N_47363);
nor U48491 (N_48491,N_46796,N_47662);
nand U48492 (N_48492,N_46563,N_47720);
or U48493 (N_48493,N_47521,N_47193);
nand U48494 (N_48494,N_46519,N_46002);
and U48495 (N_48495,N_47632,N_47707);
and U48496 (N_48496,N_47255,N_46800);
nand U48497 (N_48497,N_47564,N_46231);
nor U48498 (N_48498,N_47325,N_47035);
or U48499 (N_48499,N_46533,N_47991);
and U48500 (N_48500,N_47108,N_46788);
xnor U48501 (N_48501,N_47532,N_47477);
nand U48502 (N_48502,N_46057,N_46186);
or U48503 (N_48503,N_46629,N_46574);
or U48504 (N_48504,N_47277,N_47016);
xor U48505 (N_48505,N_46266,N_47913);
or U48506 (N_48506,N_47667,N_46942);
and U48507 (N_48507,N_47659,N_47872);
nand U48508 (N_48508,N_47341,N_47380);
nor U48509 (N_48509,N_47845,N_47653);
xor U48510 (N_48510,N_46364,N_46174);
or U48511 (N_48511,N_47650,N_47008);
nand U48512 (N_48512,N_46693,N_47004);
nand U48513 (N_48513,N_47879,N_47214);
nand U48514 (N_48514,N_47508,N_46532);
nand U48515 (N_48515,N_46027,N_46617);
and U48516 (N_48516,N_47600,N_47698);
and U48517 (N_48517,N_47590,N_46577);
nor U48518 (N_48518,N_46968,N_47100);
and U48519 (N_48519,N_46171,N_47754);
nor U48520 (N_48520,N_46207,N_47723);
nor U48521 (N_48521,N_46608,N_46872);
and U48522 (N_48522,N_47899,N_47250);
and U48523 (N_48523,N_47378,N_47296);
or U48524 (N_48524,N_46270,N_46769);
xor U48525 (N_48525,N_46437,N_46308);
and U48526 (N_48526,N_47466,N_46136);
nor U48527 (N_48527,N_46210,N_47389);
nand U48528 (N_48528,N_46471,N_47915);
and U48529 (N_48529,N_46412,N_47449);
nand U48530 (N_48530,N_46742,N_46329);
xor U48531 (N_48531,N_47131,N_46754);
or U48532 (N_48532,N_47470,N_46012);
xor U48533 (N_48533,N_47105,N_47652);
nand U48534 (N_48534,N_47878,N_47604);
xor U48535 (N_48535,N_47115,N_46812);
or U48536 (N_48536,N_47736,N_47043);
nand U48537 (N_48537,N_46924,N_46108);
nand U48538 (N_48538,N_47165,N_46099);
nand U48539 (N_48539,N_47782,N_47225);
or U48540 (N_48540,N_46569,N_46093);
nor U48541 (N_48541,N_47124,N_46673);
xor U48542 (N_48542,N_47974,N_46646);
nand U48543 (N_48543,N_46129,N_47586);
and U48544 (N_48544,N_47807,N_46929);
and U48545 (N_48545,N_47966,N_47458);
and U48546 (N_48546,N_46576,N_47293);
or U48547 (N_48547,N_46320,N_47700);
nor U48548 (N_48548,N_46765,N_46580);
or U48549 (N_48549,N_46592,N_47103);
or U48550 (N_48550,N_46980,N_46675);
nor U48551 (N_48551,N_46213,N_47633);
nor U48552 (N_48552,N_46388,N_46782);
nand U48553 (N_48553,N_47680,N_46879);
nor U48554 (N_48554,N_46846,N_47021);
or U48555 (N_48555,N_47988,N_46509);
xnor U48556 (N_48556,N_46165,N_46134);
xnor U48557 (N_48557,N_46296,N_47869);
and U48558 (N_48558,N_47641,N_46876);
or U48559 (N_48559,N_46227,N_46967);
nor U48560 (N_48560,N_47333,N_46686);
and U48561 (N_48561,N_46188,N_47465);
or U48562 (N_48562,N_46035,N_47366);
xnor U48563 (N_48563,N_46855,N_46039);
and U48564 (N_48564,N_46271,N_47397);
nor U48565 (N_48565,N_47580,N_46538);
nor U48566 (N_48566,N_47457,N_47886);
nand U48567 (N_48567,N_47298,N_46386);
and U48568 (N_48568,N_47087,N_46377);
nand U48569 (N_48569,N_46083,N_46483);
and U48570 (N_48570,N_47085,N_47745);
and U48571 (N_48571,N_47308,N_47587);
and U48572 (N_48572,N_47613,N_46000);
or U48573 (N_48573,N_46052,N_46954);
nor U48574 (N_48574,N_47727,N_47049);
nand U48575 (N_48575,N_47501,N_46817);
nor U48576 (N_48576,N_46790,N_46501);
xor U48577 (N_48577,N_46205,N_47926);
xnor U48578 (N_48578,N_46850,N_46634);
nand U48579 (N_48579,N_47476,N_47530);
nand U48580 (N_48580,N_46426,N_47388);
nand U48581 (N_48581,N_46607,N_47507);
xor U48582 (N_48582,N_46276,N_46680);
or U48583 (N_48583,N_46299,N_46964);
nand U48584 (N_48584,N_47661,N_46539);
or U48585 (N_48585,N_46087,N_47155);
xnor U48586 (N_48586,N_46297,N_47236);
xor U48587 (N_48587,N_46036,N_46147);
nand U48588 (N_48588,N_46473,N_47158);
or U48589 (N_48589,N_46865,N_46904);
or U48590 (N_48590,N_47050,N_46376);
and U48591 (N_48591,N_47446,N_46211);
xor U48592 (N_48592,N_47439,N_46514);
or U48593 (N_48593,N_47068,N_47677);
nor U48594 (N_48594,N_46247,N_46191);
nand U48595 (N_48595,N_47956,N_47478);
or U48596 (N_48596,N_47560,N_47258);
nand U48597 (N_48597,N_46187,N_46456);
nor U48598 (N_48598,N_46780,N_46462);
xor U48599 (N_48599,N_46864,N_47260);
and U48600 (N_48600,N_47649,N_47598);
xnor U48601 (N_48601,N_47626,N_47075);
nor U48602 (N_48602,N_47454,N_46753);
xnor U48603 (N_48603,N_46125,N_47630);
nand U48604 (N_48604,N_46441,N_46197);
nand U48605 (N_48605,N_46990,N_46733);
xor U48606 (N_48606,N_46614,N_46503);
or U48607 (N_48607,N_47065,N_47883);
and U48608 (N_48608,N_47304,N_46815);
or U48609 (N_48609,N_46195,N_47681);
xnor U48610 (N_48610,N_46145,N_46804);
nor U48611 (N_48611,N_46282,N_47894);
nor U48612 (N_48612,N_46067,N_46579);
xnor U48613 (N_48613,N_47808,N_47221);
and U48614 (N_48614,N_47867,N_47534);
xor U48615 (N_48615,N_47854,N_46248);
xnor U48616 (N_48616,N_46952,N_47935);
nand U48617 (N_48617,N_47014,N_47078);
xor U48618 (N_48618,N_46341,N_46708);
xor U48619 (N_48619,N_47762,N_46043);
and U48620 (N_48620,N_46799,N_46620);
xor U48621 (N_48621,N_47888,N_46898);
and U48622 (N_48622,N_46146,N_46402);
and U48623 (N_48623,N_46316,N_46218);
nor U48624 (N_48624,N_46460,N_46801);
nand U48625 (N_48625,N_46571,N_46391);
and U48626 (N_48626,N_46255,N_47201);
and U48627 (N_48627,N_47265,N_47864);
nor U48628 (N_48628,N_46606,N_47777);
xnor U48629 (N_48629,N_46694,N_47407);
or U48630 (N_48630,N_47724,N_46970);
nor U48631 (N_48631,N_46267,N_46901);
nor U48632 (N_48632,N_46401,N_46429);
nand U48633 (N_48633,N_47370,N_46896);
or U48634 (N_48634,N_46322,N_46300);
xor U48635 (N_48635,N_46774,N_46381);
nor U48636 (N_48636,N_47773,N_46570);
xnor U48637 (N_48637,N_47456,N_46823);
nand U48638 (N_48638,N_46004,N_46540);
or U48639 (N_48639,N_47931,N_46178);
xnor U48640 (N_48640,N_47627,N_47379);
or U48641 (N_48641,N_46295,N_46325);
or U48642 (N_48642,N_47920,N_46166);
or U48643 (N_48643,N_46104,N_47847);
nor U48644 (N_48644,N_46848,N_46111);
and U48645 (N_48645,N_47862,N_46584);
xnor U48646 (N_48646,N_47601,N_47373);
or U48647 (N_48647,N_46387,N_47174);
or U48648 (N_48648,N_46639,N_46144);
or U48649 (N_48649,N_46705,N_46827);
or U48650 (N_48650,N_46691,N_46353);
nand U48651 (N_48651,N_46551,N_47396);
xor U48652 (N_48652,N_46177,N_46335);
or U48653 (N_48653,N_47748,N_47765);
or U48654 (N_48654,N_47390,N_46524);
and U48655 (N_48655,N_47209,N_46837);
and U48656 (N_48656,N_47810,N_47619);
xnor U48657 (N_48657,N_46940,N_47368);
and U48658 (N_48658,N_47271,N_46996);
xnor U48659 (N_48659,N_47606,N_47579);
xor U48660 (N_48660,N_46507,N_47752);
and U48661 (N_48661,N_46819,N_47783);
and U48662 (N_48662,N_47120,N_46941);
xnor U48663 (N_48663,N_46399,N_46442);
nand U48664 (N_48664,N_46775,N_47575);
nand U48665 (N_48665,N_46419,N_46181);
or U48666 (N_48666,N_46258,N_46756);
nor U48667 (N_48667,N_47232,N_46505);
or U48668 (N_48668,N_47117,N_46470);
xnor U48669 (N_48669,N_46933,N_47805);
and U48670 (N_48670,N_47234,N_46315);
nor U48671 (N_48671,N_47393,N_47890);
xor U48672 (N_48672,N_46140,N_47411);
xnor U48673 (N_48673,N_46071,N_46305);
nand U48674 (N_48674,N_47233,N_47663);
or U48675 (N_48675,N_47873,N_47057);
xnor U48676 (N_48676,N_46877,N_47929);
nand U48677 (N_48677,N_47468,N_46168);
and U48678 (N_48678,N_47374,N_47073);
and U48679 (N_48679,N_47350,N_46317);
nand U48680 (N_48680,N_46066,N_46431);
xor U48681 (N_48681,N_46206,N_46573);
nor U48682 (N_48682,N_47079,N_47145);
and U48683 (N_48683,N_46293,N_47836);
nand U48684 (N_48684,N_46264,N_47897);
or U48685 (N_48685,N_46814,N_47045);
xnor U48686 (N_48686,N_47292,N_46238);
xnor U48687 (N_48687,N_46420,N_47437);
xnor U48688 (N_48688,N_47354,N_46077);
nor U48689 (N_48689,N_46088,N_47030);
and U48690 (N_48690,N_46726,N_47344);
nor U48691 (N_48691,N_46962,N_46212);
nand U48692 (N_48692,N_47051,N_47514);
and U48693 (N_48693,N_47009,N_47077);
nand U48694 (N_48694,N_47300,N_47968);
nor U48695 (N_48695,N_47123,N_46183);
xor U48696 (N_48696,N_46314,N_47975);
and U48697 (N_48697,N_47504,N_46874);
xnor U48698 (N_48698,N_46789,N_46504);
and U48699 (N_48699,N_47625,N_47977);
nor U48700 (N_48700,N_46809,N_47020);
and U48701 (N_48701,N_47451,N_46454);
and U48702 (N_48702,N_47853,N_46180);
and U48703 (N_48703,N_47987,N_47518);
nor U48704 (N_48704,N_46875,N_47634);
nand U48705 (N_48705,N_47005,N_47911);
nand U48706 (N_48706,N_46644,N_46286);
nor U48707 (N_48707,N_47096,N_46922);
xnor U48708 (N_48708,N_46457,N_46559);
nand U48709 (N_48709,N_47509,N_46349);
nor U48710 (N_48710,N_46204,N_47083);
and U48711 (N_48711,N_47336,N_46798);
xnor U48712 (N_48712,N_47032,N_46488);
nor U48713 (N_48713,N_46217,N_47082);
nor U48714 (N_48714,N_47811,N_47141);
or U48715 (N_48715,N_46492,N_47044);
and U48716 (N_48716,N_46628,N_46687);
nand U48717 (N_48717,N_46567,N_47849);
or U48718 (N_48718,N_46727,N_47262);
xor U48719 (N_48719,N_46118,N_47986);
xor U48720 (N_48720,N_46613,N_47058);
nand U48721 (N_48721,N_46082,N_46190);
nand U48722 (N_48722,N_46785,N_46074);
or U48723 (N_48723,N_47946,N_47160);
nand U48724 (N_48724,N_47893,N_47801);
nor U48725 (N_48725,N_46344,N_46672);
or U48726 (N_48726,N_46290,N_47706);
nor U48727 (N_48727,N_47526,N_46303);
or U48728 (N_48728,N_47609,N_46203);
nor U48729 (N_48729,N_46667,N_47732);
nand U48730 (N_48730,N_47135,N_47462);
or U48731 (N_48731,N_47343,N_47028);
or U48732 (N_48732,N_47934,N_47459);
nand U48733 (N_48733,N_47656,N_47806);
nor U48734 (N_48734,N_46603,N_47740);
or U48735 (N_48735,N_47767,N_46955);
or U48736 (N_48736,N_46268,N_46747);
nand U48737 (N_48737,N_47566,N_46991);
and U48738 (N_48738,N_47132,N_47090);
or U48739 (N_48739,N_47110,N_46920);
xor U48740 (N_48740,N_47480,N_46120);
nand U48741 (N_48741,N_46891,N_47299);
xor U48742 (N_48742,N_46662,N_46770);
nor U48743 (N_48743,N_47353,N_46416);
xnor U48744 (N_48744,N_46384,N_46246);
nor U48745 (N_48745,N_46626,N_47584);
nor U48746 (N_48746,N_46979,N_46417);
xnor U48747 (N_48747,N_47309,N_46548);
nor U48748 (N_48748,N_46982,N_46928);
and U48749 (N_48749,N_46064,N_46917);
nor U48750 (N_48750,N_47282,N_46506);
nand U48751 (N_48751,N_47955,N_46596);
nor U48752 (N_48752,N_47142,N_46400);
nand U48753 (N_48753,N_47766,N_47187);
and U48754 (N_48754,N_47162,N_46625);
or U48755 (N_48755,N_46834,N_46755);
or U48756 (N_48756,N_46499,N_47307);
and U48757 (N_48757,N_47002,N_46695);
nor U48758 (N_48758,N_47906,N_46333);
and U48759 (N_48759,N_46283,N_47010);
xnor U48760 (N_48760,N_47933,N_46945);
nand U48761 (N_48761,N_46966,N_46637);
nand U48762 (N_48762,N_47770,N_47568);
or U48763 (N_48763,N_47403,N_47944);
nor U48764 (N_48764,N_47553,N_47408);
nor U48765 (N_48765,N_47555,N_47725);
nor U48766 (N_48766,N_46362,N_47643);
nor U48767 (N_48767,N_47559,N_46757);
nand U48768 (N_48768,N_46934,N_47143);
nor U48769 (N_48769,N_46061,N_46771);
nor U48770 (N_48770,N_47239,N_46396);
nand U48771 (N_48771,N_47793,N_46101);
nor U48772 (N_48772,N_46100,N_46351);
nand U48773 (N_48773,N_47546,N_47352);
nor U48774 (N_48774,N_46302,N_46383);
xnor U48775 (N_48775,N_46511,N_47764);
and U48776 (N_48776,N_46199,N_46269);
nand U48777 (N_48777,N_47416,N_47027);
or U48778 (N_48778,N_47060,N_46925);
nand U48779 (N_48779,N_46393,N_47941);
and U48780 (N_48780,N_47497,N_47487);
and U48781 (N_48781,N_47916,N_46701);
and U48782 (N_48782,N_47376,N_47978);
nor U48783 (N_48783,N_47800,N_46016);
nor U48784 (N_48784,N_47540,N_46986);
nor U48785 (N_48785,N_46913,N_47394);
and U48786 (N_48786,N_46946,N_47022);
xor U48787 (N_48787,N_46365,N_47557);
or U48788 (N_48788,N_46717,N_46342);
and U48789 (N_48789,N_47786,N_46919);
nor U48790 (N_48790,N_46844,N_47339);
nor U48791 (N_48791,N_46128,N_46987);
xor U48792 (N_48792,N_46816,N_46472);
nand U48793 (N_48793,N_47213,N_46649);
xnor U48794 (N_48794,N_46021,N_47385);
nand U48795 (N_48795,N_46070,N_46354);
nand U48796 (N_48796,N_46030,N_47828);
nand U48797 (N_48797,N_47735,N_46477);
nand U48798 (N_48798,N_47429,N_46007);
and U48799 (N_48799,N_47316,N_46228);
nor U48800 (N_48800,N_47825,N_46718);
nor U48801 (N_48801,N_47240,N_46251);
nor U48802 (N_48802,N_47205,N_47150);
nand U48803 (N_48803,N_47990,N_47315);
xnor U48804 (N_48804,N_47163,N_46455);
nor U48805 (N_48805,N_46581,N_46510);
nand U48806 (N_48806,N_47369,N_47945);
or U48807 (N_48807,N_47151,N_46884);
xor U48808 (N_48808,N_47917,N_46597);
nor U48809 (N_48809,N_47314,N_47741);
nor U48810 (N_48810,N_47699,N_46601);
nand U48811 (N_48811,N_47402,N_46676);
or U48812 (N_48812,N_47996,N_47246);
or U48813 (N_48813,N_47778,N_46547);
or U48814 (N_48814,N_47664,N_47860);
and U48815 (N_48815,N_47692,N_47081);
nor U48816 (N_48816,N_47571,N_46003);
or U48817 (N_48817,N_47003,N_47195);
and U48818 (N_48818,N_46719,N_47809);
and U48819 (N_48819,N_46887,N_46216);
xnor U48820 (N_48820,N_46279,N_47244);
xor U48821 (N_48821,N_47775,N_47981);
and U48822 (N_48822,N_46214,N_47679);
or U48823 (N_48823,N_46638,N_47041);
xor U48824 (N_48824,N_46234,N_46761);
and U48825 (N_48825,N_47037,N_46889);
and U48826 (N_48826,N_46943,N_46363);
and U48827 (N_48827,N_46151,N_47329);
and U48828 (N_48828,N_46710,N_46831);
xor U48829 (N_48829,N_46367,N_46860);
or U48830 (N_48830,N_46054,N_47453);
xor U48831 (N_48831,N_46459,N_46023);
xnor U48832 (N_48832,N_47733,N_47128);
nor U48833 (N_48833,N_47992,N_47721);
nor U48834 (N_48834,N_47272,N_46198);
xnor U48835 (N_48835,N_47328,N_47802);
xnor U48836 (N_48836,N_46288,N_46671);
and U48837 (N_48837,N_47383,N_47932);
or U48838 (N_48838,N_47618,N_46242);
nand U48839 (N_48839,N_47269,N_46491);
and U48840 (N_48840,N_47159,N_46311);
or U48841 (N_48841,N_46861,N_46750);
xnor U48842 (N_48842,N_47312,N_47980);
nor U48843 (N_48843,N_46623,N_46274);
nand U48844 (N_48844,N_46998,N_47227);
xnor U48845 (N_48845,N_47829,N_47517);
or U48846 (N_48846,N_47178,N_47569);
and U48847 (N_48847,N_46745,N_47072);
or U48848 (N_48848,N_47624,N_46265);
xor U48849 (N_48849,N_47856,N_46161);
nand U48850 (N_48850,N_46482,N_47267);
nor U48851 (N_48851,N_46424,N_46670);
nand U48852 (N_48852,N_47761,N_47147);
xnor U48853 (N_48853,N_47467,N_47471);
nand U48854 (N_48854,N_46159,N_47539);
nand U48855 (N_48855,N_47718,N_46550);
nor U48856 (N_48856,N_47545,N_47646);
nor U48857 (N_48857,N_46502,N_47704);
and U48858 (N_48858,N_47301,N_47827);
nor U48859 (N_48859,N_46666,N_47243);
xor U48860 (N_48860,N_46900,N_46397);
nand U48861 (N_48861,N_46647,N_46868);
nand U48862 (N_48862,N_46857,N_46781);
xor U48863 (N_48863,N_47694,N_46160);
nand U48864 (N_48864,N_46724,N_46319);
nand U48865 (N_48865,N_46114,N_46610);
and U48866 (N_48866,N_46572,N_46886);
nand U48867 (N_48867,N_46703,N_46273);
nor U48868 (N_48868,N_47469,N_47550);
or U48869 (N_48869,N_46598,N_47533);
nand U48870 (N_48870,N_46097,N_46843);
or U48871 (N_48871,N_46312,N_47685);
and U48872 (N_48872,N_46130,N_46643);
nor U48873 (N_48873,N_47186,N_47543);
or U48874 (N_48874,N_47330,N_46515);
nand U48875 (N_48875,N_47970,N_46379);
xor U48876 (N_48876,N_47168,N_46866);
xor U48877 (N_48877,N_46433,N_46960);
xnor U48878 (N_48878,N_46697,N_46566);
nor U48879 (N_48879,N_47954,N_47875);
xnor U48880 (N_48880,N_47561,N_46407);
xnor U48881 (N_48881,N_47831,N_47047);
and U48882 (N_48882,N_46707,N_46122);
nand U48883 (N_48883,N_47345,N_47012);
xnor U48884 (N_48884,N_46743,N_46565);
and U48885 (N_48885,N_47435,N_47092);
nand U48886 (N_48886,N_46469,N_46909);
or U48887 (N_48887,N_47503,N_47278);
and U48888 (N_48888,N_46985,N_46395);
or U48889 (N_48889,N_47993,N_47310);
nand U48890 (N_48890,N_47146,N_47505);
nand U48891 (N_48891,N_47289,N_46916);
or U48892 (N_48892,N_47715,N_47711);
or U48893 (N_48893,N_47074,N_46591);
or U48894 (N_48894,N_46768,N_47157);
or U48895 (N_48895,N_47512,N_46905);
nand U48896 (N_48896,N_47395,N_46041);
or U48897 (N_48897,N_47717,N_46764);
or U48898 (N_48898,N_46530,N_47994);
nor U48899 (N_48899,N_46735,N_46096);
and U48900 (N_48900,N_47909,N_46220);
xor U48901 (N_48901,N_47185,N_46112);
xnor U48902 (N_48902,N_46711,N_46537);
nand U48903 (N_48903,N_46679,N_47321);
nor U48904 (N_48904,N_47231,N_47279);
xor U48905 (N_48905,N_46200,N_46158);
or U48906 (N_48906,N_46280,N_47219);
xor U48907 (N_48907,N_46558,N_46056);
nor U48908 (N_48908,N_46440,N_47848);
nor U48909 (N_48909,N_47817,N_47608);
and U48910 (N_48910,N_46261,N_47673);
or U48911 (N_48911,N_47302,N_47900);
nand U48912 (N_48912,N_47212,N_47104);
and U48913 (N_48913,N_46948,N_47332);
xnor U48914 (N_48914,N_46163,N_47855);
nand U48915 (N_48915,N_46292,N_46508);
xor U48916 (N_48916,N_47111,N_46751);
or U48917 (N_48917,N_47882,N_47846);
nor U48918 (N_48918,N_46257,N_46415);
or U48919 (N_48919,N_47516,N_47919);
and U48920 (N_48920,N_46065,N_47481);
nand U48921 (N_48921,N_47593,N_46072);
nand U48922 (N_48922,N_47400,N_46969);
or U48923 (N_48923,N_47118,N_46493);
xor U48924 (N_48924,N_47525,N_46427);
or U48925 (N_48925,N_47387,N_47774);
xnor U48926 (N_48926,N_46421,N_47814);
xor U48927 (N_48927,N_47154,N_47116);
nand U48928 (N_48928,N_46155,N_47614);
nor U48929 (N_48929,N_46031,N_47052);
and U48930 (N_48930,N_47826,N_47180);
and U48931 (N_48931,N_46778,N_46392);
nor U48932 (N_48932,N_47611,N_46102);
nand U48933 (N_48933,N_47578,N_46075);
nand U48934 (N_48934,N_47235,N_46807);
nor U48935 (N_48935,N_46044,N_47054);
nand U48936 (N_48936,N_47357,N_46736);
xnor U48937 (N_48937,N_47738,N_46345);
nand U48938 (N_48938,N_47918,N_47645);
nand U48939 (N_48939,N_47217,N_47228);
nor U48940 (N_48940,N_46926,N_47355);
and U48941 (N_48941,N_47423,N_47479);
and U48942 (N_48942,N_47554,N_46240);
and U48943 (N_48943,N_47984,N_46090);
nand U48944 (N_48944,N_46525,N_46830);
nand U48945 (N_48945,N_47181,N_47840);
xor U48946 (N_48946,N_46309,N_46912);
or U48947 (N_48947,N_47841,N_46209);
nand U48948 (N_48948,N_47697,N_47524);
or U48949 (N_48949,N_46252,N_47772);
and U48950 (N_48950,N_46026,N_47637);
and U48951 (N_48951,N_46839,N_47094);
nor U48952 (N_48952,N_47759,N_47710);
nor U48953 (N_48953,N_47818,N_46445);
or U48954 (N_48954,N_47644,N_46149);
and U48955 (N_48955,N_47015,N_47249);
nand U48956 (N_48956,N_46658,N_47842);
xor U48957 (N_48957,N_47749,N_46553);
or U48958 (N_48958,N_47797,N_46304);
and U48959 (N_48959,N_47660,N_47876);
and U48960 (N_48960,N_46977,N_46224);
nand U48961 (N_48961,N_46352,N_47930);
or U48962 (N_48962,N_46825,N_47361);
nand U48963 (N_48963,N_46959,N_47693);
xor U48964 (N_48964,N_47223,N_46895);
or U48965 (N_48965,N_47499,N_46179);
nand U48966 (N_48966,N_47798,N_46783);
nand U48967 (N_48967,N_46521,N_47844);
or U48968 (N_48968,N_46542,N_47538);
nand U48969 (N_48969,N_46291,N_47055);
nor U48970 (N_48970,N_47171,N_46883);
nor U48971 (N_48971,N_47406,N_46517);
and U48972 (N_48972,N_47588,N_46587);
nor U48973 (N_48973,N_46173,N_46069);
nor U48974 (N_48974,N_47716,N_46681);
nand U48975 (N_48975,N_46549,N_47067);
or U48976 (N_48976,N_47177,N_46260);
or U48977 (N_48977,N_46575,N_47833);
nor U48978 (N_48978,N_47281,N_47172);
or U48979 (N_48979,N_47066,N_46500);
xnor U48980 (N_48980,N_46709,N_47737);
or U48981 (N_48981,N_47106,N_47192);
nor U48982 (N_48982,N_46495,N_47520);
and U48983 (N_48983,N_46758,N_47620);
and U48984 (N_48984,N_46749,N_47420);
nor U48985 (N_48985,N_46347,N_47881);
nand U48986 (N_48986,N_46346,N_47816);
or U48987 (N_48987,N_46640,N_47405);
nand U48988 (N_48988,N_46654,N_46237);
xor U48989 (N_48989,N_46845,N_47409);
nor U48990 (N_48990,N_46313,N_46600);
or U48991 (N_48991,N_46189,N_47113);
xor U48992 (N_48992,N_46888,N_46009);
xor U48993 (N_48993,N_46461,N_46022);
xor U48994 (N_48994,N_47152,N_46599);
nor U48995 (N_48995,N_46167,N_46880);
xor U48996 (N_48996,N_47247,N_47686);
xor U48997 (N_48997,N_46230,N_46762);
xnor U48998 (N_48998,N_47887,N_46466);
or U48999 (N_48999,N_47196,N_47642);
xor U49000 (N_49000,N_46379,N_46827);
and U49001 (N_49001,N_47287,N_46476);
or U49002 (N_49002,N_46780,N_46592);
nand U49003 (N_49003,N_47962,N_47334);
nor U49004 (N_49004,N_47032,N_47297);
or U49005 (N_49005,N_47755,N_46220);
xnor U49006 (N_49006,N_46482,N_46513);
or U49007 (N_49007,N_47068,N_46401);
nand U49008 (N_49008,N_46799,N_46496);
nand U49009 (N_49009,N_47492,N_47267);
xor U49010 (N_49010,N_47177,N_46254);
xnor U49011 (N_49011,N_47602,N_46189);
and U49012 (N_49012,N_47578,N_47276);
xor U49013 (N_49013,N_47208,N_46081);
or U49014 (N_49014,N_47361,N_46360);
and U49015 (N_49015,N_46221,N_46620);
and U49016 (N_49016,N_47931,N_46658);
and U49017 (N_49017,N_47455,N_46781);
xnor U49018 (N_49018,N_47631,N_46028);
nor U49019 (N_49019,N_46711,N_46352);
and U49020 (N_49020,N_47573,N_47574);
xor U49021 (N_49021,N_46410,N_47596);
nor U49022 (N_49022,N_46812,N_47370);
xnor U49023 (N_49023,N_47395,N_47162);
nor U49024 (N_49024,N_46833,N_47566);
and U49025 (N_49025,N_47610,N_46995);
nor U49026 (N_49026,N_46310,N_47091);
or U49027 (N_49027,N_47588,N_47568);
nand U49028 (N_49028,N_46061,N_47759);
xor U49029 (N_49029,N_46768,N_47563);
xnor U49030 (N_49030,N_47745,N_47353);
or U49031 (N_49031,N_47930,N_46542);
nor U49032 (N_49032,N_47185,N_46678);
xor U49033 (N_49033,N_46111,N_46055);
xor U49034 (N_49034,N_47708,N_47934);
or U49035 (N_49035,N_47123,N_46595);
nand U49036 (N_49036,N_46008,N_47113);
and U49037 (N_49037,N_46118,N_47332);
and U49038 (N_49038,N_47742,N_46210);
xnor U49039 (N_49039,N_47433,N_46693);
xnor U49040 (N_49040,N_46389,N_47833);
xnor U49041 (N_49041,N_47153,N_47815);
and U49042 (N_49042,N_46615,N_47757);
nor U49043 (N_49043,N_47424,N_47173);
and U49044 (N_49044,N_47325,N_47511);
nand U49045 (N_49045,N_46554,N_47225);
nand U49046 (N_49046,N_46967,N_47784);
nand U49047 (N_49047,N_47293,N_47989);
xor U49048 (N_49048,N_46724,N_46268);
nand U49049 (N_49049,N_47590,N_47154);
xor U49050 (N_49050,N_47346,N_47179);
and U49051 (N_49051,N_47747,N_46850);
and U49052 (N_49052,N_46434,N_47288);
and U49053 (N_49053,N_47325,N_47639);
nand U49054 (N_49054,N_47131,N_46274);
xnor U49055 (N_49055,N_46601,N_47884);
nand U49056 (N_49056,N_46961,N_46245);
nand U49057 (N_49057,N_46372,N_46614);
or U49058 (N_49058,N_47091,N_47060);
or U49059 (N_49059,N_47093,N_46515);
or U49060 (N_49060,N_46848,N_46687);
and U49061 (N_49061,N_46412,N_47890);
and U49062 (N_49062,N_46450,N_46934);
xnor U49063 (N_49063,N_47359,N_47376);
nand U49064 (N_49064,N_46093,N_46937);
and U49065 (N_49065,N_47883,N_46600);
and U49066 (N_49066,N_47823,N_46009);
or U49067 (N_49067,N_47068,N_47487);
nand U49068 (N_49068,N_47433,N_46124);
and U49069 (N_49069,N_47169,N_47358);
or U49070 (N_49070,N_47401,N_46899);
nor U49071 (N_49071,N_47247,N_46357);
xnor U49072 (N_49072,N_47736,N_47645);
and U49073 (N_49073,N_47795,N_46926);
and U49074 (N_49074,N_46806,N_47030);
or U49075 (N_49075,N_46732,N_47235);
or U49076 (N_49076,N_47136,N_46679);
or U49077 (N_49077,N_47637,N_46656);
nand U49078 (N_49078,N_47436,N_47168);
and U49079 (N_49079,N_46195,N_46210);
nand U49080 (N_49080,N_47678,N_47997);
and U49081 (N_49081,N_46846,N_46798);
nor U49082 (N_49082,N_46413,N_46795);
xor U49083 (N_49083,N_46100,N_47865);
nand U49084 (N_49084,N_46043,N_46177);
or U49085 (N_49085,N_47502,N_47729);
or U49086 (N_49086,N_47361,N_47216);
or U49087 (N_49087,N_47115,N_46207);
or U49088 (N_49088,N_47262,N_46628);
xnor U49089 (N_49089,N_47939,N_47629);
or U49090 (N_49090,N_47286,N_46430);
nand U49091 (N_49091,N_46650,N_47658);
xnor U49092 (N_49092,N_47043,N_46976);
and U49093 (N_49093,N_47674,N_47786);
or U49094 (N_49094,N_47114,N_46928);
or U49095 (N_49095,N_47905,N_46901);
nand U49096 (N_49096,N_46350,N_46688);
nor U49097 (N_49097,N_46117,N_47327);
xor U49098 (N_49098,N_47666,N_46327);
or U49099 (N_49099,N_47467,N_46643);
or U49100 (N_49100,N_46774,N_46725);
xnor U49101 (N_49101,N_46511,N_46713);
nand U49102 (N_49102,N_47718,N_46908);
xnor U49103 (N_49103,N_47482,N_47585);
nand U49104 (N_49104,N_47778,N_46626);
nor U49105 (N_49105,N_46886,N_47555);
or U49106 (N_49106,N_46062,N_46015);
nor U49107 (N_49107,N_47349,N_47667);
and U49108 (N_49108,N_46098,N_47711);
nor U49109 (N_49109,N_47085,N_46972);
nor U49110 (N_49110,N_47250,N_47684);
xor U49111 (N_49111,N_47082,N_46052);
or U49112 (N_49112,N_47689,N_46199);
or U49113 (N_49113,N_47133,N_47977);
and U49114 (N_49114,N_46029,N_46958);
nand U49115 (N_49115,N_47029,N_46589);
or U49116 (N_49116,N_47884,N_47417);
nand U49117 (N_49117,N_46023,N_47439);
xor U49118 (N_49118,N_47158,N_46882);
nor U49119 (N_49119,N_46005,N_47450);
nor U49120 (N_49120,N_46241,N_47605);
xnor U49121 (N_49121,N_47696,N_46271);
xnor U49122 (N_49122,N_46942,N_46373);
nor U49123 (N_49123,N_46813,N_47193);
nand U49124 (N_49124,N_47055,N_46895);
or U49125 (N_49125,N_47233,N_47940);
and U49126 (N_49126,N_46545,N_47609);
xor U49127 (N_49127,N_47869,N_46389);
and U49128 (N_49128,N_46617,N_47163);
and U49129 (N_49129,N_46228,N_46494);
nor U49130 (N_49130,N_46893,N_46423);
nand U49131 (N_49131,N_46811,N_47354);
xnor U49132 (N_49132,N_46006,N_47679);
xnor U49133 (N_49133,N_47109,N_46621);
nor U49134 (N_49134,N_46067,N_46127);
xor U49135 (N_49135,N_46807,N_46279);
xnor U49136 (N_49136,N_47409,N_47301);
and U49137 (N_49137,N_47721,N_47144);
nand U49138 (N_49138,N_46200,N_47198);
xnor U49139 (N_49139,N_46814,N_46551);
and U49140 (N_49140,N_47410,N_46258);
nand U49141 (N_49141,N_47099,N_47255);
nand U49142 (N_49142,N_46635,N_47643);
or U49143 (N_49143,N_46990,N_47751);
xor U49144 (N_49144,N_47477,N_46460);
nor U49145 (N_49145,N_46657,N_46717);
xnor U49146 (N_49146,N_47607,N_47493);
nor U49147 (N_49147,N_47441,N_47195);
xor U49148 (N_49148,N_46163,N_47899);
xor U49149 (N_49149,N_47671,N_46443);
or U49150 (N_49150,N_47981,N_46630);
xor U49151 (N_49151,N_46933,N_46410);
xnor U49152 (N_49152,N_46126,N_47145);
nor U49153 (N_49153,N_46908,N_46877);
and U49154 (N_49154,N_46277,N_46915);
or U49155 (N_49155,N_46938,N_46444);
nor U49156 (N_49156,N_46971,N_47042);
nand U49157 (N_49157,N_46030,N_46435);
nor U49158 (N_49158,N_47004,N_46412);
or U49159 (N_49159,N_47987,N_47424);
xnor U49160 (N_49160,N_46915,N_46385);
nor U49161 (N_49161,N_47630,N_46755);
nor U49162 (N_49162,N_47126,N_46165);
nand U49163 (N_49163,N_47012,N_46511);
nor U49164 (N_49164,N_46163,N_46072);
and U49165 (N_49165,N_47860,N_47107);
nor U49166 (N_49166,N_47660,N_47891);
xor U49167 (N_49167,N_46820,N_46865);
nand U49168 (N_49168,N_47450,N_47937);
xor U49169 (N_49169,N_46117,N_46388);
and U49170 (N_49170,N_46718,N_47666);
or U49171 (N_49171,N_47409,N_46653);
xor U49172 (N_49172,N_47817,N_46498);
or U49173 (N_49173,N_47798,N_46010);
nand U49174 (N_49174,N_47889,N_46142);
xor U49175 (N_49175,N_46701,N_47872);
and U49176 (N_49176,N_47042,N_46142);
xnor U49177 (N_49177,N_46201,N_46261);
and U49178 (N_49178,N_47820,N_46818);
nor U49179 (N_49179,N_46709,N_46793);
and U49180 (N_49180,N_47629,N_46561);
xnor U49181 (N_49181,N_46637,N_47245);
nor U49182 (N_49182,N_46107,N_47725);
nand U49183 (N_49183,N_46497,N_46972);
or U49184 (N_49184,N_47374,N_46736);
or U49185 (N_49185,N_47850,N_47810);
xor U49186 (N_49186,N_47304,N_47975);
nor U49187 (N_49187,N_46561,N_47432);
and U49188 (N_49188,N_46096,N_47654);
nand U49189 (N_49189,N_46998,N_47880);
xor U49190 (N_49190,N_46799,N_47313);
nor U49191 (N_49191,N_46107,N_46998);
xnor U49192 (N_49192,N_47206,N_47428);
xnor U49193 (N_49193,N_46796,N_46750);
and U49194 (N_49194,N_47738,N_46690);
nor U49195 (N_49195,N_46121,N_46788);
and U49196 (N_49196,N_46619,N_47709);
xnor U49197 (N_49197,N_47044,N_46992);
and U49198 (N_49198,N_46819,N_46814);
nor U49199 (N_49199,N_46302,N_47137);
or U49200 (N_49200,N_47549,N_46756);
or U49201 (N_49201,N_47850,N_46149);
xor U49202 (N_49202,N_46138,N_47630);
and U49203 (N_49203,N_47396,N_47659);
nand U49204 (N_49204,N_46469,N_47372);
and U49205 (N_49205,N_46753,N_46189);
nand U49206 (N_49206,N_47534,N_47476);
or U49207 (N_49207,N_47673,N_46640);
and U49208 (N_49208,N_47758,N_47428);
and U49209 (N_49209,N_46681,N_46298);
and U49210 (N_49210,N_46250,N_47017);
xnor U49211 (N_49211,N_46216,N_46023);
xnor U49212 (N_49212,N_46957,N_47859);
xor U49213 (N_49213,N_47198,N_47026);
nand U49214 (N_49214,N_46486,N_47113);
nand U49215 (N_49215,N_47115,N_46971);
xnor U49216 (N_49216,N_46693,N_46490);
nand U49217 (N_49217,N_46870,N_47564);
xor U49218 (N_49218,N_46943,N_46895);
and U49219 (N_49219,N_47215,N_47013);
nand U49220 (N_49220,N_47389,N_47410);
or U49221 (N_49221,N_46411,N_47051);
and U49222 (N_49222,N_47759,N_47279);
and U49223 (N_49223,N_47847,N_47827);
and U49224 (N_49224,N_46659,N_47016);
nand U49225 (N_49225,N_47268,N_46103);
xnor U49226 (N_49226,N_46478,N_46924);
nor U49227 (N_49227,N_46011,N_47693);
nand U49228 (N_49228,N_47993,N_47458);
and U49229 (N_49229,N_46690,N_47818);
nor U49230 (N_49230,N_47925,N_46149);
or U49231 (N_49231,N_46130,N_47577);
or U49232 (N_49232,N_46073,N_47599);
nand U49233 (N_49233,N_47852,N_46400);
nor U49234 (N_49234,N_47519,N_47268);
xor U49235 (N_49235,N_46516,N_46570);
nand U49236 (N_49236,N_47349,N_46494);
or U49237 (N_49237,N_46257,N_46942);
nor U49238 (N_49238,N_47697,N_47230);
or U49239 (N_49239,N_46095,N_47022);
and U49240 (N_49240,N_46401,N_46622);
or U49241 (N_49241,N_46921,N_46722);
xor U49242 (N_49242,N_46277,N_47541);
xnor U49243 (N_49243,N_46142,N_46740);
nand U49244 (N_49244,N_47434,N_47432);
or U49245 (N_49245,N_47914,N_47946);
xor U49246 (N_49246,N_47212,N_47019);
xor U49247 (N_49247,N_46935,N_46520);
and U49248 (N_49248,N_46938,N_46108);
or U49249 (N_49249,N_46344,N_46165);
and U49250 (N_49250,N_46444,N_46607);
and U49251 (N_49251,N_46163,N_47766);
nor U49252 (N_49252,N_46219,N_47928);
or U49253 (N_49253,N_46468,N_47933);
xnor U49254 (N_49254,N_46910,N_47766);
or U49255 (N_49255,N_47496,N_47245);
and U49256 (N_49256,N_47532,N_46611);
and U49257 (N_49257,N_47643,N_46612);
nor U49258 (N_49258,N_46538,N_47769);
nand U49259 (N_49259,N_47010,N_47805);
and U49260 (N_49260,N_46472,N_47742);
xnor U49261 (N_49261,N_47893,N_47464);
or U49262 (N_49262,N_46171,N_46262);
nand U49263 (N_49263,N_46418,N_47436);
nor U49264 (N_49264,N_47621,N_47053);
nand U49265 (N_49265,N_47231,N_46036);
nand U49266 (N_49266,N_46499,N_47830);
or U49267 (N_49267,N_47608,N_47256);
xor U49268 (N_49268,N_47994,N_47433);
xor U49269 (N_49269,N_46931,N_46491);
xor U49270 (N_49270,N_46789,N_46657);
nand U49271 (N_49271,N_46520,N_46793);
and U49272 (N_49272,N_46388,N_47958);
or U49273 (N_49273,N_47864,N_47460);
and U49274 (N_49274,N_47835,N_47061);
nor U49275 (N_49275,N_47659,N_47119);
nand U49276 (N_49276,N_46877,N_47547);
nand U49277 (N_49277,N_47394,N_47504);
or U49278 (N_49278,N_46140,N_46815);
nand U49279 (N_49279,N_46750,N_46741);
nor U49280 (N_49280,N_47214,N_47094);
nor U49281 (N_49281,N_46250,N_46232);
or U49282 (N_49282,N_46136,N_46656);
nand U49283 (N_49283,N_47339,N_47948);
nor U49284 (N_49284,N_47168,N_47471);
nor U49285 (N_49285,N_47989,N_46422);
nor U49286 (N_49286,N_46079,N_46366);
and U49287 (N_49287,N_47137,N_47747);
xnor U49288 (N_49288,N_47648,N_46406);
and U49289 (N_49289,N_46545,N_46373);
xor U49290 (N_49290,N_46202,N_46595);
and U49291 (N_49291,N_46541,N_47668);
nor U49292 (N_49292,N_47771,N_46171);
nand U49293 (N_49293,N_47414,N_47544);
nor U49294 (N_49294,N_47780,N_46992);
xnor U49295 (N_49295,N_47887,N_47617);
nand U49296 (N_49296,N_46619,N_46961);
and U49297 (N_49297,N_47739,N_46757);
nand U49298 (N_49298,N_46407,N_46024);
nand U49299 (N_49299,N_46818,N_47496);
nor U49300 (N_49300,N_47198,N_46781);
or U49301 (N_49301,N_46864,N_47459);
nor U49302 (N_49302,N_47740,N_47498);
or U49303 (N_49303,N_47855,N_46756);
and U49304 (N_49304,N_47499,N_46227);
nor U49305 (N_49305,N_47473,N_47093);
nor U49306 (N_49306,N_46502,N_47127);
nor U49307 (N_49307,N_47057,N_46679);
and U49308 (N_49308,N_47652,N_47184);
nand U49309 (N_49309,N_46447,N_46609);
nor U49310 (N_49310,N_46919,N_46875);
or U49311 (N_49311,N_47076,N_46909);
and U49312 (N_49312,N_47860,N_47594);
or U49313 (N_49313,N_46499,N_46033);
or U49314 (N_49314,N_47803,N_47936);
or U49315 (N_49315,N_47849,N_46448);
xor U49316 (N_49316,N_47537,N_46600);
xor U49317 (N_49317,N_47996,N_46132);
xnor U49318 (N_49318,N_47742,N_47298);
or U49319 (N_49319,N_46260,N_47036);
and U49320 (N_49320,N_47083,N_47312);
or U49321 (N_49321,N_47479,N_47730);
and U49322 (N_49322,N_46785,N_47826);
nor U49323 (N_49323,N_46285,N_46198);
nand U49324 (N_49324,N_46951,N_47975);
nor U49325 (N_49325,N_46038,N_46934);
and U49326 (N_49326,N_47798,N_47160);
or U49327 (N_49327,N_47574,N_46950);
and U49328 (N_49328,N_46592,N_47670);
nand U49329 (N_49329,N_46494,N_46686);
or U49330 (N_49330,N_46358,N_46979);
xor U49331 (N_49331,N_46690,N_46208);
xor U49332 (N_49332,N_47548,N_47904);
or U49333 (N_49333,N_47006,N_47164);
and U49334 (N_49334,N_46889,N_47465);
nand U49335 (N_49335,N_46653,N_46487);
nand U49336 (N_49336,N_46893,N_47560);
or U49337 (N_49337,N_47110,N_47251);
nor U49338 (N_49338,N_46036,N_47124);
nand U49339 (N_49339,N_46361,N_47972);
or U49340 (N_49340,N_47118,N_46812);
xnor U49341 (N_49341,N_46088,N_47685);
xnor U49342 (N_49342,N_46755,N_47882);
nor U49343 (N_49343,N_46056,N_46614);
nand U49344 (N_49344,N_46712,N_47280);
or U49345 (N_49345,N_46748,N_46598);
nor U49346 (N_49346,N_47960,N_46215);
and U49347 (N_49347,N_46495,N_47121);
nand U49348 (N_49348,N_46024,N_46085);
or U49349 (N_49349,N_47426,N_46548);
nand U49350 (N_49350,N_47848,N_47659);
and U49351 (N_49351,N_47076,N_47317);
xor U49352 (N_49352,N_46438,N_46238);
or U49353 (N_49353,N_47256,N_46004);
or U49354 (N_49354,N_47489,N_47486);
and U49355 (N_49355,N_47334,N_47602);
xor U49356 (N_49356,N_46010,N_46717);
or U49357 (N_49357,N_46813,N_46243);
xor U49358 (N_49358,N_46733,N_46423);
and U49359 (N_49359,N_47778,N_46098);
nand U49360 (N_49360,N_46314,N_46252);
nor U49361 (N_49361,N_46316,N_47558);
nor U49362 (N_49362,N_47393,N_47773);
or U49363 (N_49363,N_46611,N_47453);
and U49364 (N_49364,N_47814,N_46373);
nor U49365 (N_49365,N_47086,N_46502);
and U49366 (N_49366,N_46999,N_46651);
nand U49367 (N_49367,N_47869,N_46079);
nor U49368 (N_49368,N_46330,N_46273);
or U49369 (N_49369,N_46410,N_47703);
nand U49370 (N_49370,N_47129,N_46616);
or U49371 (N_49371,N_47080,N_47663);
and U49372 (N_49372,N_46679,N_47259);
nor U49373 (N_49373,N_47135,N_46403);
xnor U49374 (N_49374,N_46893,N_46171);
xor U49375 (N_49375,N_47373,N_47779);
and U49376 (N_49376,N_47803,N_46747);
xnor U49377 (N_49377,N_46195,N_46499);
or U49378 (N_49378,N_47681,N_47426);
and U49379 (N_49379,N_46825,N_47485);
xor U49380 (N_49380,N_47020,N_46865);
nor U49381 (N_49381,N_47669,N_46446);
and U49382 (N_49382,N_47050,N_46575);
nor U49383 (N_49383,N_46820,N_47156);
xor U49384 (N_49384,N_47816,N_46091);
and U49385 (N_49385,N_46300,N_46845);
xnor U49386 (N_49386,N_47279,N_47129);
xor U49387 (N_49387,N_46418,N_47241);
nor U49388 (N_49388,N_46940,N_46035);
or U49389 (N_49389,N_47698,N_47674);
nand U49390 (N_49390,N_47809,N_47458);
and U49391 (N_49391,N_47530,N_46694);
xor U49392 (N_49392,N_46205,N_46262);
nand U49393 (N_49393,N_47084,N_47093);
nand U49394 (N_49394,N_47575,N_47836);
nor U49395 (N_49395,N_46300,N_46667);
or U49396 (N_49396,N_47705,N_47424);
nor U49397 (N_49397,N_47675,N_47613);
nor U49398 (N_49398,N_47226,N_46267);
and U49399 (N_49399,N_47689,N_47001);
and U49400 (N_49400,N_46167,N_46160);
and U49401 (N_49401,N_46639,N_46220);
nor U49402 (N_49402,N_46538,N_46634);
nor U49403 (N_49403,N_47155,N_47144);
nand U49404 (N_49404,N_46546,N_47044);
xnor U49405 (N_49405,N_47575,N_46429);
and U49406 (N_49406,N_47171,N_46350);
xnor U49407 (N_49407,N_47612,N_46723);
and U49408 (N_49408,N_46197,N_47697);
or U49409 (N_49409,N_47772,N_47763);
nor U49410 (N_49410,N_47590,N_47513);
and U49411 (N_49411,N_46272,N_46018);
and U49412 (N_49412,N_47964,N_46995);
nand U49413 (N_49413,N_47845,N_47984);
nor U49414 (N_49414,N_46782,N_46201);
or U49415 (N_49415,N_46430,N_46445);
and U49416 (N_49416,N_46222,N_46611);
or U49417 (N_49417,N_47710,N_46632);
nor U49418 (N_49418,N_46844,N_47932);
nor U49419 (N_49419,N_46838,N_47327);
nand U49420 (N_49420,N_46683,N_47660);
xnor U49421 (N_49421,N_47676,N_47705);
nor U49422 (N_49422,N_47223,N_46961);
nand U49423 (N_49423,N_46520,N_47342);
or U49424 (N_49424,N_46671,N_46709);
and U49425 (N_49425,N_47546,N_47138);
or U49426 (N_49426,N_46158,N_46822);
xnor U49427 (N_49427,N_46801,N_46018);
and U49428 (N_49428,N_46591,N_47526);
nand U49429 (N_49429,N_46243,N_46982);
xnor U49430 (N_49430,N_47275,N_47965);
and U49431 (N_49431,N_47842,N_47583);
xnor U49432 (N_49432,N_47146,N_46735);
or U49433 (N_49433,N_47282,N_46422);
nor U49434 (N_49434,N_47967,N_47986);
nand U49435 (N_49435,N_47969,N_47361);
nand U49436 (N_49436,N_47647,N_46275);
and U49437 (N_49437,N_47630,N_47758);
xor U49438 (N_49438,N_47777,N_47369);
nor U49439 (N_49439,N_46360,N_47411);
nor U49440 (N_49440,N_47741,N_47746);
nor U49441 (N_49441,N_47430,N_47566);
or U49442 (N_49442,N_47624,N_46739);
nor U49443 (N_49443,N_47890,N_47299);
nor U49444 (N_49444,N_46809,N_47766);
xnor U49445 (N_49445,N_47057,N_47412);
or U49446 (N_49446,N_46887,N_46498);
or U49447 (N_49447,N_47771,N_47274);
nand U49448 (N_49448,N_46840,N_46725);
nor U49449 (N_49449,N_46999,N_46706);
xor U49450 (N_49450,N_46917,N_46846);
nand U49451 (N_49451,N_47281,N_47212);
xor U49452 (N_49452,N_46821,N_47675);
and U49453 (N_49453,N_46097,N_46857);
and U49454 (N_49454,N_46182,N_46523);
nor U49455 (N_49455,N_46698,N_46525);
xor U49456 (N_49456,N_47959,N_46517);
nor U49457 (N_49457,N_46803,N_46658);
xnor U49458 (N_49458,N_47448,N_46545);
nand U49459 (N_49459,N_46489,N_46689);
nand U49460 (N_49460,N_47944,N_47408);
or U49461 (N_49461,N_46969,N_47643);
xnor U49462 (N_49462,N_47177,N_46883);
xnor U49463 (N_49463,N_46985,N_46143);
nor U49464 (N_49464,N_47313,N_46085);
and U49465 (N_49465,N_46902,N_46208);
nor U49466 (N_49466,N_47604,N_46920);
xnor U49467 (N_49467,N_46021,N_46657);
xor U49468 (N_49468,N_47751,N_46078);
and U49469 (N_49469,N_46622,N_47547);
nand U49470 (N_49470,N_47461,N_47626);
and U49471 (N_49471,N_46394,N_47648);
nor U49472 (N_49472,N_46519,N_46441);
and U49473 (N_49473,N_47223,N_46729);
nor U49474 (N_49474,N_46227,N_46453);
xnor U49475 (N_49475,N_46173,N_46231);
or U49476 (N_49476,N_47253,N_46379);
nand U49477 (N_49477,N_46676,N_46220);
xor U49478 (N_49478,N_47161,N_46388);
nand U49479 (N_49479,N_46387,N_46753);
nand U49480 (N_49480,N_47538,N_46071);
nand U49481 (N_49481,N_46959,N_47453);
and U49482 (N_49482,N_46886,N_47027);
or U49483 (N_49483,N_46680,N_47910);
xor U49484 (N_49484,N_46773,N_46035);
xnor U49485 (N_49485,N_47801,N_47952);
or U49486 (N_49486,N_46665,N_47064);
nand U49487 (N_49487,N_46729,N_47688);
and U49488 (N_49488,N_46917,N_46857);
and U49489 (N_49489,N_46440,N_46922);
nor U49490 (N_49490,N_47656,N_46700);
nand U49491 (N_49491,N_47568,N_47316);
and U49492 (N_49492,N_46523,N_46519);
nor U49493 (N_49493,N_46073,N_46178);
nand U49494 (N_49494,N_46451,N_47408);
nand U49495 (N_49495,N_46029,N_47127);
nor U49496 (N_49496,N_46185,N_46788);
xor U49497 (N_49497,N_46327,N_47237);
xnor U49498 (N_49498,N_47083,N_47762);
and U49499 (N_49499,N_46267,N_46867);
nand U49500 (N_49500,N_46853,N_46211);
nor U49501 (N_49501,N_46147,N_46306);
or U49502 (N_49502,N_47454,N_47440);
or U49503 (N_49503,N_47968,N_46675);
xor U49504 (N_49504,N_46998,N_46318);
or U49505 (N_49505,N_47845,N_46329);
nand U49506 (N_49506,N_46314,N_47347);
xor U49507 (N_49507,N_47054,N_46421);
and U49508 (N_49508,N_46101,N_47375);
nor U49509 (N_49509,N_47227,N_46454);
and U49510 (N_49510,N_47419,N_47046);
nor U49511 (N_49511,N_46947,N_47506);
or U49512 (N_49512,N_46676,N_46096);
and U49513 (N_49513,N_46452,N_46704);
nor U49514 (N_49514,N_46356,N_46104);
xor U49515 (N_49515,N_47714,N_47328);
and U49516 (N_49516,N_46595,N_46382);
nor U49517 (N_49517,N_46537,N_46862);
and U49518 (N_49518,N_46244,N_46490);
or U49519 (N_49519,N_46013,N_47214);
or U49520 (N_49520,N_46597,N_46688);
xor U49521 (N_49521,N_46427,N_46421);
xor U49522 (N_49522,N_46117,N_47621);
nand U49523 (N_49523,N_47394,N_47359);
nor U49524 (N_49524,N_46558,N_46417);
or U49525 (N_49525,N_46382,N_47910);
or U49526 (N_49526,N_46011,N_46569);
nand U49527 (N_49527,N_46702,N_46988);
xnor U49528 (N_49528,N_46520,N_47940);
or U49529 (N_49529,N_46516,N_47073);
xnor U49530 (N_49530,N_47548,N_47461);
xnor U49531 (N_49531,N_46999,N_47036);
nand U49532 (N_49532,N_47039,N_46213);
nand U49533 (N_49533,N_47029,N_47555);
nor U49534 (N_49534,N_47066,N_47912);
nand U49535 (N_49535,N_46602,N_46944);
nand U49536 (N_49536,N_46403,N_47230);
and U49537 (N_49537,N_47473,N_47618);
nor U49538 (N_49538,N_46601,N_47538);
and U49539 (N_49539,N_46319,N_46304);
or U49540 (N_49540,N_46402,N_46424);
or U49541 (N_49541,N_47940,N_47897);
and U49542 (N_49542,N_47104,N_47039);
nor U49543 (N_49543,N_46090,N_46556);
and U49544 (N_49544,N_47247,N_46117);
nor U49545 (N_49545,N_47611,N_47484);
nand U49546 (N_49546,N_46865,N_46387);
nor U49547 (N_49547,N_47462,N_47285);
xor U49548 (N_49548,N_47709,N_47048);
and U49549 (N_49549,N_47416,N_47643);
nand U49550 (N_49550,N_47371,N_47479);
xor U49551 (N_49551,N_46889,N_46963);
and U49552 (N_49552,N_47358,N_47013);
nor U49553 (N_49553,N_47688,N_47340);
nand U49554 (N_49554,N_47191,N_47257);
xnor U49555 (N_49555,N_46197,N_47994);
nand U49556 (N_49556,N_46424,N_47305);
xnor U49557 (N_49557,N_46531,N_47691);
nor U49558 (N_49558,N_46770,N_47249);
nor U49559 (N_49559,N_47311,N_47255);
xnor U49560 (N_49560,N_46487,N_46320);
or U49561 (N_49561,N_46767,N_46998);
and U49562 (N_49562,N_46304,N_46977);
nor U49563 (N_49563,N_47876,N_46243);
xor U49564 (N_49564,N_47664,N_46127);
nand U49565 (N_49565,N_46825,N_47180);
nand U49566 (N_49566,N_46370,N_47563);
nand U49567 (N_49567,N_46685,N_47049);
nor U49568 (N_49568,N_46025,N_47030);
and U49569 (N_49569,N_47988,N_47315);
xnor U49570 (N_49570,N_47939,N_46973);
nor U49571 (N_49571,N_46222,N_46740);
xnor U49572 (N_49572,N_46598,N_47187);
nor U49573 (N_49573,N_47670,N_47953);
nor U49574 (N_49574,N_46316,N_47341);
xor U49575 (N_49575,N_47318,N_47180);
or U49576 (N_49576,N_47762,N_46548);
or U49577 (N_49577,N_46578,N_47311);
nor U49578 (N_49578,N_47478,N_47326);
xor U49579 (N_49579,N_46105,N_47103);
nand U49580 (N_49580,N_46193,N_47242);
and U49581 (N_49581,N_47326,N_46835);
nand U49582 (N_49582,N_46392,N_46688);
nand U49583 (N_49583,N_46298,N_46557);
and U49584 (N_49584,N_46287,N_46599);
xor U49585 (N_49585,N_47447,N_47421);
or U49586 (N_49586,N_47650,N_46504);
xor U49587 (N_49587,N_46170,N_47096);
and U49588 (N_49588,N_47294,N_47408);
or U49589 (N_49589,N_47977,N_47382);
or U49590 (N_49590,N_46416,N_46439);
nand U49591 (N_49591,N_46676,N_47453);
xnor U49592 (N_49592,N_47235,N_47440);
or U49593 (N_49593,N_47061,N_46926);
xnor U49594 (N_49594,N_47761,N_47166);
xnor U49595 (N_49595,N_47261,N_47545);
or U49596 (N_49596,N_46363,N_47522);
nor U49597 (N_49597,N_47069,N_46622);
or U49598 (N_49598,N_46925,N_46427);
and U49599 (N_49599,N_46025,N_47602);
nand U49600 (N_49600,N_47415,N_46378);
or U49601 (N_49601,N_46996,N_47077);
and U49602 (N_49602,N_47137,N_46668);
xnor U49603 (N_49603,N_46740,N_46989);
and U49604 (N_49604,N_46863,N_47422);
and U49605 (N_49605,N_46940,N_46621);
and U49606 (N_49606,N_47656,N_47682);
xnor U49607 (N_49607,N_46026,N_47895);
and U49608 (N_49608,N_47313,N_47594);
nor U49609 (N_49609,N_47066,N_46016);
or U49610 (N_49610,N_47449,N_46249);
nor U49611 (N_49611,N_46952,N_46714);
and U49612 (N_49612,N_46368,N_47893);
nor U49613 (N_49613,N_47658,N_47037);
or U49614 (N_49614,N_46847,N_46375);
xnor U49615 (N_49615,N_47349,N_46557);
nand U49616 (N_49616,N_46859,N_46348);
or U49617 (N_49617,N_46084,N_46888);
nand U49618 (N_49618,N_46832,N_46447);
and U49619 (N_49619,N_47937,N_47336);
and U49620 (N_49620,N_46574,N_47491);
nor U49621 (N_49621,N_47196,N_47520);
xor U49622 (N_49622,N_46384,N_47060);
nor U49623 (N_49623,N_47635,N_47480);
nor U49624 (N_49624,N_47066,N_47434);
nor U49625 (N_49625,N_46338,N_46681);
xnor U49626 (N_49626,N_46428,N_47015);
xor U49627 (N_49627,N_46306,N_47421);
xnor U49628 (N_49628,N_46336,N_46775);
nand U49629 (N_49629,N_46780,N_47536);
xnor U49630 (N_49630,N_47830,N_47980);
or U49631 (N_49631,N_47463,N_47166);
nor U49632 (N_49632,N_46713,N_46389);
xnor U49633 (N_49633,N_46289,N_47370);
xnor U49634 (N_49634,N_46247,N_46619);
nand U49635 (N_49635,N_47312,N_47813);
nor U49636 (N_49636,N_47293,N_47933);
or U49637 (N_49637,N_46612,N_46873);
or U49638 (N_49638,N_46711,N_46230);
xnor U49639 (N_49639,N_47118,N_47031);
nand U49640 (N_49640,N_46105,N_46666);
and U49641 (N_49641,N_46012,N_46134);
or U49642 (N_49642,N_46281,N_46950);
nor U49643 (N_49643,N_46848,N_46544);
nand U49644 (N_49644,N_47712,N_46333);
and U49645 (N_49645,N_47010,N_47183);
nor U49646 (N_49646,N_46456,N_46305);
and U49647 (N_49647,N_46861,N_47800);
nor U49648 (N_49648,N_46168,N_46802);
xor U49649 (N_49649,N_47683,N_46476);
nand U49650 (N_49650,N_47808,N_47490);
nand U49651 (N_49651,N_47948,N_46099);
xor U49652 (N_49652,N_47072,N_46947);
nor U49653 (N_49653,N_47798,N_46781);
nor U49654 (N_49654,N_47643,N_47180);
nand U49655 (N_49655,N_46187,N_47677);
or U49656 (N_49656,N_47613,N_47990);
and U49657 (N_49657,N_47997,N_46171);
nor U49658 (N_49658,N_47861,N_47653);
and U49659 (N_49659,N_46831,N_46841);
nand U49660 (N_49660,N_47339,N_47160);
and U49661 (N_49661,N_47939,N_46785);
and U49662 (N_49662,N_46438,N_47383);
nor U49663 (N_49663,N_46192,N_47983);
xor U49664 (N_49664,N_47510,N_46505);
xor U49665 (N_49665,N_46750,N_46545);
and U49666 (N_49666,N_46172,N_46055);
nor U49667 (N_49667,N_46362,N_46216);
xnor U49668 (N_49668,N_47300,N_47866);
xnor U49669 (N_49669,N_46751,N_47683);
xor U49670 (N_49670,N_47905,N_47164);
or U49671 (N_49671,N_46118,N_46810);
xor U49672 (N_49672,N_46506,N_47195);
xor U49673 (N_49673,N_46545,N_46669);
nor U49674 (N_49674,N_47386,N_47900);
nand U49675 (N_49675,N_46288,N_46187);
or U49676 (N_49676,N_47149,N_46130);
xor U49677 (N_49677,N_47504,N_46228);
xnor U49678 (N_49678,N_47020,N_46815);
and U49679 (N_49679,N_47734,N_46851);
and U49680 (N_49680,N_47207,N_46709);
and U49681 (N_49681,N_47122,N_47078);
and U49682 (N_49682,N_46897,N_47195);
and U49683 (N_49683,N_47935,N_47369);
xor U49684 (N_49684,N_46799,N_46771);
xor U49685 (N_49685,N_47725,N_47931);
and U49686 (N_49686,N_46395,N_46575);
xor U49687 (N_49687,N_46468,N_46969);
nand U49688 (N_49688,N_46017,N_47835);
nand U49689 (N_49689,N_47390,N_46150);
xnor U49690 (N_49690,N_47835,N_47202);
or U49691 (N_49691,N_47001,N_46441);
xnor U49692 (N_49692,N_46421,N_47332);
nand U49693 (N_49693,N_47442,N_47506);
and U49694 (N_49694,N_46339,N_47191);
nand U49695 (N_49695,N_46559,N_46544);
or U49696 (N_49696,N_47158,N_47756);
and U49697 (N_49697,N_46023,N_46172);
and U49698 (N_49698,N_46505,N_46235);
or U49699 (N_49699,N_47227,N_46540);
nand U49700 (N_49700,N_47815,N_46553);
or U49701 (N_49701,N_46179,N_46432);
nand U49702 (N_49702,N_47496,N_47998);
nor U49703 (N_49703,N_46618,N_47748);
or U49704 (N_49704,N_46725,N_47646);
xor U49705 (N_49705,N_47529,N_46801);
xnor U49706 (N_49706,N_46720,N_47203);
or U49707 (N_49707,N_46917,N_47554);
xnor U49708 (N_49708,N_46489,N_46620);
or U49709 (N_49709,N_46825,N_46217);
nor U49710 (N_49710,N_47112,N_46083);
nor U49711 (N_49711,N_47198,N_46535);
xor U49712 (N_49712,N_47116,N_47644);
nand U49713 (N_49713,N_46577,N_46159);
and U49714 (N_49714,N_46525,N_46350);
or U49715 (N_49715,N_47082,N_46467);
nand U49716 (N_49716,N_47814,N_47816);
or U49717 (N_49717,N_46233,N_46791);
nor U49718 (N_49718,N_46218,N_46835);
xor U49719 (N_49719,N_46727,N_47966);
nor U49720 (N_49720,N_46590,N_46022);
or U49721 (N_49721,N_46858,N_46255);
nor U49722 (N_49722,N_47846,N_46951);
and U49723 (N_49723,N_46428,N_47849);
nor U49724 (N_49724,N_47358,N_46135);
or U49725 (N_49725,N_46042,N_46128);
xnor U49726 (N_49726,N_47973,N_47227);
nand U49727 (N_49727,N_46780,N_46737);
nor U49728 (N_49728,N_46026,N_46730);
or U49729 (N_49729,N_47569,N_47654);
and U49730 (N_49730,N_47151,N_47050);
nand U49731 (N_49731,N_47469,N_47417);
and U49732 (N_49732,N_47073,N_47588);
and U49733 (N_49733,N_47442,N_47504);
nand U49734 (N_49734,N_47079,N_46884);
or U49735 (N_49735,N_47309,N_47675);
nand U49736 (N_49736,N_47315,N_46789);
and U49737 (N_49737,N_47835,N_47988);
nand U49738 (N_49738,N_47496,N_46170);
and U49739 (N_49739,N_47267,N_46316);
xnor U49740 (N_49740,N_47531,N_46357);
nand U49741 (N_49741,N_46095,N_46649);
or U49742 (N_49742,N_46937,N_47241);
nor U49743 (N_49743,N_46741,N_46024);
and U49744 (N_49744,N_47781,N_47834);
nor U49745 (N_49745,N_46341,N_46159);
and U49746 (N_49746,N_47415,N_47782);
or U49747 (N_49747,N_46611,N_46690);
nor U49748 (N_49748,N_47588,N_47179);
xor U49749 (N_49749,N_47902,N_46896);
or U49750 (N_49750,N_47049,N_47210);
nand U49751 (N_49751,N_46010,N_47825);
xor U49752 (N_49752,N_46850,N_47330);
nand U49753 (N_49753,N_46616,N_46808);
nand U49754 (N_49754,N_47454,N_46748);
and U49755 (N_49755,N_47888,N_46789);
and U49756 (N_49756,N_46430,N_47619);
xor U49757 (N_49757,N_47602,N_47790);
nand U49758 (N_49758,N_46923,N_46676);
nand U49759 (N_49759,N_47035,N_47083);
nand U49760 (N_49760,N_46789,N_46729);
xnor U49761 (N_49761,N_47993,N_46348);
nor U49762 (N_49762,N_46282,N_46735);
or U49763 (N_49763,N_46870,N_46194);
xnor U49764 (N_49764,N_46256,N_47378);
xor U49765 (N_49765,N_47029,N_46364);
or U49766 (N_49766,N_46367,N_46243);
xnor U49767 (N_49767,N_47567,N_46819);
or U49768 (N_49768,N_46008,N_47577);
and U49769 (N_49769,N_46354,N_47970);
nand U49770 (N_49770,N_46867,N_46269);
or U49771 (N_49771,N_47431,N_47552);
nor U49772 (N_49772,N_46826,N_47446);
nand U49773 (N_49773,N_46017,N_46085);
nand U49774 (N_49774,N_46538,N_47739);
nor U49775 (N_49775,N_46569,N_46767);
nor U49776 (N_49776,N_47688,N_46328);
xnor U49777 (N_49777,N_47400,N_47030);
and U49778 (N_49778,N_47422,N_47774);
xor U49779 (N_49779,N_47241,N_46864);
and U49780 (N_49780,N_46654,N_46338);
nor U49781 (N_49781,N_46017,N_46707);
xnor U49782 (N_49782,N_47461,N_47534);
nor U49783 (N_49783,N_47317,N_46756);
nor U49784 (N_49784,N_47978,N_47339);
and U49785 (N_49785,N_47862,N_47823);
nor U49786 (N_49786,N_47915,N_46089);
nor U49787 (N_49787,N_46123,N_47111);
xnor U49788 (N_49788,N_47808,N_47238);
nor U49789 (N_49789,N_46899,N_47781);
or U49790 (N_49790,N_46864,N_47541);
nand U49791 (N_49791,N_47622,N_46557);
xnor U49792 (N_49792,N_47902,N_46561);
and U49793 (N_49793,N_46004,N_46136);
xor U49794 (N_49794,N_46861,N_46077);
and U49795 (N_49795,N_47169,N_47552);
xor U49796 (N_49796,N_47744,N_46697);
xor U49797 (N_49797,N_46238,N_47864);
and U49798 (N_49798,N_47833,N_47703);
nand U49799 (N_49799,N_46266,N_47139);
and U49800 (N_49800,N_46559,N_46680);
xnor U49801 (N_49801,N_47409,N_47926);
or U49802 (N_49802,N_47740,N_46226);
xnor U49803 (N_49803,N_47275,N_46507);
or U49804 (N_49804,N_47944,N_47892);
nand U49805 (N_49805,N_47789,N_47772);
xnor U49806 (N_49806,N_46253,N_47975);
nor U49807 (N_49807,N_47454,N_47617);
xnor U49808 (N_49808,N_46349,N_47530);
or U49809 (N_49809,N_46229,N_47137);
xor U49810 (N_49810,N_47267,N_46930);
or U49811 (N_49811,N_47227,N_47928);
xnor U49812 (N_49812,N_46709,N_47912);
or U49813 (N_49813,N_47985,N_46395);
or U49814 (N_49814,N_46227,N_46725);
nor U49815 (N_49815,N_47296,N_47308);
nand U49816 (N_49816,N_47322,N_47500);
or U49817 (N_49817,N_47948,N_46887);
nor U49818 (N_49818,N_47669,N_47670);
xnor U49819 (N_49819,N_46134,N_46488);
and U49820 (N_49820,N_47950,N_47218);
nand U49821 (N_49821,N_47571,N_46689);
xnor U49822 (N_49822,N_47181,N_46887);
and U49823 (N_49823,N_47126,N_47865);
and U49824 (N_49824,N_47351,N_46480);
or U49825 (N_49825,N_47873,N_47791);
xnor U49826 (N_49826,N_46445,N_46403);
xnor U49827 (N_49827,N_46964,N_47585);
nor U49828 (N_49828,N_46183,N_47979);
and U49829 (N_49829,N_47207,N_47740);
nor U49830 (N_49830,N_46767,N_46070);
nand U49831 (N_49831,N_46658,N_46009);
nand U49832 (N_49832,N_47297,N_46364);
xnor U49833 (N_49833,N_47134,N_46253);
nand U49834 (N_49834,N_46678,N_46651);
nand U49835 (N_49835,N_47462,N_47620);
nand U49836 (N_49836,N_47564,N_47820);
xnor U49837 (N_49837,N_46761,N_46301);
or U49838 (N_49838,N_47961,N_47566);
nor U49839 (N_49839,N_47043,N_46232);
or U49840 (N_49840,N_47510,N_47614);
nor U49841 (N_49841,N_47755,N_46994);
or U49842 (N_49842,N_47285,N_47092);
and U49843 (N_49843,N_47837,N_46099);
or U49844 (N_49844,N_47605,N_46579);
or U49845 (N_49845,N_46066,N_47455);
nor U49846 (N_49846,N_47001,N_46960);
xnor U49847 (N_49847,N_46620,N_46377);
or U49848 (N_49848,N_46446,N_47807);
nor U49849 (N_49849,N_47455,N_47188);
nand U49850 (N_49850,N_46230,N_46354);
nand U49851 (N_49851,N_46081,N_47752);
or U49852 (N_49852,N_47398,N_46321);
or U49853 (N_49853,N_46817,N_47294);
nand U49854 (N_49854,N_46510,N_46002);
xor U49855 (N_49855,N_46630,N_47501);
xnor U49856 (N_49856,N_46394,N_47515);
or U49857 (N_49857,N_46321,N_47342);
xor U49858 (N_49858,N_46730,N_46851);
nand U49859 (N_49859,N_46298,N_47262);
nor U49860 (N_49860,N_46129,N_46839);
or U49861 (N_49861,N_47517,N_47947);
nand U49862 (N_49862,N_46813,N_46084);
and U49863 (N_49863,N_47593,N_46680);
nor U49864 (N_49864,N_47095,N_47292);
nand U49865 (N_49865,N_46749,N_46804);
xnor U49866 (N_49866,N_46842,N_46392);
or U49867 (N_49867,N_47058,N_47975);
and U49868 (N_49868,N_47993,N_47044);
or U49869 (N_49869,N_46327,N_46376);
or U49870 (N_49870,N_47027,N_46911);
nand U49871 (N_49871,N_47011,N_47168);
nand U49872 (N_49872,N_46738,N_46398);
xor U49873 (N_49873,N_47921,N_47954);
nand U49874 (N_49874,N_47734,N_46753);
and U49875 (N_49875,N_47926,N_47418);
nand U49876 (N_49876,N_46490,N_47866);
nor U49877 (N_49877,N_47071,N_47587);
and U49878 (N_49878,N_47532,N_47357);
nand U49879 (N_49879,N_47424,N_46453);
nand U49880 (N_49880,N_47580,N_46464);
and U49881 (N_49881,N_47600,N_47450);
xor U49882 (N_49882,N_46583,N_46785);
or U49883 (N_49883,N_47312,N_46104);
nor U49884 (N_49884,N_47420,N_47060);
or U49885 (N_49885,N_46916,N_47433);
and U49886 (N_49886,N_46787,N_47526);
or U49887 (N_49887,N_46816,N_46612);
nand U49888 (N_49888,N_47145,N_47202);
nand U49889 (N_49889,N_47179,N_46906);
nor U49890 (N_49890,N_46895,N_46207);
nor U49891 (N_49891,N_46846,N_47386);
or U49892 (N_49892,N_47028,N_47829);
or U49893 (N_49893,N_47961,N_46433);
or U49894 (N_49894,N_47685,N_47338);
xor U49895 (N_49895,N_47966,N_47251);
nor U49896 (N_49896,N_47945,N_46087);
or U49897 (N_49897,N_47445,N_47011);
nor U49898 (N_49898,N_47739,N_46213);
nor U49899 (N_49899,N_47336,N_47303);
or U49900 (N_49900,N_46564,N_46428);
nand U49901 (N_49901,N_46548,N_47422);
nand U49902 (N_49902,N_47858,N_47859);
xor U49903 (N_49903,N_46146,N_46682);
or U49904 (N_49904,N_47808,N_47722);
nor U49905 (N_49905,N_47080,N_47266);
or U49906 (N_49906,N_47133,N_46414);
nand U49907 (N_49907,N_47353,N_46089);
and U49908 (N_49908,N_47061,N_47244);
and U49909 (N_49909,N_46321,N_46010);
xor U49910 (N_49910,N_47357,N_46200);
nor U49911 (N_49911,N_47457,N_46815);
xor U49912 (N_49912,N_47309,N_47671);
and U49913 (N_49913,N_47459,N_46855);
and U49914 (N_49914,N_46582,N_47454);
nor U49915 (N_49915,N_47831,N_46488);
nor U49916 (N_49916,N_46301,N_47245);
or U49917 (N_49917,N_47291,N_47873);
nand U49918 (N_49918,N_46413,N_47929);
xnor U49919 (N_49919,N_46716,N_47508);
nor U49920 (N_49920,N_47463,N_46994);
and U49921 (N_49921,N_46071,N_46836);
xnor U49922 (N_49922,N_47201,N_46634);
or U49923 (N_49923,N_46113,N_47805);
nand U49924 (N_49924,N_47593,N_46663);
and U49925 (N_49925,N_46444,N_47197);
nand U49926 (N_49926,N_47227,N_46857);
nand U49927 (N_49927,N_46721,N_46354);
xnor U49928 (N_49928,N_47834,N_46540);
nor U49929 (N_49929,N_47550,N_46181);
and U49930 (N_49930,N_46391,N_46589);
or U49931 (N_49931,N_46389,N_47153);
nand U49932 (N_49932,N_47313,N_46275);
and U49933 (N_49933,N_46599,N_47537);
or U49934 (N_49934,N_47925,N_46021);
nand U49935 (N_49935,N_47269,N_46475);
nor U49936 (N_49936,N_47032,N_47822);
and U49937 (N_49937,N_47335,N_46006);
and U49938 (N_49938,N_46329,N_47783);
xnor U49939 (N_49939,N_47586,N_47990);
xor U49940 (N_49940,N_47842,N_46279);
xnor U49941 (N_49941,N_46846,N_46451);
xor U49942 (N_49942,N_47614,N_47681);
nand U49943 (N_49943,N_46797,N_47275);
or U49944 (N_49944,N_47886,N_47836);
nor U49945 (N_49945,N_46930,N_46921);
and U49946 (N_49946,N_46992,N_46173);
nand U49947 (N_49947,N_47768,N_46811);
xnor U49948 (N_49948,N_47227,N_46104);
nand U49949 (N_49949,N_47293,N_46836);
nand U49950 (N_49950,N_46351,N_47505);
and U49951 (N_49951,N_46129,N_47221);
or U49952 (N_49952,N_47801,N_47614);
nand U49953 (N_49953,N_47495,N_46459);
xnor U49954 (N_49954,N_47329,N_47396);
and U49955 (N_49955,N_47346,N_46105);
or U49956 (N_49956,N_46101,N_47577);
nand U49957 (N_49957,N_46949,N_47070);
xnor U49958 (N_49958,N_46704,N_47602);
and U49959 (N_49959,N_46274,N_47576);
xor U49960 (N_49960,N_47371,N_46202);
and U49961 (N_49961,N_47102,N_47865);
or U49962 (N_49962,N_46932,N_46768);
xnor U49963 (N_49963,N_46846,N_47615);
nor U49964 (N_49964,N_47892,N_47671);
or U49965 (N_49965,N_47019,N_46455);
xnor U49966 (N_49966,N_47272,N_47869);
xnor U49967 (N_49967,N_47073,N_46598);
xor U49968 (N_49968,N_47567,N_47239);
xnor U49969 (N_49969,N_47886,N_46631);
xnor U49970 (N_49970,N_47133,N_46933);
nand U49971 (N_49971,N_46148,N_47833);
nand U49972 (N_49972,N_46492,N_47490);
or U49973 (N_49973,N_47034,N_47255);
xor U49974 (N_49974,N_47165,N_46527);
nor U49975 (N_49975,N_47773,N_47554);
nand U49976 (N_49976,N_46748,N_47602);
or U49977 (N_49977,N_46138,N_47956);
xnor U49978 (N_49978,N_47380,N_46260);
xor U49979 (N_49979,N_46061,N_47943);
and U49980 (N_49980,N_47761,N_47811);
and U49981 (N_49981,N_47115,N_47877);
xor U49982 (N_49982,N_47747,N_46427);
nand U49983 (N_49983,N_47579,N_46201);
and U49984 (N_49984,N_47628,N_46072);
nand U49985 (N_49985,N_47729,N_46537);
xor U49986 (N_49986,N_46759,N_46505);
nor U49987 (N_49987,N_47618,N_46142);
nand U49988 (N_49988,N_47714,N_47230);
nand U49989 (N_49989,N_46888,N_46367);
xnor U49990 (N_49990,N_46809,N_46475);
xnor U49991 (N_49991,N_46916,N_46019);
or U49992 (N_49992,N_47957,N_47530);
nand U49993 (N_49993,N_47196,N_47665);
and U49994 (N_49994,N_46746,N_47994);
xnor U49995 (N_49995,N_46286,N_47143);
xor U49996 (N_49996,N_46026,N_47063);
nand U49997 (N_49997,N_46718,N_47549);
xnor U49998 (N_49998,N_47951,N_47578);
xor U49999 (N_49999,N_46179,N_47323);
or UO_0 (O_0,N_49867,N_49508);
nand UO_1 (O_1,N_48416,N_48949);
and UO_2 (O_2,N_48536,N_48284);
or UO_3 (O_3,N_48187,N_49286);
and UO_4 (O_4,N_49648,N_48725);
nor UO_5 (O_5,N_48845,N_48782);
nor UO_6 (O_6,N_49160,N_49354);
and UO_7 (O_7,N_48272,N_49891);
nand UO_8 (O_8,N_49194,N_48251);
or UO_9 (O_9,N_48367,N_49726);
or UO_10 (O_10,N_48653,N_49369);
nor UO_11 (O_11,N_48194,N_48054);
or UO_12 (O_12,N_48023,N_48963);
nand UO_13 (O_13,N_49509,N_48445);
xnor UO_14 (O_14,N_49633,N_49510);
nand UO_15 (O_15,N_49703,N_49045);
xnor UO_16 (O_16,N_49756,N_49500);
or UO_17 (O_17,N_49663,N_48684);
xor UO_18 (O_18,N_49581,N_48181);
or UO_19 (O_19,N_48326,N_48928);
or UO_20 (O_20,N_48058,N_48790);
nor UO_21 (O_21,N_48084,N_48926);
nor UO_22 (O_22,N_48520,N_49124);
nand UO_23 (O_23,N_49938,N_49747);
nor UO_24 (O_24,N_49729,N_48231);
nand UO_25 (O_25,N_48991,N_48118);
xnor UO_26 (O_26,N_49682,N_48219);
nor UO_27 (O_27,N_49972,N_48702);
nand UO_28 (O_28,N_48131,N_49088);
nor UO_29 (O_29,N_48355,N_48469);
nand UO_30 (O_30,N_49477,N_49230);
or UO_31 (O_31,N_48361,N_48739);
or UO_32 (O_32,N_49568,N_48422);
and UO_33 (O_33,N_48395,N_49918);
xor UO_34 (O_34,N_48117,N_48747);
or UO_35 (O_35,N_49454,N_48444);
or UO_36 (O_36,N_48726,N_48650);
nand UO_37 (O_37,N_48070,N_48635);
and UO_38 (O_38,N_48797,N_48851);
or UO_39 (O_39,N_49292,N_48091);
nand UO_40 (O_40,N_49934,N_48749);
xnor UO_41 (O_41,N_49854,N_48573);
or UO_42 (O_42,N_48741,N_49187);
nor UO_43 (O_43,N_48254,N_48238);
xnor UO_44 (O_44,N_48850,N_48621);
xnor UO_45 (O_45,N_48654,N_49385);
xor UO_46 (O_46,N_49481,N_49212);
xnor UO_47 (O_47,N_49567,N_49936);
or UO_48 (O_48,N_48408,N_48245);
xnor UO_49 (O_49,N_49681,N_48713);
xor UO_50 (O_50,N_49724,N_49229);
or UO_51 (O_51,N_49280,N_48529);
and UO_52 (O_52,N_49422,N_48675);
or UO_53 (O_53,N_48087,N_49870);
xnor UO_54 (O_54,N_49225,N_48328);
nand UO_55 (O_55,N_48064,N_49276);
nand UO_56 (O_56,N_48802,N_48804);
and UO_57 (O_57,N_48166,N_48410);
xnor UO_58 (O_58,N_48496,N_48167);
xnor UO_59 (O_59,N_48622,N_49328);
and UO_60 (O_60,N_49907,N_49794);
xor UO_61 (O_61,N_49770,N_49498);
or UO_62 (O_62,N_49690,N_49381);
nand UO_63 (O_63,N_49522,N_49954);
and UO_64 (O_64,N_49043,N_49266);
nand UO_65 (O_65,N_49034,N_48500);
or UO_66 (O_66,N_49023,N_48729);
nor UO_67 (O_67,N_48587,N_49413);
or UO_68 (O_68,N_48705,N_48704);
nand UO_69 (O_69,N_48431,N_48210);
nand UO_70 (O_70,N_49779,N_49634);
and UO_71 (O_71,N_49470,N_49763);
nand UO_72 (O_72,N_49262,N_49988);
nand UO_73 (O_73,N_49669,N_48728);
nor UO_74 (O_74,N_49184,N_48830);
nand UO_75 (O_75,N_48967,N_48218);
and UO_76 (O_76,N_49976,N_49616);
xor UO_77 (O_77,N_48796,N_49689);
and UO_78 (O_78,N_49909,N_48304);
or UO_79 (O_79,N_49448,N_48392);
or UO_80 (O_80,N_49281,N_48885);
xor UO_81 (O_81,N_48337,N_49984);
nor UO_82 (O_82,N_49344,N_48116);
or UO_83 (O_83,N_48225,N_49569);
xor UO_84 (O_84,N_48208,N_48917);
xnor UO_85 (O_85,N_48628,N_49159);
nand UO_86 (O_86,N_48154,N_48655);
nor UO_87 (O_87,N_49817,N_49956);
nand UO_88 (O_88,N_48482,N_49391);
xor UO_89 (O_89,N_48515,N_49361);
xor UO_90 (O_90,N_48880,N_48171);
nor UO_91 (O_91,N_48932,N_49613);
or UO_92 (O_92,N_49585,N_48871);
xor UO_93 (O_93,N_49602,N_48378);
or UO_94 (O_94,N_48464,N_48756);
or UO_95 (O_95,N_48798,N_48616);
or UO_96 (O_96,N_49371,N_48459);
xor UO_97 (O_97,N_48435,N_49645);
and UO_98 (O_98,N_49624,N_49596);
or UO_99 (O_99,N_48978,N_48115);
nand UO_100 (O_100,N_48033,N_49492);
xor UO_101 (O_101,N_48402,N_48534);
nand UO_102 (O_102,N_48307,N_48130);
nor UO_103 (O_103,N_48974,N_49929);
xnor UO_104 (O_104,N_48948,N_49363);
or UO_105 (O_105,N_48132,N_49181);
or UO_106 (O_106,N_49368,N_49675);
xnor UO_107 (O_107,N_49051,N_48895);
or UO_108 (O_108,N_48062,N_48191);
xnor UO_109 (O_109,N_49557,N_48998);
nor UO_110 (O_110,N_49488,N_48386);
nor UO_111 (O_111,N_48201,N_48776);
and UO_112 (O_112,N_49902,N_49758);
or UO_113 (O_113,N_48538,N_48810);
xor UO_114 (O_114,N_49693,N_49270);
nor UO_115 (O_115,N_48585,N_48108);
nor UO_116 (O_116,N_49259,N_49534);
and UO_117 (O_117,N_48428,N_49329);
xnor UO_118 (O_118,N_48915,N_49012);
nor UO_119 (O_119,N_49582,N_49501);
nand UO_120 (O_120,N_48638,N_48504);
nand UO_121 (O_121,N_48869,N_48122);
nor UO_122 (O_122,N_49927,N_49315);
and UO_123 (O_123,N_49811,N_49153);
xnor UO_124 (O_124,N_48818,N_49904);
or UO_125 (O_125,N_48577,N_48169);
xor UO_126 (O_126,N_48902,N_49164);
and UO_127 (O_127,N_49844,N_48574);
nor UO_128 (O_128,N_49711,N_49917);
and UO_129 (O_129,N_48282,N_48965);
nor UO_130 (O_130,N_49457,N_48910);
xor UO_131 (O_131,N_49705,N_49475);
nor UO_132 (O_132,N_49482,N_48615);
or UO_133 (O_133,N_49223,N_48458);
nor UO_134 (O_134,N_48831,N_49610);
or UO_135 (O_135,N_49553,N_48786);
and UO_136 (O_136,N_49373,N_48227);
nand UO_137 (O_137,N_48452,N_48249);
and UO_138 (O_138,N_48501,N_48050);
or UO_139 (O_139,N_48485,N_49775);
or UO_140 (O_140,N_48746,N_48570);
xor UO_141 (O_141,N_48543,N_49824);
nand UO_142 (O_142,N_48761,N_49327);
or UO_143 (O_143,N_48506,N_48490);
or UO_144 (O_144,N_48987,N_49342);
xor UO_145 (O_145,N_49774,N_48723);
nor UO_146 (O_146,N_48590,N_49263);
xor UO_147 (O_147,N_49341,N_48447);
xnor UO_148 (O_148,N_49074,N_49801);
and UO_149 (O_149,N_48698,N_48614);
and UO_150 (O_150,N_48737,N_49042);
nor UO_151 (O_151,N_48305,N_49117);
and UO_152 (O_152,N_49120,N_48775);
and UO_153 (O_153,N_48806,N_48829);
and UO_154 (O_154,N_48937,N_49411);
nor UO_155 (O_155,N_49351,N_48250);
xnor UO_156 (O_156,N_49921,N_48679);
nor UO_157 (O_157,N_48891,N_49790);
or UO_158 (O_158,N_48040,N_49535);
xnor UO_159 (O_159,N_48792,N_49089);
and UO_160 (O_160,N_49502,N_48980);
or UO_161 (O_161,N_48602,N_48579);
xor UO_162 (O_162,N_48498,N_48521);
and UO_163 (O_163,N_48817,N_49220);
nor UO_164 (O_164,N_49390,N_49039);
or UO_165 (O_165,N_48027,N_49592);
nand UO_166 (O_166,N_49096,N_49456);
nor UO_167 (O_167,N_48953,N_48528);
nor UO_168 (O_168,N_49686,N_48403);
nor UO_169 (O_169,N_48732,N_49720);
nand UO_170 (O_170,N_49980,N_49838);
nor UO_171 (O_171,N_49677,N_48834);
xnor UO_172 (O_172,N_48198,N_49766);
xor UO_173 (O_173,N_49318,N_48109);
or UO_174 (O_174,N_49472,N_49551);
xor UO_175 (O_175,N_48076,N_48007);
or UO_176 (O_176,N_49440,N_49982);
nand UO_177 (O_177,N_49374,N_49486);
nor UO_178 (O_178,N_49480,N_49186);
and UO_179 (O_179,N_49673,N_49064);
nor UO_180 (O_180,N_49964,N_48913);
or UO_181 (O_181,N_49965,N_49873);
xnor UO_182 (O_182,N_48985,N_49353);
xnor UO_183 (O_183,N_48688,N_49424);
nor UO_184 (O_184,N_48778,N_48396);
xnor UO_185 (O_185,N_48886,N_48019);
nor UO_186 (O_186,N_48276,N_49886);
xnor UO_187 (O_187,N_48162,N_48486);
nor UO_188 (O_188,N_49084,N_49771);
and UO_189 (O_189,N_48677,N_49267);
and UO_190 (O_190,N_49674,N_48009);
and UO_191 (O_191,N_49310,N_49609);
and UO_192 (O_192,N_48123,N_49299);
nand UO_193 (O_193,N_49449,N_48883);
and UO_194 (O_194,N_48159,N_49442);
nor UO_195 (O_195,N_49678,N_49393);
nand UO_196 (O_196,N_49126,N_48423);
nor UO_197 (O_197,N_48964,N_48795);
nor UO_198 (O_198,N_48681,N_48363);
and UO_199 (O_199,N_48733,N_48128);
and UO_200 (O_200,N_48188,N_49887);
xor UO_201 (O_201,N_48566,N_49661);
nand UO_202 (O_202,N_48125,N_48316);
or UO_203 (O_203,N_49129,N_49130);
nand UO_204 (O_204,N_49895,N_48352);
or UO_205 (O_205,N_48645,N_49494);
and UO_206 (O_206,N_48468,N_49762);
xnor UO_207 (O_207,N_49367,N_48517);
xnor UO_208 (O_208,N_49505,N_48211);
or UO_209 (O_209,N_48551,N_48626);
nand UO_210 (O_210,N_49713,N_49311);
nor UO_211 (O_211,N_48911,N_49094);
nand UO_212 (O_212,N_48595,N_48297);
nor UO_213 (O_213,N_49836,N_48754);
nand UO_214 (O_214,N_49722,N_48526);
xor UO_215 (O_215,N_48580,N_49764);
nand UO_216 (O_216,N_49955,N_48832);
nand UO_217 (O_217,N_48757,N_48478);
xnor UO_218 (O_218,N_49086,N_48760);
nor UO_219 (O_219,N_49197,N_49666);
xnor UO_220 (O_220,N_48646,N_48596);
nand UO_221 (O_221,N_49403,N_48450);
xor UO_222 (O_222,N_49044,N_48583);
nand UO_223 (O_223,N_49316,N_49813);
and UO_224 (O_224,N_49580,N_49093);
nand UO_225 (O_225,N_49541,N_48242);
nand UO_226 (O_226,N_48800,N_49347);
and UO_227 (O_227,N_48406,N_48014);
nor UO_228 (O_228,N_48593,N_48981);
or UO_229 (O_229,N_48957,N_49721);
xnor UO_230 (O_230,N_49366,N_48714);
and UO_231 (O_231,N_49588,N_49254);
or UO_232 (O_232,N_49935,N_48335);
and UO_233 (O_233,N_48941,N_49846);
or UO_234 (O_234,N_48642,N_49405);
or UO_235 (O_235,N_48507,N_48855);
nand UO_236 (O_236,N_48460,N_48750);
nand UO_237 (O_237,N_49214,N_49123);
xnor UO_238 (O_238,N_48068,N_49389);
nor UO_239 (O_239,N_49533,N_49637);
or UO_240 (O_240,N_49060,N_49862);
or UO_241 (O_241,N_49532,N_49820);
nor UO_242 (O_242,N_49425,N_49208);
and UO_243 (O_243,N_49611,N_49450);
or UO_244 (O_244,N_48670,N_49029);
and UO_245 (O_245,N_48461,N_49105);
nor UO_246 (O_246,N_48884,N_49038);
nor UO_247 (O_247,N_48535,N_49396);
or UO_248 (O_248,N_49467,N_48073);
nor UO_249 (O_249,N_49970,N_49036);
nor UO_250 (O_250,N_49141,N_49875);
or UO_251 (O_251,N_48145,N_48755);
nand UO_252 (O_252,N_49778,N_48502);
or UO_253 (O_253,N_49925,N_49979);
xnor UO_254 (O_254,N_49167,N_49022);
or UO_255 (O_255,N_48671,N_49962);
xnor UO_256 (O_256,N_49864,N_49708);
or UO_257 (O_257,N_49204,N_48720);
nand UO_258 (O_258,N_48510,N_49843);
and UO_259 (O_259,N_49110,N_49166);
and UO_260 (O_260,N_48303,N_48481);
or UO_261 (O_261,N_49182,N_49461);
and UO_262 (O_262,N_49783,N_49590);
and UO_263 (O_263,N_48186,N_48773);
nand UO_264 (O_264,N_49848,N_48024);
and UO_265 (O_265,N_49072,N_48152);
and UO_266 (O_266,N_49899,N_48840);
nand UO_267 (O_267,N_49701,N_48893);
nor UO_268 (O_268,N_48309,N_48685);
nor UO_269 (O_269,N_48689,N_49679);
and UO_270 (O_270,N_49489,N_48793);
and UO_271 (O_271,N_48656,N_49443);
nor UO_272 (O_272,N_49728,N_49706);
or UO_273 (O_273,N_49462,N_48598);
and UO_274 (O_274,N_48427,N_49264);
xnor UO_275 (O_275,N_48041,N_48820);
nand UO_276 (O_276,N_48588,N_49868);
or UO_277 (O_277,N_48440,N_48263);
nor UO_278 (O_278,N_49221,N_48025);
and UO_279 (O_279,N_48342,N_49863);
or UO_280 (O_280,N_48925,N_49849);
nor UO_281 (O_281,N_49050,N_48940);
nand UO_282 (O_282,N_48258,N_48081);
and UO_283 (O_283,N_49526,N_48665);
xor UO_284 (O_284,N_49295,N_49750);
nand UO_285 (O_285,N_48172,N_49542);
xor UO_286 (O_286,N_49073,N_48920);
nand UO_287 (O_287,N_48686,N_49469);
nand UO_288 (O_288,N_48943,N_48697);
nand UO_289 (O_289,N_48899,N_48321);
xor UO_290 (O_290,N_48270,N_48604);
nor UO_291 (O_291,N_48098,N_49211);
xnor UO_292 (O_292,N_48256,N_49745);
or UO_293 (O_293,N_48712,N_49217);
nand UO_294 (O_294,N_48951,N_49538);
nand UO_295 (O_295,N_49807,N_48336);
nor UO_296 (O_296,N_49205,N_48105);
and UO_297 (O_297,N_48082,N_49203);
nor UO_298 (O_298,N_48822,N_49258);
nand UO_299 (O_299,N_49598,N_49122);
or UO_300 (O_300,N_48924,N_48472);
or UO_301 (O_301,N_49201,N_49268);
and UO_302 (O_302,N_49052,N_49885);
nand UO_303 (O_303,N_49736,N_48512);
or UO_304 (O_304,N_48875,N_48405);
nand UO_305 (O_305,N_48228,N_49821);
nand UO_306 (O_306,N_48962,N_49209);
and UO_307 (O_307,N_48541,N_48864);
nor UO_308 (O_308,N_49845,N_48694);
nor UO_309 (O_309,N_49439,N_49213);
or UO_310 (O_310,N_49529,N_48072);
nor UO_311 (O_311,N_49330,N_48996);
and UO_312 (O_312,N_49063,N_49339);
and UO_313 (O_313,N_49539,N_48462);
or UO_314 (O_314,N_49246,N_49438);
nor UO_315 (O_315,N_48037,N_49162);
nand UO_316 (O_316,N_49985,N_48142);
nor UO_317 (O_317,N_48323,N_49651);
nor UO_318 (O_318,N_49404,N_48966);
and UO_319 (O_319,N_49772,N_49355);
or UO_320 (O_320,N_48914,N_48079);
and UO_321 (O_321,N_49565,N_48120);
or UO_322 (O_322,N_49865,N_48660);
xor UO_323 (O_323,N_48101,N_49314);
and UO_324 (O_324,N_49697,N_49791);
or UO_325 (O_325,N_49743,N_48680);
nor UO_326 (O_326,N_48944,N_48020);
nor UO_327 (O_327,N_49635,N_49100);
nand UO_328 (O_328,N_48483,N_49386);
or UO_329 (O_329,N_49421,N_48456);
xnor UO_330 (O_330,N_48146,N_49773);
or UO_331 (O_331,N_49748,N_48357);
nand UO_332 (O_332,N_49233,N_49995);
nor UO_333 (O_333,N_48292,N_49283);
xor UO_334 (O_334,N_49629,N_48608);
and UO_335 (O_335,N_48229,N_48111);
nor UO_336 (O_336,N_48136,N_49111);
nor UO_337 (O_337,N_48542,N_49435);
nand UO_338 (O_338,N_48599,N_49804);
and UO_339 (O_339,N_49739,N_49277);
and UO_340 (O_340,N_49416,N_48266);
or UO_341 (O_341,N_48333,N_49032);
nand UO_342 (O_342,N_49654,N_48623);
or UO_343 (O_343,N_48280,N_49178);
nand UO_344 (O_344,N_49549,N_48301);
nand UO_345 (O_345,N_49253,N_49607);
and UO_346 (O_346,N_49833,N_49829);
nand UO_347 (O_347,N_49199,N_48374);
or UO_348 (O_348,N_49603,N_48351);
xnor UO_349 (O_349,N_49087,N_49615);
or UO_350 (O_350,N_48196,N_48617);
xor UO_351 (O_351,N_48185,N_49473);
or UO_352 (O_352,N_48848,N_49892);
and UO_353 (O_353,N_49382,N_48183);
nand UO_354 (O_354,N_49937,N_48678);
or UO_355 (O_355,N_49803,N_49249);
nor UO_356 (O_356,N_48466,N_49832);
nor UO_357 (O_357,N_49798,N_48824);
xnor UO_358 (O_358,N_48411,N_48212);
or UO_359 (O_359,N_49504,N_48956);
and UO_360 (O_360,N_48606,N_48373);
or UO_361 (O_361,N_48134,N_48682);
nor UO_362 (O_362,N_49888,N_48867);
nand UO_363 (O_363,N_49983,N_48426);
xor UO_364 (O_364,N_48269,N_48066);
nand UO_365 (O_365,N_49082,N_48106);
and UO_366 (O_366,N_48764,N_48572);
and UO_367 (O_367,N_48527,N_48173);
nor UO_368 (O_368,N_49586,N_49765);
and UO_369 (O_369,N_49321,N_48006);
and UO_370 (O_370,N_48611,N_48278);
nor UO_371 (O_371,N_49952,N_49282);
xnor UO_372 (O_372,N_48121,N_49752);
xor UO_373 (O_373,N_49062,N_48013);
and UO_374 (O_374,N_48390,N_49506);
xnor UO_375 (O_375,N_48176,N_49265);
nor UO_376 (O_376,N_49710,N_49175);
or UO_377 (O_377,N_49228,N_49077);
xor UO_378 (O_378,N_48257,N_49957);
and UO_379 (O_379,N_48178,N_48619);
and UO_380 (O_380,N_48222,N_49188);
and UO_381 (O_381,N_48214,N_48584);
xnor UO_382 (O_382,N_48873,N_49638);
or UO_383 (O_383,N_49780,N_49990);
or UO_384 (O_384,N_48691,N_48799);
and UO_385 (O_385,N_49147,N_48350);
xnor UO_386 (O_386,N_48644,N_49372);
nor UO_387 (O_387,N_48341,N_48837);
and UO_388 (O_388,N_49884,N_48153);
nor UO_389 (O_389,N_48938,N_48567);
and UO_390 (O_390,N_48700,N_49815);
nand UO_391 (O_391,N_48843,N_48550);
and UO_392 (O_392,N_48643,N_48407);
and UO_393 (O_393,N_49577,N_48972);
and UO_394 (O_394,N_48494,N_48971);
and UO_395 (O_395,N_48877,N_48463);
or UO_396 (O_396,N_49576,N_48988);
and UO_397 (O_397,N_49879,N_48992);
or UO_398 (O_398,N_48339,N_49628);
nand UO_399 (O_399,N_49320,N_49376);
nand UO_400 (O_400,N_48765,N_49890);
or UO_401 (O_401,N_48385,N_49966);
and UO_402 (O_402,N_48200,N_48205);
nor UO_403 (O_403,N_48375,N_49017);
and UO_404 (O_404,N_49296,N_49789);
xor UO_405 (O_405,N_48300,N_48929);
nor UO_406 (O_406,N_49973,N_49059);
xnor UO_407 (O_407,N_49643,N_49916);
nor UO_408 (O_408,N_49346,N_48711);
nor UO_409 (O_409,N_49667,N_49119);
and UO_410 (O_410,N_48630,N_49275);
and UO_411 (O_411,N_49996,N_48067);
nand UO_412 (O_412,N_48240,N_48970);
xor UO_413 (O_413,N_49731,N_49191);
and UO_414 (O_414,N_48544,N_48641);
nor UO_415 (O_415,N_49099,N_48983);
nor UO_416 (O_416,N_49026,N_48047);
or UO_417 (O_417,N_49802,N_48320);
nor UO_418 (O_418,N_48514,N_48290);
xor UO_419 (O_419,N_48138,N_48872);
nand UO_420 (O_420,N_49793,N_49685);
nand UO_421 (O_421,N_48075,N_48449);
or UO_422 (O_422,N_48184,N_49272);
or UO_423 (O_423,N_48043,N_49920);
nand UO_424 (O_424,N_48735,N_49642);
nand UO_425 (O_425,N_48492,N_48532);
xnor UO_426 (O_426,N_49035,N_49572);
nand UO_427 (O_427,N_49800,N_49759);
or UO_428 (O_428,N_48696,N_49933);
or UO_429 (O_429,N_48839,N_49410);
nor UO_430 (O_430,N_49524,N_48640);
xor UO_431 (O_431,N_48668,N_49834);
xnor UO_432 (O_432,N_48288,N_49304);
nor UO_433 (O_433,N_48564,N_49562);
and UO_434 (O_434,N_49516,N_48874);
and UO_435 (O_435,N_49195,N_48785);
xor UO_436 (O_436,N_49109,N_48224);
nand UO_437 (O_437,N_48894,N_48192);
nor UO_438 (O_438,N_49232,N_48531);
nand UO_439 (O_439,N_49046,N_48889);
nor UO_440 (O_440,N_49942,N_49788);
xor UO_441 (O_441,N_48819,N_48457);
nor UO_442 (O_442,N_49244,N_48055);
nor UO_443 (O_443,N_49139,N_48028);
xor UO_444 (O_444,N_48330,N_49977);
nor UO_445 (O_445,N_49687,N_49735);
and UO_446 (O_446,N_48661,N_48345);
or UO_447 (O_447,N_49655,N_48846);
nand UO_448 (O_448,N_48308,N_48133);
nor UO_449 (O_449,N_48513,N_49950);
nor UO_450 (O_450,N_49787,N_48744);
or UO_451 (O_451,N_48430,N_49132);
or UO_452 (O_452,N_48364,N_48495);
or UO_453 (O_453,N_49819,N_49009);
or UO_454 (O_454,N_49563,N_48721);
nand UO_455 (O_455,N_49755,N_48939);
and UO_456 (O_456,N_49154,N_49601);
or UO_457 (O_457,N_48816,N_49290);
or UO_458 (O_458,N_48904,N_48788);
or UO_459 (O_459,N_48973,N_48752);
nor UO_460 (O_460,N_48129,N_49658);
nand UO_461 (O_461,N_49600,N_49297);
nor UO_462 (O_462,N_48419,N_49608);
nand UO_463 (O_463,N_49530,N_48056);
nor UO_464 (O_464,N_49858,N_49842);
xnor UO_465 (O_465,N_48103,N_49478);
and UO_466 (O_466,N_49460,N_49792);
xor UO_467 (O_467,N_49499,N_48576);
nor UO_468 (O_468,N_48348,N_48632);
xor UO_469 (O_469,N_48354,N_48434);
xor UO_470 (O_470,N_48794,N_48859);
and UO_471 (O_471,N_49769,N_48716);
xnor UO_472 (O_472,N_49485,N_48039);
and UO_473 (O_473,N_49158,N_48969);
and UO_474 (O_474,N_48594,N_49767);
xor UO_475 (O_475,N_48935,N_49872);
and UO_476 (O_476,N_49288,N_49531);
and UO_477 (O_477,N_48399,N_48448);
nand UO_478 (O_478,N_48947,N_49627);
xor UO_479 (O_479,N_48031,N_48371);
xor UO_480 (O_480,N_49696,N_48690);
xor UO_481 (O_481,N_48801,N_48878);
xnor UO_482 (O_482,N_49649,N_49149);
and UO_483 (O_483,N_48353,N_49922);
xnor UO_484 (O_484,N_48182,N_49877);
and UO_485 (O_485,N_48847,N_48609);
nor UO_486 (O_486,N_48809,N_49219);
nand UO_487 (O_487,N_48002,N_49468);
nand UO_488 (O_488,N_49269,N_49252);
nand UO_489 (O_489,N_49647,N_49359);
and UO_490 (O_490,N_48921,N_48581);
nor UO_491 (O_491,N_49584,N_48156);
nand UO_492 (O_492,N_49869,N_49866);
nand UO_493 (O_493,N_49234,N_49702);
or UO_494 (O_494,N_48489,N_48493);
and UO_495 (O_495,N_48627,N_48658);
nor UO_496 (O_496,N_49152,N_49926);
nor UO_497 (O_497,N_49698,N_48094);
nand UO_498 (O_498,N_48724,N_49326);
or UO_499 (O_499,N_49566,N_48215);
nor UO_500 (O_500,N_49243,N_48233);
nor UO_501 (O_501,N_48557,N_48368);
and UO_502 (O_502,N_49850,N_48057);
nand UO_503 (O_503,N_49981,N_49011);
nand UO_504 (O_504,N_48090,N_49168);
and UO_505 (O_505,N_48359,N_49463);
and UO_506 (O_506,N_48223,N_49751);
nor UO_507 (O_507,N_49128,N_49010);
or UO_508 (O_508,N_48369,N_48362);
and UO_509 (O_509,N_48479,N_48900);
or UO_510 (O_510,N_49108,N_48391);
or UO_511 (O_511,N_48015,N_49969);
or UO_512 (O_512,N_49340,N_49963);
nand UO_513 (O_513,N_49594,N_48347);
or UO_514 (O_514,N_49855,N_48346);
xor UO_515 (O_515,N_49294,N_49257);
nand UO_516 (O_516,N_49928,N_48401);
and UO_517 (O_517,N_49959,N_48078);
nor UO_518 (O_518,N_49520,N_48299);
nand UO_519 (O_519,N_49156,N_49092);
and UO_520 (O_520,N_48093,N_48701);
and UO_521 (O_521,N_48340,N_48454);
nand UO_522 (O_522,N_49835,N_49694);
nor UO_523 (O_523,N_48199,N_48505);
or UO_524 (O_524,N_49967,N_49379);
and UO_525 (O_525,N_49319,N_48918);
xor UO_526 (O_526,N_48475,N_49978);
or UO_527 (O_527,N_49453,N_49727);
nor UO_528 (O_528,N_48959,N_48530);
or UO_529 (O_529,N_49619,N_49799);
nand UO_530 (O_530,N_48865,N_49431);
nand UO_531 (O_531,N_48255,N_48995);
xor UO_532 (O_532,N_48451,N_48934);
nor UO_533 (O_533,N_48112,N_49671);
nand UO_534 (O_534,N_49112,N_49881);
nor UO_535 (O_535,N_49548,N_48139);
xnor UO_536 (O_536,N_48657,N_48388);
or UO_537 (O_537,N_48387,N_48968);
nand UO_538 (O_538,N_48265,N_48163);
xnor UO_539 (O_539,N_48383,N_48734);
nand UO_540 (O_540,N_48206,N_48545);
or UO_541 (O_541,N_48999,N_48114);
nor UO_542 (O_542,N_48104,N_49349);
xor UO_543 (O_543,N_48669,N_49595);
and UO_544 (O_544,N_48180,N_48000);
nor UO_545 (O_545,N_49714,N_48907);
and UO_546 (O_546,N_48213,N_49317);
nor UO_547 (O_547,N_49636,N_48045);
or UO_548 (O_548,N_49945,N_48285);
or UO_549 (O_549,N_48327,N_48556);
xor UO_550 (O_550,N_49248,N_49560);
nor UO_551 (O_551,N_49140,N_48738);
nand UO_552 (O_552,N_49483,N_49725);
nand UO_553 (O_553,N_49515,N_48313);
or UO_554 (O_554,N_49040,N_48085);
nand UO_555 (O_555,N_49547,N_49911);
xnor UO_556 (O_556,N_48607,N_48555);
or UO_557 (O_557,N_49554,N_49527);
and UO_558 (O_558,N_49013,N_49003);
nand UO_559 (O_559,N_49900,N_48204);
and UO_560 (O_560,N_49841,N_49019);
nand UO_561 (O_561,N_48942,N_48766);
xor UO_562 (O_562,N_48620,N_49054);
nor UO_563 (O_563,N_48035,N_48216);
nor UO_564 (O_564,N_49951,N_48325);
xor UO_565 (O_565,N_49883,N_48511);
or UO_566 (O_566,N_48438,N_49777);
nor UO_567 (O_567,N_48791,N_49298);
nor UO_568 (O_568,N_48268,N_48271);
or UO_569 (O_569,N_49536,N_48663);
and UO_570 (O_570,N_48488,N_49095);
xor UO_571 (O_571,N_48262,N_49496);
xor UO_572 (O_572,N_49362,N_49027);
and UO_573 (O_573,N_49947,N_48639);
nor UO_574 (O_574,N_48961,N_49055);
and UO_575 (O_575,N_49688,N_48993);
or UO_576 (O_576,N_48687,N_48203);
and UO_577 (O_577,N_48625,N_48415);
or UO_578 (O_578,N_48896,N_48933);
nor UO_579 (O_579,N_48437,N_49753);
and UO_580 (O_580,N_49994,N_49406);
or UO_581 (O_581,N_49014,N_48239);
nand UO_582 (O_582,N_48589,N_48842);
or UO_583 (O_583,N_49174,N_48273);
nand UO_584 (O_584,N_48077,N_48591);
and UO_585 (O_585,N_49732,N_48150);
or UO_586 (O_586,N_49507,N_49901);
nand UO_587 (O_587,N_48059,N_49662);
xor UO_588 (O_588,N_48302,N_49352);
and UO_589 (O_589,N_48155,N_49737);
xor UO_590 (O_590,N_48232,N_49511);
nor UO_591 (O_591,N_49589,N_48038);
nand UO_592 (O_592,N_49550,N_49604);
nand UO_593 (O_593,N_49325,N_49617);
xor UO_594 (O_594,N_48110,N_48575);
nor UO_595 (O_595,N_48771,N_49033);
and UO_596 (O_596,N_48158,N_48770);
nand UO_597 (O_597,N_49715,N_48709);
nor UO_598 (O_598,N_49564,N_49823);
or UO_599 (O_599,N_49402,N_49144);
or UO_600 (O_600,N_49172,N_48217);
nor UO_601 (O_601,N_49704,N_49447);
and UO_602 (O_602,N_48421,N_48561);
nor UO_603 (O_603,N_49081,N_49528);
or UO_604 (O_604,N_48293,N_48813);
xnor UO_605 (O_605,N_49897,N_49303);
or UO_606 (O_606,N_48095,N_49786);
xor UO_607 (O_607,N_49430,N_48722);
xor UO_608 (O_608,N_48294,N_48772);
nand UO_609 (O_609,N_49118,N_49313);
xnor UO_610 (O_610,N_49716,N_48672);
nand UO_611 (O_611,N_48071,N_49289);
and UO_612 (O_612,N_48414,N_49242);
xor UO_613 (O_613,N_49659,N_48016);
or UO_614 (O_614,N_48693,N_48412);
and UO_615 (O_615,N_48322,N_48174);
nor UO_616 (O_616,N_48436,N_49180);
and UO_617 (O_617,N_48052,N_49670);
or UO_618 (O_618,N_49818,N_48286);
and UO_619 (O_619,N_49006,N_48659);
nor UO_620 (O_620,N_49000,N_48311);
xor UO_621 (O_621,N_49652,N_48137);
nor UO_622 (O_622,N_48870,N_49653);
nor UO_623 (O_623,N_49968,N_49631);
nand UO_624 (O_624,N_48048,N_49948);
nand UO_625 (O_625,N_49236,N_48291);
xnor UO_626 (O_626,N_48298,N_48888);
or UO_627 (O_627,N_48274,N_49332);
and UO_628 (O_628,N_49757,N_49852);
or UO_629 (O_629,N_49024,N_48148);
nand UO_630 (O_630,N_48164,N_49031);
nor UO_631 (O_631,N_48246,N_49656);
and UO_632 (O_632,N_49738,N_49004);
or UO_633 (O_633,N_48221,N_48432);
nor UO_634 (O_634,N_48624,N_49102);
or UO_635 (O_635,N_49133,N_49387);
nand UO_636 (O_636,N_48252,N_49989);
nand UO_637 (O_637,N_49207,N_48467);
and UO_638 (O_638,N_49091,N_49273);
and UO_639 (O_639,N_48613,N_48652);
or UO_640 (O_640,N_49749,N_49556);
nand UO_641 (O_641,N_49419,N_49429);
xor UO_642 (O_642,N_48241,N_49943);
and UO_643 (O_643,N_49545,N_49131);
nand UO_644 (O_644,N_48100,N_48429);
xor UO_645 (O_645,N_49812,N_49518);
nor UO_646 (O_646,N_49345,N_49910);
nor UO_647 (O_647,N_48453,N_48636);
nand UO_648 (O_648,N_49896,N_49455);
or UO_649 (O_649,N_49474,N_48080);
or UO_650 (O_650,N_49597,N_49641);
and UO_651 (O_651,N_48289,N_49579);
nand UO_652 (O_652,N_48267,N_49445);
nor UO_653 (O_653,N_49519,N_49358);
nor UO_654 (O_654,N_49007,N_49157);
nor UO_655 (O_655,N_49047,N_49552);
or UO_656 (O_656,N_49491,N_48853);
nor UO_657 (O_657,N_48381,N_49718);
xor UO_658 (O_658,N_49444,N_49388);
nor UO_659 (O_659,N_49612,N_48424);
or UO_660 (O_660,N_49898,N_48633);
xor UO_661 (O_661,N_49037,N_48860);
and UO_662 (O_662,N_48061,N_49664);
or UO_663 (O_663,N_48719,N_49660);
and UO_664 (O_664,N_48879,N_48312);
nand UO_665 (O_665,N_48844,N_49640);
xor UO_666 (O_666,N_48209,N_49744);
nand UO_667 (O_667,N_49383,N_49949);
xor UO_668 (O_668,N_49202,N_48631);
nand UO_669 (O_669,N_48476,N_48986);
nor UO_670 (O_670,N_48170,N_49781);
nor UO_671 (O_671,N_48088,N_49002);
nor UO_672 (O_672,N_49285,N_48372);
and UO_673 (O_673,N_49741,N_48127);
xnor UO_674 (O_674,N_49993,N_49441);
xor UO_675 (O_675,N_48179,N_49200);
and UO_676 (O_676,N_48673,N_48767);
nand UO_677 (O_677,N_49723,N_48662);
or UO_678 (O_678,N_48537,N_48618);
nand UO_679 (O_679,N_49874,N_49395);
and UO_680 (O_680,N_48523,N_48751);
xnor UO_681 (O_681,N_49853,N_48807);
nor UO_682 (O_682,N_48253,N_49231);
or UO_683 (O_683,N_48897,N_49370);
xnor UO_684 (O_684,N_48010,N_49049);
or UO_685 (O_685,N_48480,N_48876);
and UO_686 (O_686,N_49495,N_48086);
nor UO_687 (O_687,N_48393,N_48823);
xor UO_688 (O_688,N_49931,N_48906);
and UO_689 (O_689,N_49476,N_49903);
nand UO_690 (O_690,N_48706,N_48936);
and UO_691 (O_691,N_49250,N_48731);
nor UO_692 (O_692,N_48803,N_48260);
xor UO_693 (O_693,N_49222,N_49312);
xnor UO_694 (O_694,N_48703,N_49930);
and UO_695 (O_695,N_49115,N_49924);
xor UO_696 (O_696,N_48692,N_49138);
nand UO_697 (O_697,N_49746,N_48945);
nor UO_698 (O_698,N_49071,N_49822);
and UO_699 (O_699,N_49226,N_49971);
and UO_700 (O_700,N_49809,N_49599);
xor UO_701 (O_701,N_49365,N_48143);
xnor UO_702 (O_702,N_48954,N_49417);
nor UO_703 (O_703,N_49493,N_49754);
nand UO_704 (O_704,N_49375,N_49356);
and UO_705 (O_705,N_49058,N_48946);
or UO_706 (O_706,N_49620,N_49490);
xnor UO_707 (O_707,N_49030,N_49255);
nor UO_708 (O_708,N_48124,N_49251);
xor UO_709 (O_709,N_49065,N_48277);
and UO_710 (O_710,N_48425,N_49805);
or UO_711 (O_711,N_49908,N_49380);
or UO_712 (O_712,N_49336,N_48315);
or UO_713 (O_713,N_48560,N_49712);
nand UO_714 (O_714,N_48318,N_48890);
and UO_715 (O_715,N_49075,N_49020);
and UO_716 (O_716,N_48230,N_48168);
or UO_717 (O_717,N_49540,N_48398);
nor UO_718 (O_718,N_48826,N_48189);
nand UO_719 (O_719,N_48261,N_49169);
and UO_720 (O_720,N_49614,N_49350);
or UO_721 (O_721,N_48365,N_49625);
nor UO_722 (O_722,N_48763,N_49171);
xnor UO_723 (O_723,N_48892,N_49061);
and UO_724 (O_724,N_49503,N_49573);
and UO_725 (O_725,N_48612,N_48912);
xor UO_726 (O_726,N_49464,N_48018);
or UO_727 (O_727,N_48649,N_49459);
xor UO_728 (O_728,N_49238,N_48140);
xor UO_729 (O_729,N_49307,N_48465);
nor UO_730 (O_730,N_48854,N_49107);
nor UO_731 (O_731,N_48379,N_48667);
xnor UO_732 (O_732,N_48065,N_49070);
xor UO_733 (O_733,N_48950,N_49960);
xnor UO_734 (O_734,N_48264,N_48519);
nand UO_735 (O_735,N_48849,N_48533);
and UO_736 (O_736,N_48439,N_49512);
or UO_737 (O_737,N_49525,N_49206);
or UO_738 (O_738,N_48976,N_49008);
and UO_739 (O_739,N_49826,N_48042);
or UO_740 (O_740,N_48787,N_48144);
nand UO_741 (O_741,N_49302,N_48955);
xor UO_742 (O_742,N_49992,N_49831);
or UO_743 (O_743,N_48443,N_48742);
xor UO_744 (O_744,N_49795,N_48597);
and UO_745 (O_745,N_49256,N_48994);
and UO_746 (O_746,N_48234,N_48769);
and UO_747 (O_747,N_48758,N_48281);
nor UO_748 (O_748,N_49067,N_49090);
and UO_749 (O_749,N_49830,N_48008);
and UO_750 (O_750,N_49322,N_48279);
or UO_751 (O_751,N_48089,N_49471);
or UO_752 (O_752,N_48474,N_48409);
nor UO_753 (O_753,N_48857,N_49436);
or UO_754 (O_754,N_48699,N_48958);
or UO_755 (O_755,N_48603,N_48394);
nor UO_756 (O_756,N_48161,N_48376);
nor UO_757 (O_757,N_49622,N_48236);
nor UO_758 (O_758,N_48119,N_49392);
xor UO_759 (O_759,N_49399,N_49083);
xnor UO_760 (O_760,N_49334,N_48828);
xnor UO_761 (O_761,N_48349,N_49048);
nor UO_762 (O_762,N_49837,N_49644);
and UO_763 (O_763,N_48919,N_48861);
and UO_764 (O_764,N_48989,N_48099);
or UO_765 (O_765,N_48605,N_49555);
and UO_766 (O_766,N_48296,N_49114);
and UO_767 (O_767,N_49426,N_49810);
nor UO_768 (O_768,N_49776,N_48382);
or UO_769 (O_769,N_48433,N_49113);
nand UO_770 (O_770,N_48730,N_49423);
nor UO_771 (O_771,N_49618,N_49218);
xnor UO_772 (O_772,N_49001,N_48400);
xnor UO_773 (O_773,N_48487,N_49384);
nor UO_774 (O_774,N_49080,N_48748);
nor UO_775 (O_775,N_49151,N_48370);
xnor UO_776 (O_776,N_48317,N_48637);
nor UO_777 (O_777,N_49401,N_49097);
and UO_778 (O_778,N_49893,N_48275);
nor UO_779 (O_779,N_48982,N_49861);
or UO_780 (O_780,N_48029,N_48306);
xor UO_781 (O_781,N_48812,N_49458);
or UO_782 (O_782,N_48647,N_48442);
and UO_783 (O_783,N_49451,N_49057);
nor UO_784 (O_784,N_49717,N_48927);
nor UO_785 (O_785,N_48207,N_49974);
and UO_786 (O_786,N_48683,N_49148);
nor UO_787 (O_787,N_49940,N_48283);
xor UO_788 (O_788,N_48473,N_49015);
nand UO_789 (O_789,N_49876,N_48762);
nor UO_790 (O_790,N_48334,N_49143);
and UO_791 (O_791,N_49291,N_48774);
nor UO_792 (O_792,N_49975,N_48707);
and UO_793 (O_793,N_48553,N_48674);
xor UO_794 (O_794,N_48516,N_48343);
or UO_795 (O_795,N_48695,N_48107);
and UO_796 (O_796,N_49487,N_49127);
xnor UO_797 (O_797,N_49466,N_49446);
nor UO_798 (O_798,N_48338,N_48177);
nor UO_799 (O_799,N_48559,N_49432);
nor UO_800 (O_800,N_49245,N_48960);
nor UO_801 (O_801,N_49606,N_48314);
nor UO_802 (O_802,N_49161,N_49828);
or UO_803 (O_803,N_48060,N_49241);
or UO_804 (O_804,N_49574,N_49986);
or UO_805 (O_805,N_49215,N_48524);
or UO_806 (O_806,N_48235,N_48011);
or UO_807 (O_807,N_48868,N_48825);
xnor UO_808 (O_808,N_48053,N_48499);
or UO_809 (O_809,N_48571,N_49394);
or UO_810 (O_810,N_48471,N_49919);
and UO_811 (O_811,N_48923,N_49906);
or UO_812 (O_812,N_49224,N_48197);
xor UO_813 (O_813,N_48835,N_49571);
or UO_814 (O_814,N_48558,N_49301);
nand UO_815 (O_815,N_49761,N_48727);
xor UO_816 (O_816,N_49076,N_48717);
xnor UO_817 (O_817,N_48592,N_49235);
xnor UO_818 (O_818,N_49335,N_48838);
or UO_819 (O_819,N_49578,N_48324);
or UO_820 (O_820,N_49626,N_49558);
or UO_821 (O_821,N_48420,N_48634);
xor UO_822 (O_822,N_48165,N_49428);
or UO_823 (O_823,N_48329,N_48046);
and UO_824 (O_824,N_49177,N_49364);
nand UO_825 (O_825,N_48247,N_48413);
or UO_826 (O_826,N_48380,N_48147);
and UO_827 (O_827,N_49190,N_49544);
xnor UO_828 (O_828,N_48858,N_48141);
and UO_829 (O_829,N_49760,N_48135);
nor UO_830 (O_830,N_49279,N_48397);
nand UO_831 (O_831,N_48777,N_49953);
nor UO_832 (O_832,N_49101,N_49135);
and UO_833 (O_833,N_48578,N_49517);
or UO_834 (O_834,N_48975,N_48666);
and UO_835 (O_835,N_48331,N_49434);
and UO_836 (O_836,N_49198,N_48195);
nor UO_837 (O_837,N_49343,N_48930);
xor UO_838 (O_838,N_49103,N_49284);
and UO_839 (O_839,N_49146,N_48833);
nand UO_840 (O_840,N_48418,N_48032);
xor UO_841 (O_841,N_49709,N_48546);
and UO_842 (O_842,N_49997,N_48220);
nand UO_843 (O_843,N_48021,N_49193);
and UO_844 (O_844,N_48049,N_48901);
xnor UO_845 (O_845,N_49857,N_48708);
nand UO_846 (O_846,N_49915,N_48518);
nor UO_847 (O_847,N_48887,N_48814);
or UO_848 (O_848,N_48562,N_49418);
nor UO_849 (O_849,N_49142,N_48916);
and UO_850 (O_850,N_49145,N_49816);
and UO_851 (O_851,N_49192,N_49839);
nor UO_852 (O_852,N_49630,N_48977);
nor UO_853 (O_853,N_48001,N_49155);
or UO_854 (O_854,N_49946,N_48477);
nor UO_855 (O_855,N_48193,N_48017);
nand UO_856 (O_856,N_48753,N_49913);
nand UO_857 (O_857,N_49878,N_49360);
nand UO_858 (O_858,N_48012,N_49437);
xor UO_859 (O_859,N_49397,N_48190);
nand UO_860 (O_860,N_49665,N_49293);
xor UO_861 (O_861,N_48470,N_48175);
or UO_862 (O_862,N_49137,N_49591);
nor UO_863 (O_863,N_49639,N_49657);
nor UO_864 (O_864,N_49991,N_48126);
or UO_865 (O_865,N_49210,N_48781);
nand UO_866 (O_866,N_49987,N_49859);
or UO_867 (O_867,N_49150,N_49587);
nor UO_868 (O_868,N_49079,N_48484);
or UO_869 (O_869,N_48149,N_49537);
nor UO_870 (O_870,N_48783,N_48990);
nand UO_871 (O_871,N_48569,N_49427);
nand UO_872 (O_872,N_48931,N_48881);
xnor UO_873 (O_873,N_48287,N_49707);
or UO_874 (O_874,N_48821,N_49176);
or UO_875 (O_875,N_49814,N_48811);
xor UO_876 (O_876,N_48295,N_49905);
nor UO_877 (O_877,N_48003,N_48759);
xor UO_878 (O_878,N_49605,N_49683);
nand UO_879 (O_879,N_49078,N_49348);
xnor UO_880 (O_880,N_48805,N_49840);
xor UO_881 (O_881,N_49196,N_49583);
or UO_882 (O_882,N_48952,N_49561);
nor UO_883 (O_883,N_49337,N_49333);
nor UO_884 (O_884,N_49570,N_49623);
xor UO_885 (O_885,N_48344,N_49308);
nand UO_886 (O_886,N_49338,N_49247);
or UO_887 (O_887,N_48243,N_48074);
xor UO_888 (O_888,N_49871,N_48736);
xnor UO_889 (O_889,N_48083,N_48908);
or UO_890 (O_890,N_49808,N_49733);
and UO_891 (O_891,N_48610,N_48866);
or UO_892 (O_892,N_49378,N_49260);
nor UO_893 (O_893,N_49880,N_48548);
and UO_894 (O_894,N_49894,N_49066);
or UO_895 (O_895,N_48202,N_48898);
nor UO_896 (O_896,N_48092,N_48565);
xor UO_897 (O_897,N_48384,N_48568);
or UO_898 (O_898,N_49085,N_49240);
nand UO_899 (O_899,N_49912,N_48366);
nor UO_900 (O_900,N_48856,N_48780);
nand UO_901 (O_901,N_49415,N_48922);
nor UO_902 (O_902,N_48539,N_48836);
xnor UO_903 (O_903,N_48508,N_48446);
nor UO_904 (O_904,N_48356,N_49484);
nand UO_905 (O_905,N_49695,N_48248);
and UO_906 (O_906,N_49742,N_48417);
xor UO_907 (O_907,N_48743,N_48069);
and UO_908 (O_908,N_48863,N_49796);
nor UO_909 (O_909,N_48022,N_49409);
nand UO_910 (O_910,N_49331,N_49523);
xor UO_911 (O_911,N_48651,N_48903);
and UO_912 (O_912,N_49684,N_49400);
nand UO_913 (O_913,N_48034,N_48718);
nand UO_914 (O_914,N_49408,N_49237);
and UO_915 (O_915,N_49136,N_49125);
nand UO_916 (O_916,N_48882,N_49691);
or UO_917 (O_917,N_48151,N_49261);
xnor UO_918 (O_918,N_48740,N_48497);
xnor UO_919 (O_919,N_48789,N_49797);
nand UO_920 (O_920,N_48710,N_49740);
or UO_921 (O_921,N_48455,N_48113);
nor UO_922 (O_922,N_49170,N_49041);
or UO_923 (O_923,N_48503,N_49021);
nor UO_924 (O_924,N_48096,N_49121);
nor UO_925 (O_925,N_49768,N_49069);
nor UO_926 (O_926,N_49305,N_49407);
nand UO_927 (O_927,N_49414,N_49546);
or UO_928 (O_928,N_49961,N_48051);
xor UO_929 (O_929,N_48582,N_48044);
or UO_930 (O_930,N_48815,N_49668);
xor UO_931 (O_931,N_49521,N_49699);
nor UO_932 (O_932,N_48779,N_49827);
xor UO_933 (O_933,N_49999,N_49104);
xor UO_934 (O_934,N_49646,N_49514);
xor UO_935 (O_935,N_48036,N_48097);
nor UO_936 (O_936,N_49719,N_49497);
nand UO_937 (O_937,N_48549,N_49018);
nand UO_938 (O_938,N_48310,N_49851);
nor UO_939 (O_939,N_49882,N_49889);
and UO_940 (O_940,N_49412,N_49274);
xnor UO_941 (O_941,N_49513,N_49825);
xnor UO_942 (O_942,N_48244,N_49632);
nor UO_943 (O_943,N_49559,N_49692);
or UO_944 (O_944,N_49806,N_49183);
xor UO_945 (O_945,N_49116,N_48030);
nand UO_946 (O_946,N_48862,N_48997);
xor UO_947 (O_947,N_48601,N_49543);
nand UO_948 (O_948,N_48441,N_48491);
and UO_949 (O_949,N_49785,N_49398);
or UO_950 (O_950,N_48629,N_48404);
and UO_951 (O_951,N_49324,N_49593);
or UO_952 (O_952,N_48160,N_49860);
xnor UO_953 (O_953,N_48509,N_49165);
nand UO_954 (O_954,N_49958,N_49056);
and UO_955 (O_955,N_49784,N_48676);
and UO_956 (O_956,N_48226,N_48237);
nor UO_957 (O_957,N_48026,N_48827);
xnor UO_958 (O_958,N_49377,N_48319);
nand UO_959 (O_959,N_49098,N_49433);
xor UO_960 (O_960,N_48525,N_48979);
nor UO_961 (O_961,N_49227,N_49621);
nand UO_962 (O_962,N_48005,N_48358);
nand UO_963 (O_963,N_48332,N_49189);
and UO_964 (O_964,N_49734,N_48984);
or UO_965 (O_965,N_48715,N_49680);
nand UO_966 (O_966,N_48389,N_49025);
or UO_967 (O_967,N_49163,N_49300);
nor UO_968 (O_968,N_49700,N_48768);
nand UO_969 (O_969,N_48157,N_48648);
and UO_970 (O_970,N_49028,N_49185);
or UO_971 (O_971,N_48905,N_49005);
or UO_972 (O_972,N_49134,N_49106);
xnor UO_973 (O_973,N_49944,N_49016);
or UO_974 (O_974,N_49782,N_49939);
nand UO_975 (O_975,N_48522,N_49287);
xor UO_976 (O_976,N_48377,N_49278);
xor UO_977 (O_977,N_48841,N_48102);
or UO_978 (O_978,N_49452,N_48547);
nor UO_979 (O_979,N_49420,N_49672);
xor UO_980 (O_980,N_49179,N_49309);
nand UO_981 (O_981,N_49053,N_48784);
and UO_982 (O_982,N_49357,N_49856);
nor UO_983 (O_983,N_49173,N_49941);
nor UO_984 (O_984,N_48600,N_48004);
and UO_985 (O_985,N_48259,N_49923);
and UO_986 (O_986,N_48540,N_49068);
nor UO_987 (O_987,N_48563,N_48586);
nand UO_988 (O_988,N_49932,N_49271);
nand UO_989 (O_989,N_49730,N_49323);
nand UO_990 (O_990,N_48808,N_48909);
or UO_991 (O_991,N_48664,N_49650);
nor UO_992 (O_992,N_48745,N_49216);
xnor UO_993 (O_993,N_49479,N_49914);
and UO_994 (O_994,N_48552,N_48360);
xnor UO_995 (O_995,N_49306,N_49676);
and UO_996 (O_996,N_49998,N_49847);
nand UO_997 (O_997,N_49575,N_48063);
or UO_998 (O_998,N_49239,N_48554);
nor UO_999 (O_999,N_49465,N_48852);
nand UO_1000 (O_1000,N_48093,N_48164);
and UO_1001 (O_1001,N_49728,N_49055);
nor UO_1002 (O_1002,N_49149,N_49081);
nand UO_1003 (O_1003,N_49736,N_48728);
or UO_1004 (O_1004,N_49097,N_49789);
nand UO_1005 (O_1005,N_49770,N_48720);
or UO_1006 (O_1006,N_49926,N_48245);
xor UO_1007 (O_1007,N_49393,N_48892);
xnor UO_1008 (O_1008,N_49745,N_49262);
or UO_1009 (O_1009,N_48406,N_48796);
nor UO_1010 (O_1010,N_49613,N_49409);
xor UO_1011 (O_1011,N_48143,N_48669);
nand UO_1012 (O_1012,N_49027,N_49764);
nor UO_1013 (O_1013,N_49995,N_48737);
or UO_1014 (O_1014,N_48315,N_48429);
nor UO_1015 (O_1015,N_49802,N_49681);
xnor UO_1016 (O_1016,N_49586,N_48443);
and UO_1017 (O_1017,N_48449,N_48223);
xor UO_1018 (O_1018,N_49189,N_49262);
nor UO_1019 (O_1019,N_48373,N_48791);
nand UO_1020 (O_1020,N_48332,N_49751);
or UO_1021 (O_1021,N_48896,N_48347);
or UO_1022 (O_1022,N_48659,N_48746);
nor UO_1023 (O_1023,N_48067,N_48460);
and UO_1024 (O_1024,N_48787,N_49231);
xor UO_1025 (O_1025,N_49856,N_49685);
nor UO_1026 (O_1026,N_49211,N_48146);
and UO_1027 (O_1027,N_48929,N_48346);
nand UO_1028 (O_1028,N_48160,N_49792);
and UO_1029 (O_1029,N_48432,N_49881);
xor UO_1030 (O_1030,N_48095,N_48413);
and UO_1031 (O_1031,N_48691,N_49771);
and UO_1032 (O_1032,N_49516,N_48251);
or UO_1033 (O_1033,N_48812,N_49109);
nor UO_1034 (O_1034,N_49408,N_49688);
or UO_1035 (O_1035,N_48761,N_49185);
nand UO_1036 (O_1036,N_49852,N_49657);
xnor UO_1037 (O_1037,N_49313,N_49150);
xnor UO_1038 (O_1038,N_49780,N_48222);
nand UO_1039 (O_1039,N_49765,N_49195);
nor UO_1040 (O_1040,N_49594,N_49444);
or UO_1041 (O_1041,N_49747,N_49586);
nor UO_1042 (O_1042,N_49552,N_49990);
nor UO_1043 (O_1043,N_48140,N_49796);
or UO_1044 (O_1044,N_49108,N_48555);
xor UO_1045 (O_1045,N_49626,N_49475);
and UO_1046 (O_1046,N_49702,N_48244);
or UO_1047 (O_1047,N_49076,N_49196);
nor UO_1048 (O_1048,N_49045,N_49647);
xnor UO_1049 (O_1049,N_49334,N_49579);
or UO_1050 (O_1050,N_48086,N_48244);
nor UO_1051 (O_1051,N_48490,N_49415);
and UO_1052 (O_1052,N_48482,N_48346);
xor UO_1053 (O_1053,N_49247,N_49446);
or UO_1054 (O_1054,N_49972,N_48906);
and UO_1055 (O_1055,N_48336,N_49203);
or UO_1056 (O_1056,N_48485,N_49751);
and UO_1057 (O_1057,N_49721,N_49150);
xnor UO_1058 (O_1058,N_49256,N_49939);
or UO_1059 (O_1059,N_48916,N_49290);
nand UO_1060 (O_1060,N_49675,N_49347);
xor UO_1061 (O_1061,N_49425,N_48378);
nand UO_1062 (O_1062,N_48099,N_49876);
or UO_1063 (O_1063,N_48160,N_49473);
or UO_1064 (O_1064,N_48434,N_49693);
or UO_1065 (O_1065,N_48019,N_48740);
nor UO_1066 (O_1066,N_48700,N_48221);
and UO_1067 (O_1067,N_49843,N_49260);
nand UO_1068 (O_1068,N_48421,N_49681);
nor UO_1069 (O_1069,N_48830,N_49890);
and UO_1070 (O_1070,N_49998,N_49241);
or UO_1071 (O_1071,N_49044,N_49788);
or UO_1072 (O_1072,N_49211,N_49001);
nand UO_1073 (O_1073,N_49222,N_49114);
or UO_1074 (O_1074,N_49377,N_48292);
and UO_1075 (O_1075,N_48008,N_49432);
nor UO_1076 (O_1076,N_49617,N_49579);
and UO_1077 (O_1077,N_49696,N_48102);
nand UO_1078 (O_1078,N_49290,N_48745);
or UO_1079 (O_1079,N_48248,N_48056);
or UO_1080 (O_1080,N_48349,N_48698);
nand UO_1081 (O_1081,N_48651,N_49368);
and UO_1082 (O_1082,N_49784,N_48061);
xnor UO_1083 (O_1083,N_48664,N_49611);
and UO_1084 (O_1084,N_49836,N_48039);
xor UO_1085 (O_1085,N_48201,N_48541);
nor UO_1086 (O_1086,N_49150,N_49700);
nand UO_1087 (O_1087,N_49953,N_49127);
and UO_1088 (O_1088,N_49003,N_49951);
xnor UO_1089 (O_1089,N_48948,N_48186);
nand UO_1090 (O_1090,N_48164,N_49623);
nor UO_1091 (O_1091,N_49378,N_49040);
or UO_1092 (O_1092,N_49363,N_49017);
nor UO_1093 (O_1093,N_48089,N_49229);
xor UO_1094 (O_1094,N_49729,N_48741);
nand UO_1095 (O_1095,N_48311,N_49082);
xor UO_1096 (O_1096,N_48204,N_48942);
and UO_1097 (O_1097,N_48583,N_48140);
nand UO_1098 (O_1098,N_48325,N_49025);
and UO_1099 (O_1099,N_48597,N_49222);
xor UO_1100 (O_1100,N_49061,N_49051);
nor UO_1101 (O_1101,N_49899,N_48296);
xnor UO_1102 (O_1102,N_48220,N_49953);
nand UO_1103 (O_1103,N_48573,N_48730);
or UO_1104 (O_1104,N_49101,N_49017);
nand UO_1105 (O_1105,N_48981,N_49484);
and UO_1106 (O_1106,N_49092,N_48761);
nor UO_1107 (O_1107,N_49825,N_48361);
xor UO_1108 (O_1108,N_48791,N_48808);
xor UO_1109 (O_1109,N_48641,N_48588);
xor UO_1110 (O_1110,N_48454,N_48563);
or UO_1111 (O_1111,N_48875,N_48594);
and UO_1112 (O_1112,N_48717,N_48755);
xor UO_1113 (O_1113,N_49423,N_48702);
nor UO_1114 (O_1114,N_48412,N_48644);
or UO_1115 (O_1115,N_48116,N_49275);
nor UO_1116 (O_1116,N_49792,N_48652);
or UO_1117 (O_1117,N_49965,N_49343);
nand UO_1118 (O_1118,N_48763,N_48031);
and UO_1119 (O_1119,N_49979,N_48544);
nor UO_1120 (O_1120,N_48819,N_48790);
and UO_1121 (O_1121,N_49223,N_48816);
and UO_1122 (O_1122,N_49761,N_49010);
or UO_1123 (O_1123,N_49289,N_49473);
nor UO_1124 (O_1124,N_48978,N_49152);
or UO_1125 (O_1125,N_48055,N_49792);
or UO_1126 (O_1126,N_48916,N_49319);
nand UO_1127 (O_1127,N_48595,N_49393);
or UO_1128 (O_1128,N_49331,N_48632);
nor UO_1129 (O_1129,N_49398,N_49589);
nand UO_1130 (O_1130,N_48245,N_49795);
nand UO_1131 (O_1131,N_48007,N_48406);
nor UO_1132 (O_1132,N_48728,N_49322);
nand UO_1133 (O_1133,N_49132,N_49837);
xnor UO_1134 (O_1134,N_49222,N_48686);
and UO_1135 (O_1135,N_49667,N_49124);
and UO_1136 (O_1136,N_49716,N_49791);
and UO_1137 (O_1137,N_49354,N_49615);
or UO_1138 (O_1138,N_48040,N_49779);
nor UO_1139 (O_1139,N_48775,N_49126);
nand UO_1140 (O_1140,N_48585,N_49516);
xor UO_1141 (O_1141,N_48850,N_48342);
and UO_1142 (O_1142,N_49651,N_49099);
and UO_1143 (O_1143,N_48934,N_49576);
nand UO_1144 (O_1144,N_49962,N_48108);
nand UO_1145 (O_1145,N_49676,N_49748);
and UO_1146 (O_1146,N_49693,N_49196);
xor UO_1147 (O_1147,N_48772,N_48414);
nand UO_1148 (O_1148,N_48495,N_49910);
nand UO_1149 (O_1149,N_49561,N_48540);
nor UO_1150 (O_1150,N_49086,N_48587);
nor UO_1151 (O_1151,N_48100,N_49896);
and UO_1152 (O_1152,N_49644,N_49907);
xnor UO_1153 (O_1153,N_49076,N_49534);
xor UO_1154 (O_1154,N_48045,N_48844);
nand UO_1155 (O_1155,N_49523,N_48760);
or UO_1156 (O_1156,N_49803,N_48003);
and UO_1157 (O_1157,N_48451,N_49568);
and UO_1158 (O_1158,N_48304,N_49015);
nand UO_1159 (O_1159,N_49588,N_49115);
nor UO_1160 (O_1160,N_48734,N_49404);
nand UO_1161 (O_1161,N_48636,N_48273);
nand UO_1162 (O_1162,N_49968,N_48016);
and UO_1163 (O_1163,N_49862,N_48052);
and UO_1164 (O_1164,N_49178,N_48110);
and UO_1165 (O_1165,N_49636,N_49613);
xnor UO_1166 (O_1166,N_49758,N_48752);
or UO_1167 (O_1167,N_49379,N_49708);
nand UO_1168 (O_1168,N_48125,N_49591);
nor UO_1169 (O_1169,N_49711,N_48616);
xor UO_1170 (O_1170,N_49437,N_48206);
nand UO_1171 (O_1171,N_48392,N_48383);
nor UO_1172 (O_1172,N_49912,N_48609);
and UO_1173 (O_1173,N_48572,N_49873);
nor UO_1174 (O_1174,N_49533,N_49461);
nor UO_1175 (O_1175,N_49834,N_48505);
and UO_1176 (O_1176,N_49868,N_49148);
or UO_1177 (O_1177,N_49860,N_48732);
or UO_1178 (O_1178,N_49838,N_49482);
nand UO_1179 (O_1179,N_48353,N_49807);
nor UO_1180 (O_1180,N_48788,N_49512);
and UO_1181 (O_1181,N_49479,N_48994);
nor UO_1182 (O_1182,N_48881,N_48005);
nand UO_1183 (O_1183,N_48244,N_48051);
nand UO_1184 (O_1184,N_49937,N_48237);
and UO_1185 (O_1185,N_49802,N_48033);
and UO_1186 (O_1186,N_49571,N_49863);
nand UO_1187 (O_1187,N_49829,N_48616);
and UO_1188 (O_1188,N_49052,N_48217);
or UO_1189 (O_1189,N_48899,N_49237);
nand UO_1190 (O_1190,N_49812,N_49004);
nor UO_1191 (O_1191,N_49947,N_48875);
nand UO_1192 (O_1192,N_49691,N_49031);
or UO_1193 (O_1193,N_48999,N_49654);
or UO_1194 (O_1194,N_48570,N_48803);
xor UO_1195 (O_1195,N_48605,N_49320);
and UO_1196 (O_1196,N_48382,N_48428);
and UO_1197 (O_1197,N_48146,N_48423);
nand UO_1198 (O_1198,N_48239,N_48281);
or UO_1199 (O_1199,N_48346,N_49532);
or UO_1200 (O_1200,N_49339,N_48442);
nor UO_1201 (O_1201,N_49558,N_48305);
nand UO_1202 (O_1202,N_48817,N_49637);
nor UO_1203 (O_1203,N_49805,N_49684);
nand UO_1204 (O_1204,N_48412,N_49000);
xnor UO_1205 (O_1205,N_48105,N_49788);
nand UO_1206 (O_1206,N_48617,N_49367);
and UO_1207 (O_1207,N_49662,N_49935);
or UO_1208 (O_1208,N_48674,N_48112);
nor UO_1209 (O_1209,N_49065,N_49700);
xor UO_1210 (O_1210,N_48596,N_48918);
nand UO_1211 (O_1211,N_48266,N_48130);
xor UO_1212 (O_1212,N_49922,N_48840);
xnor UO_1213 (O_1213,N_49165,N_48582);
or UO_1214 (O_1214,N_48356,N_49797);
nand UO_1215 (O_1215,N_48795,N_48211);
xnor UO_1216 (O_1216,N_48517,N_48126);
and UO_1217 (O_1217,N_49815,N_49865);
nor UO_1218 (O_1218,N_48261,N_48000);
nor UO_1219 (O_1219,N_49093,N_49973);
nor UO_1220 (O_1220,N_48917,N_49845);
xnor UO_1221 (O_1221,N_48723,N_48550);
xnor UO_1222 (O_1222,N_49450,N_48531);
or UO_1223 (O_1223,N_48528,N_48603);
or UO_1224 (O_1224,N_49909,N_48128);
nand UO_1225 (O_1225,N_48385,N_49439);
or UO_1226 (O_1226,N_48974,N_48259);
or UO_1227 (O_1227,N_49116,N_48819);
and UO_1228 (O_1228,N_48463,N_49692);
nand UO_1229 (O_1229,N_48709,N_49746);
and UO_1230 (O_1230,N_48816,N_48705);
and UO_1231 (O_1231,N_49246,N_48898);
xor UO_1232 (O_1232,N_49567,N_48249);
xor UO_1233 (O_1233,N_48359,N_49808);
nor UO_1234 (O_1234,N_49357,N_48495);
nand UO_1235 (O_1235,N_48387,N_49701);
nand UO_1236 (O_1236,N_48946,N_48119);
nand UO_1237 (O_1237,N_49442,N_48733);
xor UO_1238 (O_1238,N_49404,N_48458);
nand UO_1239 (O_1239,N_49365,N_49125);
and UO_1240 (O_1240,N_48416,N_48298);
nand UO_1241 (O_1241,N_48961,N_49040);
nor UO_1242 (O_1242,N_48393,N_48523);
or UO_1243 (O_1243,N_49613,N_49892);
nor UO_1244 (O_1244,N_49022,N_49587);
xnor UO_1245 (O_1245,N_49082,N_49077);
xor UO_1246 (O_1246,N_48329,N_49907);
and UO_1247 (O_1247,N_48960,N_48449);
nand UO_1248 (O_1248,N_49832,N_49857);
nor UO_1249 (O_1249,N_49817,N_48247);
nand UO_1250 (O_1250,N_49845,N_48896);
or UO_1251 (O_1251,N_49338,N_48238);
and UO_1252 (O_1252,N_48027,N_49776);
and UO_1253 (O_1253,N_49723,N_48107);
nand UO_1254 (O_1254,N_49813,N_49657);
or UO_1255 (O_1255,N_49249,N_48734);
and UO_1256 (O_1256,N_49054,N_49421);
nand UO_1257 (O_1257,N_48354,N_48600);
and UO_1258 (O_1258,N_49195,N_48405);
and UO_1259 (O_1259,N_48077,N_49681);
and UO_1260 (O_1260,N_49279,N_49571);
nand UO_1261 (O_1261,N_48029,N_49296);
xnor UO_1262 (O_1262,N_49638,N_49096);
xnor UO_1263 (O_1263,N_49564,N_48524);
nor UO_1264 (O_1264,N_49389,N_49776);
or UO_1265 (O_1265,N_49213,N_49129);
nor UO_1266 (O_1266,N_49563,N_48231);
xor UO_1267 (O_1267,N_48519,N_49904);
and UO_1268 (O_1268,N_49995,N_48114);
or UO_1269 (O_1269,N_49501,N_48631);
or UO_1270 (O_1270,N_48017,N_49058);
xnor UO_1271 (O_1271,N_48786,N_49832);
nand UO_1272 (O_1272,N_48254,N_48929);
nand UO_1273 (O_1273,N_48339,N_49283);
and UO_1274 (O_1274,N_48271,N_49980);
or UO_1275 (O_1275,N_49238,N_48604);
xor UO_1276 (O_1276,N_49644,N_49688);
nor UO_1277 (O_1277,N_49784,N_49316);
nor UO_1278 (O_1278,N_49279,N_48236);
and UO_1279 (O_1279,N_49267,N_48949);
and UO_1280 (O_1280,N_48532,N_48795);
nand UO_1281 (O_1281,N_48228,N_48598);
nor UO_1282 (O_1282,N_48324,N_49775);
or UO_1283 (O_1283,N_48500,N_49411);
nor UO_1284 (O_1284,N_49221,N_49793);
and UO_1285 (O_1285,N_48987,N_48315);
nand UO_1286 (O_1286,N_48543,N_49869);
and UO_1287 (O_1287,N_48830,N_49403);
nor UO_1288 (O_1288,N_49196,N_49683);
nand UO_1289 (O_1289,N_49263,N_49793);
and UO_1290 (O_1290,N_48497,N_49048);
xor UO_1291 (O_1291,N_48949,N_49064);
or UO_1292 (O_1292,N_49172,N_49348);
nor UO_1293 (O_1293,N_49686,N_48943);
and UO_1294 (O_1294,N_48920,N_48108);
nand UO_1295 (O_1295,N_49190,N_48686);
or UO_1296 (O_1296,N_49111,N_48258);
and UO_1297 (O_1297,N_49833,N_49053);
or UO_1298 (O_1298,N_48857,N_48559);
or UO_1299 (O_1299,N_48607,N_48057);
and UO_1300 (O_1300,N_48093,N_48436);
and UO_1301 (O_1301,N_48150,N_48440);
nor UO_1302 (O_1302,N_48873,N_48719);
nand UO_1303 (O_1303,N_49650,N_49863);
nor UO_1304 (O_1304,N_48722,N_49500);
or UO_1305 (O_1305,N_48249,N_49616);
nor UO_1306 (O_1306,N_48445,N_48912);
and UO_1307 (O_1307,N_49843,N_49267);
xor UO_1308 (O_1308,N_48979,N_48485);
or UO_1309 (O_1309,N_49073,N_48518);
xnor UO_1310 (O_1310,N_48451,N_49752);
or UO_1311 (O_1311,N_49135,N_48805);
and UO_1312 (O_1312,N_48168,N_48454);
or UO_1313 (O_1313,N_48842,N_48253);
nor UO_1314 (O_1314,N_48772,N_49900);
or UO_1315 (O_1315,N_48537,N_49863);
xor UO_1316 (O_1316,N_48826,N_49885);
nand UO_1317 (O_1317,N_49402,N_48316);
and UO_1318 (O_1318,N_48057,N_49801);
xnor UO_1319 (O_1319,N_49659,N_48615);
and UO_1320 (O_1320,N_49693,N_48214);
xor UO_1321 (O_1321,N_48727,N_49277);
nand UO_1322 (O_1322,N_49910,N_48857);
and UO_1323 (O_1323,N_48633,N_49688);
and UO_1324 (O_1324,N_48643,N_48315);
or UO_1325 (O_1325,N_48945,N_49570);
nand UO_1326 (O_1326,N_48408,N_48871);
and UO_1327 (O_1327,N_49984,N_49006);
or UO_1328 (O_1328,N_48788,N_48454);
and UO_1329 (O_1329,N_49613,N_48280);
xnor UO_1330 (O_1330,N_48680,N_48900);
and UO_1331 (O_1331,N_49291,N_49490);
and UO_1332 (O_1332,N_49755,N_49938);
or UO_1333 (O_1333,N_48901,N_48863);
xnor UO_1334 (O_1334,N_48457,N_48356);
nand UO_1335 (O_1335,N_49807,N_49790);
nor UO_1336 (O_1336,N_48164,N_49227);
xor UO_1337 (O_1337,N_48658,N_49378);
or UO_1338 (O_1338,N_49954,N_49986);
and UO_1339 (O_1339,N_49604,N_49877);
xor UO_1340 (O_1340,N_49270,N_49947);
xor UO_1341 (O_1341,N_48196,N_49204);
or UO_1342 (O_1342,N_48720,N_49161);
nand UO_1343 (O_1343,N_49832,N_49508);
xnor UO_1344 (O_1344,N_49882,N_48999);
nand UO_1345 (O_1345,N_49996,N_49125);
and UO_1346 (O_1346,N_48642,N_49468);
and UO_1347 (O_1347,N_49856,N_48016);
nor UO_1348 (O_1348,N_49291,N_48235);
xnor UO_1349 (O_1349,N_48927,N_48452);
nor UO_1350 (O_1350,N_49001,N_48230);
or UO_1351 (O_1351,N_48104,N_48591);
xnor UO_1352 (O_1352,N_48474,N_48478);
nor UO_1353 (O_1353,N_48068,N_48722);
and UO_1354 (O_1354,N_49680,N_49968);
xnor UO_1355 (O_1355,N_49798,N_48460);
or UO_1356 (O_1356,N_49939,N_48628);
and UO_1357 (O_1357,N_49920,N_49157);
nand UO_1358 (O_1358,N_48030,N_48967);
or UO_1359 (O_1359,N_49698,N_48772);
nor UO_1360 (O_1360,N_48654,N_48379);
xor UO_1361 (O_1361,N_49246,N_49032);
or UO_1362 (O_1362,N_49895,N_49787);
nand UO_1363 (O_1363,N_48746,N_48045);
nor UO_1364 (O_1364,N_48866,N_48714);
nor UO_1365 (O_1365,N_49994,N_49709);
or UO_1366 (O_1366,N_48968,N_49708);
and UO_1367 (O_1367,N_48925,N_48788);
and UO_1368 (O_1368,N_48629,N_49583);
nor UO_1369 (O_1369,N_49832,N_48941);
nor UO_1370 (O_1370,N_48589,N_49739);
and UO_1371 (O_1371,N_49707,N_49808);
nand UO_1372 (O_1372,N_49452,N_49434);
and UO_1373 (O_1373,N_48584,N_49562);
or UO_1374 (O_1374,N_48098,N_48373);
or UO_1375 (O_1375,N_49831,N_49086);
or UO_1376 (O_1376,N_49835,N_49373);
nand UO_1377 (O_1377,N_48583,N_48371);
nand UO_1378 (O_1378,N_49593,N_48821);
xnor UO_1379 (O_1379,N_48734,N_49223);
and UO_1380 (O_1380,N_49923,N_49100);
xnor UO_1381 (O_1381,N_48716,N_49339);
nand UO_1382 (O_1382,N_48017,N_48359);
nand UO_1383 (O_1383,N_49390,N_48517);
xor UO_1384 (O_1384,N_48856,N_49421);
and UO_1385 (O_1385,N_49885,N_48310);
nor UO_1386 (O_1386,N_49566,N_48605);
nor UO_1387 (O_1387,N_49613,N_48249);
xor UO_1388 (O_1388,N_48309,N_49600);
and UO_1389 (O_1389,N_49125,N_48218);
and UO_1390 (O_1390,N_49627,N_48386);
and UO_1391 (O_1391,N_49155,N_49007);
and UO_1392 (O_1392,N_48312,N_48733);
or UO_1393 (O_1393,N_49121,N_49069);
nor UO_1394 (O_1394,N_49228,N_49968);
nand UO_1395 (O_1395,N_48225,N_49381);
or UO_1396 (O_1396,N_49662,N_49946);
and UO_1397 (O_1397,N_49446,N_48862);
xnor UO_1398 (O_1398,N_49227,N_48346);
and UO_1399 (O_1399,N_49531,N_48173);
and UO_1400 (O_1400,N_49958,N_49301);
xnor UO_1401 (O_1401,N_48053,N_49589);
or UO_1402 (O_1402,N_48441,N_49624);
and UO_1403 (O_1403,N_49586,N_49414);
and UO_1404 (O_1404,N_49497,N_48514);
or UO_1405 (O_1405,N_48172,N_49963);
or UO_1406 (O_1406,N_49062,N_49180);
nor UO_1407 (O_1407,N_48839,N_49781);
nor UO_1408 (O_1408,N_48922,N_48421);
nor UO_1409 (O_1409,N_48664,N_48197);
and UO_1410 (O_1410,N_48963,N_48870);
or UO_1411 (O_1411,N_49407,N_48855);
xor UO_1412 (O_1412,N_48541,N_48474);
nand UO_1413 (O_1413,N_49988,N_48141);
or UO_1414 (O_1414,N_48365,N_48054);
or UO_1415 (O_1415,N_49687,N_48387);
or UO_1416 (O_1416,N_48658,N_48706);
nand UO_1417 (O_1417,N_48498,N_48052);
or UO_1418 (O_1418,N_48772,N_49233);
nand UO_1419 (O_1419,N_49719,N_49289);
and UO_1420 (O_1420,N_49783,N_48546);
and UO_1421 (O_1421,N_48727,N_49122);
or UO_1422 (O_1422,N_49608,N_48970);
and UO_1423 (O_1423,N_48526,N_49577);
or UO_1424 (O_1424,N_48558,N_48631);
nor UO_1425 (O_1425,N_48393,N_49548);
or UO_1426 (O_1426,N_49546,N_48246);
nor UO_1427 (O_1427,N_49882,N_49393);
nand UO_1428 (O_1428,N_49708,N_48950);
and UO_1429 (O_1429,N_49492,N_48536);
nor UO_1430 (O_1430,N_48164,N_48200);
or UO_1431 (O_1431,N_49412,N_48216);
nor UO_1432 (O_1432,N_48389,N_49391);
or UO_1433 (O_1433,N_49623,N_49134);
xnor UO_1434 (O_1434,N_49430,N_49965);
nand UO_1435 (O_1435,N_49330,N_49525);
xnor UO_1436 (O_1436,N_48909,N_49005);
nand UO_1437 (O_1437,N_48318,N_48633);
and UO_1438 (O_1438,N_49449,N_48578);
or UO_1439 (O_1439,N_49213,N_48229);
or UO_1440 (O_1440,N_49461,N_49955);
and UO_1441 (O_1441,N_49310,N_49100);
nor UO_1442 (O_1442,N_49520,N_49556);
and UO_1443 (O_1443,N_48498,N_48494);
nor UO_1444 (O_1444,N_48981,N_48650);
or UO_1445 (O_1445,N_48990,N_48004);
nor UO_1446 (O_1446,N_48845,N_48383);
or UO_1447 (O_1447,N_48494,N_48350);
or UO_1448 (O_1448,N_49307,N_48851);
or UO_1449 (O_1449,N_49466,N_49018);
xor UO_1450 (O_1450,N_49638,N_49396);
nand UO_1451 (O_1451,N_48190,N_49546);
nor UO_1452 (O_1452,N_49666,N_48002);
xnor UO_1453 (O_1453,N_49503,N_49012);
nor UO_1454 (O_1454,N_49951,N_48847);
nor UO_1455 (O_1455,N_48511,N_49130);
nand UO_1456 (O_1456,N_48478,N_48547);
nor UO_1457 (O_1457,N_49880,N_49470);
or UO_1458 (O_1458,N_49195,N_49677);
or UO_1459 (O_1459,N_49628,N_48274);
xnor UO_1460 (O_1460,N_48242,N_49709);
xnor UO_1461 (O_1461,N_48477,N_49682);
or UO_1462 (O_1462,N_48180,N_48529);
nor UO_1463 (O_1463,N_49997,N_48570);
nand UO_1464 (O_1464,N_49306,N_48963);
or UO_1465 (O_1465,N_49348,N_49409);
xor UO_1466 (O_1466,N_48366,N_48653);
nor UO_1467 (O_1467,N_49626,N_49130);
or UO_1468 (O_1468,N_48711,N_48427);
xnor UO_1469 (O_1469,N_48411,N_49980);
or UO_1470 (O_1470,N_49026,N_49293);
and UO_1471 (O_1471,N_48457,N_49690);
or UO_1472 (O_1472,N_48274,N_49208);
nand UO_1473 (O_1473,N_49028,N_48832);
nor UO_1474 (O_1474,N_49953,N_48309);
nor UO_1475 (O_1475,N_49283,N_48664);
nor UO_1476 (O_1476,N_48085,N_49966);
or UO_1477 (O_1477,N_49208,N_48781);
or UO_1478 (O_1478,N_48315,N_48357);
nor UO_1479 (O_1479,N_48768,N_49023);
nand UO_1480 (O_1480,N_48877,N_48447);
or UO_1481 (O_1481,N_48116,N_48746);
nand UO_1482 (O_1482,N_48179,N_48683);
and UO_1483 (O_1483,N_48807,N_48595);
xnor UO_1484 (O_1484,N_49811,N_48605);
nand UO_1485 (O_1485,N_48444,N_48438);
or UO_1486 (O_1486,N_48031,N_49792);
and UO_1487 (O_1487,N_49552,N_48680);
or UO_1488 (O_1488,N_48194,N_49530);
or UO_1489 (O_1489,N_49286,N_49630);
or UO_1490 (O_1490,N_49840,N_48251);
nand UO_1491 (O_1491,N_48532,N_49244);
and UO_1492 (O_1492,N_49746,N_49320);
nor UO_1493 (O_1493,N_48279,N_49556);
xnor UO_1494 (O_1494,N_49892,N_49908);
and UO_1495 (O_1495,N_48740,N_49256);
or UO_1496 (O_1496,N_49413,N_48703);
or UO_1497 (O_1497,N_49620,N_48159);
nand UO_1498 (O_1498,N_49707,N_49129);
or UO_1499 (O_1499,N_48896,N_48149);
or UO_1500 (O_1500,N_49591,N_49269);
nor UO_1501 (O_1501,N_49290,N_48395);
nand UO_1502 (O_1502,N_48171,N_48916);
xor UO_1503 (O_1503,N_48015,N_49373);
and UO_1504 (O_1504,N_48336,N_49775);
and UO_1505 (O_1505,N_49953,N_48999);
or UO_1506 (O_1506,N_49743,N_48558);
or UO_1507 (O_1507,N_49654,N_48227);
nand UO_1508 (O_1508,N_49915,N_48887);
or UO_1509 (O_1509,N_49315,N_48981);
nand UO_1510 (O_1510,N_49254,N_49476);
nor UO_1511 (O_1511,N_49081,N_49933);
xor UO_1512 (O_1512,N_49350,N_49495);
nand UO_1513 (O_1513,N_49867,N_49736);
or UO_1514 (O_1514,N_49717,N_49220);
nor UO_1515 (O_1515,N_49676,N_49060);
nand UO_1516 (O_1516,N_49911,N_48363);
xnor UO_1517 (O_1517,N_48723,N_49517);
and UO_1518 (O_1518,N_48750,N_48425);
xor UO_1519 (O_1519,N_48562,N_48778);
nor UO_1520 (O_1520,N_49021,N_49152);
xor UO_1521 (O_1521,N_49496,N_48037);
and UO_1522 (O_1522,N_49197,N_49007);
xnor UO_1523 (O_1523,N_49794,N_49965);
or UO_1524 (O_1524,N_48111,N_48900);
nor UO_1525 (O_1525,N_49713,N_49545);
or UO_1526 (O_1526,N_49050,N_48187);
xnor UO_1527 (O_1527,N_48906,N_48644);
xnor UO_1528 (O_1528,N_48897,N_48401);
and UO_1529 (O_1529,N_49415,N_49130);
nor UO_1530 (O_1530,N_49053,N_48926);
nand UO_1531 (O_1531,N_48370,N_48984);
nor UO_1532 (O_1532,N_48609,N_49915);
or UO_1533 (O_1533,N_48997,N_48677);
nand UO_1534 (O_1534,N_49124,N_49242);
xnor UO_1535 (O_1535,N_49554,N_48323);
nand UO_1536 (O_1536,N_49766,N_48090);
xnor UO_1537 (O_1537,N_48308,N_48190);
xor UO_1538 (O_1538,N_48933,N_48034);
and UO_1539 (O_1539,N_48117,N_48811);
or UO_1540 (O_1540,N_49142,N_49140);
nand UO_1541 (O_1541,N_49853,N_49700);
nor UO_1542 (O_1542,N_49006,N_48808);
and UO_1543 (O_1543,N_48322,N_48585);
nand UO_1544 (O_1544,N_48729,N_49400);
nor UO_1545 (O_1545,N_48016,N_49108);
nand UO_1546 (O_1546,N_49516,N_48339);
and UO_1547 (O_1547,N_49867,N_48205);
nand UO_1548 (O_1548,N_48854,N_49495);
and UO_1549 (O_1549,N_48846,N_49649);
or UO_1550 (O_1550,N_49676,N_48099);
or UO_1551 (O_1551,N_48864,N_48570);
or UO_1552 (O_1552,N_49625,N_48429);
nor UO_1553 (O_1553,N_48136,N_49784);
or UO_1554 (O_1554,N_49900,N_48644);
nor UO_1555 (O_1555,N_49923,N_49805);
nor UO_1556 (O_1556,N_49527,N_48996);
xnor UO_1557 (O_1557,N_49370,N_48904);
xnor UO_1558 (O_1558,N_49714,N_49327);
nand UO_1559 (O_1559,N_49733,N_49393);
and UO_1560 (O_1560,N_48333,N_49735);
and UO_1561 (O_1561,N_48909,N_49909);
or UO_1562 (O_1562,N_48274,N_48206);
or UO_1563 (O_1563,N_49271,N_49924);
nand UO_1564 (O_1564,N_48778,N_48556);
xnor UO_1565 (O_1565,N_49778,N_49997);
and UO_1566 (O_1566,N_48205,N_49048);
or UO_1567 (O_1567,N_48418,N_48484);
or UO_1568 (O_1568,N_48090,N_49344);
and UO_1569 (O_1569,N_48689,N_48677);
xnor UO_1570 (O_1570,N_48538,N_49982);
nor UO_1571 (O_1571,N_48820,N_49718);
or UO_1572 (O_1572,N_48283,N_49414);
or UO_1573 (O_1573,N_48171,N_49870);
xor UO_1574 (O_1574,N_49702,N_48552);
nand UO_1575 (O_1575,N_49161,N_49405);
nor UO_1576 (O_1576,N_49672,N_49358);
or UO_1577 (O_1577,N_48462,N_49511);
xnor UO_1578 (O_1578,N_49594,N_49208);
xor UO_1579 (O_1579,N_49427,N_48290);
nand UO_1580 (O_1580,N_48602,N_49372);
nor UO_1581 (O_1581,N_49479,N_48806);
xnor UO_1582 (O_1582,N_48939,N_48997);
nand UO_1583 (O_1583,N_49342,N_49798);
or UO_1584 (O_1584,N_49920,N_49878);
nand UO_1585 (O_1585,N_48928,N_49886);
xnor UO_1586 (O_1586,N_48865,N_48713);
nand UO_1587 (O_1587,N_49908,N_49388);
and UO_1588 (O_1588,N_48711,N_49250);
and UO_1589 (O_1589,N_48998,N_48058);
and UO_1590 (O_1590,N_48699,N_49600);
nand UO_1591 (O_1591,N_49082,N_48241);
xnor UO_1592 (O_1592,N_48811,N_49387);
xor UO_1593 (O_1593,N_48179,N_48035);
or UO_1594 (O_1594,N_48193,N_48293);
xor UO_1595 (O_1595,N_48043,N_49594);
and UO_1596 (O_1596,N_48800,N_49398);
nor UO_1597 (O_1597,N_48637,N_49329);
nand UO_1598 (O_1598,N_49410,N_48033);
nor UO_1599 (O_1599,N_48340,N_49144);
or UO_1600 (O_1600,N_48977,N_49130);
or UO_1601 (O_1601,N_49001,N_48558);
xnor UO_1602 (O_1602,N_49250,N_48400);
and UO_1603 (O_1603,N_48895,N_48096);
nor UO_1604 (O_1604,N_48878,N_48080);
xor UO_1605 (O_1605,N_48686,N_49050);
or UO_1606 (O_1606,N_48600,N_48707);
nand UO_1607 (O_1607,N_49347,N_49470);
or UO_1608 (O_1608,N_49743,N_49488);
nand UO_1609 (O_1609,N_49299,N_49767);
nor UO_1610 (O_1610,N_49844,N_49204);
xor UO_1611 (O_1611,N_48013,N_48789);
nand UO_1612 (O_1612,N_48755,N_49950);
and UO_1613 (O_1613,N_48423,N_48637);
or UO_1614 (O_1614,N_48758,N_48723);
xor UO_1615 (O_1615,N_49473,N_48120);
or UO_1616 (O_1616,N_49823,N_48364);
nor UO_1617 (O_1617,N_48118,N_48472);
and UO_1618 (O_1618,N_48732,N_48898);
or UO_1619 (O_1619,N_48294,N_48015);
nor UO_1620 (O_1620,N_49861,N_48336);
xor UO_1621 (O_1621,N_49098,N_48782);
and UO_1622 (O_1622,N_49828,N_49440);
nand UO_1623 (O_1623,N_49730,N_48052);
and UO_1624 (O_1624,N_48675,N_49687);
xor UO_1625 (O_1625,N_49097,N_49424);
nand UO_1626 (O_1626,N_48518,N_49564);
or UO_1627 (O_1627,N_49759,N_48611);
or UO_1628 (O_1628,N_48731,N_49394);
xnor UO_1629 (O_1629,N_49095,N_48865);
or UO_1630 (O_1630,N_48412,N_48067);
nand UO_1631 (O_1631,N_48358,N_48562);
xnor UO_1632 (O_1632,N_48050,N_49123);
xor UO_1633 (O_1633,N_48099,N_49667);
or UO_1634 (O_1634,N_48623,N_48634);
and UO_1635 (O_1635,N_48430,N_48475);
and UO_1636 (O_1636,N_49005,N_49314);
nand UO_1637 (O_1637,N_48486,N_49408);
or UO_1638 (O_1638,N_48830,N_49413);
and UO_1639 (O_1639,N_48656,N_49777);
nand UO_1640 (O_1640,N_49236,N_49195);
nand UO_1641 (O_1641,N_49919,N_48752);
and UO_1642 (O_1642,N_49938,N_48099);
nor UO_1643 (O_1643,N_48954,N_48956);
nand UO_1644 (O_1644,N_48999,N_49486);
nor UO_1645 (O_1645,N_48435,N_49850);
xor UO_1646 (O_1646,N_49770,N_49637);
and UO_1647 (O_1647,N_48115,N_48670);
and UO_1648 (O_1648,N_48010,N_48160);
or UO_1649 (O_1649,N_48222,N_49126);
or UO_1650 (O_1650,N_49403,N_48801);
xnor UO_1651 (O_1651,N_48041,N_49709);
and UO_1652 (O_1652,N_48596,N_49965);
nor UO_1653 (O_1653,N_48144,N_49086);
nor UO_1654 (O_1654,N_48330,N_49889);
nand UO_1655 (O_1655,N_48615,N_48346);
and UO_1656 (O_1656,N_49230,N_49080);
nand UO_1657 (O_1657,N_48662,N_48231);
and UO_1658 (O_1658,N_48998,N_49244);
xnor UO_1659 (O_1659,N_49648,N_49281);
or UO_1660 (O_1660,N_48786,N_48164);
or UO_1661 (O_1661,N_49525,N_48234);
or UO_1662 (O_1662,N_48779,N_49956);
xor UO_1663 (O_1663,N_48599,N_49985);
nor UO_1664 (O_1664,N_49155,N_49359);
nor UO_1665 (O_1665,N_48631,N_48346);
xnor UO_1666 (O_1666,N_48604,N_48774);
nand UO_1667 (O_1667,N_48277,N_48547);
and UO_1668 (O_1668,N_48578,N_48349);
or UO_1669 (O_1669,N_48947,N_49068);
or UO_1670 (O_1670,N_49953,N_49112);
and UO_1671 (O_1671,N_48868,N_48237);
xor UO_1672 (O_1672,N_49287,N_48583);
nor UO_1673 (O_1673,N_49049,N_48981);
xnor UO_1674 (O_1674,N_49762,N_49099);
xor UO_1675 (O_1675,N_48761,N_48582);
and UO_1676 (O_1676,N_49800,N_49151);
and UO_1677 (O_1677,N_49700,N_48937);
xor UO_1678 (O_1678,N_49614,N_48151);
xor UO_1679 (O_1679,N_48928,N_48577);
and UO_1680 (O_1680,N_48921,N_48928);
xor UO_1681 (O_1681,N_48384,N_48591);
and UO_1682 (O_1682,N_49638,N_49210);
and UO_1683 (O_1683,N_49226,N_48948);
xor UO_1684 (O_1684,N_48996,N_48579);
nand UO_1685 (O_1685,N_48670,N_48214);
or UO_1686 (O_1686,N_49604,N_48043);
nand UO_1687 (O_1687,N_48595,N_48790);
or UO_1688 (O_1688,N_49212,N_49084);
nand UO_1689 (O_1689,N_49702,N_48305);
xor UO_1690 (O_1690,N_49182,N_49370);
nand UO_1691 (O_1691,N_49845,N_48460);
and UO_1692 (O_1692,N_48229,N_49171);
nand UO_1693 (O_1693,N_49077,N_49985);
and UO_1694 (O_1694,N_48598,N_49194);
and UO_1695 (O_1695,N_49091,N_49410);
xor UO_1696 (O_1696,N_49031,N_49273);
or UO_1697 (O_1697,N_48079,N_49010);
xor UO_1698 (O_1698,N_48933,N_48636);
nand UO_1699 (O_1699,N_48680,N_49878);
and UO_1700 (O_1700,N_49589,N_49177);
or UO_1701 (O_1701,N_48892,N_49231);
nor UO_1702 (O_1702,N_49611,N_49183);
nand UO_1703 (O_1703,N_49012,N_49790);
xnor UO_1704 (O_1704,N_48429,N_49718);
and UO_1705 (O_1705,N_49281,N_48374);
or UO_1706 (O_1706,N_48042,N_49276);
and UO_1707 (O_1707,N_49684,N_48175);
nand UO_1708 (O_1708,N_48655,N_49191);
nor UO_1709 (O_1709,N_48382,N_49714);
and UO_1710 (O_1710,N_48657,N_49409);
xor UO_1711 (O_1711,N_48646,N_48809);
xor UO_1712 (O_1712,N_48741,N_48411);
nand UO_1713 (O_1713,N_48306,N_48576);
xor UO_1714 (O_1714,N_49384,N_49680);
and UO_1715 (O_1715,N_49835,N_49023);
xnor UO_1716 (O_1716,N_48013,N_48281);
nor UO_1717 (O_1717,N_49206,N_49048);
nand UO_1718 (O_1718,N_48110,N_49071);
or UO_1719 (O_1719,N_49865,N_49137);
nand UO_1720 (O_1720,N_48505,N_48278);
nor UO_1721 (O_1721,N_49573,N_49643);
xnor UO_1722 (O_1722,N_48403,N_48668);
nor UO_1723 (O_1723,N_48120,N_49213);
nor UO_1724 (O_1724,N_49934,N_48050);
xnor UO_1725 (O_1725,N_49130,N_48849);
nand UO_1726 (O_1726,N_48215,N_49744);
or UO_1727 (O_1727,N_48204,N_48506);
nor UO_1728 (O_1728,N_49365,N_48941);
nand UO_1729 (O_1729,N_49051,N_48113);
or UO_1730 (O_1730,N_48759,N_49811);
nand UO_1731 (O_1731,N_48918,N_48855);
or UO_1732 (O_1732,N_48779,N_49196);
nand UO_1733 (O_1733,N_48140,N_48148);
nor UO_1734 (O_1734,N_48705,N_49413);
xnor UO_1735 (O_1735,N_48748,N_48708);
or UO_1736 (O_1736,N_49063,N_49424);
nor UO_1737 (O_1737,N_48404,N_48499);
nand UO_1738 (O_1738,N_48008,N_48181);
nand UO_1739 (O_1739,N_49086,N_49501);
or UO_1740 (O_1740,N_49293,N_49088);
or UO_1741 (O_1741,N_49664,N_48207);
xnor UO_1742 (O_1742,N_49406,N_49404);
nand UO_1743 (O_1743,N_48700,N_49144);
nand UO_1744 (O_1744,N_48659,N_48014);
or UO_1745 (O_1745,N_48306,N_49734);
and UO_1746 (O_1746,N_49604,N_49851);
and UO_1747 (O_1747,N_48699,N_48423);
xor UO_1748 (O_1748,N_49634,N_48142);
nand UO_1749 (O_1749,N_48522,N_48713);
or UO_1750 (O_1750,N_49580,N_48338);
xor UO_1751 (O_1751,N_48837,N_48784);
and UO_1752 (O_1752,N_48915,N_49980);
xor UO_1753 (O_1753,N_48527,N_48138);
nor UO_1754 (O_1754,N_49826,N_48952);
xnor UO_1755 (O_1755,N_48950,N_49602);
xnor UO_1756 (O_1756,N_48442,N_49489);
nand UO_1757 (O_1757,N_48706,N_49921);
or UO_1758 (O_1758,N_48675,N_48907);
nor UO_1759 (O_1759,N_48360,N_48230);
xnor UO_1760 (O_1760,N_48474,N_49433);
and UO_1761 (O_1761,N_49890,N_49033);
nor UO_1762 (O_1762,N_48894,N_48508);
nand UO_1763 (O_1763,N_48259,N_48986);
and UO_1764 (O_1764,N_49238,N_49771);
or UO_1765 (O_1765,N_49411,N_49967);
and UO_1766 (O_1766,N_49643,N_48283);
nand UO_1767 (O_1767,N_48680,N_48758);
and UO_1768 (O_1768,N_49312,N_49168);
and UO_1769 (O_1769,N_49750,N_48867);
nand UO_1770 (O_1770,N_49073,N_48015);
nor UO_1771 (O_1771,N_49754,N_48840);
or UO_1772 (O_1772,N_48342,N_48735);
or UO_1773 (O_1773,N_48583,N_48445);
nor UO_1774 (O_1774,N_49473,N_48998);
xor UO_1775 (O_1775,N_48807,N_48312);
xor UO_1776 (O_1776,N_48310,N_49840);
nor UO_1777 (O_1777,N_48495,N_48355);
or UO_1778 (O_1778,N_48343,N_48550);
nor UO_1779 (O_1779,N_48190,N_48091);
nand UO_1780 (O_1780,N_49622,N_48916);
xor UO_1781 (O_1781,N_49261,N_48072);
and UO_1782 (O_1782,N_49193,N_49379);
nor UO_1783 (O_1783,N_49731,N_49883);
xor UO_1784 (O_1784,N_49211,N_49251);
nor UO_1785 (O_1785,N_49381,N_49949);
nand UO_1786 (O_1786,N_48881,N_48992);
xor UO_1787 (O_1787,N_49923,N_48544);
nand UO_1788 (O_1788,N_48936,N_49583);
xor UO_1789 (O_1789,N_49110,N_48319);
or UO_1790 (O_1790,N_49987,N_48075);
xnor UO_1791 (O_1791,N_49327,N_48153);
or UO_1792 (O_1792,N_49353,N_48595);
nor UO_1793 (O_1793,N_48103,N_48419);
nor UO_1794 (O_1794,N_49302,N_49366);
or UO_1795 (O_1795,N_49856,N_49768);
and UO_1796 (O_1796,N_48657,N_48925);
nor UO_1797 (O_1797,N_48537,N_48778);
and UO_1798 (O_1798,N_49827,N_49157);
or UO_1799 (O_1799,N_48547,N_48168);
nor UO_1800 (O_1800,N_49455,N_49696);
or UO_1801 (O_1801,N_48335,N_49766);
and UO_1802 (O_1802,N_49497,N_49459);
nor UO_1803 (O_1803,N_48643,N_48524);
nand UO_1804 (O_1804,N_49164,N_48128);
or UO_1805 (O_1805,N_48839,N_48063);
nand UO_1806 (O_1806,N_49202,N_49520);
and UO_1807 (O_1807,N_49964,N_48282);
xnor UO_1808 (O_1808,N_49809,N_48942);
nand UO_1809 (O_1809,N_48011,N_48994);
nand UO_1810 (O_1810,N_48671,N_49892);
and UO_1811 (O_1811,N_48710,N_48630);
or UO_1812 (O_1812,N_48005,N_48685);
or UO_1813 (O_1813,N_49844,N_49748);
nor UO_1814 (O_1814,N_49117,N_48831);
or UO_1815 (O_1815,N_49651,N_48713);
or UO_1816 (O_1816,N_48734,N_49579);
or UO_1817 (O_1817,N_49014,N_49705);
and UO_1818 (O_1818,N_48700,N_49496);
nand UO_1819 (O_1819,N_48832,N_48656);
xor UO_1820 (O_1820,N_48118,N_49600);
nand UO_1821 (O_1821,N_48316,N_48481);
or UO_1822 (O_1822,N_48845,N_48948);
or UO_1823 (O_1823,N_49180,N_48019);
nand UO_1824 (O_1824,N_49076,N_48466);
or UO_1825 (O_1825,N_48567,N_49184);
nor UO_1826 (O_1826,N_49416,N_48088);
or UO_1827 (O_1827,N_49530,N_48665);
nand UO_1828 (O_1828,N_48116,N_49326);
xnor UO_1829 (O_1829,N_49603,N_49180);
xnor UO_1830 (O_1830,N_48915,N_48850);
or UO_1831 (O_1831,N_49320,N_48575);
xnor UO_1832 (O_1832,N_49075,N_49421);
and UO_1833 (O_1833,N_49920,N_49701);
nor UO_1834 (O_1834,N_48382,N_48374);
nor UO_1835 (O_1835,N_48780,N_48526);
or UO_1836 (O_1836,N_48838,N_48280);
xor UO_1837 (O_1837,N_48741,N_48149);
xor UO_1838 (O_1838,N_49613,N_49926);
and UO_1839 (O_1839,N_49481,N_49478);
nand UO_1840 (O_1840,N_48413,N_48328);
nor UO_1841 (O_1841,N_48774,N_48858);
nand UO_1842 (O_1842,N_48583,N_49776);
nor UO_1843 (O_1843,N_48570,N_48260);
or UO_1844 (O_1844,N_48952,N_48181);
nor UO_1845 (O_1845,N_49344,N_49938);
nor UO_1846 (O_1846,N_49082,N_48628);
nor UO_1847 (O_1847,N_48529,N_48286);
and UO_1848 (O_1848,N_48822,N_48276);
nor UO_1849 (O_1849,N_48604,N_48711);
xnor UO_1850 (O_1850,N_48908,N_48394);
xor UO_1851 (O_1851,N_48399,N_48311);
nor UO_1852 (O_1852,N_49755,N_49805);
xor UO_1853 (O_1853,N_48196,N_49468);
nor UO_1854 (O_1854,N_48831,N_49501);
and UO_1855 (O_1855,N_49856,N_48391);
nor UO_1856 (O_1856,N_48472,N_49967);
nor UO_1857 (O_1857,N_49856,N_49393);
and UO_1858 (O_1858,N_49138,N_48446);
xnor UO_1859 (O_1859,N_48192,N_49349);
xnor UO_1860 (O_1860,N_49683,N_48556);
nor UO_1861 (O_1861,N_48914,N_48361);
and UO_1862 (O_1862,N_48002,N_49775);
or UO_1863 (O_1863,N_49637,N_49167);
nor UO_1864 (O_1864,N_49515,N_49449);
and UO_1865 (O_1865,N_49190,N_48750);
or UO_1866 (O_1866,N_48818,N_48981);
or UO_1867 (O_1867,N_48900,N_49432);
and UO_1868 (O_1868,N_48439,N_49896);
nand UO_1869 (O_1869,N_48965,N_48202);
or UO_1870 (O_1870,N_48413,N_49259);
or UO_1871 (O_1871,N_49875,N_48233);
nor UO_1872 (O_1872,N_48794,N_49766);
nand UO_1873 (O_1873,N_48374,N_48570);
nor UO_1874 (O_1874,N_49359,N_49512);
and UO_1875 (O_1875,N_49059,N_48746);
xor UO_1876 (O_1876,N_49695,N_49823);
xor UO_1877 (O_1877,N_49547,N_49017);
or UO_1878 (O_1878,N_49022,N_48254);
and UO_1879 (O_1879,N_49014,N_48142);
and UO_1880 (O_1880,N_49846,N_48374);
xor UO_1881 (O_1881,N_48872,N_49110);
or UO_1882 (O_1882,N_48603,N_49695);
nor UO_1883 (O_1883,N_48271,N_48777);
or UO_1884 (O_1884,N_49475,N_49052);
or UO_1885 (O_1885,N_49549,N_49822);
or UO_1886 (O_1886,N_49453,N_48142);
and UO_1887 (O_1887,N_48097,N_48627);
or UO_1888 (O_1888,N_48807,N_48903);
xnor UO_1889 (O_1889,N_49752,N_48534);
nor UO_1890 (O_1890,N_48567,N_49902);
nand UO_1891 (O_1891,N_48473,N_49877);
xnor UO_1892 (O_1892,N_49720,N_49669);
xor UO_1893 (O_1893,N_48248,N_48599);
and UO_1894 (O_1894,N_48135,N_48620);
and UO_1895 (O_1895,N_49193,N_49156);
and UO_1896 (O_1896,N_49587,N_49225);
or UO_1897 (O_1897,N_49148,N_48370);
xnor UO_1898 (O_1898,N_48570,N_49994);
xnor UO_1899 (O_1899,N_49750,N_49606);
and UO_1900 (O_1900,N_49139,N_49357);
or UO_1901 (O_1901,N_48761,N_48361);
and UO_1902 (O_1902,N_49786,N_49313);
and UO_1903 (O_1903,N_49336,N_48899);
xor UO_1904 (O_1904,N_49782,N_48270);
nor UO_1905 (O_1905,N_48291,N_48222);
nand UO_1906 (O_1906,N_49692,N_49303);
nor UO_1907 (O_1907,N_49632,N_48337);
xor UO_1908 (O_1908,N_48849,N_49487);
or UO_1909 (O_1909,N_48532,N_49341);
or UO_1910 (O_1910,N_49414,N_49143);
xor UO_1911 (O_1911,N_49231,N_48206);
and UO_1912 (O_1912,N_49522,N_48802);
and UO_1913 (O_1913,N_49199,N_49110);
or UO_1914 (O_1914,N_48544,N_49215);
or UO_1915 (O_1915,N_48182,N_49690);
xor UO_1916 (O_1916,N_48320,N_48154);
nor UO_1917 (O_1917,N_49686,N_48917);
and UO_1918 (O_1918,N_49180,N_49794);
nor UO_1919 (O_1919,N_48540,N_48907);
and UO_1920 (O_1920,N_48216,N_49707);
nand UO_1921 (O_1921,N_49464,N_48090);
or UO_1922 (O_1922,N_49881,N_48974);
nand UO_1923 (O_1923,N_48430,N_49917);
nor UO_1924 (O_1924,N_48190,N_48412);
xor UO_1925 (O_1925,N_49308,N_48355);
or UO_1926 (O_1926,N_49287,N_49895);
nand UO_1927 (O_1927,N_49976,N_49431);
nand UO_1928 (O_1928,N_49190,N_48476);
nand UO_1929 (O_1929,N_49386,N_48436);
xnor UO_1930 (O_1930,N_49637,N_48089);
and UO_1931 (O_1931,N_48759,N_49620);
and UO_1932 (O_1932,N_48898,N_48259);
nor UO_1933 (O_1933,N_48545,N_48736);
or UO_1934 (O_1934,N_48185,N_48992);
xor UO_1935 (O_1935,N_49142,N_49199);
nor UO_1936 (O_1936,N_48697,N_48302);
nor UO_1937 (O_1937,N_48217,N_48872);
and UO_1938 (O_1938,N_48908,N_49204);
and UO_1939 (O_1939,N_48524,N_49667);
and UO_1940 (O_1940,N_48164,N_48779);
nand UO_1941 (O_1941,N_48365,N_48171);
or UO_1942 (O_1942,N_48611,N_48978);
or UO_1943 (O_1943,N_48805,N_49679);
nor UO_1944 (O_1944,N_49648,N_49231);
nand UO_1945 (O_1945,N_49538,N_48144);
or UO_1946 (O_1946,N_49728,N_48903);
or UO_1947 (O_1947,N_49362,N_48577);
and UO_1948 (O_1948,N_48568,N_49028);
nand UO_1949 (O_1949,N_48351,N_49434);
xor UO_1950 (O_1950,N_49982,N_49862);
or UO_1951 (O_1951,N_49828,N_49136);
or UO_1952 (O_1952,N_49405,N_49878);
or UO_1953 (O_1953,N_48626,N_49381);
xnor UO_1954 (O_1954,N_49981,N_48504);
nand UO_1955 (O_1955,N_48280,N_49595);
xor UO_1956 (O_1956,N_49480,N_48487);
nand UO_1957 (O_1957,N_49868,N_48372);
or UO_1958 (O_1958,N_48164,N_48386);
or UO_1959 (O_1959,N_49738,N_49917);
and UO_1960 (O_1960,N_48413,N_48091);
nor UO_1961 (O_1961,N_48943,N_49813);
xnor UO_1962 (O_1962,N_49235,N_49872);
or UO_1963 (O_1963,N_49476,N_48112);
and UO_1964 (O_1964,N_48925,N_48153);
or UO_1965 (O_1965,N_49403,N_48376);
and UO_1966 (O_1966,N_49051,N_48031);
or UO_1967 (O_1967,N_49543,N_48242);
and UO_1968 (O_1968,N_48163,N_48712);
or UO_1969 (O_1969,N_49358,N_48194);
xor UO_1970 (O_1970,N_48448,N_49431);
nand UO_1971 (O_1971,N_49261,N_49600);
and UO_1972 (O_1972,N_49768,N_48604);
and UO_1973 (O_1973,N_49913,N_48216);
nor UO_1974 (O_1974,N_49272,N_48986);
and UO_1975 (O_1975,N_49072,N_48611);
xnor UO_1976 (O_1976,N_48600,N_49695);
or UO_1977 (O_1977,N_49907,N_48944);
and UO_1978 (O_1978,N_48932,N_49787);
and UO_1979 (O_1979,N_49709,N_49497);
nand UO_1980 (O_1980,N_48261,N_48460);
xnor UO_1981 (O_1981,N_48497,N_48166);
nor UO_1982 (O_1982,N_48257,N_48757);
nand UO_1983 (O_1983,N_49851,N_49655);
xor UO_1984 (O_1984,N_49372,N_49890);
nand UO_1985 (O_1985,N_49859,N_49356);
nor UO_1986 (O_1986,N_49971,N_48376);
nand UO_1987 (O_1987,N_48392,N_49342);
nor UO_1988 (O_1988,N_49391,N_49253);
nand UO_1989 (O_1989,N_48182,N_48711);
or UO_1990 (O_1990,N_48864,N_49340);
and UO_1991 (O_1991,N_48298,N_48854);
and UO_1992 (O_1992,N_48659,N_48418);
xor UO_1993 (O_1993,N_48503,N_48791);
xnor UO_1994 (O_1994,N_48695,N_49030);
xor UO_1995 (O_1995,N_49586,N_49577);
and UO_1996 (O_1996,N_48295,N_49452);
and UO_1997 (O_1997,N_48422,N_48160);
nor UO_1998 (O_1998,N_48763,N_48438);
xor UO_1999 (O_1999,N_48668,N_49314);
and UO_2000 (O_2000,N_49183,N_48669);
nand UO_2001 (O_2001,N_49528,N_49883);
xor UO_2002 (O_2002,N_48114,N_49083);
or UO_2003 (O_2003,N_48616,N_48786);
nand UO_2004 (O_2004,N_49034,N_49923);
nor UO_2005 (O_2005,N_49212,N_48484);
nor UO_2006 (O_2006,N_49952,N_49861);
or UO_2007 (O_2007,N_48541,N_48786);
nor UO_2008 (O_2008,N_48635,N_48275);
nand UO_2009 (O_2009,N_49404,N_48497);
and UO_2010 (O_2010,N_48441,N_48197);
or UO_2011 (O_2011,N_49722,N_48403);
nor UO_2012 (O_2012,N_49565,N_48756);
nor UO_2013 (O_2013,N_49819,N_49541);
nor UO_2014 (O_2014,N_49861,N_48748);
nor UO_2015 (O_2015,N_48801,N_49334);
nand UO_2016 (O_2016,N_49708,N_49919);
nand UO_2017 (O_2017,N_49402,N_49908);
nor UO_2018 (O_2018,N_48490,N_48556);
and UO_2019 (O_2019,N_48920,N_48816);
xor UO_2020 (O_2020,N_49131,N_49294);
and UO_2021 (O_2021,N_49507,N_48397);
nor UO_2022 (O_2022,N_48960,N_48376);
nand UO_2023 (O_2023,N_49822,N_48860);
and UO_2024 (O_2024,N_49488,N_48998);
nor UO_2025 (O_2025,N_49396,N_48879);
or UO_2026 (O_2026,N_49000,N_49291);
nor UO_2027 (O_2027,N_49709,N_49349);
or UO_2028 (O_2028,N_48591,N_49421);
and UO_2029 (O_2029,N_48180,N_49627);
xnor UO_2030 (O_2030,N_49252,N_48289);
nor UO_2031 (O_2031,N_48714,N_49785);
nor UO_2032 (O_2032,N_48484,N_49110);
nand UO_2033 (O_2033,N_49714,N_49770);
nand UO_2034 (O_2034,N_49230,N_49122);
and UO_2035 (O_2035,N_49835,N_49433);
xor UO_2036 (O_2036,N_49144,N_49212);
and UO_2037 (O_2037,N_48974,N_49135);
and UO_2038 (O_2038,N_49973,N_49992);
nor UO_2039 (O_2039,N_48800,N_48158);
and UO_2040 (O_2040,N_48994,N_49219);
or UO_2041 (O_2041,N_49967,N_48956);
nand UO_2042 (O_2042,N_48098,N_48820);
nor UO_2043 (O_2043,N_48758,N_49803);
xnor UO_2044 (O_2044,N_49045,N_49091);
and UO_2045 (O_2045,N_48179,N_48028);
or UO_2046 (O_2046,N_48360,N_49369);
or UO_2047 (O_2047,N_48561,N_48787);
or UO_2048 (O_2048,N_48639,N_49167);
xnor UO_2049 (O_2049,N_48125,N_48757);
or UO_2050 (O_2050,N_48725,N_49751);
or UO_2051 (O_2051,N_48640,N_49421);
xor UO_2052 (O_2052,N_48946,N_49391);
nor UO_2053 (O_2053,N_49715,N_49531);
nor UO_2054 (O_2054,N_48862,N_49043);
nand UO_2055 (O_2055,N_48293,N_48695);
nand UO_2056 (O_2056,N_49673,N_49408);
nor UO_2057 (O_2057,N_48574,N_48528);
nand UO_2058 (O_2058,N_49820,N_49563);
nor UO_2059 (O_2059,N_48436,N_48085);
nor UO_2060 (O_2060,N_49421,N_49230);
nor UO_2061 (O_2061,N_49669,N_49128);
nor UO_2062 (O_2062,N_49498,N_49526);
nand UO_2063 (O_2063,N_48633,N_49694);
and UO_2064 (O_2064,N_49235,N_48746);
and UO_2065 (O_2065,N_48121,N_49747);
or UO_2066 (O_2066,N_48358,N_48898);
nand UO_2067 (O_2067,N_49156,N_48736);
nand UO_2068 (O_2068,N_48288,N_49676);
or UO_2069 (O_2069,N_49799,N_48533);
and UO_2070 (O_2070,N_49531,N_48629);
or UO_2071 (O_2071,N_48212,N_49747);
or UO_2072 (O_2072,N_48019,N_49036);
nand UO_2073 (O_2073,N_48933,N_49068);
nor UO_2074 (O_2074,N_49898,N_49799);
or UO_2075 (O_2075,N_48277,N_49565);
and UO_2076 (O_2076,N_49203,N_49196);
or UO_2077 (O_2077,N_49745,N_48406);
nor UO_2078 (O_2078,N_49071,N_49372);
nor UO_2079 (O_2079,N_49550,N_48956);
nand UO_2080 (O_2080,N_48102,N_48579);
nand UO_2081 (O_2081,N_48020,N_49728);
and UO_2082 (O_2082,N_49404,N_48199);
and UO_2083 (O_2083,N_48431,N_48066);
xnor UO_2084 (O_2084,N_48409,N_49099);
or UO_2085 (O_2085,N_49558,N_48377);
or UO_2086 (O_2086,N_49058,N_49709);
and UO_2087 (O_2087,N_48907,N_48910);
and UO_2088 (O_2088,N_49944,N_49899);
nand UO_2089 (O_2089,N_49601,N_48944);
nor UO_2090 (O_2090,N_49852,N_48594);
or UO_2091 (O_2091,N_48647,N_48553);
or UO_2092 (O_2092,N_48309,N_48782);
and UO_2093 (O_2093,N_49224,N_48213);
or UO_2094 (O_2094,N_48725,N_49248);
nand UO_2095 (O_2095,N_48198,N_49735);
or UO_2096 (O_2096,N_49530,N_48704);
and UO_2097 (O_2097,N_49934,N_49546);
and UO_2098 (O_2098,N_49086,N_48209);
nand UO_2099 (O_2099,N_48622,N_49799);
and UO_2100 (O_2100,N_49567,N_49275);
nand UO_2101 (O_2101,N_49875,N_48279);
nand UO_2102 (O_2102,N_49463,N_49053);
nor UO_2103 (O_2103,N_49783,N_49364);
nand UO_2104 (O_2104,N_49131,N_48864);
and UO_2105 (O_2105,N_48370,N_49138);
nor UO_2106 (O_2106,N_49573,N_49357);
nand UO_2107 (O_2107,N_48166,N_49333);
nand UO_2108 (O_2108,N_48599,N_49009);
xor UO_2109 (O_2109,N_49515,N_48782);
nor UO_2110 (O_2110,N_48168,N_48535);
or UO_2111 (O_2111,N_49509,N_48020);
nor UO_2112 (O_2112,N_48154,N_49575);
and UO_2113 (O_2113,N_49553,N_49700);
xor UO_2114 (O_2114,N_49670,N_48213);
nand UO_2115 (O_2115,N_49596,N_49313);
xnor UO_2116 (O_2116,N_49505,N_49027);
or UO_2117 (O_2117,N_49736,N_49904);
nand UO_2118 (O_2118,N_49140,N_49272);
or UO_2119 (O_2119,N_48596,N_48716);
xnor UO_2120 (O_2120,N_49182,N_49204);
nand UO_2121 (O_2121,N_48861,N_49614);
nand UO_2122 (O_2122,N_48197,N_49391);
and UO_2123 (O_2123,N_48723,N_49167);
and UO_2124 (O_2124,N_48545,N_49542);
or UO_2125 (O_2125,N_48521,N_48091);
nand UO_2126 (O_2126,N_48366,N_48843);
and UO_2127 (O_2127,N_49174,N_48549);
nor UO_2128 (O_2128,N_48651,N_49828);
nor UO_2129 (O_2129,N_49438,N_48787);
nand UO_2130 (O_2130,N_48839,N_48348);
nor UO_2131 (O_2131,N_48382,N_49720);
nand UO_2132 (O_2132,N_48370,N_48649);
and UO_2133 (O_2133,N_48824,N_49467);
or UO_2134 (O_2134,N_48329,N_48420);
nor UO_2135 (O_2135,N_49576,N_48939);
nand UO_2136 (O_2136,N_49497,N_48836);
xnor UO_2137 (O_2137,N_48289,N_48684);
nand UO_2138 (O_2138,N_49264,N_49339);
nor UO_2139 (O_2139,N_49791,N_49317);
nand UO_2140 (O_2140,N_49109,N_48754);
or UO_2141 (O_2141,N_49703,N_48654);
nand UO_2142 (O_2142,N_48513,N_48878);
or UO_2143 (O_2143,N_48454,N_48339);
xor UO_2144 (O_2144,N_49323,N_48173);
and UO_2145 (O_2145,N_48970,N_48331);
and UO_2146 (O_2146,N_49585,N_48167);
or UO_2147 (O_2147,N_49904,N_49066);
nor UO_2148 (O_2148,N_49552,N_48577);
and UO_2149 (O_2149,N_48555,N_49088);
or UO_2150 (O_2150,N_48411,N_48906);
and UO_2151 (O_2151,N_49327,N_49141);
nand UO_2152 (O_2152,N_48029,N_49442);
or UO_2153 (O_2153,N_49290,N_48802);
and UO_2154 (O_2154,N_49002,N_49409);
and UO_2155 (O_2155,N_49790,N_48762);
and UO_2156 (O_2156,N_49002,N_48593);
and UO_2157 (O_2157,N_48357,N_48624);
nand UO_2158 (O_2158,N_49335,N_49940);
nor UO_2159 (O_2159,N_48163,N_48741);
nor UO_2160 (O_2160,N_49903,N_48188);
nand UO_2161 (O_2161,N_49630,N_49536);
and UO_2162 (O_2162,N_48213,N_49037);
xnor UO_2163 (O_2163,N_49838,N_48108);
and UO_2164 (O_2164,N_48773,N_48172);
nand UO_2165 (O_2165,N_49359,N_48417);
nand UO_2166 (O_2166,N_49922,N_49342);
or UO_2167 (O_2167,N_49010,N_49264);
nor UO_2168 (O_2168,N_49329,N_48487);
nand UO_2169 (O_2169,N_49375,N_48109);
nand UO_2170 (O_2170,N_49210,N_48275);
nand UO_2171 (O_2171,N_48388,N_48459);
nor UO_2172 (O_2172,N_48813,N_48380);
nand UO_2173 (O_2173,N_48305,N_49760);
nand UO_2174 (O_2174,N_49505,N_48458);
nor UO_2175 (O_2175,N_49860,N_48779);
nor UO_2176 (O_2176,N_49874,N_49528);
and UO_2177 (O_2177,N_48829,N_49152);
xor UO_2178 (O_2178,N_48946,N_48824);
nand UO_2179 (O_2179,N_48188,N_49627);
nand UO_2180 (O_2180,N_48630,N_49360);
nor UO_2181 (O_2181,N_48597,N_48118);
nand UO_2182 (O_2182,N_49808,N_49558);
nor UO_2183 (O_2183,N_49063,N_48588);
and UO_2184 (O_2184,N_48537,N_49192);
nand UO_2185 (O_2185,N_48026,N_48393);
nor UO_2186 (O_2186,N_48090,N_49916);
or UO_2187 (O_2187,N_49931,N_49879);
or UO_2188 (O_2188,N_49658,N_49971);
xor UO_2189 (O_2189,N_48879,N_48996);
nor UO_2190 (O_2190,N_49697,N_49366);
nor UO_2191 (O_2191,N_48254,N_49119);
or UO_2192 (O_2192,N_48125,N_48627);
nand UO_2193 (O_2193,N_49777,N_48068);
or UO_2194 (O_2194,N_48084,N_48976);
nand UO_2195 (O_2195,N_49616,N_49365);
nand UO_2196 (O_2196,N_49576,N_49524);
or UO_2197 (O_2197,N_49531,N_49579);
and UO_2198 (O_2198,N_48201,N_49126);
and UO_2199 (O_2199,N_49998,N_48511);
or UO_2200 (O_2200,N_48273,N_48341);
nand UO_2201 (O_2201,N_48518,N_48059);
nor UO_2202 (O_2202,N_48352,N_48804);
nand UO_2203 (O_2203,N_48277,N_49126);
xor UO_2204 (O_2204,N_48189,N_49719);
and UO_2205 (O_2205,N_49677,N_49620);
or UO_2206 (O_2206,N_49994,N_48965);
xnor UO_2207 (O_2207,N_48448,N_48774);
nand UO_2208 (O_2208,N_48146,N_48815);
and UO_2209 (O_2209,N_48941,N_49648);
nand UO_2210 (O_2210,N_49597,N_49564);
xor UO_2211 (O_2211,N_49274,N_49401);
and UO_2212 (O_2212,N_49281,N_48728);
xnor UO_2213 (O_2213,N_49191,N_49189);
or UO_2214 (O_2214,N_48102,N_48774);
or UO_2215 (O_2215,N_48602,N_48824);
or UO_2216 (O_2216,N_48720,N_48443);
and UO_2217 (O_2217,N_48974,N_49210);
nand UO_2218 (O_2218,N_49616,N_49304);
nor UO_2219 (O_2219,N_49360,N_49104);
and UO_2220 (O_2220,N_49726,N_49508);
nand UO_2221 (O_2221,N_48099,N_49227);
xnor UO_2222 (O_2222,N_48778,N_49112);
or UO_2223 (O_2223,N_48893,N_48357);
xnor UO_2224 (O_2224,N_49616,N_48272);
and UO_2225 (O_2225,N_49220,N_49835);
nand UO_2226 (O_2226,N_48278,N_48011);
nor UO_2227 (O_2227,N_48595,N_49832);
and UO_2228 (O_2228,N_49106,N_49756);
nand UO_2229 (O_2229,N_49962,N_49735);
or UO_2230 (O_2230,N_49645,N_48203);
nand UO_2231 (O_2231,N_48945,N_48232);
nand UO_2232 (O_2232,N_48598,N_48305);
nor UO_2233 (O_2233,N_49893,N_48659);
xor UO_2234 (O_2234,N_49190,N_49944);
nand UO_2235 (O_2235,N_49232,N_49229);
nand UO_2236 (O_2236,N_49517,N_49921);
and UO_2237 (O_2237,N_48179,N_48919);
or UO_2238 (O_2238,N_48622,N_48066);
xnor UO_2239 (O_2239,N_48476,N_49310);
xor UO_2240 (O_2240,N_49176,N_48790);
xnor UO_2241 (O_2241,N_48334,N_48496);
and UO_2242 (O_2242,N_49910,N_49904);
or UO_2243 (O_2243,N_48160,N_49890);
nand UO_2244 (O_2244,N_48853,N_48616);
and UO_2245 (O_2245,N_49881,N_49850);
nor UO_2246 (O_2246,N_49715,N_48380);
nor UO_2247 (O_2247,N_48553,N_48769);
xnor UO_2248 (O_2248,N_48839,N_48952);
and UO_2249 (O_2249,N_49018,N_48830);
or UO_2250 (O_2250,N_48327,N_49547);
xor UO_2251 (O_2251,N_48660,N_49632);
or UO_2252 (O_2252,N_49292,N_48525);
nand UO_2253 (O_2253,N_48716,N_48936);
nand UO_2254 (O_2254,N_48607,N_49104);
and UO_2255 (O_2255,N_49135,N_49634);
xor UO_2256 (O_2256,N_49434,N_48577);
nand UO_2257 (O_2257,N_49396,N_49145);
nand UO_2258 (O_2258,N_49947,N_48052);
or UO_2259 (O_2259,N_48984,N_49272);
or UO_2260 (O_2260,N_48532,N_48242);
or UO_2261 (O_2261,N_49526,N_49804);
and UO_2262 (O_2262,N_49490,N_49994);
nor UO_2263 (O_2263,N_49133,N_48599);
xnor UO_2264 (O_2264,N_49288,N_49652);
nor UO_2265 (O_2265,N_48443,N_49433);
nor UO_2266 (O_2266,N_48017,N_48771);
nand UO_2267 (O_2267,N_49663,N_48679);
nor UO_2268 (O_2268,N_49045,N_49458);
xor UO_2269 (O_2269,N_48399,N_49379);
nor UO_2270 (O_2270,N_48494,N_48571);
xor UO_2271 (O_2271,N_48770,N_49033);
or UO_2272 (O_2272,N_48675,N_48625);
nand UO_2273 (O_2273,N_48073,N_48150);
nor UO_2274 (O_2274,N_48673,N_49143);
or UO_2275 (O_2275,N_49604,N_49219);
xor UO_2276 (O_2276,N_49728,N_49316);
or UO_2277 (O_2277,N_49479,N_48518);
nand UO_2278 (O_2278,N_48383,N_48662);
or UO_2279 (O_2279,N_49307,N_48290);
nand UO_2280 (O_2280,N_48372,N_49166);
nand UO_2281 (O_2281,N_49497,N_48393);
nor UO_2282 (O_2282,N_48471,N_49326);
and UO_2283 (O_2283,N_49194,N_48762);
or UO_2284 (O_2284,N_48635,N_49946);
and UO_2285 (O_2285,N_49508,N_49598);
nand UO_2286 (O_2286,N_49657,N_49332);
xnor UO_2287 (O_2287,N_49653,N_48170);
and UO_2288 (O_2288,N_49576,N_49122);
and UO_2289 (O_2289,N_48747,N_48017);
or UO_2290 (O_2290,N_48448,N_49855);
or UO_2291 (O_2291,N_49339,N_49097);
or UO_2292 (O_2292,N_48078,N_49930);
and UO_2293 (O_2293,N_49900,N_48035);
or UO_2294 (O_2294,N_49807,N_48091);
xnor UO_2295 (O_2295,N_49316,N_49101);
nand UO_2296 (O_2296,N_49715,N_48421);
and UO_2297 (O_2297,N_49293,N_48598);
nand UO_2298 (O_2298,N_49594,N_48147);
and UO_2299 (O_2299,N_48591,N_49078);
nand UO_2300 (O_2300,N_48052,N_49553);
or UO_2301 (O_2301,N_48032,N_49832);
and UO_2302 (O_2302,N_49179,N_48195);
nor UO_2303 (O_2303,N_49157,N_49665);
xnor UO_2304 (O_2304,N_49692,N_48485);
or UO_2305 (O_2305,N_49732,N_48446);
nor UO_2306 (O_2306,N_48324,N_49484);
xnor UO_2307 (O_2307,N_48630,N_48355);
nand UO_2308 (O_2308,N_49331,N_49719);
nand UO_2309 (O_2309,N_49368,N_48711);
and UO_2310 (O_2310,N_48257,N_48449);
and UO_2311 (O_2311,N_48219,N_48712);
and UO_2312 (O_2312,N_48350,N_48504);
nand UO_2313 (O_2313,N_48248,N_49315);
and UO_2314 (O_2314,N_49163,N_49288);
nand UO_2315 (O_2315,N_49406,N_48876);
or UO_2316 (O_2316,N_49759,N_48260);
nor UO_2317 (O_2317,N_49221,N_49783);
nor UO_2318 (O_2318,N_48040,N_49594);
or UO_2319 (O_2319,N_48863,N_48044);
and UO_2320 (O_2320,N_49991,N_48495);
and UO_2321 (O_2321,N_48411,N_49475);
xnor UO_2322 (O_2322,N_49704,N_48999);
nor UO_2323 (O_2323,N_49130,N_48033);
nor UO_2324 (O_2324,N_48179,N_49111);
nand UO_2325 (O_2325,N_49705,N_48546);
nand UO_2326 (O_2326,N_48263,N_48288);
nor UO_2327 (O_2327,N_48266,N_48730);
nand UO_2328 (O_2328,N_49116,N_49512);
xor UO_2329 (O_2329,N_49612,N_48845);
nand UO_2330 (O_2330,N_48581,N_49974);
and UO_2331 (O_2331,N_49721,N_49583);
nor UO_2332 (O_2332,N_48103,N_48715);
nor UO_2333 (O_2333,N_48171,N_49416);
and UO_2334 (O_2334,N_48384,N_48726);
and UO_2335 (O_2335,N_48497,N_48627);
xor UO_2336 (O_2336,N_49532,N_48039);
and UO_2337 (O_2337,N_49813,N_49628);
nor UO_2338 (O_2338,N_48499,N_49566);
and UO_2339 (O_2339,N_49901,N_49605);
and UO_2340 (O_2340,N_48680,N_48205);
xnor UO_2341 (O_2341,N_49603,N_49868);
xor UO_2342 (O_2342,N_49214,N_48376);
and UO_2343 (O_2343,N_49782,N_48110);
or UO_2344 (O_2344,N_48816,N_48349);
xnor UO_2345 (O_2345,N_48612,N_48903);
nor UO_2346 (O_2346,N_49727,N_48777);
nand UO_2347 (O_2347,N_49311,N_48818);
xor UO_2348 (O_2348,N_49597,N_48803);
or UO_2349 (O_2349,N_49431,N_48014);
nor UO_2350 (O_2350,N_49942,N_49277);
nor UO_2351 (O_2351,N_49068,N_48354);
xor UO_2352 (O_2352,N_48780,N_48737);
or UO_2353 (O_2353,N_49476,N_49160);
and UO_2354 (O_2354,N_48132,N_48615);
and UO_2355 (O_2355,N_49083,N_48138);
or UO_2356 (O_2356,N_48666,N_49040);
nand UO_2357 (O_2357,N_49878,N_48327);
nand UO_2358 (O_2358,N_48596,N_49464);
xnor UO_2359 (O_2359,N_49029,N_48502);
and UO_2360 (O_2360,N_48039,N_48229);
and UO_2361 (O_2361,N_49615,N_49361);
or UO_2362 (O_2362,N_48843,N_48303);
nand UO_2363 (O_2363,N_48444,N_49316);
nand UO_2364 (O_2364,N_48037,N_48406);
or UO_2365 (O_2365,N_48553,N_48081);
or UO_2366 (O_2366,N_48522,N_49841);
nor UO_2367 (O_2367,N_49049,N_48800);
nand UO_2368 (O_2368,N_49669,N_48656);
or UO_2369 (O_2369,N_48803,N_49640);
nor UO_2370 (O_2370,N_48103,N_49943);
nor UO_2371 (O_2371,N_48564,N_48625);
and UO_2372 (O_2372,N_49680,N_48829);
and UO_2373 (O_2373,N_49479,N_49733);
nor UO_2374 (O_2374,N_49322,N_48712);
nor UO_2375 (O_2375,N_48250,N_49977);
nand UO_2376 (O_2376,N_48180,N_48079);
nand UO_2377 (O_2377,N_48832,N_49356);
xor UO_2378 (O_2378,N_49390,N_49783);
xnor UO_2379 (O_2379,N_49972,N_48337);
or UO_2380 (O_2380,N_48261,N_48076);
nand UO_2381 (O_2381,N_48269,N_48572);
and UO_2382 (O_2382,N_49017,N_49577);
nor UO_2383 (O_2383,N_48829,N_49644);
xor UO_2384 (O_2384,N_49373,N_49942);
xor UO_2385 (O_2385,N_48780,N_49291);
nand UO_2386 (O_2386,N_48580,N_49736);
xor UO_2387 (O_2387,N_49512,N_48941);
and UO_2388 (O_2388,N_48346,N_48807);
nor UO_2389 (O_2389,N_48203,N_48595);
and UO_2390 (O_2390,N_49521,N_48298);
xor UO_2391 (O_2391,N_48593,N_48454);
xnor UO_2392 (O_2392,N_48885,N_48997);
and UO_2393 (O_2393,N_48868,N_49147);
nand UO_2394 (O_2394,N_48654,N_49190);
xnor UO_2395 (O_2395,N_48847,N_48234);
or UO_2396 (O_2396,N_49769,N_49024);
xnor UO_2397 (O_2397,N_49974,N_49967);
nand UO_2398 (O_2398,N_49941,N_49222);
or UO_2399 (O_2399,N_48918,N_49375);
nor UO_2400 (O_2400,N_48606,N_48125);
nand UO_2401 (O_2401,N_48086,N_48308);
nor UO_2402 (O_2402,N_48228,N_48269);
xor UO_2403 (O_2403,N_49240,N_49629);
nor UO_2404 (O_2404,N_48589,N_49150);
nor UO_2405 (O_2405,N_48385,N_49956);
and UO_2406 (O_2406,N_48372,N_48105);
nor UO_2407 (O_2407,N_48549,N_48069);
nand UO_2408 (O_2408,N_49729,N_49397);
or UO_2409 (O_2409,N_48427,N_48835);
nor UO_2410 (O_2410,N_49090,N_48389);
xor UO_2411 (O_2411,N_48270,N_49598);
and UO_2412 (O_2412,N_49723,N_49106);
nor UO_2413 (O_2413,N_49443,N_49705);
xnor UO_2414 (O_2414,N_49943,N_49633);
and UO_2415 (O_2415,N_49302,N_48239);
or UO_2416 (O_2416,N_48883,N_48401);
nor UO_2417 (O_2417,N_48194,N_49979);
nor UO_2418 (O_2418,N_48823,N_49650);
and UO_2419 (O_2419,N_48895,N_48580);
and UO_2420 (O_2420,N_48205,N_48772);
nor UO_2421 (O_2421,N_49382,N_49016);
xnor UO_2422 (O_2422,N_48165,N_48669);
and UO_2423 (O_2423,N_49096,N_49474);
or UO_2424 (O_2424,N_49591,N_49126);
nand UO_2425 (O_2425,N_49153,N_48734);
nand UO_2426 (O_2426,N_48551,N_49124);
or UO_2427 (O_2427,N_49188,N_49126);
nand UO_2428 (O_2428,N_49740,N_49090);
xnor UO_2429 (O_2429,N_48093,N_48261);
or UO_2430 (O_2430,N_48050,N_48253);
nand UO_2431 (O_2431,N_48674,N_49747);
xnor UO_2432 (O_2432,N_49013,N_48850);
nand UO_2433 (O_2433,N_48945,N_48121);
xnor UO_2434 (O_2434,N_48178,N_49224);
and UO_2435 (O_2435,N_49217,N_48634);
xor UO_2436 (O_2436,N_49248,N_48009);
nand UO_2437 (O_2437,N_49748,N_49316);
or UO_2438 (O_2438,N_48622,N_48702);
xnor UO_2439 (O_2439,N_48222,N_48868);
nor UO_2440 (O_2440,N_49498,N_49173);
nand UO_2441 (O_2441,N_49276,N_49169);
nor UO_2442 (O_2442,N_48348,N_48746);
or UO_2443 (O_2443,N_48427,N_48020);
nor UO_2444 (O_2444,N_49117,N_48594);
nand UO_2445 (O_2445,N_48365,N_49515);
xnor UO_2446 (O_2446,N_49056,N_48221);
or UO_2447 (O_2447,N_48736,N_49677);
nand UO_2448 (O_2448,N_48653,N_49606);
or UO_2449 (O_2449,N_49546,N_48022);
or UO_2450 (O_2450,N_49889,N_48173);
or UO_2451 (O_2451,N_49793,N_49932);
nand UO_2452 (O_2452,N_49380,N_49090);
nor UO_2453 (O_2453,N_49585,N_48944);
nand UO_2454 (O_2454,N_49296,N_48243);
and UO_2455 (O_2455,N_49440,N_49911);
nor UO_2456 (O_2456,N_49462,N_48620);
nor UO_2457 (O_2457,N_49783,N_49633);
or UO_2458 (O_2458,N_49064,N_48100);
and UO_2459 (O_2459,N_49968,N_49080);
and UO_2460 (O_2460,N_48960,N_48658);
or UO_2461 (O_2461,N_49504,N_49339);
and UO_2462 (O_2462,N_49941,N_49879);
nor UO_2463 (O_2463,N_48116,N_48782);
nor UO_2464 (O_2464,N_48419,N_49350);
and UO_2465 (O_2465,N_48388,N_48687);
and UO_2466 (O_2466,N_49973,N_48949);
and UO_2467 (O_2467,N_48123,N_49307);
nand UO_2468 (O_2468,N_48294,N_48191);
or UO_2469 (O_2469,N_48153,N_48421);
and UO_2470 (O_2470,N_49391,N_49121);
nand UO_2471 (O_2471,N_48118,N_48997);
xor UO_2472 (O_2472,N_49846,N_48763);
or UO_2473 (O_2473,N_48112,N_49047);
nand UO_2474 (O_2474,N_49657,N_49492);
or UO_2475 (O_2475,N_48547,N_48283);
nand UO_2476 (O_2476,N_49342,N_49542);
xor UO_2477 (O_2477,N_48198,N_49770);
nor UO_2478 (O_2478,N_49717,N_49410);
nor UO_2479 (O_2479,N_49061,N_49363);
and UO_2480 (O_2480,N_48752,N_48352);
or UO_2481 (O_2481,N_49316,N_49137);
nor UO_2482 (O_2482,N_49734,N_49092);
or UO_2483 (O_2483,N_49815,N_49413);
nor UO_2484 (O_2484,N_48382,N_48160);
nor UO_2485 (O_2485,N_49509,N_49810);
and UO_2486 (O_2486,N_49977,N_48178);
xor UO_2487 (O_2487,N_49549,N_49247);
nand UO_2488 (O_2488,N_48873,N_48750);
nor UO_2489 (O_2489,N_49771,N_49653);
nor UO_2490 (O_2490,N_48842,N_49014);
nand UO_2491 (O_2491,N_48696,N_49525);
or UO_2492 (O_2492,N_48356,N_48406);
and UO_2493 (O_2493,N_49516,N_49800);
or UO_2494 (O_2494,N_48975,N_48683);
nor UO_2495 (O_2495,N_48684,N_49462);
and UO_2496 (O_2496,N_49556,N_48002);
xnor UO_2497 (O_2497,N_48390,N_49947);
nand UO_2498 (O_2498,N_48370,N_49942);
or UO_2499 (O_2499,N_49363,N_48491);
or UO_2500 (O_2500,N_49098,N_49674);
nor UO_2501 (O_2501,N_48312,N_48830);
and UO_2502 (O_2502,N_49531,N_48087);
and UO_2503 (O_2503,N_48861,N_49662);
nor UO_2504 (O_2504,N_48546,N_49040);
and UO_2505 (O_2505,N_48882,N_48273);
and UO_2506 (O_2506,N_49983,N_49854);
nor UO_2507 (O_2507,N_48415,N_48136);
and UO_2508 (O_2508,N_48286,N_48152);
nand UO_2509 (O_2509,N_49218,N_49929);
and UO_2510 (O_2510,N_49752,N_49156);
nand UO_2511 (O_2511,N_49329,N_48887);
xnor UO_2512 (O_2512,N_48315,N_49827);
xnor UO_2513 (O_2513,N_48230,N_48647);
nor UO_2514 (O_2514,N_49745,N_49382);
or UO_2515 (O_2515,N_48181,N_49361);
xor UO_2516 (O_2516,N_49857,N_48874);
nor UO_2517 (O_2517,N_49432,N_48007);
xnor UO_2518 (O_2518,N_49624,N_48366);
nand UO_2519 (O_2519,N_49670,N_49589);
xnor UO_2520 (O_2520,N_49428,N_48188);
and UO_2521 (O_2521,N_48181,N_49979);
nand UO_2522 (O_2522,N_48489,N_49946);
nor UO_2523 (O_2523,N_48258,N_49346);
and UO_2524 (O_2524,N_49500,N_49775);
nor UO_2525 (O_2525,N_49941,N_48222);
nor UO_2526 (O_2526,N_48542,N_48920);
xor UO_2527 (O_2527,N_48817,N_49495);
and UO_2528 (O_2528,N_49841,N_49970);
or UO_2529 (O_2529,N_48631,N_49982);
nor UO_2530 (O_2530,N_49325,N_48162);
xor UO_2531 (O_2531,N_48367,N_49086);
and UO_2532 (O_2532,N_49253,N_48379);
or UO_2533 (O_2533,N_48595,N_48086);
xnor UO_2534 (O_2534,N_49583,N_48250);
nor UO_2535 (O_2535,N_49342,N_49064);
or UO_2536 (O_2536,N_49199,N_48697);
and UO_2537 (O_2537,N_48263,N_49484);
xnor UO_2538 (O_2538,N_48578,N_49465);
or UO_2539 (O_2539,N_49977,N_49685);
nand UO_2540 (O_2540,N_48593,N_49161);
xnor UO_2541 (O_2541,N_49022,N_48022);
xnor UO_2542 (O_2542,N_49450,N_48360);
nor UO_2543 (O_2543,N_49509,N_49349);
and UO_2544 (O_2544,N_48370,N_49022);
nand UO_2545 (O_2545,N_48266,N_49599);
and UO_2546 (O_2546,N_49670,N_49920);
nand UO_2547 (O_2547,N_49602,N_49836);
nand UO_2548 (O_2548,N_49977,N_49136);
and UO_2549 (O_2549,N_48028,N_48120);
and UO_2550 (O_2550,N_48689,N_49375);
or UO_2551 (O_2551,N_49355,N_49987);
and UO_2552 (O_2552,N_48578,N_49217);
or UO_2553 (O_2553,N_49868,N_49018);
or UO_2554 (O_2554,N_48050,N_48645);
xor UO_2555 (O_2555,N_49145,N_49274);
and UO_2556 (O_2556,N_48695,N_48984);
and UO_2557 (O_2557,N_49347,N_49201);
or UO_2558 (O_2558,N_48320,N_49517);
nor UO_2559 (O_2559,N_48164,N_49235);
nand UO_2560 (O_2560,N_49533,N_48781);
xor UO_2561 (O_2561,N_49170,N_48937);
nand UO_2562 (O_2562,N_48322,N_49018);
nor UO_2563 (O_2563,N_48382,N_48746);
nor UO_2564 (O_2564,N_49015,N_48515);
or UO_2565 (O_2565,N_48956,N_49413);
nand UO_2566 (O_2566,N_48350,N_48868);
nand UO_2567 (O_2567,N_48015,N_49832);
nor UO_2568 (O_2568,N_49523,N_48464);
xor UO_2569 (O_2569,N_48219,N_49143);
xor UO_2570 (O_2570,N_49792,N_49780);
nor UO_2571 (O_2571,N_49583,N_48560);
nor UO_2572 (O_2572,N_48682,N_49353);
or UO_2573 (O_2573,N_49964,N_49455);
and UO_2574 (O_2574,N_48863,N_48795);
nand UO_2575 (O_2575,N_49944,N_48729);
nand UO_2576 (O_2576,N_48913,N_48543);
nor UO_2577 (O_2577,N_48307,N_48956);
nor UO_2578 (O_2578,N_48983,N_48271);
xnor UO_2579 (O_2579,N_49815,N_48020);
and UO_2580 (O_2580,N_48337,N_49974);
or UO_2581 (O_2581,N_48978,N_49233);
xnor UO_2582 (O_2582,N_48324,N_48575);
nor UO_2583 (O_2583,N_49431,N_49724);
nand UO_2584 (O_2584,N_49291,N_49656);
or UO_2585 (O_2585,N_49643,N_49836);
or UO_2586 (O_2586,N_48371,N_48204);
nand UO_2587 (O_2587,N_48161,N_48715);
xor UO_2588 (O_2588,N_49192,N_48206);
xnor UO_2589 (O_2589,N_49915,N_49293);
nand UO_2590 (O_2590,N_48096,N_48664);
or UO_2591 (O_2591,N_49769,N_48890);
xor UO_2592 (O_2592,N_49025,N_48501);
and UO_2593 (O_2593,N_48909,N_48132);
or UO_2594 (O_2594,N_48820,N_49949);
and UO_2595 (O_2595,N_49854,N_48552);
xor UO_2596 (O_2596,N_48853,N_48492);
xor UO_2597 (O_2597,N_49106,N_49614);
and UO_2598 (O_2598,N_49368,N_48600);
xnor UO_2599 (O_2599,N_49413,N_48541);
nor UO_2600 (O_2600,N_48835,N_49223);
nor UO_2601 (O_2601,N_48918,N_48829);
nand UO_2602 (O_2602,N_49137,N_48958);
and UO_2603 (O_2603,N_48637,N_49085);
or UO_2604 (O_2604,N_48491,N_49124);
nand UO_2605 (O_2605,N_49456,N_48299);
xnor UO_2606 (O_2606,N_49540,N_49220);
and UO_2607 (O_2607,N_49269,N_48901);
nand UO_2608 (O_2608,N_48144,N_48747);
or UO_2609 (O_2609,N_48270,N_49678);
nor UO_2610 (O_2610,N_49196,N_48890);
or UO_2611 (O_2611,N_49431,N_48559);
nor UO_2612 (O_2612,N_48449,N_49297);
or UO_2613 (O_2613,N_49265,N_49865);
nand UO_2614 (O_2614,N_48235,N_49979);
or UO_2615 (O_2615,N_48936,N_48077);
nor UO_2616 (O_2616,N_49802,N_49130);
xor UO_2617 (O_2617,N_48779,N_49554);
nand UO_2618 (O_2618,N_49128,N_48912);
nand UO_2619 (O_2619,N_48032,N_49789);
or UO_2620 (O_2620,N_48845,N_49371);
xor UO_2621 (O_2621,N_49121,N_49368);
or UO_2622 (O_2622,N_48684,N_48643);
xnor UO_2623 (O_2623,N_48100,N_49815);
xor UO_2624 (O_2624,N_49888,N_48312);
and UO_2625 (O_2625,N_49703,N_48508);
or UO_2626 (O_2626,N_48299,N_48479);
nand UO_2627 (O_2627,N_48742,N_48215);
and UO_2628 (O_2628,N_48757,N_48987);
nand UO_2629 (O_2629,N_49407,N_49222);
nand UO_2630 (O_2630,N_48498,N_48639);
xor UO_2631 (O_2631,N_48837,N_49740);
nand UO_2632 (O_2632,N_49988,N_49145);
or UO_2633 (O_2633,N_49911,N_48503);
and UO_2634 (O_2634,N_49033,N_48493);
nor UO_2635 (O_2635,N_49171,N_48181);
xor UO_2636 (O_2636,N_48898,N_49484);
or UO_2637 (O_2637,N_48892,N_48280);
and UO_2638 (O_2638,N_48363,N_48227);
nand UO_2639 (O_2639,N_49727,N_49100);
or UO_2640 (O_2640,N_49592,N_48310);
and UO_2641 (O_2641,N_48531,N_49996);
nand UO_2642 (O_2642,N_48683,N_48162);
or UO_2643 (O_2643,N_49636,N_49236);
nand UO_2644 (O_2644,N_49081,N_49068);
nor UO_2645 (O_2645,N_48113,N_48504);
xor UO_2646 (O_2646,N_48401,N_49858);
and UO_2647 (O_2647,N_48601,N_49847);
xor UO_2648 (O_2648,N_49220,N_48267);
xor UO_2649 (O_2649,N_48305,N_49336);
nand UO_2650 (O_2650,N_48249,N_48925);
nand UO_2651 (O_2651,N_48617,N_49780);
nand UO_2652 (O_2652,N_48845,N_48063);
and UO_2653 (O_2653,N_49305,N_48975);
nor UO_2654 (O_2654,N_48610,N_49902);
nor UO_2655 (O_2655,N_49250,N_49647);
or UO_2656 (O_2656,N_48858,N_49088);
or UO_2657 (O_2657,N_48316,N_49739);
nand UO_2658 (O_2658,N_49544,N_48810);
and UO_2659 (O_2659,N_48524,N_48346);
nand UO_2660 (O_2660,N_48996,N_48790);
and UO_2661 (O_2661,N_48717,N_49707);
nand UO_2662 (O_2662,N_49327,N_48400);
and UO_2663 (O_2663,N_49396,N_48265);
or UO_2664 (O_2664,N_49847,N_48596);
xnor UO_2665 (O_2665,N_49873,N_49595);
and UO_2666 (O_2666,N_48735,N_49597);
xor UO_2667 (O_2667,N_49981,N_49920);
nor UO_2668 (O_2668,N_49651,N_48695);
xnor UO_2669 (O_2669,N_48853,N_49890);
xnor UO_2670 (O_2670,N_49284,N_48783);
or UO_2671 (O_2671,N_48199,N_48263);
xor UO_2672 (O_2672,N_48768,N_49495);
and UO_2673 (O_2673,N_48549,N_49430);
xnor UO_2674 (O_2674,N_49835,N_49019);
xor UO_2675 (O_2675,N_49649,N_48285);
nor UO_2676 (O_2676,N_48909,N_49623);
and UO_2677 (O_2677,N_48469,N_49407);
and UO_2678 (O_2678,N_48708,N_49996);
xnor UO_2679 (O_2679,N_49524,N_49102);
xnor UO_2680 (O_2680,N_48424,N_49085);
nor UO_2681 (O_2681,N_49819,N_49889);
and UO_2682 (O_2682,N_49750,N_49188);
xnor UO_2683 (O_2683,N_48085,N_48364);
xnor UO_2684 (O_2684,N_48463,N_49875);
nor UO_2685 (O_2685,N_49240,N_48675);
or UO_2686 (O_2686,N_49916,N_48503);
nand UO_2687 (O_2687,N_49594,N_49577);
or UO_2688 (O_2688,N_49420,N_49166);
or UO_2689 (O_2689,N_49138,N_49211);
and UO_2690 (O_2690,N_49758,N_49031);
and UO_2691 (O_2691,N_48057,N_49409);
or UO_2692 (O_2692,N_48776,N_48240);
xor UO_2693 (O_2693,N_49451,N_48646);
or UO_2694 (O_2694,N_49931,N_49189);
xor UO_2695 (O_2695,N_49639,N_48137);
and UO_2696 (O_2696,N_48542,N_49209);
nand UO_2697 (O_2697,N_48935,N_48510);
xnor UO_2698 (O_2698,N_49456,N_49487);
nand UO_2699 (O_2699,N_49959,N_48813);
xor UO_2700 (O_2700,N_48122,N_48257);
xnor UO_2701 (O_2701,N_48398,N_49344);
or UO_2702 (O_2702,N_49456,N_48349);
and UO_2703 (O_2703,N_49467,N_48555);
or UO_2704 (O_2704,N_49136,N_48168);
and UO_2705 (O_2705,N_48059,N_49888);
and UO_2706 (O_2706,N_49539,N_49075);
xor UO_2707 (O_2707,N_49622,N_48959);
nand UO_2708 (O_2708,N_48003,N_48274);
nor UO_2709 (O_2709,N_49306,N_48022);
xor UO_2710 (O_2710,N_48132,N_49984);
and UO_2711 (O_2711,N_48647,N_49203);
and UO_2712 (O_2712,N_48865,N_49782);
xnor UO_2713 (O_2713,N_49989,N_49908);
or UO_2714 (O_2714,N_48223,N_49345);
nor UO_2715 (O_2715,N_49460,N_49083);
and UO_2716 (O_2716,N_49362,N_49254);
nand UO_2717 (O_2717,N_49646,N_49324);
or UO_2718 (O_2718,N_48006,N_49279);
and UO_2719 (O_2719,N_49176,N_49025);
and UO_2720 (O_2720,N_48609,N_49923);
nand UO_2721 (O_2721,N_48475,N_48640);
and UO_2722 (O_2722,N_49631,N_49951);
or UO_2723 (O_2723,N_48512,N_49184);
nand UO_2724 (O_2724,N_49797,N_49053);
xor UO_2725 (O_2725,N_49125,N_49392);
xor UO_2726 (O_2726,N_49049,N_49696);
or UO_2727 (O_2727,N_49872,N_49680);
and UO_2728 (O_2728,N_48216,N_48869);
xnor UO_2729 (O_2729,N_48833,N_48631);
nor UO_2730 (O_2730,N_48097,N_48399);
nor UO_2731 (O_2731,N_48383,N_49308);
or UO_2732 (O_2732,N_49304,N_48639);
nand UO_2733 (O_2733,N_48199,N_49164);
nand UO_2734 (O_2734,N_48702,N_48390);
or UO_2735 (O_2735,N_48052,N_49162);
xnor UO_2736 (O_2736,N_49460,N_49465);
xnor UO_2737 (O_2737,N_48479,N_49246);
nor UO_2738 (O_2738,N_48850,N_49227);
nand UO_2739 (O_2739,N_49331,N_49693);
xnor UO_2740 (O_2740,N_48157,N_49654);
and UO_2741 (O_2741,N_49360,N_49252);
and UO_2742 (O_2742,N_49565,N_48270);
nor UO_2743 (O_2743,N_48712,N_48001);
or UO_2744 (O_2744,N_48680,N_48643);
or UO_2745 (O_2745,N_49133,N_49694);
xnor UO_2746 (O_2746,N_49490,N_49876);
and UO_2747 (O_2747,N_49263,N_48270);
or UO_2748 (O_2748,N_49158,N_48086);
nand UO_2749 (O_2749,N_49423,N_49530);
nand UO_2750 (O_2750,N_48360,N_48683);
and UO_2751 (O_2751,N_48951,N_49206);
nand UO_2752 (O_2752,N_49422,N_48401);
or UO_2753 (O_2753,N_48998,N_48796);
and UO_2754 (O_2754,N_49323,N_49286);
nand UO_2755 (O_2755,N_49571,N_49023);
nor UO_2756 (O_2756,N_48927,N_48027);
or UO_2757 (O_2757,N_49307,N_49722);
and UO_2758 (O_2758,N_49878,N_48814);
nor UO_2759 (O_2759,N_49885,N_49863);
or UO_2760 (O_2760,N_49032,N_48801);
and UO_2761 (O_2761,N_48979,N_49575);
and UO_2762 (O_2762,N_48823,N_48516);
nor UO_2763 (O_2763,N_49325,N_48345);
or UO_2764 (O_2764,N_49781,N_48739);
xnor UO_2765 (O_2765,N_49305,N_49658);
or UO_2766 (O_2766,N_48304,N_49166);
nand UO_2767 (O_2767,N_48203,N_49991);
xor UO_2768 (O_2768,N_49488,N_48521);
xnor UO_2769 (O_2769,N_49758,N_49742);
and UO_2770 (O_2770,N_48897,N_49228);
nor UO_2771 (O_2771,N_48386,N_48694);
nand UO_2772 (O_2772,N_48773,N_48428);
xnor UO_2773 (O_2773,N_48939,N_49112);
or UO_2774 (O_2774,N_49985,N_49949);
nor UO_2775 (O_2775,N_48350,N_49209);
and UO_2776 (O_2776,N_48885,N_48257);
and UO_2777 (O_2777,N_48750,N_49350);
xor UO_2778 (O_2778,N_49965,N_49135);
and UO_2779 (O_2779,N_49586,N_48665);
nand UO_2780 (O_2780,N_49942,N_49289);
and UO_2781 (O_2781,N_48107,N_48265);
nand UO_2782 (O_2782,N_49556,N_48963);
nand UO_2783 (O_2783,N_49347,N_49370);
xnor UO_2784 (O_2784,N_48573,N_49628);
and UO_2785 (O_2785,N_48232,N_48406);
xnor UO_2786 (O_2786,N_49622,N_48323);
nor UO_2787 (O_2787,N_49746,N_49389);
or UO_2788 (O_2788,N_48158,N_49591);
nor UO_2789 (O_2789,N_48883,N_48412);
or UO_2790 (O_2790,N_49711,N_48623);
or UO_2791 (O_2791,N_48108,N_48592);
nand UO_2792 (O_2792,N_48569,N_48521);
xnor UO_2793 (O_2793,N_49893,N_48177);
xnor UO_2794 (O_2794,N_49824,N_49799);
xnor UO_2795 (O_2795,N_49702,N_49032);
nand UO_2796 (O_2796,N_49910,N_49900);
or UO_2797 (O_2797,N_49353,N_49087);
nor UO_2798 (O_2798,N_49372,N_49142);
nand UO_2799 (O_2799,N_48265,N_48551);
and UO_2800 (O_2800,N_49319,N_48907);
or UO_2801 (O_2801,N_49737,N_49450);
nor UO_2802 (O_2802,N_49002,N_49530);
nand UO_2803 (O_2803,N_49747,N_48234);
xor UO_2804 (O_2804,N_49709,N_49264);
nand UO_2805 (O_2805,N_49991,N_48830);
nand UO_2806 (O_2806,N_49645,N_49620);
xnor UO_2807 (O_2807,N_48834,N_48056);
xnor UO_2808 (O_2808,N_49063,N_49529);
nand UO_2809 (O_2809,N_49214,N_48314);
nand UO_2810 (O_2810,N_49410,N_48491);
xnor UO_2811 (O_2811,N_49012,N_48573);
or UO_2812 (O_2812,N_49337,N_49971);
nand UO_2813 (O_2813,N_48531,N_49321);
or UO_2814 (O_2814,N_49332,N_48050);
nand UO_2815 (O_2815,N_48945,N_49722);
and UO_2816 (O_2816,N_49228,N_48578);
or UO_2817 (O_2817,N_48073,N_49985);
xor UO_2818 (O_2818,N_49031,N_49699);
or UO_2819 (O_2819,N_48197,N_49603);
nand UO_2820 (O_2820,N_49810,N_49244);
and UO_2821 (O_2821,N_48049,N_48944);
or UO_2822 (O_2822,N_48463,N_48542);
and UO_2823 (O_2823,N_49941,N_49875);
or UO_2824 (O_2824,N_48813,N_48560);
nand UO_2825 (O_2825,N_48001,N_49897);
nand UO_2826 (O_2826,N_49429,N_48391);
and UO_2827 (O_2827,N_49066,N_49780);
xnor UO_2828 (O_2828,N_48325,N_49054);
nor UO_2829 (O_2829,N_49286,N_49926);
nor UO_2830 (O_2830,N_49054,N_48319);
and UO_2831 (O_2831,N_48029,N_49828);
nor UO_2832 (O_2832,N_48661,N_49736);
and UO_2833 (O_2833,N_49495,N_49142);
nand UO_2834 (O_2834,N_49476,N_49677);
and UO_2835 (O_2835,N_49212,N_49044);
and UO_2836 (O_2836,N_48874,N_49867);
nand UO_2837 (O_2837,N_49175,N_49188);
xor UO_2838 (O_2838,N_49882,N_49047);
and UO_2839 (O_2839,N_49044,N_48128);
xor UO_2840 (O_2840,N_49117,N_49355);
or UO_2841 (O_2841,N_49177,N_49088);
nor UO_2842 (O_2842,N_49535,N_48582);
xnor UO_2843 (O_2843,N_49582,N_48644);
nand UO_2844 (O_2844,N_48903,N_48087);
xor UO_2845 (O_2845,N_48692,N_48445);
xnor UO_2846 (O_2846,N_48744,N_49758);
and UO_2847 (O_2847,N_48310,N_48657);
nand UO_2848 (O_2848,N_48534,N_49683);
and UO_2849 (O_2849,N_48796,N_48528);
xor UO_2850 (O_2850,N_48424,N_49520);
or UO_2851 (O_2851,N_49182,N_48261);
or UO_2852 (O_2852,N_49969,N_49423);
xnor UO_2853 (O_2853,N_48822,N_49351);
nand UO_2854 (O_2854,N_49406,N_49632);
xor UO_2855 (O_2855,N_48795,N_48016);
and UO_2856 (O_2856,N_49125,N_48462);
and UO_2857 (O_2857,N_48003,N_49425);
or UO_2858 (O_2858,N_48743,N_49812);
and UO_2859 (O_2859,N_48796,N_49125);
xor UO_2860 (O_2860,N_48338,N_48959);
nor UO_2861 (O_2861,N_48731,N_48391);
or UO_2862 (O_2862,N_49348,N_49744);
and UO_2863 (O_2863,N_48735,N_49192);
and UO_2864 (O_2864,N_48887,N_48256);
nand UO_2865 (O_2865,N_48549,N_48736);
or UO_2866 (O_2866,N_48009,N_48830);
and UO_2867 (O_2867,N_49354,N_49592);
nand UO_2868 (O_2868,N_49569,N_49650);
xnor UO_2869 (O_2869,N_49144,N_49863);
nor UO_2870 (O_2870,N_48544,N_49241);
and UO_2871 (O_2871,N_49131,N_48984);
nand UO_2872 (O_2872,N_48326,N_49928);
and UO_2873 (O_2873,N_48192,N_49182);
nand UO_2874 (O_2874,N_49200,N_48121);
xor UO_2875 (O_2875,N_48287,N_49591);
or UO_2876 (O_2876,N_48367,N_49634);
or UO_2877 (O_2877,N_48191,N_48844);
or UO_2878 (O_2878,N_49643,N_49909);
and UO_2879 (O_2879,N_49482,N_48346);
or UO_2880 (O_2880,N_49499,N_48070);
or UO_2881 (O_2881,N_49816,N_49553);
nand UO_2882 (O_2882,N_48393,N_48822);
or UO_2883 (O_2883,N_48306,N_49971);
nor UO_2884 (O_2884,N_48008,N_49732);
nor UO_2885 (O_2885,N_49361,N_48476);
xnor UO_2886 (O_2886,N_49750,N_48685);
xor UO_2887 (O_2887,N_49432,N_49414);
or UO_2888 (O_2888,N_49840,N_49229);
nand UO_2889 (O_2889,N_48647,N_49776);
or UO_2890 (O_2890,N_49749,N_48915);
and UO_2891 (O_2891,N_48206,N_48143);
xor UO_2892 (O_2892,N_48733,N_49983);
nor UO_2893 (O_2893,N_49787,N_48102);
xor UO_2894 (O_2894,N_49164,N_49991);
nor UO_2895 (O_2895,N_49464,N_48622);
xnor UO_2896 (O_2896,N_49351,N_48338);
or UO_2897 (O_2897,N_48658,N_48782);
nand UO_2898 (O_2898,N_48427,N_48100);
and UO_2899 (O_2899,N_48731,N_48169);
xor UO_2900 (O_2900,N_49911,N_49172);
nor UO_2901 (O_2901,N_48573,N_49396);
nor UO_2902 (O_2902,N_49490,N_49606);
xnor UO_2903 (O_2903,N_49012,N_48148);
or UO_2904 (O_2904,N_49205,N_49516);
or UO_2905 (O_2905,N_48214,N_48448);
and UO_2906 (O_2906,N_49444,N_49401);
nand UO_2907 (O_2907,N_49172,N_49107);
nor UO_2908 (O_2908,N_48720,N_48694);
or UO_2909 (O_2909,N_49800,N_48184);
nor UO_2910 (O_2910,N_49887,N_49868);
nand UO_2911 (O_2911,N_49701,N_49224);
nor UO_2912 (O_2912,N_48801,N_48570);
nand UO_2913 (O_2913,N_48774,N_49755);
nor UO_2914 (O_2914,N_49343,N_48675);
nor UO_2915 (O_2915,N_49909,N_49700);
or UO_2916 (O_2916,N_49260,N_49774);
nor UO_2917 (O_2917,N_48147,N_49595);
nor UO_2918 (O_2918,N_49271,N_49077);
nand UO_2919 (O_2919,N_48212,N_49285);
and UO_2920 (O_2920,N_48626,N_49048);
and UO_2921 (O_2921,N_48457,N_48023);
or UO_2922 (O_2922,N_49026,N_49852);
or UO_2923 (O_2923,N_49845,N_49574);
or UO_2924 (O_2924,N_48104,N_48712);
xor UO_2925 (O_2925,N_48958,N_49498);
nor UO_2926 (O_2926,N_49578,N_48834);
xnor UO_2927 (O_2927,N_48883,N_49815);
xnor UO_2928 (O_2928,N_49207,N_48206);
or UO_2929 (O_2929,N_48265,N_48998);
or UO_2930 (O_2930,N_49950,N_49254);
or UO_2931 (O_2931,N_48218,N_49201);
nand UO_2932 (O_2932,N_48695,N_49347);
or UO_2933 (O_2933,N_49387,N_49361);
nor UO_2934 (O_2934,N_49351,N_48258);
nand UO_2935 (O_2935,N_49141,N_49761);
nor UO_2936 (O_2936,N_49865,N_48264);
and UO_2937 (O_2937,N_49897,N_49028);
or UO_2938 (O_2938,N_49448,N_49011);
nand UO_2939 (O_2939,N_48386,N_48721);
and UO_2940 (O_2940,N_48176,N_48168);
and UO_2941 (O_2941,N_48965,N_48200);
nor UO_2942 (O_2942,N_48625,N_48413);
xor UO_2943 (O_2943,N_48949,N_48846);
and UO_2944 (O_2944,N_49204,N_48540);
nor UO_2945 (O_2945,N_48108,N_49253);
and UO_2946 (O_2946,N_49973,N_49721);
nand UO_2947 (O_2947,N_48357,N_48350);
nor UO_2948 (O_2948,N_49341,N_49990);
nor UO_2949 (O_2949,N_49155,N_48747);
or UO_2950 (O_2950,N_49404,N_49413);
and UO_2951 (O_2951,N_49532,N_48655);
nor UO_2952 (O_2952,N_48671,N_49047);
and UO_2953 (O_2953,N_49432,N_48450);
and UO_2954 (O_2954,N_48035,N_48922);
and UO_2955 (O_2955,N_49888,N_48988);
nor UO_2956 (O_2956,N_49797,N_48504);
xnor UO_2957 (O_2957,N_49688,N_49641);
and UO_2958 (O_2958,N_48505,N_49674);
or UO_2959 (O_2959,N_49774,N_49183);
xor UO_2960 (O_2960,N_48800,N_49165);
and UO_2961 (O_2961,N_49050,N_48350);
nand UO_2962 (O_2962,N_48755,N_49892);
nor UO_2963 (O_2963,N_48737,N_48817);
or UO_2964 (O_2964,N_49418,N_49991);
and UO_2965 (O_2965,N_49744,N_48684);
and UO_2966 (O_2966,N_49717,N_48421);
and UO_2967 (O_2967,N_49949,N_48416);
or UO_2968 (O_2968,N_48323,N_49527);
xor UO_2969 (O_2969,N_48475,N_48628);
nor UO_2970 (O_2970,N_48364,N_48055);
xor UO_2971 (O_2971,N_48500,N_48925);
or UO_2972 (O_2972,N_49128,N_48334);
nor UO_2973 (O_2973,N_49042,N_49534);
nor UO_2974 (O_2974,N_49299,N_49978);
and UO_2975 (O_2975,N_49837,N_48690);
nor UO_2976 (O_2976,N_49998,N_49417);
or UO_2977 (O_2977,N_49890,N_48103);
xor UO_2978 (O_2978,N_49481,N_49409);
xor UO_2979 (O_2979,N_48697,N_49870);
xor UO_2980 (O_2980,N_49643,N_49008);
xnor UO_2981 (O_2981,N_49038,N_49027);
and UO_2982 (O_2982,N_49459,N_48593);
or UO_2983 (O_2983,N_49272,N_48815);
nor UO_2984 (O_2984,N_49199,N_48541);
nand UO_2985 (O_2985,N_49886,N_49180);
or UO_2986 (O_2986,N_49252,N_49085);
nand UO_2987 (O_2987,N_49439,N_48829);
nor UO_2988 (O_2988,N_48749,N_48521);
xnor UO_2989 (O_2989,N_49827,N_49431);
xor UO_2990 (O_2990,N_48365,N_49521);
nor UO_2991 (O_2991,N_49530,N_49337);
nand UO_2992 (O_2992,N_48837,N_48914);
or UO_2993 (O_2993,N_49982,N_49816);
or UO_2994 (O_2994,N_49572,N_49754);
xor UO_2995 (O_2995,N_48695,N_49403);
xnor UO_2996 (O_2996,N_49977,N_49526);
and UO_2997 (O_2997,N_49493,N_48151);
nor UO_2998 (O_2998,N_48445,N_48178);
xnor UO_2999 (O_2999,N_48627,N_48990);
nand UO_3000 (O_3000,N_49967,N_49420);
nor UO_3001 (O_3001,N_48829,N_48312);
or UO_3002 (O_3002,N_48530,N_49198);
nor UO_3003 (O_3003,N_49277,N_48130);
nor UO_3004 (O_3004,N_48475,N_49561);
nand UO_3005 (O_3005,N_49921,N_49235);
nor UO_3006 (O_3006,N_49174,N_48477);
xor UO_3007 (O_3007,N_49976,N_49219);
and UO_3008 (O_3008,N_49084,N_49408);
xnor UO_3009 (O_3009,N_48753,N_48404);
nor UO_3010 (O_3010,N_48835,N_49975);
or UO_3011 (O_3011,N_48023,N_49542);
nand UO_3012 (O_3012,N_49583,N_48692);
nor UO_3013 (O_3013,N_49545,N_48440);
and UO_3014 (O_3014,N_48907,N_48165);
xnor UO_3015 (O_3015,N_48256,N_49908);
or UO_3016 (O_3016,N_49521,N_48535);
and UO_3017 (O_3017,N_49304,N_49055);
and UO_3018 (O_3018,N_48745,N_48182);
nor UO_3019 (O_3019,N_48793,N_49380);
nor UO_3020 (O_3020,N_48754,N_48960);
or UO_3021 (O_3021,N_48988,N_48134);
and UO_3022 (O_3022,N_49584,N_48581);
and UO_3023 (O_3023,N_49183,N_49161);
or UO_3024 (O_3024,N_48264,N_48375);
nand UO_3025 (O_3025,N_49666,N_48103);
and UO_3026 (O_3026,N_48937,N_48845);
nand UO_3027 (O_3027,N_48507,N_49197);
nand UO_3028 (O_3028,N_48528,N_49899);
nor UO_3029 (O_3029,N_49905,N_49890);
and UO_3030 (O_3030,N_49916,N_49566);
and UO_3031 (O_3031,N_49379,N_48503);
nand UO_3032 (O_3032,N_49015,N_49370);
nor UO_3033 (O_3033,N_48602,N_48654);
nand UO_3034 (O_3034,N_49624,N_49991);
or UO_3035 (O_3035,N_49021,N_48428);
and UO_3036 (O_3036,N_48515,N_49366);
or UO_3037 (O_3037,N_49250,N_48375);
nor UO_3038 (O_3038,N_48550,N_49595);
and UO_3039 (O_3039,N_49090,N_49933);
xor UO_3040 (O_3040,N_48585,N_49209);
or UO_3041 (O_3041,N_49383,N_48811);
nor UO_3042 (O_3042,N_48820,N_48185);
and UO_3043 (O_3043,N_48807,N_49329);
and UO_3044 (O_3044,N_48712,N_48562);
nand UO_3045 (O_3045,N_48534,N_49789);
or UO_3046 (O_3046,N_48501,N_48838);
nand UO_3047 (O_3047,N_49495,N_49995);
nand UO_3048 (O_3048,N_48899,N_49984);
or UO_3049 (O_3049,N_49645,N_48651);
and UO_3050 (O_3050,N_49331,N_48977);
nand UO_3051 (O_3051,N_49365,N_48802);
or UO_3052 (O_3052,N_49720,N_49909);
nor UO_3053 (O_3053,N_49287,N_49105);
nand UO_3054 (O_3054,N_49298,N_48573);
nand UO_3055 (O_3055,N_48991,N_49412);
xnor UO_3056 (O_3056,N_48440,N_49381);
nor UO_3057 (O_3057,N_48159,N_48247);
nor UO_3058 (O_3058,N_49594,N_48251);
and UO_3059 (O_3059,N_48036,N_48370);
nand UO_3060 (O_3060,N_48455,N_49224);
xnor UO_3061 (O_3061,N_48675,N_48354);
nor UO_3062 (O_3062,N_49553,N_49614);
or UO_3063 (O_3063,N_49171,N_48052);
nand UO_3064 (O_3064,N_49816,N_49693);
or UO_3065 (O_3065,N_48292,N_49366);
or UO_3066 (O_3066,N_48586,N_49592);
or UO_3067 (O_3067,N_49382,N_49966);
xor UO_3068 (O_3068,N_49547,N_49126);
nand UO_3069 (O_3069,N_49819,N_49011);
nor UO_3070 (O_3070,N_48393,N_49183);
nor UO_3071 (O_3071,N_48543,N_48521);
nor UO_3072 (O_3072,N_48231,N_48601);
or UO_3073 (O_3073,N_48180,N_48519);
nand UO_3074 (O_3074,N_49881,N_48106);
nor UO_3075 (O_3075,N_48466,N_48486);
and UO_3076 (O_3076,N_49751,N_49385);
and UO_3077 (O_3077,N_48256,N_49194);
nor UO_3078 (O_3078,N_48779,N_48741);
nand UO_3079 (O_3079,N_48621,N_48322);
xor UO_3080 (O_3080,N_48546,N_48814);
and UO_3081 (O_3081,N_49123,N_48875);
and UO_3082 (O_3082,N_49960,N_48260);
nor UO_3083 (O_3083,N_49129,N_49170);
nor UO_3084 (O_3084,N_49886,N_48419);
nor UO_3085 (O_3085,N_49057,N_48926);
or UO_3086 (O_3086,N_48246,N_48521);
xor UO_3087 (O_3087,N_48890,N_49351);
nand UO_3088 (O_3088,N_49331,N_48928);
or UO_3089 (O_3089,N_49204,N_49040);
nand UO_3090 (O_3090,N_48675,N_49285);
nor UO_3091 (O_3091,N_48341,N_49597);
and UO_3092 (O_3092,N_49711,N_48093);
nor UO_3093 (O_3093,N_49236,N_49662);
and UO_3094 (O_3094,N_48046,N_48897);
or UO_3095 (O_3095,N_48806,N_49075);
nand UO_3096 (O_3096,N_48665,N_48779);
xnor UO_3097 (O_3097,N_49064,N_49383);
or UO_3098 (O_3098,N_48317,N_48888);
xnor UO_3099 (O_3099,N_49196,N_49818);
or UO_3100 (O_3100,N_49630,N_48075);
nand UO_3101 (O_3101,N_49107,N_49336);
nand UO_3102 (O_3102,N_48826,N_49628);
and UO_3103 (O_3103,N_49720,N_49857);
nor UO_3104 (O_3104,N_49095,N_49580);
or UO_3105 (O_3105,N_49803,N_49742);
xor UO_3106 (O_3106,N_48881,N_48575);
or UO_3107 (O_3107,N_48196,N_49331);
nor UO_3108 (O_3108,N_48947,N_49386);
and UO_3109 (O_3109,N_49716,N_49289);
and UO_3110 (O_3110,N_49790,N_49147);
nand UO_3111 (O_3111,N_48787,N_49952);
nor UO_3112 (O_3112,N_49288,N_48319);
or UO_3113 (O_3113,N_49653,N_48720);
xor UO_3114 (O_3114,N_48081,N_49834);
or UO_3115 (O_3115,N_49192,N_49462);
and UO_3116 (O_3116,N_49335,N_49309);
xnor UO_3117 (O_3117,N_49858,N_49850);
nor UO_3118 (O_3118,N_48500,N_49388);
xor UO_3119 (O_3119,N_48941,N_49940);
or UO_3120 (O_3120,N_49958,N_49562);
and UO_3121 (O_3121,N_48871,N_49175);
nand UO_3122 (O_3122,N_49800,N_48596);
and UO_3123 (O_3123,N_49653,N_48641);
or UO_3124 (O_3124,N_49254,N_48963);
xnor UO_3125 (O_3125,N_49963,N_49689);
xnor UO_3126 (O_3126,N_48766,N_49571);
nand UO_3127 (O_3127,N_49168,N_49895);
and UO_3128 (O_3128,N_49742,N_48368);
nor UO_3129 (O_3129,N_49793,N_48220);
nor UO_3130 (O_3130,N_49562,N_49625);
xnor UO_3131 (O_3131,N_49206,N_48485);
nand UO_3132 (O_3132,N_48664,N_49017);
xor UO_3133 (O_3133,N_49293,N_49380);
nand UO_3134 (O_3134,N_48048,N_49799);
nor UO_3135 (O_3135,N_49640,N_49798);
nand UO_3136 (O_3136,N_48099,N_49250);
or UO_3137 (O_3137,N_48026,N_49509);
xor UO_3138 (O_3138,N_48234,N_48439);
and UO_3139 (O_3139,N_49611,N_49182);
xor UO_3140 (O_3140,N_49566,N_49866);
xor UO_3141 (O_3141,N_49490,N_49748);
or UO_3142 (O_3142,N_49735,N_49823);
xor UO_3143 (O_3143,N_49573,N_48761);
nand UO_3144 (O_3144,N_48826,N_48684);
nand UO_3145 (O_3145,N_49185,N_48725);
xnor UO_3146 (O_3146,N_48130,N_49628);
and UO_3147 (O_3147,N_48310,N_48465);
nor UO_3148 (O_3148,N_48892,N_49305);
nor UO_3149 (O_3149,N_49958,N_48431);
and UO_3150 (O_3150,N_48590,N_49620);
nor UO_3151 (O_3151,N_48725,N_49689);
nand UO_3152 (O_3152,N_48901,N_48824);
or UO_3153 (O_3153,N_48702,N_49275);
or UO_3154 (O_3154,N_48784,N_49346);
xnor UO_3155 (O_3155,N_48792,N_49973);
or UO_3156 (O_3156,N_48926,N_48704);
or UO_3157 (O_3157,N_48305,N_48481);
and UO_3158 (O_3158,N_49530,N_49414);
or UO_3159 (O_3159,N_48244,N_48908);
nor UO_3160 (O_3160,N_48359,N_48995);
and UO_3161 (O_3161,N_48406,N_49679);
nand UO_3162 (O_3162,N_48167,N_48250);
and UO_3163 (O_3163,N_49761,N_48049);
or UO_3164 (O_3164,N_49431,N_49487);
and UO_3165 (O_3165,N_49878,N_48978);
nand UO_3166 (O_3166,N_48874,N_48901);
and UO_3167 (O_3167,N_48379,N_48846);
nand UO_3168 (O_3168,N_48604,N_48327);
and UO_3169 (O_3169,N_49302,N_48429);
and UO_3170 (O_3170,N_49290,N_48544);
xnor UO_3171 (O_3171,N_48226,N_49856);
nor UO_3172 (O_3172,N_48049,N_48785);
nor UO_3173 (O_3173,N_49647,N_48571);
or UO_3174 (O_3174,N_48123,N_48650);
nor UO_3175 (O_3175,N_48132,N_48726);
xnor UO_3176 (O_3176,N_49193,N_49819);
and UO_3177 (O_3177,N_48524,N_48982);
nand UO_3178 (O_3178,N_48632,N_48639);
and UO_3179 (O_3179,N_48627,N_49775);
xor UO_3180 (O_3180,N_48753,N_48825);
or UO_3181 (O_3181,N_48597,N_48580);
nor UO_3182 (O_3182,N_49494,N_49722);
or UO_3183 (O_3183,N_49656,N_48701);
nand UO_3184 (O_3184,N_49409,N_49140);
nor UO_3185 (O_3185,N_48703,N_49575);
nor UO_3186 (O_3186,N_48104,N_48286);
nor UO_3187 (O_3187,N_48011,N_48480);
or UO_3188 (O_3188,N_49657,N_49929);
nor UO_3189 (O_3189,N_49402,N_49233);
or UO_3190 (O_3190,N_49289,N_48572);
nand UO_3191 (O_3191,N_49824,N_48940);
nor UO_3192 (O_3192,N_49972,N_48744);
and UO_3193 (O_3193,N_48265,N_49390);
nand UO_3194 (O_3194,N_48577,N_49000);
xor UO_3195 (O_3195,N_48474,N_48521);
and UO_3196 (O_3196,N_49110,N_49008);
or UO_3197 (O_3197,N_49324,N_49755);
nor UO_3198 (O_3198,N_49728,N_48346);
and UO_3199 (O_3199,N_49645,N_49335);
nand UO_3200 (O_3200,N_48832,N_49212);
and UO_3201 (O_3201,N_48242,N_49708);
nor UO_3202 (O_3202,N_49187,N_48296);
nor UO_3203 (O_3203,N_49438,N_49839);
nor UO_3204 (O_3204,N_49011,N_49551);
xor UO_3205 (O_3205,N_48119,N_49756);
and UO_3206 (O_3206,N_48846,N_49985);
nor UO_3207 (O_3207,N_48280,N_49149);
nor UO_3208 (O_3208,N_48362,N_49095);
xnor UO_3209 (O_3209,N_48742,N_48346);
or UO_3210 (O_3210,N_48657,N_49487);
and UO_3211 (O_3211,N_49477,N_48775);
nand UO_3212 (O_3212,N_48139,N_49795);
or UO_3213 (O_3213,N_48936,N_48823);
nand UO_3214 (O_3214,N_48820,N_48853);
or UO_3215 (O_3215,N_49365,N_48564);
nor UO_3216 (O_3216,N_48219,N_48962);
nor UO_3217 (O_3217,N_49556,N_48488);
nand UO_3218 (O_3218,N_48925,N_49596);
or UO_3219 (O_3219,N_49560,N_48514);
or UO_3220 (O_3220,N_48434,N_48050);
nand UO_3221 (O_3221,N_49325,N_49361);
xor UO_3222 (O_3222,N_48263,N_48528);
or UO_3223 (O_3223,N_49876,N_48441);
and UO_3224 (O_3224,N_49119,N_48497);
nor UO_3225 (O_3225,N_48692,N_48707);
xnor UO_3226 (O_3226,N_49209,N_48559);
xnor UO_3227 (O_3227,N_48389,N_49052);
nor UO_3228 (O_3228,N_49421,N_48057);
or UO_3229 (O_3229,N_48798,N_49034);
xnor UO_3230 (O_3230,N_49299,N_48889);
or UO_3231 (O_3231,N_48342,N_48734);
and UO_3232 (O_3232,N_49017,N_49367);
nor UO_3233 (O_3233,N_49501,N_49776);
nand UO_3234 (O_3234,N_49785,N_48243);
nand UO_3235 (O_3235,N_49058,N_48953);
and UO_3236 (O_3236,N_49281,N_48387);
nor UO_3237 (O_3237,N_49379,N_49158);
or UO_3238 (O_3238,N_49615,N_48318);
and UO_3239 (O_3239,N_48683,N_49905);
and UO_3240 (O_3240,N_49114,N_48796);
nor UO_3241 (O_3241,N_48627,N_49818);
and UO_3242 (O_3242,N_49239,N_49116);
or UO_3243 (O_3243,N_49404,N_48863);
or UO_3244 (O_3244,N_48793,N_49534);
nor UO_3245 (O_3245,N_48037,N_48731);
xor UO_3246 (O_3246,N_48398,N_48930);
nand UO_3247 (O_3247,N_48542,N_48638);
nor UO_3248 (O_3248,N_49430,N_48573);
and UO_3249 (O_3249,N_48873,N_48211);
nand UO_3250 (O_3250,N_49887,N_49540);
or UO_3251 (O_3251,N_49910,N_49290);
and UO_3252 (O_3252,N_48344,N_49124);
or UO_3253 (O_3253,N_48941,N_48736);
and UO_3254 (O_3254,N_49139,N_49959);
nor UO_3255 (O_3255,N_49663,N_49025);
nor UO_3256 (O_3256,N_48656,N_48540);
xnor UO_3257 (O_3257,N_48014,N_49667);
or UO_3258 (O_3258,N_49980,N_49687);
nor UO_3259 (O_3259,N_48949,N_48099);
and UO_3260 (O_3260,N_48116,N_48380);
or UO_3261 (O_3261,N_49349,N_48893);
and UO_3262 (O_3262,N_48602,N_49918);
xor UO_3263 (O_3263,N_48787,N_49436);
nand UO_3264 (O_3264,N_48390,N_48344);
or UO_3265 (O_3265,N_48910,N_49120);
and UO_3266 (O_3266,N_49682,N_48839);
and UO_3267 (O_3267,N_48858,N_49180);
nor UO_3268 (O_3268,N_48260,N_48763);
nor UO_3269 (O_3269,N_48610,N_49910);
xor UO_3270 (O_3270,N_49037,N_48019);
nand UO_3271 (O_3271,N_49279,N_49858);
and UO_3272 (O_3272,N_48661,N_49797);
nor UO_3273 (O_3273,N_48855,N_49913);
xnor UO_3274 (O_3274,N_49028,N_49887);
or UO_3275 (O_3275,N_49658,N_48429);
nor UO_3276 (O_3276,N_48251,N_49983);
or UO_3277 (O_3277,N_48052,N_48036);
xnor UO_3278 (O_3278,N_49170,N_48074);
or UO_3279 (O_3279,N_48528,N_48420);
or UO_3280 (O_3280,N_48419,N_49716);
xnor UO_3281 (O_3281,N_49519,N_49897);
and UO_3282 (O_3282,N_49933,N_49120);
nand UO_3283 (O_3283,N_48709,N_48202);
and UO_3284 (O_3284,N_48032,N_49604);
xnor UO_3285 (O_3285,N_49688,N_49262);
nand UO_3286 (O_3286,N_49316,N_49861);
nand UO_3287 (O_3287,N_48014,N_48393);
and UO_3288 (O_3288,N_49249,N_48553);
and UO_3289 (O_3289,N_48300,N_49562);
and UO_3290 (O_3290,N_49219,N_49210);
nor UO_3291 (O_3291,N_48143,N_49093);
or UO_3292 (O_3292,N_48784,N_49638);
nand UO_3293 (O_3293,N_49780,N_49702);
nor UO_3294 (O_3294,N_49284,N_49628);
or UO_3295 (O_3295,N_49136,N_48445);
xnor UO_3296 (O_3296,N_48796,N_49896);
nor UO_3297 (O_3297,N_48854,N_48960);
xnor UO_3298 (O_3298,N_48156,N_48596);
xor UO_3299 (O_3299,N_49700,N_49502);
or UO_3300 (O_3300,N_48302,N_48071);
xnor UO_3301 (O_3301,N_49399,N_48951);
or UO_3302 (O_3302,N_48215,N_49408);
nand UO_3303 (O_3303,N_48092,N_49596);
nand UO_3304 (O_3304,N_48199,N_48493);
or UO_3305 (O_3305,N_48125,N_49666);
and UO_3306 (O_3306,N_49094,N_49468);
nor UO_3307 (O_3307,N_49850,N_49018);
nand UO_3308 (O_3308,N_49803,N_48949);
nand UO_3309 (O_3309,N_48664,N_48591);
or UO_3310 (O_3310,N_49789,N_48635);
xor UO_3311 (O_3311,N_49137,N_49154);
nand UO_3312 (O_3312,N_49214,N_48196);
nand UO_3313 (O_3313,N_49766,N_49830);
or UO_3314 (O_3314,N_48926,N_48073);
and UO_3315 (O_3315,N_49813,N_48148);
or UO_3316 (O_3316,N_48575,N_48449);
or UO_3317 (O_3317,N_48780,N_48148);
and UO_3318 (O_3318,N_49693,N_48971);
xnor UO_3319 (O_3319,N_48370,N_49642);
or UO_3320 (O_3320,N_49048,N_48198);
nand UO_3321 (O_3321,N_48351,N_49468);
nand UO_3322 (O_3322,N_49384,N_49265);
xor UO_3323 (O_3323,N_49388,N_48222);
or UO_3324 (O_3324,N_48838,N_48067);
nor UO_3325 (O_3325,N_48944,N_49166);
nor UO_3326 (O_3326,N_49372,N_48389);
nor UO_3327 (O_3327,N_48180,N_49108);
xnor UO_3328 (O_3328,N_49576,N_48590);
nand UO_3329 (O_3329,N_48170,N_49431);
xnor UO_3330 (O_3330,N_49752,N_48353);
and UO_3331 (O_3331,N_48609,N_48749);
and UO_3332 (O_3332,N_48079,N_48832);
nor UO_3333 (O_3333,N_48684,N_49050);
or UO_3334 (O_3334,N_49028,N_48479);
and UO_3335 (O_3335,N_49117,N_49213);
or UO_3336 (O_3336,N_48827,N_49333);
xnor UO_3337 (O_3337,N_48357,N_49658);
xor UO_3338 (O_3338,N_48189,N_48807);
xnor UO_3339 (O_3339,N_48777,N_49249);
and UO_3340 (O_3340,N_49377,N_49618);
nand UO_3341 (O_3341,N_49234,N_48642);
nand UO_3342 (O_3342,N_48303,N_48989);
or UO_3343 (O_3343,N_49799,N_48092);
and UO_3344 (O_3344,N_48824,N_48749);
nand UO_3345 (O_3345,N_48120,N_49358);
nand UO_3346 (O_3346,N_48305,N_48820);
xnor UO_3347 (O_3347,N_48099,N_48100);
or UO_3348 (O_3348,N_49208,N_48659);
nor UO_3349 (O_3349,N_48300,N_48438);
xnor UO_3350 (O_3350,N_49089,N_49226);
or UO_3351 (O_3351,N_48332,N_49287);
nand UO_3352 (O_3352,N_49880,N_49870);
nand UO_3353 (O_3353,N_48612,N_49878);
nand UO_3354 (O_3354,N_48081,N_48660);
or UO_3355 (O_3355,N_49897,N_49195);
and UO_3356 (O_3356,N_48665,N_48407);
and UO_3357 (O_3357,N_49195,N_48851);
xnor UO_3358 (O_3358,N_49737,N_49840);
xor UO_3359 (O_3359,N_48141,N_48414);
xor UO_3360 (O_3360,N_49624,N_48668);
nand UO_3361 (O_3361,N_48656,N_49355);
xor UO_3362 (O_3362,N_49046,N_48963);
or UO_3363 (O_3363,N_48741,N_49881);
xor UO_3364 (O_3364,N_48213,N_48626);
xor UO_3365 (O_3365,N_48971,N_48493);
nor UO_3366 (O_3366,N_49011,N_48734);
xor UO_3367 (O_3367,N_48974,N_48447);
nor UO_3368 (O_3368,N_49370,N_48177);
xor UO_3369 (O_3369,N_48033,N_49739);
xor UO_3370 (O_3370,N_49406,N_48598);
nand UO_3371 (O_3371,N_49353,N_49847);
nor UO_3372 (O_3372,N_48305,N_49038);
xor UO_3373 (O_3373,N_48009,N_49379);
and UO_3374 (O_3374,N_49110,N_49610);
nand UO_3375 (O_3375,N_48254,N_49950);
nand UO_3376 (O_3376,N_49659,N_49522);
xnor UO_3377 (O_3377,N_49467,N_48588);
nor UO_3378 (O_3378,N_48147,N_48081);
and UO_3379 (O_3379,N_48638,N_48777);
xnor UO_3380 (O_3380,N_49790,N_48602);
xnor UO_3381 (O_3381,N_48208,N_48634);
or UO_3382 (O_3382,N_48702,N_48680);
or UO_3383 (O_3383,N_48596,N_49433);
xor UO_3384 (O_3384,N_48062,N_49726);
nand UO_3385 (O_3385,N_48988,N_49520);
or UO_3386 (O_3386,N_48687,N_49863);
and UO_3387 (O_3387,N_49609,N_49406);
xnor UO_3388 (O_3388,N_48598,N_48745);
nor UO_3389 (O_3389,N_48879,N_49687);
nand UO_3390 (O_3390,N_48206,N_48323);
and UO_3391 (O_3391,N_49337,N_49286);
or UO_3392 (O_3392,N_48706,N_49783);
or UO_3393 (O_3393,N_49872,N_49242);
and UO_3394 (O_3394,N_49544,N_49601);
nor UO_3395 (O_3395,N_49021,N_49291);
or UO_3396 (O_3396,N_49741,N_49499);
nand UO_3397 (O_3397,N_48728,N_48692);
nand UO_3398 (O_3398,N_48653,N_49003);
xnor UO_3399 (O_3399,N_48199,N_48733);
xor UO_3400 (O_3400,N_48695,N_49979);
nand UO_3401 (O_3401,N_49120,N_48268);
nor UO_3402 (O_3402,N_49132,N_49090);
and UO_3403 (O_3403,N_48473,N_49269);
nor UO_3404 (O_3404,N_49467,N_49353);
and UO_3405 (O_3405,N_49363,N_48418);
and UO_3406 (O_3406,N_48704,N_49599);
nor UO_3407 (O_3407,N_48791,N_48205);
or UO_3408 (O_3408,N_49014,N_48517);
xor UO_3409 (O_3409,N_49092,N_49555);
nand UO_3410 (O_3410,N_49993,N_48178);
and UO_3411 (O_3411,N_48384,N_49584);
nor UO_3412 (O_3412,N_48982,N_48918);
or UO_3413 (O_3413,N_48992,N_48933);
nor UO_3414 (O_3414,N_48542,N_49359);
xor UO_3415 (O_3415,N_48304,N_48550);
or UO_3416 (O_3416,N_48617,N_48632);
and UO_3417 (O_3417,N_49910,N_49621);
and UO_3418 (O_3418,N_48228,N_49483);
xor UO_3419 (O_3419,N_49039,N_49513);
nor UO_3420 (O_3420,N_49997,N_48678);
xor UO_3421 (O_3421,N_48169,N_49950);
xor UO_3422 (O_3422,N_48299,N_49867);
and UO_3423 (O_3423,N_49181,N_49302);
or UO_3424 (O_3424,N_48394,N_48595);
or UO_3425 (O_3425,N_49636,N_48691);
and UO_3426 (O_3426,N_48727,N_49794);
xnor UO_3427 (O_3427,N_49963,N_48403);
nor UO_3428 (O_3428,N_49517,N_49728);
nand UO_3429 (O_3429,N_49471,N_48019);
nor UO_3430 (O_3430,N_48998,N_49531);
or UO_3431 (O_3431,N_49292,N_48123);
and UO_3432 (O_3432,N_49038,N_48603);
xnor UO_3433 (O_3433,N_49266,N_48888);
xor UO_3434 (O_3434,N_48190,N_48136);
and UO_3435 (O_3435,N_49120,N_48431);
xnor UO_3436 (O_3436,N_48697,N_48310);
nor UO_3437 (O_3437,N_49187,N_48436);
xnor UO_3438 (O_3438,N_49807,N_49188);
nand UO_3439 (O_3439,N_49057,N_48443);
nor UO_3440 (O_3440,N_49244,N_49798);
xor UO_3441 (O_3441,N_49995,N_48312);
or UO_3442 (O_3442,N_48341,N_49723);
nand UO_3443 (O_3443,N_49052,N_48068);
nand UO_3444 (O_3444,N_49046,N_48174);
nor UO_3445 (O_3445,N_48499,N_49200);
or UO_3446 (O_3446,N_48941,N_48550);
nand UO_3447 (O_3447,N_49815,N_49224);
or UO_3448 (O_3448,N_49436,N_48793);
nor UO_3449 (O_3449,N_48018,N_48782);
and UO_3450 (O_3450,N_49400,N_48533);
nand UO_3451 (O_3451,N_48274,N_48425);
xor UO_3452 (O_3452,N_49799,N_49903);
nand UO_3453 (O_3453,N_48804,N_48275);
xnor UO_3454 (O_3454,N_48061,N_49650);
nor UO_3455 (O_3455,N_48552,N_49362);
xor UO_3456 (O_3456,N_49935,N_48589);
xor UO_3457 (O_3457,N_49387,N_49407);
xnor UO_3458 (O_3458,N_49300,N_49951);
nor UO_3459 (O_3459,N_49489,N_48885);
or UO_3460 (O_3460,N_49863,N_48560);
xor UO_3461 (O_3461,N_49865,N_49347);
xnor UO_3462 (O_3462,N_48340,N_48043);
nand UO_3463 (O_3463,N_49695,N_48130);
and UO_3464 (O_3464,N_48635,N_49085);
nand UO_3465 (O_3465,N_49545,N_49053);
and UO_3466 (O_3466,N_49096,N_49859);
nand UO_3467 (O_3467,N_48058,N_48096);
nor UO_3468 (O_3468,N_48569,N_49227);
xor UO_3469 (O_3469,N_49493,N_49185);
and UO_3470 (O_3470,N_49340,N_48397);
nand UO_3471 (O_3471,N_49386,N_49398);
nor UO_3472 (O_3472,N_49877,N_48342);
and UO_3473 (O_3473,N_48513,N_49122);
and UO_3474 (O_3474,N_48441,N_49119);
or UO_3475 (O_3475,N_49994,N_49966);
xor UO_3476 (O_3476,N_48012,N_49634);
and UO_3477 (O_3477,N_48489,N_48882);
xor UO_3478 (O_3478,N_48621,N_48023);
or UO_3479 (O_3479,N_49997,N_49281);
nor UO_3480 (O_3480,N_49100,N_49746);
xnor UO_3481 (O_3481,N_49126,N_49783);
nor UO_3482 (O_3482,N_49002,N_49613);
or UO_3483 (O_3483,N_49695,N_49700);
nand UO_3484 (O_3484,N_48026,N_48372);
and UO_3485 (O_3485,N_49290,N_48356);
xnor UO_3486 (O_3486,N_48917,N_49138);
or UO_3487 (O_3487,N_49999,N_49804);
and UO_3488 (O_3488,N_48327,N_48174);
and UO_3489 (O_3489,N_48822,N_49741);
nand UO_3490 (O_3490,N_49230,N_48498);
nor UO_3491 (O_3491,N_48913,N_48579);
and UO_3492 (O_3492,N_49012,N_49267);
and UO_3493 (O_3493,N_49435,N_49083);
nor UO_3494 (O_3494,N_49870,N_49420);
or UO_3495 (O_3495,N_48490,N_48263);
xnor UO_3496 (O_3496,N_48893,N_48745);
or UO_3497 (O_3497,N_49189,N_49342);
xor UO_3498 (O_3498,N_48434,N_49075);
nand UO_3499 (O_3499,N_49374,N_49770);
or UO_3500 (O_3500,N_49032,N_48826);
nand UO_3501 (O_3501,N_49274,N_48557);
xnor UO_3502 (O_3502,N_48786,N_49849);
nor UO_3503 (O_3503,N_48694,N_49180);
or UO_3504 (O_3504,N_48712,N_49671);
nor UO_3505 (O_3505,N_49430,N_49872);
xnor UO_3506 (O_3506,N_49095,N_49113);
and UO_3507 (O_3507,N_48283,N_48791);
or UO_3508 (O_3508,N_49800,N_49011);
nand UO_3509 (O_3509,N_49673,N_49755);
nand UO_3510 (O_3510,N_49697,N_49156);
or UO_3511 (O_3511,N_48071,N_49267);
xnor UO_3512 (O_3512,N_48879,N_48429);
and UO_3513 (O_3513,N_49977,N_48672);
nor UO_3514 (O_3514,N_49402,N_49245);
nand UO_3515 (O_3515,N_49947,N_49744);
or UO_3516 (O_3516,N_49807,N_49832);
and UO_3517 (O_3517,N_49840,N_49859);
nor UO_3518 (O_3518,N_49659,N_48186);
nor UO_3519 (O_3519,N_48060,N_48978);
xor UO_3520 (O_3520,N_48742,N_48285);
or UO_3521 (O_3521,N_48207,N_49516);
nand UO_3522 (O_3522,N_48910,N_48569);
and UO_3523 (O_3523,N_48119,N_49344);
xnor UO_3524 (O_3524,N_49530,N_48659);
nand UO_3525 (O_3525,N_48776,N_49896);
and UO_3526 (O_3526,N_48900,N_48537);
or UO_3527 (O_3527,N_48146,N_48271);
xor UO_3528 (O_3528,N_49002,N_48214);
xnor UO_3529 (O_3529,N_48644,N_49986);
or UO_3530 (O_3530,N_49650,N_49760);
and UO_3531 (O_3531,N_48640,N_49217);
or UO_3532 (O_3532,N_48795,N_48223);
xor UO_3533 (O_3533,N_48987,N_48506);
and UO_3534 (O_3534,N_49213,N_49903);
and UO_3535 (O_3535,N_48094,N_48163);
and UO_3536 (O_3536,N_48548,N_49793);
nand UO_3537 (O_3537,N_48260,N_48764);
or UO_3538 (O_3538,N_48489,N_49604);
or UO_3539 (O_3539,N_49475,N_49188);
xnor UO_3540 (O_3540,N_49729,N_49444);
or UO_3541 (O_3541,N_48917,N_49782);
nor UO_3542 (O_3542,N_49956,N_48813);
nand UO_3543 (O_3543,N_49376,N_49467);
nor UO_3544 (O_3544,N_48940,N_49767);
and UO_3545 (O_3545,N_49558,N_48014);
nand UO_3546 (O_3546,N_49286,N_49546);
and UO_3547 (O_3547,N_49001,N_49264);
and UO_3548 (O_3548,N_49270,N_48736);
xor UO_3549 (O_3549,N_48474,N_49947);
nor UO_3550 (O_3550,N_48872,N_48163);
xnor UO_3551 (O_3551,N_48509,N_49756);
nand UO_3552 (O_3552,N_49935,N_49839);
nand UO_3553 (O_3553,N_49596,N_48321);
nor UO_3554 (O_3554,N_48550,N_49127);
nand UO_3555 (O_3555,N_48162,N_48139);
and UO_3556 (O_3556,N_48486,N_49276);
or UO_3557 (O_3557,N_48068,N_49818);
or UO_3558 (O_3558,N_49311,N_49993);
nand UO_3559 (O_3559,N_49058,N_48181);
nor UO_3560 (O_3560,N_49873,N_49127);
and UO_3561 (O_3561,N_48710,N_48298);
and UO_3562 (O_3562,N_48223,N_49012);
nor UO_3563 (O_3563,N_49664,N_48941);
and UO_3564 (O_3564,N_49013,N_48007);
and UO_3565 (O_3565,N_49733,N_49056);
nor UO_3566 (O_3566,N_48079,N_48465);
nand UO_3567 (O_3567,N_48813,N_48538);
nor UO_3568 (O_3568,N_48935,N_49376);
nand UO_3569 (O_3569,N_48600,N_49366);
and UO_3570 (O_3570,N_49317,N_49121);
nand UO_3571 (O_3571,N_49596,N_48823);
and UO_3572 (O_3572,N_49006,N_48394);
nand UO_3573 (O_3573,N_48995,N_49135);
or UO_3574 (O_3574,N_48063,N_49686);
xor UO_3575 (O_3575,N_49415,N_48324);
nor UO_3576 (O_3576,N_49568,N_49578);
nand UO_3577 (O_3577,N_49620,N_49919);
nand UO_3578 (O_3578,N_48543,N_48177);
or UO_3579 (O_3579,N_48871,N_48265);
xnor UO_3580 (O_3580,N_48982,N_48969);
xor UO_3581 (O_3581,N_48341,N_49122);
or UO_3582 (O_3582,N_49074,N_48406);
and UO_3583 (O_3583,N_49924,N_49845);
nand UO_3584 (O_3584,N_48541,N_49270);
xor UO_3585 (O_3585,N_48558,N_49204);
or UO_3586 (O_3586,N_49135,N_48313);
xnor UO_3587 (O_3587,N_49391,N_49928);
and UO_3588 (O_3588,N_48714,N_48806);
and UO_3589 (O_3589,N_49882,N_49959);
nor UO_3590 (O_3590,N_48040,N_48211);
nor UO_3591 (O_3591,N_49234,N_48437);
or UO_3592 (O_3592,N_48731,N_48541);
and UO_3593 (O_3593,N_48942,N_49107);
xor UO_3594 (O_3594,N_49975,N_48724);
nor UO_3595 (O_3595,N_48155,N_48847);
nor UO_3596 (O_3596,N_48778,N_49532);
nand UO_3597 (O_3597,N_48736,N_48622);
xor UO_3598 (O_3598,N_49670,N_48269);
and UO_3599 (O_3599,N_48365,N_49581);
or UO_3600 (O_3600,N_49125,N_48509);
or UO_3601 (O_3601,N_49933,N_49591);
xor UO_3602 (O_3602,N_48285,N_48446);
and UO_3603 (O_3603,N_49106,N_49192);
nor UO_3604 (O_3604,N_48597,N_48658);
nor UO_3605 (O_3605,N_48254,N_48239);
or UO_3606 (O_3606,N_49235,N_49605);
nand UO_3607 (O_3607,N_49161,N_48012);
or UO_3608 (O_3608,N_49906,N_49496);
xor UO_3609 (O_3609,N_48092,N_49806);
or UO_3610 (O_3610,N_48616,N_48160);
nor UO_3611 (O_3611,N_48152,N_49232);
nand UO_3612 (O_3612,N_48801,N_48176);
nor UO_3613 (O_3613,N_49044,N_49465);
nor UO_3614 (O_3614,N_48330,N_49809);
or UO_3615 (O_3615,N_49601,N_49011);
xor UO_3616 (O_3616,N_49338,N_48898);
xnor UO_3617 (O_3617,N_48704,N_48994);
xnor UO_3618 (O_3618,N_49954,N_49346);
nand UO_3619 (O_3619,N_49245,N_48293);
nor UO_3620 (O_3620,N_49733,N_49815);
xnor UO_3621 (O_3621,N_49117,N_48451);
nor UO_3622 (O_3622,N_49724,N_48468);
nand UO_3623 (O_3623,N_49789,N_48476);
or UO_3624 (O_3624,N_48270,N_49463);
nand UO_3625 (O_3625,N_48117,N_49258);
nor UO_3626 (O_3626,N_48387,N_48912);
xor UO_3627 (O_3627,N_48245,N_48946);
xor UO_3628 (O_3628,N_49533,N_49090);
nor UO_3629 (O_3629,N_49032,N_49845);
nand UO_3630 (O_3630,N_49534,N_49932);
or UO_3631 (O_3631,N_49052,N_48154);
nand UO_3632 (O_3632,N_48058,N_49357);
nand UO_3633 (O_3633,N_48946,N_48641);
nand UO_3634 (O_3634,N_48848,N_48724);
or UO_3635 (O_3635,N_49952,N_48205);
nand UO_3636 (O_3636,N_48429,N_49817);
nand UO_3637 (O_3637,N_48345,N_49880);
xor UO_3638 (O_3638,N_48347,N_49177);
nand UO_3639 (O_3639,N_48968,N_49580);
or UO_3640 (O_3640,N_48011,N_49065);
nand UO_3641 (O_3641,N_48163,N_48115);
or UO_3642 (O_3642,N_49843,N_49386);
nand UO_3643 (O_3643,N_49046,N_49238);
and UO_3644 (O_3644,N_48461,N_49918);
xor UO_3645 (O_3645,N_49915,N_48605);
xnor UO_3646 (O_3646,N_48703,N_48784);
nand UO_3647 (O_3647,N_49467,N_48796);
or UO_3648 (O_3648,N_49366,N_49424);
nor UO_3649 (O_3649,N_48162,N_48645);
xor UO_3650 (O_3650,N_49103,N_49162);
nand UO_3651 (O_3651,N_48363,N_48006);
or UO_3652 (O_3652,N_48860,N_49490);
nand UO_3653 (O_3653,N_49464,N_48899);
xnor UO_3654 (O_3654,N_49462,N_49928);
and UO_3655 (O_3655,N_48345,N_48135);
nor UO_3656 (O_3656,N_49713,N_48603);
and UO_3657 (O_3657,N_49356,N_48670);
nor UO_3658 (O_3658,N_49444,N_48239);
nand UO_3659 (O_3659,N_48087,N_48121);
nand UO_3660 (O_3660,N_48562,N_48323);
nor UO_3661 (O_3661,N_48484,N_48054);
and UO_3662 (O_3662,N_48114,N_49379);
xor UO_3663 (O_3663,N_49002,N_48639);
and UO_3664 (O_3664,N_48347,N_49682);
or UO_3665 (O_3665,N_48040,N_49317);
or UO_3666 (O_3666,N_48605,N_49788);
or UO_3667 (O_3667,N_48224,N_48802);
or UO_3668 (O_3668,N_49966,N_49875);
or UO_3669 (O_3669,N_49228,N_49182);
nand UO_3670 (O_3670,N_48541,N_49075);
nor UO_3671 (O_3671,N_49493,N_48738);
nand UO_3672 (O_3672,N_49972,N_49502);
and UO_3673 (O_3673,N_48780,N_48486);
nand UO_3674 (O_3674,N_48085,N_49404);
nor UO_3675 (O_3675,N_49691,N_49425);
or UO_3676 (O_3676,N_48056,N_48741);
nor UO_3677 (O_3677,N_49686,N_48387);
xnor UO_3678 (O_3678,N_48333,N_48943);
and UO_3679 (O_3679,N_49831,N_48121);
and UO_3680 (O_3680,N_49392,N_49663);
nor UO_3681 (O_3681,N_49402,N_48903);
xor UO_3682 (O_3682,N_48005,N_49226);
xor UO_3683 (O_3683,N_48236,N_48412);
xor UO_3684 (O_3684,N_49774,N_48473);
nor UO_3685 (O_3685,N_48504,N_48161);
nand UO_3686 (O_3686,N_49870,N_48865);
xnor UO_3687 (O_3687,N_49024,N_49323);
or UO_3688 (O_3688,N_49581,N_49970);
and UO_3689 (O_3689,N_48136,N_48441);
nand UO_3690 (O_3690,N_48657,N_49821);
or UO_3691 (O_3691,N_48785,N_48279);
or UO_3692 (O_3692,N_49234,N_48169);
or UO_3693 (O_3693,N_49782,N_48462);
xnor UO_3694 (O_3694,N_48562,N_49951);
and UO_3695 (O_3695,N_49216,N_49318);
nor UO_3696 (O_3696,N_48435,N_48969);
nand UO_3697 (O_3697,N_48195,N_49005);
or UO_3698 (O_3698,N_49431,N_49926);
and UO_3699 (O_3699,N_49002,N_48645);
or UO_3700 (O_3700,N_49761,N_48892);
and UO_3701 (O_3701,N_48618,N_48473);
xnor UO_3702 (O_3702,N_49408,N_48831);
or UO_3703 (O_3703,N_49457,N_49390);
and UO_3704 (O_3704,N_49401,N_49302);
and UO_3705 (O_3705,N_49385,N_48463);
nand UO_3706 (O_3706,N_49838,N_49760);
and UO_3707 (O_3707,N_49213,N_49380);
nor UO_3708 (O_3708,N_48435,N_49787);
or UO_3709 (O_3709,N_48531,N_48154);
and UO_3710 (O_3710,N_49323,N_48285);
xor UO_3711 (O_3711,N_48032,N_49809);
or UO_3712 (O_3712,N_49106,N_48142);
and UO_3713 (O_3713,N_49374,N_49651);
or UO_3714 (O_3714,N_48695,N_49412);
and UO_3715 (O_3715,N_48993,N_49814);
and UO_3716 (O_3716,N_48579,N_49506);
nand UO_3717 (O_3717,N_49257,N_49986);
nand UO_3718 (O_3718,N_49497,N_48405);
or UO_3719 (O_3719,N_48306,N_49499);
and UO_3720 (O_3720,N_48139,N_49504);
xnor UO_3721 (O_3721,N_48482,N_48952);
xor UO_3722 (O_3722,N_49847,N_48290);
or UO_3723 (O_3723,N_48298,N_49041);
xnor UO_3724 (O_3724,N_48962,N_48380);
or UO_3725 (O_3725,N_48994,N_49607);
nand UO_3726 (O_3726,N_48745,N_49058);
xnor UO_3727 (O_3727,N_48209,N_48774);
and UO_3728 (O_3728,N_48141,N_49749);
xor UO_3729 (O_3729,N_48410,N_49239);
nor UO_3730 (O_3730,N_49097,N_48739);
xnor UO_3731 (O_3731,N_48508,N_49426);
and UO_3732 (O_3732,N_48606,N_49497);
nand UO_3733 (O_3733,N_49727,N_49949);
nand UO_3734 (O_3734,N_48319,N_49323);
and UO_3735 (O_3735,N_48926,N_48234);
and UO_3736 (O_3736,N_49015,N_49443);
nand UO_3737 (O_3737,N_48431,N_48922);
nor UO_3738 (O_3738,N_49259,N_48723);
nand UO_3739 (O_3739,N_48913,N_48149);
nor UO_3740 (O_3740,N_48650,N_49522);
nand UO_3741 (O_3741,N_48363,N_49326);
nand UO_3742 (O_3742,N_49657,N_49696);
xor UO_3743 (O_3743,N_49602,N_49022);
nor UO_3744 (O_3744,N_49946,N_48897);
xnor UO_3745 (O_3745,N_48931,N_48523);
nor UO_3746 (O_3746,N_49627,N_48763);
xnor UO_3747 (O_3747,N_49806,N_49467);
nor UO_3748 (O_3748,N_48482,N_48168);
nor UO_3749 (O_3749,N_49506,N_48402);
nor UO_3750 (O_3750,N_48221,N_48544);
xnor UO_3751 (O_3751,N_48220,N_49297);
nand UO_3752 (O_3752,N_48736,N_49305);
xor UO_3753 (O_3753,N_48226,N_49793);
nand UO_3754 (O_3754,N_48332,N_48191);
and UO_3755 (O_3755,N_48693,N_49557);
nand UO_3756 (O_3756,N_49716,N_48808);
or UO_3757 (O_3757,N_48149,N_48558);
and UO_3758 (O_3758,N_49418,N_48806);
or UO_3759 (O_3759,N_49059,N_48361);
xnor UO_3760 (O_3760,N_48542,N_48264);
and UO_3761 (O_3761,N_48132,N_49400);
xor UO_3762 (O_3762,N_49705,N_48473);
or UO_3763 (O_3763,N_48242,N_48837);
nor UO_3764 (O_3764,N_48212,N_49576);
or UO_3765 (O_3765,N_49502,N_49722);
and UO_3766 (O_3766,N_49649,N_48391);
nor UO_3767 (O_3767,N_48588,N_48922);
nand UO_3768 (O_3768,N_48187,N_49318);
and UO_3769 (O_3769,N_48976,N_48992);
and UO_3770 (O_3770,N_48539,N_48237);
nor UO_3771 (O_3771,N_49560,N_49348);
and UO_3772 (O_3772,N_49448,N_48372);
or UO_3773 (O_3773,N_48432,N_49234);
xor UO_3774 (O_3774,N_49365,N_48405);
nor UO_3775 (O_3775,N_49343,N_48740);
nand UO_3776 (O_3776,N_49533,N_49706);
or UO_3777 (O_3777,N_48025,N_49289);
nor UO_3778 (O_3778,N_49001,N_48353);
xnor UO_3779 (O_3779,N_49479,N_49827);
nor UO_3780 (O_3780,N_48344,N_48172);
nand UO_3781 (O_3781,N_48106,N_49018);
nor UO_3782 (O_3782,N_48863,N_49142);
and UO_3783 (O_3783,N_49949,N_48281);
and UO_3784 (O_3784,N_49846,N_49185);
nor UO_3785 (O_3785,N_49196,N_49324);
xnor UO_3786 (O_3786,N_49662,N_49852);
nand UO_3787 (O_3787,N_48168,N_49228);
xor UO_3788 (O_3788,N_48908,N_48461);
or UO_3789 (O_3789,N_49605,N_49563);
or UO_3790 (O_3790,N_49583,N_48167);
nand UO_3791 (O_3791,N_48968,N_49261);
and UO_3792 (O_3792,N_49376,N_49791);
nand UO_3793 (O_3793,N_49240,N_49207);
and UO_3794 (O_3794,N_48647,N_49518);
and UO_3795 (O_3795,N_49333,N_48232);
xor UO_3796 (O_3796,N_49619,N_49241);
xor UO_3797 (O_3797,N_48032,N_49131);
or UO_3798 (O_3798,N_48244,N_49362);
xnor UO_3799 (O_3799,N_48542,N_48408);
xnor UO_3800 (O_3800,N_48402,N_48056);
nand UO_3801 (O_3801,N_49862,N_49202);
nand UO_3802 (O_3802,N_49601,N_49836);
xnor UO_3803 (O_3803,N_49697,N_48445);
nor UO_3804 (O_3804,N_48158,N_49461);
nand UO_3805 (O_3805,N_48203,N_49712);
nor UO_3806 (O_3806,N_49871,N_48051);
nand UO_3807 (O_3807,N_49146,N_48942);
xor UO_3808 (O_3808,N_49747,N_48706);
and UO_3809 (O_3809,N_48406,N_49607);
nor UO_3810 (O_3810,N_49217,N_49368);
xnor UO_3811 (O_3811,N_49358,N_49934);
nand UO_3812 (O_3812,N_48432,N_48107);
xnor UO_3813 (O_3813,N_48560,N_48916);
xor UO_3814 (O_3814,N_48800,N_49343);
or UO_3815 (O_3815,N_48947,N_49171);
nor UO_3816 (O_3816,N_49890,N_48407);
xnor UO_3817 (O_3817,N_48565,N_49592);
or UO_3818 (O_3818,N_49511,N_48573);
and UO_3819 (O_3819,N_49648,N_49642);
nor UO_3820 (O_3820,N_49307,N_48149);
nor UO_3821 (O_3821,N_49300,N_48354);
nor UO_3822 (O_3822,N_48279,N_48274);
or UO_3823 (O_3823,N_49026,N_49321);
nor UO_3824 (O_3824,N_48313,N_49079);
nand UO_3825 (O_3825,N_49620,N_49825);
nor UO_3826 (O_3826,N_48115,N_49484);
xnor UO_3827 (O_3827,N_49138,N_48233);
nand UO_3828 (O_3828,N_49981,N_49795);
and UO_3829 (O_3829,N_49653,N_49200);
nand UO_3830 (O_3830,N_49492,N_48657);
nand UO_3831 (O_3831,N_48024,N_49380);
or UO_3832 (O_3832,N_48552,N_48608);
nand UO_3833 (O_3833,N_48289,N_48832);
nor UO_3834 (O_3834,N_49186,N_49936);
xnor UO_3835 (O_3835,N_48987,N_49252);
and UO_3836 (O_3836,N_49149,N_48266);
xor UO_3837 (O_3837,N_48987,N_48937);
nor UO_3838 (O_3838,N_48985,N_49155);
nor UO_3839 (O_3839,N_49378,N_49203);
or UO_3840 (O_3840,N_48111,N_48429);
or UO_3841 (O_3841,N_49597,N_49599);
and UO_3842 (O_3842,N_48379,N_48059);
nor UO_3843 (O_3843,N_48717,N_48386);
xor UO_3844 (O_3844,N_49643,N_48210);
or UO_3845 (O_3845,N_49765,N_48834);
nand UO_3846 (O_3846,N_48500,N_49291);
xor UO_3847 (O_3847,N_48631,N_48735);
xor UO_3848 (O_3848,N_48800,N_49991);
nand UO_3849 (O_3849,N_49161,N_48083);
and UO_3850 (O_3850,N_49528,N_49200);
or UO_3851 (O_3851,N_49305,N_49421);
or UO_3852 (O_3852,N_49018,N_49531);
nor UO_3853 (O_3853,N_49058,N_48431);
xnor UO_3854 (O_3854,N_48789,N_49710);
and UO_3855 (O_3855,N_48861,N_49861);
xor UO_3856 (O_3856,N_48670,N_48507);
nand UO_3857 (O_3857,N_48626,N_48351);
and UO_3858 (O_3858,N_49333,N_49484);
nor UO_3859 (O_3859,N_48363,N_49927);
nand UO_3860 (O_3860,N_49471,N_49207);
and UO_3861 (O_3861,N_48622,N_48110);
or UO_3862 (O_3862,N_49403,N_48731);
nor UO_3863 (O_3863,N_49986,N_48470);
xnor UO_3864 (O_3864,N_48997,N_48565);
or UO_3865 (O_3865,N_48010,N_48120);
and UO_3866 (O_3866,N_49125,N_49370);
and UO_3867 (O_3867,N_48404,N_49681);
xor UO_3868 (O_3868,N_48007,N_48448);
xor UO_3869 (O_3869,N_48874,N_48109);
and UO_3870 (O_3870,N_48014,N_49810);
xor UO_3871 (O_3871,N_48806,N_49690);
nor UO_3872 (O_3872,N_48473,N_48020);
and UO_3873 (O_3873,N_48445,N_48977);
nand UO_3874 (O_3874,N_49279,N_48941);
and UO_3875 (O_3875,N_49052,N_49445);
or UO_3876 (O_3876,N_49246,N_49487);
xnor UO_3877 (O_3877,N_48448,N_49956);
nor UO_3878 (O_3878,N_48976,N_49278);
nor UO_3879 (O_3879,N_49014,N_48537);
and UO_3880 (O_3880,N_49836,N_48917);
and UO_3881 (O_3881,N_49351,N_48870);
and UO_3882 (O_3882,N_48720,N_48848);
nand UO_3883 (O_3883,N_48219,N_49543);
nor UO_3884 (O_3884,N_48589,N_48332);
or UO_3885 (O_3885,N_49955,N_48020);
xor UO_3886 (O_3886,N_48020,N_49128);
nor UO_3887 (O_3887,N_49402,N_49699);
xnor UO_3888 (O_3888,N_48881,N_48986);
xnor UO_3889 (O_3889,N_48574,N_48066);
nand UO_3890 (O_3890,N_48273,N_49459);
nor UO_3891 (O_3891,N_49681,N_49042);
and UO_3892 (O_3892,N_48921,N_49684);
nor UO_3893 (O_3893,N_49614,N_48203);
xor UO_3894 (O_3894,N_49959,N_48741);
nor UO_3895 (O_3895,N_49270,N_48457);
nor UO_3896 (O_3896,N_49089,N_48519);
nor UO_3897 (O_3897,N_49455,N_49161);
nor UO_3898 (O_3898,N_48025,N_48485);
and UO_3899 (O_3899,N_48377,N_48913);
and UO_3900 (O_3900,N_48293,N_48044);
xnor UO_3901 (O_3901,N_48846,N_49428);
nand UO_3902 (O_3902,N_49520,N_48575);
xor UO_3903 (O_3903,N_48501,N_49673);
nor UO_3904 (O_3904,N_49298,N_49838);
xor UO_3905 (O_3905,N_48708,N_48232);
nor UO_3906 (O_3906,N_49843,N_49060);
and UO_3907 (O_3907,N_49970,N_49202);
nand UO_3908 (O_3908,N_49012,N_48282);
nand UO_3909 (O_3909,N_49184,N_49946);
or UO_3910 (O_3910,N_48783,N_48589);
or UO_3911 (O_3911,N_48473,N_48940);
nor UO_3912 (O_3912,N_48621,N_48145);
nor UO_3913 (O_3913,N_49701,N_49829);
or UO_3914 (O_3914,N_49054,N_49432);
nor UO_3915 (O_3915,N_48993,N_49568);
nor UO_3916 (O_3916,N_49928,N_49777);
xnor UO_3917 (O_3917,N_48775,N_48226);
nor UO_3918 (O_3918,N_49997,N_49789);
and UO_3919 (O_3919,N_48057,N_49910);
or UO_3920 (O_3920,N_48505,N_49533);
nand UO_3921 (O_3921,N_48142,N_49189);
nor UO_3922 (O_3922,N_49394,N_48066);
nand UO_3923 (O_3923,N_49348,N_48499);
or UO_3924 (O_3924,N_49550,N_49427);
xor UO_3925 (O_3925,N_49318,N_49958);
or UO_3926 (O_3926,N_48524,N_49921);
or UO_3927 (O_3927,N_48680,N_48736);
nor UO_3928 (O_3928,N_49807,N_49521);
xor UO_3929 (O_3929,N_48175,N_49790);
or UO_3930 (O_3930,N_49413,N_49276);
nor UO_3931 (O_3931,N_48907,N_48068);
xnor UO_3932 (O_3932,N_49424,N_49121);
nor UO_3933 (O_3933,N_49204,N_49101);
or UO_3934 (O_3934,N_48616,N_48780);
nor UO_3935 (O_3935,N_49654,N_48168);
nor UO_3936 (O_3936,N_48697,N_48046);
nand UO_3937 (O_3937,N_49275,N_49042);
xnor UO_3938 (O_3938,N_49680,N_49866);
nand UO_3939 (O_3939,N_48307,N_48783);
nand UO_3940 (O_3940,N_49620,N_48184);
nand UO_3941 (O_3941,N_49893,N_48607);
nor UO_3942 (O_3942,N_48392,N_49278);
or UO_3943 (O_3943,N_48718,N_49561);
nor UO_3944 (O_3944,N_49800,N_49138);
xnor UO_3945 (O_3945,N_49711,N_48235);
nand UO_3946 (O_3946,N_49748,N_48181);
or UO_3947 (O_3947,N_48043,N_49830);
and UO_3948 (O_3948,N_48493,N_49300);
and UO_3949 (O_3949,N_48886,N_48630);
or UO_3950 (O_3950,N_48385,N_49709);
nor UO_3951 (O_3951,N_49051,N_48129);
or UO_3952 (O_3952,N_48201,N_49929);
xor UO_3953 (O_3953,N_48906,N_49977);
nand UO_3954 (O_3954,N_48141,N_49134);
or UO_3955 (O_3955,N_49367,N_48204);
nand UO_3956 (O_3956,N_48448,N_49191);
nor UO_3957 (O_3957,N_48938,N_48283);
or UO_3958 (O_3958,N_49944,N_48510);
or UO_3959 (O_3959,N_48802,N_49984);
and UO_3960 (O_3960,N_48840,N_49691);
and UO_3961 (O_3961,N_49021,N_49402);
xnor UO_3962 (O_3962,N_48506,N_49400);
xnor UO_3963 (O_3963,N_48402,N_48113);
xnor UO_3964 (O_3964,N_49817,N_48946);
nand UO_3965 (O_3965,N_49441,N_49967);
nor UO_3966 (O_3966,N_49725,N_49630);
and UO_3967 (O_3967,N_48688,N_48142);
or UO_3968 (O_3968,N_49938,N_49688);
or UO_3969 (O_3969,N_48927,N_48594);
nand UO_3970 (O_3970,N_48623,N_48502);
nand UO_3971 (O_3971,N_49678,N_49980);
nor UO_3972 (O_3972,N_49237,N_49215);
or UO_3973 (O_3973,N_48985,N_48730);
xnor UO_3974 (O_3974,N_48729,N_49533);
or UO_3975 (O_3975,N_49594,N_49777);
or UO_3976 (O_3976,N_48914,N_48378);
and UO_3977 (O_3977,N_49593,N_48948);
and UO_3978 (O_3978,N_49441,N_48689);
or UO_3979 (O_3979,N_49028,N_48232);
nor UO_3980 (O_3980,N_48100,N_48379);
nor UO_3981 (O_3981,N_48330,N_49744);
xor UO_3982 (O_3982,N_49024,N_48163);
or UO_3983 (O_3983,N_49704,N_49285);
nor UO_3984 (O_3984,N_49490,N_48314);
xor UO_3985 (O_3985,N_48785,N_48412);
nand UO_3986 (O_3986,N_49488,N_48393);
nand UO_3987 (O_3987,N_49599,N_48563);
or UO_3988 (O_3988,N_49881,N_49704);
xnor UO_3989 (O_3989,N_49193,N_49283);
or UO_3990 (O_3990,N_49626,N_49514);
nand UO_3991 (O_3991,N_49260,N_48433);
xnor UO_3992 (O_3992,N_49456,N_49977);
and UO_3993 (O_3993,N_48392,N_48624);
xnor UO_3994 (O_3994,N_48555,N_48092);
nor UO_3995 (O_3995,N_49938,N_49645);
or UO_3996 (O_3996,N_48803,N_48454);
and UO_3997 (O_3997,N_48892,N_49924);
nand UO_3998 (O_3998,N_49217,N_49762);
nand UO_3999 (O_3999,N_48084,N_49699);
xor UO_4000 (O_4000,N_49922,N_48521);
and UO_4001 (O_4001,N_49501,N_49137);
nor UO_4002 (O_4002,N_48063,N_48854);
nand UO_4003 (O_4003,N_49744,N_48457);
nor UO_4004 (O_4004,N_48689,N_49871);
nor UO_4005 (O_4005,N_48257,N_48361);
and UO_4006 (O_4006,N_48175,N_49570);
nor UO_4007 (O_4007,N_48263,N_48219);
and UO_4008 (O_4008,N_48228,N_49432);
or UO_4009 (O_4009,N_49713,N_49091);
nor UO_4010 (O_4010,N_49398,N_49845);
and UO_4011 (O_4011,N_48353,N_49848);
nor UO_4012 (O_4012,N_49832,N_49283);
nand UO_4013 (O_4013,N_48717,N_49849);
nand UO_4014 (O_4014,N_48283,N_48810);
and UO_4015 (O_4015,N_49123,N_49239);
and UO_4016 (O_4016,N_49766,N_48761);
nor UO_4017 (O_4017,N_48691,N_49000);
and UO_4018 (O_4018,N_49772,N_49433);
or UO_4019 (O_4019,N_49557,N_49891);
nand UO_4020 (O_4020,N_49661,N_48540);
nand UO_4021 (O_4021,N_49266,N_48538);
or UO_4022 (O_4022,N_49188,N_48128);
nand UO_4023 (O_4023,N_49149,N_48670);
and UO_4024 (O_4024,N_49466,N_49059);
nor UO_4025 (O_4025,N_49740,N_48131);
nand UO_4026 (O_4026,N_48985,N_49015);
nor UO_4027 (O_4027,N_48005,N_48048);
nor UO_4028 (O_4028,N_48153,N_48365);
and UO_4029 (O_4029,N_49188,N_49943);
and UO_4030 (O_4030,N_49097,N_48923);
nand UO_4031 (O_4031,N_49415,N_48395);
or UO_4032 (O_4032,N_49990,N_48446);
xnor UO_4033 (O_4033,N_49936,N_48880);
or UO_4034 (O_4034,N_49181,N_49378);
nand UO_4035 (O_4035,N_49082,N_49148);
and UO_4036 (O_4036,N_48814,N_48730);
nor UO_4037 (O_4037,N_49176,N_49752);
or UO_4038 (O_4038,N_48765,N_48987);
nor UO_4039 (O_4039,N_48710,N_49897);
nor UO_4040 (O_4040,N_48875,N_49820);
xnor UO_4041 (O_4041,N_49865,N_48918);
xor UO_4042 (O_4042,N_48099,N_49089);
xor UO_4043 (O_4043,N_48120,N_49357);
nand UO_4044 (O_4044,N_48668,N_49928);
xnor UO_4045 (O_4045,N_48302,N_48762);
and UO_4046 (O_4046,N_48791,N_48688);
nand UO_4047 (O_4047,N_49475,N_48159);
nand UO_4048 (O_4048,N_48154,N_48167);
or UO_4049 (O_4049,N_48173,N_49534);
or UO_4050 (O_4050,N_49267,N_48955);
and UO_4051 (O_4051,N_49078,N_49956);
or UO_4052 (O_4052,N_48204,N_49177);
or UO_4053 (O_4053,N_49248,N_49531);
nor UO_4054 (O_4054,N_48494,N_49310);
or UO_4055 (O_4055,N_49595,N_48437);
or UO_4056 (O_4056,N_49957,N_48113);
nor UO_4057 (O_4057,N_48496,N_48125);
and UO_4058 (O_4058,N_49316,N_49318);
or UO_4059 (O_4059,N_48925,N_48122);
nand UO_4060 (O_4060,N_48673,N_49127);
and UO_4061 (O_4061,N_48189,N_48282);
and UO_4062 (O_4062,N_48581,N_48505);
xnor UO_4063 (O_4063,N_49512,N_48683);
or UO_4064 (O_4064,N_49081,N_48045);
nor UO_4065 (O_4065,N_49128,N_49872);
xnor UO_4066 (O_4066,N_48509,N_49854);
or UO_4067 (O_4067,N_49360,N_49085);
nand UO_4068 (O_4068,N_48187,N_48347);
xor UO_4069 (O_4069,N_49621,N_49648);
nand UO_4070 (O_4070,N_48756,N_49555);
nor UO_4071 (O_4071,N_48381,N_48843);
xor UO_4072 (O_4072,N_48041,N_48403);
and UO_4073 (O_4073,N_49193,N_49123);
or UO_4074 (O_4074,N_49214,N_48122);
and UO_4075 (O_4075,N_49461,N_48293);
nor UO_4076 (O_4076,N_48443,N_49041);
nor UO_4077 (O_4077,N_49684,N_48844);
xor UO_4078 (O_4078,N_48286,N_49010);
xnor UO_4079 (O_4079,N_49312,N_49202);
xor UO_4080 (O_4080,N_48373,N_49330);
nor UO_4081 (O_4081,N_49753,N_48552);
or UO_4082 (O_4082,N_49601,N_49051);
nor UO_4083 (O_4083,N_49581,N_48984);
nand UO_4084 (O_4084,N_49461,N_49039);
xnor UO_4085 (O_4085,N_49097,N_49446);
or UO_4086 (O_4086,N_49855,N_48497);
and UO_4087 (O_4087,N_49445,N_48579);
xor UO_4088 (O_4088,N_49692,N_48819);
or UO_4089 (O_4089,N_49028,N_48585);
xor UO_4090 (O_4090,N_49127,N_49210);
nand UO_4091 (O_4091,N_49653,N_49168);
nand UO_4092 (O_4092,N_48371,N_48290);
or UO_4093 (O_4093,N_48338,N_48423);
nand UO_4094 (O_4094,N_48298,N_48850);
or UO_4095 (O_4095,N_49792,N_49197);
xor UO_4096 (O_4096,N_49397,N_48640);
or UO_4097 (O_4097,N_49693,N_49920);
and UO_4098 (O_4098,N_49141,N_48488);
nor UO_4099 (O_4099,N_49775,N_49361);
and UO_4100 (O_4100,N_48067,N_48223);
nand UO_4101 (O_4101,N_49794,N_49982);
nor UO_4102 (O_4102,N_49318,N_49507);
or UO_4103 (O_4103,N_48476,N_48332);
xor UO_4104 (O_4104,N_48477,N_48432);
and UO_4105 (O_4105,N_49661,N_49855);
nor UO_4106 (O_4106,N_48463,N_49782);
nor UO_4107 (O_4107,N_49074,N_49718);
nand UO_4108 (O_4108,N_48793,N_48904);
or UO_4109 (O_4109,N_49699,N_48010);
xnor UO_4110 (O_4110,N_48776,N_48854);
or UO_4111 (O_4111,N_49805,N_48443);
or UO_4112 (O_4112,N_49873,N_49316);
and UO_4113 (O_4113,N_48978,N_48534);
nand UO_4114 (O_4114,N_48373,N_48223);
xor UO_4115 (O_4115,N_49142,N_48765);
xnor UO_4116 (O_4116,N_48744,N_49987);
or UO_4117 (O_4117,N_49126,N_48731);
nand UO_4118 (O_4118,N_49408,N_49316);
or UO_4119 (O_4119,N_48720,N_48141);
nand UO_4120 (O_4120,N_48621,N_49859);
or UO_4121 (O_4121,N_49686,N_48123);
and UO_4122 (O_4122,N_48106,N_48665);
xor UO_4123 (O_4123,N_48301,N_49159);
or UO_4124 (O_4124,N_48717,N_49815);
or UO_4125 (O_4125,N_49191,N_49560);
nor UO_4126 (O_4126,N_48939,N_48678);
and UO_4127 (O_4127,N_49849,N_49779);
xor UO_4128 (O_4128,N_48043,N_48808);
nor UO_4129 (O_4129,N_49775,N_49750);
nor UO_4130 (O_4130,N_48750,N_49941);
or UO_4131 (O_4131,N_48417,N_48191);
and UO_4132 (O_4132,N_48636,N_48483);
xnor UO_4133 (O_4133,N_48780,N_48397);
or UO_4134 (O_4134,N_48414,N_49978);
and UO_4135 (O_4135,N_48675,N_49322);
nand UO_4136 (O_4136,N_48677,N_48617);
or UO_4137 (O_4137,N_49990,N_49095);
and UO_4138 (O_4138,N_49219,N_48478);
and UO_4139 (O_4139,N_49955,N_49568);
nand UO_4140 (O_4140,N_48816,N_49734);
and UO_4141 (O_4141,N_49205,N_49705);
nor UO_4142 (O_4142,N_48655,N_49743);
and UO_4143 (O_4143,N_49690,N_49473);
nand UO_4144 (O_4144,N_49274,N_48363);
and UO_4145 (O_4145,N_48960,N_49709);
and UO_4146 (O_4146,N_49710,N_49206);
xnor UO_4147 (O_4147,N_48102,N_49027);
and UO_4148 (O_4148,N_48261,N_49436);
or UO_4149 (O_4149,N_49145,N_49179);
or UO_4150 (O_4150,N_49578,N_48069);
nor UO_4151 (O_4151,N_49366,N_48909);
nand UO_4152 (O_4152,N_48583,N_49386);
nand UO_4153 (O_4153,N_49401,N_49921);
or UO_4154 (O_4154,N_49390,N_48234);
and UO_4155 (O_4155,N_48975,N_48591);
or UO_4156 (O_4156,N_48209,N_49991);
nand UO_4157 (O_4157,N_49386,N_49879);
nor UO_4158 (O_4158,N_49256,N_48824);
nor UO_4159 (O_4159,N_48145,N_48029);
or UO_4160 (O_4160,N_49375,N_49001);
or UO_4161 (O_4161,N_49641,N_49138);
nor UO_4162 (O_4162,N_49792,N_49401);
xnor UO_4163 (O_4163,N_48708,N_49458);
nor UO_4164 (O_4164,N_49921,N_48086);
and UO_4165 (O_4165,N_48963,N_49725);
or UO_4166 (O_4166,N_49013,N_48098);
nor UO_4167 (O_4167,N_48276,N_48282);
or UO_4168 (O_4168,N_49380,N_48947);
or UO_4169 (O_4169,N_48867,N_49412);
or UO_4170 (O_4170,N_49697,N_48472);
and UO_4171 (O_4171,N_49706,N_49223);
or UO_4172 (O_4172,N_49069,N_48689);
nor UO_4173 (O_4173,N_49904,N_49258);
nand UO_4174 (O_4174,N_49202,N_48323);
and UO_4175 (O_4175,N_48651,N_49038);
and UO_4176 (O_4176,N_48588,N_48600);
and UO_4177 (O_4177,N_48464,N_49209);
or UO_4178 (O_4178,N_49348,N_49554);
xor UO_4179 (O_4179,N_49339,N_49267);
or UO_4180 (O_4180,N_49237,N_48115);
nand UO_4181 (O_4181,N_49939,N_48126);
or UO_4182 (O_4182,N_49807,N_48226);
nand UO_4183 (O_4183,N_48306,N_49370);
or UO_4184 (O_4184,N_49282,N_48863);
nor UO_4185 (O_4185,N_48804,N_49834);
xnor UO_4186 (O_4186,N_49598,N_48883);
nor UO_4187 (O_4187,N_48719,N_49984);
or UO_4188 (O_4188,N_48458,N_49102);
and UO_4189 (O_4189,N_48230,N_49583);
xnor UO_4190 (O_4190,N_49362,N_49019);
xor UO_4191 (O_4191,N_48351,N_49062);
and UO_4192 (O_4192,N_48814,N_48425);
and UO_4193 (O_4193,N_49542,N_49410);
nand UO_4194 (O_4194,N_49540,N_48860);
and UO_4195 (O_4195,N_48196,N_49393);
nand UO_4196 (O_4196,N_48779,N_48125);
xor UO_4197 (O_4197,N_48315,N_48790);
and UO_4198 (O_4198,N_48064,N_48744);
and UO_4199 (O_4199,N_48862,N_48150);
nor UO_4200 (O_4200,N_48380,N_48124);
or UO_4201 (O_4201,N_49622,N_48987);
or UO_4202 (O_4202,N_48999,N_48460);
and UO_4203 (O_4203,N_48930,N_48102);
xnor UO_4204 (O_4204,N_49541,N_48192);
nand UO_4205 (O_4205,N_49515,N_48303);
or UO_4206 (O_4206,N_49143,N_48741);
nand UO_4207 (O_4207,N_48805,N_48189);
and UO_4208 (O_4208,N_49236,N_48719);
nand UO_4209 (O_4209,N_48580,N_48460);
xnor UO_4210 (O_4210,N_49220,N_49576);
xor UO_4211 (O_4211,N_48262,N_49075);
xnor UO_4212 (O_4212,N_49147,N_48953);
nor UO_4213 (O_4213,N_48246,N_48819);
and UO_4214 (O_4214,N_49132,N_49442);
or UO_4215 (O_4215,N_49782,N_49096);
xor UO_4216 (O_4216,N_48896,N_49236);
xnor UO_4217 (O_4217,N_49635,N_49139);
and UO_4218 (O_4218,N_49289,N_49759);
or UO_4219 (O_4219,N_48928,N_49946);
or UO_4220 (O_4220,N_49168,N_48673);
xor UO_4221 (O_4221,N_48902,N_49096);
and UO_4222 (O_4222,N_49189,N_49901);
nor UO_4223 (O_4223,N_49075,N_48783);
or UO_4224 (O_4224,N_49911,N_49154);
and UO_4225 (O_4225,N_48610,N_48493);
nand UO_4226 (O_4226,N_49958,N_48397);
nor UO_4227 (O_4227,N_49010,N_49876);
nor UO_4228 (O_4228,N_49794,N_49934);
xor UO_4229 (O_4229,N_48526,N_49418);
xnor UO_4230 (O_4230,N_48322,N_48402);
or UO_4231 (O_4231,N_48936,N_49674);
or UO_4232 (O_4232,N_48271,N_48747);
and UO_4233 (O_4233,N_49405,N_49000);
and UO_4234 (O_4234,N_49606,N_49155);
nor UO_4235 (O_4235,N_48025,N_48813);
nand UO_4236 (O_4236,N_49179,N_49150);
or UO_4237 (O_4237,N_49547,N_49705);
nand UO_4238 (O_4238,N_49326,N_48702);
nor UO_4239 (O_4239,N_49948,N_49017);
nor UO_4240 (O_4240,N_49905,N_48976);
nor UO_4241 (O_4241,N_48375,N_48314);
and UO_4242 (O_4242,N_49274,N_48166);
or UO_4243 (O_4243,N_49595,N_48547);
nand UO_4244 (O_4244,N_49522,N_49510);
nor UO_4245 (O_4245,N_49611,N_48621);
or UO_4246 (O_4246,N_48542,N_49221);
and UO_4247 (O_4247,N_48503,N_48868);
nand UO_4248 (O_4248,N_48069,N_48789);
or UO_4249 (O_4249,N_49234,N_48816);
and UO_4250 (O_4250,N_49050,N_49236);
xnor UO_4251 (O_4251,N_48355,N_48962);
nand UO_4252 (O_4252,N_48047,N_49313);
xor UO_4253 (O_4253,N_49997,N_49305);
xor UO_4254 (O_4254,N_49497,N_48876);
and UO_4255 (O_4255,N_49228,N_48037);
or UO_4256 (O_4256,N_48209,N_48553);
or UO_4257 (O_4257,N_49324,N_49202);
or UO_4258 (O_4258,N_48923,N_48524);
or UO_4259 (O_4259,N_49225,N_48627);
and UO_4260 (O_4260,N_48437,N_48383);
xor UO_4261 (O_4261,N_48969,N_49047);
nand UO_4262 (O_4262,N_49781,N_49999);
nor UO_4263 (O_4263,N_49409,N_49596);
nand UO_4264 (O_4264,N_48414,N_48957);
nor UO_4265 (O_4265,N_48374,N_48878);
and UO_4266 (O_4266,N_48438,N_48459);
nand UO_4267 (O_4267,N_48719,N_49126);
xnor UO_4268 (O_4268,N_48633,N_48284);
nor UO_4269 (O_4269,N_49967,N_49634);
nand UO_4270 (O_4270,N_48142,N_49302);
nand UO_4271 (O_4271,N_49845,N_48824);
or UO_4272 (O_4272,N_48143,N_48502);
or UO_4273 (O_4273,N_48081,N_48160);
nor UO_4274 (O_4274,N_49519,N_49244);
or UO_4275 (O_4275,N_49068,N_49724);
nor UO_4276 (O_4276,N_49026,N_49770);
nand UO_4277 (O_4277,N_49979,N_48302);
nand UO_4278 (O_4278,N_48879,N_48393);
nand UO_4279 (O_4279,N_48330,N_49697);
or UO_4280 (O_4280,N_49670,N_48715);
nand UO_4281 (O_4281,N_49309,N_49004);
or UO_4282 (O_4282,N_49847,N_49966);
or UO_4283 (O_4283,N_49323,N_49592);
nor UO_4284 (O_4284,N_48183,N_49598);
or UO_4285 (O_4285,N_48766,N_49147);
nand UO_4286 (O_4286,N_49993,N_48238);
and UO_4287 (O_4287,N_48684,N_49080);
nor UO_4288 (O_4288,N_48058,N_48633);
or UO_4289 (O_4289,N_48252,N_49505);
and UO_4290 (O_4290,N_49861,N_48284);
xnor UO_4291 (O_4291,N_48161,N_49708);
nor UO_4292 (O_4292,N_49077,N_49093);
xnor UO_4293 (O_4293,N_49377,N_48425);
xor UO_4294 (O_4294,N_48981,N_49828);
xnor UO_4295 (O_4295,N_48588,N_48047);
nor UO_4296 (O_4296,N_49438,N_49307);
nand UO_4297 (O_4297,N_49636,N_49154);
nand UO_4298 (O_4298,N_49153,N_49076);
nor UO_4299 (O_4299,N_48649,N_48905);
nand UO_4300 (O_4300,N_49098,N_48719);
nand UO_4301 (O_4301,N_48319,N_48041);
nand UO_4302 (O_4302,N_48986,N_49382);
xnor UO_4303 (O_4303,N_48509,N_48097);
or UO_4304 (O_4304,N_49936,N_48268);
nor UO_4305 (O_4305,N_49642,N_49327);
nor UO_4306 (O_4306,N_49561,N_48410);
and UO_4307 (O_4307,N_49141,N_48501);
and UO_4308 (O_4308,N_49531,N_48222);
nor UO_4309 (O_4309,N_48202,N_48329);
nand UO_4310 (O_4310,N_48691,N_49995);
nor UO_4311 (O_4311,N_48412,N_49588);
xnor UO_4312 (O_4312,N_48854,N_48492);
nand UO_4313 (O_4313,N_48883,N_49029);
and UO_4314 (O_4314,N_48289,N_48606);
and UO_4315 (O_4315,N_49551,N_48969);
xnor UO_4316 (O_4316,N_49049,N_49008);
nor UO_4317 (O_4317,N_48930,N_48925);
and UO_4318 (O_4318,N_48875,N_49795);
xor UO_4319 (O_4319,N_48771,N_49528);
xnor UO_4320 (O_4320,N_49099,N_48921);
xor UO_4321 (O_4321,N_48181,N_49811);
nor UO_4322 (O_4322,N_49301,N_49936);
and UO_4323 (O_4323,N_48656,N_49183);
nor UO_4324 (O_4324,N_48647,N_49166);
nor UO_4325 (O_4325,N_49309,N_49250);
nand UO_4326 (O_4326,N_49723,N_49348);
xnor UO_4327 (O_4327,N_48024,N_49847);
xnor UO_4328 (O_4328,N_48520,N_49943);
or UO_4329 (O_4329,N_49393,N_49452);
xor UO_4330 (O_4330,N_48608,N_48546);
or UO_4331 (O_4331,N_49624,N_49843);
nor UO_4332 (O_4332,N_48339,N_49087);
xnor UO_4333 (O_4333,N_48414,N_49955);
xnor UO_4334 (O_4334,N_49288,N_49384);
and UO_4335 (O_4335,N_49352,N_48206);
nor UO_4336 (O_4336,N_48702,N_48325);
xnor UO_4337 (O_4337,N_49775,N_48651);
and UO_4338 (O_4338,N_48792,N_48536);
xor UO_4339 (O_4339,N_48706,N_49120);
nor UO_4340 (O_4340,N_48660,N_49697);
and UO_4341 (O_4341,N_49438,N_49576);
xor UO_4342 (O_4342,N_49907,N_48078);
nor UO_4343 (O_4343,N_49014,N_49494);
nand UO_4344 (O_4344,N_48353,N_48343);
xnor UO_4345 (O_4345,N_48662,N_48408);
xnor UO_4346 (O_4346,N_48723,N_49057);
nand UO_4347 (O_4347,N_49086,N_49853);
and UO_4348 (O_4348,N_48580,N_49805);
nor UO_4349 (O_4349,N_49746,N_49551);
or UO_4350 (O_4350,N_48502,N_49670);
xor UO_4351 (O_4351,N_49367,N_49266);
nor UO_4352 (O_4352,N_49529,N_49656);
or UO_4353 (O_4353,N_48764,N_48220);
and UO_4354 (O_4354,N_49802,N_49525);
or UO_4355 (O_4355,N_49405,N_49616);
nand UO_4356 (O_4356,N_48528,N_49947);
and UO_4357 (O_4357,N_48472,N_49074);
nand UO_4358 (O_4358,N_49217,N_49130);
xnor UO_4359 (O_4359,N_48550,N_49427);
nand UO_4360 (O_4360,N_49423,N_48032);
or UO_4361 (O_4361,N_48454,N_49026);
or UO_4362 (O_4362,N_49715,N_48725);
and UO_4363 (O_4363,N_49137,N_49227);
and UO_4364 (O_4364,N_48040,N_48453);
and UO_4365 (O_4365,N_48201,N_48023);
nand UO_4366 (O_4366,N_48332,N_48463);
nor UO_4367 (O_4367,N_48468,N_48840);
nor UO_4368 (O_4368,N_48829,N_48405);
xnor UO_4369 (O_4369,N_48327,N_49791);
nand UO_4370 (O_4370,N_49663,N_49544);
and UO_4371 (O_4371,N_49261,N_49284);
xnor UO_4372 (O_4372,N_49362,N_49198);
or UO_4373 (O_4373,N_48395,N_48893);
nor UO_4374 (O_4374,N_49813,N_49565);
nand UO_4375 (O_4375,N_49817,N_48438);
or UO_4376 (O_4376,N_49110,N_48532);
xnor UO_4377 (O_4377,N_49755,N_49109);
nand UO_4378 (O_4378,N_49513,N_48119);
or UO_4379 (O_4379,N_48941,N_49475);
nand UO_4380 (O_4380,N_48861,N_48576);
nor UO_4381 (O_4381,N_48253,N_48063);
nor UO_4382 (O_4382,N_49544,N_48666);
and UO_4383 (O_4383,N_48782,N_48146);
xor UO_4384 (O_4384,N_49700,N_48823);
xor UO_4385 (O_4385,N_49788,N_48701);
nand UO_4386 (O_4386,N_49310,N_48232);
xor UO_4387 (O_4387,N_48843,N_49015);
or UO_4388 (O_4388,N_49018,N_48229);
or UO_4389 (O_4389,N_48656,N_48307);
or UO_4390 (O_4390,N_48615,N_48117);
and UO_4391 (O_4391,N_48413,N_49307);
nor UO_4392 (O_4392,N_49864,N_48438);
nand UO_4393 (O_4393,N_48932,N_48113);
xnor UO_4394 (O_4394,N_48571,N_49684);
or UO_4395 (O_4395,N_49501,N_48435);
nor UO_4396 (O_4396,N_49655,N_49449);
nor UO_4397 (O_4397,N_49813,N_49387);
xor UO_4398 (O_4398,N_48913,N_48070);
and UO_4399 (O_4399,N_48054,N_48052);
or UO_4400 (O_4400,N_49109,N_49050);
nand UO_4401 (O_4401,N_48125,N_48185);
nor UO_4402 (O_4402,N_49253,N_49390);
or UO_4403 (O_4403,N_48236,N_49024);
or UO_4404 (O_4404,N_49729,N_48310);
and UO_4405 (O_4405,N_49866,N_49718);
nor UO_4406 (O_4406,N_48506,N_49830);
and UO_4407 (O_4407,N_49767,N_49173);
and UO_4408 (O_4408,N_49893,N_49977);
nor UO_4409 (O_4409,N_48389,N_48039);
nor UO_4410 (O_4410,N_48060,N_48529);
nand UO_4411 (O_4411,N_48744,N_49548);
and UO_4412 (O_4412,N_48873,N_48916);
nor UO_4413 (O_4413,N_48678,N_48258);
or UO_4414 (O_4414,N_49336,N_49815);
xor UO_4415 (O_4415,N_48641,N_49454);
xnor UO_4416 (O_4416,N_48145,N_48483);
or UO_4417 (O_4417,N_49171,N_49607);
xnor UO_4418 (O_4418,N_48218,N_49801);
nor UO_4419 (O_4419,N_49592,N_49058);
nor UO_4420 (O_4420,N_49733,N_49404);
nand UO_4421 (O_4421,N_48784,N_48369);
or UO_4422 (O_4422,N_48047,N_49346);
or UO_4423 (O_4423,N_49856,N_48850);
or UO_4424 (O_4424,N_48480,N_49088);
nor UO_4425 (O_4425,N_49561,N_48079);
and UO_4426 (O_4426,N_48386,N_48892);
and UO_4427 (O_4427,N_49308,N_48675);
and UO_4428 (O_4428,N_48379,N_48425);
and UO_4429 (O_4429,N_48435,N_48211);
and UO_4430 (O_4430,N_49848,N_48959);
nor UO_4431 (O_4431,N_48740,N_49712);
nor UO_4432 (O_4432,N_48688,N_49830);
or UO_4433 (O_4433,N_48739,N_49507);
and UO_4434 (O_4434,N_48456,N_48656);
nor UO_4435 (O_4435,N_48531,N_48905);
or UO_4436 (O_4436,N_48960,N_48545);
xnor UO_4437 (O_4437,N_49894,N_48949);
and UO_4438 (O_4438,N_49988,N_48404);
and UO_4439 (O_4439,N_49832,N_49699);
and UO_4440 (O_4440,N_48137,N_49897);
nand UO_4441 (O_4441,N_48961,N_49703);
or UO_4442 (O_4442,N_48124,N_48505);
and UO_4443 (O_4443,N_48633,N_49358);
or UO_4444 (O_4444,N_48024,N_49188);
nand UO_4445 (O_4445,N_48660,N_49184);
nand UO_4446 (O_4446,N_48748,N_49062);
nor UO_4447 (O_4447,N_49367,N_48703);
and UO_4448 (O_4448,N_48679,N_49215);
or UO_4449 (O_4449,N_49265,N_48708);
and UO_4450 (O_4450,N_48787,N_48502);
nand UO_4451 (O_4451,N_49722,N_49521);
nor UO_4452 (O_4452,N_49173,N_49973);
nand UO_4453 (O_4453,N_48275,N_48012);
xor UO_4454 (O_4454,N_49662,N_48767);
and UO_4455 (O_4455,N_48449,N_49605);
nand UO_4456 (O_4456,N_48413,N_49202);
nand UO_4457 (O_4457,N_48118,N_48944);
xor UO_4458 (O_4458,N_48671,N_48451);
nand UO_4459 (O_4459,N_49980,N_49677);
nor UO_4460 (O_4460,N_49264,N_48102);
nand UO_4461 (O_4461,N_49939,N_49185);
nor UO_4462 (O_4462,N_49713,N_48664);
nor UO_4463 (O_4463,N_49472,N_49933);
or UO_4464 (O_4464,N_48968,N_48717);
xnor UO_4465 (O_4465,N_49911,N_48262);
and UO_4466 (O_4466,N_49033,N_49924);
and UO_4467 (O_4467,N_49393,N_49837);
nor UO_4468 (O_4468,N_49058,N_48444);
and UO_4469 (O_4469,N_49945,N_49914);
nor UO_4470 (O_4470,N_49473,N_49375);
nor UO_4471 (O_4471,N_48005,N_49138);
xor UO_4472 (O_4472,N_49694,N_49293);
and UO_4473 (O_4473,N_49785,N_49858);
and UO_4474 (O_4474,N_49809,N_49151);
nand UO_4475 (O_4475,N_48589,N_49818);
or UO_4476 (O_4476,N_48349,N_48951);
xnor UO_4477 (O_4477,N_49841,N_48581);
nor UO_4478 (O_4478,N_48454,N_49308);
or UO_4479 (O_4479,N_48829,N_48159);
nor UO_4480 (O_4480,N_49273,N_49262);
or UO_4481 (O_4481,N_48584,N_49716);
or UO_4482 (O_4482,N_49530,N_49891);
nand UO_4483 (O_4483,N_49361,N_49751);
xnor UO_4484 (O_4484,N_48786,N_49736);
nor UO_4485 (O_4485,N_49254,N_49809);
xor UO_4486 (O_4486,N_48215,N_49205);
xnor UO_4487 (O_4487,N_49194,N_48800);
nand UO_4488 (O_4488,N_49110,N_48139);
nand UO_4489 (O_4489,N_48816,N_49945);
nor UO_4490 (O_4490,N_49025,N_48083);
or UO_4491 (O_4491,N_48975,N_49912);
nor UO_4492 (O_4492,N_49511,N_49374);
xor UO_4493 (O_4493,N_49263,N_48664);
xnor UO_4494 (O_4494,N_48540,N_49844);
or UO_4495 (O_4495,N_49602,N_48104);
xor UO_4496 (O_4496,N_49656,N_49674);
nor UO_4497 (O_4497,N_48855,N_49463);
xor UO_4498 (O_4498,N_49016,N_48587);
or UO_4499 (O_4499,N_48789,N_48525);
nand UO_4500 (O_4500,N_48746,N_49665);
or UO_4501 (O_4501,N_49010,N_49485);
nor UO_4502 (O_4502,N_49624,N_48677);
nand UO_4503 (O_4503,N_49173,N_49692);
or UO_4504 (O_4504,N_48931,N_48128);
nand UO_4505 (O_4505,N_48369,N_49027);
and UO_4506 (O_4506,N_49270,N_48630);
nor UO_4507 (O_4507,N_48472,N_48531);
nand UO_4508 (O_4508,N_49351,N_49234);
nor UO_4509 (O_4509,N_49251,N_48929);
xnor UO_4510 (O_4510,N_48282,N_48100);
nor UO_4511 (O_4511,N_48953,N_48937);
nor UO_4512 (O_4512,N_48535,N_48120);
nand UO_4513 (O_4513,N_48686,N_49320);
or UO_4514 (O_4514,N_49503,N_49469);
xnor UO_4515 (O_4515,N_48889,N_49055);
nand UO_4516 (O_4516,N_48007,N_48804);
or UO_4517 (O_4517,N_49376,N_49702);
xor UO_4518 (O_4518,N_48076,N_49492);
and UO_4519 (O_4519,N_49611,N_48422);
xnor UO_4520 (O_4520,N_49420,N_49422);
and UO_4521 (O_4521,N_48070,N_49783);
nand UO_4522 (O_4522,N_48228,N_49588);
nand UO_4523 (O_4523,N_49893,N_48818);
or UO_4524 (O_4524,N_49566,N_49908);
or UO_4525 (O_4525,N_49166,N_48423);
and UO_4526 (O_4526,N_48691,N_49398);
or UO_4527 (O_4527,N_49331,N_49488);
xnor UO_4528 (O_4528,N_48193,N_49906);
or UO_4529 (O_4529,N_49829,N_49229);
and UO_4530 (O_4530,N_48959,N_49963);
xor UO_4531 (O_4531,N_49248,N_48799);
nor UO_4532 (O_4532,N_49278,N_49485);
or UO_4533 (O_4533,N_48230,N_49121);
nand UO_4534 (O_4534,N_49070,N_49935);
and UO_4535 (O_4535,N_49618,N_49407);
and UO_4536 (O_4536,N_48752,N_48181);
nor UO_4537 (O_4537,N_49074,N_49731);
nor UO_4538 (O_4538,N_49438,N_48680);
xor UO_4539 (O_4539,N_49649,N_48055);
xnor UO_4540 (O_4540,N_48772,N_48673);
and UO_4541 (O_4541,N_49193,N_48944);
xor UO_4542 (O_4542,N_49690,N_48479);
xor UO_4543 (O_4543,N_48159,N_49575);
and UO_4544 (O_4544,N_48594,N_49618);
nor UO_4545 (O_4545,N_48951,N_48158);
or UO_4546 (O_4546,N_48398,N_49842);
or UO_4547 (O_4547,N_48946,N_49031);
nor UO_4548 (O_4548,N_49497,N_49375);
or UO_4549 (O_4549,N_49669,N_48635);
xor UO_4550 (O_4550,N_48058,N_48032);
or UO_4551 (O_4551,N_48876,N_49928);
xnor UO_4552 (O_4552,N_48652,N_48367);
xnor UO_4553 (O_4553,N_48773,N_49292);
or UO_4554 (O_4554,N_48015,N_48537);
xor UO_4555 (O_4555,N_48218,N_49734);
and UO_4556 (O_4556,N_49487,N_49360);
xnor UO_4557 (O_4557,N_49662,N_49385);
and UO_4558 (O_4558,N_48819,N_48024);
or UO_4559 (O_4559,N_49875,N_49958);
nor UO_4560 (O_4560,N_49521,N_49826);
or UO_4561 (O_4561,N_49612,N_49927);
and UO_4562 (O_4562,N_48523,N_49125);
nor UO_4563 (O_4563,N_48265,N_49527);
nand UO_4564 (O_4564,N_48294,N_49143);
and UO_4565 (O_4565,N_49549,N_48134);
or UO_4566 (O_4566,N_49272,N_48233);
and UO_4567 (O_4567,N_48389,N_49704);
nand UO_4568 (O_4568,N_48083,N_48322);
nor UO_4569 (O_4569,N_48487,N_48100);
or UO_4570 (O_4570,N_49247,N_49753);
nor UO_4571 (O_4571,N_48644,N_48524);
nand UO_4572 (O_4572,N_49371,N_49564);
nor UO_4573 (O_4573,N_49588,N_48287);
nand UO_4574 (O_4574,N_49572,N_49548);
nand UO_4575 (O_4575,N_48743,N_49658);
xnor UO_4576 (O_4576,N_48675,N_49863);
or UO_4577 (O_4577,N_49655,N_48314);
nor UO_4578 (O_4578,N_48636,N_48447);
nand UO_4579 (O_4579,N_48250,N_49136);
or UO_4580 (O_4580,N_49585,N_48981);
xnor UO_4581 (O_4581,N_49242,N_49258);
or UO_4582 (O_4582,N_48646,N_49426);
and UO_4583 (O_4583,N_48414,N_48334);
nand UO_4584 (O_4584,N_49174,N_49965);
nand UO_4585 (O_4585,N_49692,N_49413);
or UO_4586 (O_4586,N_49525,N_49597);
or UO_4587 (O_4587,N_49720,N_48779);
nand UO_4588 (O_4588,N_48773,N_48420);
xor UO_4589 (O_4589,N_49005,N_48241);
nand UO_4590 (O_4590,N_48044,N_48611);
xnor UO_4591 (O_4591,N_49629,N_48017);
or UO_4592 (O_4592,N_48504,N_49827);
and UO_4593 (O_4593,N_48592,N_48307);
xnor UO_4594 (O_4594,N_49285,N_48629);
xnor UO_4595 (O_4595,N_49160,N_48144);
nand UO_4596 (O_4596,N_49531,N_48609);
or UO_4597 (O_4597,N_49346,N_48159);
or UO_4598 (O_4598,N_48065,N_49778);
xor UO_4599 (O_4599,N_49628,N_48860);
and UO_4600 (O_4600,N_48647,N_49425);
xor UO_4601 (O_4601,N_48083,N_48781);
xnor UO_4602 (O_4602,N_48007,N_49111);
and UO_4603 (O_4603,N_49516,N_48143);
nand UO_4604 (O_4604,N_48268,N_49106);
or UO_4605 (O_4605,N_49561,N_48055);
or UO_4606 (O_4606,N_48297,N_49055);
xnor UO_4607 (O_4607,N_49214,N_49401);
or UO_4608 (O_4608,N_49166,N_49236);
xnor UO_4609 (O_4609,N_49591,N_49529);
or UO_4610 (O_4610,N_48471,N_48240);
nand UO_4611 (O_4611,N_49427,N_49973);
nor UO_4612 (O_4612,N_48178,N_49257);
nand UO_4613 (O_4613,N_49043,N_48749);
nor UO_4614 (O_4614,N_48074,N_49651);
and UO_4615 (O_4615,N_49587,N_49784);
xor UO_4616 (O_4616,N_49590,N_48564);
xor UO_4617 (O_4617,N_49355,N_49626);
xor UO_4618 (O_4618,N_48519,N_49260);
or UO_4619 (O_4619,N_49051,N_48026);
and UO_4620 (O_4620,N_48646,N_48005);
xnor UO_4621 (O_4621,N_48810,N_48944);
nor UO_4622 (O_4622,N_48450,N_49653);
nor UO_4623 (O_4623,N_49110,N_49019);
nand UO_4624 (O_4624,N_48303,N_48305);
nor UO_4625 (O_4625,N_48713,N_48675);
or UO_4626 (O_4626,N_48439,N_48082);
nor UO_4627 (O_4627,N_49530,N_49468);
nand UO_4628 (O_4628,N_49085,N_48157);
and UO_4629 (O_4629,N_49388,N_48903);
and UO_4630 (O_4630,N_48917,N_48579);
or UO_4631 (O_4631,N_48162,N_48170);
xnor UO_4632 (O_4632,N_49161,N_49384);
xor UO_4633 (O_4633,N_48394,N_48856);
xnor UO_4634 (O_4634,N_48911,N_48233);
nor UO_4635 (O_4635,N_48295,N_48956);
or UO_4636 (O_4636,N_48015,N_48213);
nor UO_4637 (O_4637,N_48148,N_49760);
xor UO_4638 (O_4638,N_49496,N_48175);
or UO_4639 (O_4639,N_48225,N_49059);
and UO_4640 (O_4640,N_48154,N_49133);
and UO_4641 (O_4641,N_49037,N_48522);
or UO_4642 (O_4642,N_49007,N_49024);
nor UO_4643 (O_4643,N_48567,N_48925);
nor UO_4644 (O_4644,N_49668,N_49364);
and UO_4645 (O_4645,N_48331,N_49009);
nand UO_4646 (O_4646,N_48602,N_48599);
nor UO_4647 (O_4647,N_49620,N_49423);
nor UO_4648 (O_4648,N_49098,N_49118);
xor UO_4649 (O_4649,N_48239,N_49901);
and UO_4650 (O_4650,N_49294,N_48667);
nor UO_4651 (O_4651,N_49946,N_49548);
or UO_4652 (O_4652,N_49305,N_48130);
and UO_4653 (O_4653,N_49709,N_49914);
and UO_4654 (O_4654,N_49769,N_49748);
nor UO_4655 (O_4655,N_49055,N_48388);
xor UO_4656 (O_4656,N_48049,N_48701);
xnor UO_4657 (O_4657,N_49978,N_48788);
or UO_4658 (O_4658,N_48740,N_49324);
and UO_4659 (O_4659,N_49908,N_49006);
or UO_4660 (O_4660,N_49202,N_49577);
xnor UO_4661 (O_4661,N_48206,N_48337);
or UO_4662 (O_4662,N_49346,N_49892);
xor UO_4663 (O_4663,N_48066,N_48074);
or UO_4664 (O_4664,N_48967,N_49605);
nand UO_4665 (O_4665,N_49577,N_49548);
nand UO_4666 (O_4666,N_48910,N_49506);
and UO_4667 (O_4667,N_48873,N_48654);
xnor UO_4668 (O_4668,N_48990,N_48291);
xnor UO_4669 (O_4669,N_49339,N_49390);
xor UO_4670 (O_4670,N_49747,N_49594);
xor UO_4671 (O_4671,N_48460,N_48135);
and UO_4672 (O_4672,N_49945,N_48645);
or UO_4673 (O_4673,N_49027,N_48432);
or UO_4674 (O_4674,N_49482,N_48195);
or UO_4675 (O_4675,N_48446,N_48573);
nand UO_4676 (O_4676,N_49049,N_48449);
nor UO_4677 (O_4677,N_49585,N_49711);
nor UO_4678 (O_4678,N_49652,N_49807);
nand UO_4679 (O_4679,N_48668,N_49469);
nor UO_4680 (O_4680,N_48801,N_48803);
or UO_4681 (O_4681,N_49810,N_49762);
nor UO_4682 (O_4682,N_49595,N_48405);
nand UO_4683 (O_4683,N_49377,N_49089);
xor UO_4684 (O_4684,N_49674,N_48243);
nand UO_4685 (O_4685,N_49502,N_49049);
xnor UO_4686 (O_4686,N_48428,N_49095);
nand UO_4687 (O_4687,N_49219,N_48935);
nor UO_4688 (O_4688,N_48081,N_48326);
and UO_4689 (O_4689,N_48315,N_49980);
or UO_4690 (O_4690,N_49244,N_48922);
nor UO_4691 (O_4691,N_48498,N_49695);
xor UO_4692 (O_4692,N_49974,N_48173);
xor UO_4693 (O_4693,N_48264,N_48922);
nor UO_4694 (O_4694,N_48960,N_49802);
and UO_4695 (O_4695,N_48084,N_48699);
and UO_4696 (O_4696,N_49432,N_48003);
xor UO_4697 (O_4697,N_48552,N_48567);
nand UO_4698 (O_4698,N_48042,N_49432);
nor UO_4699 (O_4699,N_49478,N_49900);
nor UO_4700 (O_4700,N_49175,N_48944);
xor UO_4701 (O_4701,N_49846,N_49841);
nor UO_4702 (O_4702,N_48302,N_49172);
xor UO_4703 (O_4703,N_48035,N_49355);
nor UO_4704 (O_4704,N_49481,N_48637);
or UO_4705 (O_4705,N_49635,N_48723);
nand UO_4706 (O_4706,N_48618,N_49644);
nand UO_4707 (O_4707,N_49518,N_49893);
and UO_4708 (O_4708,N_48191,N_48988);
nand UO_4709 (O_4709,N_48605,N_49134);
nand UO_4710 (O_4710,N_49164,N_48276);
nor UO_4711 (O_4711,N_48566,N_48875);
nor UO_4712 (O_4712,N_48295,N_49913);
or UO_4713 (O_4713,N_49616,N_48835);
nor UO_4714 (O_4714,N_48762,N_48372);
and UO_4715 (O_4715,N_49735,N_48804);
nand UO_4716 (O_4716,N_49431,N_48971);
nand UO_4717 (O_4717,N_49644,N_48005);
xnor UO_4718 (O_4718,N_49142,N_48860);
and UO_4719 (O_4719,N_49612,N_49761);
xnor UO_4720 (O_4720,N_49516,N_48421);
or UO_4721 (O_4721,N_49075,N_48071);
nand UO_4722 (O_4722,N_48889,N_48146);
nor UO_4723 (O_4723,N_48393,N_48543);
and UO_4724 (O_4724,N_49117,N_49423);
nand UO_4725 (O_4725,N_48431,N_49391);
nor UO_4726 (O_4726,N_48852,N_48085);
nand UO_4727 (O_4727,N_48909,N_48254);
nand UO_4728 (O_4728,N_48552,N_48494);
and UO_4729 (O_4729,N_49550,N_48442);
or UO_4730 (O_4730,N_49445,N_49969);
and UO_4731 (O_4731,N_48915,N_48102);
xor UO_4732 (O_4732,N_48824,N_48173);
xor UO_4733 (O_4733,N_48685,N_49281);
and UO_4734 (O_4734,N_49537,N_49493);
nor UO_4735 (O_4735,N_49325,N_48214);
nor UO_4736 (O_4736,N_48858,N_48618);
nor UO_4737 (O_4737,N_49181,N_48126);
nor UO_4738 (O_4738,N_49446,N_48530);
nand UO_4739 (O_4739,N_48997,N_48102);
or UO_4740 (O_4740,N_48261,N_49258);
xnor UO_4741 (O_4741,N_49800,N_49936);
or UO_4742 (O_4742,N_49851,N_48095);
nand UO_4743 (O_4743,N_48219,N_49899);
and UO_4744 (O_4744,N_48704,N_49965);
or UO_4745 (O_4745,N_49803,N_48552);
or UO_4746 (O_4746,N_48764,N_49044);
and UO_4747 (O_4747,N_48590,N_48637);
xor UO_4748 (O_4748,N_48119,N_49071);
nand UO_4749 (O_4749,N_49278,N_49912);
nor UO_4750 (O_4750,N_49577,N_49171);
nand UO_4751 (O_4751,N_48385,N_48854);
or UO_4752 (O_4752,N_49460,N_49677);
and UO_4753 (O_4753,N_48411,N_49173);
xor UO_4754 (O_4754,N_48706,N_49317);
nor UO_4755 (O_4755,N_48113,N_48108);
or UO_4756 (O_4756,N_48863,N_48085);
nor UO_4757 (O_4757,N_49894,N_49542);
xor UO_4758 (O_4758,N_48639,N_48939);
xnor UO_4759 (O_4759,N_48905,N_48693);
and UO_4760 (O_4760,N_49991,N_48829);
nor UO_4761 (O_4761,N_48603,N_48818);
and UO_4762 (O_4762,N_49042,N_48084);
and UO_4763 (O_4763,N_49719,N_49905);
xor UO_4764 (O_4764,N_49957,N_49540);
xor UO_4765 (O_4765,N_48680,N_49497);
xnor UO_4766 (O_4766,N_49727,N_48805);
xnor UO_4767 (O_4767,N_49739,N_48608);
nor UO_4768 (O_4768,N_49914,N_48418);
or UO_4769 (O_4769,N_49859,N_48767);
nand UO_4770 (O_4770,N_48599,N_48526);
and UO_4771 (O_4771,N_49177,N_48564);
xor UO_4772 (O_4772,N_48082,N_49114);
nand UO_4773 (O_4773,N_48497,N_48620);
and UO_4774 (O_4774,N_49120,N_49292);
or UO_4775 (O_4775,N_48836,N_49648);
nand UO_4776 (O_4776,N_49985,N_48670);
or UO_4777 (O_4777,N_49162,N_48408);
nand UO_4778 (O_4778,N_49701,N_48872);
nand UO_4779 (O_4779,N_49689,N_48194);
nor UO_4780 (O_4780,N_49942,N_49370);
or UO_4781 (O_4781,N_49759,N_49225);
or UO_4782 (O_4782,N_48538,N_49771);
nor UO_4783 (O_4783,N_49634,N_48934);
nor UO_4784 (O_4784,N_49052,N_48463);
xnor UO_4785 (O_4785,N_49519,N_48641);
or UO_4786 (O_4786,N_48326,N_49908);
nand UO_4787 (O_4787,N_48995,N_48290);
and UO_4788 (O_4788,N_49153,N_49854);
or UO_4789 (O_4789,N_48342,N_48350);
xor UO_4790 (O_4790,N_49824,N_49696);
nand UO_4791 (O_4791,N_48147,N_49933);
nor UO_4792 (O_4792,N_48883,N_49627);
and UO_4793 (O_4793,N_48209,N_49014);
or UO_4794 (O_4794,N_48879,N_48726);
nand UO_4795 (O_4795,N_48144,N_48958);
nor UO_4796 (O_4796,N_49461,N_49704);
and UO_4797 (O_4797,N_49745,N_48219);
nand UO_4798 (O_4798,N_48675,N_48931);
or UO_4799 (O_4799,N_49142,N_49024);
xor UO_4800 (O_4800,N_48728,N_48290);
or UO_4801 (O_4801,N_48257,N_48988);
xor UO_4802 (O_4802,N_48506,N_49470);
or UO_4803 (O_4803,N_49188,N_49676);
nand UO_4804 (O_4804,N_48610,N_48226);
nand UO_4805 (O_4805,N_48400,N_48662);
xor UO_4806 (O_4806,N_48942,N_49379);
xor UO_4807 (O_4807,N_48334,N_49393);
and UO_4808 (O_4808,N_49692,N_49984);
or UO_4809 (O_4809,N_48776,N_49171);
nor UO_4810 (O_4810,N_48715,N_48523);
xor UO_4811 (O_4811,N_48860,N_49295);
nand UO_4812 (O_4812,N_48242,N_49295);
nand UO_4813 (O_4813,N_48457,N_49570);
xnor UO_4814 (O_4814,N_48181,N_49005);
xnor UO_4815 (O_4815,N_49187,N_49549);
nor UO_4816 (O_4816,N_49837,N_49074);
or UO_4817 (O_4817,N_48688,N_49411);
xor UO_4818 (O_4818,N_49378,N_48735);
or UO_4819 (O_4819,N_48311,N_48946);
or UO_4820 (O_4820,N_49981,N_48522);
xnor UO_4821 (O_4821,N_48599,N_49816);
and UO_4822 (O_4822,N_48654,N_48730);
and UO_4823 (O_4823,N_49379,N_49230);
nor UO_4824 (O_4824,N_48180,N_48541);
nor UO_4825 (O_4825,N_48356,N_48709);
nor UO_4826 (O_4826,N_48858,N_49224);
nand UO_4827 (O_4827,N_48307,N_48896);
nor UO_4828 (O_4828,N_49642,N_49190);
nor UO_4829 (O_4829,N_48756,N_48309);
and UO_4830 (O_4830,N_49460,N_48385);
xor UO_4831 (O_4831,N_48396,N_49544);
xnor UO_4832 (O_4832,N_48039,N_49409);
or UO_4833 (O_4833,N_49184,N_48052);
nand UO_4834 (O_4834,N_49519,N_49388);
or UO_4835 (O_4835,N_49406,N_48429);
or UO_4836 (O_4836,N_49350,N_49923);
or UO_4837 (O_4837,N_49323,N_48491);
and UO_4838 (O_4838,N_48406,N_49042);
xor UO_4839 (O_4839,N_48680,N_48521);
nor UO_4840 (O_4840,N_48877,N_49216);
nand UO_4841 (O_4841,N_49672,N_49189);
xor UO_4842 (O_4842,N_49013,N_48525);
or UO_4843 (O_4843,N_49682,N_49254);
nand UO_4844 (O_4844,N_48055,N_48994);
and UO_4845 (O_4845,N_48602,N_48506);
and UO_4846 (O_4846,N_49503,N_49033);
nand UO_4847 (O_4847,N_49174,N_49010);
nor UO_4848 (O_4848,N_48108,N_49853);
or UO_4849 (O_4849,N_48378,N_49606);
or UO_4850 (O_4850,N_48778,N_48356);
nand UO_4851 (O_4851,N_48436,N_49612);
nor UO_4852 (O_4852,N_48443,N_48783);
and UO_4853 (O_4853,N_49730,N_49449);
nand UO_4854 (O_4854,N_48748,N_48864);
nor UO_4855 (O_4855,N_49699,N_49230);
xnor UO_4856 (O_4856,N_49832,N_48038);
nand UO_4857 (O_4857,N_48966,N_48621);
and UO_4858 (O_4858,N_49261,N_49344);
and UO_4859 (O_4859,N_48023,N_49125);
xnor UO_4860 (O_4860,N_48661,N_48690);
xor UO_4861 (O_4861,N_49837,N_48759);
and UO_4862 (O_4862,N_49294,N_49016);
xor UO_4863 (O_4863,N_48798,N_48780);
nand UO_4864 (O_4864,N_48613,N_48847);
or UO_4865 (O_4865,N_49255,N_49509);
nor UO_4866 (O_4866,N_48912,N_49823);
or UO_4867 (O_4867,N_49211,N_48695);
nand UO_4868 (O_4868,N_49070,N_49150);
xor UO_4869 (O_4869,N_49989,N_48168);
xnor UO_4870 (O_4870,N_49729,N_48255);
nor UO_4871 (O_4871,N_48286,N_48173);
or UO_4872 (O_4872,N_49659,N_48698);
or UO_4873 (O_4873,N_48120,N_48405);
and UO_4874 (O_4874,N_48804,N_49956);
nand UO_4875 (O_4875,N_48188,N_49477);
nand UO_4876 (O_4876,N_48523,N_49974);
nand UO_4877 (O_4877,N_49771,N_48808);
or UO_4878 (O_4878,N_49941,N_49600);
xor UO_4879 (O_4879,N_49269,N_49993);
xor UO_4880 (O_4880,N_48868,N_49780);
or UO_4881 (O_4881,N_49907,N_49175);
nor UO_4882 (O_4882,N_49731,N_49382);
and UO_4883 (O_4883,N_49513,N_48735);
or UO_4884 (O_4884,N_49052,N_49458);
or UO_4885 (O_4885,N_48819,N_49117);
nor UO_4886 (O_4886,N_48500,N_49837);
or UO_4887 (O_4887,N_49301,N_49912);
or UO_4888 (O_4888,N_49116,N_49683);
nand UO_4889 (O_4889,N_48871,N_49365);
and UO_4890 (O_4890,N_49182,N_48188);
xor UO_4891 (O_4891,N_49705,N_49714);
or UO_4892 (O_4892,N_48158,N_49213);
xnor UO_4893 (O_4893,N_49606,N_49262);
and UO_4894 (O_4894,N_48378,N_49556);
and UO_4895 (O_4895,N_48617,N_49786);
nor UO_4896 (O_4896,N_48818,N_49923);
or UO_4897 (O_4897,N_48829,N_49359);
and UO_4898 (O_4898,N_48862,N_48619);
or UO_4899 (O_4899,N_49709,N_48363);
xor UO_4900 (O_4900,N_49065,N_49780);
xnor UO_4901 (O_4901,N_49928,N_49912);
xor UO_4902 (O_4902,N_48627,N_49645);
and UO_4903 (O_4903,N_49796,N_49723);
or UO_4904 (O_4904,N_48797,N_49842);
and UO_4905 (O_4905,N_48147,N_48394);
and UO_4906 (O_4906,N_48191,N_48183);
nor UO_4907 (O_4907,N_49929,N_48933);
and UO_4908 (O_4908,N_48704,N_49704);
nor UO_4909 (O_4909,N_49226,N_48707);
nand UO_4910 (O_4910,N_48136,N_49615);
nand UO_4911 (O_4911,N_49788,N_48606);
nand UO_4912 (O_4912,N_49586,N_49659);
xnor UO_4913 (O_4913,N_48918,N_49246);
xor UO_4914 (O_4914,N_49342,N_49356);
and UO_4915 (O_4915,N_48444,N_49581);
nor UO_4916 (O_4916,N_49085,N_49779);
nor UO_4917 (O_4917,N_49529,N_48148);
nand UO_4918 (O_4918,N_48285,N_49037);
and UO_4919 (O_4919,N_49354,N_49515);
xnor UO_4920 (O_4920,N_48881,N_48973);
xnor UO_4921 (O_4921,N_49830,N_49907);
nor UO_4922 (O_4922,N_48085,N_49810);
nor UO_4923 (O_4923,N_48007,N_49648);
xor UO_4924 (O_4924,N_48571,N_48438);
and UO_4925 (O_4925,N_49228,N_48674);
and UO_4926 (O_4926,N_49402,N_48901);
nand UO_4927 (O_4927,N_48148,N_48081);
or UO_4928 (O_4928,N_48955,N_48344);
xnor UO_4929 (O_4929,N_49150,N_49898);
nor UO_4930 (O_4930,N_49637,N_49332);
nor UO_4931 (O_4931,N_48250,N_48536);
and UO_4932 (O_4932,N_49125,N_48032);
nor UO_4933 (O_4933,N_49903,N_49069);
and UO_4934 (O_4934,N_49322,N_49352);
xnor UO_4935 (O_4935,N_49568,N_49752);
xor UO_4936 (O_4936,N_49350,N_49022);
nor UO_4937 (O_4937,N_49262,N_49899);
xnor UO_4938 (O_4938,N_49841,N_49827);
nor UO_4939 (O_4939,N_49326,N_48679);
nand UO_4940 (O_4940,N_49305,N_48665);
nor UO_4941 (O_4941,N_48408,N_49358);
xor UO_4942 (O_4942,N_49118,N_48731);
or UO_4943 (O_4943,N_49658,N_48846);
and UO_4944 (O_4944,N_48052,N_48972);
and UO_4945 (O_4945,N_48149,N_48232);
or UO_4946 (O_4946,N_49298,N_48866);
or UO_4947 (O_4947,N_48163,N_49768);
xor UO_4948 (O_4948,N_48354,N_49267);
nand UO_4949 (O_4949,N_49644,N_48773);
and UO_4950 (O_4950,N_49131,N_49044);
xor UO_4951 (O_4951,N_48025,N_49721);
nor UO_4952 (O_4952,N_48738,N_48093);
nand UO_4953 (O_4953,N_49936,N_48871);
nor UO_4954 (O_4954,N_48736,N_48282);
or UO_4955 (O_4955,N_49803,N_49910);
or UO_4956 (O_4956,N_48330,N_49590);
or UO_4957 (O_4957,N_48343,N_49430);
nand UO_4958 (O_4958,N_49384,N_49859);
or UO_4959 (O_4959,N_49777,N_48452);
and UO_4960 (O_4960,N_49489,N_48459);
or UO_4961 (O_4961,N_49844,N_48081);
nand UO_4962 (O_4962,N_49697,N_48152);
nand UO_4963 (O_4963,N_49411,N_49381);
xor UO_4964 (O_4964,N_49967,N_49283);
or UO_4965 (O_4965,N_49258,N_49395);
or UO_4966 (O_4966,N_49630,N_48636);
xnor UO_4967 (O_4967,N_49418,N_49098);
nand UO_4968 (O_4968,N_49582,N_49811);
and UO_4969 (O_4969,N_49553,N_49363);
or UO_4970 (O_4970,N_49930,N_49676);
nand UO_4971 (O_4971,N_48192,N_49978);
and UO_4972 (O_4972,N_48949,N_48402);
nor UO_4973 (O_4973,N_49099,N_49318);
or UO_4974 (O_4974,N_48934,N_49659);
xnor UO_4975 (O_4975,N_49178,N_48736);
xnor UO_4976 (O_4976,N_49359,N_49657);
or UO_4977 (O_4977,N_49634,N_49381);
and UO_4978 (O_4978,N_49554,N_49166);
or UO_4979 (O_4979,N_49499,N_48455);
xnor UO_4980 (O_4980,N_48585,N_48471);
xor UO_4981 (O_4981,N_49350,N_49529);
nand UO_4982 (O_4982,N_48223,N_48492);
and UO_4983 (O_4983,N_49423,N_49964);
nand UO_4984 (O_4984,N_48626,N_48487);
or UO_4985 (O_4985,N_48521,N_49396);
nand UO_4986 (O_4986,N_49294,N_48131);
nor UO_4987 (O_4987,N_49720,N_48792);
or UO_4988 (O_4988,N_48673,N_48364);
nand UO_4989 (O_4989,N_49709,N_48778);
nand UO_4990 (O_4990,N_49445,N_49954);
nand UO_4991 (O_4991,N_48552,N_48139);
and UO_4992 (O_4992,N_48388,N_49974);
nor UO_4993 (O_4993,N_49408,N_49396);
nand UO_4994 (O_4994,N_49461,N_48614);
and UO_4995 (O_4995,N_48007,N_49805);
or UO_4996 (O_4996,N_48963,N_49527);
or UO_4997 (O_4997,N_49470,N_48911);
nand UO_4998 (O_4998,N_48802,N_48065);
nor UO_4999 (O_4999,N_49233,N_48051);
endmodule