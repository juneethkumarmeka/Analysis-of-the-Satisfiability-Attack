module basic_3000_30000_3500_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_2212,In_2925);
nor U1 (N_1,In_1096,In_38);
xnor U2 (N_2,In_2539,In_446);
xor U3 (N_3,In_2301,In_2841);
and U4 (N_4,In_1929,In_1425);
nor U5 (N_5,In_1370,In_2486);
xor U6 (N_6,In_925,In_1439);
and U7 (N_7,In_2970,In_963);
and U8 (N_8,In_669,In_1377);
or U9 (N_9,In_2251,In_442);
nor U10 (N_10,In_1864,In_843);
xor U11 (N_11,In_2609,In_198);
nor U12 (N_12,In_2821,In_291);
nor U13 (N_13,In_2046,In_1114);
or U14 (N_14,In_2109,In_1450);
nand U15 (N_15,In_801,In_2271);
nand U16 (N_16,In_2913,In_650);
or U17 (N_17,In_1239,In_1782);
xor U18 (N_18,In_601,In_2685);
and U19 (N_19,In_826,In_350);
nor U20 (N_20,In_1493,In_1479);
nand U21 (N_21,In_1170,In_2324);
or U22 (N_22,In_1834,In_1332);
nor U23 (N_23,In_2371,In_1651);
and U24 (N_24,In_978,In_1243);
or U25 (N_25,In_2388,In_961);
and U26 (N_26,In_1870,In_492);
nand U27 (N_27,In_1944,In_2876);
or U28 (N_28,In_932,In_441);
nand U29 (N_29,In_1320,In_1552);
nor U30 (N_30,In_1793,In_2911);
or U31 (N_31,In_2089,In_1165);
or U32 (N_32,In_2559,In_2941);
and U33 (N_33,In_677,In_1211);
or U34 (N_34,In_2160,In_2590);
nand U35 (N_35,In_829,In_1836);
nand U36 (N_36,In_981,In_1732);
or U37 (N_37,In_1542,In_634);
xor U38 (N_38,In_1945,In_1956);
xor U39 (N_39,In_233,In_400);
and U40 (N_40,In_2740,In_950);
nor U41 (N_41,In_2723,In_444);
or U42 (N_42,In_1185,In_1041);
nand U43 (N_43,In_311,In_782);
xor U44 (N_44,In_1666,In_1058);
xor U45 (N_45,In_2581,In_384);
xor U46 (N_46,In_1759,In_287);
or U47 (N_47,In_2368,In_2191);
or U48 (N_48,In_520,In_1531);
and U49 (N_49,In_566,In_183);
nor U50 (N_50,In_2446,In_652);
nor U51 (N_51,In_153,In_416);
or U52 (N_52,In_2727,In_2679);
nor U53 (N_53,In_1478,In_791);
or U54 (N_54,In_1973,In_1275);
xor U55 (N_55,In_748,In_1324);
xor U56 (N_56,In_1491,In_2257);
nand U57 (N_57,In_1704,In_2783);
and U58 (N_58,In_1691,In_2489);
nand U59 (N_59,In_1757,In_2756);
and U60 (N_60,In_1700,In_429);
xor U61 (N_61,In_1517,In_1045);
and U62 (N_62,In_832,In_513);
nand U63 (N_63,In_1784,In_1534);
nor U64 (N_64,In_2432,In_1141);
nand U65 (N_65,In_1481,In_1507);
and U66 (N_66,In_2347,In_1786);
nand U67 (N_67,In_2107,In_1317);
nor U68 (N_68,In_2282,In_600);
and U69 (N_69,In_468,In_2648);
xor U70 (N_70,In_2292,In_2782);
xor U71 (N_71,In_277,In_435);
and U72 (N_72,In_2550,In_1803);
nor U73 (N_73,In_2203,In_1471);
and U74 (N_74,In_649,In_2562);
and U75 (N_75,In_860,In_973);
xor U76 (N_76,In_2080,In_583);
or U77 (N_77,In_2015,In_1915);
or U78 (N_78,In_2653,In_1184);
xnor U79 (N_79,In_316,In_1730);
and U80 (N_80,In_1909,In_684);
nand U81 (N_81,In_466,In_642);
nor U82 (N_82,In_2177,In_521);
nor U83 (N_83,In_575,In_1011);
nor U84 (N_84,In_1035,In_63);
or U85 (N_85,In_2595,In_536);
nor U86 (N_86,In_2423,In_798);
xor U87 (N_87,In_2376,In_681);
or U88 (N_88,In_1105,In_2289);
nor U89 (N_89,In_2554,In_909);
or U90 (N_90,In_215,In_850);
and U91 (N_91,In_592,In_2773);
nor U92 (N_92,In_2403,In_1416);
nor U93 (N_93,In_990,In_1348);
or U94 (N_94,In_1843,In_2885);
or U95 (N_95,In_2457,In_1496);
nor U96 (N_96,In_1910,In_1971);
xnor U97 (N_97,In_1128,In_879);
nor U98 (N_98,In_122,In_313);
nor U99 (N_99,In_2240,In_2641);
or U100 (N_100,In_1998,In_2130);
nor U101 (N_101,In_2897,In_2220);
nor U102 (N_102,In_2448,In_643);
or U103 (N_103,In_565,In_2778);
and U104 (N_104,In_2419,In_703);
nand U105 (N_105,In_528,In_1350);
or U106 (N_106,In_896,In_2620);
xnor U107 (N_107,In_646,In_2495);
nand U108 (N_108,In_827,In_1925);
nor U109 (N_109,In_705,In_1596);
nor U110 (N_110,In_498,In_469);
or U111 (N_111,In_953,In_1231);
or U112 (N_112,In_814,In_2334);
nor U113 (N_113,In_2823,In_2933);
or U114 (N_114,In_2771,In_1619);
nor U115 (N_115,In_542,In_1225);
or U116 (N_116,In_785,In_2031);
and U117 (N_117,In_1993,In_2901);
nand U118 (N_118,In_1095,In_2165);
and U119 (N_119,In_2296,In_1374);
or U120 (N_120,In_151,In_1183);
nand U121 (N_121,In_201,In_1790);
nand U122 (N_122,In_2494,In_719);
or U123 (N_123,In_1187,In_998);
or U124 (N_124,In_1381,In_424);
and U125 (N_125,In_1369,In_647);
nand U126 (N_126,In_1553,In_1076);
nand U127 (N_127,In_1411,In_955);
xor U128 (N_128,In_1598,In_1193);
and U129 (N_129,In_2988,In_172);
or U130 (N_130,In_2365,In_91);
nor U131 (N_131,In_1281,In_1140);
or U132 (N_132,In_2711,In_1712);
nor U133 (N_133,In_1030,In_554);
or U134 (N_134,In_1622,In_2444);
nor U135 (N_135,In_1389,In_659);
nand U136 (N_136,In_1477,In_480);
and U137 (N_137,In_2518,In_1714);
and U138 (N_138,In_2415,In_1671);
nand U139 (N_139,In_2230,In_2318);
or U140 (N_140,In_377,In_2081);
nor U141 (N_141,In_2317,In_132);
and U142 (N_142,In_1357,In_837);
nand U143 (N_143,In_784,In_988);
xor U144 (N_144,In_1037,In_1807);
nor U145 (N_145,In_247,In_2927);
or U146 (N_146,In_1875,In_1069);
and U147 (N_147,In_1126,In_1075);
xnor U148 (N_148,In_49,In_2017);
nand U149 (N_149,In_2760,In_569);
nor U150 (N_150,In_1716,In_572);
and U151 (N_151,In_629,In_2661);
and U152 (N_152,In_2038,In_1489);
or U153 (N_153,In_506,In_2302);
or U154 (N_154,In_1982,In_2255);
or U155 (N_155,In_974,In_1868);
nand U156 (N_156,In_2267,In_694);
or U157 (N_157,In_2052,In_337);
nand U158 (N_158,In_617,In_2976);
and U159 (N_159,In_1558,In_1609);
nand U160 (N_160,In_2682,In_81);
nand U161 (N_161,In_486,In_2849);
nand U162 (N_162,In_2853,In_396);
nand U163 (N_163,In_2537,In_1541);
or U164 (N_164,In_181,In_1023);
nand U165 (N_165,In_1194,In_2630);
or U166 (N_166,In_2542,In_2796);
xor U167 (N_167,In_892,In_2894);
nor U168 (N_168,In_1575,In_574);
nand U169 (N_169,In_1897,In_1113);
nor U170 (N_170,In_2684,In_718);
nor U171 (N_171,In_1431,In_2065);
and U172 (N_172,In_2755,In_361);
and U173 (N_173,In_2026,In_0);
nor U174 (N_174,In_500,In_1046);
and U175 (N_175,In_1146,In_744);
and U176 (N_176,In_1607,In_640);
xor U177 (N_177,In_149,In_1571);
and U178 (N_178,In_353,In_787);
nor U179 (N_179,In_983,In_678);
nand U180 (N_180,In_2739,In_1545);
and U181 (N_181,In_2944,In_2263);
or U182 (N_182,In_2831,In_2131);
or U183 (N_183,In_2034,In_2409);
nand U184 (N_184,In_912,In_2435);
nor U185 (N_185,In_2604,In_937);
or U186 (N_186,In_872,In_1846);
or U187 (N_187,In_1959,In_530);
xor U188 (N_188,In_1401,In_1436);
xnor U189 (N_189,In_1572,In_1195);
nor U190 (N_190,In_1829,In_779);
nand U191 (N_191,In_940,In_2055);
and U192 (N_192,In_2442,In_2173);
or U193 (N_193,In_2624,In_227);
or U194 (N_194,In_2150,In_2380);
or U195 (N_195,In_481,In_224);
nand U196 (N_196,In_2651,In_944);
nor U197 (N_197,In_1343,In_1640);
nand U198 (N_198,In_387,In_495);
nor U199 (N_199,In_1620,In_1678);
or U200 (N_200,In_2361,In_2087);
or U201 (N_201,In_2708,In_366);
nor U202 (N_202,In_2765,In_1778);
xnor U203 (N_203,In_2033,In_380);
and U204 (N_204,In_1287,In_645);
nand U205 (N_205,In_44,In_76);
and U206 (N_206,In_50,In_715);
nand U207 (N_207,In_173,In_1798);
or U208 (N_208,In_2623,In_2504);
xor U209 (N_209,In_1990,In_1991);
nand U210 (N_210,In_1688,In_2654);
xnor U211 (N_211,In_2304,In_2837);
or U212 (N_212,In_2071,In_222);
nor U213 (N_213,In_1301,In_630);
nor U214 (N_214,In_2709,In_1877);
nor U215 (N_215,In_2194,In_1053);
nand U216 (N_216,In_2186,In_2519);
nand U217 (N_217,In_2333,In_450);
nor U218 (N_218,In_231,In_1881);
or U219 (N_219,In_2279,In_2450);
nand U220 (N_220,In_2642,In_516);
nor U221 (N_221,In_317,In_2346);
nor U222 (N_222,In_31,In_1858);
nand U223 (N_223,In_2445,In_840);
xor U224 (N_224,In_2068,In_2557);
nand U225 (N_225,In_1524,In_1890);
or U226 (N_226,In_1862,In_1682);
nand U227 (N_227,In_199,In_1335);
nor U228 (N_228,In_1373,In_2994);
nand U229 (N_229,In_917,In_1551);
and U230 (N_230,In_1634,In_831);
nand U231 (N_231,In_891,In_56);
and U232 (N_232,In_2511,In_662);
nand U233 (N_233,In_807,In_2284);
nor U234 (N_234,In_2319,In_2433);
and U235 (N_235,In_1774,In_914);
nand U236 (N_236,In_476,In_2366);
and U237 (N_237,In_1060,In_557);
nor U238 (N_238,In_1801,In_2949);
and U239 (N_239,In_460,In_1197);
and U240 (N_240,In_924,In_1333);
and U241 (N_241,In_939,In_293);
and U242 (N_242,In_2962,In_1444);
or U243 (N_243,In_2427,In_2585);
xor U244 (N_244,In_2076,In_186);
nand U245 (N_245,In_376,In_398);
or U246 (N_246,In_2352,In_26);
xnor U247 (N_247,In_1957,In_1254);
xor U248 (N_248,In_1339,In_1380);
xor U249 (N_249,In_138,In_663);
xnor U250 (N_250,In_2592,In_2938);
nor U251 (N_251,In_1931,In_1021);
nor U252 (N_252,In_676,In_1417);
and U253 (N_253,In_168,In_1302);
nor U254 (N_254,In_323,In_544);
and U255 (N_255,In_688,In_2514);
xnor U256 (N_256,In_329,In_2422);
xnor U257 (N_257,In_2695,In_1364);
or U258 (N_258,In_2386,In_561);
xnor U259 (N_259,In_1675,In_263);
xor U260 (N_260,In_1916,In_618);
nand U261 (N_261,In_2159,In_1894);
xor U262 (N_262,In_1448,In_1887);
nor U263 (N_263,In_810,In_698);
or U264 (N_264,In_237,In_2232);
and U265 (N_265,In_300,In_123);
and U266 (N_266,In_1074,In_274);
xnor U267 (N_267,In_88,In_711);
nand U268 (N_268,In_2873,In_1300);
nor U269 (N_269,In_2155,In_304);
or U270 (N_270,In_1528,In_1735);
xnor U271 (N_271,In_2209,In_704);
nor U272 (N_272,In_2090,In_1564);
and U273 (N_273,In_484,In_1777);
nand U274 (N_274,In_2407,In_1372);
or U275 (N_275,In_527,In_2474);
nand U276 (N_276,In_2016,In_2568);
nor U277 (N_277,In_1748,In_755);
nor U278 (N_278,In_2919,In_695);
or U279 (N_279,In_182,In_1307);
and U280 (N_280,In_1950,In_2461);
nand U281 (N_281,In_2729,In_2245);
nor U282 (N_282,In_994,In_33);
nand U283 (N_283,In_202,In_603);
nand U284 (N_284,In_2656,In_760);
nor U285 (N_285,In_675,In_142);
xor U286 (N_286,In_1669,In_1476);
nor U287 (N_287,In_60,In_1);
nor U288 (N_288,In_318,In_217);
or U289 (N_289,In_1192,In_2691);
nor U290 (N_290,In_1336,In_401);
xor U291 (N_291,In_1563,In_1226);
or U292 (N_292,In_1340,In_620);
and U293 (N_293,In_1158,In_434);
nor U294 (N_294,In_1198,In_1821);
nand U295 (N_295,In_2971,In_1454);
or U296 (N_296,In_2965,In_2753);
or U297 (N_297,In_1181,In_1326);
xor U298 (N_298,In_1539,In_1762);
nand U299 (N_299,In_644,In_1008);
or U300 (N_300,In_1772,In_2992);
nor U301 (N_301,In_2589,In_365);
or U302 (N_302,In_1808,In_1133);
nor U303 (N_303,In_864,In_325);
or U304 (N_304,In_221,In_1050);
xnor U305 (N_305,In_518,In_1854);
or U306 (N_306,In_587,In_1690);
and U307 (N_307,In_577,In_2847);
or U308 (N_308,In_911,In_2587);
nor U309 (N_309,In_1831,In_562);
or U310 (N_310,In_626,In_2775);
nand U311 (N_311,In_1764,In_2548);
xnor U312 (N_312,In_369,In_858);
nand U313 (N_313,In_427,In_1015);
nor U314 (N_314,In_1721,In_1227);
xnor U315 (N_315,In_2921,In_930);
nor U316 (N_316,In_2694,In_2698);
xnor U317 (N_317,In_1093,In_452);
nor U318 (N_318,In_1588,In_373);
nand U319 (N_319,In_975,In_242);
and U320 (N_320,In_598,In_1153);
or U321 (N_321,In_1718,In_1086);
or U322 (N_322,In_514,In_706);
and U323 (N_323,In_2225,In_220);
xor U324 (N_324,In_1160,In_721);
nand U325 (N_325,In_2106,In_195);
and U326 (N_326,In_2686,In_730);
and U327 (N_327,In_470,In_1665);
xnor U328 (N_328,In_893,In_2275);
and U329 (N_329,In_2268,In_156);
nand U330 (N_330,In_1070,In_942);
or U331 (N_331,In_1889,In_728);
xor U332 (N_332,In_1487,In_1648);
nand U333 (N_333,In_352,In_1310);
nor U334 (N_334,In_1771,In_1986);
nand U335 (N_335,In_41,In_1724);
nand U336 (N_336,In_2234,In_2597);
xnor U337 (N_337,In_2963,In_949);
xnor U338 (N_338,In_2036,In_2241);
nor U339 (N_339,In_2216,In_2822);
xnor U340 (N_340,In_1149,In_295);
nor U341 (N_341,In_2930,In_2824);
xnor U342 (N_342,In_2002,In_1804);
and U343 (N_343,In_2382,In_73);
or U344 (N_344,In_261,In_2561);
nand U345 (N_345,In_1662,In_1510);
and U346 (N_346,In_2731,In_2337);
or U347 (N_347,In_1446,In_64);
or U348 (N_348,In_815,In_1544);
or U349 (N_349,In_2136,In_2598);
nor U350 (N_350,In_797,In_2336);
and U351 (N_351,In_2198,In_581);
nor U352 (N_352,In_1178,In_2270);
and U353 (N_353,In_1328,In_2861);
nor U354 (N_354,In_239,In_1162);
and U355 (N_355,In_1610,In_2061);
nand U356 (N_356,In_821,In_2816);
and U357 (N_357,In_1382,In_1750);
nor U358 (N_358,In_2190,In_1294);
nor U359 (N_359,In_2870,In_2488);
nor U360 (N_360,In_1345,In_83);
nand U361 (N_361,In_2811,In_667);
nand U362 (N_362,In_1584,In_2468);
nor U363 (N_363,In_2817,In_596);
nor U364 (N_364,In_2794,In_1896);
and U365 (N_365,In_737,In_2758);
xor U366 (N_366,In_1430,In_5);
and U367 (N_367,In_1422,In_2785);
nand U368 (N_368,In_1859,In_2582);
and U369 (N_369,In_2132,In_2842);
xor U370 (N_370,In_943,In_1681);
xor U371 (N_371,In_1535,In_2535);
and U372 (N_372,In_1562,In_1802);
nor U373 (N_373,In_1822,In_631);
nor U374 (N_374,In_2395,In_1592);
xnor U375 (N_375,In_1776,In_2156);
xor U376 (N_376,In_1670,In_1710);
nand U377 (N_377,In_2262,In_2835);
or U378 (N_378,In_1039,In_59);
nand U379 (N_379,In_19,In_2780);
nand U380 (N_380,In_1219,In_2142);
or U381 (N_381,In_2907,In_1832);
nor U382 (N_382,In_1623,In_2238);
xnor U383 (N_383,In_2871,In_1511);
xor U384 (N_384,In_1933,In_1267);
xor U385 (N_385,In_2573,In_1943);
nor U386 (N_386,In_1787,In_2869);
or U387 (N_387,In_1080,In_364);
xor U388 (N_388,In_747,In_2223);
and U389 (N_389,In_1636,In_795);
nand U390 (N_390,In_1576,In_2144);
or U391 (N_391,In_1561,In_97);
nand U392 (N_392,In_1898,In_576);
nand U393 (N_393,In_2506,In_1375);
and U394 (N_394,In_30,In_870);
nand U395 (N_395,In_1988,In_457);
nand U396 (N_396,In_2168,In_1861);
and U397 (N_397,In_2717,In_1961);
nand U398 (N_398,In_1118,In_550);
nor U399 (N_399,In_2863,In_2985);
xnor U400 (N_400,In_2400,In_2607);
nor U401 (N_401,In_1215,In_894);
nor U402 (N_402,In_40,In_16);
and U403 (N_403,In_580,In_1135);
nand U404 (N_404,In_1498,In_420);
or U405 (N_405,In_612,In_62);
nand U406 (N_406,In_573,In_2786);
and U407 (N_407,In_547,In_1465);
nor U408 (N_408,In_1924,In_929);
and U409 (N_409,In_1617,In_2341);
and U410 (N_410,In_2097,In_2533);
xnor U411 (N_411,In_2233,In_2452);
xnor U412 (N_412,In_866,In_970);
and U413 (N_413,In_2390,In_2021);
nor U414 (N_414,In_1547,In_388);
xor U415 (N_415,In_472,In_2252);
xnor U416 (N_416,In_1627,In_18);
xnor U417 (N_417,In_413,In_1155);
xor U418 (N_418,In_2274,In_701);
nand U419 (N_419,In_133,In_855);
or U420 (N_420,In_2636,In_349);
or U421 (N_421,In_691,In_2261);
and U422 (N_422,In_2955,In_1108);
and U423 (N_423,In_2877,In_184);
xor U424 (N_424,In_406,In_226);
nor U425 (N_425,In_1191,In_1674);
nor U426 (N_426,In_2772,In_2044);
or U427 (N_427,In_2627,In_1720);
xor U428 (N_428,In_430,In_121);
nand U429 (N_429,In_2354,In_1205);
or U430 (N_430,In_757,In_991);
nand U431 (N_431,In_382,In_1233);
and U432 (N_432,In_979,In_2664);
xor U433 (N_433,In_1996,In_2544);
nor U434 (N_434,In_2683,In_2690);
xnor U435 (N_435,In_363,In_1272);
nand U436 (N_436,In_214,In_1999);
xnor U437 (N_437,In_273,In_1519);
and U438 (N_438,In_79,In_2974);
xor U439 (N_439,In_607,In_1441);
xnor U440 (N_440,In_2666,In_2312);
xor U441 (N_441,In_1156,In_2472);
or U442 (N_442,In_657,In_179);
and U443 (N_443,In_1811,In_1927);
xnor U444 (N_444,In_2171,In_2309);
xnor U445 (N_445,In_584,In_1819);
nand U446 (N_446,In_2175,In_2037);
and U447 (N_447,In_913,In_1055);
nand U448 (N_448,In_1523,In_2072);
or U449 (N_449,In_2655,In_543);
nand U450 (N_450,In_232,In_2688);
and U451 (N_451,In_69,In_1034);
nand U452 (N_452,In_188,In_799);
xnor U453 (N_453,In_2040,In_1376);
xor U454 (N_454,In_1794,In_283);
or U455 (N_455,In_2558,In_504);
xnor U456 (N_456,In_822,In_2411);
nand U457 (N_457,In_881,In_1270);
or U458 (N_458,In_271,In_1680);
nand U459 (N_459,In_1560,In_1161);
nand U460 (N_460,In_2538,In_833);
or U461 (N_461,In_882,In_1365);
nand U462 (N_462,In_507,In_1390);
or U463 (N_463,In_1483,In_889);
nand U464 (N_464,In_1084,In_432);
and U465 (N_465,In_1785,In_1687);
nor U466 (N_466,In_1362,In_651);
nand U467 (N_467,In_604,In_347);
and U468 (N_468,In_1739,In_1813);
xnor U469 (N_469,In_7,In_1447);
nor U470 (N_470,In_2769,In_1438);
or U471 (N_471,In_2250,In_2328);
nand U472 (N_472,In_2237,In_260);
nand U473 (N_473,In_236,In_2143);
and U474 (N_474,In_1077,In_2594);
xor U475 (N_475,In_116,In_2121);
or U476 (N_476,In_2622,In_2702);
and U477 (N_477,In_2918,In_137);
nor U478 (N_478,In_1157,In_599);
nand U479 (N_479,In_686,In_2798);
or U480 (N_480,In_1013,In_102);
nor U481 (N_481,In_1130,In_878);
and U482 (N_482,In_6,In_2266);
and U483 (N_483,In_1286,In_2219);
nand U484 (N_484,In_210,In_2952);
nand U485 (N_485,In_811,In_559);
and U486 (N_486,In_2524,In_964);
nor U487 (N_487,In_796,In_1460);
nand U488 (N_488,In_284,In_1906);
nor U489 (N_489,In_741,In_423);
and U490 (N_490,In_2942,In_2193);
and U491 (N_491,In_2172,In_608);
and U492 (N_492,In_2868,In_258);
nand U493 (N_493,In_1975,In_453);
or U494 (N_494,In_1468,In_1679);
xnor U495 (N_495,In_697,In_905);
nand U496 (N_496,In_370,In_1512);
nand U497 (N_497,In_926,In_2619);
xnor U498 (N_498,In_473,In_1625);
nor U499 (N_499,In_1432,In_722);
nand U500 (N_500,In_1017,In_1079);
xnor U501 (N_501,In_1304,In_749);
and U502 (N_502,In_250,In_65);
nor U503 (N_503,In_1694,In_1189);
xnor U504 (N_504,In_605,In_545);
xor U505 (N_505,In_1760,In_969);
or U506 (N_506,In_750,In_282);
and U507 (N_507,In_971,In_769);
nor U508 (N_508,In_1089,In_1914);
or U509 (N_509,In_192,In_2096);
nor U510 (N_510,In_2222,In_2946);
nand U511 (N_511,In_1057,In_1921);
nor U512 (N_512,In_2560,In_2665);
xnor U513 (N_513,In_2881,In_431);
xnor U514 (N_514,In_2520,In_2351);
or U515 (N_515,In_729,In_1061);
nand U516 (N_516,In_2088,In_1632);
xor U517 (N_517,In_1685,In_1062);
or U518 (N_518,In_1860,In_415);
and U519 (N_519,In_2936,In_789);
xor U520 (N_520,In_463,In_1400);
xnor U521 (N_521,In_803,In_1779);
nand U522 (N_522,In_2093,In_2313);
or U523 (N_523,In_511,In_292);
or U524 (N_524,In_2905,In_129);
and U525 (N_525,In_2205,In_2164);
nand U526 (N_526,In_857,In_24);
xor U527 (N_527,In_1800,In_1415);
nand U528 (N_528,In_134,In_2118);
or U529 (N_529,In_1565,In_1965);
and U530 (N_530,In_624,In_1752);
xnor U531 (N_531,In_1395,In_1518);
nand U532 (N_532,In_160,In_2588);
xnor U533 (N_533,In_2526,In_2948);
nand U534 (N_534,In_1245,In_1863);
xor U535 (N_535,In_374,In_209);
nor U536 (N_536,In_526,In_1989);
or U537 (N_537,In_2105,In_538);
and U538 (N_538,In_42,In_164);
and U539 (N_539,In_1516,In_394);
nor U540 (N_540,In_117,In_1009);
nor U541 (N_541,In_1812,In_2991);
and U542 (N_542,In_1878,In_2153);
or U543 (N_543,In_895,In_1246);
and U544 (N_544,In_421,In_635);
or U545 (N_545,In_1182,In_93);
xor U546 (N_546,In_2424,In_1816);
nand U547 (N_547,In_96,In_1919);
and U548 (N_548,In_1209,In_1744);
nor U549 (N_549,In_461,In_1977);
nand U550 (N_550,In_793,In_1653);
nand U551 (N_551,In_679,In_410);
xor U552 (N_552,In_1824,In_1384);
nor U553 (N_553,In_1148,In_2350);
xnor U554 (N_554,In_1538,In_853);
or U555 (N_555,In_1164,In_86);
and U556 (N_556,In_2699,In_2633);
and U557 (N_557,In_501,In_708);
nand U558 (N_558,In_1463,In_609);
nand U559 (N_559,In_834,In_1913);
xor U560 (N_560,In_12,In_321);
nand U561 (N_561,In_1667,In_2966);
nand U562 (N_562,In_2864,In_2467);
or U563 (N_563,In_55,In_713);
or U564 (N_564,In_1120,In_510);
nand U565 (N_565,In_1367,In_1885);
and U566 (N_566,In_2332,In_2384);
nor U567 (N_567,In_331,In_2889);
or U568 (N_568,In_252,In_606);
nand U569 (N_569,In_1329,In_262);
xnor U570 (N_570,In_1492,In_2712);
nand U571 (N_571,In_2206,In_2355);
or U572 (N_572,In_2123,In_67);
nand U573 (N_573,In_595,In_2492);
xnor U574 (N_574,In_82,In_2957);
nor U575 (N_575,In_1936,In_2269);
and U576 (N_576,In_1385,In_1536);
xor U577 (N_577,In_2327,In_848);
or U578 (N_578,In_245,In_2054);
nand U579 (N_579,In_960,In_2812);
nand U580 (N_580,In_1044,In_2827);
or U581 (N_581,In_2904,In_2744);
nand U582 (N_582,In_2362,In_1692);
and U583 (N_583,In_278,In_2977);
and U584 (N_584,In_1566,In_2405);
nor U585 (N_585,In_2483,In_1085);
nand U586 (N_586,In_1856,In_2387);
nor U587 (N_587,In_1488,In_191);
nand U588 (N_588,In_2989,In_2416);
or U589 (N_589,In_2441,In_1229);
nor U590 (N_590,In_471,In_2928);
nor U591 (N_591,In_267,In_2613);
and U592 (N_592,In_2874,In_1773);
or U593 (N_593,In_2050,In_2116);
or U594 (N_594,In_2998,In_792);
nand U595 (N_595,In_1673,In_1255);
xor U596 (N_596,In_946,In_493);
and U597 (N_597,In_1949,In_2133);
xnor U598 (N_598,In_27,In_166);
and U599 (N_599,In_1527,In_1847);
or U600 (N_600,In_2724,In_1263);
nor U601 (N_601,In_2845,In_1026);
or U602 (N_602,In_302,In_1048);
or U603 (N_603,In_594,In_1984);
xor U604 (N_604,In_2049,In_982);
or U605 (N_605,In_2343,In_2496);
nor U606 (N_606,In_1960,In_391);
nor U607 (N_607,In_654,In_658);
nor U608 (N_608,In_1292,In_2129);
xnor U609 (N_609,In_477,In_360);
nor U610 (N_610,In_1112,In_2809);
and U611 (N_611,In_1188,In_2465);
nand U612 (N_612,In_754,In_1749);
nand U613 (N_613,In_2791,In_2126);
xor U614 (N_614,In_2398,In_541);
nand U615 (N_615,In_1223,In_2378);
and U616 (N_616,In_1024,In_655);
nand U617 (N_617,In_2438,In_1761);
and U618 (N_618,In_2197,In_1284);
xor U619 (N_619,In_2990,In_1727);
and U620 (N_620,In_2242,In_505);
or U621 (N_621,In_1805,In_2789);
nand U622 (N_622,In_1795,In_2968);
xnor U623 (N_623,In_319,In_2001);
or U624 (N_624,In_1791,In_333);
xor U625 (N_625,In_1388,In_2202);
or U626 (N_626,In_2675,In_2000);
nor U627 (N_627,In_1792,In_1337);
or U628 (N_628,In_2618,In_208);
nor U629 (N_629,In_2576,In_809);
and U630 (N_630,In_1851,In_1419);
nand U631 (N_631,In_225,In_1063);
nand U632 (N_632,In_2074,In_2063);
and U633 (N_633,In_1305,In_934);
nor U634 (N_634,In_120,In_2578);
xnor U635 (N_635,In_2638,In_1279);
nand U636 (N_636,In_2418,In_2714);
and U637 (N_637,In_171,In_2855);
xnor U638 (N_638,In_1293,In_485);
xor U639 (N_639,In_2022,In_1296);
xor U640 (N_640,In_2315,In_1289);
and U641 (N_641,In_1297,In_2883);
xor U642 (N_642,In_1404,In_2570);
nand U643 (N_643,In_1259,In_614);
or U644 (N_644,In_412,In_2999);
or U645 (N_645,In_2208,In_841);
nand U646 (N_646,In_588,In_1139);
or U647 (N_647,In_2793,In_602);
and U648 (N_648,In_2053,In_2852);
xnor U649 (N_649,In_838,In_2295);
or U650 (N_650,In_692,In_1515);
xor U651 (N_651,In_2064,In_1942);
nand U652 (N_652,In_1591,In_1010);
and U653 (N_653,In_2961,In_2389);
or U654 (N_654,In_2029,In_636);
xor U655 (N_655,In_1767,In_354);
xnor U656 (N_656,In_2947,In_752);
nor U657 (N_657,In_2872,In_1230);
and U658 (N_658,In_918,In_1940);
xor U659 (N_659,In_2843,In_962);
xor U660 (N_660,In_1503,In_1758);
or U661 (N_661,In_2425,In_147);
nand U662 (N_662,In_1125,In_2606);
nor U663 (N_663,In_119,In_1845);
xor U664 (N_664,In_2857,In_494);
nor U665 (N_665,In_2272,In_2285);
and U666 (N_666,In_2476,In_2147);
and U667 (N_667,In_2982,In_957);
or U668 (N_668,In_1078,In_2480);
nor U669 (N_669,In_2331,In_1299);
nor U670 (N_670,In_700,In_131);
and U671 (N_671,In_357,In_1589);
nand U672 (N_672,In_1064,In_1360);
or U673 (N_673,In_2804,In_2807);
and U674 (N_674,In_997,In_758);
or U675 (N_675,In_519,In_1399);
nand U676 (N_676,In_2640,In_1445);
xnor U677 (N_677,In_475,In_1091);
or U678 (N_678,In_1893,In_1452);
and U679 (N_679,In_255,In_2715);
or U680 (N_680,In_847,In_800);
nor U681 (N_681,In_1261,In_61);
nand U682 (N_682,In_1796,In_448);
nor U683 (N_683,In_861,In_393);
nand U684 (N_684,In_13,In_296);
nor U685 (N_685,In_2657,In_2085);
or U686 (N_686,In_1809,In_1731);
and U687 (N_687,In_984,In_1235);
or U688 (N_688,In_639,In_371);
or U689 (N_689,In_1283,In_2579);
or U690 (N_690,In_1213,In_1322);
nor U691 (N_691,In_2737,In_2484);
or U692 (N_692,In_1769,In_2443);
nor U693 (N_693,In_1012,In_144);
xor U694 (N_694,In_656,In_1006);
nand U695 (N_695,In_1269,In_458);
or U696 (N_696,In_1599,In_2629);
and U697 (N_697,In_52,In_1788);
xor U698 (N_698,In_1618,In_2886);
or U699 (N_699,In_1175,In_2658);
xor U700 (N_700,In_1455,In_1964);
or U701 (N_701,In_976,In_2108);
or U702 (N_702,In_1865,In_196);
and U703 (N_703,In_696,In_1746);
or U704 (N_704,In_717,In_1608);
nand U705 (N_705,In_1497,In_956);
or U706 (N_706,In_1657,In_2751);
or U707 (N_707,In_109,In_2082);
or U708 (N_708,In_1733,In_2227);
xnor U709 (N_709,In_941,In_1948);
and U710 (N_710,In_1038,In_670);
nand U711 (N_711,In_1765,In_1241);
xor U712 (N_712,In_551,In_390);
nor U713 (N_713,In_178,In_2099);
and U714 (N_714,In_1974,In_2521);
xor U715 (N_715,In_2134,In_2353);
or U716 (N_716,In_1888,In_2950);
xnor U717 (N_717,In_411,In_727);
nand U718 (N_718,In_1216,In_2276);
or U719 (N_719,In_320,In_1051);
xnor U720 (N_720,In_1123,In_2226);
or U721 (N_721,In_673,In_842);
nor U722 (N_722,In_2004,In_1107);
xor U723 (N_723,In_2057,In_1351);
xnor U724 (N_724,In_2677,In_344);
nand U725 (N_725,In_1546,In_2569);
and U726 (N_726,In_615,In_2149);
and U727 (N_727,In_1319,In_2420);
nor U728 (N_728,In_1014,In_1457);
nand U729 (N_729,In_2231,In_2338);
xor U730 (N_730,In_338,In_1614);
nor U731 (N_731,In_2672,In_508);
nand U732 (N_732,In_1616,In_1111);
or U733 (N_733,In_2605,In_1451);
nand U734 (N_734,In_1533,In_1783);
and U735 (N_735,In_336,In_230);
or U736 (N_736,In_2704,In_1273);
xnor U737 (N_737,In_2908,In_666);
xor U738 (N_738,In_1100,In_883);
nand U739 (N_739,In_2635,In_2719);
xnor U740 (N_740,In_244,In_437);
nor U741 (N_741,In_2490,In_383);
nor U742 (N_742,In_1594,In_1696);
xnor U743 (N_743,In_2286,In_359);
and U744 (N_744,In_2545,In_1082);
and U745 (N_745,In_2014,In_2617);
nand U746 (N_746,In_653,In_303);
nor U747 (N_747,In_127,In_1876);
nor U748 (N_748,In_2323,In_2615);
and U749 (N_749,In_1347,In_2187);
or U750 (N_750,In_1409,In_2290);
or U751 (N_751,In_844,In_294);
nand U752 (N_752,In_770,In_2148);
xnor U753 (N_753,In_805,In_378);
and U754 (N_754,In_381,In_582);
and U755 (N_755,In_2459,In_2283);
or U756 (N_756,In_2436,In_2100);
nand U757 (N_757,In_180,In_958);
nor U758 (N_758,In_959,In_1649);
nand U759 (N_759,In_496,In_2880);
nor U760 (N_760,In_2763,In_43);
nand U761 (N_761,In_622,In_2030);
xnor U762 (N_762,In_1462,In_1972);
nor U763 (N_763,In_2645,In_1738);
and U764 (N_764,In_2707,In_2732);
and U765 (N_765,In_235,In_2377);
or U766 (N_766,In_2358,In_1701);
nor U767 (N_767,In_1568,In_916);
nor U768 (N_768,In_935,In_140);
nor U769 (N_769,In_2614,In_2278);
or U770 (N_770,In_205,In_1309);
nor U771 (N_771,In_254,In_890);
and U772 (N_772,In_671,In_2701);
and U773 (N_773,In_517,In_2784);
and U774 (N_774,In_2246,In_264);
xor U775 (N_775,In_2095,In_2273);
nand U776 (N_776,In_2580,In_2048);
nand U777 (N_777,In_788,In_1857);
xnor U778 (N_778,In_2632,In_491);
xnor U779 (N_779,In_552,In_330);
xnor U780 (N_780,In_780,In_308);
or U781 (N_781,In_269,In_902);
nand U782 (N_782,In_2596,In_1935);
and U783 (N_783,In_915,In_1799);
nor U784 (N_784,In_2764,In_57);
nand U785 (N_785,In_2047,In_1655);
nand U786 (N_786,In_560,In_2900);
and U787 (N_787,In_2487,In_2035);
nand U788 (N_788,In_2532,In_920);
xor U789 (N_789,In_2909,In_499);
nand U790 (N_790,In_854,In_356);
nor U791 (N_791,In_2541,In_2503);
or U792 (N_792,In_1131,In_2722);
nor U793 (N_793,In_1838,In_2349);
xor U794 (N_794,In_1490,In_972);
nand U795 (N_795,In_2608,In_2958);
nor U796 (N_796,In_1751,In_1664);
nand U797 (N_797,In_1201,In_425);
nand U798 (N_798,In_2196,In_2953);
xor U799 (N_799,In_1094,In_835);
or U800 (N_800,In_781,In_951);
and U801 (N_801,In_1007,In_1650);
nand U802 (N_802,In_1569,In_2996);
and U803 (N_803,In_2104,In_743);
nand U804 (N_804,In_1265,In_1699);
nand U805 (N_805,In_2253,In_2528);
and U806 (N_806,In_2135,In_2920);
xor U807 (N_807,In_641,In_1081);
and U808 (N_808,In_1473,In_53);
or U809 (N_809,In_2010,In_2599);
nor U810 (N_810,In_845,In_487);
and U811 (N_811,In_1427,In_92);
and U812 (N_812,In_1387,In_689);
nand U813 (N_813,In_29,In_702);
xor U814 (N_814,In_875,In_279);
xor U815 (N_815,In_90,In_58);
and U816 (N_816,In_2670,In_483);
and U817 (N_817,In_996,In_871);
nor U818 (N_818,In_2757,In_2215);
and U819 (N_819,In_2829,In_111);
xor U820 (N_820,In_819,In_2980);
xor U821 (N_821,In_426,In_2826);
or U822 (N_822,In_2127,In_2491);
xnor U823 (N_823,In_1207,In_2111);
and U824 (N_824,In_1018,In_289);
nand U825 (N_825,In_2455,In_1208);
nor U826 (N_826,In_1250,In_1453);
xnor U827 (N_827,In_1180,In_343);
nand U828 (N_828,In_17,In_1740);
nand U829 (N_829,In_852,In_778);
nand U830 (N_830,In_2512,In_768);
nor U831 (N_831,In_1358,In_68);
nand U832 (N_832,In_1966,In_1312);
nand U833 (N_833,In_1825,In_1978);
and U834 (N_834,In_625,In_107);
nand U835 (N_835,In_2181,In_95);
and U836 (N_836,In_2611,In_1049);
nand U837 (N_837,In_489,In_1036);
and U838 (N_838,In_2750,In_1855);
and U839 (N_839,In_2774,In_1780);
or U840 (N_840,In_2882,In_2553);
nor U841 (N_841,In_2045,In_128);
and U842 (N_842,In_2531,In_1520);
xnor U843 (N_843,In_328,In_2348);
or U844 (N_844,In_23,In_897);
nor U845 (N_845,In_334,In_1658);
nand U846 (N_846,In_2929,In_418);
nor U847 (N_847,In_2426,In_2373);
or U848 (N_848,In_1525,In_206);
nor U849 (N_849,In_2102,In_2204);
or U850 (N_850,In_585,In_1695);
xnor U851 (N_851,In_405,In_1019);
or U852 (N_852,In_189,In_351);
and U853 (N_853,In_2244,In_1349);
or U854 (N_854,In_464,In_2369);
xnor U855 (N_855,In_1656,In_1257);
nand U856 (N_856,In_1001,In_933);
nor U857 (N_857,In_2516,In_2981);
xor U858 (N_858,In_802,In_2603);
xor U859 (N_859,In_1321,In_2066);
or U860 (N_860,In_98,In_75);
nand U861 (N_861,In_2954,In_2140);
nand U862 (N_862,In_1706,In_1025);
xor U863 (N_863,In_813,In_690);
nand U864 (N_864,In_2043,In_2571);
nand U865 (N_865,In_229,In_1248);
or U866 (N_866,In_2248,In_1886);
nor U867 (N_867,In_1844,In_2379);
nor U868 (N_868,In_1177,In_1042);
xor U869 (N_869,In_555,In_512);
xnor U870 (N_870,In_2830,In_1702);
nand U871 (N_871,In_2865,In_1456);
and U872 (N_872,In_2466,In_2254);
and U873 (N_873,In_1725,In_1615);
and U874 (N_874,In_2828,In_571);
xor U875 (N_875,In_1059,In_1236);
nand U876 (N_876,In_2124,In_2820);
nor U877 (N_877,In_2051,In_502);
or U878 (N_878,In_1461,In_2460);
nor U879 (N_879,In_2482,In_2264);
nand U880 (N_880,In_456,In_1124);
nor U881 (N_881,In_1147,In_2703);
nand U882 (N_882,In_1022,In_1522);
or U883 (N_883,In_141,In_80);
or U884 (N_884,In_2819,In_1661);
xor U885 (N_885,In_2462,In_1573);
and U886 (N_886,In_2179,In_549);
and U887 (N_887,In_399,In_1981);
nand U888 (N_888,In_1282,In_2025);
xor U889 (N_889,In_2978,In_286);
nor U890 (N_890,In_738,In_2434);
and U891 (N_891,In_868,In_445);
or U892 (N_892,In_2878,In_1150);
xor U893 (N_893,In_818,In_1753);
or U894 (N_894,In_1693,In_1741);
nand U895 (N_895,In_2891,In_2114);
and U896 (N_896,In_1869,In_115);
xnor U897 (N_897,In_2860,In_2833);
or U898 (N_898,In_2265,In_169);
or U899 (N_899,In_2940,In_265);
xor U900 (N_900,In_1506,In_355);
or U901 (N_901,In_1970,In_154);
nand U902 (N_902,In_368,In_1923);
xor U903 (N_903,In_808,In_1396);
nand U904 (N_904,In_2217,In_2814);
xnor U905 (N_905,In_1203,In_2899);
nor U906 (N_906,In_1828,In_823);
or U907 (N_907,In_1559,In_693);
and U908 (N_908,In_877,In_2027);
nand U909 (N_909,In_1848,In_777);
nand U910 (N_910,In_1826,In_2840);
and U911 (N_911,In_1880,In_2236);
or U912 (N_912,In_1494,In_2602);
nand U913 (N_913,In_1806,In_2360);
or U914 (N_914,In_1303,In_2803);
or U915 (N_915,In_2776,In_2359);
nor U916 (N_916,In_433,In_2993);
nor U917 (N_917,In_1132,In_2738);
nor U918 (N_918,In_938,In_2330);
or U919 (N_919,In_2335,In_348);
and U920 (N_920,In_2326,In_1850);
or U921 (N_921,In_1938,In_2188);
xnor U922 (N_922,In_2094,In_1402);
nor U923 (N_923,In_1295,In_1839);
nand U924 (N_924,In_2471,In_1548);
nor U925 (N_925,In_2801,In_2414);
nor U926 (N_926,In_1905,In_103);
xnor U927 (N_927,In_2009,In_509);
nand U928 (N_928,In_207,In_567);
xor U929 (N_929,In_999,In_1501);
and U930 (N_930,In_2761,In_765);
nor U931 (N_931,In_1144,In_2696);
and U932 (N_932,In_440,In_2910);
nand U933 (N_933,In_1603,In_1557);
or U934 (N_934,In_1403,In_2056);
xnor U935 (N_935,In_1842,In_2200);
or U936 (N_936,In_1711,In_266);
or U937 (N_937,In_709,In_307);
xor U938 (N_938,In_28,In_2166);
and U939 (N_939,In_419,In_1280);
nand U940 (N_940,In_1707,In_1371);
nor U941 (N_941,In_1734,In_1683);
nor U942 (N_942,In_212,In_1217);
nor U943 (N_943,In_948,In_2591);
nor U944 (N_944,In_1142,In_2916);
and U945 (N_945,In_2572,In_1097);
or U946 (N_946,In_859,In_2329);
nor U947 (N_947,In_1033,In_1621);
or U948 (N_948,In_2507,In_240);
xnor U949 (N_949,In_1138,In_849);
and U950 (N_950,In_219,In_794);
xor U951 (N_951,In_1449,In_1630);
or U952 (N_952,In_2287,In_2391);
and U953 (N_953,In_1629,In_1052);
xnor U954 (N_954,In_2668,In_2059);
nor U955 (N_955,In_967,In_2728);
or U956 (N_956,In_2084,In_922);
or U957 (N_957,In_324,In_680);
nand U958 (N_958,In_1072,In_1443);
nand U959 (N_959,In_2800,In_1171);
and U960 (N_960,In_281,In_1628);
nor U961 (N_961,In_1073,In_2898);
or U962 (N_962,In_2943,In_1334);
nand U963 (N_963,In_759,In_1412);
and U964 (N_964,In_2481,In_2451);
nor U965 (N_965,In_306,In_2399);
or U966 (N_966,In_2357,In_2600);
and U967 (N_967,In_1994,In_94);
nor U968 (N_968,In_816,In_1756);
nand U969 (N_969,In_1871,In_1726);
nand U970 (N_970,In_2429,In_22);
nor U971 (N_971,In_2787,In_2374);
and U972 (N_972,In_1660,In_1763);
and U973 (N_973,In_1434,In_2007);
and U974 (N_974,In_2967,In_2734);
and U975 (N_975,In_2844,In_2410);
nor U976 (N_976,In_358,In_746);
xor U977 (N_977,In_2667,In_2939);
xnor U978 (N_978,In_2396,In_2401);
nand U979 (N_979,In_1997,In_1379);
xor U980 (N_980,In_1323,In_1247);
xor U981 (N_981,In_2705,In_1366);
nor U982 (N_982,In_248,In_2687);
or U983 (N_983,In_761,In_297);
and U984 (N_984,In_312,In_627);
xor U985 (N_985,In_2229,In_2612);
and U986 (N_986,In_2372,In_2862);
and U987 (N_987,In_2639,In_32);
nor U988 (N_988,In_2839,In_764);
and U989 (N_989,In_404,In_1641);
and U990 (N_990,In_2383,In_1736);
nand U991 (N_991,In_125,In_1327);
xnor U992 (N_992,In_885,In_2086);
and U993 (N_993,In_1987,In_1912);
xnor U994 (N_994,In_1068,In_417);
and U995 (N_995,In_776,In_1676);
or U996 (N_996,In_2437,In_234);
or U997 (N_997,In_2945,In_683);
nand U998 (N_998,In_1952,In_2028);
and U999 (N_999,In_2119,In_2397);
xnor U1000 (N_1000,In_1098,In_1315);
and U1001 (N_1001,In_986,In_1413);
or U1002 (N_1002,In_1238,In_533);
nand U1003 (N_1003,In_568,In_1908);
and U1004 (N_1004,In_157,In_1837);
xor U1005 (N_1005,In_786,In_1087);
nor U1006 (N_1006,In_37,In_2174);
or U1007 (N_1007,In_1717,In_1145);
and U1008 (N_1008,In_1420,In_2797);
nor U1009 (N_1009,In_459,In_766);
xor U1010 (N_1010,In_1918,In_1677);
and U1011 (N_1011,In_1612,In_1004);
nand U1012 (N_1012,In_395,In_2912);
nor U1013 (N_1013,In_1249,In_1930);
nor U1014 (N_1014,In_1278,In_2243);
nor U1015 (N_1015,In_342,In_2593);
and U1016 (N_1016,In_2019,In_309);
nor U1017 (N_1017,In_1827,In_249);
or U1018 (N_1018,In_908,In_280);
nand U1019 (N_1019,In_87,In_176);
nand U1020 (N_1020,In_2062,In_1256);
and U1021 (N_1021,In_327,In_385);
and U1022 (N_1022,In_2616,In_1143);
nand U1023 (N_1023,In_2154,In_1586);
or U1024 (N_1024,In_1242,In_1104);
nor U1025 (N_1025,In_2563,In_2128);
nand U1026 (N_1026,In_2367,In_1065);
xor U1027 (N_1027,In_1567,In_165);
nor U1028 (N_1028,In_2726,In_326);
nor U1029 (N_1029,In_1313,In_672);
nand U1030 (N_1030,In_1031,In_100);
or U1031 (N_1031,In_736,In_2502);
nor U1032 (N_1032,In_2935,In_1597);
or U1033 (N_1033,In_2479,In_632);
nand U1034 (N_1034,In_1266,In_1101);
or U1035 (N_1035,In_2306,In_2693);
and U1036 (N_1036,In_1840,In_2370);
xor U1037 (N_1037,In_1768,In_1407);
nand U1038 (N_1038,In_735,In_1437);
nand U1039 (N_1039,In_2628,In_1635);
nor U1040 (N_1040,In_1581,In_2091);
and U1041 (N_1041,In_2473,In_1815);
and U1042 (N_1042,In_2180,In_888);
nand U1043 (N_1043,In_2777,In_1686);
or U1044 (N_1044,In_2184,In_2649);
xor U1045 (N_1045,In_1713,In_112);
or U1046 (N_1046,In_989,In_1979);
or U1047 (N_1047,In_2601,In_2960);
or U1048 (N_1048,In_272,In_2903);
nand U1049 (N_1049,In_2888,In_2463);
and U1050 (N_1050,In_2277,In_873);
nor U1051 (N_1051,In_197,In_397);
nand U1052 (N_1052,In_2176,In_2730);
and U1053 (N_1053,In_1823,In_2926);
xnor U1054 (N_1054,In_931,In_1781);
nand U1055 (N_1055,In_1529,In_824);
nor U1056 (N_1056,In_927,In_1102);
nor U1057 (N_1057,In_1937,In_532);
xor U1058 (N_1058,In_613,In_288);
nand U1059 (N_1059,In_2674,In_2626);
or U1060 (N_1060,In_1288,In_2513);
or U1061 (N_1061,In_1423,In_2320);
and U1062 (N_1062,In_1106,In_621);
xnor U1063 (N_1063,In_1421,In_563);
or U1064 (N_1064,In_2192,In_1129);
xnor U1065 (N_1065,In_732,In_1134);
nor U1066 (N_1066,In_9,In_2469);
nand U1067 (N_1067,In_2316,In_2973);
or U1068 (N_1068,In_1891,In_716);
and U1069 (N_1069,In_2152,In_161);
or U1070 (N_1070,In_1550,In_1330);
and U1071 (N_1071,In_919,In_707);
or U1072 (N_1072,In_2075,In_1742);
nor U1073 (N_1073,In_170,In_2145);
or U1074 (N_1074,In_1167,In_315);
and U1075 (N_1075,In_2112,In_1251);
or U1076 (N_1076,In_136,In_162);
nor U1077 (N_1077,In_2497,In_619);
nor U1078 (N_1078,In_699,In_2733);
and U1079 (N_1079,In_305,In_1470);
nor U1080 (N_1080,In_290,In_99);
nand U1081 (N_1081,In_1122,In_2498);
or U1082 (N_1082,In_720,In_223);
or U1083 (N_1083,In_465,In_1818);
or U1084 (N_1084,In_1901,In_2385);
xnor U1085 (N_1085,In_2749,In_2625);
xor U1086 (N_1086,In_2005,In_839);
nand U1087 (N_1087,In_1088,In_1775);
xnor U1088 (N_1088,In_1932,In_851);
and U1089 (N_1089,In_2915,In_1426);
and U1090 (N_1090,In_2530,In_1316);
and U1091 (N_1091,In_2832,In_2984);
nand U1092 (N_1092,In_2207,In_1268);
nor U1093 (N_1093,In_455,In_106);
or U1094 (N_1094,In_1495,In_1587);
or U1095 (N_1095,In_593,In_1442);
xnor U1096 (N_1096,In_1090,In_2914);
xor U1097 (N_1097,In_2069,In_1951);
xor U1098 (N_1098,In_2151,In_804);
and U1099 (N_1099,In_1976,In_159);
xor U1100 (N_1100,In_146,In_1353);
or U1101 (N_1101,In_1405,In_2508);
nand U1102 (N_1102,In_812,In_310);
and U1103 (N_1103,In_2766,In_1613);
or U1104 (N_1104,In_1127,In_771);
xor U1105 (N_1105,In_2141,In_2846);
or U1106 (N_1106,In_1639,In_2110);
nor U1107 (N_1107,In_2713,In_2808);
xor U1108 (N_1108,In_2975,In_1593);
xnor U1109 (N_1109,In_2813,In_1647);
or U1110 (N_1110,In_2161,In_1895);
nand U1111 (N_1111,In_1016,In_21);
xnor U1112 (N_1112,In_586,In_2013);
xnor U1113 (N_1113,In_2681,In_2663);
nor U1114 (N_1114,In_2260,In_534);
and U1115 (N_1115,In_820,In_921);
nor U1116 (N_1116,In_1502,In_2644);
nor U1117 (N_1117,In_1355,In_2098);
and U1118 (N_1118,In_2167,In_977);
or U1119 (N_1119,In_1900,In_2637);
and U1120 (N_1120,In_2195,In_1504);
nor U1121 (N_1121,In_488,In_2157);
and U1122 (N_1122,In_1318,In_564);
and U1123 (N_1123,In_1841,In_1505);
xnor U1124 (N_1124,In_723,In_1770);
and U1125 (N_1125,In_2893,In_2169);
and U1126 (N_1126,In_923,In_2182);
xnor U1127 (N_1127,In_2762,In_2342);
nor U1128 (N_1128,In_1220,In_2662);
xnor U1129 (N_1129,In_314,In_2745);
or U1130 (N_1130,In_135,In_579);
nand U1131 (N_1131,In_2856,In_525);
and U1132 (N_1132,In_1083,In_72);
and U1133 (N_1133,In_1645,In_1595);
nand U1134 (N_1134,In_2475,In_2079);
nand U1135 (N_1135,In_1480,In_1532);
nand U1136 (N_1136,In_402,In_1537);
nand U1137 (N_1137,In_1264,In_428);
and U1138 (N_1138,In_158,In_285);
nand U1139 (N_1139,In_740,In_2643);
nand U1140 (N_1140,In_1747,In_623);
nand U1141 (N_1141,In_529,In_1224);
nor U1142 (N_1142,In_762,In_1985);
xor U1143 (N_1143,In_34,In_301);
nand U1144 (N_1144,In_70,In_1969);
and U1145 (N_1145,In_1392,In_2951);
xor U1146 (N_1146,In_980,In_1884);
nor U1147 (N_1147,In_1152,In_856);
or U1148 (N_1148,In_2499,In_1137);
nor U1149 (N_1149,In_1954,In_2478);
and U1150 (N_1150,In_2892,In_2454);
xnor U1151 (N_1151,In_1797,In_1398);
nand U1152 (N_1152,In_490,In_2555);
nor U1153 (N_1153,In_1383,In_503);
xnor U1154 (N_1154,In_2439,In_1356);
nand U1155 (N_1155,In_228,In_556);
nor U1156 (N_1156,In_1833,In_539);
nand U1157 (N_1157,In_1291,In_482);
nand U1158 (N_1158,In_1429,In_1154);
nand U1159 (N_1159,In_616,In_1737);
nand U1160 (N_1160,In_863,In_443);
xnor U1161 (N_1161,In_1314,In_590);
or U1162 (N_1162,In_447,In_2);
nor U1163 (N_1163,In_1212,In_1585);
nand U1164 (N_1164,In_276,In_322);
nor U1165 (N_1165,In_1928,In_449);
and U1166 (N_1166,In_1240,In_389);
nand U1167 (N_1167,In_884,In_886);
and U1168 (N_1168,In_1967,In_1883);
or U1169 (N_1169,In_2525,In_2392);
nor U1170 (N_1170,In_118,In_1947);
nor U1171 (N_1171,In_589,In_54);
or U1172 (N_1172,In_1459,In_243);
nor U1173 (N_1173,In_1472,In_2344);
nor U1174 (N_1174,In_2546,In_20);
xnor U1175 (N_1175,In_2408,In_887);
nand U1176 (N_1176,In_2549,In_4);
or U1177 (N_1177,In_1672,In_2583);
and U1178 (N_1178,In_2294,In_1346);
nor U1179 (N_1179,In_2522,In_1485);
nand U1180 (N_1180,In_2447,In_1331);
nor U1181 (N_1181,In_436,In_2556);
xnor U1182 (N_1182,In_2854,In_2895);
xnor U1183 (N_1183,In_1222,In_2956);
or U1184 (N_1184,In_867,In_1066);
and U1185 (N_1185,In_2077,In_174);
xor U1186 (N_1186,In_2884,In_1556);
nand U1187 (N_1187,In_85,In_2647);
nor U1188 (N_1188,In_1397,In_438);
xnor U1189 (N_1189,In_1391,In_403);
nand U1190 (N_1190,In_2851,In_2340);
xor U1191 (N_1191,In_2564,In_253);
or U1192 (N_1192,In_2321,In_48);
xnor U1193 (N_1193,In_78,In_257);
nand U1194 (N_1194,In_497,In_2485);
xnor U1195 (N_1195,In_1577,In_1308);
and U1196 (N_1196,In_77,In_1980);
and U1197 (N_1197,In_194,In_836);
or U1198 (N_1198,In_724,In_1054);
or U1199 (N_1199,In_340,In_84);
nand U1200 (N_1200,In_2818,In_335);
nand U1201 (N_1201,In_1032,In_1467);
nor U1202 (N_1202,In_1466,In_2239);
or U1203 (N_1203,In_638,In_2345);
nand U1204 (N_1204,In_2402,In_2917);
and U1205 (N_1205,In_2565,In_2375);
nand U1206 (N_1206,In_1196,In_660);
or U1207 (N_1207,In_904,In_1766);
xor U1208 (N_1208,In_3,In_1814);
or U1209 (N_1209,In_2011,In_2906);
nand U1210 (N_1210,In_1199,In_2440);
and U1211 (N_1211,In_1210,In_1879);
and U1212 (N_1212,In_1631,In_467);
and U1213 (N_1213,In_1830,In_114);
or U1214 (N_1214,In_2754,In_2720);
and U1215 (N_1215,In_2523,In_108);
xor U1216 (N_1216,In_2867,In_2183);
nand U1217 (N_1217,In_2834,In_954);
and U1218 (N_1218,In_1474,In_1424);
or U1219 (N_1219,In_1611,In_2987);
nand U1220 (N_1220,In_1703,In_2650);
nand U1221 (N_1221,In_1464,In_830);
xor U1222 (N_1222,In_846,In_2281);
nor U1223 (N_1223,In_407,In_1698);
and U1224 (N_1224,In_2959,In_1172);
and U1225 (N_1225,In_341,In_45);
or U1226 (N_1226,In_2838,In_2023);
and U1227 (N_1227,In_775,In_1244);
nor U1228 (N_1228,In_2536,In_1116);
nand U1229 (N_1229,In_869,In_2567);
and U1230 (N_1230,In_1902,In_1554);
nand U1231 (N_1231,In_1325,In_1168);
nor U1232 (N_1232,In_1602,In_2117);
or U1233 (N_1233,In_910,In_1817);
nor U1234 (N_1234,In_1754,In_2552);
or U1235 (N_1235,In_1440,In_1500);
or U1236 (N_1236,In_1027,In_1968);
and U1237 (N_1237,In_2449,In_2505);
or U1238 (N_1238,In_2802,In_1258);
xor U1239 (N_1239,In_710,In_2634);
nand U1240 (N_1240,In_1159,In_2020);
and U1241 (N_1241,In_216,In_1722);
or U1242 (N_1242,In_874,In_89);
and U1243 (N_1243,In_2716,In_346);
nand U1244 (N_1244,In_1574,In_1200);
nor U1245 (N_1245,In_664,In_1354);
nor U1246 (N_1246,In_2070,In_1508);
or U1247 (N_1247,In_2510,In_1911);
xnor U1248 (N_1248,In_2185,In_145);
nor U1249 (N_1249,In_386,In_451);
and U1250 (N_1250,In_2527,In_2747);
or U1251 (N_1251,In_1056,In_2464);
and U1252 (N_1252,In_2058,In_2887);
nor U1253 (N_1253,In_2660,In_454);
nand U1254 (N_1254,In_2697,In_372);
nand U1255 (N_1255,In_1958,In_1290);
or U1256 (N_1256,In_2018,In_1386);
xnor U1257 (N_1257,In_2456,In_712);
nor U1258 (N_1258,In_1202,In_1029);
nand U1259 (N_1259,In_2676,In_2235);
xnor U1260 (N_1260,In_2413,In_1922);
nor U1261 (N_1261,In_2858,In_2743);
nor U1262 (N_1262,In_422,In_2735);
xor U1263 (N_1263,In_2280,In_2859);
and U1264 (N_1264,In_1067,In_1276);
or U1265 (N_1265,In_1363,In_1852);
and U1266 (N_1266,In_2659,In_2363);
nor U1267 (N_1267,In_2574,In_1237);
or U1268 (N_1268,In_190,In_339);
nand U1269 (N_1269,In_825,In_2247);
nand U1270 (N_1270,In_1428,In_1934);
nand U1271 (N_1271,In_806,In_1190);
nor U1272 (N_1272,In_39,In_46);
nor U1273 (N_1273,In_2394,In_177);
xnor U1274 (N_1274,In_104,In_1136);
nand U1275 (N_1275,In_2879,In_2748);
xnor U1276 (N_1276,In_1186,In_1174);
and U1277 (N_1277,In_1917,In_880);
and U1278 (N_1278,In_71,In_828);
nand U1279 (N_1279,In_367,In_1393);
and U1280 (N_1280,In_2024,In_790);
xor U1281 (N_1281,In_2083,In_2850);
xor U1282 (N_1282,In_578,In_2534);
xnor U1283 (N_1283,In_362,In_2997);
xor U1284 (N_1284,In_238,In_139);
and U1285 (N_1285,In_2115,In_2790);
or U1286 (N_1286,In_2692,In_2258);
nor U1287 (N_1287,In_992,In_259);
nand U1288 (N_1288,In_2032,In_2073);
and U1289 (N_1289,In_2039,In_1513);
xnor U1290 (N_1290,In_2700,In_2146);
and U1291 (N_1291,In_1115,In_150);
xnor U1292 (N_1292,In_2741,In_685);
or U1293 (N_1293,In_1646,In_1435);
nand U1294 (N_1294,In_1020,In_2300);
xnor U1295 (N_1295,In_2932,In_2902);
nor U1296 (N_1296,In_1475,In_110);
nand U1297 (N_1297,In_1482,In_163);
nor U1298 (N_1298,In_1003,In_591);
and U1299 (N_1299,In_903,In_478);
nor U1300 (N_1300,In_2678,In_2163);
and U1301 (N_1301,In_531,In_2768);
nor U1302 (N_1302,In_1578,In_1708);
nand U1303 (N_1303,In_11,In_611);
nand U1304 (N_1304,In_2431,In_1920);
or U1305 (N_1305,In_774,In_1179);
or U1306 (N_1306,In_2139,In_409);
nand U1307 (N_1307,In_515,In_2673);
or U1308 (N_1308,In_2836,In_345);
nor U1309 (N_1309,In_241,In_2509);
nor U1310 (N_1310,In_152,In_2671);
nor U1311 (N_1311,In_1361,In_35);
nand U1312 (N_1312,In_1642,In_751);
nor U1313 (N_1313,In_1151,In_2428);
nand U1314 (N_1314,In_1874,In_682);
xnor U1315 (N_1315,In_1406,In_2113);
nand U1316 (N_1316,In_2792,In_2256);
nand U1317 (N_1317,In_2199,In_2979);
and U1318 (N_1318,In_2964,In_218);
and U1319 (N_1319,In_1099,In_1955);
or U1320 (N_1320,In_1176,In_597);
or U1321 (N_1321,In_865,In_2746);
nand U1322 (N_1322,In_1028,In_2825);
or U1323 (N_1323,In_1643,In_2221);
xnor U1324 (N_1324,In_966,In_628);
nand U1325 (N_1325,In_213,In_74);
nand U1326 (N_1326,In_2299,In_2325);
or U1327 (N_1327,In_2983,In_379);
and U1328 (N_1328,In_25,In_1526);
xnor U1329 (N_1329,In_901,In_1092);
or U1330 (N_1330,In_2458,In_1663);
or U1331 (N_1331,In_1983,In_2249);
nor U1332 (N_1332,In_1169,In_2652);
nor U1333 (N_1333,In_270,In_1234);
nand U1334 (N_1334,In_633,In_2779);
nor U1335 (N_1335,In_1604,In_1232);
and U1336 (N_1336,In_1206,In_2575);
or U1337 (N_1337,In_1953,In_2810);
nand U1338 (N_1338,In_1946,In_1218);
nor U1339 (N_1339,In_2259,In_1810);
nor U1340 (N_1340,In_648,In_2969);
xor U1341 (N_1341,In_1723,In_540);
xor U1342 (N_1342,In_2078,In_1486);
nand U1343 (N_1343,In_1540,In_1040);
nand U1344 (N_1344,In_2610,In_1606);
xnor U1345 (N_1345,In_15,In_105);
nand U1346 (N_1346,In_1872,In_66);
or U1347 (N_1347,In_2924,In_2138);
nor U1348 (N_1348,In_1904,In_1684);
xnor U1349 (N_1349,In_773,In_408);
nand U1350 (N_1350,In_251,In_1907);
and U1351 (N_1351,In_1652,In_2515);
nor U1352 (N_1352,In_1820,In_1110);
xnor U1353 (N_1353,In_2934,In_2759);
nand U1354 (N_1354,In_1298,In_1583);
xor U1355 (N_1355,In_1047,In_2178);
xnor U1356 (N_1356,In_203,In_1414);
or U1357 (N_1357,In_1359,In_2453);
or U1358 (N_1358,In_1121,In_907);
xnor U1359 (N_1359,In_2815,In_2214);
nor U1360 (N_1360,In_1311,In_2158);
nand U1361 (N_1361,In_2228,In_185);
xnor U1362 (N_1362,In_2101,In_155);
nand U1363 (N_1363,In_2213,In_763);
and U1364 (N_1364,In_1600,In_2421);
nand U1365 (N_1365,In_899,In_1644);
nand U1366 (N_1366,In_1637,In_1605);
nor U1367 (N_1367,In_535,In_2517);
and U1368 (N_1368,In_714,In_1715);
xor U1369 (N_1369,In_2972,In_2931);
nor U1370 (N_1370,In_876,In_126);
and U1371 (N_1371,In_375,In_200);
nor U1372 (N_1372,In_523,In_439);
xnor U1373 (N_1373,In_2003,In_1043);
and U1374 (N_1374,In_2577,In_1719);
nand U1375 (N_1375,In_1109,In_2393);
or U1376 (N_1376,In_1433,In_817);
xor U1377 (N_1377,In_2631,In_947);
or U1378 (N_1378,In_1002,In_1274);
or U1379 (N_1379,In_965,In_985);
and U1380 (N_1380,In_2339,In_1071);
xor U1381 (N_1381,In_1338,In_1899);
nand U1382 (N_1382,In_731,In_2162);
nand U1383 (N_1383,In_2725,In_637);
nor U1384 (N_1384,In_1378,In_1410);
nand U1385 (N_1385,In_2669,In_1277);
and U1386 (N_1386,In_2896,In_1654);
xor U1387 (N_1387,In_392,In_124);
nand U1388 (N_1388,In_1000,In_928);
or U1389 (N_1389,In_1689,In_14);
xor U1390 (N_1390,In_898,In_661);
and U1391 (N_1391,In_2866,In_1253);
and U1392 (N_1392,In_2092,In_1992);
nand U1393 (N_1393,In_2706,In_1469);
nand U1394 (N_1394,In_1728,In_2308);
and U1395 (N_1395,In_756,In_2224);
nor U1396 (N_1396,In_995,In_570);
nor U1397 (N_1397,In_2799,In_726);
nor U1398 (N_1398,In_1514,In_2875);
and U1399 (N_1399,In_1306,In_739);
xor U1400 (N_1400,In_767,In_2770);
xnor U1401 (N_1401,In_1745,In_414);
nand U1402 (N_1402,In_130,In_204);
nand U1403 (N_1403,In_1204,In_2210);
nor U1404 (N_1404,In_2298,In_1705);
and U1405 (N_1405,In_2500,In_1499);
or U1406 (N_1406,In_2584,In_275);
and U1407 (N_1407,In_1543,In_1103);
or U1408 (N_1408,In_2470,In_2012);
xor U1409 (N_1409,In_1262,In_1633);
and U1410 (N_1410,In_175,In_299);
and U1411 (N_1411,In_1659,In_1285);
or U1412 (N_1412,In_783,In_10);
nand U1413 (N_1413,In_772,In_1962);
nand U1414 (N_1414,In_2122,In_1394);
nor U1415 (N_1415,In_462,In_1555);
nor U1416 (N_1416,In_2293,In_1580);
and U1417 (N_1417,In_1344,In_2430);
and U1418 (N_1418,In_668,In_2986);
and U1419 (N_1419,In_1853,In_1521);
nor U1420 (N_1420,In_2125,In_36);
nand U1421 (N_1421,In_2621,In_1939);
xnor U1422 (N_1422,In_2189,In_1867);
nor U1423 (N_1423,In_1590,In_952);
or U1424 (N_1424,In_1173,In_2540);
nor U1425 (N_1425,In_2404,In_968);
xnor U1426 (N_1426,In_1214,In_1352);
and U1427 (N_1427,In_1729,In_987);
nor U1428 (N_1428,In_2381,In_862);
nand U1429 (N_1429,In_193,In_2303);
and U1430 (N_1430,In_2406,In_674);
and U1431 (N_1431,In_1626,In_1941);
xnor U1432 (N_1432,In_2305,In_742);
nor U1433 (N_1433,In_2501,In_2718);
xor U1434 (N_1434,In_2736,In_2137);
nand U1435 (N_1435,In_1601,In_2551);
xnor U1436 (N_1436,In_1252,In_548);
or U1437 (N_1437,In_2170,In_2890);
or U1438 (N_1438,In_1408,In_1755);
or U1439 (N_1439,In_479,In_1341);
nand U1440 (N_1440,In_1163,In_1368);
nor U1441 (N_1441,In_1849,In_474);
nand U1442 (N_1442,In_1697,In_2937);
nand U1443 (N_1443,In_1530,In_2297);
nor U1444 (N_1444,In_1882,In_2417);
or U1445 (N_1445,In_2721,In_2291);
xor U1446 (N_1446,In_2742,In_1926);
and U1447 (N_1447,In_1638,In_2008);
and U1448 (N_1448,In_1005,In_256);
nor U1449 (N_1449,In_2288,In_734);
nor U1450 (N_1450,In_211,In_2211);
nand U1451 (N_1451,In_1509,In_558);
xnor U1452 (N_1452,In_113,In_2586);
nor U1453 (N_1453,In_753,In_546);
nand U1454 (N_1454,In_733,In_522);
xor U1455 (N_1455,In_1789,In_1221);
nand U1456 (N_1456,In_725,In_936);
nand U1457 (N_1457,In_2680,In_1892);
xor U1458 (N_1458,In_2543,In_945);
or U1459 (N_1459,In_2103,In_2041);
and U1460 (N_1460,In_2322,In_1260);
nor U1461 (N_1461,In_900,In_8);
nand U1462 (N_1462,In_610,In_2307);
or U1463 (N_1463,In_1484,In_2788);
nand U1464 (N_1464,In_993,In_1570);
or U1465 (N_1465,In_1582,In_1866);
nor U1466 (N_1466,In_2529,In_246);
or U1467 (N_1467,In_2364,In_2042);
nor U1468 (N_1468,In_537,In_745);
and U1469 (N_1469,In_1271,In_2356);
or U1470 (N_1470,In_1709,In_2767);
and U1471 (N_1471,In_553,In_1117);
nand U1472 (N_1472,In_1995,In_1418);
or U1473 (N_1473,In_268,In_2477);
and U1474 (N_1474,In_1342,In_2805);
nor U1475 (N_1475,In_2314,In_2067);
and U1476 (N_1476,In_1743,In_2781);
or U1477 (N_1477,In_2995,In_298);
xor U1478 (N_1478,In_2646,In_2923);
nor U1479 (N_1479,In_2412,In_148);
xor U1480 (N_1480,In_2566,In_2006);
nor U1481 (N_1481,In_2493,In_47);
or U1482 (N_1482,In_665,In_1549);
and U1483 (N_1483,In_906,In_1835);
and U1484 (N_1484,In_2848,In_2922);
and U1485 (N_1485,In_1963,In_1624);
nand U1486 (N_1486,In_51,In_2689);
nand U1487 (N_1487,In_187,In_2311);
nand U1488 (N_1488,In_687,In_2120);
nor U1489 (N_1489,In_101,In_2060);
or U1490 (N_1490,In_2806,In_1903);
xor U1491 (N_1491,In_1166,In_1668);
nand U1492 (N_1492,In_143,In_2310);
nand U1493 (N_1493,In_1579,In_332);
nor U1494 (N_1494,In_2547,In_2201);
and U1495 (N_1495,In_2218,In_524);
or U1496 (N_1496,In_2710,In_167);
or U1497 (N_1497,In_2795,In_1458);
nor U1498 (N_1498,In_1228,In_1119);
nand U1499 (N_1499,In_1873,In_2752);
and U1500 (N_1500,In_706,In_2757);
nand U1501 (N_1501,In_2750,In_2393);
nor U1502 (N_1502,In_922,In_461);
xor U1503 (N_1503,In_2039,In_1982);
and U1504 (N_1504,In_2183,In_1411);
or U1505 (N_1505,In_1879,In_869);
and U1506 (N_1506,In_198,In_1434);
and U1507 (N_1507,In_1209,In_862);
and U1508 (N_1508,In_1968,In_1601);
nand U1509 (N_1509,In_1662,In_2585);
or U1510 (N_1510,In_2731,In_1268);
and U1511 (N_1511,In_2021,In_643);
and U1512 (N_1512,In_1002,In_1956);
nand U1513 (N_1513,In_2338,In_1245);
or U1514 (N_1514,In_2144,In_703);
and U1515 (N_1515,In_2558,In_2624);
nand U1516 (N_1516,In_842,In_865);
or U1517 (N_1517,In_2530,In_2912);
and U1518 (N_1518,In_1568,In_2356);
or U1519 (N_1519,In_538,In_782);
and U1520 (N_1520,In_461,In_1492);
and U1521 (N_1521,In_1597,In_1837);
nand U1522 (N_1522,In_2443,In_2139);
or U1523 (N_1523,In_269,In_30);
or U1524 (N_1524,In_1736,In_2568);
xor U1525 (N_1525,In_311,In_143);
nor U1526 (N_1526,In_869,In_1035);
or U1527 (N_1527,In_963,In_1420);
xnor U1528 (N_1528,In_819,In_15);
or U1529 (N_1529,In_1448,In_2310);
nor U1530 (N_1530,In_603,In_2103);
xnor U1531 (N_1531,In_2861,In_939);
and U1532 (N_1532,In_145,In_876);
or U1533 (N_1533,In_2539,In_1733);
nor U1534 (N_1534,In_1398,In_2111);
or U1535 (N_1535,In_2165,In_200);
or U1536 (N_1536,In_1672,In_2455);
xor U1537 (N_1537,In_2205,In_1055);
nor U1538 (N_1538,In_1450,In_218);
and U1539 (N_1539,In_1522,In_1930);
or U1540 (N_1540,In_1368,In_2966);
nand U1541 (N_1541,In_1376,In_960);
or U1542 (N_1542,In_1498,In_2191);
or U1543 (N_1543,In_2544,In_2373);
nand U1544 (N_1544,In_1231,In_2232);
or U1545 (N_1545,In_224,In_2304);
or U1546 (N_1546,In_2152,In_2153);
nand U1547 (N_1547,In_2054,In_1853);
or U1548 (N_1548,In_2121,In_2281);
and U1549 (N_1549,In_914,In_385);
xnor U1550 (N_1550,In_372,In_1257);
nor U1551 (N_1551,In_536,In_970);
or U1552 (N_1552,In_1434,In_620);
nor U1553 (N_1553,In_2472,In_112);
or U1554 (N_1554,In_2865,In_2601);
nor U1555 (N_1555,In_1983,In_481);
xnor U1556 (N_1556,In_280,In_901);
or U1557 (N_1557,In_2369,In_1599);
nor U1558 (N_1558,In_2710,In_90);
xnor U1559 (N_1559,In_2228,In_2451);
or U1560 (N_1560,In_2740,In_467);
nor U1561 (N_1561,In_2421,In_1907);
nor U1562 (N_1562,In_2727,In_522);
nand U1563 (N_1563,In_2603,In_2952);
nor U1564 (N_1564,In_1835,In_2274);
xnor U1565 (N_1565,In_1802,In_1825);
xor U1566 (N_1566,In_392,In_1621);
or U1567 (N_1567,In_485,In_1027);
xnor U1568 (N_1568,In_504,In_1743);
and U1569 (N_1569,In_2430,In_2092);
xnor U1570 (N_1570,In_1510,In_1177);
and U1571 (N_1571,In_1245,In_2777);
xnor U1572 (N_1572,In_2801,In_2519);
xor U1573 (N_1573,In_677,In_1841);
or U1574 (N_1574,In_2223,In_2074);
xor U1575 (N_1575,In_2945,In_2439);
xnor U1576 (N_1576,In_2971,In_1368);
nand U1577 (N_1577,In_1173,In_1713);
xor U1578 (N_1578,In_1672,In_1220);
or U1579 (N_1579,In_2260,In_480);
xnor U1580 (N_1580,In_146,In_2695);
xor U1581 (N_1581,In_738,In_25);
or U1582 (N_1582,In_2694,In_364);
or U1583 (N_1583,In_2448,In_2699);
or U1584 (N_1584,In_2714,In_537);
nand U1585 (N_1585,In_413,In_1222);
nand U1586 (N_1586,In_599,In_1690);
nand U1587 (N_1587,In_838,In_327);
or U1588 (N_1588,In_2507,In_1385);
and U1589 (N_1589,In_1020,In_1055);
xor U1590 (N_1590,In_96,In_2878);
nor U1591 (N_1591,In_2205,In_1351);
xnor U1592 (N_1592,In_2135,In_1856);
or U1593 (N_1593,In_424,In_656);
and U1594 (N_1594,In_1292,In_1);
nand U1595 (N_1595,In_1355,In_2222);
and U1596 (N_1596,In_1798,In_1474);
or U1597 (N_1597,In_2842,In_1960);
xor U1598 (N_1598,In_282,In_2927);
xnor U1599 (N_1599,In_1205,In_493);
or U1600 (N_1600,In_1747,In_176);
and U1601 (N_1601,In_1583,In_425);
xor U1602 (N_1602,In_2422,In_1828);
nand U1603 (N_1603,In_2617,In_2577);
nor U1604 (N_1604,In_2489,In_2347);
nor U1605 (N_1605,In_2510,In_690);
nand U1606 (N_1606,In_2706,In_1287);
nand U1607 (N_1607,In_1050,In_566);
nor U1608 (N_1608,In_955,In_1561);
xnor U1609 (N_1609,In_438,In_2566);
nand U1610 (N_1610,In_847,In_2054);
nand U1611 (N_1611,In_2263,In_2553);
or U1612 (N_1612,In_2069,In_210);
nor U1613 (N_1613,In_2819,In_292);
xor U1614 (N_1614,In_2359,In_2632);
nor U1615 (N_1615,In_2149,In_1337);
nand U1616 (N_1616,In_1177,In_2106);
or U1617 (N_1617,In_2210,In_558);
xor U1618 (N_1618,In_416,In_1811);
and U1619 (N_1619,In_152,In_648);
and U1620 (N_1620,In_1538,In_2326);
and U1621 (N_1621,In_2375,In_1916);
xnor U1622 (N_1622,In_2548,In_2063);
xnor U1623 (N_1623,In_729,In_1878);
or U1624 (N_1624,In_2389,In_18);
nand U1625 (N_1625,In_2973,In_1928);
and U1626 (N_1626,In_822,In_2782);
or U1627 (N_1627,In_166,In_475);
nand U1628 (N_1628,In_669,In_1911);
nand U1629 (N_1629,In_768,In_2014);
or U1630 (N_1630,In_1420,In_1551);
nand U1631 (N_1631,In_1974,In_1992);
or U1632 (N_1632,In_947,In_2413);
nor U1633 (N_1633,In_2852,In_1599);
nor U1634 (N_1634,In_1905,In_1459);
or U1635 (N_1635,In_1986,In_1249);
nand U1636 (N_1636,In_919,In_2828);
or U1637 (N_1637,In_109,In_2248);
and U1638 (N_1638,In_614,In_387);
nor U1639 (N_1639,In_1681,In_2627);
or U1640 (N_1640,In_2575,In_2564);
nor U1641 (N_1641,In_101,In_2827);
or U1642 (N_1642,In_2337,In_1408);
nor U1643 (N_1643,In_858,In_1030);
xnor U1644 (N_1644,In_2246,In_1433);
and U1645 (N_1645,In_2802,In_1476);
and U1646 (N_1646,In_2042,In_746);
nand U1647 (N_1647,In_783,In_1017);
xnor U1648 (N_1648,In_1773,In_1379);
and U1649 (N_1649,In_1676,In_469);
nor U1650 (N_1650,In_28,In_1081);
or U1651 (N_1651,In_2287,In_2892);
or U1652 (N_1652,In_1154,In_505);
xnor U1653 (N_1653,In_390,In_2890);
or U1654 (N_1654,In_2655,In_1733);
and U1655 (N_1655,In_1990,In_304);
or U1656 (N_1656,In_57,In_714);
and U1657 (N_1657,In_1954,In_2977);
xnor U1658 (N_1658,In_2047,In_891);
nand U1659 (N_1659,In_1746,In_687);
xor U1660 (N_1660,In_1276,In_2029);
xnor U1661 (N_1661,In_769,In_2535);
or U1662 (N_1662,In_2437,In_795);
nor U1663 (N_1663,In_1060,In_178);
nor U1664 (N_1664,In_1770,In_1456);
nand U1665 (N_1665,In_482,In_2281);
nor U1666 (N_1666,In_2831,In_2053);
xor U1667 (N_1667,In_1229,In_1339);
and U1668 (N_1668,In_341,In_1749);
nor U1669 (N_1669,In_1338,In_2310);
xnor U1670 (N_1670,In_1277,In_1027);
or U1671 (N_1671,In_1176,In_396);
or U1672 (N_1672,In_2003,In_2717);
nor U1673 (N_1673,In_195,In_2539);
nor U1674 (N_1674,In_2649,In_896);
and U1675 (N_1675,In_77,In_306);
or U1676 (N_1676,In_766,In_106);
and U1677 (N_1677,In_2318,In_2881);
xor U1678 (N_1678,In_1954,In_152);
or U1679 (N_1679,In_2484,In_783);
and U1680 (N_1680,In_1728,In_651);
nand U1681 (N_1681,In_785,In_2330);
or U1682 (N_1682,In_1527,In_1043);
nor U1683 (N_1683,In_2698,In_2783);
and U1684 (N_1684,In_1913,In_763);
or U1685 (N_1685,In_567,In_2383);
and U1686 (N_1686,In_2004,In_1437);
nor U1687 (N_1687,In_1656,In_707);
or U1688 (N_1688,In_624,In_1883);
nor U1689 (N_1689,In_207,In_1664);
and U1690 (N_1690,In_1353,In_1792);
xor U1691 (N_1691,In_2591,In_2670);
nor U1692 (N_1692,In_1945,In_2480);
nor U1693 (N_1693,In_2679,In_1332);
nor U1694 (N_1694,In_2859,In_2589);
xor U1695 (N_1695,In_533,In_833);
xor U1696 (N_1696,In_728,In_2027);
or U1697 (N_1697,In_2407,In_2759);
and U1698 (N_1698,In_965,In_2308);
xor U1699 (N_1699,In_2059,In_1930);
or U1700 (N_1700,In_1936,In_1649);
nand U1701 (N_1701,In_1154,In_1283);
nand U1702 (N_1702,In_2538,In_608);
and U1703 (N_1703,In_631,In_1452);
nand U1704 (N_1704,In_1198,In_372);
and U1705 (N_1705,In_541,In_66);
nor U1706 (N_1706,In_2198,In_2865);
xor U1707 (N_1707,In_1669,In_1596);
nor U1708 (N_1708,In_1336,In_2140);
nor U1709 (N_1709,In_2501,In_1397);
xnor U1710 (N_1710,In_1944,In_2352);
or U1711 (N_1711,In_1571,In_2298);
and U1712 (N_1712,In_1423,In_1628);
or U1713 (N_1713,In_523,In_2375);
or U1714 (N_1714,In_856,In_936);
xor U1715 (N_1715,In_1020,In_2564);
nor U1716 (N_1716,In_2194,In_1196);
or U1717 (N_1717,In_1808,In_742);
or U1718 (N_1718,In_2301,In_2655);
xnor U1719 (N_1719,In_321,In_701);
or U1720 (N_1720,In_704,In_1466);
or U1721 (N_1721,In_790,In_2751);
or U1722 (N_1722,In_670,In_1408);
nand U1723 (N_1723,In_2368,In_1508);
or U1724 (N_1724,In_2755,In_695);
and U1725 (N_1725,In_446,In_1290);
or U1726 (N_1726,In_513,In_1278);
or U1727 (N_1727,In_2570,In_2013);
or U1728 (N_1728,In_739,In_2844);
nor U1729 (N_1729,In_462,In_2495);
and U1730 (N_1730,In_179,In_2853);
or U1731 (N_1731,In_2398,In_1818);
xnor U1732 (N_1732,In_1911,In_980);
or U1733 (N_1733,In_1122,In_1200);
nor U1734 (N_1734,In_1216,In_1474);
and U1735 (N_1735,In_198,In_661);
or U1736 (N_1736,In_618,In_715);
and U1737 (N_1737,In_2517,In_920);
and U1738 (N_1738,In_2954,In_1891);
or U1739 (N_1739,In_1223,In_2865);
or U1740 (N_1740,In_2923,In_51);
nand U1741 (N_1741,In_2847,In_2987);
and U1742 (N_1742,In_1352,In_1242);
nand U1743 (N_1743,In_2860,In_2906);
nor U1744 (N_1744,In_453,In_304);
or U1745 (N_1745,In_2563,In_140);
and U1746 (N_1746,In_2555,In_803);
or U1747 (N_1747,In_1928,In_2480);
xor U1748 (N_1748,In_21,In_1624);
xor U1749 (N_1749,In_2924,In_2986);
xor U1750 (N_1750,In_2853,In_330);
or U1751 (N_1751,In_2276,In_844);
nand U1752 (N_1752,In_2243,In_2823);
nand U1753 (N_1753,In_2294,In_2043);
and U1754 (N_1754,In_1439,In_1585);
nor U1755 (N_1755,In_1314,In_1531);
xnor U1756 (N_1756,In_2977,In_260);
nand U1757 (N_1757,In_1645,In_525);
xor U1758 (N_1758,In_1210,In_1634);
nand U1759 (N_1759,In_2970,In_2640);
or U1760 (N_1760,In_1778,In_684);
xor U1761 (N_1761,In_2815,In_701);
nor U1762 (N_1762,In_726,In_2781);
or U1763 (N_1763,In_713,In_1636);
and U1764 (N_1764,In_326,In_1769);
xnor U1765 (N_1765,In_97,In_2836);
and U1766 (N_1766,In_927,In_332);
or U1767 (N_1767,In_1115,In_874);
nand U1768 (N_1768,In_1341,In_1361);
nor U1769 (N_1769,In_2974,In_1087);
nor U1770 (N_1770,In_729,In_1074);
or U1771 (N_1771,In_599,In_1676);
or U1772 (N_1772,In_2354,In_2900);
nand U1773 (N_1773,In_440,In_345);
xnor U1774 (N_1774,In_1878,In_2637);
xnor U1775 (N_1775,In_299,In_1193);
and U1776 (N_1776,In_1759,In_1483);
xnor U1777 (N_1777,In_328,In_2832);
nor U1778 (N_1778,In_2789,In_505);
nor U1779 (N_1779,In_622,In_888);
xor U1780 (N_1780,In_1408,In_1467);
nor U1781 (N_1781,In_876,In_138);
nand U1782 (N_1782,In_304,In_2648);
nor U1783 (N_1783,In_1288,In_686);
xor U1784 (N_1784,In_171,In_1099);
or U1785 (N_1785,In_2278,In_512);
or U1786 (N_1786,In_926,In_642);
nand U1787 (N_1787,In_2562,In_2284);
xor U1788 (N_1788,In_881,In_1706);
nor U1789 (N_1789,In_1897,In_2086);
xnor U1790 (N_1790,In_346,In_1945);
xnor U1791 (N_1791,In_2790,In_1613);
and U1792 (N_1792,In_514,In_1059);
or U1793 (N_1793,In_1200,In_2936);
and U1794 (N_1794,In_1337,In_1027);
nor U1795 (N_1795,In_119,In_231);
xnor U1796 (N_1796,In_1945,In_267);
xor U1797 (N_1797,In_298,In_1656);
xor U1798 (N_1798,In_1141,In_2743);
and U1799 (N_1799,In_1694,In_153);
and U1800 (N_1800,In_1000,In_2070);
xnor U1801 (N_1801,In_2992,In_191);
or U1802 (N_1802,In_1247,In_308);
xor U1803 (N_1803,In_1645,In_489);
nor U1804 (N_1804,In_2579,In_1814);
or U1805 (N_1805,In_2713,In_1042);
and U1806 (N_1806,In_523,In_2830);
nand U1807 (N_1807,In_379,In_611);
or U1808 (N_1808,In_1064,In_2188);
or U1809 (N_1809,In_2241,In_1133);
and U1810 (N_1810,In_1161,In_1770);
xor U1811 (N_1811,In_2565,In_1787);
or U1812 (N_1812,In_2743,In_1324);
and U1813 (N_1813,In_109,In_602);
nor U1814 (N_1814,In_1128,In_1513);
and U1815 (N_1815,In_47,In_2674);
nor U1816 (N_1816,In_2725,In_194);
nand U1817 (N_1817,In_2487,In_2998);
and U1818 (N_1818,In_2875,In_803);
and U1819 (N_1819,In_1346,In_1034);
nor U1820 (N_1820,In_858,In_2650);
nor U1821 (N_1821,In_2538,In_2854);
or U1822 (N_1822,In_416,In_1012);
or U1823 (N_1823,In_1882,In_2347);
nand U1824 (N_1824,In_2267,In_726);
and U1825 (N_1825,In_1604,In_896);
or U1826 (N_1826,In_548,In_442);
nor U1827 (N_1827,In_1141,In_615);
nor U1828 (N_1828,In_411,In_2825);
or U1829 (N_1829,In_1407,In_32);
nand U1830 (N_1830,In_1245,In_1556);
xnor U1831 (N_1831,In_1984,In_704);
nor U1832 (N_1832,In_1633,In_1691);
and U1833 (N_1833,In_2175,In_2044);
xnor U1834 (N_1834,In_1661,In_2696);
or U1835 (N_1835,In_395,In_85);
or U1836 (N_1836,In_634,In_696);
nand U1837 (N_1837,In_2164,In_2503);
xnor U1838 (N_1838,In_19,In_735);
and U1839 (N_1839,In_2173,In_899);
or U1840 (N_1840,In_597,In_545);
nor U1841 (N_1841,In_2501,In_2420);
and U1842 (N_1842,In_1192,In_1296);
xor U1843 (N_1843,In_2582,In_221);
or U1844 (N_1844,In_546,In_1233);
nand U1845 (N_1845,In_1282,In_647);
or U1846 (N_1846,In_2991,In_2692);
xor U1847 (N_1847,In_1723,In_1875);
or U1848 (N_1848,In_2602,In_2738);
xnor U1849 (N_1849,In_1905,In_1121);
nand U1850 (N_1850,In_1092,In_2714);
nor U1851 (N_1851,In_2255,In_2258);
and U1852 (N_1852,In_2980,In_433);
and U1853 (N_1853,In_2895,In_1413);
nor U1854 (N_1854,In_955,In_351);
nor U1855 (N_1855,In_1755,In_368);
xor U1856 (N_1856,In_795,In_2807);
and U1857 (N_1857,In_145,In_2493);
xor U1858 (N_1858,In_1793,In_2009);
nor U1859 (N_1859,In_362,In_1415);
nor U1860 (N_1860,In_100,In_2861);
or U1861 (N_1861,In_2172,In_337);
nand U1862 (N_1862,In_373,In_339);
nor U1863 (N_1863,In_1379,In_1785);
or U1864 (N_1864,In_2439,In_639);
xnor U1865 (N_1865,In_1465,In_2943);
nand U1866 (N_1866,In_2600,In_1545);
or U1867 (N_1867,In_472,In_2565);
nand U1868 (N_1868,In_1069,In_224);
nand U1869 (N_1869,In_611,In_2908);
and U1870 (N_1870,In_567,In_2461);
nor U1871 (N_1871,In_1039,In_2238);
nor U1872 (N_1872,In_1110,In_184);
or U1873 (N_1873,In_1540,In_164);
and U1874 (N_1874,In_477,In_171);
or U1875 (N_1875,In_1155,In_301);
and U1876 (N_1876,In_511,In_2889);
nand U1877 (N_1877,In_1253,In_1460);
nor U1878 (N_1878,In_2655,In_160);
and U1879 (N_1879,In_1092,In_1387);
xor U1880 (N_1880,In_520,In_1468);
nor U1881 (N_1881,In_1284,In_2434);
nand U1882 (N_1882,In_1396,In_2687);
xnor U1883 (N_1883,In_917,In_1124);
nand U1884 (N_1884,In_2747,In_146);
nand U1885 (N_1885,In_2976,In_419);
and U1886 (N_1886,In_2757,In_2161);
nor U1887 (N_1887,In_42,In_2793);
nor U1888 (N_1888,In_1135,In_534);
and U1889 (N_1889,In_2144,In_841);
nand U1890 (N_1890,In_948,In_1511);
xor U1891 (N_1891,In_1111,In_461);
nor U1892 (N_1892,In_1749,In_1531);
or U1893 (N_1893,In_1822,In_817);
and U1894 (N_1894,In_1631,In_2170);
and U1895 (N_1895,In_858,In_1889);
and U1896 (N_1896,In_893,In_1569);
nor U1897 (N_1897,In_211,In_1884);
nor U1898 (N_1898,In_551,In_948);
or U1899 (N_1899,In_2560,In_905);
xor U1900 (N_1900,In_634,In_1923);
nor U1901 (N_1901,In_2011,In_1906);
nand U1902 (N_1902,In_1194,In_1898);
xnor U1903 (N_1903,In_2755,In_800);
and U1904 (N_1904,In_1308,In_2653);
nor U1905 (N_1905,In_1513,In_1326);
or U1906 (N_1906,In_2553,In_1436);
nand U1907 (N_1907,In_390,In_779);
or U1908 (N_1908,In_1192,In_2894);
or U1909 (N_1909,In_1267,In_864);
nor U1910 (N_1910,In_34,In_2850);
nor U1911 (N_1911,In_158,In_1619);
or U1912 (N_1912,In_849,In_298);
and U1913 (N_1913,In_837,In_339);
and U1914 (N_1914,In_1948,In_360);
nand U1915 (N_1915,In_712,In_1122);
and U1916 (N_1916,In_2896,In_2079);
and U1917 (N_1917,In_150,In_1376);
and U1918 (N_1918,In_1420,In_285);
or U1919 (N_1919,In_1024,In_416);
xnor U1920 (N_1920,In_626,In_1171);
nor U1921 (N_1921,In_2761,In_2731);
nor U1922 (N_1922,In_2674,In_514);
nand U1923 (N_1923,In_1540,In_560);
nand U1924 (N_1924,In_2155,In_2973);
and U1925 (N_1925,In_1742,In_641);
xnor U1926 (N_1926,In_1566,In_795);
nand U1927 (N_1927,In_1891,In_2112);
and U1928 (N_1928,In_2807,In_236);
nand U1929 (N_1929,In_1030,In_397);
or U1930 (N_1930,In_2567,In_2179);
nor U1931 (N_1931,In_1401,In_2284);
and U1932 (N_1932,In_1509,In_2868);
and U1933 (N_1933,In_2966,In_1806);
nand U1934 (N_1934,In_2404,In_681);
and U1935 (N_1935,In_219,In_1960);
nor U1936 (N_1936,In_1776,In_2175);
nand U1937 (N_1937,In_2964,In_2411);
and U1938 (N_1938,In_1460,In_1912);
and U1939 (N_1939,In_695,In_2077);
nor U1940 (N_1940,In_221,In_1583);
xnor U1941 (N_1941,In_2912,In_1898);
xnor U1942 (N_1942,In_2103,In_1969);
nor U1943 (N_1943,In_2597,In_151);
and U1944 (N_1944,In_241,In_1489);
and U1945 (N_1945,In_885,In_309);
or U1946 (N_1946,In_2854,In_1752);
nor U1947 (N_1947,In_244,In_1819);
xor U1948 (N_1948,In_2322,In_762);
nand U1949 (N_1949,In_86,In_2647);
nand U1950 (N_1950,In_2564,In_766);
and U1951 (N_1951,In_1786,In_1446);
and U1952 (N_1952,In_2872,In_2967);
nor U1953 (N_1953,In_1847,In_715);
nor U1954 (N_1954,In_335,In_1661);
and U1955 (N_1955,In_654,In_2079);
nand U1956 (N_1956,In_857,In_1674);
and U1957 (N_1957,In_556,In_2038);
nand U1958 (N_1958,In_2772,In_2963);
nor U1959 (N_1959,In_1367,In_2466);
and U1960 (N_1960,In_195,In_484);
nor U1961 (N_1961,In_1095,In_2277);
nand U1962 (N_1962,In_2485,In_1207);
or U1963 (N_1963,In_2464,In_2637);
nand U1964 (N_1964,In_1538,In_2445);
and U1965 (N_1965,In_2164,In_2105);
nor U1966 (N_1966,In_2283,In_656);
nand U1967 (N_1967,In_505,In_2359);
nand U1968 (N_1968,In_2529,In_477);
or U1969 (N_1969,In_428,In_514);
nand U1970 (N_1970,In_866,In_482);
or U1971 (N_1971,In_1481,In_1617);
or U1972 (N_1972,In_2536,In_2939);
and U1973 (N_1973,In_2388,In_2175);
nor U1974 (N_1974,In_282,In_429);
nor U1975 (N_1975,In_1640,In_1471);
nand U1976 (N_1976,In_673,In_249);
nor U1977 (N_1977,In_1273,In_360);
and U1978 (N_1978,In_2198,In_1387);
nand U1979 (N_1979,In_2370,In_2203);
and U1980 (N_1980,In_1225,In_2314);
xor U1981 (N_1981,In_115,In_114);
xnor U1982 (N_1982,In_1599,In_127);
nor U1983 (N_1983,In_1585,In_556);
or U1984 (N_1984,In_2428,In_239);
xor U1985 (N_1985,In_251,In_2107);
nor U1986 (N_1986,In_2893,In_600);
nor U1987 (N_1987,In_1299,In_1726);
and U1988 (N_1988,In_1678,In_2876);
and U1989 (N_1989,In_1835,In_2925);
and U1990 (N_1990,In_2202,In_2900);
nor U1991 (N_1991,In_365,In_2510);
nand U1992 (N_1992,In_2919,In_1177);
and U1993 (N_1993,In_1841,In_367);
nor U1994 (N_1994,In_1192,In_545);
nand U1995 (N_1995,In_1393,In_498);
or U1996 (N_1996,In_2527,In_1245);
nor U1997 (N_1997,In_1605,In_523);
xor U1998 (N_1998,In_1229,In_2698);
nand U1999 (N_1999,In_2079,In_2821);
xnor U2000 (N_2000,In_2061,In_2047);
xor U2001 (N_2001,In_1643,In_2559);
or U2002 (N_2002,In_216,In_794);
or U2003 (N_2003,In_2627,In_673);
and U2004 (N_2004,In_2498,In_172);
nand U2005 (N_2005,In_1526,In_547);
or U2006 (N_2006,In_334,In_1173);
and U2007 (N_2007,In_1120,In_492);
nor U2008 (N_2008,In_2573,In_401);
and U2009 (N_2009,In_1027,In_1877);
or U2010 (N_2010,In_2861,In_760);
nand U2011 (N_2011,In_1781,In_2584);
and U2012 (N_2012,In_1965,In_1777);
and U2013 (N_2013,In_1659,In_2737);
or U2014 (N_2014,In_1179,In_783);
or U2015 (N_2015,In_2202,In_100);
or U2016 (N_2016,In_2973,In_952);
xnor U2017 (N_2017,In_1897,In_843);
and U2018 (N_2018,In_2864,In_990);
nand U2019 (N_2019,In_2076,In_1367);
or U2020 (N_2020,In_1747,In_644);
and U2021 (N_2021,In_2225,In_915);
nand U2022 (N_2022,In_346,In_2918);
nor U2023 (N_2023,In_2266,In_636);
nand U2024 (N_2024,In_402,In_914);
xnor U2025 (N_2025,In_269,In_2239);
xor U2026 (N_2026,In_2447,In_2586);
or U2027 (N_2027,In_22,In_2900);
or U2028 (N_2028,In_133,In_966);
nand U2029 (N_2029,In_2806,In_2111);
nand U2030 (N_2030,In_1823,In_1967);
or U2031 (N_2031,In_2903,In_486);
and U2032 (N_2032,In_895,In_466);
nand U2033 (N_2033,In_1144,In_737);
nand U2034 (N_2034,In_878,In_12);
or U2035 (N_2035,In_259,In_2468);
and U2036 (N_2036,In_506,In_2971);
nor U2037 (N_2037,In_1514,In_1995);
and U2038 (N_2038,In_2840,In_2656);
nand U2039 (N_2039,In_2513,In_570);
or U2040 (N_2040,In_1915,In_2572);
or U2041 (N_2041,In_1789,In_403);
nand U2042 (N_2042,In_473,In_1466);
xnor U2043 (N_2043,In_2502,In_242);
and U2044 (N_2044,In_2717,In_789);
and U2045 (N_2045,In_2143,In_596);
nand U2046 (N_2046,In_457,In_1736);
xor U2047 (N_2047,In_1326,In_436);
or U2048 (N_2048,In_1864,In_2887);
nor U2049 (N_2049,In_1693,In_2197);
nand U2050 (N_2050,In_2680,In_60);
and U2051 (N_2051,In_2075,In_389);
nor U2052 (N_2052,In_854,In_627);
xnor U2053 (N_2053,In_1996,In_325);
and U2054 (N_2054,In_2728,In_906);
or U2055 (N_2055,In_1444,In_540);
nand U2056 (N_2056,In_1936,In_2813);
nor U2057 (N_2057,In_570,In_1278);
and U2058 (N_2058,In_1954,In_2834);
or U2059 (N_2059,In_2005,In_1269);
nor U2060 (N_2060,In_372,In_1233);
and U2061 (N_2061,In_2720,In_377);
nor U2062 (N_2062,In_1511,In_2114);
or U2063 (N_2063,In_1737,In_1456);
nor U2064 (N_2064,In_1974,In_2967);
xor U2065 (N_2065,In_1409,In_2263);
xor U2066 (N_2066,In_944,In_2227);
nand U2067 (N_2067,In_2279,In_882);
xnor U2068 (N_2068,In_2226,In_2578);
nand U2069 (N_2069,In_1500,In_552);
nand U2070 (N_2070,In_168,In_1369);
or U2071 (N_2071,In_2899,In_1634);
or U2072 (N_2072,In_2862,In_411);
and U2073 (N_2073,In_2142,In_2013);
nand U2074 (N_2074,In_2696,In_1127);
xnor U2075 (N_2075,In_425,In_926);
and U2076 (N_2076,In_2529,In_2095);
xor U2077 (N_2077,In_997,In_1149);
and U2078 (N_2078,In_1216,In_779);
or U2079 (N_2079,In_1013,In_2492);
xor U2080 (N_2080,In_1996,In_215);
and U2081 (N_2081,In_966,In_2385);
xnor U2082 (N_2082,In_1495,In_1674);
nand U2083 (N_2083,In_2882,In_1289);
or U2084 (N_2084,In_962,In_2995);
and U2085 (N_2085,In_120,In_1275);
and U2086 (N_2086,In_2632,In_1319);
nor U2087 (N_2087,In_1976,In_1470);
nor U2088 (N_2088,In_862,In_2229);
or U2089 (N_2089,In_7,In_2777);
nand U2090 (N_2090,In_577,In_2030);
nor U2091 (N_2091,In_1292,In_449);
xor U2092 (N_2092,In_2046,In_2380);
xor U2093 (N_2093,In_765,In_2894);
nand U2094 (N_2094,In_2261,In_2789);
xnor U2095 (N_2095,In_1005,In_2489);
xnor U2096 (N_2096,In_57,In_2225);
nand U2097 (N_2097,In_2495,In_994);
nand U2098 (N_2098,In_1791,In_495);
nor U2099 (N_2099,In_964,In_1935);
nand U2100 (N_2100,In_1799,In_1579);
xor U2101 (N_2101,In_2041,In_2491);
nand U2102 (N_2102,In_1697,In_2172);
nor U2103 (N_2103,In_854,In_927);
or U2104 (N_2104,In_1862,In_960);
xnor U2105 (N_2105,In_2672,In_2808);
nor U2106 (N_2106,In_2769,In_1069);
xor U2107 (N_2107,In_2938,In_1562);
and U2108 (N_2108,In_112,In_968);
and U2109 (N_2109,In_2368,In_560);
and U2110 (N_2110,In_924,In_1632);
xnor U2111 (N_2111,In_1871,In_2178);
xnor U2112 (N_2112,In_504,In_2024);
or U2113 (N_2113,In_662,In_2603);
and U2114 (N_2114,In_2768,In_2957);
xnor U2115 (N_2115,In_2961,In_935);
xor U2116 (N_2116,In_429,In_1679);
nor U2117 (N_2117,In_1822,In_792);
and U2118 (N_2118,In_2736,In_190);
or U2119 (N_2119,In_2410,In_2264);
nand U2120 (N_2120,In_1149,In_869);
or U2121 (N_2121,In_2522,In_2639);
or U2122 (N_2122,In_2079,In_1262);
or U2123 (N_2123,In_803,In_363);
nor U2124 (N_2124,In_2157,In_1744);
nand U2125 (N_2125,In_849,In_2704);
and U2126 (N_2126,In_1991,In_698);
or U2127 (N_2127,In_1941,In_1078);
nand U2128 (N_2128,In_2422,In_2873);
and U2129 (N_2129,In_255,In_2286);
or U2130 (N_2130,In_721,In_2627);
or U2131 (N_2131,In_1632,In_264);
nand U2132 (N_2132,In_684,In_2433);
and U2133 (N_2133,In_893,In_395);
nor U2134 (N_2134,In_2688,In_2257);
nor U2135 (N_2135,In_2019,In_1984);
or U2136 (N_2136,In_1301,In_2102);
nor U2137 (N_2137,In_239,In_966);
nand U2138 (N_2138,In_646,In_654);
xnor U2139 (N_2139,In_1221,In_1553);
xnor U2140 (N_2140,In_2760,In_1549);
xor U2141 (N_2141,In_2782,In_568);
nand U2142 (N_2142,In_636,In_1522);
or U2143 (N_2143,In_2857,In_2968);
or U2144 (N_2144,In_2645,In_1751);
or U2145 (N_2145,In_2789,In_883);
or U2146 (N_2146,In_2295,In_1503);
and U2147 (N_2147,In_133,In_774);
and U2148 (N_2148,In_2157,In_957);
nor U2149 (N_2149,In_2313,In_75);
nor U2150 (N_2150,In_2240,In_2957);
and U2151 (N_2151,In_1507,In_1891);
or U2152 (N_2152,In_2853,In_468);
nor U2153 (N_2153,In_2806,In_545);
xnor U2154 (N_2154,In_808,In_1299);
nor U2155 (N_2155,In_622,In_2192);
nor U2156 (N_2156,In_893,In_561);
nor U2157 (N_2157,In_651,In_2466);
xnor U2158 (N_2158,In_356,In_1012);
and U2159 (N_2159,In_2268,In_149);
nand U2160 (N_2160,In_2725,In_2890);
or U2161 (N_2161,In_1968,In_577);
xnor U2162 (N_2162,In_2934,In_2292);
nand U2163 (N_2163,In_2076,In_1948);
nand U2164 (N_2164,In_1135,In_2774);
nor U2165 (N_2165,In_2155,In_1481);
and U2166 (N_2166,In_2659,In_1188);
or U2167 (N_2167,In_164,In_1967);
nand U2168 (N_2168,In_1356,In_1995);
and U2169 (N_2169,In_1783,In_2457);
nand U2170 (N_2170,In_1174,In_1024);
nor U2171 (N_2171,In_2532,In_2919);
nor U2172 (N_2172,In_1152,In_707);
nor U2173 (N_2173,In_631,In_2823);
nor U2174 (N_2174,In_1513,In_2546);
or U2175 (N_2175,In_2296,In_1392);
nor U2176 (N_2176,In_1560,In_2807);
and U2177 (N_2177,In_1799,In_978);
nand U2178 (N_2178,In_1500,In_2339);
or U2179 (N_2179,In_1370,In_457);
xnor U2180 (N_2180,In_959,In_1293);
nor U2181 (N_2181,In_2324,In_692);
xnor U2182 (N_2182,In_731,In_787);
and U2183 (N_2183,In_2682,In_2387);
xor U2184 (N_2184,In_380,In_1305);
nand U2185 (N_2185,In_658,In_1345);
or U2186 (N_2186,In_1309,In_1564);
nor U2187 (N_2187,In_2616,In_936);
nor U2188 (N_2188,In_448,In_2484);
and U2189 (N_2189,In_839,In_1828);
nand U2190 (N_2190,In_1716,In_1774);
xor U2191 (N_2191,In_2571,In_1905);
and U2192 (N_2192,In_951,In_1316);
or U2193 (N_2193,In_417,In_55);
xnor U2194 (N_2194,In_1549,In_2913);
and U2195 (N_2195,In_165,In_2363);
nor U2196 (N_2196,In_2268,In_1373);
nor U2197 (N_2197,In_2385,In_1639);
nand U2198 (N_2198,In_2643,In_734);
or U2199 (N_2199,In_734,In_127);
nand U2200 (N_2200,In_174,In_1804);
xnor U2201 (N_2201,In_798,In_6);
nor U2202 (N_2202,In_2995,In_493);
xnor U2203 (N_2203,In_2683,In_1208);
or U2204 (N_2204,In_1245,In_1749);
xor U2205 (N_2205,In_482,In_1739);
nor U2206 (N_2206,In_2742,In_2734);
nor U2207 (N_2207,In_2436,In_1665);
or U2208 (N_2208,In_2200,In_2758);
xor U2209 (N_2209,In_1797,In_1853);
or U2210 (N_2210,In_640,In_1421);
nand U2211 (N_2211,In_1914,In_208);
nand U2212 (N_2212,In_148,In_2975);
nor U2213 (N_2213,In_543,In_2147);
nor U2214 (N_2214,In_320,In_2674);
and U2215 (N_2215,In_438,In_1260);
nor U2216 (N_2216,In_251,In_2946);
and U2217 (N_2217,In_2892,In_2930);
nor U2218 (N_2218,In_1412,In_2939);
xor U2219 (N_2219,In_2851,In_2577);
xnor U2220 (N_2220,In_827,In_2353);
nand U2221 (N_2221,In_2535,In_2975);
or U2222 (N_2222,In_696,In_2515);
or U2223 (N_2223,In_1359,In_2014);
xor U2224 (N_2224,In_2621,In_1559);
nor U2225 (N_2225,In_246,In_2533);
nor U2226 (N_2226,In_2012,In_2932);
and U2227 (N_2227,In_2127,In_2272);
nor U2228 (N_2228,In_192,In_2025);
nand U2229 (N_2229,In_1751,In_713);
nor U2230 (N_2230,In_2185,In_2634);
xnor U2231 (N_2231,In_2184,In_1556);
xor U2232 (N_2232,In_1914,In_1928);
nor U2233 (N_2233,In_1250,In_541);
or U2234 (N_2234,In_2793,In_1581);
nor U2235 (N_2235,In_2367,In_312);
and U2236 (N_2236,In_949,In_1679);
xor U2237 (N_2237,In_2457,In_1531);
or U2238 (N_2238,In_2315,In_1203);
or U2239 (N_2239,In_2742,In_678);
nor U2240 (N_2240,In_1978,In_2805);
xnor U2241 (N_2241,In_2164,In_1188);
xor U2242 (N_2242,In_689,In_1853);
xnor U2243 (N_2243,In_271,In_1651);
xnor U2244 (N_2244,In_192,In_159);
and U2245 (N_2245,In_468,In_1769);
and U2246 (N_2246,In_555,In_854);
nand U2247 (N_2247,In_1885,In_659);
or U2248 (N_2248,In_832,In_1940);
xnor U2249 (N_2249,In_549,In_1814);
nor U2250 (N_2250,In_954,In_1322);
or U2251 (N_2251,In_2847,In_1831);
nand U2252 (N_2252,In_2460,In_2683);
nand U2253 (N_2253,In_534,In_153);
and U2254 (N_2254,In_1727,In_1250);
nand U2255 (N_2255,In_1908,In_1633);
or U2256 (N_2256,In_1448,In_1799);
or U2257 (N_2257,In_1185,In_1296);
and U2258 (N_2258,In_686,In_2290);
xnor U2259 (N_2259,In_774,In_2609);
nand U2260 (N_2260,In_2784,In_2553);
and U2261 (N_2261,In_753,In_2870);
nor U2262 (N_2262,In_2841,In_1808);
nor U2263 (N_2263,In_759,In_2717);
xnor U2264 (N_2264,In_2142,In_2269);
nand U2265 (N_2265,In_2841,In_2313);
or U2266 (N_2266,In_2630,In_2421);
nand U2267 (N_2267,In_2144,In_2896);
nand U2268 (N_2268,In_2259,In_412);
or U2269 (N_2269,In_610,In_2105);
xnor U2270 (N_2270,In_342,In_229);
nand U2271 (N_2271,In_2254,In_2257);
nand U2272 (N_2272,In_154,In_765);
and U2273 (N_2273,In_597,In_586);
and U2274 (N_2274,In_143,In_1920);
nor U2275 (N_2275,In_2152,In_1648);
or U2276 (N_2276,In_1121,In_1519);
nand U2277 (N_2277,In_2071,In_250);
xnor U2278 (N_2278,In_121,In_1125);
nor U2279 (N_2279,In_1716,In_299);
nand U2280 (N_2280,In_2388,In_741);
nand U2281 (N_2281,In_2158,In_1221);
nor U2282 (N_2282,In_866,In_860);
and U2283 (N_2283,In_2654,In_2737);
and U2284 (N_2284,In_1920,In_1633);
xor U2285 (N_2285,In_840,In_552);
and U2286 (N_2286,In_1621,In_103);
xor U2287 (N_2287,In_390,In_2811);
and U2288 (N_2288,In_1843,In_1014);
nor U2289 (N_2289,In_1766,In_1758);
nor U2290 (N_2290,In_2764,In_1513);
xor U2291 (N_2291,In_2025,In_1122);
xnor U2292 (N_2292,In_208,In_2861);
nor U2293 (N_2293,In_2906,In_559);
nand U2294 (N_2294,In_2010,In_2595);
xnor U2295 (N_2295,In_124,In_1930);
xnor U2296 (N_2296,In_766,In_1348);
nand U2297 (N_2297,In_2822,In_2941);
or U2298 (N_2298,In_493,In_2001);
or U2299 (N_2299,In_2883,In_980);
nor U2300 (N_2300,In_1111,In_2295);
or U2301 (N_2301,In_2029,In_1122);
or U2302 (N_2302,In_2539,In_1076);
nor U2303 (N_2303,In_257,In_379);
and U2304 (N_2304,In_2101,In_707);
xor U2305 (N_2305,In_2791,In_2655);
xor U2306 (N_2306,In_2066,In_1516);
and U2307 (N_2307,In_2932,In_49);
xor U2308 (N_2308,In_2371,In_297);
or U2309 (N_2309,In_1386,In_1565);
and U2310 (N_2310,In_2697,In_1056);
nor U2311 (N_2311,In_1552,In_258);
nand U2312 (N_2312,In_2029,In_250);
nand U2313 (N_2313,In_81,In_1542);
or U2314 (N_2314,In_1445,In_1511);
nor U2315 (N_2315,In_597,In_377);
nor U2316 (N_2316,In_2949,In_1218);
and U2317 (N_2317,In_2526,In_326);
nor U2318 (N_2318,In_2092,In_570);
and U2319 (N_2319,In_1214,In_150);
nor U2320 (N_2320,In_1181,In_2909);
nand U2321 (N_2321,In_1511,In_1042);
nand U2322 (N_2322,In_655,In_2836);
nand U2323 (N_2323,In_1234,In_220);
xor U2324 (N_2324,In_75,In_1862);
nand U2325 (N_2325,In_2129,In_225);
nor U2326 (N_2326,In_1923,In_2708);
xor U2327 (N_2327,In_543,In_1978);
nor U2328 (N_2328,In_179,In_2616);
xnor U2329 (N_2329,In_1321,In_1219);
xnor U2330 (N_2330,In_1569,In_2390);
nor U2331 (N_2331,In_165,In_2876);
or U2332 (N_2332,In_1783,In_2231);
and U2333 (N_2333,In_1901,In_2502);
xor U2334 (N_2334,In_789,In_2293);
and U2335 (N_2335,In_1129,In_2082);
xnor U2336 (N_2336,In_2310,In_2119);
nand U2337 (N_2337,In_2886,In_2611);
xor U2338 (N_2338,In_1521,In_2827);
or U2339 (N_2339,In_2875,In_1820);
or U2340 (N_2340,In_1305,In_2848);
xnor U2341 (N_2341,In_1016,In_1270);
nand U2342 (N_2342,In_843,In_565);
and U2343 (N_2343,In_1516,In_1247);
or U2344 (N_2344,In_2171,In_871);
or U2345 (N_2345,In_1158,In_2537);
nor U2346 (N_2346,In_695,In_745);
and U2347 (N_2347,In_861,In_2256);
and U2348 (N_2348,In_1549,In_2477);
xor U2349 (N_2349,In_669,In_1087);
xor U2350 (N_2350,In_836,In_75);
xnor U2351 (N_2351,In_1400,In_1712);
xnor U2352 (N_2352,In_2633,In_982);
xor U2353 (N_2353,In_709,In_2075);
and U2354 (N_2354,In_1223,In_1204);
nand U2355 (N_2355,In_1660,In_2136);
and U2356 (N_2356,In_2448,In_2122);
nand U2357 (N_2357,In_2266,In_1709);
or U2358 (N_2358,In_454,In_1997);
nor U2359 (N_2359,In_1384,In_1323);
or U2360 (N_2360,In_483,In_2051);
or U2361 (N_2361,In_1501,In_2285);
xnor U2362 (N_2362,In_2242,In_2420);
and U2363 (N_2363,In_646,In_1504);
and U2364 (N_2364,In_229,In_1853);
xnor U2365 (N_2365,In_2780,In_686);
nand U2366 (N_2366,In_2506,In_1949);
and U2367 (N_2367,In_2940,In_2203);
nand U2368 (N_2368,In_1736,In_1959);
nor U2369 (N_2369,In_795,In_2100);
nor U2370 (N_2370,In_342,In_161);
and U2371 (N_2371,In_2964,In_1242);
nand U2372 (N_2372,In_1611,In_2583);
nand U2373 (N_2373,In_122,In_974);
xnor U2374 (N_2374,In_2908,In_274);
and U2375 (N_2375,In_2508,In_2120);
or U2376 (N_2376,In_1628,In_495);
nor U2377 (N_2377,In_1399,In_2675);
xnor U2378 (N_2378,In_2853,In_719);
xnor U2379 (N_2379,In_1228,In_639);
and U2380 (N_2380,In_2992,In_1974);
nor U2381 (N_2381,In_2738,In_9);
nor U2382 (N_2382,In_457,In_2591);
nand U2383 (N_2383,In_1531,In_2348);
nand U2384 (N_2384,In_1263,In_1071);
nor U2385 (N_2385,In_688,In_1731);
nand U2386 (N_2386,In_2878,In_1159);
nor U2387 (N_2387,In_998,In_2629);
nand U2388 (N_2388,In_2986,In_1232);
and U2389 (N_2389,In_382,In_1995);
xnor U2390 (N_2390,In_1501,In_138);
and U2391 (N_2391,In_1066,In_1668);
nor U2392 (N_2392,In_1145,In_605);
or U2393 (N_2393,In_1550,In_781);
xor U2394 (N_2394,In_1808,In_277);
and U2395 (N_2395,In_663,In_401);
or U2396 (N_2396,In_1349,In_157);
or U2397 (N_2397,In_1332,In_1404);
nand U2398 (N_2398,In_1557,In_1552);
xor U2399 (N_2399,In_461,In_2150);
nand U2400 (N_2400,In_546,In_1109);
nand U2401 (N_2401,In_1671,In_1974);
and U2402 (N_2402,In_2729,In_2138);
xnor U2403 (N_2403,In_488,In_294);
xor U2404 (N_2404,In_2394,In_449);
and U2405 (N_2405,In_1948,In_801);
xor U2406 (N_2406,In_2807,In_2826);
xnor U2407 (N_2407,In_386,In_1810);
or U2408 (N_2408,In_669,In_1920);
and U2409 (N_2409,In_2581,In_2005);
nand U2410 (N_2410,In_1277,In_1947);
or U2411 (N_2411,In_333,In_2352);
and U2412 (N_2412,In_1540,In_2449);
or U2413 (N_2413,In_2259,In_1592);
or U2414 (N_2414,In_1277,In_1901);
nand U2415 (N_2415,In_1757,In_138);
nand U2416 (N_2416,In_1747,In_419);
or U2417 (N_2417,In_2994,In_425);
or U2418 (N_2418,In_389,In_2174);
and U2419 (N_2419,In_2512,In_2202);
xor U2420 (N_2420,In_1433,In_1067);
xor U2421 (N_2421,In_2713,In_2100);
nand U2422 (N_2422,In_1814,In_534);
nor U2423 (N_2423,In_1194,In_2911);
nand U2424 (N_2424,In_2377,In_1035);
or U2425 (N_2425,In_2102,In_818);
nand U2426 (N_2426,In_958,In_2285);
or U2427 (N_2427,In_1904,In_2857);
nor U2428 (N_2428,In_585,In_2005);
and U2429 (N_2429,In_2,In_1151);
nor U2430 (N_2430,In_2729,In_104);
and U2431 (N_2431,In_1894,In_1226);
nand U2432 (N_2432,In_845,In_137);
or U2433 (N_2433,In_185,In_1031);
xnor U2434 (N_2434,In_2605,In_2264);
or U2435 (N_2435,In_226,In_614);
nand U2436 (N_2436,In_2905,In_2961);
nand U2437 (N_2437,In_1960,In_2948);
nand U2438 (N_2438,In_1519,In_2647);
and U2439 (N_2439,In_1759,In_1613);
and U2440 (N_2440,In_882,In_2314);
xor U2441 (N_2441,In_849,In_593);
nand U2442 (N_2442,In_2236,In_2264);
nand U2443 (N_2443,In_1200,In_2394);
xnor U2444 (N_2444,In_639,In_2812);
and U2445 (N_2445,In_417,In_537);
nand U2446 (N_2446,In_1376,In_531);
nor U2447 (N_2447,In_2409,In_1143);
xor U2448 (N_2448,In_866,In_2283);
xor U2449 (N_2449,In_1537,In_997);
and U2450 (N_2450,In_2848,In_1866);
or U2451 (N_2451,In_144,In_2900);
xnor U2452 (N_2452,In_2629,In_2584);
or U2453 (N_2453,In_239,In_2577);
and U2454 (N_2454,In_2674,In_1462);
or U2455 (N_2455,In_1336,In_653);
nand U2456 (N_2456,In_90,In_857);
xor U2457 (N_2457,In_1996,In_2605);
nor U2458 (N_2458,In_940,In_116);
or U2459 (N_2459,In_2996,In_2359);
and U2460 (N_2460,In_766,In_702);
and U2461 (N_2461,In_2775,In_551);
and U2462 (N_2462,In_661,In_2790);
and U2463 (N_2463,In_1026,In_662);
nand U2464 (N_2464,In_1460,In_1295);
and U2465 (N_2465,In_463,In_1937);
nor U2466 (N_2466,In_2362,In_1798);
and U2467 (N_2467,In_2021,In_1366);
nand U2468 (N_2468,In_95,In_1274);
nand U2469 (N_2469,In_1018,In_616);
nor U2470 (N_2470,In_2155,In_888);
and U2471 (N_2471,In_30,In_1267);
xnor U2472 (N_2472,In_1875,In_1228);
nor U2473 (N_2473,In_405,In_296);
and U2474 (N_2474,In_1114,In_960);
or U2475 (N_2475,In_863,In_1051);
and U2476 (N_2476,In_1188,In_2876);
nor U2477 (N_2477,In_1244,In_2754);
nand U2478 (N_2478,In_1049,In_581);
xor U2479 (N_2479,In_1164,In_2669);
and U2480 (N_2480,In_1387,In_2098);
nor U2481 (N_2481,In_138,In_1891);
or U2482 (N_2482,In_726,In_680);
and U2483 (N_2483,In_1936,In_1094);
nor U2484 (N_2484,In_2994,In_110);
nand U2485 (N_2485,In_1598,In_2998);
and U2486 (N_2486,In_2705,In_1193);
nor U2487 (N_2487,In_441,In_1262);
or U2488 (N_2488,In_348,In_2814);
nand U2489 (N_2489,In_1841,In_1677);
xor U2490 (N_2490,In_1965,In_2158);
nand U2491 (N_2491,In_1063,In_648);
nand U2492 (N_2492,In_1107,In_2824);
and U2493 (N_2493,In_789,In_67);
or U2494 (N_2494,In_1226,In_1019);
or U2495 (N_2495,In_2040,In_2547);
or U2496 (N_2496,In_586,In_1809);
nor U2497 (N_2497,In_1442,In_620);
or U2498 (N_2498,In_388,In_191);
or U2499 (N_2499,In_2759,In_908);
or U2500 (N_2500,In_1750,In_958);
xnor U2501 (N_2501,In_90,In_2600);
nand U2502 (N_2502,In_356,In_2632);
xnor U2503 (N_2503,In_2573,In_45);
nor U2504 (N_2504,In_2901,In_840);
nand U2505 (N_2505,In_1559,In_1881);
xnor U2506 (N_2506,In_2836,In_2811);
nand U2507 (N_2507,In_2256,In_816);
nor U2508 (N_2508,In_1987,In_516);
nand U2509 (N_2509,In_1669,In_2920);
xnor U2510 (N_2510,In_2034,In_667);
or U2511 (N_2511,In_4,In_516);
nand U2512 (N_2512,In_1026,In_589);
xnor U2513 (N_2513,In_1267,In_2403);
and U2514 (N_2514,In_2051,In_2997);
nand U2515 (N_2515,In_99,In_276);
and U2516 (N_2516,In_547,In_6);
nand U2517 (N_2517,In_58,In_2675);
nor U2518 (N_2518,In_1947,In_1631);
or U2519 (N_2519,In_2586,In_979);
and U2520 (N_2520,In_2099,In_2920);
xnor U2521 (N_2521,In_2070,In_1873);
nor U2522 (N_2522,In_2347,In_339);
or U2523 (N_2523,In_544,In_1921);
nand U2524 (N_2524,In_2727,In_1086);
xnor U2525 (N_2525,In_142,In_1271);
nor U2526 (N_2526,In_1105,In_2610);
and U2527 (N_2527,In_746,In_1615);
or U2528 (N_2528,In_2212,In_2293);
or U2529 (N_2529,In_2804,In_5);
and U2530 (N_2530,In_1968,In_2736);
xnor U2531 (N_2531,In_2036,In_5);
or U2532 (N_2532,In_726,In_1154);
nand U2533 (N_2533,In_2659,In_1525);
nand U2534 (N_2534,In_2589,In_2380);
or U2535 (N_2535,In_1537,In_2118);
xor U2536 (N_2536,In_2487,In_1335);
or U2537 (N_2537,In_2683,In_788);
nand U2538 (N_2538,In_2018,In_2718);
nor U2539 (N_2539,In_1243,In_1947);
or U2540 (N_2540,In_1653,In_2117);
nand U2541 (N_2541,In_737,In_2650);
or U2542 (N_2542,In_2228,In_650);
nor U2543 (N_2543,In_2758,In_265);
xor U2544 (N_2544,In_556,In_489);
xor U2545 (N_2545,In_1248,In_531);
xor U2546 (N_2546,In_407,In_1768);
or U2547 (N_2547,In_816,In_2041);
xor U2548 (N_2548,In_2728,In_2944);
or U2549 (N_2549,In_461,In_1766);
and U2550 (N_2550,In_1280,In_1565);
nand U2551 (N_2551,In_2938,In_200);
nand U2552 (N_2552,In_2341,In_1015);
nor U2553 (N_2553,In_2785,In_1056);
xnor U2554 (N_2554,In_469,In_1034);
nand U2555 (N_2555,In_1266,In_1461);
nand U2556 (N_2556,In_2509,In_1299);
xor U2557 (N_2557,In_2387,In_537);
xor U2558 (N_2558,In_2595,In_573);
or U2559 (N_2559,In_614,In_1953);
xnor U2560 (N_2560,In_166,In_1631);
or U2561 (N_2561,In_1675,In_2176);
nor U2562 (N_2562,In_441,In_1280);
nand U2563 (N_2563,In_214,In_517);
and U2564 (N_2564,In_478,In_1394);
xor U2565 (N_2565,In_1340,In_172);
nand U2566 (N_2566,In_4,In_2507);
nor U2567 (N_2567,In_2128,In_1464);
or U2568 (N_2568,In_222,In_2373);
and U2569 (N_2569,In_1635,In_725);
nor U2570 (N_2570,In_1863,In_2228);
nor U2571 (N_2571,In_494,In_724);
nor U2572 (N_2572,In_473,In_1312);
nor U2573 (N_2573,In_1825,In_1200);
nor U2574 (N_2574,In_1850,In_562);
or U2575 (N_2575,In_1859,In_782);
nand U2576 (N_2576,In_2982,In_301);
nand U2577 (N_2577,In_2336,In_2276);
nand U2578 (N_2578,In_2711,In_1830);
nor U2579 (N_2579,In_2849,In_1467);
nand U2580 (N_2580,In_2217,In_1405);
nand U2581 (N_2581,In_1281,In_1003);
nor U2582 (N_2582,In_1643,In_1036);
nand U2583 (N_2583,In_1727,In_2561);
or U2584 (N_2584,In_369,In_1909);
xor U2585 (N_2585,In_2787,In_90);
nand U2586 (N_2586,In_1861,In_1062);
or U2587 (N_2587,In_2809,In_799);
nand U2588 (N_2588,In_1832,In_640);
xor U2589 (N_2589,In_1972,In_1960);
or U2590 (N_2590,In_2042,In_1539);
xor U2591 (N_2591,In_305,In_1081);
or U2592 (N_2592,In_2851,In_2988);
and U2593 (N_2593,In_2990,In_1640);
and U2594 (N_2594,In_2214,In_2008);
or U2595 (N_2595,In_1697,In_1277);
nor U2596 (N_2596,In_1096,In_1125);
nor U2597 (N_2597,In_13,In_653);
and U2598 (N_2598,In_1046,In_877);
or U2599 (N_2599,In_124,In_2245);
or U2600 (N_2600,In_2431,In_115);
nand U2601 (N_2601,In_1184,In_1276);
nand U2602 (N_2602,In_2310,In_130);
xnor U2603 (N_2603,In_254,In_2512);
and U2604 (N_2604,In_971,In_1931);
nand U2605 (N_2605,In_382,In_1531);
xor U2606 (N_2606,In_133,In_1386);
nor U2607 (N_2607,In_597,In_770);
and U2608 (N_2608,In_2870,In_1253);
xnor U2609 (N_2609,In_1046,In_649);
and U2610 (N_2610,In_1541,In_1502);
nand U2611 (N_2611,In_2231,In_1538);
or U2612 (N_2612,In_623,In_1591);
xor U2613 (N_2613,In_2234,In_1224);
xor U2614 (N_2614,In_939,In_2013);
xnor U2615 (N_2615,In_2107,In_1916);
nor U2616 (N_2616,In_583,In_198);
or U2617 (N_2617,In_1013,In_816);
nor U2618 (N_2618,In_901,In_649);
and U2619 (N_2619,In_2391,In_894);
or U2620 (N_2620,In_2638,In_769);
or U2621 (N_2621,In_101,In_1100);
nand U2622 (N_2622,In_2497,In_2056);
xor U2623 (N_2623,In_2373,In_2788);
nor U2624 (N_2624,In_488,In_1623);
or U2625 (N_2625,In_1870,In_101);
and U2626 (N_2626,In_1269,In_2106);
and U2627 (N_2627,In_413,In_1497);
nor U2628 (N_2628,In_290,In_2662);
and U2629 (N_2629,In_919,In_1509);
xor U2630 (N_2630,In_798,In_2240);
xnor U2631 (N_2631,In_117,In_2412);
or U2632 (N_2632,In_555,In_2230);
and U2633 (N_2633,In_239,In_1745);
or U2634 (N_2634,In_1422,In_9);
and U2635 (N_2635,In_2919,In_1913);
xnor U2636 (N_2636,In_2821,In_1089);
nor U2637 (N_2637,In_1062,In_1114);
or U2638 (N_2638,In_2298,In_445);
nand U2639 (N_2639,In_2392,In_78);
nand U2640 (N_2640,In_2094,In_329);
nor U2641 (N_2641,In_1178,In_1233);
and U2642 (N_2642,In_2573,In_1029);
or U2643 (N_2643,In_854,In_1967);
nor U2644 (N_2644,In_2654,In_837);
nor U2645 (N_2645,In_356,In_121);
nand U2646 (N_2646,In_954,In_1996);
or U2647 (N_2647,In_1179,In_1686);
xnor U2648 (N_2648,In_1604,In_2291);
or U2649 (N_2649,In_2556,In_2249);
nor U2650 (N_2650,In_682,In_563);
and U2651 (N_2651,In_361,In_1861);
nand U2652 (N_2652,In_1966,In_975);
nor U2653 (N_2653,In_82,In_2807);
and U2654 (N_2654,In_1762,In_868);
nand U2655 (N_2655,In_762,In_2939);
or U2656 (N_2656,In_1435,In_155);
nand U2657 (N_2657,In_267,In_1717);
and U2658 (N_2658,In_2864,In_414);
nor U2659 (N_2659,In_1941,In_2349);
or U2660 (N_2660,In_1664,In_414);
or U2661 (N_2661,In_2101,In_2468);
nor U2662 (N_2662,In_1272,In_2230);
and U2663 (N_2663,In_1305,In_66);
nand U2664 (N_2664,In_2850,In_1169);
or U2665 (N_2665,In_1432,In_580);
and U2666 (N_2666,In_84,In_2466);
xor U2667 (N_2667,In_2515,In_2491);
or U2668 (N_2668,In_2238,In_2404);
and U2669 (N_2669,In_1361,In_298);
xor U2670 (N_2670,In_1068,In_691);
nor U2671 (N_2671,In_2102,In_1087);
xor U2672 (N_2672,In_2951,In_2670);
or U2673 (N_2673,In_497,In_2419);
or U2674 (N_2674,In_145,In_110);
xor U2675 (N_2675,In_856,In_1880);
or U2676 (N_2676,In_2464,In_2285);
xnor U2677 (N_2677,In_897,In_1509);
xnor U2678 (N_2678,In_2315,In_1965);
and U2679 (N_2679,In_99,In_496);
nor U2680 (N_2680,In_2287,In_244);
and U2681 (N_2681,In_2086,In_2171);
or U2682 (N_2682,In_112,In_434);
xnor U2683 (N_2683,In_1783,In_917);
xnor U2684 (N_2684,In_2365,In_1485);
and U2685 (N_2685,In_1084,In_1966);
nand U2686 (N_2686,In_406,In_1423);
and U2687 (N_2687,In_1120,In_307);
nor U2688 (N_2688,In_1669,In_1069);
xnor U2689 (N_2689,In_2611,In_2849);
nand U2690 (N_2690,In_1766,In_2207);
nand U2691 (N_2691,In_1910,In_2545);
and U2692 (N_2692,In_1977,In_1540);
nand U2693 (N_2693,In_1310,In_2840);
nor U2694 (N_2694,In_880,In_288);
or U2695 (N_2695,In_487,In_2695);
xnor U2696 (N_2696,In_2681,In_2543);
and U2697 (N_2697,In_2940,In_851);
or U2698 (N_2698,In_2135,In_1836);
or U2699 (N_2699,In_492,In_909);
xor U2700 (N_2700,In_2482,In_1635);
xor U2701 (N_2701,In_1305,In_2289);
nand U2702 (N_2702,In_2777,In_2557);
nand U2703 (N_2703,In_2862,In_1066);
nor U2704 (N_2704,In_2775,In_1863);
or U2705 (N_2705,In_1699,In_419);
xor U2706 (N_2706,In_694,In_2512);
or U2707 (N_2707,In_2459,In_816);
xnor U2708 (N_2708,In_1309,In_339);
or U2709 (N_2709,In_2618,In_2102);
and U2710 (N_2710,In_1824,In_1130);
xnor U2711 (N_2711,In_630,In_875);
nand U2712 (N_2712,In_322,In_340);
or U2713 (N_2713,In_1607,In_2683);
nor U2714 (N_2714,In_2401,In_1243);
nand U2715 (N_2715,In_2558,In_676);
nor U2716 (N_2716,In_2437,In_1794);
and U2717 (N_2717,In_820,In_1991);
nor U2718 (N_2718,In_2494,In_2613);
nand U2719 (N_2719,In_2328,In_1684);
and U2720 (N_2720,In_2128,In_2488);
xor U2721 (N_2721,In_2144,In_2977);
nand U2722 (N_2722,In_2162,In_2620);
nand U2723 (N_2723,In_2196,In_2767);
and U2724 (N_2724,In_1377,In_2702);
and U2725 (N_2725,In_2455,In_1377);
or U2726 (N_2726,In_1521,In_2730);
xnor U2727 (N_2727,In_2829,In_545);
nor U2728 (N_2728,In_374,In_1073);
xnor U2729 (N_2729,In_625,In_2269);
and U2730 (N_2730,In_2901,In_2929);
or U2731 (N_2731,In_2343,In_1321);
or U2732 (N_2732,In_1210,In_2228);
xnor U2733 (N_2733,In_1919,In_839);
xnor U2734 (N_2734,In_133,In_2790);
xor U2735 (N_2735,In_236,In_577);
or U2736 (N_2736,In_672,In_833);
and U2737 (N_2737,In_679,In_1676);
nor U2738 (N_2738,In_2289,In_1921);
and U2739 (N_2739,In_2650,In_752);
xor U2740 (N_2740,In_1718,In_882);
xnor U2741 (N_2741,In_2517,In_1001);
xor U2742 (N_2742,In_245,In_2662);
nand U2743 (N_2743,In_2740,In_1547);
nand U2744 (N_2744,In_157,In_2640);
nand U2745 (N_2745,In_2098,In_558);
nor U2746 (N_2746,In_2356,In_1465);
xor U2747 (N_2747,In_2632,In_1410);
xor U2748 (N_2748,In_517,In_998);
nand U2749 (N_2749,In_2049,In_2167);
or U2750 (N_2750,In_2289,In_2664);
and U2751 (N_2751,In_2087,In_2811);
and U2752 (N_2752,In_2647,In_630);
or U2753 (N_2753,In_319,In_2996);
xnor U2754 (N_2754,In_2384,In_2934);
nor U2755 (N_2755,In_1060,In_2969);
or U2756 (N_2756,In_2576,In_779);
xnor U2757 (N_2757,In_2205,In_1478);
and U2758 (N_2758,In_1142,In_457);
and U2759 (N_2759,In_531,In_295);
nor U2760 (N_2760,In_2649,In_1422);
nor U2761 (N_2761,In_609,In_2665);
and U2762 (N_2762,In_439,In_1209);
xnor U2763 (N_2763,In_93,In_611);
or U2764 (N_2764,In_2510,In_1882);
nand U2765 (N_2765,In_312,In_2854);
nand U2766 (N_2766,In_2917,In_1583);
and U2767 (N_2767,In_1408,In_2014);
or U2768 (N_2768,In_522,In_2688);
or U2769 (N_2769,In_961,In_770);
and U2770 (N_2770,In_1536,In_1726);
and U2771 (N_2771,In_30,In_704);
and U2772 (N_2772,In_1636,In_2909);
and U2773 (N_2773,In_1711,In_2240);
and U2774 (N_2774,In_589,In_1147);
and U2775 (N_2775,In_2134,In_1841);
xnor U2776 (N_2776,In_732,In_2923);
or U2777 (N_2777,In_1671,In_2465);
or U2778 (N_2778,In_1807,In_1196);
nor U2779 (N_2779,In_1024,In_861);
and U2780 (N_2780,In_23,In_277);
nand U2781 (N_2781,In_2374,In_1018);
or U2782 (N_2782,In_313,In_2449);
and U2783 (N_2783,In_1406,In_1518);
and U2784 (N_2784,In_178,In_1318);
nor U2785 (N_2785,In_2865,In_1200);
xor U2786 (N_2786,In_2049,In_406);
xnor U2787 (N_2787,In_1281,In_2969);
nand U2788 (N_2788,In_630,In_18);
xnor U2789 (N_2789,In_1215,In_667);
nor U2790 (N_2790,In_510,In_1647);
nand U2791 (N_2791,In_2881,In_520);
nor U2792 (N_2792,In_1532,In_366);
or U2793 (N_2793,In_1030,In_1038);
or U2794 (N_2794,In_2534,In_588);
nor U2795 (N_2795,In_1154,In_419);
and U2796 (N_2796,In_1720,In_523);
nand U2797 (N_2797,In_2224,In_697);
nor U2798 (N_2798,In_2435,In_540);
and U2799 (N_2799,In_1198,In_2758);
nor U2800 (N_2800,In_554,In_2452);
and U2801 (N_2801,In_211,In_2977);
nor U2802 (N_2802,In_1290,In_602);
and U2803 (N_2803,In_899,In_1557);
nor U2804 (N_2804,In_2919,In_428);
or U2805 (N_2805,In_1018,In_2431);
or U2806 (N_2806,In_917,In_2133);
nor U2807 (N_2807,In_796,In_2933);
xnor U2808 (N_2808,In_29,In_1346);
and U2809 (N_2809,In_1674,In_1522);
nand U2810 (N_2810,In_2036,In_1368);
nand U2811 (N_2811,In_1063,In_363);
nor U2812 (N_2812,In_2390,In_2681);
nand U2813 (N_2813,In_1813,In_49);
or U2814 (N_2814,In_2718,In_105);
nand U2815 (N_2815,In_902,In_313);
nor U2816 (N_2816,In_337,In_2688);
or U2817 (N_2817,In_662,In_467);
nor U2818 (N_2818,In_2170,In_975);
or U2819 (N_2819,In_1538,In_1796);
and U2820 (N_2820,In_2118,In_218);
and U2821 (N_2821,In_1960,In_2969);
nand U2822 (N_2822,In_2834,In_339);
or U2823 (N_2823,In_1254,In_2054);
nand U2824 (N_2824,In_2412,In_36);
and U2825 (N_2825,In_716,In_1861);
xor U2826 (N_2826,In_1708,In_1866);
or U2827 (N_2827,In_2411,In_545);
nand U2828 (N_2828,In_1857,In_1079);
xor U2829 (N_2829,In_1376,In_2154);
and U2830 (N_2830,In_1674,In_2074);
and U2831 (N_2831,In_1872,In_126);
nand U2832 (N_2832,In_464,In_2691);
xor U2833 (N_2833,In_2072,In_1263);
nand U2834 (N_2834,In_1146,In_1490);
xor U2835 (N_2835,In_2871,In_2151);
and U2836 (N_2836,In_335,In_1565);
nor U2837 (N_2837,In_2179,In_2329);
nand U2838 (N_2838,In_1788,In_1781);
or U2839 (N_2839,In_2192,In_2485);
xnor U2840 (N_2840,In_1432,In_2968);
nor U2841 (N_2841,In_2412,In_535);
nor U2842 (N_2842,In_2494,In_605);
or U2843 (N_2843,In_1935,In_2972);
and U2844 (N_2844,In_1341,In_2422);
xnor U2845 (N_2845,In_1737,In_1851);
nor U2846 (N_2846,In_2982,In_636);
or U2847 (N_2847,In_386,In_1357);
nand U2848 (N_2848,In_1618,In_2716);
or U2849 (N_2849,In_2525,In_2150);
nor U2850 (N_2850,In_2523,In_1026);
nand U2851 (N_2851,In_933,In_2749);
and U2852 (N_2852,In_201,In_566);
and U2853 (N_2853,In_258,In_2681);
nand U2854 (N_2854,In_2259,In_886);
and U2855 (N_2855,In_985,In_264);
or U2856 (N_2856,In_2507,In_926);
or U2857 (N_2857,In_2684,In_1498);
nand U2858 (N_2858,In_2600,In_1325);
xor U2859 (N_2859,In_503,In_1347);
and U2860 (N_2860,In_2373,In_442);
or U2861 (N_2861,In_1958,In_2746);
xnor U2862 (N_2862,In_950,In_979);
nand U2863 (N_2863,In_2120,In_2777);
nand U2864 (N_2864,In_2878,In_2810);
nand U2865 (N_2865,In_1643,In_536);
or U2866 (N_2866,In_2400,In_2300);
nand U2867 (N_2867,In_2826,In_556);
and U2868 (N_2868,In_1098,In_942);
and U2869 (N_2869,In_481,In_1036);
and U2870 (N_2870,In_2654,In_1348);
nand U2871 (N_2871,In_1535,In_327);
xor U2872 (N_2872,In_151,In_55);
xor U2873 (N_2873,In_2523,In_873);
and U2874 (N_2874,In_2931,In_2571);
or U2875 (N_2875,In_235,In_2626);
or U2876 (N_2876,In_1207,In_1887);
xor U2877 (N_2877,In_2007,In_1781);
nand U2878 (N_2878,In_968,In_760);
nand U2879 (N_2879,In_2873,In_1453);
or U2880 (N_2880,In_196,In_1710);
nand U2881 (N_2881,In_150,In_70);
nand U2882 (N_2882,In_146,In_2880);
nand U2883 (N_2883,In_636,In_2488);
nor U2884 (N_2884,In_2220,In_142);
and U2885 (N_2885,In_2962,In_2324);
or U2886 (N_2886,In_131,In_2832);
nor U2887 (N_2887,In_667,In_2456);
nand U2888 (N_2888,In_8,In_2827);
or U2889 (N_2889,In_89,In_1024);
or U2890 (N_2890,In_2679,In_2410);
or U2891 (N_2891,In_497,In_2587);
nor U2892 (N_2892,In_2981,In_605);
and U2893 (N_2893,In_1654,In_1886);
or U2894 (N_2894,In_157,In_2204);
xor U2895 (N_2895,In_22,In_1045);
nor U2896 (N_2896,In_1757,In_779);
and U2897 (N_2897,In_1707,In_2006);
nor U2898 (N_2898,In_2478,In_2791);
and U2899 (N_2899,In_2494,In_320);
or U2900 (N_2900,In_236,In_934);
nand U2901 (N_2901,In_1805,In_1803);
or U2902 (N_2902,In_493,In_2115);
and U2903 (N_2903,In_2038,In_131);
nor U2904 (N_2904,In_269,In_1427);
nor U2905 (N_2905,In_1139,In_2615);
and U2906 (N_2906,In_2555,In_391);
or U2907 (N_2907,In_1202,In_505);
nand U2908 (N_2908,In_1676,In_2272);
and U2909 (N_2909,In_330,In_749);
nor U2910 (N_2910,In_1637,In_2725);
or U2911 (N_2911,In_854,In_583);
or U2912 (N_2912,In_2558,In_2187);
xor U2913 (N_2913,In_481,In_529);
nand U2914 (N_2914,In_1971,In_1024);
and U2915 (N_2915,In_2394,In_1517);
nand U2916 (N_2916,In_1192,In_1285);
nand U2917 (N_2917,In_2200,In_1311);
nor U2918 (N_2918,In_401,In_2614);
nor U2919 (N_2919,In_1092,In_1895);
xnor U2920 (N_2920,In_1881,In_2108);
or U2921 (N_2921,In_818,In_95);
nand U2922 (N_2922,In_2406,In_2351);
and U2923 (N_2923,In_292,In_2743);
or U2924 (N_2924,In_2788,In_1052);
or U2925 (N_2925,In_271,In_984);
xor U2926 (N_2926,In_702,In_2929);
nor U2927 (N_2927,In_1646,In_655);
nor U2928 (N_2928,In_1186,In_1354);
xnor U2929 (N_2929,In_2299,In_2248);
xor U2930 (N_2930,In_690,In_1253);
or U2931 (N_2931,In_1496,In_723);
and U2932 (N_2932,In_1715,In_1124);
nor U2933 (N_2933,In_39,In_499);
nor U2934 (N_2934,In_1541,In_1493);
or U2935 (N_2935,In_2720,In_2846);
and U2936 (N_2936,In_1680,In_1013);
nor U2937 (N_2937,In_1935,In_56);
xnor U2938 (N_2938,In_59,In_1711);
xnor U2939 (N_2939,In_1738,In_795);
nand U2940 (N_2940,In_2458,In_1170);
or U2941 (N_2941,In_2722,In_2588);
nand U2942 (N_2942,In_2426,In_2780);
nand U2943 (N_2943,In_1909,In_1844);
nand U2944 (N_2944,In_220,In_1712);
and U2945 (N_2945,In_2302,In_1005);
xnor U2946 (N_2946,In_2560,In_2375);
and U2947 (N_2947,In_694,In_2980);
and U2948 (N_2948,In_2054,In_218);
nand U2949 (N_2949,In_2428,In_455);
and U2950 (N_2950,In_2125,In_2311);
xnor U2951 (N_2951,In_709,In_1132);
nor U2952 (N_2952,In_359,In_1357);
nand U2953 (N_2953,In_994,In_2580);
nand U2954 (N_2954,In_374,In_2297);
xnor U2955 (N_2955,In_1560,In_1063);
or U2956 (N_2956,In_1668,In_529);
and U2957 (N_2957,In_2808,In_554);
or U2958 (N_2958,In_2013,In_2130);
and U2959 (N_2959,In_2273,In_371);
or U2960 (N_2960,In_1530,In_661);
xor U2961 (N_2961,In_756,In_2295);
nor U2962 (N_2962,In_2215,In_1681);
and U2963 (N_2963,In_2254,In_2425);
or U2964 (N_2964,In_2640,In_384);
nor U2965 (N_2965,In_1800,In_670);
xor U2966 (N_2966,In_2046,In_2501);
nor U2967 (N_2967,In_1007,In_2167);
and U2968 (N_2968,In_1911,In_2384);
or U2969 (N_2969,In_1416,In_823);
and U2970 (N_2970,In_2316,In_116);
xnor U2971 (N_2971,In_2584,In_1720);
nor U2972 (N_2972,In_2963,In_1109);
and U2973 (N_2973,In_2143,In_612);
and U2974 (N_2974,In_2428,In_2719);
or U2975 (N_2975,In_604,In_253);
or U2976 (N_2976,In_2697,In_1909);
xnor U2977 (N_2977,In_2719,In_1900);
xor U2978 (N_2978,In_2787,In_2207);
nand U2979 (N_2979,In_812,In_132);
xor U2980 (N_2980,In_455,In_1791);
nor U2981 (N_2981,In_955,In_1888);
nor U2982 (N_2982,In_632,In_572);
nor U2983 (N_2983,In_312,In_1905);
nor U2984 (N_2984,In_1817,In_2811);
or U2985 (N_2985,In_1837,In_474);
nand U2986 (N_2986,In_2506,In_625);
xnor U2987 (N_2987,In_2376,In_1078);
xnor U2988 (N_2988,In_1960,In_1237);
xnor U2989 (N_2989,In_1112,In_1876);
or U2990 (N_2990,In_1168,In_1921);
nor U2991 (N_2991,In_2247,In_2870);
nor U2992 (N_2992,In_2871,In_2565);
nor U2993 (N_2993,In_2754,In_2734);
and U2994 (N_2994,In_127,In_905);
or U2995 (N_2995,In_882,In_1905);
and U2996 (N_2996,In_761,In_461);
xor U2997 (N_2997,In_1909,In_1104);
or U2998 (N_2998,In_1840,In_2330);
xnor U2999 (N_2999,In_651,In_2138);
and U3000 (N_3000,In_2962,In_1604);
nor U3001 (N_3001,In_471,In_882);
nand U3002 (N_3002,In_2364,In_6);
xnor U3003 (N_3003,In_2289,In_2743);
nand U3004 (N_3004,In_72,In_312);
nand U3005 (N_3005,In_2644,In_1039);
and U3006 (N_3006,In_576,In_1677);
and U3007 (N_3007,In_2119,In_2016);
nand U3008 (N_3008,In_2114,In_759);
or U3009 (N_3009,In_1042,In_1954);
or U3010 (N_3010,In_147,In_1901);
nor U3011 (N_3011,In_871,In_438);
or U3012 (N_3012,In_702,In_2467);
nand U3013 (N_3013,In_1228,In_1022);
xor U3014 (N_3014,In_244,In_1545);
xnor U3015 (N_3015,In_239,In_2431);
and U3016 (N_3016,In_956,In_1398);
xor U3017 (N_3017,In_203,In_1757);
and U3018 (N_3018,In_2102,In_2101);
and U3019 (N_3019,In_654,In_2714);
nand U3020 (N_3020,In_2903,In_957);
and U3021 (N_3021,In_553,In_2392);
nand U3022 (N_3022,In_2593,In_77);
nor U3023 (N_3023,In_1637,In_1585);
and U3024 (N_3024,In_1217,In_2802);
xnor U3025 (N_3025,In_1898,In_2357);
or U3026 (N_3026,In_244,In_2076);
nor U3027 (N_3027,In_1337,In_680);
or U3028 (N_3028,In_846,In_209);
xor U3029 (N_3029,In_2683,In_1123);
nand U3030 (N_3030,In_2462,In_245);
and U3031 (N_3031,In_1666,In_2018);
or U3032 (N_3032,In_368,In_684);
or U3033 (N_3033,In_2549,In_1169);
nand U3034 (N_3034,In_391,In_859);
or U3035 (N_3035,In_377,In_2709);
or U3036 (N_3036,In_2483,In_2825);
nand U3037 (N_3037,In_2113,In_1467);
xnor U3038 (N_3038,In_2416,In_1235);
and U3039 (N_3039,In_674,In_998);
nor U3040 (N_3040,In_746,In_1703);
nand U3041 (N_3041,In_2253,In_15);
nand U3042 (N_3042,In_1731,In_1014);
or U3043 (N_3043,In_146,In_2374);
nor U3044 (N_3044,In_2772,In_362);
nor U3045 (N_3045,In_1405,In_187);
or U3046 (N_3046,In_2019,In_1891);
and U3047 (N_3047,In_2534,In_315);
and U3048 (N_3048,In_242,In_426);
and U3049 (N_3049,In_1787,In_2960);
and U3050 (N_3050,In_2385,In_277);
or U3051 (N_3051,In_1652,In_1359);
nand U3052 (N_3052,In_325,In_707);
or U3053 (N_3053,In_229,In_1741);
nor U3054 (N_3054,In_433,In_1348);
xor U3055 (N_3055,In_2446,In_1376);
nand U3056 (N_3056,In_1599,In_622);
nor U3057 (N_3057,In_921,In_2269);
nor U3058 (N_3058,In_35,In_1391);
or U3059 (N_3059,In_2406,In_2922);
xnor U3060 (N_3060,In_2087,In_1528);
nand U3061 (N_3061,In_1336,In_1797);
and U3062 (N_3062,In_819,In_1063);
nand U3063 (N_3063,In_442,In_1482);
or U3064 (N_3064,In_2178,In_1367);
or U3065 (N_3065,In_2676,In_1902);
xnor U3066 (N_3066,In_1262,In_2084);
or U3067 (N_3067,In_2134,In_2338);
nor U3068 (N_3068,In_1538,In_2045);
nor U3069 (N_3069,In_323,In_2366);
nor U3070 (N_3070,In_1143,In_2910);
and U3071 (N_3071,In_1545,In_420);
or U3072 (N_3072,In_2917,In_1040);
nor U3073 (N_3073,In_563,In_1824);
or U3074 (N_3074,In_426,In_2624);
and U3075 (N_3075,In_1778,In_762);
or U3076 (N_3076,In_2866,In_2171);
nand U3077 (N_3077,In_2348,In_78);
nand U3078 (N_3078,In_735,In_1478);
and U3079 (N_3079,In_1440,In_1297);
and U3080 (N_3080,In_2065,In_720);
and U3081 (N_3081,In_626,In_1770);
nor U3082 (N_3082,In_53,In_7);
and U3083 (N_3083,In_1532,In_1582);
or U3084 (N_3084,In_645,In_1854);
nor U3085 (N_3085,In_838,In_21);
xnor U3086 (N_3086,In_884,In_608);
nor U3087 (N_3087,In_2279,In_2656);
nor U3088 (N_3088,In_1725,In_2037);
nor U3089 (N_3089,In_1547,In_1796);
and U3090 (N_3090,In_2973,In_2280);
nand U3091 (N_3091,In_2697,In_728);
xor U3092 (N_3092,In_893,In_2106);
and U3093 (N_3093,In_126,In_2894);
nand U3094 (N_3094,In_85,In_1244);
nand U3095 (N_3095,In_2457,In_1412);
xnor U3096 (N_3096,In_1144,In_1897);
or U3097 (N_3097,In_2346,In_446);
xor U3098 (N_3098,In_1057,In_381);
and U3099 (N_3099,In_1709,In_342);
and U3100 (N_3100,In_458,In_2309);
nand U3101 (N_3101,In_2054,In_1709);
and U3102 (N_3102,In_2128,In_2978);
nor U3103 (N_3103,In_2733,In_2545);
or U3104 (N_3104,In_1451,In_1484);
xor U3105 (N_3105,In_1307,In_78);
nor U3106 (N_3106,In_2422,In_1823);
and U3107 (N_3107,In_344,In_2025);
nor U3108 (N_3108,In_696,In_2794);
and U3109 (N_3109,In_113,In_2909);
nand U3110 (N_3110,In_2663,In_932);
xor U3111 (N_3111,In_2728,In_1280);
xnor U3112 (N_3112,In_1819,In_1664);
or U3113 (N_3113,In_2822,In_661);
or U3114 (N_3114,In_2490,In_884);
nand U3115 (N_3115,In_1198,In_1660);
or U3116 (N_3116,In_2569,In_537);
or U3117 (N_3117,In_142,In_2746);
or U3118 (N_3118,In_900,In_1200);
or U3119 (N_3119,In_101,In_22);
or U3120 (N_3120,In_2331,In_2783);
or U3121 (N_3121,In_13,In_66);
and U3122 (N_3122,In_105,In_847);
or U3123 (N_3123,In_13,In_1243);
nor U3124 (N_3124,In_363,In_2640);
and U3125 (N_3125,In_2079,In_2310);
xnor U3126 (N_3126,In_930,In_1924);
nor U3127 (N_3127,In_756,In_1779);
nor U3128 (N_3128,In_392,In_320);
nand U3129 (N_3129,In_367,In_2231);
and U3130 (N_3130,In_1472,In_2486);
nand U3131 (N_3131,In_2472,In_1598);
nor U3132 (N_3132,In_2410,In_2860);
nor U3133 (N_3133,In_374,In_2420);
or U3134 (N_3134,In_1728,In_191);
xnor U3135 (N_3135,In_157,In_704);
nor U3136 (N_3136,In_2521,In_1645);
and U3137 (N_3137,In_148,In_964);
nor U3138 (N_3138,In_2180,In_837);
nor U3139 (N_3139,In_2905,In_2654);
or U3140 (N_3140,In_1042,In_42);
xor U3141 (N_3141,In_730,In_2451);
nand U3142 (N_3142,In_549,In_1265);
nand U3143 (N_3143,In_450,In_2980);
xor U3144 (N_3144,In_845,In_787);
nor U3145 (N_3145,In_2108,In_1979);
xnor U3146 (N_3146,In_2862,In_1629);
or U3147 (N_3147,In_2505,In_2775);
nand U3148 (N_3148,In_2204,In_207);
xor U3149 (N_3149,In_2036,In_165);
or U3150 (N_3150,In_2469,In_1926);
xnor U3151 (N_3151,In_1451,In_1656);
or U3152 (N_3152,In_1364,In_218);
and U3153 (N_3153,In_187,In_2577);
nor U3154 (N_3154,In_717,In_681);
xor U3155 (N_3155,In_1187,In_2766);
nor U3156 (N_3156,In_2576,In_2282);
nand U3157 (N_3157,In_2528,In_2721);
xor U3158 (N_3158,In_2979,In_1540);
xnor U3159 (N_3159,In_473,In_1386);
nor U3160 (N_3160,In_357,In_1697);
nor U3161 (N_3161,In_272,In_72);
and U3162 (N_3162,In_2111,In_1238);
or U3163 (N_3163,In_2591,In_1531);
or U3164 (N_3164,In_803,In_2600);
or U3165 (N_3165,In_66,In_2600);
nand U3166 (N_3166,In_1134,In_2940);
and U3167 (N_3167,In_816,In_1114);
or U3168 (N_3168,In_1206,In_1352);
or U3169 (N_3169,In_2446,In_119);
nand U3170 (N_3170,In_1199,In_2519);
nor U3171 (N_3171,In_2406,In_2517);
and U3172 (N_3172,In_369,In_2280);
and U3173 (N_3173,In_1749,In_584);
nand U3174 (N_3174,In_1553,In_1631);
or U3175 (N_3175,In_2768,In_2333);
nor U3176 (N_3176,In_2115,In_377);
xor U3177 (N_3177,In_2380,In_430);
nand U3178 (N_3178,In_1329,In_2649);
nand U3179 (N_3179,In_1317,In_568);
or U3180 (N_3180,In_1248,In_2145);
nand U3181 (N_3181,In_486,In_2811);
nor U3182 (N_3182,In_2623,In_1879);
nand U3183 (N_3183,In_35,In_808);
or U3184 (N_3184,In_2825,In_909);
and U3185 (N_3185,In_1136,In_1431);
or U3186 (N_3186,In_1819,In_1631);
and U3187 (N_3187,In_1566,In_238);
xnor U3188 (N_3188,In_1887,In_242);
and U3189 (N_3189,In_1930,In_2882);
nand U3190 (N_3190,In_1954,In_15);
nor U3191 (N_3191,In_1319,In_2503);
xor U3192 (N_3192,In_1911,In_40);
xor U3193 (N_3193,In_1083,In_1828);
nand U3194 (N_3194,In_1446,In_1310);
nor U3195 (N_3195,In_2715,In_794);
nor U3196 (N_3196,In_1123,In_396);
nand U3197 (N_3197,In_509,In_1174);
xor U3198 (N_3198,In_2109,In_2966);
and U3199 (N_3199,In_2912,In_1399);
or U3200 (N_3200,In_210,In_1240);
nor U3201 (N_3201,In_1248,In_1600);
nand U3202 (N_3202,In_1169,In_162);
nor U3203 (N_3203,In_137,In_1388);
nor U3204 (N_3204,In_2182,In_2956);
nand U3205 (N_3205,In_84,In_2788);
nor U3206 (N_3206,In_1310,In_2952);
nand U3207 (N_3207,In_2540,In_1482);
xnor U3208 (N_3208,In_359,In_573);
xnor U3209 (N_3209,In_1538,In_1058);
or U3210 (N_3210,In_2481,In_1283);
xor U3211 (N_3211,In_1772,In_2548);
nor U3212 (N_3212,In_1401,In_190);
and U3213 (N_3213,In_2483,In_1678);
or U3214 (N_3214,In_2920,In_242);
and U3215 (N_3215,In_1756,In_2278);
or U3216 (N_3216,In_1142,In_2028);
nor U3217 (N_3217,In_114,In_341);
and U3218 (N_3218,In_1934,In_515);
and U3219 (N_3219,In_467,In_221);
or U3220 (N_3220,In_786,In_2354);
and U3221 (N_3221,In_2101,In_1078);
nand U3222 (N_3222,In_1687,In_148);
nor U3223 (N_3223,In_1963,In_2220);
and U3224 (N_3224,In_1893,In_2801);
nand U3225 (N_3225,In_1522,In_1068);
nor U3226 (N_3226,In_1953,In_157);
nand U3227 (N_3227,In_431,In_1910);
and U3228 (N_3228,In_2256,In_2933);
nand U3229 (N_3229,In_854,In_1774);
nand U3230 (N_3230,In_906,In_261);
nand U3231 (N_3231,In_2039,In_1029);
nor U3232 (N_3232,In_194,In_408);
nor U3233 (N_3233,In_158,In_232);
and U3234 (N_3234,In_2767,In_2891);
nor U3235 (N_3235,In_2231,In_2161);
and U3236 (N_3236,In_273,In_2625);
and U3237 (N_3237,In_2644,In_405);
or U3238 (N_3238,In_1743,In_1417);
nand U3239 (N_3239,In_991,In_313);
nand U3240 (N_3240,In_1970,In_774);
nor U3241 (N_3241,In_535,In_890);
nor U3242 (N_3242,In_384,In_2336);
and U3243 (N_3243,In_1882,In_2816);
xnor U3244 (N_3244,In_2687,In_2764);
or U3245 (N_3245,In_1820,In_988);
or U3246 (N_3246,In_2119,In_488);
xor U3247 (N_3247,In_46,In_2045);
and U3248 (N_3248,In_2606,In_2642);
nand U3249 (N_3249,In_305,In_189);
or U3250 (N_3250,In_1172,In_115);
xnor U3251 (N_3251,In_1194,In_1456);
nor U3252 (N_3252,In_2610,In_1471);
or U3253 (N_3253,In_2538,In_1308);
nor U3254 (N_3254,In_900,In_1520);
and U3255 (N_3255,In_875,In_1009);
nor U3256 (N_3256,In_1808,In_103);
xor U3257 (N_3257,In_707,In_1116);
nor U3258 (N_3258,In_33,In_1542);
nor U3259 (N_3259,In_2547,In_693);
xor U3260 (N_3260,In_1176,In_1718);
xnor U3261 (N_3261,In_1395,In_820);
or U3262 (N_3262,In_2742,In_2699);
and U3263 (N_3263,In_172,In_2523);
and U3264 (N_3264,In_1705,In_1158);
or U3265 (N_3265,In_2190,In_2470);
nor U3266 (N_3266,In_2075,In_1708);
xor U3267 (N_3267,In_544,In_735);
and U3268 (N_3268,In_2058,In_2705);
nand U3269 (N_3269,In_379,In_1151);
nor U3270 (N_3270,In_1640,In_871);
nor U3271 (N_3271,In_150,In_127);
and U3272 (N_3272,In_2587,In_2795);
or U3273 (N_3273,In_594,In_2953);
xnor U3274 (N_3274,In_1735,In_1979);
xnor U3275 (N_3275,In_1505,In_2268);
nor U3276 (N_3276,In_1741,In_997);
or U3277 (N_3277,In_2985,In_1542);
nor U3278 (N_3278,In_2122,In_1950);
xnor U3279 (N_3279,In_812,In_159);
nand U3280 (N_3280,In_2547,In_911);
nor U3281 (N_3281,In_1671,In_471);
xor U3282 (N_3282,In_1531,In_191);
and U3283 (N_3283,In_457,In_1291);
nand U3284 (N_3284,In_767,In_151);
nor U3285 (N_3285,In_935,In_596);
nor U3286 (N_3286,In_3,In_2454);
and U3287 (N_3287,In_1030,In_2389);
nand U3288 (N_3288,In_2546,In_119);
nor U3289 (N_3289,In_1359,In_1307);
and U3290 (N_3290,In_2250,In_1512);
nand U3291 (N_3291,In_1031,In_2012);
xor U3292 (N_3292,In_471,In_2077);
or U3293 (N_3293,In_474,In_2315);
and U3294 (N_3294,In_1496,In_587);
xor U3295 (N_3295,In_2926,In_172);
xnor U3296 (N_3296,In_2125,In_101);
nor U3297 (N_3297,In_1105,In_1644);
or U3298 (N_3298,In_1129,In_429);
and U3299 (N_3299,In_2457,In_729);
xnor U3300 (N_3300,In_2725,In_1680);
nor U3301 (N_3301,In_1945,In_2301);
and U3302 (N_3302,In_945,In_1370);
and U3303 (N_3303,In_2229,In_2809);
and U3304 (N_3304,In_2936,In_96);
xnor U3305 (N_3305,In_1618,In_2365);
nand U3306 (N_3306,In_2449,In_609);
nor U3307 (N_3307,In_677,In_657);
xnor U3308 (N_3308,In_893,In_2445);
and U3309 (N_3309,In_2818,In_1444);
nor U3310 (N_3310,In_2169,In_2726);
nor U3311 (N_3311,In_1644,In_2649);
xor U3312 (N_3312,In_2863,In_41);
nand U3313 (N_3313,In_2321,In_1786);
nor U3314 (N_3314,In_1492,In_828);
or U3315 (N_3315,In_2242,In_2803);
nor U3316 (N_3316,In_1553,In_1220);
nand U3317 (N_3317,In_1280,In_523);
or U3318 (N_3318,In_520,In_962);
or U3319 (N_3319,In_257,In_2516);
nor U3320 (N_3320,In_932,In_1913);
nand U3321 (N_3321,In_49,In_713);
xor U3322 (N_3322,In_1789,In_2478);
nand U3323 (N_3323,In_1457,In_2805);
or U3324 (N_3324,In_295,In_1400);
and U3325 (N_3325,In_2982,In_2393);
and U3326 (N_3326,In_2574,In_1076);
and U3327 (N_3327,In_2887,In_1699);
or U3328 (N_3328,In_361,In_2703);
nand U3329 (N_3329,In_1347,In_658);
or U3330 (N_3330,In_644,In_2257);
xor U3331 (N_3331,In_140,In_2471);
xnor U3332 (N_3332,In_277,In_2117);
xnor U3333 (N_3333,In_1702,In_1755);
or U3334 (N_3334,In_2509,In_2798);
or U3335 (N_3335,In_219,In_978);
nor U3336 (N_3336,In_1100,In_2165);
or U3337 (N_3337,In_2891,In_1158);
xor U3338 (N_3338,In_1334,In_1167);
nand U3339 (N_3339,In_1630,In_2795);
and U3340 (N_3340,In_596,In_2818);
xor U3341 (N_3341,In_1591,In_2796);
or U3342 (N_3342,In_1005,In_1404);
and U3343 (N_3343,In_2946,In_1042);
nand U3344 (N_3344,In_1281,In_992);
or U3345 (N_3345,In_2067,In_2828);
nand U3346 (N_3346,In_2464,In_1057);
or U3347 (N_3347,In_619,In_1282);
and U3348 (N_3348,In_2492,In_1216);
nand U3349 (N_3349,In_1720,In_2817);
nand U3350 (N_3350,In_1533,In_2174);
and U3351 (N_3351,In_1539,In_2165);
or U3352 (N_3352,In_374,In_677);
xor U3353 (N_3353,In_1163,In_1525);
or U3354 (N_3354,In_2623,In_1367);
or U3355 (N_3355,In_2935,In_2013);
nor U3356 (N_3356,In_1013,In_1953);
or U3357 (N_3357,In_378,In_2639);
nor U3358 (N_3358,In_488,In_610);
nor U3359 (N_3359,In_1371,In_2435);
or U3360 (N_3360,In_2434,In_1105);
nor U3361 (N_3361,In_334,In_847);
nor U3362 (N_3362,In_2630,In_33);
and U3363 (N_3363,In_2908,In_175);
and U3364 (N_3364,In_2278,In_365);
nor U3365 (N_3365,In_724,In_356);
xor U3366 (N_3366,In_1846,In_2369);
nand U3367 (N_3367,In_448,In_1071);
and U3368 (N_3368,In_1872,In_2105);
xor U3369 (N_3369,In_1783,In_1662);
and U3370 (N_3370,In_39,In_614);
nand U3371 (N_3371,In_1170,In_569);
xnor U3372 (N_3372,In_1220,In_102);
nor U3373 (N_3373,In_2658,In_269);
nand U3374 (N_3374,In_1901,In_1838);
nor U3375 (N_3375,In_2108,In_2076);
nor U3376 (N_3376,In_1512,In_1616);
nor U3377 (N_3377,In_2779,In_1018);
and U3378 (N_3378,In_138,In_1623);
and U3379 (N_3379,In_1964,In_2076);
nor U3380 (N_3380,In_768,In_81);
and U3381 (N_3381,In_751,In_2046);
xnor U3382 (N_3382,In_662,In_1904);
and U3383 (N_3383,In_2872,In_2792);
and U3384 (N_3384,In_1963,In_2466);
nand U3385 (N_3385,In_1682,In_1482);
nor U3386 (N_3386,In_2277,In_1470);
and U3387 (N_3387,In_458,In_1849);
nand U3388 (N_3388,In_2333,In_1833);
nor U3389 (N_3389,In_2549,In_1170);
and U3390 (N_3390,In_2868,In_2685);
and U3391 (N_3391,In_852,In_1477);
or U3392 (N_3392,In_1013,In_1994);
xnor U3393 (N_3393,In_1947,In_1739);
nand U3394 (N_3394,In_319,In_1516);
or U3395 (N_3395,In_1175,In_365);
nor U3396 (N_3396,In_2303,In_2462);
nor U3397 (N_3397,In_317,In_2214);
or U3398 (N_3398,In_426,In_77);
or U3399 (N_3399,In_306,In_1599);
nand U3400 (N_3400,In_1416,In_2779);
nand U3401 (N_3401,In_1223,In_866);
or U3402 (N_3402,In_405,In_2221);
nand U3403 (N_3403,In_2545,In_2295);
xnor U3404 (N_3404,In_2176,In_482);
or U3405 (N_3405,In_1555,In_425);
xnor U3406 (N_3406,In_2380,In_1921);
or U3407 (N_3407,In_321,In_108);
or U3408 (N_3408,In_2475,In_2269);
nor U3409 (N_3409,In_988,In_1151);
xor U3410 (N_3410,In_2090,In_2050);
and U3411 (N_3411,In_1958,In_1831);
nor U3412 (N_3412,In_1734,In_1441);
or U3413 (N_3413,In_753,In_1283);
or U3414 (N_3414,In_2939,In_795);
or U3415 (N_3415,In_1958,In_1033);
nand U3416 (N_3416,In_292,In_2783);
and U3417 (N_3417,In_1304,In_2159);
xor U3418 (N_3418,In_1977,In_1976);
xnor U3419 (N_3419,In_2414,In_2024);
nand U3420 (N_3420,In_2178,In_983);
or U3421 (N_3421,In_154,In_465);
and U3422 (N_3422,In_1624,In_2777);
xnor U3423 (N_3423,In_2066,In_2985);
xnor U3424 (N_3424,In_1031,In_1785);
and U3425 (N_3425,In_122,In_1344);
or U3426 (N_3426,In_480,In_251);
nand U3427 (N_3427,In_560,In_2450);
xor U3428 (N_3428,In_1530,In_2833);
xor U3429 (N_3429,In_1403,In_529);
or U3430 (N_3430,In_1568,In_1947);
or U3431 (N_3431,In_384,In_1950);
nor U3432 (N_3432,In_210,In_220);
xnor U3433 (N_3433,In_1209,In_1811);
or U3434 (N_3434,In_1238,In_2590);
nor U3435 (N_3435,In_2492,In_1808);
nand U3436 (N_3436,In_2094,In_256);
or U3437 (N_3437,In_2970,In_2376);
or U3438 (N_3438,In_762,In_1952);
nand U3439 (N_3439,In_2600,In_2835);
nand U3440 (N_3440,In_458,In_270);
nand U3441 (N_3441,In_686,In_2544);
or U3442 (N_3442,In_1939,In_254);
and U3443 (N_3443,In_2155,In_82);
xnor U3444 (N_3444,In_686,In_217);
and U3445 (N_3445,In_2898,In_1695);
nand U3446 (N_3446,In_1226,In_2921);
nor U3447 (N_3447,In_2889,In_1172);
nand U3448 (N_3448,In_648,In_625);
nand U3449 (N_3449,In_238,In_130);
nand U3450 (N_3450,In_2169,In_1907);
xor U3451 (N_3451,In_2730,In_2555);
and U3452 (N_3452,In_489,In_2496);
nor U3453 (N_3453,In_756,In_1673);
and U3454 (N_3454,In_1879,In_2397);
xor U3455 (N_3455,In_1134,In_883);
nor U3456 (N_3456,In_535,In_2671);
nor U3457 (N_3457,In_1688,In_2326);
nor U3458 (N_3458,In_1831,In_975);
nand U3459 (N_3459,In_1703,In_924);
and U3460 (N_3460,In_2073,In_2126);
and U3461 (N_3461,In_702,In_1081);
xor U3462 (N_3462,In_2465,In_553);
and U3463 (N_3463,In_164,In_2205);
xor U3464 (N_3464,In_595,In_1747);
xor U3465 (N_3465,In_2351,In_523);
nand U3466 (N_3466,In_124,In_2152);
nor U3467 (N_3467,In_2371,In_128);
or U3468 (N_3468,In_1662,In_2187);
xor U3469 (N_3469,In_2875,In_2989);
nor U3470 (N_3470,In_565,In_2318);
nand U3471 (N_3471,In_841,In_1270);
nor U3472 (N_3472,In_2092,In_2296);
nand U3473 (N_3473,In_1862,In_839);
or U3474 (N_3474,In_684,In_2787);
xor U3475 (N_3475,In_1564,In_1056);
and U3476 (N_3476,In_1611,In_1269);
nand U3477 (N_3477,In_284,In_1512);
nor U3478 (N_3478,In_1630,In_563);
nor U3479 (N_3479,In_241,In_497);
xnor U3480 (N_3480,In_1576,In_2619);
or U3481 (N_3481,In_2226,In_359);
nand U3482 (N_3482,In_1997,In_1519);
or U3483 (N_3483,In_1196,In_2256);
nor U3484 (N_3484,In_92,In_123);
nor U3485 (N_3485,In_1403,In_1207);
and U3486 (N_3486,In_85,In_1533);
xnor U3487 (N_3487,In_348,In_2103);
xnor U3488 (N_3488,In_2294,In_1644);
nor U3489 (N_3489,In_770,In_254);
or U3490 (N_3490,In_940,In_2722);
or U3491 (N_3491,In_237,In_2947);
nand U3492 (N_3492,In_646,In_1890);
nand U3493 (N_3493,In_1822,In_2694);
and U3494 (N_3494,In_715,In_1937);
or U3495 (N_3495,In_562,In_797);
nand U3496 (N_3496,In_2979,In_2419);
nand U3497 (N_3497,In_1110,In_851);
nor U3498 (N_3498,In_1587,In_2158);
nor U3499 (N_3499,In_533,In_2327);
and U3500 (N_3500,In_2658,In_790);
nand U3501 (N_3501,In_2908,In_901);
nor U3502 (N_3502,In_2891,In_763);
xor U3503 (N_3503,In_1033,In_616);
xor U3504 (N_3504,In_570,In_1443);
nor U3505 (N_3505,In_478,In_52);
nor U3506 (N_3506,In_941,In_2587);
or U3507 (N_3507,In_347,In_1476);
nor U3508 (N_3508,In_2192,In_909);
or U3509 (N_3509,In_1912,In_594);
or U3510 (N_3510,In_996,In_75);
nand U3511 (N_3511,In_1027,In_462);
xor U3512 (N_3512,In_1207,In_2275);
xnor U3513 (N_3513,In_118,In_263);
nand U3514 (N_3514,In_2169,In_1040);
nand U3515 (N_3515,In_318,In_63);
and U3516 (N_3516,In_2662,In_391);
nand U3517 (N_3517,In_1449,In_2382);
nand U3518 (N_3518,In_2305,In_740);
and U3519 (N_3519,In_2606,In_2987);
nand U3520 (N_3520,In_459,In_453);
xor U3521 (N_3521,In_638,In_486);
nand U3522 (N_3522,In_2555,In_2142);
or U3523 (N_3523,In_599,In_289);
nand U3524 (N_3524,In_957,In_668);
and U3525 (N_3525,In_2155,In_162);
xnor U3526 (N_3526,In_2359,In_2703);
and U3527 (N_3527,In_2576,In_2394);
nor U3528 (N_3528,In_2563,In_2238);
nand U3529 (N_3529,In_1917,In_2393);
and U3530 (N_3530,In_2173,In_485);
and U3531 (N_3531,In_2927,In_1611);
nor U3532 (N_3532,In_2000,In_821);
nor U3533 (N_3533,In_1247,In_1253);
and U3534 (N_3534,In_154,In_1183);
or U3535 (N_3535,In_2198,In_372);
xor U3536 (N_3536,In_1962,In_357);
or U3537 (N_3537,In_1952,In_2677);
xor U3538 (N_3538,In_319,In_1432);
or U3539 (N_3539,In_570,In_1537);
nand U3540 (N_3540,In_1878,In_2015);
nor U3541 (N_3541,In_412,In_2217);
nor U3542 (N_3542,In_2836,In_2662);
and U3543 (N_3543,In_131,In_1000);
and U3544 (N_3544,In_1412,In_1808);
or U3545 (N_3545,In_1991,In_2502);
and U3546 (N_3546,In_371,In_444);
or U3547 (N_3547,In_1433,In_2826);
or U3548 (N_3548,In_2214,In_498);
nand U3549 (N_3549,In_2094,In_2767);
nor U3550 (N_3550,In_67,In_2866);
nor U3551 (N_3551,In_2947,In_319);
or U3552 (N_3552,In_1458,In_2268);
nor U3553 (N_3553,In_395,In_1141);
or U3554 (N_3554,In_2839,In_2824);
xnor U3555 (N_3555,In_2584,In_764);
or U3556 (N_3556,In_2371,In_362);
or U3557 (N_3557,In_2742,In_1556);
and U3558 (N_3558,In_2747,In_80);
nor U3559 (N_3559,In_1174,In_1590);
or U3560 (N_3560,In_1274,In_1693);
xor U3561 (N_3561,In_1803,In_972);
or U3562 (N_3562,In_1521,In_800);
and U3563 (N_3563,In_2493,In_2745);
and U3564 (N_3564,In_1947,In_2894);
or U3565 (N_3565,In_1134,In_1226);
or U3566 (N_3566,In_1861,In_2833);
xnor U3567 (N_3567,In_2790,In_1942);
nand U3568 (N_3568,In_462,In_2036);
nor U3569 (N_3569,In_1650,In_1374);
xnor U3570 (N_3570,In_159,In_1332);
xnor U3571 (N_3571,In_223,In_1793);
and U3572 (N_3572,In_2384,In_2650);
xnor U3573 (N_3573,In_2973,In_2682);
xor U3574 (N_3574,In_273,In_2156);
nor U3575 (N_3575,In_1639,In_2004);
xnor U3576 (N_3576,In_1092,In_1996);
nor U3577 (N_3577,In_18,In_2076);
and U3578 (N_3578,In_1876,In_2883);
nand U3579 (N_3579,In_1572,In_402);
xor U3580 (N_3580,In_1492,In_636);
xor U3581 (N_3581,In_125,In_623);
nor U3582 (N_3582,In_2294,In_2163);
or U3583 (N_3583,In_1262,In_1742);
and U3584 (N_3584,In_2226,In_1801);
or U3585 (N_3585,In_149,In_2165);
nor U3586 (N_3586,In_2694,In_2391);
and U3587 (N_3587,In_435,In_2146);
nand U3588 (N_3588,In_1353,In_2963);
and U3589 (N_3589,In_490,In_613);
nand U3590 (N_3590,In_1925,In_1849);
and U3591 (N_3591,In_1769,In_2380);
nand U3592 (N_3592,In_2600,In_2065);
and U3593 (N_3593,In_1285,In_1898);
nand U3594 (N_3594,In_208,In_1844);
or U3595 (N_3595,In_2819,In_2614);
xnor U3596 (N_3596,In_1007,In_1806);
nor U3597 (N_3597,In_2608,In_261);
or U3598 (N_3598,In_65,In_103);
or U3599 (N_3599,In_1186,In_2922);
xor U3600 (N_3600,In_1517,In_1961);
xor U3601 (N_3601,In_1473,In_2102);
nor U3602 (N_3602,In_2683,In_1487);
xnor U3603 (N_3603,In_99,In_2056);
xor U3604 (N_3604,In_2577,In_672);
nand U3605 (N_3605,In_1414,In_315);
nor U3606 (N_3606,In_2825,In_1713);
nand U3607 (N_3607,In_2057,In_1590);
or U3608 (N_3608,In_514,In_991);
nor U3609 (N_3609,In_1505,In_808);
and U3610 (N_3610,In_2831,In_1875);
nor U3611 (N_3611,In_382,In_1352);
and U3612 (N_3612,In_2281,In_1118);
or U3613 (N_3613,In_159,In_409);
xnor U3614 (N_3614,In_1031,In_2405);
and U3615 (N_3615,In_2591,In_1349);
or U3616 (N_3616,In_223,In_686);
nor U3617 (N_3617,In_1936,In_482);
or U3618 (N_3618,In_2733,In_320);
nand U3619 (N_3619,In_1078,In_1781);
xnor U3620 (N_3620,In_2155,In_2769);
or U3621 (N_3621,In_2888,In_759);
nor U3622 (N_3622,In_394,In_102);
xnor U3623 (N_3623,In_1717,In_13);
and U3624 (N_3624,In_1576,In_1229);
nor U3625 (N_3625,In_2714,In_2916);
or U3626 (N_3626,In_2923,In_2150);
nor U3627 (N_3627,In_2854,In_2812);
nor U3628 (N_3628,In_7,In_1701);
and U3629 (N_3629,In_2124,In_2516);
or U3630 (N_3630,In_758,In_2657);
xor U3631 (N_3631,In_2269,In_2725);
xor U3632 (N_3632,In_929,In_619);
nor U3633 (N_3633,In_1289,In_2149);
xor U3634 (N_3634,In_1133,In_635);
nor U3635 (N_3635,In_513,In_1477);
or U3636 (N_3636,In_1346,In_2707);
or U3637 (N_3637,In_111,In_1430);
and U3638 (N_3638,In_23,In_980);
nand U3639 (N_3639,In_2601,In_2487);
and U3640 (N_3640,In_1151,In_1072);
nand U3641 (N_3641,In_2592,In_966);
xnor U3642 (N_3642,In_418,In_493);
xnor U3643 (N_3643,In_760,In_1654);
nand U3644 (N_3644,In_179,In_2850);
nor U3645 (N_3645,In_702,In_689);
nand U3646 (N_3646,In_1469,In_1665);
nor U3647 (N_3647,In_2940,In_1934);
nor U3648 (N_3648,In_2666,In_2213);
nor U3649 (N_3649,In_1603,In_1035);
and U3650 (N_3650,In_1646,In_1015);
nand U3651 (N_3651,In_861,In_282);
nand U3652 (N_3652,In_2104,In_2240);
nand U3653 (N_3653,In_515,In_1177);
xnor U3654 (N_3654,In_2221,In_228);
and U3655 (N_3655,In_1601,In_1235);
or U3656 (N_3656,In_533,In_2236);
nor U3657 (N_3657,In_20,In_2605);
nand U3658 (N_3658,In_1396,In_2014);
xor U3659 (N_3659,In_2273,In_2741);
xnor U3660 (N_3660,In_1601,In_1647);
nand U3661 (N_3661,In_343,In_2707);
nor U3662 (N_3662,In_2124,In_2714);
or U3663 (N_3663,In_481,In_1921);
and U3664 (N_3664,In_2157,In_2640);
or U3665 (N_3665,In_2368,In_1294);
nor U3666 (N_3666,In_2110,In_1567);
nor U3667 (N_3667,In_731,In_2805);
xnor U3668 (N_3668,In_2876,In_116);
nor U3669 (N_3669,In_647,In_2276);
nor U3670 (N_3670,In_1581,In_1450);
xor U3671 (N_3671,In_2422,In_1352);
or U3672 (N_3672,In_592,In_82);
nor U3673 (N_3673,In_1400,In_221);
and U3674 (N_3674,In_2637,In_77);
and U3675 (N_3675,In_1528,In_2762);
nand U3676 (N_3676,In_1674,In_122);
nor U3677 (N_3677,In_1462,In_2344);
or U3678 (N_3678,In_1905,In_1807);
or U3679 (N_3679,In_794,In_314);
nand U3680 (N_3680,In_2833,In_658);
xor U3681 (N_3681,In_584,In_42);
xor U3682 (N_3682,In_1704,In_2804);
nand U3683 (N_3683,In_2428,In_987);
and U3684 (N_3684,In_2628,In_2264);
nand U3685 (N_3685,In_1939,In_1049);
and U3686 (N_3686,In_2507,In_1695);
or U3687 (N_3687,In_360,In_1931);
xnor U3688 (N_3688,In_907,In_1844);
and U3689 (N_3689,In_941,In_1962);
and U3690 (N_3690,In_1401,In_1665);
and U3691 (N_3691,In_2404,In_1956);
xor U3692 (N_3692,In_1963,In_1636);
and U3693 (N_3693,In_2030,In_849);
xnor U3694 (N_3694,In_473,In_167);
nor U3695 (N_3695,In_2224,In_677);
nand U3696 (N_3696,In_1833,In_1904);
xor U3697 (N_3697,In_682,In_240);
and U3698 (N_3698,In_2116,In_349);
or U3699 (N_3699,In_1970,In_2722);
and U3700 (N_3700,In_427,In_2838);
nor U3701 (N_3701,In_1133,In_302);
or U3702 (N_3702,In_1329,In_446);
and U3703 (N_3703,In_2334,In_2153);
nor U3704 (N_3704,In_1863,In_1855);
nor U3705 (N_3705,In_2769,In_1665);
or U3706 (N_3706,In_1414,In_323);
xor U3707 (N_3707,In_911,In_1524);
nand U3708 (N_3708,In_1839,In_956);
and U3709 (N_3709,In_1833,In_2547);
or U3710 (N_3710,In_1578,In_2528);
or U3711 (N_3711,In_2613,In_1047);
and U3712 (N_3712,In_246,In_145);
xnor U3713 (N_3713,In_2,In_2667);
nor U3714 (N_3714,In_2256,In_1462);
nor U3715 (N_3715,In_1981,In_1156);
nand U3716 (N_3716,In_585,In_179);
nand U3717 (N_3717,In_2940,In_2299);
and U3718 (N_3718,In_3,In_2455);
xor U3719 (N_3719,In_335,In_2811);
and U3720 (N_3720,In_439,In_2516);
nor U3721 (N_3721,In_1392,In_632);
and U3722 (N_3722,In_637,In_2996);
nand U3723 (N_3723,In_566,In_1552);
and U3724 (N_3724,In_2459,In_963);
and U3725 (N_3725,In_895,In_344);
xor U3726 (N_3726,In_632,In_2226);
and U3727 (N_3727,In_2585,In_2353);
or U3728 (N_3728,In_1915,In_1185);
or U3729 (N_3729,In_1408,In_362);
or U3730 (N_3730,In_1201,In_323);
and U3731 (N_3731,In_561,In_1980);
and U3732 (N_3732,In_2760,In_1623);
nor U3733 (N_3733,In_1145,In_616);
nor U3734 (N_3734,In_932,In_2171);
nor U3735 (N_3735,In_707,In_100);
or U3736 (N_3736,In_806,In_2777);
nor U3737 (N_3737,In_1081,In_1293);
and U3738 (N_3738,In_1930,In_2440);
and U3739 (N_3739,In_363,In_2080);
xor U3740 (N_3740,In_1908,In_767);
xnor U3741 (N_3741,In_574,In_587);
and U3742 (N_3742,In_764,In_462);
nand U3743 (N_3743,In_576,In_1556);
or U3744 (N_3744,In_1832,In_2445);
and U3745 (N_3745,In_517,In_409);
xnor U3746 (N_3746,In_2778,In_1580);
nand U3747 (N_3747,In_1786,In_248);
nand U3748 (N_3748,In_2868,In_2604);
or U3749 (N_3749,In_104,In_1989);
nand U3750 (N_3750,In_2201,In_835);
and U3751 (N_3751,In_1340,In_2566);
or U3752 (N_3752,In_1045,In_906);
nand U3753 (N_3753,In_2425,In_2711);
or U3754 (N_3754,In_2028,In_2024);
nor U3755 (N_3755,In_1211,In_2281);
nand U3756 (N_3756,In_1318,In_751);
xor U3757 (N_3757,In_1239,In_953);
nor U3758 (N_3758,In_2418,In_2655);
nor U3759 (N_3759,In_2828,In_671);
or U3760 (N_3760,In_1076,In_810);
and U3761 (N_3761,In_2581,In_1509);
xor U3762 (N_3762,In_2914,In_2151);
or U3763 (N_3763,In_972,In_1554);
nor U3764 (N_3764,In_1420,In_1986);
xnor U3765 (N_3765,In_1123,In_2534);
nand U3766 (N_3766,In_2184,In_2636);
or U3767 (N_3767,In_144,In_2675);
or U3768 (N_3768,In_1908,In_2796);
and U3769 (N_3769,In_2301,In_2642);
nand U3770 (N_3770,In_679,In_243);
nand U3771 (N_3771,In_2021,In_1666);
or U3772 (N_3772,In_1747,In_2660);
nor U3773 (N_3773,In_1755,In_2586);
nor U3774 (N_3774,In_1079,In_1132);
or U3775 (N_3775,In_319,In_2897);
xor U3776 (N_3776,In_2965,In_2554);
and U3777 (N_3777,In_1378,In_445);
xor U3778 (N_3778,In_938,In_1767);
and U3779 (N_3779,In_2584,In_1316);
xor U3780 (N_3780,In_963,In_2894);
nor U3781 (N_3781,In_2049,In_677);
and U3782 (N_3782,In_1926,In_1091);
nor U3783 (N_3783,In_2758,In_1691);
xor U3784 (N_3784,In_1087,In_743);
nand U3785 (N_3785,In_1555,In_2762);
or U3786 (N_3786,In_980,In_1384);
nor U3787 (N_3787,In_2422,In_219);
nor U3788 (N_3788,In_184,In_2332);
and U3789 (N_3789,In_256,In_2828);
and U3790 (N_3790,In_1507,In_2721);
or U3791 (N_3791,In_1029,In_474);
or U3792 (N_3792,In_921,In_2007);
xor U3793 (N_3793,In_1653,In_2636);
and U3794 (N_3794,In_1774,In_2803);
nand U3795 (N_3795,In_1346,In_511);
and U3796 (N_3796,In_2445,In_1638);
nor U3797 (N_3797,In_2077,In_1755);
or U3798 (N_3798,In_994,In_505);
nand U3799 (N_3799,In_1909,In_2494);
nor U3800 (N_3800,In_801,In_574);
nor U3801 (N_3801,In_2031,In_1521);
or U3802 (N_3802,In_1530,In_2367);
and U3803 (N_3803,In_246,In_2026);
xor U3804 (N_3804,In_927,In_1421);
nor U3805 (N_3805,In_796,In_2450);
nand U3806 (N_3806,In_1605,In_324);
and U3807 (N_3807,In_2113,In_861);
nor U3808 (N_3808,In_465,In_129);
or U3809 (N_3809,In_2244,In_916);
and U3810 (N_3810,In_1921,In_1646);
or U3811 (N_3811,In_1797,In_1295);
or U3812 (N_3812,In_946,In_2336);
and U3813 (N_3813,In_222,In_1355);
nor U3814 (N_3814,In_2417,In_1149);
and U3815 (N_3815,In_2038,In_2299);
or U3816 (N_3816,In_1174,In_556);
and U3817 (N_3817,In_176,In_1307);
or U3818 (N_3818,In_1121,In_470);
xor U3819 (N_3819,In_2207,In_499);
and U3820 (N_3820,In_2420,In_2815);
nand U3821 (N_3821,In_381,In_1208);
nand U3822 (N_3822,In_918,In_2496);
and U3823 (N_3823,In_1359,In_86);
nor U3824 (N_3824,In_922,In_752);
or U3825 (N_3825,In_1192,In_357);
xnor U3826 (N_3826,In_1667,In_1151);
xor U3827 (N_3827,In_651,In_2519);
and U3828 (N_3828,In_2755,In_1123);
or U3829 (N_3829,In_1707,In_371);
and U3830 (N_3830,In_52,In_2152);
xnor U3831 (N_3831,In_593,In_1315);
nand U3832 (N_3832,In_1896,In_360);
and U3833 (N_3833,In_266,In_2736);
nand U3834 (N_3834,In_2922,In_507);
nor U3835 (N_3835,In_871,In_868);
and U3836 (N_3836,In_1521,In_482);
and U3837 (N_3837,In_1050,In_703);
or U3838 (N_3838,In_897,In_2795);
nand U3839 (N_3839,In_2851,In_1557);
nor U3840 (N_3840,In_1960,In_723);
nand U3841 (N_3841,In_1144,In_886);
and U3842 (N_3842,In_450,In_1241);
xnor U3843 (N_3843,In_2661,In_2442);
nand U3844 (N_3844,In_631,In_2323);
or U3845 (N_3845,In_1912,In_1211);
or U3846 (N_3846,In_2250,In_2500);
nor U3847 (N_3847,In_2602,In_2459);
nand U3848 (N_3848,In_918,In_2708);
xnor U3849 (N_3849,In_1190,In_1900);
or U3850 (N_3850,In_2011,In_2316);
nor U3851 (N_3851,In_290,In_1599);
or U3852 (N_3852,In_1419,In_2504);
nor U3853 (N_3853,In_1070,In_200);
and U3854 (N_3854,In_116,In_106);
nor U3855 (N_3855,In_2770,In_906);
nand U3856 (N_3856,In_1507,In_2781);
xor U3857 (N_3857,In_1871,In_1734);
xnor U3858 (N_3858,In_500,In_2927);
nor U3859 (N_3859,In_2462,In_1659);
nor U3860 (N_3860,In_966,In_2728);
xor U3861 (N_3861,In_363,In_2585);
nor U3862 (N_3862,In_2034,In_2152);
or U3863 (N_3863,In_991,In_2200);
nor U3864 (N_3864,In_914,In_1915);
nand U3865 (N_3865,In_200,In_1869);
nand U3866 (N_3866,In_2876,In_1025);
nor U3867 (N_3867,In_2148,In_170);
nor U3868 (N_3868,In_101,In_243);
and U3869 (N_3869,In_669,In_2811);
and U3870 (N_3870,In_824,In_361);
or U3871 (N_3871,In_1512,In_2456);
and U3872 (N_3872,In_1979,In_1339);
or U3873 (N_3873,In_1762,In_167);
nand U3874 (N_3874,In_1806,In_546);
xor U3875 (N_3875,In_1007,In_1608);
nor U3876 (N_3876,In_375,In_1144);
nor U3877 (N_3877,In_2560,In_377);
xor U3878 (N_3878,In_420,In_2995);
nor U3879 (N_3879,In_325,In_1404);
or U3880 (N_3880,In_2555,In_264);
and U3881 (N_3881,In_1467,In_150);
and U3882 (N_3882,In_1563,In_1352);
nor U3883 (N_3883,In_2248,In_2955);
nor U3884 (N_3884,In_855,In_2345);
xor U3885 (N_3885,In_2195,In_2513);
and U3886 (N_3886,In_1889,In_1942);
and U3887 (N_3887,In_2621,In_194);
xnor U3888 (N_3888,In_1355,In_1321);
nand U3889 (N_3889,In_1872,In_1727);
and U3890 (N_3890,In_1613,In_134);
nand U3891 (N_3891,In_839,In_2041);
or U3892 (N_3892,In_1155,In_1655);
xor U3893 (N_3893,In_1835,In_1482);
nand U3894 (N_3894,In_2236,In_1155);
nand U3895 (N_3895,In_1444,In_625);
nor U3896 (N_3896,In_2911,In_2960);
and U3897 (N_3897,In_2679,In_2870);
xnor U3898 (N_3898,In_161,In_2398);
nor U3899 (N_3899,In_2711,In_588);
xor U3900 (N_3900,In_556,In_2236);
or U3901 (N_3901,In_232,In_716);
or U3902 (N_3902,In_2702,In_1877);
and U3903 (N_3903,In_1610,In_2176);
nand U3904 (N_3904,In_128,In_2804);
nand U3905 (N_3905,In_2950,In_198);
xnor U3906 (N_3906,In_313,In_645);
or U3907 (N_3907,In_853,In_2189);
nand U3908 (N_3908,In_1974,In_1158);
xor U3909 (N_3909,In_2614,In_2764);
xnor U3910 (N_3910,In_1181,In_2111);
or U3911 (N_3911,In_2149,In_1748);
or U3912 (N_3912,In_2381,In_1778);
or U3913 (N_3913,In_1721,In_1851);
nand U3914 (N_3914,In_2413,In_1859);
and U3915 (N_3915,In_1047,In_1623);
xor U3916 (N_3916,In_1830,In_815);
and U3917 (N_3917,In_1205,In_531);
xor U3918 (N_3918,In_1419,In_683);
or U3919 (N_3919,In_1131,In_2092);
xor U3920 (N_3920,In_2955,In_958);
and U3921 (N_3921,In_1923,In_1685);
nor U3922 (N_3922,In_2379,In_328);
and U3923 (N_3923,In_521,In_1824);
nor U3924 (N_3924,In_1405,In_1111);
or U3925 (N_3925,In_253,In_1688);
nand U3926 (N_3926,In_1271,In_1837);
nor U3927 (N_3927,In_2615,In_368);
xnor U3928 (N_3928,In_606,In_2205);
nor U3929 (N_3929,In_1203,In_786);
nand U3930 (N_3930,In_207,In_89);
nor U3931 (N_3931,In_1482,In_2374);
nand U3932 (N_3932,In_2446,In_715);
xnor U3933 (N_3933,In_2393,In_1993);
nand U3934 (N_3934,In_840,In_1963);
or U3935 (N_3935,In_2682,In_273);
and U3936 (N_3936,In_1094,In_2014);
nand U3937 (N_3937,In_150,In_1100);
nand U3938 (N_3938,In_692,In_262);
or U3939 (N_3939,In_551,In_369);
nand U3940 (N_3940,In_271,In_985);
and U3941 (N_3941,In_1404,In_549);
and U3942 (N_3942,In_2047,In_1803);
nand U3943 (N_3943,In_1021,In_1035);
nand U3944 (N_3944,In_1281,In_36);
and U3945 (N_3945,In_1437,In_122);
xnor U3946 (N_3946,In_1520,In_2819);
and U3947 (N_3947,In_1827,In_637);
or U3948 (N_3948,In_1830,In_2643);
xnor U3949 (N_3949,In_1820,In_597);
nand U3950 (N_3950,In_2602,In_1482);
nand U3951 (N_3951,In_144,In_550);
and U3952 (N_3952,In_1527,In_826);
xnor U3953 (N_3953,In_2845,In_1027);
nor U3954 (N_3954,In_1242,In_263);
nand U3955 (N_3955,In_2459,In_765);
or U3956 (N_3956,In_1565,In_2339);
and U3957 (N_3957,In_94,In_2136);
nor U3958 (N_3958,In_1926,In_11);
or U3959 (N_3959,In_696,In_3);
or U3960 (N_3960,In_2506,In_1242);
nor U3961 (N_3961,In_2629,In_969);
or U3962 (N_3962,In_1230,In_1565);
xnor U3963 (N_3963,In_418,In_513);
xor U3964 (N_3964,In_2737,In_1452);
or U3965 (N_3965,In_2458,In_1238);
or U3966 (N_3966,In_2120,In_1298);
nor U3967 (N_3967,In_1980,In_1164);
or U3968 (N_3968,In_505,In_2993);
and U3969 (N_3969,In_2861,In_2267);
and U3970 (N_3970,In_1388,In_912);
or U3971 (N_3971,In_896,In_1850);
nor U3972 (N_3972,In_1414,In_2129);
and U3973 (N_3973,In_2397,In_1550);
nor U3974 (N_3974,In_346,In_1563);
and U3975 (N_3975,In_696,In_2774);
xnor U3976 (N_3976,In_2349,In_357);
xor U3977 (N_3977,In_2437,In_499);
or U3978 (N_3978,In_2856,In_118);
nor U3979 (N_3979,In_2514,In_2631);
or U3980 (N_3980,In_2562,In_1254);
or U3981 (N_3981,In_679,In_2104);
or U3982 (N_3982,In_1868,In_208);
and U3983 (N_3983,In_1079,In_142);
and U3984 (N_3984,In_478,In_1297);
xnor U3985 (N_3985,In_1304,In_2862);
nor U3986 (N_3986,In_1935,In_597);
xor U3987 (N_3987,In_916,In_2179);
nand U3988 (N_3988,In_1486,In_2721);
xor U3989 (N_3989,In_2992,In_2040);
nor U3990 (N_3990,In_677,In_1887);
and U3991 (N_3991,In_2106,In_760);
and U3992 (N_3992,In_2984,In_195);
xnor U3993 (N_3993,In_1174,In_1961);
or U3994 (N_3994,In_1132,In_2688);
nand U3995 (N_3995,In_2779,In_1847);
and U3996 (N_3996,In_1975,In_2287);
or U3997 (N_3997,In_1079,In_1236);
xnor U3998 (N_3998,In_634,In_924);
xor U3999 (N_3999,In_1510,In_929);
nor U4000 (N_4000,In_2602,In_2319);
nor U4001 (N_4001,In_535,In_2806);
or U4002 (N_4002,In_2994,In_1385);
nor U4003 (N_4003,In_1534,In_568);
xor U4004 (N_4004,In_1520,In_1549);
and U4005 (N_4005,In_117,In_39);
nand U4006 (N_4006,In_1297,In_2469);
nor U4007 (N_4007,In_1895,In_1109);
and U4008 (N_4008,In_2596,In_2128);
and U4009 (N_4009,In_498,In_100);
and U4010 (N_4010,In_94,In_1763);
and U4011 (N_4011,In_463,In_2857);
nand U4012 (N_4012,In_680,In_128);
and U4013 (N_4013,In_1772,In_1734);
nor U4014 (N_4014,In_781,In_1555);
xor U4015 (N_4015,In_2292,In_881);
nand U4016 (N_4016,In_2969,In_2072);
nor U4017 (N_4017,In_1167,In_2201);
or U4018 (N_4018,In_579,In_2200);
xor U4019 (N_4019,In_96,In_1567);
nor U4020 (N_4020,In_1542,In_2508);
nand U4021 (N_4021,In_648,In_962);
and U4022 (N_4022,In_352,In_83);
and U4023 (N_4023,In_273,In_1505);
and U4024 (N_4024,In_841,In_2841);
or U4025 (N_4025,In_2154,In_212);
nor U4026 (N_4026,In_1165,In_2920);
nor U4027 (N_4027,In_2149,In_310);
and U4028 (N_4028,In_1905,In_842);
nand U4029 (N_4029,In_2241,In_1833);
or U4030 (N_4030,In_1883,In_2842);
or U4031 (N_4031,In_475,In_177);
or U4032 (N_4032,In_1455,In_1835);
or U4033 (N_4033,In_2958,In_332);
nor U4034 (N_4034,In_2980,In_1318);
nor U4035 (N_4035,In_1709,In_1930);
or U4036 (N_4036,In_1226,In_2845);
or U4037 (N_4037,In_2922,In_823);
xor U4038 (N_4038,In_522,In_2951);
xor U4039 (N_4039,In_918,In_2352);
nand U4040 (N_4040,In_2277,In_1558);
nor U4041 (N_4041,In_1838,In_672);
or U4042 (N_4042,In_2664,In_1904);
nor U4043 (N_4043,In_425,In_2289);
nand U4044 (N_4044,In_1858,In_2325);
nor U4045 (N_4045,In_50,In_1395);
or U4046 (N_4046,In_2227,In_1684);
xor U4047 (N_4047,In_2430,In_200);
xor U4048 (N_4048,In_1879,In_2925);
and U4049 (N_4049,In_2174,In_2087);
nor U4050 (N_4050,In_129,In_2816);
and U4051 (N_4051,In_88,In_198);
or U4052 (N_4052,In_1321,In_1822);
nor U4053 (N_4053,In_2607,In_929);
nand U4054 (N_4054,In_2481,In_1966);
nor U4055 (N_4055,In_1762,In_2550);
or U4056 (N_4056,In_273,In_2644);
nand U4057 (N_4057,In_928,In_124);
nor U4058 (N_4058,In_2528,In_2641);
nand U4059 (N_4059,In_2154,In_2348);
or U4060 (N_4060,In_2133,In_738);
and U4061 (N_4061,In_461,In_1613);
nor U4062 (N_4062,In_1287,In_2080);
nor U4063 (N_4063,In_2941,In_559);
nor U4064 (N_4064,In_1980,In_599);
nor U4065 (N_4065,In_204,In_2267);
nand U4066 (N_4066,In_2882,In_691);
nor U4067 (N_4067,In_2839,In_2428);
nor U4068 (N_4068,In_1591,In_238);
or U4069 (N_4069,In_460,In_461);
and U4070 (N_4070,In_1203,In_848);
xor U4071 (N_4071,In_692,In_690);
nand U4072 (N_4072,In_1010,In_252);
xnor U4073 (N_4073,In_2078,In_1230);
and U4074 (N_4074,In_1687,In_495);
nand U4075 (N_4075,In_637,In_461);
or U4076 (N_4076,In_1258,In_1983);
and U4077 (N_4077,In_2011,In_173);
nand U4078 (N_4078,In_758,In_2514);
nand U4079 (N_4079,In_2586,In_501);
or U4080 (N_4080,In_1042,In_2948);
xnor U4081 (N_4081,In_1610,In_706);
nand U4082 (N_4082,In_936,In_990);
nor U4083 (N_4083,In_2042,In_2652);
nand U4084 (N_4084,In_2458,In_2855);
nand U4085 (N_4085,In_1323,In_1463);
nor U4086 (N_4086,In_1829,In_1386);
nand U4087 (N_4087,In_1650,In_1704);
xnor U4088 (N_4088,In_1170,In_2495);
nor U4089 (N_4089,In_1434,In_1765);
or U4090 (N_4090,In_1791,In_1612);
or U4091 (N_4091,In_368,In_117);
xnor U4092 (N_4092,In_1020,In_1078);
nand U4093 (N_4093,In_1874,In_1618);
nand U4094 (N_4094,In_283,In_1459);
nor U4095 (N_4095,In_2231,In_2040);
or U4096 (N_4096,In_2500,In_1456);
xnor U4097 (N_4097,In_198,In_1885);
nor U4098 (N_4098,In_1895,In_2515);
nand U4099 (N_4099,In_451,In_1317);
nand U4100 (N_4100,In_45,In_1013);
xor U4101 (N_4101,In_1779,In_2742);
xnor U4102 (N_4102,In_242,In_2596);
nand U4103 (N_4103,In_955,In_772);
nand U4104 (N_4104,In_2481,In_1207);
and U4105 (N_4105,In_2685,In_423);
and U4106 (N_4106,In_2224,In_2270);
or U4107 (N_4107,In_535,In_2247);
and U4108 (N_4108,In_2599,In_1507);
nor U4109 (N_4109,In_784,In_2444);
or U4110 (N_4110,In_151,In_2555);
xor U4111 (N_4111,In_1667,In_1535);
nand U4112 (N_4112,In_63,In_1183);
xnor U4113 (N_4113,In_20,In_266);
and U4114 (N_4114,In_2684,In_2099);
nand U4115 (N_4115,In_629,In_670);
nor U4116 (N_4116,In_1730,In_114);
nand U4117 (N_4117,In_1746,In_710);
and U4118 (N_4118,In_2313,In_2904);
and U4119 (N_4119,In_1273,In_1447);
xnor U4120 (N_4120,In_2985,In_217);
nand U4121 (N_4121,In_196,In_2250);
and U4122 (N_4122,In_1127,In_774);
nor U4123 (N_4123,In_392,In_1383);
or U4124 (N_4124,In_681,In_1769);
and U4125 (N_4125,In_45,In_912);
nand U4126 (N_4126,In_2339,In_2853);
nor U4127 (N_4127,In_2898,In_1253);
or U4128 (N_4128,In_122,In_2412);
nand U4129 (N_4129,In_1572,In_638);
nand U4130 (N_4130,In_2867,In_2605);
xor U4131 (N_4131,In_2896,In_2050);
and U4132 (N_4132,In_1515,In_1949);
xnor U4133 (N_4133,In_2329,In_906);
nand U4134 (N_4134,In_488,In_1972);
or U4135 (N_4135,In_2682,In_170);
nand U4136 (N_4136,In_2679,In_2394);
or U4137 (N_4137,In_2816,In_2876);
or U4138 (N_4138,In_2285,In_2363);
and U4139 (N_4139,In_2472,In_535);
or U4140 (N_4140,In_2516,In_2997);
or U4141 (N_4141,In_1857,In_1933);
or U4142 (N_4142,In_2297,In_2259);
or U4143 (N_4143,In_2132,In_1751);
xnor U4144 (N_4144,In_820,In_428);
xnor U4145 (N_4145,In_2135,In_231);
nand U4146 (N_4146,In_2073,In_1357);
xor U4147 (N_4147,In_1680,In_2306);
nand U4148 (N_4148,In_2745,In_2301);
or U4149 (N_4149,In_1265,In_2522);
nand U4150 (N_4150,In_37,In_818);
xnor U4151 (N_4151,In_62,In_362);
xor U4152 (N_4152,In_1012,In_134);
and U4153 (N_4153,In_99,In_416);
nor U4154 (N_4154,In_402,In_1493);
xnor U4155 (N_4155,In_1890,In_1987);
or U4156 (N_4156,In_1210,In_2110);
nand U4157 (N_4157,In_616,In_1911);
nand U4158 (N_4158,In_1222,In_2609);
or U4159 (N_4159,In_1793,In_2852);
nor U4160 (N_4160,In_1824,In_1944);
nor U4161 (N_4161,In_2277,In_1975);
and U4162 (N_4162,In_1769,In_271);
nor U4163 (N_4163,In_899,In_2418);
and U4164 (N_4164,In_73,In_1025);
or U4165 (N_4165,In_1650,In_2749);
and U4166 (N_4166,In_143,In_242);
and U4167 (N_4167,In_1182,In_587);
nor U4168 (N_4168,In_2481,In_1452);
xnor U4169 (N_4169,In_2436,In_2202);
nand U4170 (N_4170,In_2446,In_1691);
xor U4171 (N_4171,In_865,In_342);
or U4172 (N_4172,In_2114,In_787);
and U4173 (N_4173,In_951,In_1300);
xnor U4174 (N_4174,In_1615,In_1851);
nand U4175 (N_4175,In_1041,In_1621);
nand U4176 (N_4176,In_1657,In_732);
nor U4177 (N_4177,In_1639,In_2379);
nand U4178 (N_4178,In_2827,In_1450);
or U4179 (N_4179,In_774,In_2361);
xor U4180 (N_4180,In_2641,In_2625);
nor U4181 (N_4181,In_245,In_1469);
and U4182 (N_4182,In_944,In_497);
nand U4183 (N_4183,In_854,In_2697);
nand U4184 (N_4184,In_1064,In_1626);
nand U4185 (N_4185,In_1694,In_531);
xor U4186 (N_4186,In_333,In_2518);
xor U4187 (N_4187,In_2874,In_2619);
nand U4188 (N_4188,In_327,In_333);
or U4189 (N_4189,In_1660,In_186);
nor U4190 (N_4190,In_2283,In_1576);
or U4191 (N_4191,In_819,In_2056);
and U4192 (N_4192,In_1278,In_2198);
and U4193 (N_4193,In_1207,In_861);
or U4194 (N_4194,In_1395,In_1476);
and U4195 (N_4195,In_2558,In_1753);
nor U4196 (N_4196,In_2976,In_117);
xnor U4197 (N_4197,In_1849,In_1102);
nor U4198 (N_4198,In_2193,In_1097);
xnor U4199 (N_4199,In_744,In_2620);
nand U4200 (N_4200,In_2770,In_1910);
xor U4201 (N_4201,In_1472,In_918);
xor U4202 (N_4202,In_1432,In_753);
or U4203 (N_4203,In_2909,In_190);
or U4204 (N_4204,In_1121,In_2443);
xnor U4205 (N_4205,In_295,In_1524);
nand U4206 (N_4206,In_1682,In_2098);
nor U4207 (N_4207,In_109,In_1664);
or U4208 (N_4208,In_2520,In_1419);
nor U4209 (N_4209,In_2444,In_892);
or U4210 (N_4210,In_458,In_488);
nand U4211 (N_4211,In_154,In_1803);
xnor U4212 (N_4212,In_733,In_1501);
xor U4213 (N_4213,In_728,In_993);
and U4214 (N_4214,In_87,In_1240);
or U4215 (N_4215,In_1668,In_80);
nor U4216 (N_4216,In_1725,In_1326);
nand U4217 (N_4217,In_1787,In_975);
xor U4218 (N_4218,In_529,In_2657);
and U4219 (N_4219,In_2441,In_1326);
or U4220 (N_4220,In_970,In_1143);
or U4221 (N_4221,In_1289,In_2067);
nand U4222 (N_4222,In_1927,In_492);
and U4223 (N_4223,In_2644,In_553);
or U4224 (N_4224,In_1242,In_931);
or U4225 (N_4225,In_1790,In_2184);
nor U4226 (N_4226,In_154,In_2017);
nor U4227 (N_4227,In_2462,In_2629);
nor U4228 (N_4228,In_2345,In_1815);
nor U4229 (N_4229,In_2481,In_2997);
xnor U4230 (N_4230,In_2881,In_1368);
and U4231 (N_4231,In_1944,In_1067);
nor U4232 (N_4232,In_2433,In_504);
or U4233 (N_4233,In_1403,In_1904);
or U4234 (N_4234,In_263,In_489);
and U4235 (N_4235,In_981,In_729);
nor U4236 (N_4236,In_2681,In_386);
nand U4237 (N_4237,In_2868,In_1834);
or U4238 (N_4238,In_2619,In_200);
and U4239 (N_4239,In_1536,In_1187);
or U4240 (N_4240,In_884,In_2760);
xor U4241 (N_4241,In_808,In_2566);
xnor U4242 (N_4242,In_362,In_434);
or U4243 (N_4243,In_2702,In_923);
nor U4244 (N_4244,In_477,In_1344);
xor U4245 (N_4245,In_1876,In_1731);
nand U4246 (N_4246,In_2712,In_2226);
xor U4247 (N_4247,In_920,In_1708);
or U4248 (N_4248,In_2998,In_1911);
nor U4249 (N_4249,In_508,In_1754);
and U4250 (N_4250,In_2703,In_1551);
nand U4251 (N_4251,In_984,In_2996);
xnor U4252 (N_4252,In_1848,In_2529);
and U4253 (N_4253,In_2238,In_2117);
nor U4254 (N_4254,In_659,In_2903);
and U4255 (N_4255,In_1921,In_2475);
or U4256 (N_4256,In_2697,In_2658);
and U4257 (N_4257,In_2135,In_2042);
nand U4258 (N_4258,In_1418,In_2416);
and U4259 (N_4259,In_623,In_2892);
or U4260 (N_4260,In_714,In_1501);
and U4261 (N_4261,In_634,In_2727);
nor U4262 (N_4262,In_2302,In_479);
nand U4263 (N_4263,In_2818,In_2025);
nand U4264 (N_4264,In_1985,In_300);
or U4265 (N_4265,In_667,In_1627);
xnor U4266 (N_4266,In_164,In_1168);
nor U4267 (N_4267,In_1777,In_911);
nor U4268 (N_4268,In_2284,In_2130);
xor U4269 (N_4269,In_815,In_786);
and U4270 (N_4270,In_1442,In_1582);
nand U4271 (N_4271,In_768,In_2334);
nor U4272 (N_4272,In_1172,In_879);
nor U4273 (N_4273,In_2632,In_1022);
xor U4274 (N_4274,In_243,In_2731);
or U4275 (N_4275,In_392,In_27);
and U4276 (N_4276,In_1501,In_1743);
xnor U4277 (N_4277,In_2804,In_1020);
nand U4278 (N_4278,In_2859,In_2959);
or U4279 (N_4279,In_1791,In_686);
or U4280 (N_4280,In_926,In_155);
nor U4281 (N_4281,In_2487,In_2308);
and U4282 (N_4282,In_1912,In_516);
nor U4283 (N_4283,In_2687,In_380);
or U4284 (N_4284,In_666,In_2442);
and U4285 (N_4285,In_760,In_1214);
xnor U4286 (N_4286,In_2258,In_1247);
nand U4287 (N_4287,In_1230,In_188);
or U4288 (N_4288,In_1230,In_1753);
nor U4289 (N_4289,In_849,In_2776);
or U4290 (N_4290,In_1057,In_1560);
nand U4291 (N_4291,In_19,In_997);
nor U4292 (N_4292,In_2322,In_2151);
xor U4293 (N_4293,In_1365,In_277);
nand U4294 (N_4294,In_998,In_618);
nand U4295 (N_4295,In_2618,In_971);
or U4296 (N_4296,In_1301,In_2900);
xor U4297 (N_4297,In_25,In_2394);
or U4298 (N_4298,In_2238,In_1821);
nor U4299 (N_4299,In_273,In_323);
and U4300 (N_4300,In_2339,In_1825);
nor U4301 (N_4301,In_838,In_2057);
and U4302 (N_4302,In_969,In_2025);
xnor U4303 (N_4303,In_1660,In_2721);
nor U4304 (N_4304,In_1706,In_742);
and U4305 (N_4305,In_1091,In_1942);
nor U4306 (N_4306,In_125,In_814);
nor U4307 (N_4307,In_4,In_2128);
nand U4308 (N_4308,In_1646,In_546);
nand U4309 (N_4309,In_115,In_182);
and U4310 (N_4310,In_1195,In_2385);
or U4311 (N_4311,In_2012,In_2434);
or U4312 (N_4312,In_2991,In_2634);
nor U4313 (N_4313,In_1949,In_1224);
nor U4314 (N_4314,In_642,In_1020);
xnor U4315 (N_4315,In_791,In_1471);
xor U4316 (N_4316,In_2902,In_1732);
and U4317 (N_4317,In_1202,In_169);
or U4318 (N_4318,In_2834,In_797);
nand U4319 (N_4319,In_362,In_2074);
nand U4320 (N_4320,In_464,In_1368);
or U4321 (N_4321,In_2152,In_1144);
nor U4322 (N_4322,In_1988,In_2025);
nand U4323 (N_4323,In_2814,In_2114);
and U4324 (N_4324,In_1481,In_683);
xnor U4325 (N_4325,In_2527,In_2321);
nand U4326 (N_4326,In_143,In_2316);
xnor U4327 (N_4327,In_1113,In_2343);
nand U4328 (N_4328,In_688,In_2310);
nor U4329 (N_4329,In_417,In_1426);
nand U4330 (N_4330,In_2117,In_821);
xor U4331 (N_4331,In_2798,In_1637);
nand U4332 (N_4332,In_107,In_814);
or U4333 (N_4333,In_2871,In_1525);
and U4334 (N_4334,In_762,In_2546);
nand U4335 (N_4335,In_2165,In_2813);
or U4336 (N_4336,In_671,In_336);
nor U4337 (N_4337,In_2088,In_1208);
or U4338 (N_4338,In_2870,In_107);
or U4339 (N_4339,In_584,In_162);
or U4340 (N_4340,In_717,In_1853);
nor U4341 (N_4341,In_2671,In_2596);
nor U4342 (N_4342,In_1209,In_739);
xnor U4343 (N_4343,In_851,In_1475);
nand U4344 (N_4344,In_11,In_157);
or U4345 (N_4345,In_2302,In_1333);
and U4346 (N_4346,In_283,In_357);
nor U4347 (N_4347,In_2186,In_2654);
and U4348 (N_4348,In_1238,In_378);
nand U4349 (N_4349,In_2090,In_1094);
nor U4350 (N_4350,In_2895,In_1077);
nand U4351 (N_4351,In_708,In_1881);
or U4352 (N_4352,In_1998,In_194);
and U4353 (N_4353,In_1354,In_2821);
xor U4354 (N_4354,In_515,In_908);
nor U4355 (N_4355,In_1350,In_365);
nand U4356 (N_4356,In_803,In_2182);
nor U4357 (N_4357,In_1257,In_35);
or U4358 (N_4358,In_373,In_2742);
xnor U4359 (N_4359,In_2078,In_1299);
or U4360 (N_4360,In_1680,In_947);
nand U4361 (N_4361,In_1872,In_2887);
nor U4362 (N_4362,In_2963,In_1248);
nand U4363 (N_4363,In_1681,In_2754);
xnor U4364 (N_4364,In_2254,In_676);
xnor U4365 (N_4365,In_1872,In_2917);
nor U4366 (N_4366,In_1987,In_2502);
nand U4367 (N_4367,In_1421,In_2355);
or U4368 (N_4368,In_1198,In_1668);
xor U4369 (N_4369,In_1480,In_314);
nor U4370 (N_4370,In_2348,In_2924);
xnor U4371 (N_4371,In_555,In_315);
or U4372 (N_4372,In_1985,In_1467);
nand U4373 (N_4373,In_816,In_2122);
and U4374 (N_4374,In_2313,In_1749);
and U4375 (N_4375,In_1974,In_713);
and U4376 (N_4376,In_2968,In_1519);
or U4377 (N_4377,In_62,In_792);
and U4378 (N_4378,In_1987,In_2537);
xnor U4379 (N_4379,In_838,In_1902);
and U4380 (N_4380,In_792,In_597);
nand U4381 (N_4381,In_1714,In_745);
nand U4382 (N_4382,In_1700,In_2219);
or U4383 (N_4383,In_928,In_444);
and U4384 (N_4384,In_1229,In_249);
nand U4385 (N_4385,In_1859,In_141);
nand U4386 (N_4386,In_2777,In_1754);
nand U4387 (N_4387,In_2160,In_1481);
xnor U4388 (N_4388,In_2151,In_719);
nand U4389 (N_4389,In_1931,In_1059);
xnor U4390 (N_4390,In_319,In_2814);
xnor U4391 (N_4391,In_1962,In_7);
nor U4392 (N_4392,In_868,In_1425);
or U4393 (N_4393,In_1980,In_1813);
nand U4394 (N_4394,In_2930,In_60);
xnor U4395 (N_4395,In_1454,In_706);
nand U4396 (N_4396,In_2951,In_650);
nand U4397 (N_4397,In_529,In_182);
xor U4398 (N_4398,In_2797,In_552);
and U4399 (N_4399,In_1943,In_2088);
or U4400 (N_4400,In_1628,In_1878);
and U4401 (N_4401,In_2458,In_246);
xor U4402 (N_4402,In_774,In_20);
nor U4403 (N_4403,In_2975,In_1033);
or U4404 (N_4404,In_2887,In_489);
and U4405 (N_4405,In_1395,In_780);
nor U4406 (N_4406,In_976,In_657);
and U4407 (N_4407,In_2417,In_121);
or U4408 (N_4408,In_1076,In_210);
or U4409 (N_4409,In_1792,In_269);
xor U4410 (N_4410,In_13,In_465);
or U4411 (N_4411,In_1349,In_638);
or U4412 (N_4412,In_2355,In_1123);
and U4413 (N_4413,In_2131,In_2505);
nor U4414 (N_4414,In_1859,In_2898);
or U4415 (N_4415,In_1190,In_684);
xor U4416 (N_4416,In_917,In_2660);
nor U4417 (N_4417,In_1673,In_1845);
and U4418 (N_4418,In_1942,In_1524);
or U4419 (N_4419,In_2156,In_2017);
nand U4420 (N_4420,In_1321,In_2571);
and U4421 (N_4421,In_882,In_1538);
nor U4422 (N_4422,In_2825,In_693);
and U4423 (N_4423,In_505,In_1319);
or U4424 (N_4424,In_2597,In_1689);
and U4425 (N_4425,In_775,In_2088);
nand U4426 (N_4426,In_1070,In_583);
xnor U4427 (N_4427,In_1374,In_2997);
or U4428 (N_4428,In_2526,In_566);
nor U4429 (N_4429,In_2299,In_2216);
or U4430 (N_4430,In_2350,In_686);
nor U4431 (N_4431,In_798,In_2954);
and U4432 (N_4432,In_1609,In_863);
and U4433 (N_4433,In_2027,In_2261);
nand U4434 (N_4434,In_1510,In_1020);
xor U4435 (N_4435,In_154,In_1286);
nor U4436 (N_4436,In_545,In_800);
and U4437 (N_4437,In_2241,In_1635);
nor U4438 (N_4438,In_360,In_2114);
nor U4439 (N_4439,In_751,In_1955);
xor U4440 (N_4440,In_590,In_1058);
nand U4441 (N_4441,In_289,In_2451);
xnor U4442 (N_4442,In_1693,In_1074);
nand U4443 (N_4443,In_2857,In_2226);
or U4444 (N_4444,In_1545,In_1129);
nand U4445 (N_4445,In_1086,In_2370);
nor U4446 (N_4446,In_2564,In_2507);
xnor U4447 (N_4447,In_1109,In_336);
or U4448 (N_4448,In_19,In_292);
nor U4449 (N_4449,In_621,In_1163);
xnor U4450 (N_4450,In_1789,In_2609);
nor U4451 (N_4451,In_1176,In_1816);
and U4452 (N_4452,In_655,In_2699);
xor U4453 (N_4453,In_1709,In_588);
or U4454 (N_4454,In_2420,In_2013);
nor U4455 (N_4455,In_1510,In_202);
nor U4456 (N_4456,In_2378,In_471);
or U4457 (N_4457,In_2934,In_2415);
nor U4458 (N_4458,In_714,In_1999);
xnor U4459 (N_4459,In_2199,In_2766);
xor U4460 (N_4460,In_2893,In_1950);
or U4461 (N_4461,In_764,In_2524);
xnor U4462 (N_4462,In_734,In_2956);
nand U4463 (N_4463,In_1120,In_537);
and U4464 (N_4464,In_505,In_541);
nand U4465 (N_4465,In_1573,In_1334);
nor U4466 (N_4466,In_1722,In_679);
and U4467 (N_4467,In_990,In_1952);
or U4468 (N_4468,In_2603,In_1515);
nand U4469 (N_4469,In_2230,In_2011);
xor U4470 (N_4470,In_1190,In_1518);
nor U4471 (N_4471,In_1036,In_1085);
or U4472 (N_4472,In_571,In_1512);
or U4473 (N_4473,In_162,In_1218);
nand U4474 (N_4474,In_1929,In_687);
nor U4475 (N_4475,In_1734,In_24);
and U4476 (N_4476,In_733,In_1947);
or U4477 (N_4477,In_1295,In_2129);
nor U4478 (N_4478,In_1073,In_1405);
xnor U4479 (N_4479,In_2776,In_795);
nand U4480 (N_4480,In_239,In_121);
or U4481 (N_4481,In_2769,In_718);
or U4482 (N_4482,In_624,In_1238);
and U4483 (N_4483,In_1055,In_1548);
nor U4484 (N_4484,In_662,In_2453);
and U4485 (N_4485,In_694,In_2997);
and U4486 (N_4486,In_1253,In_2241);
and U4487 (N_4487,In_839,In_352);
nand U4488 (N_4488,In_164,In_2216);
and U4489 (N_4489,In_241,In_386);
or U4490 (N_4490,In_2705,In_2178);
and U4491 (N_4491,In_2200,In_1169);
xor U4492 (N_4492,In_686,In_1924);
nand U4493 (N_4493,In_1879,In_1160);
and U4494 (N_4494,In_762,In_2040);
xnor U4495 (N_4495,In_1236,In_87);
xor U4496 (N_4496,In_2672,In_1385);
and U4497 (N_4497,In_97,In_934);
nor U4498 (N_4498,In_1210,In_2662);
or U4499 (N_4499,In_1796,In_1936);
nor U4500 (N_4500,In_2839,In_1323);
and U4501 (N_4501,In_1834,In_1420);
nand U4502 (N_4502,In_1494,In_933);
nand U4503 (N_4503,In_1435,In_2584);
nand U4504 (N_4504,In_2552,In_423);
or U4505 (N_4505,In_556,In_2076);
nand U4506 (N_4506,In_187,In_2628);
nand U4507 (N_4507,In_2332,In_1543);
nor U4508 (N_4508,In_163,In_2330);
nand U4509 (N_4509,In_642,In_283);
and U4510 (N_4510,In_2545,In_2131);
nand U4511 (N_4511,In_1961,In_167);
xor U4512 (N_4512,In_2848,In_1741);
xnor U4513 (N_4513,In_2932,In_2535);
or U4514 (N_4514,In_2443,In_1244);
and U4515 (N_4515,In_529,In_1010);
and U4516 (N_4516,In_928,In_1209);
or U4517 (N_4517,In_2619,In_876);
and U4518 (N_4518,In_986,In_2812);
xor U4519 (N_4519,In_2862,In_741);
nor U4520 (N_4520,In_1301,In_721);
nand U4521 (N_4521,In_2945,In_1446);
or U4522 (N_4522,In_2990,In_1702);
xor U4523 (N_4523,In_2385,In_1535);
xnor U4524 (N_4524,In_2279,In_96);
xor U4525 (N_4525,In_1285,In_1045);
nand U4526 (N_4526,In_1417,In_1725);
xor U4527 (N_4527,In_2228,In_1382);
or U4528 (N_4528,In_1719,In_2482);
or U4529 (N_4529,In_2423,In_1895);
or U4530 (N_4530,In_1704,In_1179);
or U4531 (N_4531,In_1280,In_484);
nand U4532 (N_4532,In_1960,In_2877);
or U4533 (N_4533,In_2229,In_1028);
or U4534 (N_4534,In_110,In_1585);
nor U4535 (N_4535,In_114,In_169);
xor U4536 (N_4536,In_970,In_2629);
and U4537 (N_4537,In_1418,In_2339);
nor U4538 (N_4538,In_1979,In_112);
nand U4539 (N_4539,In_773,In_1659);
xnor U4540 (N_4540,In_1144,In_399);
nor U4541 (N_4541,In_2759,In_958);
xor U4542 (N_4542,In_2490,In_416);
nand U4543 (N_4543,In_975,In_2974);
and U4544 (N_4544,In_1575,In_148);
nor U4545 (N_4545,In_1078,In_937);
and U4546 (N_4546,In_2066,In_2301);
and U4547 (N_4547,In_1046,In_715);
xnor U4548 (N_4548,In_1888,In_2445);
nand U4549 (N_4549,In_2046,In_984);
or U4550 (N_4550,In_922,In_680);
or U4551 (N_4551,In_1566,In_130);
nor U4552 (N_4552,In_2000,In_2913);
xnor U4553 (N_4553,In_1450,In_2012);
nor U4554 (N_4554,In_2681,In_1023);
nor U4555 (N_4555,In_271,In_2298);
nand U4556 (N_4556,In_2468,In_966);
or U4557 (N_4557,In_1548,In_2001);
and U4558 (N_4558,In_956,In_2362);
nor U4559 (N_4559,In_365,In_1728);
nand U4560 (N_4560,In_1319,In_488);
nor U4561 (N_4561,In_1548,In_2208);
xnor U4562 (N_4562,In_890,In_1534);
nand U4563 (N_4563,In_2673,In_2801);
xor U4564 (N_4564,In_2574,In_1745);
nor U4565 (N_4565,In_1221,In_2250);
and U4566 (N_4566,In_1835,In_1238);
nand U4567 (N_4567,In_2885,In_2999);
nor U4568 (N_4568,In_1010,In_2272);
xnor U4569 (N_4569,In_2186,In_2020);
and U4570 (N_4570,In_1245,In_945);
nand U4571 (N_4571,In_2507,In_61);
and U4572 (N_4572,In_2767,In_447);
or U4573 (N_4573,In_1546,In_116);
and U4574 (N_4574,In_2514,In_1344);
nand U4575 (N_4575,In_1231,In_1743);
xnor U4576 (N_4576,In_1686,In_10);
or U4577 (N_4577,In_2620,In_2769);
nor U4578 (N_4578,In_2131,In_2479);
xnor U4579 (N_4579,In_2515,In_2388);
and U4580 (N_4580,In_829,In_68);
xnor U4581 (N_4581,In_447,In_706);
xnor U4582 (N_4582,In_91,In_2175);
or U4583 (N_4583,In_2172,In_1948);
nor U4584 (N_4584,In_834,In_1947);
nor U4585 (N_4585,In_1387,In_782);
and U4586 (N_4586,In_2521,In_908);
or U4587 (N_4587,In_2095,In_1572);
nand U4588 (N_4588,In_2737,In_1890);
and U4589 (N_4589,In_855,In_160);
nor U4590 (N_4590,In_1579,In_2530);
nand U4591 (N_4591,In_1151,In_166);
nor U4592 (N_4592,In_727,In_1169);
nor U4593 (N_4593,In_194,In_865);
and U4594 (N_4594,In_961,In_2531);
xor U4595 (N_4595,In_2605,In_485);
and U4596 (N_4596,In_288,In_329);
and U4597 (N_4597,In_423,In_1994);
or U4598 (N_4598,In_862,In_2444);
and U4599 (N_4599,In_1417,In_1774);
nor U4600 (N_4600,In_261,In_1030);
nand U4601 (N_4601,In_1626,In_773);
and U4602 (N_4602,In_2018,In_749);
nor U4603 (N_4603,In_1690,In_1469);
nand U4604 (N_4604,In_833,In_2968);
or U4605 (N_4605,In_2255,In_2320);
and U4606 (N_4606,In_1195,In_2232);
xnor U4607 (N_4607,In_85,In_2784);
or U4608 (N_4608,In_1847,In_1568);
nor U4609 (N_4609,In_2705,In_604);
and U4610 (N_4610,In_163,In_2750);
nand U4611 (N_4611,In_2336,In_1315);
xor U4612 (N_4612,In_2946,In_1652);
nand U4613 (N_4613,In_2893,In_2964);
and U4614 (N_4614,In_330,In_121);
nand U4615 (N_4615,In_61,In_2329);
and U4616 (N_4616,In_267,In_1021);
xor U4617 (N_4617,In_976,In_1900);
nand U4618 (N_4618,In_2586,In_669);
and U4619 (N_4619,In_1405,In_1923);
nor U4620 (N_4620,In_1419,In_244);
and U4621 (N_4621,In_1346,In_2416);
or U4622 (N_4622,In_10,In_1216);
and U4623 (N_4623,In_2951,In_180);
and U4624 (N_4624,In_562,In_805);
and U4625 (N_4625,In_2366,In_1724);
nor U4626 (N_4626,In_346,In_2984);
and U4627 (N_4627,In_1779,In_1551);
or U4628 (N_4628,In_2764,In_1167);
nand U4629 (N_4629,In_904,In_2041);
or U4630 (N_4630,In_694,In_1404);
nor U4631 (N_4631,In_706,In_1569);
or U4632 (N_4632,In_1285,In_1963);
or U4633 (N_4633,In_389,In_810);
or U4634 (N_4634,In_1164,In_282);
and U4635 (N_4635,In_957,In_2402);
and U4636 (N_4636,In_952,In_1990);
xor U4637 (N_4637,In_1141,In_2979);
nor U4638 (N_4638,In_1024,In_1642);
and U4639 (N_4639,In_1417,In_1269);
nand U4640 (N_4640,In_1503,In_776);
and U4641 (N_4641,In_81,In_591);
xor U4642 (N_4642,In_2277,In_194);
nor U4643 (N_4643,In_2183,In_1320);
xnor U4644 (N_4644,In_2894,In_2892);
nor U4645 (N_4645,In_2093,In_2092);
xor U4646 (N_4646,In_451,In_1983);
nor U4647 (N_4647,In_145,In_2388);
nor U4648 (N_4648,In_2155,In_912);
or U4649 (N_4649,In_695,In_2035);
or U4650 (N_4650,In_2633,In_2829);
nor U4651 (N_4651,In_2084,In_1566);
nor U4652 (N_4652,In_2379,In_1091);
xnor U4653 (N_4653,In_1539,In_2996);
xnor U4654 (N_4654,In_2985,In_156);
nor U4655 (N_4655,In_2339,In_2258);
xnor U4656 (N_4656,In_2660,In_843);
nor U4657 (N_4657,In_273,In_2033);
nand U4658 (N_4658,In_163,In_697);
xnor U4659 (N_4659,In_2307,In_665);
or U4660 (N_4660,In_1986,In_54);
xnor U4661 (N_4661,In_147,In_734);
xor U4662 (N_4662,In_529,In_1819);
xor U4663 (N_4663,In_789,In_1894);
nand U4664 (N_4664,In_1038,In_2705);
and U4665 (N_4665,In_1599,In_1712);
nand U4666 (N_4666,In_2022,In_2871);
or U4667 (N_4667,In_2095,In_543);
or U4668 (N_4668,In_2308,In_243);
nand U4669 (N_4669,In_638,In_558);
nor U4670 (N_4670,In_670,In_1814);
nor U4671 (N_4671,In_887,In_861);
nand U4672 (N_4672,In_1093,In_976);
and U4673 (N_4673,In_23,In_1442);
nor U4674 (N_4674,In_2783,In_2967);
nand U4675 (N_4675,In_539,In_2571);
and U4676 (N_4676,In_650,In_494);
or U4677 (N_4677,In_2481,In_371);
xnor U4678 (N_4678,In_623,In_2751);
or U4679 (N_4679,In_2110,In_2551);
xor U4680 (N_4680,In_2340,In_2988);
nor U4681 (N_4681,In_2838,In_806);
and U4682 (N_4682,In_1621,In_1970);
or U4683 (N_4683,In_520,In_2074);
xor U4684 (N_4684,In_2433,In_13);
or U4685 (N_4685,In_1496,In_731);
or U4686 (N_4686,In_753,In_1118);
or U4687 (N_4687,In_2141,In_798);
or U4688 (N_4688,In_1261,In_93);
nand U4689 (N_4689,In_1769,In_1017);
nand U4690 (N_4690,In_2353,In_337);
nand U4691 (N_4691,In_2692,In_504);
nand U4692 (N_4692,In_1543,In_1442);
xor U4693 (N_4693,In_602,In_1661);
nand U4694 (N_4694,In_2643,In_1157);
or U4695 (N_4695,In_1930,In_2623);
nor U4696 (N_4696,In_2779,In_295);
nand U4697 (N_4697,In_2651,In_1906);
xnor U4698 (N_4698,In_98,In_1642);
xnor U4699 (N_4699,In_1971,In_1134);
and U4700 (N_4700,In_2534,In_803);
nor U4701 (N_4701,In_332,In_1845);
nand U4702 (N_4702,In_1912,In_1689);
xor U4703 (N_4703,In_675,In_974);
nand U4704 (N_4704,In_210,In_616);
and U4705 (N_4705,In_2983,In_1622);
or U4706 (N_4706,In_2302,In_1031);
or U4707 (N_4707,In_2495,In_13);
xnor U4708 (N_4708,In_1623,In_2261);
nor U4709 (N_4709,In_1023,In_1752);
or U4710 (N_4710,In_1198,In_1129);
nand U4711 (N_4711,In_2235,In_623);
nand U4712 (N_4712,In_2161,In_1034);
nand U4713 (N_4713,In_1022,In_1608);
xnor U4714 (N_4714,In_978,In_1301);
nand U4715 (N_4715,In_2737,In_411);
xnor U4716 (N_4716,In_1012,In_589);
and U4717 (N_4717,In_940,In_599);
or U4718 (N_4718,In_1185,In_2072);
xor U4719 (N_4719,In_1389,In_1495);
or U4720 (N_4720,In_716,In_2836);
nor U4721 (N_4721,In_2286,In_66);
nor U4722 (N_4722,In_2236,In_1037);
and U4723 (N_4723,In_556,In_1477);
nand U4724 (N_4724,In_2103,In_988);
and U4725 (N_4725,In_2193,In_969);
nor U4726 (N_4726,In_2685,In_2148);
xnor U4727 (N_4727,In_2497,In_2208);
nor U4728 (N_4728,In_1271,In_850);
xor U4729 (N_4729,In_360,In_1145);
nor U4730 (N_4730,In_325,In_678);
nand U4731 (N_4731,In_333,In_2647);
and U4732 (N_4732,In_2385,In_1752);
nor U4733 (N_4733,In_2538,In_1755);
nand U4734 (N_4734,In_2297,In_801);
nor U4735 (N_4735,In_496,In_2087);
or U4736 (N_4736,In_1995,In_2731);
xnor U4737 (N_4737,In_2998,In_1976);
xor U4738 (N_4738,In_2456,In_86);
xor U4739 (N_4739,In_2888,In_1147);
nand U4740 (N_4740,In_22,In_1232);
or U4741 (N_4741,In_1633,In_164);
xor U4742 (N_4742,In_1836,In_1076);
or U4743 (N_4743,In_1285,In_2355);
xnor U4744 (N_4744,In_975,In_1172);
and U4745 (N_4745,In_2836,In_2998);
or U4746 (N_4746,In_2866,In_1866);
xnor U4747 (N_4747,In_1471,In_1540);
or U4748 (N_4748,In_920,In_2998);
xor U4749 (N_4749,In_607,In_2969);
xnor U4750 (N_4750,In_2572,In_2605);
nor U4751 (N_4751,In_1692,In_1820);
xnor U4752 (N_4752,In_682,In_414);
nand U4753 (N_4753,In_157,In_819);
nand U4754 (N_4754,In_2770,In_2581);
nand U4755 (N_4755,In_2606,In_640);
nand U4756 (N_4756,In_1661,In_1013);
xor U4757 (N_4757,In_1250,In_1614);
nand U4758 (N_4758,In_2143,In_1160);
and U4759 (N_4759,In_459,In_2107);
or U4760 (N_4760,In_2443,In_1046);
nor U4761 (N_4761,In_1789,In_327);
xor U4762 (N_4762,In_2059,In_360);
and U4763 (N_4763,In_2899,In_2867);
nand U4764 (N_4764,In_2676,In_2188);
and U4765 (N_4765,In_2234,In_30);
and U4766 (N_4766,In_2506,In_251);
xnor U4767 (N_4767,In_1050,In_2940);
nor U4768 (N_4768,In_2133,In_1772);
and U4769 (N_4769,In_2954,In_2759);
or U4770 (N_4770,In_1483,In_1231);
or U4771 (N_4771,In_2378,In_1001);
or U4772 (N_4772,In_1956,In_1073);
nand U4773 (N_4773,In_2910,In_1491);
and U4774 (N_4774,In_1164,In_982);
xor U4775 (N_4775,In_1412,In_1008);
or U4776 (N_4776,In_2422,In_1733);
or U4777 (N_4777,In_5,In_1060);
nor U4778 (N_4778,In_1551,In_119);
xnor U4779 (N_4779,In_1374,In_1556);
nor U4780 (N_4780,In_344,In_1546);
or U4781 (N_4781,In_2497,In_2556);
and U4782 (N_4782,In_368,In_2317);
nand U4783 (N_4783,In_1112,In_2339);
xnor U4784 (N_4784,In_620,In_1482);
nor U4785 (N_4785,In_2483,In_2836);
nand U4786 (N_4786,In_184,In_1779);
nor U4787 (N_4787,In_1577,In_2498);
nand U4788 (N_4788,In_175,In_2416);
nand U4789 (N_4789,In_1382,In_2184);
nor U4790 (N_4790,In_861,In_495);
nor U4791 (N_4791,In_1435,In_348);
nor U4792 (N_4792,In_1792,In_279);
and U4793 (N_4793,In_2026,In_601);
xor U4794 (N_4794,In_1866,In_1153);
nand U4795 (N_4795,In_904,In_226);
nor U4796 (N_4796,In_367,In_2921);
and U4797 (N_4797,In_2476,In_2408);
nor U4798 (N_4798,In_1862,In_2489);
xor U4799 (N_4799,In_1800,In_1986);
and U4800 (N_4800,In_1680,In_1830);
nand U4801 (N_4801,In_442,In_899);
xor U4802 (N_4802,In_345,In_2194);
nor U4803 (N_4803,In_2990,In_2092);
xnor U4804 (N_4804,In_2236,In_358);
xor U4805 (N_4805,In_427,In_2893);
nand U4806 (N_4806,In_1608,In_1120);
and U4807 (N_4807,In_2500,In_2814);
xnor U4808 (N_4808,In_1786,In_2766);
xor U4809 (N_4809,In_1620,In_1351);
nand U4810 (N_4810,In_2780,In_960);
and U4811 (N_4811,In_2518,In_1258);
nand U4812 (N_4812,In_2244,In_621);
nor U4813 (N_4813,In_2665,In_2092);
xnor U4814 (N_4814,In_14,In_278);
and U4815 (N_4815,In_1790,In_1442);
nor U4816 (N_4816,In_2274,In_361);
or U4817 (N_4817,In_98,In_697);
nor U4818 (N_4818,In_37,In_1352);
nor U4819 (N_4819,In_1654,In_2518);
nor U4820 (N_4820,In_1077,In_1516);
or U4821 (N_4821,In_2756,In_1225);
or U4822 (N_4822,In_480,In_1285);
and U4823 (N_4823,In_1557,In_1400);
and U4824 (N_4824,In_799,In_2274);
or U4825 (N_4825,In_2542,In_1407);
nor U4826 (N_4826,In_1409,In_1965);
and U4827 (N_4827,In_358,In_2497);
nor U4828 (N_4828,In_1167,In_1702);
nand U4829 (N_4829,In_1901,In_1141);
nor U4830 (N_4830,In_1109,In_2898);
nor U4831 (N_4831,In_1890,In_671);
and U4832 (N_4832,In_696,In_2885);
nand U4833 (N_4833,In_1679,In_1020);
and U4834 (N_4834,In_1191,In_2239);
nor U4835 (N_4835,In_1589,In_1865);
nand U4836 (N_4836,In_276,In_142);
or U4837 (N_4837,In_1883,In_1102);
xor U4838 (N_4838,In_1244,In_1038);
nor U4839 (N_4839,In_294,In_1605);
or U4840 (N_4840,In_2946,In_2836);
and U4841 (N_4841,In_2108,In_2239);
or U4842 (N_4842,In_1779,In_1546);
and U4843 (N_4843,In_2813,In_1543);
and U4844 (N_4844,In_2972,In_2164);
nor U4845 (N_4845,In_490,In_1079);
and U4846 (N_4846,In_666,In_2792);
or U4847 (N_4847,In_2104,In_1202);
xor U4848 (N_4848,In_515,In_1806);
nor U4849 (N_4849,In_2758,In_1478);
or U4850 (N_4850,In_674,In_761);
nand U4851 (N_4851,In_1139,In_557);
nor U4852 (N_4852,In_1197,In_1535);
nand U4853 (N_4853,In_997,In_2295);
nand U4854 (N_4854,In_569,In_768);
xor U4855 (N_4855,In_461,In_2586);
nand U4856 (N_4856,In_2637,In_2061);
xor U4857 (N_4857,In_1321,In_2259);
xor U4858 (N_4858,In_1219,In_2489);
xor U4859 (N_4859,In_1726,In_2242);
xnor U4860 (N_4860,In_1022,In_1749);
nor U4861 (N_4861,In_1056,In_2810);
and U4862 (N_4862,In_2959,In_2021);
xnor U4863 (N_4863,In_1190,In_2232);
xnor U4864 (N_4864,In_2935,In_625);
nand U4865 (N_4865,In_1915,In_2632);
and U4866 (N_4866,In_551,In_1903);
nand U4867 (N_4867,In_1782,In_2304);
xor U4868 (N_4868,In_1951,In_1077);
and U4869 (N_4869,In_2859,In_309);
or U4870 (N_4870,In_1516,In_2550);
xor U4871 (N_4871,In_2099,In_453);
or U4872 (N_4872,In_492,In_2619);
and U4873 (N_4873,In_1718,In_2921);
or U4874 (N_4874,In_1284,In_1240);
xnor U4875 (N_4875,In_2221,In_1595);
xor U4876 (N_4876,In_2285,In_550);
and U4877 (N_4877,In_1658,In_728);
and U4878 (N_4878,In_1367,In_1279);
nor U4879 (N_4879,In_2509,In_1307);
or U4880 (N_4880,In_467,In_983);
xnor U4881 (N_4881,In_168,In_258);
and U4882 (N_4882,In_657,In_1005);
and U4883 (N_4883,In_399,In_783);
nand U4884 (N_4884,In_671,In_2451);
xnor U4885 (N_4885,In_2257,In_2311);
or U4886 (N_4886,In_885,In_1590);
xor U4887 (N_4887,In_1604,In_243);
nor U4888 (N_4888,In_2494,In_2556);
nand U4889 (N_4889,In_803,In_2134);
or U4890 (N_4890,In_932,In_640);
or U4891 (N_4891,In_1925,In_1342);
or U4892 (N_4892,In_1990,In_825);
or U4893 (N_4893,In_990,In_2684);
nand U4894 (N_4894,In_1108,In_813);
nor U4895 (N_4895,In_2461,In_1710);
xor U4896 (N_4896,In_924,In_1021);
xor U4897 (N_4897,In_2041,In_2465);
and U4898 (N_4898,In_2344,In_1427);
nand U4899 (N_4899,In_2094,In_2658);
nor U4900 (N_4900,In_1381,In_656);
or U4901 (N_4901,In_1634,In_508);
and U4902 (N_4902,In_621,In_928);
and U4903 (N_4903,In_937,In_1660);
xnor U4904 (N_4904,In_560,In_2150);
or U4905 (N_4905,In_2801,In_2161);
nor U4906 (N_4906,In_1849,In_413);
xnor U4907 (N_4907,In_1324,In_1658);
or U4908 (N_4908,In_2582,In_796);
or U4909 (N_4909,In_2034,In_1893);
and U4910 (N_4910,In_2696,In_2212);
xor U4911 (N_4911,In_1962,In_2806);
nand U4912 (N_4912,In_773,In_2775);
and U4913 (N_4913,In_2620,In_438);
and U4914 (N_4914,In_2796,In_2394);
or U4915 (N_4915,In_1118,In_19);
nand U4916 (N_4916,In_945,In_2977);
or U4917 (N_4917,In_2946,In_2462);
nand U4918 (N_4918,In_2301,In_1001);
and U4919 (N_4919,In_52,In_130);
nand U4920 (N_4920,In_1482,In_413);
nand U4921 (N_4921,In_2793,In_2288);
or U4922 (N_4922,In_1578,In_1403);
xnor U4923 (N_4923,In_2727,In_1820);
nor U4924 (N_4924,In_1435,In_1964);
nand U4925 (N_4925,In_1148,In_1398);
nor U4926 (N_4926,In_808,In_1163);
nor U4927 (N_4927,In_1838,In_284);
xnor U4928 (N_4928,In_1675,In_2736);
and U4929 (N_4929,In_380,In_1064);
or U4930 (N_4930,In_2034,In_2809);
or U4931 (N_4931,In_1476,In_758);
nand U4932 (N_4932,In_1703,In_82);
or U4933 (N_4933,In_2496,In_2792);
xor U4934 (N_4934,In_2695,In_367);
or U4935 (N_4935,In_413,In_2109);
or U4936 (N_4936,In_228,In_491);
xnor U4937 (N_4937,In_2550,In_381);
or U4938 (N_4938,In_2550,In_2492);
nor U4939 (N_4939,In_2183,In_2516);
nor U4940 (N_4940,In_322,In_1472);
or U4941 (N_4941,In_587,In_522);
nor U4942 (N_4942,In_1453,In_2553);
xor U4943 (N_4943,In_2544,In_956);
or U4944 (N_4944,In_2604,In_849);
nand U4945 (N_4945,In_1751,In_2458);
nand U4946 (N_4946,In_115,In_2059);
xor U4947 (N_4947,In_2778,In_1560);
nand U4948 (N_4948,In_1070,In_198);
and U4949 (N_4949,In_430,In_1861);
xor U4950 (N_4950,In_1908,In_86);
nor U4951 (N_4951,In_1637,In_846);
xor U4952 (N_4952,In_1954,In_2014);
and U4953 (N_4953,In_203,In_1430);
xnor U4954 (N_4954,In_2788,In_211);
nand U4955 (N_4955,In_977,In_741);
nor U4956 (N_4956,In_1436,In_798);
xnor U4957 (N_4957,In_2807,In_2859);
nand U4958 (N_4958,In_455,In_2407);
xor U4959 (N_4959,In_2111,In_1185);
nor U4960 (N_4960,In_2013,In_879);
and U4961 (N_4961,In_1568,In_327);
or U4962 (N_4962,In_2711,In_1040);
or U4963 (N_4963,In_540,In_2665);
and U4964 (N_4964,In_100,In_2756);
xor U4965 (N_4965,In_1605,In_1075);
and U4966 (N_4966,In_2418,In_2504);
nand U4967 (N_4967,In_629,In_2324);
or U4968 (N_4968,In_1459,In_2215);
xnor U4969 (N_4969,In_769,In_2630);
nand U4970 (N_4970,In_368,In_1287);
or U4971 (N_4971,In_2563,In_1357);
nor U4972 (N_4972,In_726,In_2286);
nand U4973 (N_4973,In_2343,In_1517);
nor U4974 (N_4974,In_2139,In_519);
nand U4975 (N_4975,In_1028,In_961);
or U4976 (N_4976,In_1444,In_942);
and U4977 (N_4977,In_1404,In_1399);
or U4978 (N_4978,In_525,In_289);
xor U4979 (N_4979,In_476,In_2103);
xor U4980 (N_4980,In_1858,In_2313);
nand U4981 (N_4981,In_893,In_607);
and U4982 (N_4982,In_1842,In_249);
nor U4983 (N_4983,In_1115,In_1692);
and U4984 (N_4984,In_207,In_794);
or U4985 (N_4985,In_9,In_3);
nor U4986 (N_4986,In_1436,In_809);
or U4987 (N_4987,In_1193,In_1751);
or U4988 (N_4988,In_2807,In_2501);
xnor U4989 (N_4989,In_2431,In_2062);
nand U4990 (N_4990,In_769,In_2546);
xor U4991 (N_4991,In_2139,In_918);
xor U4992 (N_4992,In_2584,In_2884);
nor U4993 (N_4993,In_893,In_542);
and U4994 (N_4994,In_1754,In_1821);
or U4995 (N_4995,In_1407,In_2364);
and U4996 (N_4996,In_351,In_59);
xor U4997 (N_4997,In_660,In_954);
and U4998 (N_4998,In_153,In_1925);
or U4999 (N_4999,In_1472,In_1621);
and U5000 (N_5000,In_215,In_1736);
nor U5001 (N_5001,In_2101,In_1584);
nor U5002 (N_5002,In_402,In_1970);
nand U5003 (N_5003,In_2880,In_1593);
nor U5004 (N_5004,In_101,In_948);
xnor U5005 (N_5005,In_2916,In_520);
nand U5006 (N_5006,In_2431,In_2375);
nor U5007 (N_5007,In_1461,In_531);
xnor U5008 (N_5008,In_2147,In_332);
and U5009 (N_5009,In_1655,In_412);
xor U5010 (N_5010,In_1458,In_786);
or U5011 (N_5011,In_66,In_335);
xor U5012 (N_5012,In_1148,In_1408);
xor U5013 (N_5013,In_2506,In_2827);
nor U5014 (N_5014,In_1218,In_875);
xor U5015 (N_5015,In_1926,In_252);
xnor U5016 (N_5016,In_166,In_923);
or U5017 (N_5017,In_2595,In_112);
nand U5018 (N_5018,In_2002,In_871);
or U5019 (N_5019,In_1221,In_1741);
nand U5020 (N_5020,In_2780,In_2038);
xnor U5021 (N_5021,In_755,In_1626);
or U5022 (N_5022,In_1689,In_461);
nand U5023 (N_5023,In_195,In_609);
xor U5024 (N_5024,In_1710,In_710);
nand U5025 (N_5025,In_2192,In_1998);
or U5026 (N_5026,In_2031,In_2735);
nand U5027 (N_5027,In_369,In_74);
or U5028 (N_5028,In_1664,In_2444);
nor U5029 (N_5029,In_726,In_2789);
xor U5030 (N_5030,In_2865,In_2622);
and U5031 (N_5031,In_1694,In_1482);
or U5032 (N_5032,In_1558,In_377);
or U5033 (N_5033,In_2826,In_534);
and U5034 (N_5034,In_2322,In_878);
or U5035 (N_5035,In_1970,In_531);
xnor U5036 (N_5036,In_2933,In_2826);
or U5037 (N_5037,In_784,In_130);
nor U5038 (N_5038,In_1346,In_586);
nand U5039 (N_5039,In_2816,In_2922);
xor U5040 (N_5040,In_385,In_2547);
or U5041 (N_5041,In_1548,In_1407);
nor U5042 (N_5042,In_2282,In_2248);
and U5043 (N_5043,In_1000,In_1410);
or U5044 (N_5044,In_1667,In_2131);
nor U5045 (N_5045,In_923,In_14);
and U5046 (N_5046,In_2109,In_840);
and U5047 (N_5047,In_2886,In_2055);
nand U5048 (N_5048,In_119,In_390);
or U5049 (N_5049,In_1620,In_1452);
nor U5050 (N_5050,In_2244,In_822);
xor U5051 (N_5051,In_408,In_1035);
nor U5052 (N_5052,In_2009,In_612);
and U5053 (N_5053,In_37,In_581);
or U5054 (N_5054,In_2427,In_2646);
and U5055 (N_5055,In_2271,In_2822);
nand U5056 (N_5056,In_896,In_2002);
nand U5057 (N_5057,In_1465,In_1519);
nor U5058 (N_5058,In_1127,In_102);
nor U5059 (N_5059,In_1580,In_770);
nand U5060 (N_5060,In_2317,In_272);
nand U5061 (N_5061,In_1109,In_245);
or U5062 (N_5062,In_628,In_1788);
or U5063 (N_5063,In_389,In_321);
or U5064 (N_5064,In_2219,In_2202);
and U5065 (N_5065,In_543,In_2832);
and U5066 (N_5066,In_737,In_2485);
or U5067 (N_5067,In_2545,In_670);
or U5068 (N_5068,In_1276,In_1634);
nand U5069 (N_5069,In_1866,In_1139);
or U5070 (N_5070,In_1694,In_2180);
nand U5071 (N_5071,In_393,In_446);
or U5072 (N_5072,In_222,In_191);
nor U5073 (N_5073,In_264,In_458);
and U5074 (N_5074,In_2516,In_245);
and U5075 (N_5075,In_670,In_520);
nand U5076 (N_5076,In_419,In_448);
nor U5077 (N_5077,In_2725,In_2964);
or U5078 (N_5078,In_1743,In_1775);
xnor U5079 (N_5079,In_349,In_952);
or U5080 (N_5080,In_1044,In_1830);
xnor U5081 (N_5081,In_2413,In_2627);
or U5082 (N_5082,In_2988,In_2825);
xnor U5083 (N_5083,In_566,In_1785);
nor U5084 (N_5084,In_2744,In_2772);
and U5085 (N_5085,In_2366,In_2810);
nor U5086 (N_5086,In_718,In_1798);
and U5087 (N_5087,In_2089,In_2061);
xor U5088 (N_5088,In_1139,In_2195);
nand U5089 (N_5089,In_2808,In_919);
xnor U5090 (N_5090,In_300,In_2133);
and U5091 (N_5091,In_2987,In_101);
xnor U5092 (N_5092,In_580,In_1224);
nor U5093 (N_5093,In_649,In_2067);
nor U5094 (N_5094,In_2894,In_2015);
and U5095 (N_5095,In_1672,In_2327);
and U5096 (N_5096,In_2028,In_610);
nand U5097 (N_5097,In_2365,In_2232);
nand U5098 (N_5098,In_1845,In_948);
nand U5099 (N_5099,In_1577,In_221);
nand U5100 (N_5100,In_806,In_997);
xnor U5101 (N_5101,In_2669,In_281);
and U5102 (N_5102,In_1316,In_1933);
and U5103 (N_5103,In_1970,In_427);
nand U5104 (N_5104,In_487,In_378);
xor U5105 (N_5105,In_2377,In_1574);
nor U5106 (N_5106,In_78,In_943);
nor U5107 (N_5107,In_1299,In_2804);
nor U5108 (N_5108,In_1611,In_71);
or U5109 (N_5109,In_416,In_1722);
or U5110 (N_5110,In_2867,In_1378);
and U5111 (N_5111,In_2431,In_2193);
or U5112 (N_5112,In_865,In_38);
or U5113 (N_5113,In_1269,In_1905);
xnor U5114 (N_5114,In_2272,In_2661);
nand U5115 (N_5115,In_125,In_955);
nand U5116 (N_5116,In_985,In_679);
nor U5117 (N_5117,In_1922,In_2222);
and U5118 (N_5118,In_2152,In_1118);
and U5119 (N_5119,In_1693,In_725);
or U5120 (N_5120,In_1824,In_1729);
nor U5121 (N_5121,In_282,In_2420);
or U5122 (N_5122,In_2171,In_2029);
nand U5123 (N_5123,In_1870,In_2710);
xnor U5124 (N_5124,In_337,In_288);
xnor U5125 (N_5125,In_329,In_1965);
or U5126 (N_5126,In_525,In_35);
and U5127 (N_5127,In_1444,In_2748);
or U5128 (N_5128,In_905,In_554);
or U5129 (N_5129,In_1071,In_1606);
or U5130 (N_5130,In_357,In_1595);
and U5131 (N_5131,In_1681,In_1743);
xnor U5132 (N_5132,In_2730,In_811);
nand U5133 (N_5133,In_479,In_2130);
or U5134 (N_5134,In_72,In_392);
or U5135 (N_5135,In_416,In_2097);
xnor U5136 (N_5136,In_2959,In_1594);
xnor U5137 (N_5137,In_898,In_2857);
and U5138 (N_5138,In_2602,In_1003);
and U5139 (N_5139,In_339,In_1383);
nor U5140 (N_5140,In_1399,In_227);
nor U5141 (N_5141,In_1826,In_831);
and U5142 (N_5142,In_1408,In_2254);
xor U5143 (N_5143,In_614,In_929);
nor U5144 (N_5144,In_2941,In_1375);
xnor U5145 (N_5145,In_845,In_2048);
and U5146 (N_5146,In_186,In_1980);
or U5147 (N_5147,In_2295,In_2999);
nand U5148 (N_5148,In_1266,In_2954);
xor U5149 (N_5149,In_2437,In_651);
and U5150 (N_5150,In_858,In_1005);
nor U5151 (N_5151,In_244,In_1227);
nor U5152 (N_5152,In_249,In_894);
nand U5153 (N_5153,In_191,In_1677);
nor U5154 (N_5154,In_1619,In_2110);
xnor U5155 (N_5155,In_13,In_912);
nor U5156 (N_5156,In_116,In_2596);
nor U5157 (N_5157,In_36,In_1128);
and U5158 (N_5158,In_2124,In_386);
or U5159 (N_5159,In_2289,In_2275);
or U5160 (N_5160,In_2498,In_2738);
or U5161 (N_5161,In_2064,In_2349);
xor U5162 (N_5162,In_991,In_2724);
nor U5163 (N_5163,In_2445,In_1269);
or U5164 (N_5164,In_2770,In_462);
xor U5165 (N_5165,In_2545,In_2973);
and U5166 (N_5166,In_630,In_1350);
xnor U5167 (N_5167,In_967,In_2875);
xor U5168 (N_5168,In_2794,In_2660);
nand U5169 (N_5169,In_1738,In_639);
or U5170 (N_5170,In_268,In_864);
or U5171 (N_5171,In_2442,In_1589);
or U5172 (N_5172,In_88,In_2444);
xnor U5173 (N_5173,In_2362,In_2965);
xnor U5174 (N_5174,In_2111,In_989);
xnor U5175 (N_5175,In_171,In_942);
or U5176 (N_5176,In_194,In_685);
or U5177 (N_5177,In_1447,In_2860);
xnor U5178 (N_5178,In_2687,In_31);
nor U5179 (N_5179,In_498,In_450);
nor U5180 (N_5180,In_814,In_2498);
and U5181 (N_5181,In_79,In_105);
xor U5182 (N_5182,In_726,In_2169);
nand U5183 (N_5183,In_1595,In_1048);
nand U5184 (N_5184,In_1203,In_267);
xor U5185 (N_5185,In_2750,In_1152);
nand U5186 (N_5186,In_716,In_2729);
or U5187 (N_5187,In_2807,In_1336);
and U5188 (N_5188,In_1718,In_1027);
and U5189 (N_5189,In_264,In_1091);
or U5190 (N_5190,In_945,In_658);
nand U5191 (N_5191,In_1592,In_2777);
or U5192 (N_5192,In_1520,In_884);
nor U5193 (N_5193,In_1459,In_2121);
or U5194 (N_5194,In_729,In_1644);
or U5195 (N_5195,In_633,In_2835);
xor U5196 (N_5196,In_884,In_1325);
nand U5197 (N_5197,In_1155,In_937);
xnor U5198 (N_5198,In_1220,In_335);
and U5199 (N_5199,In_346,In_1028);
xnor U5200 (N_5200,In_2703,In_75);
nand U5201 (N_5201,In_1140,In_1100);
xor U5202 (N_5202,In_1518,In_2965);
or U5203 (N_5203,In_210,In_1345);
or U5204 (N_5204,In_600,In_1904);
xor U5205 (N_5205,In_761,In_1260);
nor U5206 (N_5206,In_922,In_2204);
nor U5207 (N_5207,In_1060,In_603);
xnor U5208 (N_5208,In_1071,In_1549);
xor U5209 (N_5209,In_214,In_2183);
nand U5210 (N_5210,In_102,In_315);
nor U5211 (N_5211,In_2954,In_1422);
xor U5212 (N_5212,In_631,In_2884);
and U5213 (N_5213,In_1512,In_2908);
and U5214 (N_5214,In_1191,In_369);
and U5215 (N_5215,In_1903,In_1403);
and U5216 (N_5216,In_1884,In_1274);
nor U5217 (N_5217,In_613,In_1589);
nor U5218 (N_5218,In_1988,In_1750);
xor U5219 (N_5219,In_224,In_2490);
and U5220 (N_5220,In_2546,In_1597);
nand U5221 (N_5221,In_153,In_1649);
xnor U5222 (N_5222,In_672,In_2204);
nand U5223 (N_5223,In_115,In_2709);
nor U5224 (N_5224,In_48,In_1565);
nor U5225 (N_5225,In_2987,In_1976);
nand U5226 (N_5226,In_1187,In_2308);
and U5227 (N_5227,In_735,In_2719);
or U5228 (N_5228,In_2371,In_1896);
and U5229 (N_5229,In_611,In_2572);
nor U5230 (N_5230,In_46,In_577);
xor U5231 (N_5231,In_2524,In_138);
nor U5232 (N_5232,In_1937,In_468);
and U5233 (N_5233,In_428,In_1318);
nand U5234 (N_5234,In_1347,In_209);
xor U5235 (N_5235,In_318,In_1455);
nand U5236 (N_5236,In_1340,In_2520);
and U5237 (N_5237,In_1551,In_1450);
and U5238 (N_5238,In_2455,In_2980);
nor U5239 (N_5239,In_1389,In_1729);
nor U5240 (N_5240,In_468,In_194);
and U5241 (N_5241,In_954,In_355);
nor U5242 (N_5242,In_2783,In_934);
or U5243 (N_5243,In_43,In_978);
nand U5244 (N_5244,In_539,In_953);
nand U5245 (N_5245,In_2269,In_215);
nand U5246 (N_5246,In_2241,In_1761);
or U5247 (N_5247,In_519,In_323);
or U5248 (N_5248,In_1782,In_2032);
nor U5249 (N_5249,In_1362,In_54);
nor U5250 (N_5250,In_207,In_507);
xor U5251 (N_5251,In_673,In_1147);
nor U5252 (N_5252,In_1261,In_1992);
or U5253 (N_5253,In_930,In_425);
and U5254 (N_5254,In_2996,In_808);
nand U5255 (N_5255,In_2061,In_2112);
or U5256 (N_5256,In_605,In_382);
and U5257 (N_5257,In_714,In_1336);
and U5258 (N_5258,In_2389,In_727);
or U5259 (N_5259,In_1073,In_166);
nand U5260 (N_5260,In_302,In_274);
nand U5261 (N_5261,In_2569,In_1272);
nor U5262 (N_5262,In_624,In_2056);
xor U5263 (N_5263,In_1789,In_509);
or U5264 (N_5264,In_403,In_2228);
and U5265 (N_5265,In_6,In_1839);
nand U5266 (N_5266,In_2604,In_2970);
and U5267 (N_5267,In_1017,In_251);
nor U5268 (N_5268,In_1710,In_306);
nor U5269 (N_5269,In_918,In_1859);
and U5270 (N_5270,In_1850,In_2886);
nor U5271 (N_5271,In_1931,In_2275);
nand U5272 (N_5272,In_2596,In_1828);
nor U5273 (N_5273,In_954,In_1901);
nand U5274 (N_5274,In_2944,In_1737);
and U5275 (N_5275,In_416,In_1258);
or U5276 (N_5276,In_2135,In_363);
xor U5277 (N_5277,In_1460,In_1527);
nor U5278 (N_5278,In_1658,In_2420);
or U5279 (N_5279,In_341,In_235);
or U5280 (N_5280,In_1541,In_1358);
xnor U5281 (N_5281,In_1945,In_2527);
and U5282 (N_5282,In_1143,In_276);
nand U5283 (N_5283,In_2709,In_1328);
nor U5284 (N_5284,In_2220,In_2645);
nand U5285 (N_5285,In_1683,In_1707);
nand U5286 (N_5286,In_2118,In_1782);
xor U5287 (N_5287,In_2349,In_1095);
or U5288 (N_5288,In_2893,In_89);
nor U5289 (N_5289,In_552,In_1082);
nand U5290 (N_5290,In_2983,In_578);
nand U5291 (N_5291,In_2196,In_2720);
xnor U5292 (N_5292,In_358,In_670);
or U5293 (N_5293,In_591,In_579);
xor U5294 (N_5294,In_1930,In_2024);
nand U5295 (N_5295,In_54,In_847);
xnor U5296 (N_5296,In_2626,In_2689);
nor U5297 (N_5297,In_2428,In_1237);
or U5298 (N_5298,In_2219,In_1832);
or U5299 (N_5299,In_1062,In_1855);
nand U5300 (N_5300,In_2426,In_2502);
or U5301 (N_5301,In_2398,In_2660);
nand U5302 (N_5302,In_2701,In_1710);
xor U5303 (N_5303,In_65,In_2787);
nand U5304 (N_5304,In_1821,In_135);
or U5305 (N_5305,In_914,In_2339);
xor U5306 (N_5306,In_1794,In_2599);
and U5307 (N_5307,In_937,In_1209);
or U5308 (N_5308,In_2592,In_1908);
or U5309 (N_5309,In_130,In_55);
or U5310 (N_5310,In_736,In_364);
xnor U5311 (N_5311,In_556,In_2017);
nand U5312 (N_5312,In_1941,In_1567);
nand U5313 (N_5313,In_340,In_2771);
nor U5314 (N_5314,In_2113,In_459);
nor U5315 (N_5315,In_1883,In_2049);
nor U5316 (N_5316,In_2601,In_152);
xor U5317 (N_5317,In_2643,In_798);
xor U5318 (N_5318,In_500,In_2071);
and U5319 (N_5319,In_2692,In_831);
xnor U5320 (N_5320,In_330,In_1575);
nand U5321 (N_5321,In_1564,In_1469);
nand U5322 (N_5322,In_832,In_2588);
nor U5323 (N_5323,In_1876,In_1266);
nand U5324 (N_5324,In_1933,In_792);
nand U5325 (N_5325,In_1086,In_1285);
and U5326 (N_5326,In_2464,In_1885);
xnor U5327 (N_5327,In_2064,In_2617);
xnor U5328 (N_5328,In_2203,In_2216);
or U5329 (N_5329,In_246,In_1442);
nand U5330 (N_5330,In_254,In_999);
nand U5331 (N_5331,In_2050,In_1272);
or U5332 (N_5332,In_1603,In_1394);
and U5333 (N_5333,In_1759,In_537);
nor U5334 (N_5334,In_2484,In_2660);
nor U5335 (N_5335,In_452,In_1328);
xnor U5336 (N_5336,In_2652,In_2037);
nor U5337 (N_5337,In_2025,In_537);
or U5338 (N_5338,In_1658,In_2151);
xor U5339 (N_5339,In_1385,In_2885);
xnor U5340 (N_5340,In_1324,In_2493);
nor U5341 (N_5341,In_2397,In_1539);
nor U5342 (N_5342,In_2568,In_2962);
nor U5343 (N_5343,In_1552,In_2316);
nand U5344 (N_5344,In_2483,In_1977);
nand U5345 (N_5345,In_1065,In_1791);
nand U5346 (N_5346,In_2563,In_599);
or U5347 (N_5347,In_2231,In_223);
xor U5348 (N_5348,In_77,In_107);
or U5349 (N_5349,In_531,In_1607);
or U5350 (N_5350,In_1737,In_1347);
or U5351 (N_5351,In_793,In_735);
nand U5352 (N_5352,In_1339,In_2745);
nand U5353 (N_5353,In_1072,In_1680);
nand U5354 (N_5354,In_599,In_2488);
and U5355 (N_5355,In_896,In_1478);
or U5356 (N_5356,In_1683,In_2873);
nand U5357 (N_5357,In_1119,In_81);
or U5358 (N_5358,In_2275,In_1084);
or U5359 (N_5359,In_2600,In_697);
and U5360 (N_5360,In_1352,In_2439);
nand U5361 (N_5361,In_815,In_2149);
or U5362 (N_5362,In_291,In_433);
nor U5363 (N_5363,In_225,In_657);
nand U5364 (N_5364,In_823,In_2538);
nor U5365 (N_5365,In_1581,In_1209);
or U5366 (N_5366,In_184,In_162);
or U5367 (N_5367,In_810,In_791);
and U5368 (N_5368,In_2629,In_302);
nand U5369 (N_5369,In_586,In_1418);
or U5370 (N_5370,In_853,In_1334);
and U5371 (N_5371,In_78,In_2790);
nand U5372 (N_5372,In_1068,In_1779);
and U5373 (N_5373,In_2366,In_944);
xor U5374 (N_5374,In_2810,In_327);
nor U5375 (N_5375,In_2881,In_1959);
and U5376 (N_5376,In_1302,In_2625);
or U5377 (N_5377,In_2103,In_1137);
or U5378 (N_5378,In_2146,In_458);
nand U5379 (N_5379,In_2033,In_1307);
nor U5380 (N_5380,In_1487,In_1725);
and U5381 (N_5381,In_1241,In_1311);
and U5382 (N_5382,In_2369,In_959);
nor U5383 (N_5383,In_1054,In_2478);
nand U5384 (N_5384,In_1186,In_1360);
xor U5385 (N_5385,In_1264,In_1901);
and U5386 (N_5386,In_724,In_1888);
and U5387 (N_5387,In_335,In_2961);
nand U5388 (N_5388,In_982,In_19);
and U5389 (N_5389,In_600,In_889);
or U5390 (N_5390,In_196,In_412);
nand U5391 (N_5391,In_785,In_376);
nor U5392 (N_5392,In_1995,In_2082);
nor U5393 (N_5393,In_2939,In_330);
nand U5394 (N_5394,In_1629,In_1479);
nor U5395 (N_5395,In_487,In_1123);
or U5396 (N_5396,In_66,In_1269);
and U5397 (N_5397,In_286,In_2452);
or U5398 (N_5398,In_1777,In_2387);
and U5399 (N_5399,In_1346,In_2909);
and U5400 (N_5400,In_1223,In_1091);
xnor U5401 (N_5401,In_1878,In_574);
nand U5402 (N_5402,In_13,In_350);
and U5403 (N_5403,In_188,In_84);
or U5404 (N_5404,In_1735,In_1338);
or U5405 (N_5405,In_2028,In_1545);
or U5406 (N_5406,In_1055,In_430);
or U5407 (N_5407,In_43,In_2980);
and U5408 (N_5408,In_1064,In_2152);
nor U5409 (N_5409,In_2718,In_256);
or U5410 (N_5410,In_1011,In_1429);
xor U5411 (N_5411,In_255,In_973);
nor U5412 (N_5412,In_1844,In_1362);
nor U5413 (N_5413,In_270,In_199);
or U5414 (N_5414,In_1036,In_2396);
and U5415 (N_5415,In_1825,In_1953);
nand U5416 (N_5416,In_2263,In_1649);
or U5417 (N_5417,In_1465,In_1798);
nor U5418 (N_5418,In_2411,In_46);
and U5419 (N_5419,In_578,In_1159);
or U5420 (N_5420,In_2206,In_11);
or U5421 (N_5421,In_2507,In_455);
nor U5422 (N_5422,In_2323,In_2879);
and U5423 (N_5423,In_2806,In_782);
xor U5424 (N_5424,In_443,In_1890);
nand U5425 (N_5425,In_1317,In_1163);
or U5426 (N_5426,In_2404,In_1129);
and U5427 (N_5427,In_2447,In_1986);
xor U5428 (N_5428,In_442,In_2821);
nand U5429 (N_5429,In_2385,In_2831);
nand U5430 (N_5430,In_667,In_291);
nand U5431 (N_5431,In_241,In_875);
or U5432 (N_5432,In_1515,In_440);
or U5433 (N_5433,In_2993,In_1886);
nor U5434 (N_5434,In_657,In_1543);
nor U5435 (N_5435,In_2292,In_698);
xor U5436 (N_5436,In_1387,In_1957);
or U5437 (N_5437,In_442,In_2920);
or U5438 (N_5438,In_2205,In_1616);
nand U5439 (N_5439,In_2955,In_42);
or U5440 (N_5440,In_1055,In_937);
or U5441 (N_5441,In_467,In_289);
or U5442 (N_5442,In_2057,In_2486);
or U5443 (N_5443,In_2129,In_2583);
nand U5444 (N_5444,In_123,In_2655);
nor U5445 (N_5445,In_1986,In_1263);
and U5446 (N_5446,In_679,In_1537);
nand U5447 (N_5447,In_1166,In_458);
nand U5448 (N_5448,In_747,In_1088);
nand U5449 (N_5449,In_1435,In_233);
or U5450 (N_5450,In_58,In_1982);
xor U5451 (N_5451,In_2806,In_1849);
and U5452 (N_5452,In_629,In_1643);
nand U5453 (N_5453,In_485,In_388);
nor U5454 (N_5454,In_450,In_798);
xnor U5455 (N_5455,In_2004,In_1688);
and U5456 (N_5456,In_815,In_2195);
nand U5457 (N_5457,In_202,In_107);
or U5458 (N_5458,In_489,In_1724);
and U5459 (N_5459,In_2398,In_1942);
and U5460 (N_5460,In_1520,In_2550);
nor U5461 (N_5461,In_1249,In_1305);
or U5462 (N_5462,In_1796,In_1739);
xor U5463 (N_5463,In_320,In_2136);
nor U5464 (N_5464,In_2970,In_1421);
nor U5465 (N_5465,In_911,In_2830);
and U5466 (N_5466,In_2528,In_2642);
nand U5467 (N_5467,In_2254,In_1377);
nor U5468 (N_5468,In_1601,In_2571);
or U5469 (N_5469,In_2954,In_112);
xnor U5470 (N_5470,In_1663,In_1262);
xor U5471 (N_5471,In_160,In_1386);
or U5472 (N_5472,In_1528,In_2309);
nand U5473 (N_5473,In_2305,In_448);
or U5474 (N_5474,In_2903,In_960);
xnor U5475 (N_5475,In_1606,In_713);
and U5476 (N_5476,In_1413,In_75);
nand U5477 (N_5477,In_2547,In_2);
xnor U5478 (N_5478,In_1935,In_459);
and U5479 (N_5479,In_23,In_726);
xnor U5480 (N_5480,In_2149,In_1009);
and U5481 (N_5481,In_193,In_2014);
nand U5482 (N_5482,In_76,In_2481);
and U5483 (N_5483,In_335,In_2282);
and U5484 (N_5484,In_1943,In_1845);
or U5485 (N_5485,In_2736,In_523);
xor U5486 (N_5486,In_324,In_1631);
or U5487 (N_5487,In_2351,In_2596);
xnor U5488 (N_5488,In_2053,In_95);
or U5489 (N_5489,In_2698,In_477);
nand U5490 (N_5490,In_2429,In_1920);
nand U5491 (N_5491,In_2748,In_2105);
or U5492 (N_5492,In_2604,In_286);
or U5493 (N_5493,In_619,In_1101);
nor U5494 (N_5494,In_416,In_1987);
and U5495 (N_5495,In_266,In_1220);
or U5496 (N_5496,In_1159,In_566);
and U5497 (N_5497,In_302,In_2415);
and U5498 (N_5498,In_2192,In_590);
or U5499 (N_5499,In_1669,In_1408);
xor U5500 (N_5500,In_1863,In_2046);
xor U5501 (N_5501,In_2252,In_1575);
and U5502 (N_5502,In_594,In_1793);
nor U5503 (N_5503,In_1643,In_1946);
and U5504 (N_5504,In_2231,In_1007);
nor U5505 (N_5505,In_1164,In_334);
xor U5506 (N_5506,In_608,In_854);
xor U5507 (N_5507,In_1785,In_1836);
nand U5508 (N_5508,In_2553,In_2386);
and U5509 (N_5509,In_1297,In_100);
nand U5510 (N_5510,In_146,In_2694);
nand U5511 (N_5511,In_2942,In_276);
nand U5512 (N_5512,In_1515,In_1208);
or U5513 (N_5513,In_1043,In_2985);
xnor U5514 (N_5514,In_2511,In_133);
nor U5515 (N_5515,In_1122,In_2970);
or U5516 (N_5516,In_2572,In_2565);
nand U5517 (N_5517,In_1878,In_1569);
nand U5518 (N_5518,In_850,In_1324);
xnor U5519 (N_5519,In_1529,In_2272);
nand U5520 (N_5520,In_2095,In_2691);
and U5521 (N_5521,In_1346,In_1019);
nand U5522 (N_5522,In_868,In_475);
and U5523 (N_5523,In_1457,In_144);
nand U5524 (N_5524,In_1440,In_1753);
or U5525 (N_5525,In_1592,In_1414);
nor U5526 (N_5526,In_2136,In_1873);
and U5527 (N_5527,In_210,In_2990);
nand U5528 (N_5528,In_2072,In_2330);
and U5529 (N_5529,In_2345,In_381);
and U5530 (N_5530,In_1895,In_184);
nand U5531 (N_5531,In_2640,In_2044);
nor U5532 (N_5532,In_1226,In_147);
and U5533 (N_5533,In_810,In_1234);
and U5534 (N_5534,In_1612,In_371);
nand U5535 (N_5535,In_843,In_2785);
nand U5536 (N_5536,In_282,In_2056);
or U5537 (N_5537,In_1354,In_254);
and U5538 (N_5538,In_2417,In_2027);
nand U5539 (N_5539,In_2294,In_428);
xnor U5540 (N_5540,In_1396,In_24);
nand U5541 (N_5541,In_806,In_758);
nor U5542 (N_5542,In_2925,In_332);
or U5543 (N_5543,In_1113,In_1277);
and U5544 (N_5544,In_1966,In_2991);
and U5545 (N_5545,In_1406,In_376);
or U5546 (N_5546,In_2004,In_1102);
xor U5547 (N_5547,In_2731,In_2083);
nor U5548 (N_5548,In_1986,In_1922);
nand U5549 (N_5549,In_869,In_473);
or U5550 (N_5550,In_2361,In_910);
or U5551 (N_5551,In_39,In_2675);
and U5552 (N_5552,In_2317,In_1107);
and U5553 (N_5553,In_1837,In_640);
and U5554 (N_5554,In_49,In_230);
nor U5555 (N_5555,In_615,In_2590);
nor U5556 (N_5556,In_2015,In_1558);
or U5557 (N_5557,In_779,In_2160);
nor U5558 (N_5558,In_2928,In_1610);
or U5559 (N_5559,In_351,In_937);
nand U5560 (N_5560,In_609,In_1016);
xor U5561 (N_5561,In_2079,In_2827);
or U5562 (N_5562,In_2679,In_2396);
nand U5563 (N_5563,In_2678,In_620);
xnor U5564 (N_5564,In_1642,In_2305);
and U5565 (N_5565,In_1635,In_745);
and U5566 (N_5566,In_552,In_2941);
nor U5567 (N_5567,In_2811,In_2669);
xor U5568 (N_5568,In_130,In_1496);
nor U5569 (N_5569,In_2684,In_1904);
nand U5570 (N_5570,In_773,In_1297);
nor U5571 (N_5571,In_1768,In_1153);
nor U5572 (N_5572,In_1565,In_2333);
and U5573 (N_5573,In_2809,In_2789);
or U5574 (N_5574,In_2147,In_1908);
nand U5575 (N_5575,In_2408,In_1706);
nor U5576 (N_5576,In_1457,In_1376);
nand U5577 (N_5577,In_2499,In_1394);
and U5578 (N_5578,In_2874,In_1366);
xor U5579 (N_5579,In_929,In_1598);
xnor U5580 (N_5580,In_1136,In_191);
nor U5581 (N_5581,In_2239,In_2749);
xor U5582 (N_5582,In_2522,In_2017);
nor U5583 (N_5583,In_81,In_348);
xor U5584 (N_5584,In_2412,In_2247);
xnor U5585 (N_5585,In_845,In_990);
or U5586 (N_5586,In_1139,In_2419);
or U5587 (N_5587,In_444,In_2581);
nor U5588 (N_5588,In_422,In_1334);
xnor U5589 (N_5589,In_951,In_1183);
nand U5590 (N_5590,In_1300,In_22);
and U5591 (N_5591,In_2528,In_2220);
nand U5592 (N_5592,In_203,In_1701);
nor U5593 (N_5593,In_2708,In_686);
and U5594 (N_5594,In_2254,In_352);
xor U5595 (N_5595,In_1506,In_2287);
or U5596 (N_5596,In_2686,In_2366);
nand U5597 (N_5597,In_17,In_1753);
or U5598 (N_5598,In_753,In_2822);
xor U5599 (N_5599,In_2574,In_1811);
xor U5600 (N_5600,In_1350,In_2195);
nor U5601 (N_5601,In_2049,In_2899);
or U5602 (N_5602,In_519,In_45);
or U5603 (N_5603,In_609,In_495);
xnor U5604 (N_5604,In_2146,In_2202);
xnor U5605 (N_5605,In_133,In_40);
nor U5606 (N_5606,In_2891,In_1776);
or U5607 (N_5607,In_2419,In_1121);
nand U5608 (N_5608,In_2997,In_1106);
nor U5609 (N_5609,In_1685,In_147);
and U5610 (N_5610,In_933,In_2380);
nor U5611 (N_5611,In_1639,In_275);
xnor U5612 (N_5612,In_1349,In_1964);
and U5613 (N_5613,In_1810,In_531);
nor U5614 (N_5614,In_1271,In_1176);
xor U5615 (N_5615,In_2796,In_1004);
and U5616 (N_5616,In_2339,In_385);
nor U5617 (N_5617,In_1213,In_2117);
and U5618 (N_5618,In_543,In_553);
xnor U5619 (N_5619,In_579,In_364);
and U5620 (N_5620,In_762,In_421);
nand U5621 (N_5621,In_1906,In_2032);
nor U5622 (N_5622,In_2897,In_2327);
nand U5623 (N_5623,In_2704,In_1094);
nor U5624 (N_5624,In_2092,In_121);
and U5625 (N_5625,In_2939,In_1212);
xor U5626 (N_5626,In_2457,In_1221);
or U5627 (N_5627,In_918,In_2977);
nor U5628 (N_5628,In_2397,In_1814);
and U5629 (N_5629,In_2372,In_273);
nand U5630 (N_5630,In_205,In_1447);
and U5631 (N_5631,In_2988,In_129);
or U5632 (N_5632,In_1957,In_962);
xnor U5633 (N_5633,In_2754,In_1146);
and U5634 (N_5634,In_2928,In_1153);
or U5635 (N_5635,In_2597,In_118);
nand U5636 (N_5636,In_1413,In_1605);
and U5637 (N_5637,In_2854,In_86);
nand U5638 (N_5638,In_1536,In_1695);
nand U5639 (N_5639,In_1088,In_2998);
nand U5640 (N_5640,In_973,In_2940);
nand U5641 (N_5641,In_1256,In_2523);
xor U5642 (N_5642,In_2597,In_2878);
nand U5643 (N_5643,In_1789,In_1988);
nor U5644 (N_5644,In_1171,In_2825);
or U5645 (N_5645,In_2182,In_2660);
or U5646 (N_5646,In_542,In_2470);
or U5647 (N_5647,In_2134,In_1431);
or U5648 (N_5648,In_2092,In_2280);
and U5649 (N_5649,In_1331,In_891);
nand U5650 (N_5650,In_1512,In_1114);
nand U5651 (N_5651,In_1409,In_57);
nand U5652 (N_5652,In_389,In_1050);
and U5653 (N_5653,In_2300,In_1818);
xnor U5654 (N_5654,In_1443,In_1604);
nor U5655 (N_5655,In_2367,In_797);
nand U5656 (N_5656,In_2175,In_421);
xor U5657 (N_5657,In_1457,In_2321);
nor U5658 (N_5658,In_29,In_2133);
or U5659 (N_5659,In_1695,In_776);
xor U5660 (N_5660,In_1458,In_37);
nand U5661 (N_5661,In_1816,In_642);
nand U5662 (N_5662,In_165,In_2633);
and U5663 (N_5663,In_342,In_2229);
nor U5664 (N_5664,In_2373,In_664);
xnor U5665 (N_5665,In_1904,In_2190);
or U5666 (N_5666,In_1398,In_2309);
nand U5667 (N_5667,In_1860,In_976);
nor U5668 (N_5668,In_752,In_294);
and U5669 (N_5669,In_287,In_109);
xor U5670 (N_5670,In_1341,In_609);
and U5671 (N_5671,In_967,In_1340);
xnor U5672 (N_5672,In_260,In_124);
nor U5673 (N_5673,In_1597,In_2499);
nor U5674 (N_5674,In_421,In_298);
or U5675 (N_5675,In_824,In_546);
nand U5676 (N_5676,In_813,In_509);
nand U5677 (N_5677,In_2178,In_1584);
and U5678 (N_5678,In_153,In_2539);
and U5679 (N_5679,In_2750,In_509);
xor U5680 (N_5680,In_1746,In_733);
and U5681 (N_5681,In_1057,In_2004);
nand U5682 (N_5682,In_1720,In_551);
and U5683 (N_5683,In_1436,In_960);
or U5684 (N_5684,In_2268,In_1890);
xnor U5685 (N_5685,In_1482,In_1612);
nand U5686 (N_5686,In_2342,In_1485);
nand U5687 (N_5687,In_135,In_162);
nand U5688 (N_5688,In_402,In_2196);
xor U5689 (N_5689,In_1121,In_1133);
or U5690 (N_5690,In_754,In_1361);
xor U5691 (N_5691,In_2988,In_2922);
nor U5692 (N_5692,In_2329,In_1816);
or U5693 (N_5693,In_2146,In_126);
or U5694 (N_5694,In_2035,In_1052);
nor U5695 (N_5695,In_2264,In_2577);
xor U5696 (N_5696,In_939,In_944);
or U5697 (N_5697,In_108,In_2569);
nand U5698 (N_5698,In_1044,In_2882);
and U5699 (N_5699,In_389,In_1380);
xor U5700 (N_5700,In_1568,In_2222);
nand U5701 (N_5701,In_1045,In_549);
nand U5702 (N_5702,In_2860,In_2039);
or U5703 (N_5703,In_1903,In_1930);
nand U5704 (N_5704,In_2436,In_163);
or U5705 (N_5705,In_2880,In_130);
or U5706 (N_5706,In_155,In_2065);
and U5707 (N_5707,In_2581,In_1438);
xnor U5708 (N_5708,In_1283,In_53);
nor U5709 (N_5709,In_1959,In_1061);
nor U5710 (N_5710,In_1586,In_1757);
xor U5711 (N_5711,In_997,In_1068);
xnor U5712 (N_5712,In_582,In_723);
nand U5713 (N_5713,In_105,In_476);
nor U5714 (N_5714,In_2479,In_327);
nand U5715 (N_5715,In_1504,In_2099);
xnor U5716 (N_5716,In_869,In_341);
nand U5717 (N_5717,In_1626,In_30);
nor U5718 (N_5718,In_2733,In_849);
nor U5719 (N_5719,In_458,In_1300);
or U5720 (N_5720,In_702,In_2121);
nand U5721 (N_5721,In_2838,In_864);
xor U5722 (N_5722,In_134,In_790);
and U5723 (N_5723,In_1318,In_2251);
nor U5724 (N_5724,In_2399,In_345);
and U5725 (N_5725,In_2744,In_102);
and U5726 (N_5726,In_1064,In_1013);
nor U5727 (N_5727,In_1489,In_2173);
and U5728 (N_5728,In_413,In_1879);
or U5729 (N_5729,In_101,In_683);
xor U5730 (N_5730,In_2145,In_319);
nand U5731 (N_5731,In_330,In_649);
nor U5732 (N_5732,In_1986,In_2260);
xor U5733 (N_5733,In_1877,In_1824);
or U5734 (N_5734,In_820,In_2954);
nor U5735 (N_5735,In_388,In_1802);
nand U5736 (N_5736,In_980,In_1696);
or U5737 (N_5737,In_2990,In_2749);
or U5738 (N_5738,In_1238,In_143);
and U5739 (N_5739,In_1297,In_1231);
xor U5740 (N_5740,In_742,In_2602);
or U5741 (N_5741,In_605,In_926);
nor U5742 (N_5742,In_2707,In_903);
or U5743 (N_5743,In_499,In_2141);
nand U5744 (N_5744,In_2411,In_1040);
and U5745 (N_5745,In_2301,In_340);
xnor U5746 (N_5746,In_1625,In_253);
or U5747 (N_5747,In_757,In_2106);
or U5748 (N_5748,In_2938,In_1304);
xnor U5749 (N_5749,In_1130,In_2141);
nand U5750 (N_5750,In_762,In_163);
xor U5751 (N_5751,In_1327,In_161);
xnor U5752 (N_5752,In_1030,In_2337);
or U5753 (N_5753,In_1989,In_802);
or U5754 (N_5754,In_2584,In_125);
and U5755 (N_5755,In_786,In_2805);
nor U5756 (N_5756,In_2297,In_367);
nor U5757 (N_5757,In_1857,In_1248);
or U5758 (N_5758,In_397,In_2116);
nand U5759 (N_5759,In_2192,In_2538);
xnor U5760 (N_5760,In_2653,In_594);
xnor U5761 (N_5761,In_1780,In_661);
xnor U5762 (N_5762,In_2315,In_2633);
nand U5763 (N_5763,In_1548,In_183);
xor U5764 (N_5764,In_1421,In_2632);
nor U5765 (N_5765,In_213,In_2490);
nor U5766 (N_5766,In_1768,In_1920);
or U5767 (N_5767,In_1795,In_1062);
xnor U5768 (N_5768,In_1518,In_1972);
xor U5769 (N_5769,In_1853,In_1578);
or U5770 (N_5770,In_2776,In_1260);
xor U5771 (N_5771,In_2344,In_2123);
or U5772 (N_5772,In_2236,In_1120);
nand U5773 (N_5773,In_421,In_996);
nor U5774 (N_5774,In_868,In_2821);
xor U5775 (N_5775,In_467,In_978);
and U5776 (N_5776,In_1708,In_2750);
xor U5777 (N_5777,In_1246,In_1704);
xor U5778 (N_5778,In_148,In_226);
or U5779 (N_5779,In_1938,In_2013);
or U5780 (N_5780,In_1690,In_1303);
and U5781 (N_5781,In_1312,In_45);
xor U5782 (N_5782,In_1895,In_1609);
or U5783 (N_5783,In_884,In_825);
nor U5784 (N_5784,In_1388,In_2503);
xnor U5785 (N_5785,In_624,In_2172);
nor U5786 (N_5786,In_1376,In_656);
nand U5787 (N_5787,In_1063,In_1046);
xor U5788 (N_5788,In_2800,In_394);
and U5789 (N_5789,In_936,In_1458);
nand U5790 (N_5790,In_1055,In_1994);
nor U5791 (N_5791,In_793,In_2659);
and U5792 (N_5792,In_248,In_2070);
nand U5793 (N_5793,In_1970,In_1649);
or U5794 (N_5794,In_2091,In_2648);
and U5795 (N_5795,In_1398,In_573);
and U5796 (N_5796,In_2252,In_1473);
and U5797 (N_5797,In_445,In_2580);
nand U5798 (N_5798,In_1818,In_1655);
nand U5799 (N_5799,In_2009,In_833);
nor U5800 (N_5800,In_2768,In_1607);
nand U5801 (N_5801,In_867,In_2952);
nor U5802 (N_5802,In_647,In_473);
nand U5803 (N_5803,In_540,In_691);
and U5804 (N_5804,In_1887,In_417);
and U5805 (N_5805,In_82,In_1574);
nor U5806 (N_5806,In_346,In_1273);
nand U5807 (N_5807,In_555,In_2827);
xnor U5808 (N_5808,In_799,In_1823);
or U5809 (N_5809,In_2908,In_888);
xor U5810 (N_5810,In_774,In_338);
or U5811 (N_5811,In_28,In_2590);
nand U5812 (N_5812,In_91,In_395);
or U5813 (N_5813,In_2909,In_697);
xor U5814 (N_5814,In_59,In_1341);
nor U5815 (N_5815,In_1638,In_2258);
xnor U5816 (N_5816,In_259,In_2491);
nor U5817 (N_5817,In_1067,In_1170);
nand U5818 (N_5818,In_1146,In_570);
xor U5819 (N_5819,In_1288,In_2977);
or U5820 (N_5820,In_835,In_2534);
nand U5821 (N_5821,In_1370,In_1387);
or U5822 (N_5822,In_308,In_1537);
xnor U5823 (N_5823,In_1877,In_1057);
or U5824 (N_5824,In_670,In_712);
xor U5825 (N_5825,In_2429,In_2909);
and U5826 (N_5826,In_1599,In_935);
xnor U5827 (N_5827,In_2122,In_1404);
nand U5828 (N_5828,In_1256,In_706);
or U5829 (N_5829,In_1936,In_741);
and U5830 (N_5830,In_1000,In_1407);
nor U5831 (N_5831,In_410,In_2601);
xor U5832 (N_5832,In_2413,In_1215);
nand U5833 (N_5833,In_2980,In_773);
xor U5834 (N_5834,In_467,In_2844);
nand U5835 (N_5835,In_2890,In_2102);
or U5836 (N_5836,In_2098,In_172);
xor U5837 (N_5837,In_2631,In_349);
xnor U5838 (N_5838,In_1064,In_1722);
or U5839 (N_5839,In_1194,In_1411);
nor U5840 (N_5840,In_2358,In_644);
xnor U5841 (N_5841,In_113,In_546);
xor U5842 (N_5842,In_1215,In_2410);
xnor U5843 (N_5843,In_1104,In_2532);
or U5844 (N_5844,In_2203,In_886);
nand U5845 (N_5845,In_803,In_2460);
and U5846 (N_5846,In_1570,In_852);
nand U5847 (N_5847,In_1402,In_1062);
and U5848 (N_5848,In_154,In_92);
nor U5849 (N_5849,In_627,In_695);
nand U5850 (N_5850,In_1872,In_1326);
nand U5851 (N_5851,In_2743,In_414);
nor U5852 (N_5852,In_2991,In_517);
nor U5853 (N_5853,In_2185,In_306);
or U5854 (N_5854,In_991,In_778);
nor U5855 (N_5855,In_2289,In_651);
nand U5856 (N_5856,In_542,In_1187);
nor U5857 (N_5857,In_1323,In_1862);
xnor U5858 (N_5858,In_1441,In_2020);
xor U5859 (N_5859,In_1025,In_627);
nand U5860 (N_5860,In_2525,In_2087);
and U5861 (N_5861,In_1577,In_1776);
and U5862 (N_5862,In_1251,In_1886);
nand U5863 (N_5863,In_1902,In_2109);
nand U5864 (N_5864,In_1266,In_2891);
or U5865 (N_5865,In_2828,In_231);
or U5866 (N_5866,In_1861,In_1433);
and U5867 (N_5867,In_1859,In_2427);
nand U5868 (N_5868,In_1373,In_2893);
and U5869 (N_5869,In_600,In_66);
nand U5870 (N_5870,In_2734,In_443);
and U5871 (N_5871,In_1272,In_2267);
nand U5872 (N_5872,In_1186,In_1697);
nand U5873 (N_5873,In_2701,In_1932);
or U5874 (N_5874,In_1428,In_223);
xor U5875 (N_5875,In_1805,In_1930);
and U5876 (N_5876,In_2143,In_1109);
and U5877 (N_5877,In_2233,In_232);
xor U5878 (N_5878,In_653,In_18);
and U5879 (N_5879,In_1928,In_2274);
nand U5880 (N_5880,In_246,In_1746);
and U5881 (N_5881,In_2657,In_543);
and U5882 (N_5882,In_975,In_136);
nor U5883 (N_5883,In_2761,In_881);
and U5884 (N_5884,In_2886,In_2487);
nor U5885 (N_5885,In_226,In_906);
and U5886 (N_5886,In_1843,In_1840);
or U5887 (N_5887,In_340,In_1407);
nand U5888 (N_5888,In_979,In_46);
nor U5889 (N_5889,In_747,In_2129);
xor U5890 (N_5890,In_1431,In_41);
or U5891 (N_5891,In_1711,In_2691);
or U5892 (N_5892,In_1024,In_1819);
and U5893 (N_5893,In_2830,In_1545);
and U5894 (N_5894,In_1620,In_2117);
and U5895 (N_5895,In_169,In_2453);
nor U5896 (N_5896,In_2621,In_2098);
and U5897 (N_5897,In_1412,In_2701);
xor U5898 (N_5898,In_1660,In_2944);
and U5899 (N_5899,In_1725,In_2566);
xnor U5900 (N_5900,In_1687,In_2100);
nand U5901 (N_5901,In_982,In_67);
and U5902 (N_5902,In_2119,In_739);
xnor U5903 (N_5903,In_438,In_1875);
nand U5904 (N_5904,In_2907,In_930);
xnor U5905 (N_5905,In_1286,In_1441);
nor U5906 (N_5906,In_2325,In_1088);
or U5907 (N_5907,In_958,In_1411);
or U5908 (N_5908,In_2573,In_1306);
or U5909 (N_5909,In_152,In_451);
xor U5910 (N_5910,In_2621,In_722);
nor U5911 (N_5911,In_419,In_418);
or U5912 (N_5912,In_903,In_542);
xnor U5913 (N_5913,In_1719,In_1813);
nand U5914 (N_5914,In_2844,In_1120);
nor U5915 (N_5915,In_1402,In_1846);
nor U5916 (N_5916,In_2850,In_2040);
or U5917 (N_5917,In_84,In_119);
nor U5918 (N_5918,In_397,In_1103);
or U5919 (N_5919,In_1010,In_2172);
and U5920 (N_5920,In_190,In_1118);
nand U5921 (N_5921,In_310,In_2034);
xnor U5922 (N_5922,In_851,In_1178);
or U5923 (N_5923,In_2177,In_1625);
and U5924 (N_5924,In_1700,In_1046);
or U5925 (N_5925,In_1467,In_2947);
xor U5926 (N_5926,In_2076,In_111);
nor U5927 (N_5927,In_1831,In_1653);
xnor U5928 (N_5928,In_2094,In_1561);
nor U5929 (N_5929,In_284,In_1152);
and U5930 (N_5930,In_2332,In_990);
nor U5931 (N_5931,In_268,In_900);
xor U5932 (N_5932,In_2384,In_1193);
and U5933 (N_5933,In_1585,In_889);
or U5934 (N_5934,In_2357,In_1615);
nand U5935 (N_5935,In_710,In_2318);
nor U5936 (N_5936,In_1516,In_1602);
xor U5937 (N_5937,In_2646,In_2445);
nand U5938 (N_5938,In_208,In_1424);
and U5939 (N_5939,In_2520,In_758);
xor U5940 (N_5940,In_51,In_2412);
xor U5941 (N_5941,In_1249,In_1748);
nand U5942 (N_5942,In_2230,In_311);
nor U5943 (N_5943,In_2800,In_2490);
nor U5944 (N_5944,In_2933,In_2497);
or U5945 (N_5945,In_2092,In_994);
and U5946 (N_5946,In_2951,In_1584);
and U5947 (N_5947,In_375,In_192);
or U5948 (N_5948,In_2517,In_2798);
xnor U5949 (N_5949,In_271,In_1785);
nor U5950 (N_5950,In_2440,In_742);
or U5951 (N_5951,In_2154,In_1677);
and U5952 (N_5952,In_571,In_248);
and U5953 (N_5953,In_2146,In_2820);
nor U5954 (N_5954,In_1630,In_361);
xnor U5955 (N_5955,In_1382,In_2093);
or U5956 (N_5956,In_2970,In_1552);
and U5957 (N_5957,In_1126,In_2983);
nor U5958 (N_5958,In_2637,In_739);
nand U5959 (N_5959,In_2941,In_785);
nor U5960 (N_5960,In_1550,In_2571);
and U5961 (N_5961,In_1398,In_2797);
nand U5962 (N_5962,In_1059,In_2239);
nand U5963 (N_5963,In_2836,In_1246);
xor U5964 (N_5964,In_1614,In_199);
xnor U5965 (N_5965,In_1823,In_1352);
and U5966 (N_5966,In_2441,In_1634);
nand U5967 (N_5967,In_2777,In_906);
and U5968 (N_5968,In_128,In_604);
nand U5969 (N_5969,In_2255,In_1386);
or U5970 (N_5970,In_1135,In_2554);
and U5971 (N_5971,In_2534,In_1920);
xnor U5972 (N_5972,In_1781,In_2167);
nand U5973 (N_5973,In_1313,In_2738);
nor U5974 (N_5974,In_385,In_137);
nand U5975 (N_5975,In_623,In_2786);
nand U5976 (N_5976,In_2859,In_515);
or U5977 (N_5977,In_1961,In_2865);
nand U5978 (N_5978,In_2602,In_2850);
or U5979 (N_5979,In_736,In_2376);
nand U5980 (N_5980,In_1935,In_2597);
xnor U5981 (N_5981,In_843,In_708);
nor U5982 (N_5982,In_186,In_328);
or U5983 (N_5983,In_435,In_555);
or U5984 (N_5984,In_750,In_1480);
xor U5985 (N_5985,In_530,In_787);
or U5986 (N_5986,In_1642,In_2519);
and U5987 (N_5987,In_1615,In_1164);
nand U5988 (N_5988,In_980,In_2981);
and U5989 (N_5989,In_1691,In_1099);
and U5990 (N_5990,In_1349,In_2922);
xor U5991 (N_5991,In_2331,In_1980);
nand U5992 (N_5992,In_94,In_1466);
nor U5993 (N_5993,In_2695,In_1894);
nand U5994 (N_5994,In_2220,In_957);
or U5995 (N_5995,In_2592,In_1389);
xor U5996 (N_5996,In_746,In_1967);
or U5997 (N_5997,In_2345,In_2050);
nand U5998 (N_5998,In_95,In_1926);
xor U5999 (N_5999,In_1265,In_286);
nand U6000 (N_6000,N_75,N_2956);
and U6001 (N_6001,N_2376,N_4974);
xnor U6002 (N_6002,N_1631,N_2096);
or U6003 (N_6003,N_3912,N_5267);
and U6004 (N_6004,N_4638,N_162);
and U6005 (N_6005,N_5473,N_671);
or U6006 (N_6006,N_3900,N_637);
nor U6007 (N_6007,N_2188,N_1825);
xor U6008 (N_6008,N_5263,N_232);
or U6009 (N_6009,N_1413,N_1209);
nand U6010 (N_6010,N_3632,N_5002);
nor U6011 (N_6011,N_2467,N_1777);
xnor U6012 (N_6012,N_1228,N_73);
xor U6013 (N_6013,N_2700,N_1215);
nand U6014 (N_6014,N_4990,N_4634);
and U6015 (N_6015,N_5174,N_93);
nor U6016 (N_6016,N_5551,N_5776);
nor U6017 (N_6017,N_4439,N_5412);
and U6018 (N_6018,N_5980,N_4779);
xnor U6019 (N_6019,N_1294,N_2248);
nor U6020 (N_6020,N_5246,N_3621);
xnor U6021 (N_6021,N_1977,N_1478);
and U6022 (N_6022,N_5569,N_5889);
and U6023 (N_6023,N_1578,N_3490);
nor U6024 (N_6024,N_3322,N_1856);
and U6025 (N_6025,N_4329,N_4695);
nand U6026 (N_6026,N_5760,N_2309);
xnor U6027 (N_6027,N_439,N_1296);
nand U6028 (N_6028,N_137,N_5527);
nand U6029 (N_6029,N_5710,N_5395);
xor U6030 (N_6030,N_5753,N_5008);
nand U6031 (N_6031,N_4840,N_2354);
nand U6032 (N_6032,N_3595,N_4622);
nand U6033 (N_6033,N_5319,N_1256);
xnor U6034 (N_6034,N_2415,N_5368);
or U6035 (N_6035,N_1269,N_4501);
nand U6036 (N_6036,N_1684,N_5846);
or U6037 (N_6037,N_355,N_451);
xor U6038 (N_6038,N_1210,N_1696);
and U6039 (N_6039,N_3399,N_5700);
nand U6040 (N_6040,N_3010,N_4631);
nor U6041 (N_6041,N_1423,N_2298);
or U6042 (N_6042,N_5391,N_4288);
nor U6043 (N_6043,N_2689,N_2133);
and U6044 (N_6044,N_2773,N_793);
and U6045 (N_6045,N_5245,N_1634);
and U6046 (N_6046,N_4188,N_3069);
nor U6047 (N_6047,N_4552,N_5287);
or U6048 (N_6048,N_1870,N_5484);
nor U6049 (N_6049,N_362,N_836);
nor U6050 (N_6050,N_672,N_3519);
xor U6051 (N_6051,N_5979,N_4221);
nand U6052 (N_6052,N_1197,N_3169);
xor U6053 (N_6053,N_3601,N_4740);
nor U6054 (N_6054,N_3123,N_4906);
xnor U6055 (N_6055,N_5497,N_1276);
or U6056 (N_6056,N_2134,N_771);
nand U6057 (N_6057,N_1953,N_558);
nor U6058 (N_6058,N_2375,N_859);
and U6059 (N_6059,N_1122,N_201);
nor U6060 (N_6060,N_3866,N_3369);
xnor U6061 (N_6061,N_995,N_5148);
xnor U6062 (N_6062,N_4332,N_5370);
nand U6063 (N_6063,N_5439,N_2783);
or U6064 (N_6064,N_2486,N_1657);
or U6065 (N_6065,N_1848,N_4294);
or U6066 (N_6066,N_5805,N_1692);
nand U6067 (N_6067,N_2110,N_5378);
nor U6068 (N_6068,N_833,N_1568);
xor U6069 (N_6069,N_516,N_5790);
xnor U6070 (N_6070,N_4451,N_2211);
or U6071 (N_6071,N_3861,N_3032);
and U6072 (N_6072,N_208,N_2328);
xor U6073 (N_6073,N_3363,N_4937);
and U6074 (N_6074,N_1698,N_2823);
nand U6075 (N_6075,N_938,N_329);
xnor U6076 (N_6076,N_2901,N_2348);
and U6077 (N_6077,N_97,N_1690);
and U6078 (N_6078,N_2013,N_102);
and U6079 (N_6079,N_5019,N_1791);
nand U6080 (N_6080,N_2666,N_2144);
or U6081 (N_6081,N_3258,N_2829);
or U6082 (N_6082,N_2231,N_5662);
nor U6083 (N_6083,N_3250,N_4104);
nand U6084 (N_6084,N_1409,N_392);
xor U6085 (N_6085,N_4762,N_5879);
nand U6086 (N_6086,N_4599,N_86);
and U6087 (N_6087,N_1166,N_565);
or U6088 (N_6088,N_4434,N_522);
xor U6089 (N_6089,N_5336,N_5464);
xnor U6090 (N_6090,N_2766,N_3193);
nor U6091 (N_6091,N_986,N_3437);
nand U6092 (N_6092,N_3092,N_3965);
and U6093 (N_6093,N_5356,N_1818);
nand U6094 (N_6094,N_3626,N_2218);
nor U6095 (N_6095,N_4083,N_3035);
xor U6096 (N_6096,N_4930,N_3966);
or U6097 (N_6097,N_4203,N_5639);
or U6098 (N_6098,N_2526,N_4777);
xor U6099 (N_6099,N_34,N_730);
or U6100 (N_6100,N_4935,N_1061);
nand U6101 (N_6101,N_4729,N_2191);
or U6102 (N_6102,N_1934,N_925);
nand U6103 (N_6103,N_726,N_3722);
xor U6104 (N_6104,N_3124,N_3941);
or U6105 (N_6105,N_3862,N_2304);
and U6106 (N_6106,N_3885,N_3260);
and U6107 (N_6107,N_3378,N_582);
and U6108 (N_6108,N_3677,N_687);
and U6109 (N_6109,N_385,N_5036);
xor U6110 (N_6110,N_2314,N_3096);
xor U6111 (N_6111,N_4184,N_4485);
nand U6112 (N_6112,N_56,N_9);
nand U6113 (N_6113,N_2488,N_4367);
nor U6114 (N_6114,N_2186,N_510);
and U6115 (N_6115,N_3738,N_4009);
or U6116 (N_6116,N_4281,N_394);
xnor U6117 (N_6117,N_5306,N_689);
and U6118 (N_6118,N_300,N_5567);
nor U6119 (N_6119,N_2305,N_1198);
xor U6120 (N_6120,N_5146,N_2598);
nand U6121 (N_6121,N_5178,N_1862);
or U6122 (N_6122,N_5027,N_3132);
xor U6123 (N_6123,N_3120,N_1574);
nand U6124 (N_6124,N_3434,N_5703);
nor U6125 (N_6125,N_409,N_5965);
or U6126 (N_6126,N_4385,N_4889);
xor U6127 (N_6127,N_5562,N_732);
nor U6128 (N_6128,N_2262,N_2953);
xor U6129 (N_6129,N_3975,N_1567);
xor U6130 (N_6130,N_1648,N_3864);
nor U6131 (N_6131,N_1318,N_2960);
nor U6132 (N_6132,N_2241,N_3960);
nand U6133 (N_6133,N_1199,N_3526);
nor U6134 (N_6134,N_377,N_5883);
or U6135 (N_6135,N_5611,N_560);
xor U6136 (N_6136,N_684,N_5067);
and U6137 (N_6137,N_5949,N_928);
nor U6138 (N_6138,N_3175,N_353);
xnor U6139 (N_6139,N_4261,N_2642);
xor U6140 (N_6140,N_2476,N_973);
or U6141 (N_6141,N_1007,N_996);
nand U6142 (N_6142,N_1216,N_5574);
nor U6143 (N_6143,N_2919,N_4972);
nand U6144 (N_6144,N_1487,N_1201);
nand U6145 (N_6145,N_3304,N_4956);
nand U6146 (N_6146,N_2817,N_2914);
nand U6147 (N_6147,N_317,N_3908);
xor U6148 (N_6148,N_4021,N_3167);
xor U6149 (N_6149,N_2145,N_2871);
xor U6150 (N_6150,N_248,N_5234);
nand U6151 (N_6151,N_1405,N_4269);
and U6152 (N_6152,N_4005,N_1400);
nand U6153 (N_6153,N_890,N_1456);
xor U6154 (N_6154,N_1165,N_2189);
nor U6155 (N_6155,N_153,N_524);
xor U6156 (N_6156,N_4119,N_3054);
xnor U6157 (N_6157,N_2838,N_4460);
and U6158 (N_6158,N_2475,N_5612);
nand U6159 (N_6159,N_4846,N_847);
nand U6160 (N_6160,N_1247,N_1855);
nor U6161 (N_6161,N_5162,N_2224);
nand U6162 (N_6162,N_1143,N_354);
xnor U6163 (N_6163,N_3223,N_3221);
nand U6164 (N_6164,N_1939,N_5720);
nand U6165 (N_6165,N_5255,N_5559);
nand U6166 (N_6166,N_1974,N_674);
or U6167 (N_6167,N_5777,N_4257);
nand U6168 (N_6168,N_2843,N_5424);
xor U6169 (N_6169,N_5219,N_1011);
nor U6170 (N_6170,N_4939,N_4016);
nor U6171 (N_6171,N_3265,N_2353);
nor U6172 (N_6172,N_111,N_3334);
and U6173 (N_6173,N_2331,N_4076);
and U6174 (N_6174,N_2251,N_5359);
nand U6175 (N_6175,N_90,N_1685);
nor U6176 (N_6176,N_1493,N_4093);
nor U6177 (N_6177,N_1618,N_76);
and U6178 (N_6178,N_2935,N_4966);
xor U6179 (N_6179,N_3452,N_1438);
xnor U6180 (N_6180,N_1901,N_5414);
nor U6181 (N_6181,N_1367,N_783);
nand U6182 (N_6182,N_5322,N_2485);
nor U6183 (N_6183,N_1879,N_432);
nor U6184 (N_6184,N_2284,N_1859);
or U6185 (N_6185,N_2289,N_3114);
nand U6186 (N_6186,N_677,N_4399);
nor U6187 (N_6187,N_2882,N_830);
xnor U6188 (N_6188,N_4994,N_4763);
and U6189 (N_6189,N_3176,N_5990);
xor U6190 (N_6190,N_1333,N_4621);
and U6191 (N_6191,N_3263,N_1611);
or U6192 (N_6192,N_1086,N_262);
xnor U6193 (N_6193,N_3471,N_3292);
or U6194 (N_6194,N_5375,N_5515);
or U6195 (N_6195,N_515,N_5108);
or U6196 (N_6196,N_323,N_3234);
and U6197 (N_6197,N_4308,N_5230);
nor U6198 (N_6198,N_888,N_1945);
or U6199 (N_6199,N_4550,N_1768);
xor U6200 (N_6200,N_3492,N_3660);
and U6201 (N_6201,N_4409,N_4461);
and U6202 (N_6202,N_2761,N_1919);
and U6203 (N_6203,N_4857,N_2259);
and U6204 (N_6204,N_5817,N_2732);
or U6205 (N_6205,N_3565,N_1436);
and U6206 (N_6206,N_4751,N_1668);
nand U6207 (N_6207,N_2809,N_1226);
and U6208 (N_6208,N_3614,N_4917);
nand U6209 (N_6209,N_4125,N_1561);
nand U6210 (N_6210,N_3443,N_923);
and U6211 (N_6211,N_1569,N_2932);
nand U6212 (N_6212,N_612,N_4060);
or U6213 (N_6213,N_1620,N_1681);
or U6214 (N_6214,N_5792,N_1356);
nor U6215 (N_6215,N_4747,N_2789);
nand U6216 (N_6216,N_761,N_872);
nor U6217 (N_6217,N_4391,N_246);
or U6218 (N_6218,N_3371,N_4481);
xor U6219 (N_6219,N_107,N_1036);
nand U6220 (N_6220,N_4977,N_1653);
or U6221 (N_6221,N_4120,N_5663);
xor U6222 (N_6222,N_1120,N_1765);
or U6223 (N_6223,N_4144,N_1520);
nand U6224 (N_6224,N_1164,N_4472);
xnor U6225 (N_6225,N_5182,N_5010);
nand U6226 (N_6226,N_4275,N_5093);
or U6227 (N_6227,N_927,N_2473);
nand U6228 (N_6228,N_5962,N_957);
nor U6229 (N_6229,N_3217,N_2551);
xor U6230 (N_6230,N_3920,N_3629);
nand U6231 (N_6231,N_3529,N_3302);
xnor U6232 (N_6232,N_3773,N_636);
and U6233 (N_6233,N_1665,N_3098);
or U6234 (N_6234,N_4244,N_4771);
nor U6235 (N_6235,N_3473,N_4051);
or U6236 (N_6236,N_184,N_3744);
nor U6237 (N_6237,N_3026,N_5112);
or U6238 (N_6238,N_325,N_1630);
or U6239 (N_6239,N_3774,N_5077);
and U6240 (N_6240,N_588,N_3706);
nor U6241 (N_6241,N_4231,N_4013);
nand U6242 (N_6242,N_4830,N_2942);
and U6243 (N_6243,N_3600,N_5111);
nand U6244 (N_6244,N_537,N_2496);
xor U6245 (N_6245,N_3528,N_2084);
or U6246 (N_6246,N_1337,N_2061);
nand U6247 (N_6247,N_2280,N_4158);
nand U6248 (N_6248,N_750,N_2012);
nor U6249 (N_6249,N_5795,N_873);
and U6250 (N_6250,N_3802,N_3838);
or U6251 (N_6251,N_5429,N_5731);
nor U6252 (N_6252,N_4339,N_406);
xnor U6253 (N_6253,N_2612,N_5049);
xnor U6254 (N_6254,N_5051,N_757);
nor U6255 (N_6255,N_5915,N_1846);
nor U6256 (N_6256,N_1180,N_2320);
or U6257 (N_6257,N_843,N_4671);
nand U6258 (N_6258,N_2604,N_2132);
or U6259 (N_6259,N_768,N_2812);
or U6260 (N_6260,N_1625,N_5475);
nand U6261 (N_6261,N_5939,N_1524);
or U6262 (N_6262,N_1959,N_5593);
nand U6263 (N_6263,N_2039,N_2107);
nor U6264 (N_6264,N_5105,N_4784);
xnor U6265 (N_6265,N_5940,N_5625);
xor U6266 (N_6266,N_5344,N_5571);
nor U6267 (N_6267,N_3983,N_5706);
and U6268 (N_6268,N_4558,N_949);
or U6269 (N_6269,N_1457,N_414);
nor U6270 (N_6270,N_2811,N_1956);
xor U6271 (N_6271,N_1471,N_940);
and U6272 (N_6272,N_5269,N_2835);
nor U6273 (N_6273,N_4183,N_2694);
nand U6274 (N_6274,N_5589,N_4877);
nand U6275 (N_6275,N_2899,N_3927);
nand U6276 (N_6276,N_770,N_3429);
nand U6277 (N_6277,N_3758,N_2387);
or U6278 (N_6278,N_3638,N_3256);
or U6279 (N_6279,N_5839,N_3571);
and U6280 (N_6280,N_3532,N_965);
or U6281 (N_6281,N_2401,N_5914);
and U6282 (N_6282,N_742,N_5156);
xor U6283 (N_6283,N_4794,N_1327);
and U6284 (N_6284,N_3561,N_3654);
nand U6285 (N_6285,N_4851,N_1663);
xnor U6286 (N_6286,N_2322,N_5975);
nand U6287 (N_6287,N_3757,N_549);
nand U6288 (N_6288,N_1763,N_1809);
xnor U6289 (N_6289,N_1640,N_5153);
xnor U6290 (N_6290,N_4343,N_1897);
xor U6291 (N_6291,N_488,N_3649);
nor U6292 (N_6292,N_2067,N_4646);
nand U6293 (N_6293,N_4727,N_3008);
and U6294 (N_6294,N_3984,N_5404);
or U6295 (N_6295,N_1860,N_1651);
xnor U6296 (N_6296,N_4145,N_2009);
or U6297 (N_6297,N_849,N_1037);
nor U6298 (N_6298,N_4697,N_4664);
xor U6299 (N_6299,N_1417,N_4443);
and U6300 (N_6300,N_1711,N_5582);
nand U6301 (N_6301,N_2862,N_4881);
xnor U6302 (N_6302,N_1056,N_980);
and U6303 (N_6303,N_3714,N_5808);
xor U6304 (N_6304,N_4704,N_5550);
or U6305 (N_6305,N_1767,N_2661);
xor U6306 (N_6306,N_2866,N_5807);
nor U6307 (N_6307,N_1713,N_5691);
nor U6308 (N_6308,N_3659,N_1093);
nor U6309 (N_6309,N_917,N_5953);
and U6310 (N_6310,N_1552,N_4876);
nor U6311 (N_6311,N_4571,N_5159);
and U6312 (N_6312,N_4041,N_4225);
xnor U6313 (N_6313,N_5436,N_920);
xnor U6314 (N_6314,N_803,N_3786);
nor U6315 (N_6315,N_1116,N_4369);
nand U6316 (N_6316,N_1957,N_4624);
and U6317 (N_6317,N_992,N_790);
and U6318 (N_6318,N_5573,N_3266);
xnor U6319 (N_6319,N_4644,N_5561);
nor U6320 (N_6320,N_2435,N_498);
nor U6321 (N_6321,N_283,N_3921);
xnor U6322 (N_6322,N_2423,N_1499);
nand U6323 (N_6323,N_5856,N_5062);
nand U6324 (N_6324,N_2492,N_1124);
and U6325 (N_6325,N_642,N_2454);
nand U6326 (N_6326,N_975,N_4315);
or U6327 (N_6327,N_4819,N_3997);
and U6328 (N_6328,N_5614,N_2257);
nor U6329 (N_6329,N_39,N_2026);
xnor U6330 (N_6330,N_1264,N_3577);
xor U6331 (N_6331,N_1947,N_4642);
nor U6332 (N_6332,N_500,N_2710);
or U6333 (N_6333,N_471,N_5781);
nand U6334 (N_6334,N_1322,N_1677);
nand U6335 (N_6335,N_974,N_3582);
or U6336 (N_6336,N_2460,N_2287);
or U6337 (N_6337,N_669,N_100);
or U6338 (N_6338,N_4864,N_1971);
nand U6339 (N_6339,N_1381,N_5798);
nor U6340 (N_6340,N_4064,N_3350);
nand U6341 (N_6341,N_5125,N_4098);
nand U6342 (N_6342,N_3890,N_3592);
nor U6343 (N_6343,N_2464,N_4709);
xor U6344 (N_6344,N_3606,N_5673);
and U6345 (N_6345,N_5615,N_1310);
and U6346 (N_6346,N_5283,N_249);
nor U6347 (N_6347,N_4605,N_4252);
and U6348 (N_6348,N_4038,N_3243);
or U6349 (N_6349,N_2250,N_5860);
or U6350 (N_6350,N_16,N_132);
xnor U6351 (N_6351,N_2265,N_3464);
or U6352 (N_6352,N_5769,N_5348);
nand U6353 (N_6353,N_5849,N_505);
nand U6354 (N_6354,N_2137,N_5528);
xor U6355 (N_6355,N_2640,N_800);
nand U6356 (N_6356,N_3374,N_4015);
nand U6357 (N_6357,N_3916,N_2426);
xnor U6358 (N_6358,N_4742,N_3871);
nand U6359 (N_6359,N_5435,N_1410);
xnor U6360 (N_6360,N_3537,N_2714);
xor U6361 (N_6361,N_2610,N_752);
or U6362 (N_6362,N_881,N_3299);
nor U6363 (N_6363,N_3127,N_3988);
xnor U6364 (N_6364,N_2957,N_1909);
and U6365 (N_6365,N_2119,N_460);
nor U6366 (N_6366,N_1539,N_4173);
and U6367 (N_6367,N_2905,N_5232);
nand U6368 (N_6368,N_3116,N_804);
or U6369 (N_6369,N_2283,N_1760);
or U6370 (N_6370,N_2540,N_2611);
xnor U6371 (N_6371,N_5481,N_3849);
nand U6372 (N_6372,N_5568,N_4473);
or U6373 (N_6373,N_415,N_542);
and U6374 (N_6374,N_2839,N_5303);
or U6375 (N_6375,N_901,N_1761);
xnor U6376 (N_6376,N_1710,N_5324);
or U6377 (N_6377,N_4087,N_3663);
nor U6378 (N_6378,N_5823,N_2742);
xnor U6379 (N_6379,N_2529,N_5534);
or U6380 (N_6380,N_2748,N_3959);
xor U6381 (N_6381,N_1770,N_4874);
nor U6382 (N_6382,N_3465,N_1741);
xnor U6383 (N_6383,N_4816,N_517);
and U6384 (N_6384,N_2541,N_5835);
and U6385 (N_6385,N_80,N_4302);
or U6386 (N_6386,N_5327,N_1251);
and U6387 (N_6387,N_2066,N_1834);
or U6388 (N_6388,N_356,N_1683);
nor U6389 (N_6389,N_5422,N_3228);
or U6390 (N_6390,N_1387,N_3919);
nand U6391 (N_6391,N_3824,N_4475);
or U6392 (N_6392,N_2542,N_3767);
nand U6393 (N_6393,N_919,N_4833);
nand U6394 (N_6394,N_3589,N_1272);
or U6395 (N_6395,N_663,N_5367);
or U6396 (N_6396,N_1597,N_204);
or U6397 (N_6397,N_3605,N_4625);
and U6398 (N_6398,N_580,N_5253);
or U6399 (N_6399,N_703,N_5423);
nand U6400 (N_6400,N_3311,N_2318);
and U6401 (N_6401,N_2365,N_3544);
nor U6402 (N_6402,N_5305,N_1259);
and U6403 (N_6403,N_5821,N_278);
nor U6404 (N_6404,N_2254,N_5759);
nand U6405 (N_6405,N_1288,N_519);
nand U6406 (N_6406,N_4116,N_1397);
xor U6407 (N_6407,N_4483,N_478);
nand U6408 (N_6408,N_3355,N_4335);
xor U6409 (N_6409,N_328,N_879);
and U6410 (N_6410,N_3238,N_4871);
or U6411 (N_6411,N_3005,N_74);
or U6412 (N_6412,N_1549,N_5969);
or U6413 (N_6413,N_3891,N_3090);
and U6414 (N_6414,N_2726,N_3220);
nor U6415 (N_6415,N_3349,N_1283);
or U6416 (N_6416,N_3109,N_1884);
nor U6417 (N_6417,N_4793,N_1488);
nor U6418 (N_6418,N_1350,N_2692);
nor U6419 (N_6419,N_434,N_4907);
xnor U6420 (N_6420,N_1428,N_3889);
or U6421 (N_6421,N_340,N_2069);
and U6422 (N_6422,N_1641,N_2493);
xnor U6423 (N_6423,N_130,N_5413);
and U6424 (N_6424,N_2758,N_615);
xnor U6425 (N_6425,N_991,N_452);
xor U6426 (N_6426,N_1078,N_5024);
nor U6427 (N_6427,N_960,N_5878);
nand U6428 (N_6428,N_5836,N_1720);
or U6429 (N_6429,N_1261,N_2185);
or U6430 (N_6430,N_1700,N_2018);
nor U6431 (N_6431,N_2272,N_1654);
xnor U6432 (N_6432,N_84,N_1718);
nor U6433 (N_6433,N_4326,N_692);
nand U6434 (N_6434,N_3268,N_4345);
and U6435 (N_6435,N_455,N_2778);
nor U6436 (N_6436,N_5818,N_2444);
or U6437 (N_6437,N_3209,N_4542);
nand U6438 (N_6438,N_1298,N_655);
and U6439 (N_6439,N_1095,N_1090);
nand U6440 (N_6440,N_393,N_5671);
and U6441 (N_6441,N_3475,N_5207);
nand U6442 (N_6442,N_2215,N_1195);
xnor U6443 (N_6443,N_5983,N_711);
or U6444 (N_6444,N_1923,N_5124);
nand U6445 (N_6445,N_3608,N_5552);
xor U6446 (N_6446,N_5934,N_2856);
xnor U6447 (N_6447,N_4702,N_345);
nand U6448 (N_6448,N_5160,N_122);
nor U6449 (N_6449,N_3668,N_719);
and U6450 (N_6450,N_2507,N_5736);
xnor U6451 (N_6451,N_5901,N_2436);
nor U6452 (N_6452,N_3236,N_3763);
nor U6453 (N_6453,N_1058,N_2774);
or U6454 (N_6454,N_5627,N_3827);
and U6455 (N_6455,N_5987,N_3836);
and U6456 (N_6456,N_5674,N_2317);
or U6457 (N_6457,N_2765,N_1238);
xnor U6458 (N_6458,N_54,N_3195);
nand U6459 (N_6459,N_1032,N_3692);
nor U6460 (N_6460,N_1332,N_1338);
nor U6461 (N_6461,N_950,N_366);
and U6462 (N_6462,N_5091,N_4821);
or U6463 (N_6463,N_5985,N_5684);
nor U6464 (N_6464,N_5456,N_1925);
nor U6465 (N_6465,N_2762,N_405);
nor U6466 (N_6466,N_511,N_3548);
and U6467 (N_6467,N_5782,N_2879);
or U6468 (N_6468,N_4814,N_4682);
and U6469 (N_6469,N_2196,N_1542);
and U6470 (N_6470,N_4359,N_210);
or U6471 (N_6471,N_1723,N_5678);
or U6472 (N_6472,N_5623,N_1729);
nor U6473 (N_6473,N_2414,N_413);
nor U6474 (N_6474,N_1573,N_4528);
xnor U6475 (N_6475,N_3103,N_1759);
xnor U6476 (N_6476,N_4506,N_1406);
and U6477 (N_6477,N_2421,N_3314);
nand U6478 (N_6478,N_2588,N_5604);
and U6479 (N_6479,N_2617,N_2124);
or U6480 (N_6480,N_1798,N_4151);
or U6481 (N_6481,N_1015,N_5923);
and U6482 (N_6482,N_2977,N_3359);
nand U6483 (N_6483,N_5351,N_5932);
nand U6484 (N_6484,N_427,N_4560);
nand U6485 (N_6485,N_307,N_5911);
nand U6486 (N_6486,N_4324,N_2845);
nand U6487 (N_6487,N_2563,N_4892);
nor U6488 (N_6488,N_2213,N_5730);
xor U6489 (N_6489,N_3695,N_3460);
xor U6490 (N_6490,N_705,N_2915);
nor U6491 (N_6491,N_5804,N_1324);
and U6492 (N_6492,N_2759,N_1949);
nor U6493 (N_6493,N_5610,N_361);
nor U6494 (N_6494,N_2308,N_3915);
nand U6495 (N_6495,N_2357,N_4245);
or U6496 (N_6496,N_155,N_2913);
xnor U6497 (N_6497,N_104,N_5310);
xnor U6498 (N_6498,N_4731,N_4594);
and U6499 (N_6499,N_5080,N_4662);
nor U6500 (N_6500,N_2951,N_556);
and U6501 (N_6501,N_5974,N_4216);
nand U6502 (N_6502,N_2535,N_2567);
xor U6503 (N_6503,N_4898,N_5084);
nand U6504 (N_6504,N_5972,N_2249);
and U6505 (N_6505,N_2349,N_5756);
nor U6506 (N_6506,N_2029,N_1747);
xnor U6507 (N_6507,N_4698,N_499);
or U6508 (N_6508,N_4757,N_3515);
xor U6509 (N_6509,N_3701,N_3556);
and U6510 (N_6510,N_4578,N_2665);
and U6511 (N_6511,N_2115,N_4008);
nand U6512 (N_6512,N_2345,N_3211);
or U6513 (N_6513,N_1186,N_5921);
nor U6514 (N_6514,N_5815,N_3807);
nand U6515 (N_6515,N_2657,N_268);
nor U6516 (N_6516,N_2083,N_331);
nand U6517 (N_6517,N_697,N_976);
nor U6518 (N_6518,N_4810,N_5301);
nand U6519 (N_6519,N_495,N_1054);
xor U6520 (N_6520,N_4787,N_3046);
and U6521 (N_6521,N_5167,N_3888);
and U6522 (N_6522,N_3724,N_5579);
nor U6523 (N_6523,N_2232,N_2453);
or U6524 (N_6524,N_2489,N_2312);
xnor U6525 (N_6525,N_1613,N_4557);
and U6526 (N_6526,N_1751,N_5712);
nand U6527 (N_6527,N_189,N_5591);
nor U6528 (N_6528,N_1986,N_388);
and U6529 (N_6529,N_2568,N_3930);
nand U6530 (N_6530,N_4386,N_5029);
nand U6531 (N_6531,N_1583,N_5938);
xnor U6532 (N_6532,N_1148,N_2854);
or U6533 (N_6533,N_3168,N_1498);
and U6534 (N_6534,N_2499,N_2670);
and U6535 (N_6535,N_2530,N_1132);
nand U6536 (N_6536,N_187,N_3316);
nand U6537 (N_6537,N_2350,N_2021);
xor U6538 (N_6538,N_827,N_5605);
nand U6539 (N_6539,N_4659,N_3403);
xor U6540 (N_6540,N_3653,N_2219);
xor U6541 (N_6541,N_5284,N_4541);
and U6542 (N_6542,N_3157,N_4786);
xnor U6543 (N_6543,N_17,N_5544);
and U6544 (N_6544,N_3164,N_2374);
nor U6545 (N_6545,N_3410,N_1541);
nor U6546 (N_6546,N_583,N_2303);
or U6547 (N_6547,N_4209,N_5026);
and U6548 (N_6548,N_3611,N_2474);
or U6549 (N_6549,N_1721,N_4572);
nor U6550 (N_6550,N_4983,N_2908);
nor U6551 (N_6551,N_4129,N_2141);
nand U6552 (N_6552,N_1755,N_4897);
and U6553 (N_6553,N_2457,N_4053);
and U6554 (N_6554,N_621,N_1246);
nor U6555 (N_6555,N_1212,N_2577);
or U6556 (N_6556,N_889,N_3448);
nand U6557 (N_6557,N_3257,N_2652);
nand U6558 (N_6558,N_5332,N_971);
xnor U6559 (N_6559,N_2204,N_3187);
nor U6560 (N_6560,N_138,N_2991);
or U6561 (N_6561,N_2878,N_1485);
or U6562 (N_6562,N_215,N_1109);
xor U6563 (N_6563,N_182,N_1494);
and U6564 (N_6564,N_5176,N_5236);
and U6565 (N_6565,N_3541,N_929);
xor U6566 (N_6566,N_2886,N_5387);
or U6567 (N_6567,N_1068,N_239);
xnor U6568 (N_6568,N_247,N_575);
xor U6569 (N_6569,N_2355,N_4878);
xor U6570 (N_6570,N_2220,N_5063);
and U6571 (N_6571,N_3514,N_3141);
nor U6572 (N_6572,N_1534,N_5247);
and U6573 (N_6573,N_1894,N_877);
nand U6574 (N_6574,N_3368,N_5169);
nor U6575 (N_6575,N_5383,N_1173);
nor U6576 (N_6576,N_4651,N_4573);
xnor U6577 (N_6577,N_5150,N_3341);
nor U6578 (N_6578,N_5364,N_3790);
xnor U6579 (N_6579,N_2070,N_4860);
nor U6580 (N_6580,N_2597,N_2150);
xor U6581 (N_6581,N_3093,N_2389);
and U6582 (N_6582,N_2086,N_2931);
or U6583 (N_6583,N_5199,N_2082);
and U6584 (N_6584,N_5813,N_475);
nand U6585 (N_6585,N_381,N_106);
or U6586 (N_6586,N_2638,N_3754);
xor U6587 (N_6587,N_1140,N_4527);
nor U6588 (N_6588,N_846,N_4420);
or U6589 (N_6589,N_3558,N_1952);
xnor U6590 (N_6590,N_1598,N_5127);
and U6591 (N_6591,N_1865,N_1800);
xor U6592 (N_6592,N_5157,N_1447);
nand U6593 (N_6593,N_1468,N_64);
and U6594 (N_6594,N_2025,N_4135);
nor U6595 (N_6595,N_1245,N_3749);
or U6596 (N_6596,N_648,N_5099);
nor U6597 (N_6597,N_4012,N_4312);
and U6598 (N_6598,N_2586,N_797);
nand U6599 (N_6599,N_3297,N_3731);
nor U6600 (N_6600,N_3992,N_4039);
and U6601 (N_6601,N_3237,N_4118);
or U6602 (N_6602,N_4303,N_1817);
or U6603 (N_6603,N_98,N_2771);
nor U6604 (N_6604,N_914,N_3881);
xor U6605 (N_6605,N_24,N_1847);
and U6606 (N_6606,N_1887,N_379);
and U6607 (N_6607,N_2757,N_5225);
nand U6608 (N_6608,N_428,N_3310);
xnor U6609 (N_6609,N_124,N_4791);
and U6610 (N_6610,N_3761,N_989);
nand U6611 (N_6611,N_5704,N_3696);
nand U6612 (N_6612,N_4946,N_2966);
nand U6613 (N_6613,N_2619,N_3624);
or U6614 (N_6614,N_4724,N_1652);
nor U6615 (N_6615,N_4054,N_4719);
nand U6616 (N_6616,N_1548,N_3408);
and U6617 (N_6617,N_1983,N_5347);
and U6618 (N_6618,N_2352,N_4568);
and U6619 (N_6619,N_2596,N_1948);
nor U6620 (N_6620,N_5449,N_3906);
nand U6621 (N_6621,N_3907,N_224);
nand U6622 (N_6622,N_2669,N_5362);
xor U6623 (N_6623,N_1273,N_5374);
xor U6624 (N_6624,N_2266,N_4411);
nand U6625 (N_6625,N_2920,N_2092);
nand U6626 (N_6626,N_948,N_4358);
and U6627 (N_6627,N_2902,N_1980);
nand U6628 (N_6628,N_5330,N_1207);
nor U6629 (N_6629,N_823,N_4371);
nor U6630 (N_6630,N_1523,N_469);
xnor U6631 (N_6631,N_5621,N_5014);
nand U6632 (N_6632,N_3137,N_2857);
xor U6633 (N_6633,N_252,N_4912);
and U6634 (N_6634,N_2667,N_1411);
or U6635 (N_6635,N_2122,N_2593);
nor U6636 (N_6636,N_982,N_3099);
xnor U6637 (N_6637,N_4139,N_2654);
and U6638 (N_6638,N_2471,N_2998);
xnor U6639 (N_6639,N_4000,N_3112);
nor U6640 (N_6640,N_5771,N_1267);
or U6641 (N_6641,N_3777,N_22);
nand U6642 (N_6642,N_363,N_26);
xor U6643 (N_6643,N_3402,N_3886);
nand U6644 (N_6644,N_1973,N_2344);
xor U6645 (N_6645,N_375,N_5406);
and U6646 (N_6646,N_5812,N_2978);
and U6647 (N_6647,N_5187,N_2851);
nor U6648 (N_6648,N_1257,N_685);
nor U6649 (N_6649,N_1138,N_1535);
or U6650 (N_6650,N_5851,N_5810);
or U6651 (N_6651,N_1135,N_3230);
or U6652 (N_6652,N_2909,N_2643);
and U6653 (N_6653,N_3521,N_3661);
nand U6654 (N_6654,N_170,N_3972);
and U6655 (N_6655,N_1857,N_270);
and U6656 (N_6656,N_4641,N_5055);
nor U6657 (N_6657,N_3647,N_2672);
nor U6658 (N_6658,N_5743,N_3075);
xnor U6659 (N_6659,N_444,N_3644);
or U6660 (N_6660,N_310,N_4467);
nor U6661 (N_6661,N_3159,N_3152);
or U6662 (N_6662,N_4480,N_3779);
nand U6663 (N_6663,N_1566,N_4337);
and U6664 (N_6664,N_1014,N_4272);
xor U6665 (N_6665,N_5496,N_3513);
and U6666 (N_6666,N_3004,N_4091);
and U6667 (N_6667,N_5829,N_4141);
and U6668 (N_6668,N_1915,N_4859);
or U6669 (N_6669,N_5126,N_1098);
or U6670 (N_6670,N_1395,N_978);
xnor U6671 (N_6671,N_3950,N_1740);
xnor U6672 (N_6672,N_3699,N_2227);
xnor U6673 (N_6673,N_3043,N_2383);
or U6674 (N_6674,N_3524,N_2849);
or U6675 (N_6675,N_5493,N_4370);
nor U6676 (N_6676,N_2199,N_2688);
or U6677 (N_6677,N_391,N_5694);
and U6678 (N_6678,N_3106,N_41);
or U6679 (N_6679,N_5098,N_4354);
and U6680 (N_6680,N_4344,N_2295);
xnor U6681 (N_6681,N_2707,N_4404);
and U6682 (N_6682,N_352,N_1811);
nor U6683 (N_6683,N_274,N_4538);
xnor U6684 (N_6684,N_3356,N_4749);
nand U6685 (N_6685,N_3946,N_1530);
or U6686 (N_6686,N_2217,N_3675);
and U6687 (N_6687,N_5842,N_4523);
or U6688 (N_6688,N_5827,N_4843);
or U6689 (N_6689,N_5622,N_206);
and U6690 (N_6690,N_1850,N_1204);
xor U6691 (N_6691,N_3769,N_5913);
nand U6692 (N_6692,N_955,N_3436);
xor U6693 (N_6693,N_5905,N_778);
xor U6694 (N_6694,N_3361,N_4736);
xnor U6695 (N_6695,N_2859,N_298);
and U6696 (N_6696,N_5007,N_125);
nor U6697 (N_6697,N_3181,N_4804);
xor U6698 (N_6698,N_3598,N_5039);
or U6699 (N_6699,N_4365,N_733);
nand U6700 (N_6700,N_857,N_2425);
nand U6701 (N_6701,N_3657,N_4375);
nand U6702 (N_6702,N_4580,N_1353);
xnor U6703 (N_6703,N_734,N_3451);
or U6704 (N_6704,N_5843,N_1179);
xor U6705 (N_6705,N_5458,N_2051);
nand U6706 (N_6706,N_1,N_1780);
and U6707 (N_6707,N_1679,N_1906);
nand U6708 (N_6708,N_2651,N_3926);
nor U6709 (N_6709,N_3380,N_3282);
and U6710 (N_6710,N_376,N_4915);
and U6711 (N_6711,N_1984,N_3755);
and U6712 (N_6712,N_3840,N_2623);
and U6713 (N_6713,N_3583,N_1152);
and U6714 (N_6714,N_1737,N_5064);
nor U6715 (N_6715,N_1946,N_2833);
or U6716 (N_6716,N_700,N_5747);
and U6717 (N_6717,N_3364,N_5186);
nand U6718 (N_6718,N_1790,N_745);
and U6719 (N_6719,N_373,N_4903);
nand U6720 (N_6720,N_5050,N_401);
and U6721 (N_6721,N_5648,N_2687);
xnor U6722 (N_6722,N_2068,N_4926);
xnor U6723 (N_6723,N_1486,N_1743);
or U6724 (N_6724,N_1933,N_3549);
or U6725 (N_6725,N_1803,N_767);
xnor U6726 (N_6726,N_3839,N_4368);
nand U6727 (N_6727,N_2721,N_319);
and U6728 (N_6728,N_2292,N_289);
nor U6729 (N_6729,N_4705,N_1013);
nor U6730 (N_6730,N_1635,N_675);
nor U6731 (N_6731,N_4142,N_1810);
nand U6732 (N_6732,N_5685,N_78);
nand U6733 (N_6733,N_4925,N_390);
nand U6734 (N_6734,N_2403,N_3478);
nor U6735 (N_6735,N_3252,N_5196);
and U6736 (N_6736,N_3856,N_855);
nor U6737 (N_6737,N_3142,N_1155);
nand U6738 (N_6738,N_4507,N_1000);
xnor U6739 (N_6739,N_1105,N_3367);
nand U6740 (N_6740,N_2558,N_5242);
or U6741 (N_6741,N_3625,N_4088);
xor U6742 (N_6742,N_904,N_459);
and U6743 (N_6743,N_46,N_2979);
nand U6744 (N_6744,N_431,N_527);
or U6745 (N_6745,N_2959,N_4462);
and U6746 (N_6746,N_4962,N_5483);
and U6747 (N_6747,N_3053,N_4271);
and U6748 (N_6748,N_5956,N_4640);
and U6749 (N_6749,N_1392,N_598);
and U6750 (N_6750,N_3705,N_3887);
nand U6751 (N_6751,N_1188,N_2136);
or U6752 (N_6752,N_5554,N_195);
nor U6753 (N_6753,N_3486,N_2827);
nand U6754 (N_6754,N_3918,N_3493);
or U6755 (N_6755,N_2163,N_5106);
nand U6756 (N_6756,N_1094,N_1500);
and U6757 (N_6757,N_5392,N_5906);
or U6758 (N_6758,N_4201,N_953);
nand U6759 (N_6759,N_5608,N_2585);
xor U6760 (N_6760,N_4685,N_3222);
nand U6761 (N_6761,N_4498,N_1473);
nor U6762 (N_6762,N_1529,N_1505);
nand U6763 (N_6763,N_2921,N_5396);
nand U6764 (N_6764,N_234,N_437);
and U6765 (N_6765,N_4208,N_680);
or U6766 (N_6766,N_2152,N_4613);
nor U6767 (N_6767,N_1328,N_322);
nand U6768 (N_6768,N_5741,N_1043);
or U6769 (N_6769,N_2552,N_2711);
xor U6770 (N_6770,N_4995,N_4159);
xor U6771 (N_6771,N_120,N_2801);
nand U6772 (N_6772,N_4658,N_2207);
and U6773 (N_6773,N_320,N_3284);
nand U6774 (N_6774,N_1682,N_3634);
nand U6775 (N_6775,N_1374,N_3148);
and U6776 (N_6776,N_2575,N_3765);
xor U6777 (N_6777,N_5733,N_1220);
xor U6778 (N_6778,N_2169,N_5037);
and U6779 (N_6779,N_5686,N_1060);
xor U6780 (N_6780,N_4520,N_316);
or U6781 (N_6781,N_5945,N_4808);
nand U6782 (N_6782,N_5624,N_4073);
nor U6783 (N_6783,N_1227,N_810);
xnor U6784 (N_6784,N_1293,N_555);
and U6785 (N_6785,N_237,N_841);
and U6786 (N_6786,N_3775,N_5787);
nand U6787 (N_6787,N_5390,N_3791);
xnor U6788 (N_6788,N_5556,N_1582);
or U6789 (N_6789,N_3693,N_372);
nor U6790 (N_6790,N_1039,N_5012);
and U6791 (N_6791,N_5718,N_383);
nor U6792 (N_6792,N_4361,N_5060);
nor U6793 (N_6793,N_1225,N_3752);
xor U6794 (N_6794,N_4026,N_1063);
nand U6795 (N_6795,N_209,N_4495);
xor U6796 (N_6796,N_50,N_5546);
and U6797 (N_6797,N_2553,N_2723);
and U6798 (N_6798,N_2660,N_424);
nor U6799 (N_6799,N_5926,N_4024);
nand U6800 (N_6800,N_1123,N_5352);
nor U6801 (N_6801,N_1268,N_1329);
nor U6802 (N_6802,N_1988,N_1291);
nor U6803 (N_6803,N_1176,N_5518);
or U6804 (N_6804,N_4400,N_4459);
and U6805 (N_6805,N_2539,N_3848);
or U6806 (N_6806,N_599,N_1205);
nor U6807 (N_6807,N_1435,N_3196);
nor U6808 (N_6808,N_337,N_32);
and U6809 (N_6809,N_4147,N_507);
and U6810 (N_6810,N_1444,N_1900);
nand U6811 (N_6811,N_72,N_2749);
or U6812 (N_6812,N_1836,N_2698);
or U6813 (N_6813,N_2434,N_2256);
nor U6814 (N_6814,N_2999,N_4295);
nor U6815 (N_6815,N_1875,N_5188);
and U6816 (N_6816,N_2573,N_5655);
and U6817 (N_6817,N_4427,N_922);
and U6818 (N_6818,N_2176,N_1145);
xnor U6819 (N_6819,N_5003,N_787);
and U6820 (N_6820,N_3427,N_3409);
or U6821 (N_6821,N_464,N_5031);
xnor U6822 (N_6822,N_5758,N_173);
nand U6823 (N_6823,N_1448,N_443);
nor U6824 (N_6824,N_186,N_656);
and U6825 (N_6825,N_4957,N_466);
xnor U6826 (N_6826,N_338,N_5948);
nand U6827 (N_6827,N_1987,N_4853);
nand U6828 (N_6828,N_1290,N_893);
xor U6829 (N_6829,N_5056,N_4306);
xnor U6830 (N_6830,N_3850,N_4728);
nor U6831 (N_6831,N_4469,N_2116);
xnor U6832 (N_6832,N_4772,N_3557);
or U6833 (N_6833,N_5498,N_2469);
nand U6834 (N_6834,N_1701,N_5198);
and U6835 (N_6835,N_4077,N_2121);
nand U6836 (N_6836,N_1966,N_2524);
xor U6837 (N_6837,N_1576,N_2715);
nor U6838 (N_6838,N_3831,N_4489);
nand U6839 (N_6839,N_4206,N_3305);
nand U6840 (N_6840,N_962,N_3423);
nand U6841 (N_6841,N_5780,N_2875);
or U6842 (N_6842,N_5005,N_1252);
xor U6843 (N_6843,N_1311,N_410);
and U6844 (N_6844,N_2739,N_3318);
xnor U6845 (N_6845,N_535,N_1289);
and U6846 (N_6846,N_759,N_3772);
and U6847 (N_6847,N_1807,N_3003);
and U6848 (N_6848,N_1872,N_343);
or U6849 (N_6849,N_2546,N_2613);
nand U6850 (N_6850,N_1624,N_5858);
xnor U6851 (N_6851,N_4942,N_3447);
nor U6852 (N_6852,N_351,N_2709);
xnor U6853 (N_6853,N_4899,N_473);
xnor U6854 (N_6854,N_1234,N_2428);
nand U6855 (N_6855,N_3275,N_3672);
or U6856 (N_6856,N_3279,N_762);
or U6857 (N_6857,N_3235,N_1602);
or U6858 (N_6858,N_1334,N_5749);
or U6859 (N_6859,N_1804,N_4812);
xnor U6860 (N_6860,N_2171,N_4327);
nand U6861 (N_6861,N_5581,N_5788);
and U6862 (N_6862,N_5935,N_2745);
and U6863 (N_6863,N_4497,N_3588);
nor U6864 (N_6864,N_5669,N_5928);
nand U6865 (N_6865,N_1680,N_509);
and U6866 (N_6866,N_4268,N_1231);
or U6867 (N_6867,N_4233,N_2060);
and U6868 (N_6868,N_845,N_2336);
xnor U6869 (N_6869,N_2673,N_4122);
xor U6870 (N_6870,N_5337,N_2294);
xor U6871 (N_6871,N_4955,N_2699);
and U6872 (N_6872,N_5488,N_1295);
xnor U6873 (N_6873,N_5875,N_3956);
nor U6874 (N_6874,N_1981,N_3795);
nand U6875 (N_6875,N_5087,N_4811);
nand U6876 (N_6876,N_3119,N_3023);
xnor U6877 (N_6877,N_3902,N_4928);
and U6878 (N_6878,N_4867,N_924);
xnor U6879 (N_6879,N_3129,N_1614);
nor U6880 (N_6880,N_3426,N_4547);
or U6881 (N_6881,N_1712,N_290);
nor U6882 (N_6882,N_3233,N_5532);
or U6883 (N_6883,N_5081,N_1315);
nor U6884 (N_6884,N_562,N_2646);
and U6885 (N_6885,N_5831,N_676);
nor U6886 (N_6886,N_765,N_2011);
and U6887 (N_6887,N_1131,N_4865);
nor U6888 (N_6888,N_4178,N_4788);
or U6889 (N_6889,N_910,N_2872);
or U6890 (N_6890,N_2351,N_5372);
nor U6891 (N_6891,N_3205,N_40);
and U6892 (N_6892,N_176,N_1472);
and U6893 (N_6893,N_1795,N_3563);
nand U6894 (N_6894,N_5477,N_2948);
and U6895 (N_6895,N_5313,N_3736);
nor U6896 (N_6896,N_744,N_597);
or U6897 (N_6897,N_2776,N_4850);
or U6898 (N_6898,N_1189,N_2702);
or U6899 (N_6899,N_2341,N_5393);
nor U6900 (N_6900,N_2200,N_2779);
and U6901 (N_6901,N_5834,N_2035);
nor U6902 (N_6902,N_4065,N_3594);
xor U6903 (N_6903,N_3851,N_3165);
xnor U6904 (N_6904,N_5806,N_1935);
nand U6905 (N_6905,N_219,N_4562);
or U6906 (N_6906,N_2030,N_1321);
and U6907 (N_6907,N_4979,N_2390);
nand U6908 (N_6908,N_5457,N_3747);
xnor U6909 (N_6909,N_2730,N_1829);
and U6910 (N_6910,N_2085,N_3002);
xnor U6911 (N_6911,N_4106,N_1206);
nand U6912 (N_6912,N_1174,N_1788);
or U6913 (N_6913,N_3999,N_2881);
nor U6914 (N_6914,N_5223,N_2140);
or U6915 (N_6915,N_4396,N_5045);
nand U6916 (N_6916,N_1589,N_2716);
nor U6917 (N_6917,N_4305,N_156);
and U6918 (N_6918,N_5292,N_4290);
and U6919 (N_6919,N_5767,N_5213);
and U6920 (N_6920,N_1170,N_2797);
or U6921 (N_6921,N_2164,N_1158);
nand U6922 (N_6922,N_961,N_3071);
nor U6923 (N_6923,N_4107,N_3704);
xnor U6924 (N_6924,N_493,N_3457);
and U6925 (N_6925,N_1218,N_4432);
nand U6926 (N_6926,N_1714,N_5547);
and U6927 (N_6927,N_3750,N_4200);
and U6928 (N_6928,N_5872,N_717);
or U6929 (N_6929,N_2740,N_344);
and U6930 (N_6930,N_826,N_4818);
or U6931 (N_6931,N_1644,N_3425);
xor U6932 (N_6932,N_2521,N_5331);
or U6933 (N_6933,N_2052,N_3462);
nand U6934 (N_6934,N_5785,N_4049);
and U6935 (N_6935,N_4463,N_1732);
and U6936 (N_6936,N_2465,N_866);
and U6937 (N_6937,N_4470,N_5251);
or U6938 (N_6938,N_3785,N_450);
and U6939 (N_6939,N_1142,N_3709);
and U6940 (N_6940,N_1483,N_131);
nor U6941 (N_6941,N_5200,N_2903);
or U6942 (N_6942,N_3485,N_3715);
nand U6943 (N_6943,N_4214,N_2327);
or U6944 (N_6944,N_435,N_3825);
nor U6945 (N_6945,N_821,N_2388);
and U6946 (N_6946,N_3045,N_1408);
nand U6947 (N_6947,N_4040,N_2703);
xor U6948 (N_6948,N_3698,N_1031);
xor U6949 (N_6949,N_3014,N_5893);
and U6950 (N_6950,N_5832,N_609);
and U6951 (N_6951,N_746,N_4920);
nand U6952 (N_6952,N_2805,N_5408);
or U6953 (N_6953,N_725,N_2214);
and U6954 (N_6954,N_4117,N_3333);
xor U6955 (N_6955,N_3082,N_1434);
or U6956 (N_6956,N_1262,N_3384);
or U6957 (N_6957,N_4519,N_149);
nor U6958 (N_6958,N_5100,N_3012);
or U6959 (N_6959,N_2258,N_110);
and U6960 (N_6960,N_4629,N_5418);
and U6961 (N_6961,N_2372,N_1057);
nand U6962 (N_6962,N_2609,N_165);
nor U6963 (N_6963,N_4575,N_4169);
and U6964 (N_6964,N_1782,N_2691);
and U6965 (N_6965,N_1167,N_5877);
or U6966 (N_6966,N_589,N_1661);
nor U6967 (N_6967,N_151,N_2015);
nand U6968 (N_6968,N_2988,N_2206);
or U6969 (N_6969,N_5626,N_3903);
nand U6970 (N_6970,N_1129,N_2382);
nand U6971 (N_6971,N_1642,N_3841);
and U6972 (N_6972,N_4389,N_5235);
and U6973 (N_6973,N_3742,N_2293);
or U6974 (N_6974,N_3671,N_664);
nor U6975 (N_6975,N_3658,N_190);
and U6976 (N_6976,N_3799,N_2794);
and U6977 (N_6977,N_3084,N_4700);
nand U6978 (N_6978,N_4328,N_2024);
or U6979 (N_6979,N_2570,N_3746);
xnor U6980 (N_6980,N_754,N_243);
and U6981 (N_6981,N_4477,N_433);
nand U6982 (N_6982,N_3301,N_5398);
nor U6983 (N_6983,N_3844,N_2362);
and U6984 (N_6984,N_83,N_569);
xor U6985 (N_6985,N_2307,N_1437);
xnor U6986 (N_6986,N_4334,N_3197);
and U6987 (N_6987,N_2095,N_3433);
and U6988 (N_6988,N_5042,N_220);
xnor U6989 (N_6989,N_3734,N_5679);
or U6990 (N_6990,N_1233,N_4342);
and U6991 (N_6991,N_1612,N_5462);
xnor U6992 (N_6992,N_3879,N_3554);
xor U6993 (N_6993,N_5564,N_5116);
nand U6994 (N_6994,N_5964,N_5907);
xor U6995 (N_6995,N_5784,N_4249);
and U6996 (N_6996,N_4100,N_964);
nor U6997 (N_6997,N_1786,N_1601);
and U6998 (N_6998,N_1728,N_4609);
xnor U6999 (N_6999,N_5664,N_2744);
nand U7000 (N_7000,N_1756,N_3272);
nand U7001 (N_7001,N_492,N_3837);
or U7002 (N_7002,N_4199,N_4392);
nand U7003 (N_7003,N_2561,N_5727);
nand U7004 (N_7004,N_2910,N_2438);
nor U7005 (N_7005,N_788,N_2441);
or U7006 (N_7006,N_454,N_4894);
xor U7007 (N_7007,N_3110,N_3179);
nor U7008 (N_7008,N_1475,N_4366);
nand U7009 (N_7009,N_2267,N_57);
nand U7010 (N_7010,N_3271,N_3444);
nand U7011 (N_7011,N_4044,N_912);
xor U7012 (N_7012,N_1431,N_2777);
and U7013 (N_7013,N_1594,N_5680);
nand U7014 (N_7014,N_2056,N_5034);
xnor U7015 (N_7015,N_2595,N_5307);
nand U7016 (N_7016,N_4378,N_4929);
or U7017 (N_7017,N_3140,N_5376);
xnor U7018 (N_7018,N_2182,N_3778);
and U7019 (N_7019,N_256,N_3913);
and U7020 (N_7020,N_99,N_5701);
or U7021 (N_7021,N_5489,N_4037);
xor U7022 (N_7022,N_4155,N_2161);
or U7023 (N_7023,N_2967,N_728);
and U7024 (N_7024,N_1526,N_3454);
nor U7025 (N_7025,N_1596,N_1347);
nor U7026 (N_7026,N_2876,N_4796);
or U7027 (N_7027,N_5260,N_5389);
or U7028 (N_7028,N_2236,N_2046);
xnor U7029 (N_7029,N_2461,N_212);
nor U7030 (N_7030,N_4565,N_5994);
and U7031 (N_7031,N_3494,N_3076);
nor U7032 (N_7032,N_4316,N_5193);
and U7033 (N_7033,N_436,N_1912);
nor U7034 (N_7034,N_4759,N_4300);
nand U7035 (N_7035,N_4529,N_958);
and U7036 (N_7036,N_28,N_1831);
nand U7037 (N_7037,N_5619,N_4254);
or U7038 (N_7038,N_4061,N_3456);
xnor U7039 (N_7039,N_688,N_3463);
nor U7040 (N_7040,N_2746,N_4491);
xnor U7041 (N_7041,N_4256,N_5855);
nor U7042 (N_7042,N_313,N_1326);
and U7043 (N_7043,N_1600,N_4760);
and U7044 (N_7044,N_563,N_276);
nor U7045 (N_7045,N_1162,N_244);
and U7046 (N_7046,N_4235,N_611);
and U7047 (N_7047,N_2187,N_5342);
nand U7048 (N_7048,N_2027,N_3685);
or U7049 (N_7049,N_2040,N_1280);
xnor U7050 (N_7050,N_5930,N_741);
xor U7051 (N_7051,N_1970,N_3977);
nor U7052 (N_7052,N_2166,N_1643);
nand U7053 (N_7053,N_1610,N_1838);
and U7054 (N_7054,N_5555,N_2480);
nand U7055 (N_7055,N_3564,N_3335);
nor U7056 (N_7056,N_341,N_3809);
nand U7057 (N_7057,N_2080,N_421);
xnor U7058 (N_7058,N_2940,N_4032);
xnor U7059 (N_7059,N_1733,N_886);
or U7060 (N_7060,N_5101,N_5714);
xor U7061 (N_7061,N_1961,N_2574);
or U7062 (N_7062,N_3669,N_5020);
xnor U7063 (N_7063,N_4931,N_2239);
nand U7064 (N_7064,N_4603,N_27);
nor U7065 (N_7065,N_4207,N_3139);
xnor U7066 (N_7066,N_292,N_4425);
nor U7067 (N_7067,N_1401,N_4802);
and U7068 (N_7068,N_4504,N_2183);
nand U7069 (N_7069,N_1854,N_851);
and U7070 (N_7070,N_5038,N_3800);
or U7071 (N_7071,N_225,N_966);
nor U7072 (N_7072,N_735,N_5654);
or U7073 (N_7073,N_813,N_3893);
nand U7074 (N_7074,N_5558,N_5241);
and U7075 (N_7075,N_3030,N_1232);
or U7076 (N_7076,N_4959,N_3804);
nand U7077 (N_7077,N_1521,N_5638);
nor U7078 (N_7078,N_2321,N_5809);
or U7079 (N_7079,N_5864,N_5640);
nand U7080 (N_7080,N_3126,N_1028);
xor U7081 (N_7081,N_3283,N_4589);
or U7082 (N_7082,N_163,N_8);
xor U7083 (N_7083,N_2753,N_1399);
nand U7084 (N_7084,N_269,N_1927);
xnor U7085 (N_7085,N_1588,N_3718);
or U7086 (N_7086,N_139,N_3870);
or U7087 (N_7087,N_4297,N_2106);
and U7088 (N_7088,N_2032,N_916);
nor U7089 (N_7089,N_5583,N_5646);
nor U7090 (N_7090,N_2798,N_4554);
or U7091 (N_7091,N_3944,N_2731);
or U7092 (N_7092,N_1097,N_5887);
or U7093 (N_7093,N_4424,N_4555);
or U7094 (N_7094,N_1429,N_308);
and U7095 (N_7095,N_3108,N_476);
xnor U7096 (N_7096,N_1128,N_2884);
and U7097 (N_7097,N_694,N_3874);
nand U7098 (N_7098,N_2143,N_3185);
or U7099 (N_7099,N_5959,N_1509);
nor U7100 (N_7100,N_934,N_275);
nor U7101 (N_7101,N_1813,N_185);
and U7102 (N_7102,N_5577,N_780);
or U7103 (N_7103,N_3604,N_2071);
xnor U7104 (N_7104,N_3994,N_3496);
nor U7105 (N_7105,N_1066,N_5522);
xnor U7106 (N_7106,N_4017,N_5201);
nor U7107 (N_7107,N_5229,N_2162);
nand U7108 (N_7108,N_2579,N_2138);
or U7109 (N_7109,N_2495,N_627);
nand U7110 (N_7110,N_2523,N_605);
nand U7111 (N_7111,N_5035,N_3914);
or U7112 (N_7112,N_2118,N_3793);
and U7113 (N_7113,N_4707,N_2433);
nand U7114 (N_7114,N_2059,N_3990);
or U7115 (N_7115,N_2146,N_1554);
or U7116 (N_7116,N_3683,N_3635);
nand U7117 (N_7117,N_4373,N_2506);
and U7118 (N_7118,N_3896,N_5967);
xor U7119 (N_7119,N_5361,N_1719);
nand U7120 (N_7120,N_2173,N_4822);
xor U7121 (N_7121,N_324,N_3607);
and U7122 (N_7122,N_4110,N_279);
xnor U7123 (N_7123,N_1745,N_2028);
xor U7124 (N_7124,N_5998,N_848);
nand U7125 (N_7125,N_5531,N_2100);
xnor U7126 (N_7126,N_825,N_5570);
nor U7127 (N_7127,N_419,N_5656);
nor U7128 (N_7128,N_1636,N_4953);
or U7129 (N_7129,N_1543,N_3467);
xnor U7130 (N_7130,N_245,N_4773);
xnor U7131 (N_7131,N_5587,N_4314);
xor U7132 (N_7132,N_4287,N_3375);
xnor U7133 (N_7133,N_3495,N_4277);
xnor U7134 (N_7134,N_5563,N_3599);
nor U7135 (N_7135,N_4170,N_2622);
nor U7136 (N_7136,N_2602,N_903);
or U7137 (N_7137,N_81,N_4236);
and U7138 (N_7138,N_2768,N_1565);
nor U7139 (N_7139,N_1258,N_3413);
or U7140 (N_7140,N_5463,N_47);
or U7141 (N_7141,N_5256,N_5312);
and U7142 (N_7142,N_3432,N_3194);
xor U7143 (N_7143,N_2825,N_3530);
nor U7144 (N_7144,N_4998,N_1271);
nand U7145 (N_7145,N_193,N_291);
xor U7146 (N_7146,N_2420,N_2413);
xnor U7147 (N_7147,N_2101,N_4213);
nand U7148 (N_7148,N_4774,N_4265);
and U7149 (N_7149,N_5265,N_1202);
nand U7150 (N_7150,N_5797,N_468);
xnor U7151 (N_7151,N_4108,N_3146);
nor U7152 (N_7152,N_164,N_1689);
nor U7153 (N_7153,N_1802,N_3244);
nand U7154 (N_7154,N_2822,N_267);
and U7155 (N_7155,N_3089,N_4050);
and U7156 (N_7156,N_2394,N_4893);
nor U7157 (N_7157,N_937,N_2358);
and U7158 (N_7158,N_1622,N_82);
and U7159 (N_7159,N_3202,N_4712);
nand U7160 (N_7160,N_853,N_5816);
nor U7161 (N_7161,N_1866,N_5135);
or U7162 (N_7162,N_909,N_4886);
nor U7163 (N_7163,N_2212,N_2725);
nand U7164 (N_7164,N_2562,N_4232);
nor U7165 (N_7165,N_147,N_3925);
nand U7166 (N_7166,N_58,N_3042);
nand U7167 (N_7167,N_3218,N_4267);
xnor U7168 (N_7168,N_2468,N_2965);
and U7169 (N_7169,N_3174,N_5896);
or U7170 (N_7170,N_3155,N_5237);
xnor U7171 (N_7171,N_4453,N_4084);
nand U7172 (N_7172,N_4114,N_5961);
nand U7173 (N_7173,N_2005,N_3107);
nand U7174 (N_7174,N_5885,N_2277);
xor U7175 (N_7175,N_5596,N_1842);
nand U7176 (N_7176,N_2371,N_860);
or U7177 (N_7177,N_1511,N_5212);
nor U7178 (N_7178,N_4006,N_870);
and U7179 (N_7179,N_123,N_2990);
nand U7180 (N_7180,N_818,N_4493);
and U7181 (N_7181,N_5226,N_4633);
and U7182 (N_7182,N_1918,N_5320);
and U7183 (N_7183,N_5141,N_2343);
xor U7184 (N_7184,N_5764,N_2463);
nor U7185 (N_7185,N_3270,N_4732);
xor U7186 (N_7186,N_2511,N_4340);
xor U7187 (N_7187,N_907,N_4701);
nand U7188 (N_7188,N_1175,N_4514);
nor U7189 (N_7189,N_1112,N_2898);
and U7190 (N_7190,N_4444,N_312);
nand U7191 (N_7191,N_2151,N_3418);
nand U7192 (N_7192,N_5294,N_4815);
or U7193 (N_7193,N_590,N_2058);
and U7194 (N_7194,N_370,N_5128);
or U7195 (N_7195,N_1442,N_2270);
xnor U7196 (N_7196,N_2385,N_2587);
xor U7197 (N_7197,N_2681,N_5446);
nor U7198 (N_7198,N_4419,N_4849);
or U7199 (N_7199,N_602,N_5912);
nand U7200 (N_7200,N_5766,N_3676);
xor U7201 (N_7201,N_3177,N_3954);
or U7202 (N_7202,N_2923,N_4007);
nand U7203 (N_7203,N_4259,N_2243);
and U7204 (N_7204,N_4765,N_3694);
and U7205 (N_7205,N_2031,N_2108);
nand U7206 (N_7206,N_160,N_743);
nor U7207 (N_7207,N_1002,N_3111);
and U7208 (N_7208,N_5709,N_4918);
nand U7209 (N_7209,N_4789,N_1213);
nor U7210 (N_7210,N_3814,N_2361);
or U7211 (N_7211,N_1407,N_2201);
nor U7212 (N_7212,N_4204,N_5138);
nand U7213 (N_7213,N_502,N_3204);
nand U7214 (N_7214,N_5740,N_4611);
and U7215 (N_7215,N_607,N_5214);
and U7216 (N_7216,N_4681,N_1133);
nor U7217 (N_7217,N_2400,N_335);
xnor U7218 (N_7218,N_2004,N_5848);
nor U7219 (N_7219,N_3360,N_1470);
and U7220 (N_7220,N_4941,N_1744);
or U7221 (N_7221,N_5592,N_1746);
nand U7222 (N_7222,N_1194,N_5239);
nor U7223 (N_7223,N_4689,N_1025);
nor U7224 (N_7224,N_216,N_2252);
or U7225 (N_7225,N_2527,N_3006);
xor U7226 (N_7226,N_1826,N_4304);
nor U7227 (N_7227,N_868,N_3247);
xnor U7228 (N_7228,N_670,N_1623);
nor U7229 (N_7229,N_2041,N_3828);
nand U7230 (N_7230,N_3859,N_2452);
and U7231 (N_7231,N_5431,N_2550);
nor U7232 (N_7232,N_1766,N_667);
or U7233 (N_7233,N_1038,N_3041);
nor U7234 (N_7234,N_228,N_4202);
and U7235 (N_7235,N_3581,N_4778);
xor U7236 (N_7236,N_1477,N_89);
nor U7237 (N_7237,N_1221,N_400);
and U7238 (N_7238,N_4668,N_1581);
or U7239 (N_7239,N_4152,N_2557);
or U7240 (N_7240,N_867,N_559);
xor U7241 (N_7241,N_4680,N_4363);
or U7242 (N_7242,N_229,N_200);
nor U7243 (N_7243,N_2569,N_4845);
nor U7244 (N_7244,N_3681,N_1100);
nand U7245 (N_7245,N_5526,N_2288);
and U7246 (N_7246,N_4074,N_4748);
and U7247 (N_7247,N_1895,N_696);
or U7248 (N_7248,N_4847,N_640);
and U7249 (N_7249,N_2659,N_280);
xnor U7250 (N_7250,N_1647,N_3033);
nand U7251 (N_7251,N_1864,N_4672);
xor U7252 (N_7252,N_4058,N_263);
nor U7253 (N_7253,N_4258,N_4713);
nand U7254 (N_7254,N_706,N_3947);
or U7255 (N_7255,N_3337,N_619);
xor U7256 (N_7256,N_4932,N_4949);
nand U7257 (N_7257,N_3324,N_2858);
nor U7258 (N_7258,N_5113,N_2792);
nor U7259 (N_7259,N_4505,N_4683);
xnor U7260 (N_7260,N_4952,N_2044);
nor U7261 (N_7261,N_3048,N_1671);
or U7262 (N_7262,N_5161,N_1415);
nor U7263 (N_7263,N_5163,N_3477);
or U7264 (N_7264,N_2335,N_2177);
and U7265 (N_7265,N_4869,N_5172);
and U7266 (N_7266,N_51,N_686);
nand U7267 (N_7267,N_5,N_666);
and U7268 (N_7268,N_3397,N_763);
and U7269 (N_7269,N_4988,N_3121);
nand U7270 (N_7270,N_1306,N_2772);
or U7271 (N_7271,N_4014,N_5068);
or U7272 (N_7272,N_1699,N_3884);
nor U7273 (N_7273,N_3136,N_2995);
and U7274 (N_7274,N_1785,N_491);
and U7275 (N_7275,N_5250,N_4113);
nand U7276 (N_7276,N_3287,N_342);
nor U7277 (N_7277,N_5909,N_1183);
nor U7278 (N_7278,N_3531,N_3948);
xor U7279 (N_7279,N_5401,N_5861);
xnor U7280 (N_7280,N_3331,N_548);
nand U7281 (N_7281,N_5264,N_5025);
nand U7282 (N_7282,N_799,N_2234);
nor U7283 (N_7283,N_5041,N_5826);
and U7284 (N_7284,N_981,N_1362);
nor U7285 (N_7285,N_2629,N_5775);
xnor U7286 (N_7286,N_4584,N_4743);
or U7287 (N_7287,N_347,N_3213);
nand U7288 (N_7288,N_4655,N_1001);
or U7289 (N_7289,N_4336,N_181);
or U7290 (N_7290,N_4744,N_4197);
or U7291 (N_7291,N_1905,N_37);
and U7292 (N_7292,N_3508,N_5417);
nor U7293 (N_7293,N_2897,N_3697);
and U7294 (N_7294,N_2238,N_33);
and U7295 (N_7295,N_3569,N_2253);
or U7296 (N_7296,N_4924,N_772);
xnor U7297 (N_7297,N_2179,N_250);
or U7298 (N_7298,N_2786,N_5588);
and U7299 (N_7299,N_1968,N_1736);
or U7300 (N_7300,N_834,N_2606);
xor U7301 (N_7301,N_5951,N_2918);
nor U7302 (N_7302,N_755,N_4435);
nor U7303 (N_7303,N_382,N_1605);
xnor U7304 (N_7304,N_1070,N_5636);
and U7305 (N_7305,N_4364,N_727);
and U7306 (N_7306,N_3342,N_223);
xnor U7307 (N_7307,N_2081,N_3989);
nand U7308 (N_7308,N_2581,N_5958);
nand U7309 (N_7309,N_1515,N_5989);
or U7310 (N_7310,N_871,N_5954);
or U7311 (N_7311,N_2057,N_1999);
xor U7312 (N_7312,N_1911,N_1580);
and U7313 (N_7313,N_3585,N_945);
nor U7314 (N_7314,N_1119,N_3590);
nand U7315 (N_7315,N_947,N_4381);
and U7316 (N_7316,N_5254,N_4610);
nand U7317 (N_7317,N_994,N_2533);
nand U7318 (N_7318,N_3440,N_4164);
xor U7319 (N_7319,N_4508,N_1079);
nor U7320 (N_7320,N_4330,N_4805);
nor U7321 (N_7321,N_2938,N_2178);
xnor U7322 (N_7322,N_5419,N_4596);
and U7323 (N_7323,N_5382,N_4360);
or U7324 (N_7324,N_2724,N_3711);
nor U7325 (N_7325,N_528,N_2356);
and U7326 (N_7326,N_2456,N_5285);
xnor U7327 (N_7327,N_327,N_4943);
or U7328 (N_7328,N_4293,N_3843);
or U7329 (N_7329,N_5661,N_5281);
and U7330 (N_7330,N_2844,N_5649);
nand U7331 (N_7331,N_1960,N_4934);
nor U7332 (N_7332,N_1892,N_2407);
and U7333 (N_7333,N_2502,N_3855);
xnor U7334 (N_7334,N_3573,N_3484);
nor U7335 (N_7335,N_371,N_3060);
or U7336 (N_7336,N_4518,N_4048);
xor U7337 (N_7337,N_5575,N_3000);
nor U7338 (N_7338,N_1924,N_2367);
nand U7339 (N_7339,N_3832,N_4321);
xor U7340 (N_7340,N_812,N_273);
nor U7341 (N_7341,N_4067,N_3226);
nand U7342 (N_7342,N_942,N_828);
and U7343 (N_7343,N_5388,N_1102);
and U7344 (N_7344,N_5366,N_632);
nor U7345 (N_7345,N_2065,N_5793);
nor U7346 (N_7346,N_1670,N_5837);
xnor U7347 (N_7347,N_467,N_4488);
nand U7348 (N_7348,N_1376,N_4168);
or U7349 (N_7349,N_2720,N_4464);
or U7350 (N_7350,N_5043,N_2338);
nand U7351 (N_7351,N_174,N_5936);
xor U7352 (N_7352,N_3348,N_623);
and U7353 (N_7353,N_4895,N_5862);
or U7354 (N_7354,N_654,N_1508);
nor U7355 (N_7355,N_5869,N_418);
xnor U7356 (N_7356,N_15,N_2063);
xor U7357 (N_7357,N_984,N_4828);
or U7358 (N_7358,N_2576,N_2968);
or U7359 (N_7359,N_2603,N_3553);
or U7360 (N_7360,N_5380,N_5601);
and U7361 (N_7361,N_3325,N_251);
nand U7362 (N_7362,N_4717,N_5976);
and U7363 (N_7363,N_4652,N_5110);
and U7364 (N_7364,N_2770,N_3357);
and U7365 (N_7365,N_2880,N_3015);
or U7366 (N_7366,N_5880,N_5001);
nor U7367 (N_7367,N_2993,N_1380);
xnor U7368 (N_7368,N_779,N_1708);
xnor U7369 (N_7369,N_2727,N_91);
nand U7370 (N_7370,N_3725,N_3819);
nor U7371 (N_7371,N_523,N_161);
or U7372 (N_7372,N_2695,N_3506);
nand U7373 (N_7373,N_1722,N_5076);
nor U7374 (N_7374,N_486,N_4056);
nand U7375 (N_7375,N_1460,N_1147);
xnor U7376 (N_7376,N_5147,N_5672);
xnor U7377 (N_7377,N_3538,N_3013);
nor U7378 (N_7378,N_5197,N_1553);
xor U7379 (N_7379,N_4068,N_5659);
or U7380 (N_7380,N_1816,N_5323);
or U7381 (N_7381,N_1538,N_3062);
nor U7382 (N_7382,N_5154,N_3296);
or U7383 (N_7383,N_474,N_2398);
nand U7384 (N_7384,N_2290,N_2006);
nand U7385 (N_7385,N_3122,N_1481);
and U7386 (N_7386,N_4080,N_3379);
nor U7387 (N_7387,N_2937,N_295);
or U7388 (N_7388,N_584,N_3381);
and U7389 (N_7389,N_5218,N_5397);
nand U7390 (N_7390,N_2752,N_5379);
nor U7391 (N_7391,N_3149,N_3469);
nand U7392 (N_7392,N_784,N_2016);
and U7393 (N_7393,N_2892,N_3210);
nor U7394 (N_7394,N_2364,N_3666);
xor U7395 (N_7395,N_1352,N_4583);
or U7396 (N_7396,N_1853,N_4229);
nand U7397 (N_7397,N_1815,N_882);
and U7398 (N_7398,N_1287,N_3520);
or U7399 (N_7399,N_5870,N_3446);
nor U7400 (N_7400,N_3,N_1830);
xnor U7401 (N_7401,N_5018,N_1354);
xor U7402 (N_7402,N_3939,N_5073);
and U7403 (N_7403,N_1877,N_4134);
nor U7404 (N_7404,N_4066,N_3293);
and U7405 (N_7405,N_2980,N_2153);
nand U7406 (N_7406,N_5548,N_3512);
or U7407 (N_7407,N_5407,N_4820);
and U7408 (N_7408,N_4982,N_2738);
and U7409 (N_7409,N_3424,N_5286);
nand U7410 (N_7410,N_140,N_1867);
nor U7411 (N_7411,N_2451,N_4639);
or U7412 (N_7412,N_1965,N_95);
or U7413 (N_7413,N_5120,N_2271);
nor U7414 (N_7414,N_1035,N_521);
nor U7415 (N_7415,N_158,N_1419);
and U7416 (N_7416,N_1638,N_769);
and U7417 (N_7417,N_1008,N_801);
and U7418 (N_7418,N_2633,N_4753);
xnor U7419 (N_7419,N_4243,N_5293);
xnor U7420 (N_7420,N_1404,N_1517);
or U7421 (N_7421,N_4447,N_3808);
nand U7422 (N_7422,N_4004,N_1081);
or U7423 (N_7423,N_1331,N_3771);
nor U7424 (N_7424,N_634,N_1302);
or U7425 (N_7425,N_2683,N_1253);
nor U7426 (N_7426,N_2064,N_3732);
nand U7427 (N_7427,N_1773,N_1373);
or U7428 (N_7428,N_5131,N_2556);
xnor U7429 (N_7429,N_96,N_1938);
nand U7430 (N_7430,N_2865,N_1752);
nor U7431 (N_7431,N_5290,N_5888);
and U7432 (N_7432,N_4734,N_4666);
nand U7433 (N_7433,N_4582,N_802);
nor U7434 (N_7434,N_3726,N_4379);
xnor U7435 (N_7435,N_3656,N_1263);
nor U7436 (N_7436,N_2286,N_4530);
or U7437 (N_7437,N_5333,N_5708);
xor U7438 (N_7438,N_4094,N_5047);
nand U7439 (N_7439,N_5204,N_3145);
xnor U7440 (N_7440,N_4111,N_3780);
and U7441 (N_7441,N_3655,N_5430);
nand U7442 (N_7442,N_1669,N_2127);
or U7443 (N_7443,N_1519,N_1940);
or U7444 (N_7444,N_253,N_3125);
and U7445 (N_7445,N_129,N_4417);
or U7446 (N_7446,N_3065,N_2363);
or U7447 (N_7447,N_4132,N_3386);
and U7448 (N_7448,N_2824,N_213);
nor U7449 (N_7449,N_913,N_3794);
xor U7450 (N_7450,N_758,N_1908);
xor U7451 (N_7451,N_332,N_2868);
xor U7452 (N_7452,N_5642,N_60);
and U7453 (N_7453,N_2194,N_3362);
and U7454 (N_7454,N_4062,N_3052);
nor U7455 (N_7455,N_4397,N_1440);
and U7456 (N_7456,N_2830,N_2368);
nand U7457 (N_7457,N_2818,N_3680);
and U7458 (N_7458,N_3579,N_3385);
or U7459 (N_7459,N_931,N_5599);
or U7460 (N_7460,N_5066,N_3894);
nor U7461 (N_7461,N_23,N_4081);
or U7462 (N_7462,N_5238,N_2528);
xor U7463 (N_7463,N_314,N_3171);
and U7464 (N_7464,N_159,N_2329);
nand U7465 (N_7465,N_4176,N_3286);
nor U7466 (N_7466,N_5632,N_682);
or U7467 (N_7467,N_5136,N_2245);
or U7468 (N_7468,N_426,N_1184);
nand U7469 (N_7469,N_4085,N_1005);
xor U7470 (N_7470,N_1134,N_3940);
nor U7471 (N_7471,N_177,N_5745);
or U7472 (N_7472,N_5516,N_3466);
nand U7473 (N_7473,N_2442,N_2379);
or U7474 (N_7474,N_2947,N_167);
or U7475 (N_7475,N_3482,N_4179);
nand U7476 (N_7476,N_5021,N_1881);
nand U7477 (N_7477,N_1003,N_2690);
nor U7478 (N_7478,N_3138,N_5689);
nand U7479 (N_7479,N_1978,N_2325);
xnor U7480 (N_7480,N_4919,N_2233);
xnor U7481 (N_7481,N_4047,N_5184);
xor U7482 (N_7482,N_2810,N_4215);
and U7483 (N_7483,N_1888,N_2599);
nand U7484 (N_7484,N_3798,N_3593);
nand U7485 (N_7485,N_5166,N_3617);
nand U7486 (N_7486,N_887,N_4099);
or U7487 (N_7487,N_3461,N_3648);
or U7488 (N_7488,N_2589,N_103);
or U7489 (N_7489,N_551,N_5543);
nor U7490 (N_7490,N_629,N_2846);
nand U7491 (N_7491,N_3022,N_5086);
or U7492 (N_7492,N_5028,N_3783);
or U7493 (N_7493,N_1320,N_5107);
nand U7494 (N_7494,N_5519,N_5530);
xor U7495 (N_7495,N_2174,N_4296);
or U7496 (N_7496,N_348,N_3442);
and U7497 (N_7497,N_3796,N_3074);
nor U7498 (N_7498,N_255,N_2984);
nor U7499 (N_7499,N_3343,N_645);
nand U7500 (N_7500,N_4884,N_4730);
or U7501 (N_7501,N_1789,N_1667);
xnor U7502 (N_7502,N_5015,N_1579);
or U7503 (N_7503,N_1382,N_3347);
nand U7504 (N_7504,N_2693,N_3631);
xor U7505 (N_7505,N_1664,N_544);
and U7506 (N_7506,N_3309,N_5635);
nand U7507 (N_7507,N_5867,N_5692);
nor U7508 (N_7508,N_1629,N_5993);
nor U7509 (N_7509,N_112,N_3147);
and U7510 (N_7510,N_2148,N_5158);
nor U7511 (N_7511,N_2840,N_4559);
or U7512 (N_7512,N_3815,N_2225);
and U7513 (N_7513,N_396,N_2519);
and U7514 (N_7514,N_2621,N_4105);
xnor U7515 (N_7515,N_1275,N_3488);
nand U7516 (N_7516,N_2605,N_2128);
nand U7517 (N_7517,N_3294,N_3068);
nand U7518 (N_7518,N_4870,N_4607);
nand U7519 (N_7519,N_5217,N_214);
and U7520 (N_7520,N_4964,N_2701);
nor U7521 (N_7521,N_321,N_3400);
and U7522 (N_7522,N_1069,N_2123);
nand U7523 (N_7523,N_150,N_5085);
or U7524 (N_7524,N_1550,N_5402);
nor U7525 (N_7525,N_2301,N_578);
and U7526 (N_7526,N_1033,N_5773);
nor U7527 (N_7527,N_5707,N_5434);
or U7528 (N_7528,N_3415,N_4531);
xnor U7529 (N_7529,N_4001,N_3422);
and U7530 (N_7530,N_4936,N_3664);
nand U7531 (N_7531,N_1026,N_265);
xnor U7532 (N_7532,N_3932,N_5854);
and U7533 (N_7533,N_3937,N_3616);
nor U7534 (N_7534,N_2168,N_1103);
nor U7535 (N_7535,N_286,N_3445);
nand U7536 (N_7536,N_764,N_3533);
xor U7537 (N_7537,N_2974,N_5865);
xnor U7538 (N_7538,N_5074,N_5384);
or U7539 (N_7539,N_3216,N_3214);
xnor U7540 (N_7540,N_5715,N_3037);
nand U7541 (N_7541,N_4333,N_3419);
xnor U7542 (N_7542,N_4474,N_1146);
and U7543 (N_7543,N_42,N_1455);
and U7544 (N_7544,N_4721,N_1709);
or U7545 (N_7545,N_2996,N_811);
or U7546 (N_7546,N_3651,N_1958);
or U7547 (N_7547,N_1771,N_3610);
xnor U7548 (N_7548,N_3801,N_302);
nand U7549 (N_7549,N_2156,N_3803);
xor U7550 (N_7550,N_1858,N_3439);
nor U7551 (N_7551,N_4798,N_2544);
nor U7552 (N_7552,N_1615,N_5868);
and U7553 (N_7553,N_4174,N_69);
xor U7554 (N_7554,N_1883,N_1609);
xor U7555 (N_7555,N_5565,N_2337);
or U7556 (N_7556,N_5726,N_1849);
and U7557 (N_7557,N_2282,N_5641);
or U7558 (N_7558,N_4635,N_85);
and U7559 (N_7559,N_4019,N_422);
and U7560 (N_7560,N_4566,N_175);
and U7561 (N_7561,N_1357,N_2647);
nand U7562 (N_7562,N_1255,N_5416);
nor U7563 (N_7563,N_4548,N_3991);
nand U7564 (N_7564,N_5668,N_188);
or U7565 (N_7565,N_5121,N_808);
nand U7566 (N_7566,N_963,N_4126);
nand U7567 (N_7567,N_604,N_1312);
nand U7568 (N_7568,N_4563,N_816);
xor U7569 (N_7569,N_3830,N_3818);
nor U7570 (N_7570,N_2538,N_5357);
nor U7571 (N_7571,N_1230,N_1898);
and U7572 (N_7572,N_3047,N_2625);
nand U7573 (N_7573,N_4289,N_724);
or U7574 (N_7574,N_4362,N_1735);
or U7575 (N_7575,N_94,N_2741);
or U7576 (N_7576,N_3904,N_3895);
nand U7577 (N_7577,N_3865,N_591);
xnor U7578 (N_7578,N_4567,N_5104);
or U7579 (N_7579,N_1989,N_1157);
or U7580 (N_7580,N_1851,N_2181);
nor U7581 (N_7581,N_3401,N_1707);
and U7582 (N_7582,N_5946,N_2230);
nand U7583 (N_7583,N_5602,N_5190);
nor U7584 (N_7584,N_785,N_977);
or U7585 (N_7585,N_1812,N_4211);
xnor U7586 (N_7586,N_4986,N_5742);
xnor U7587 (N_7587,N_4210,N_3863);
nand U7588 (N_7588,N_4858,N_5925);
or U7589 (N_7589,N_2649,N_1260);
nand U7590 (N_7590,N_5600,N_3212);
nand U7591 (N_7591,N_1319,N_5377);
or U7592 (N_7592,N_4205,N_4323);
nor U7593 (N_7593,N_1159,N_1893);
xor U7594 (N_7594,N_3707,N_4023);
nand U7595 (N_7595,N_2048,N_1277);
nor U7596 (N_7596,N_2020,N_3180);
xor U7597 (N_7597,N_5433,N_1108);
or U7598 (N_7598,N_658,N_3239);
nand U7599 (N_7599,N_601,N_822);
xor U7600 (N_7600,N_31,N_3787);
and U7601 (N_7601,N_1991,N_3200);
nand U7602 (N_7602,N_1823,N_2210);
and U7603 (N_7603,N_5195,N_1403);
xor U7604 (N_7604,N_5739,N_1558);
nand U7605 (N_7605,N_3852,N_4887);
and U7606 (N_7606,N_3953,N_113);
nand U7607 (N_7607,N_258,N_4980);
nand U7608 (N_7608,N_3072,N_1190);
xnor U7609 (N_7609,N_4150,N_1336);
nor U7610 (N_7610,N_554,N_3280);
nand U7611 (N_7611,N_2054,N_136);
and U7612 (N_7612,N_4544,N_2793);
or U7613 (N_7613,N_1393,N_5317);
nand U7614 (N_7614,N_4855,N_4502);
and U7615 (N_7615,N_2501,N_4755);
or U7616 (N_7616,N_5468,N_2747);
xor U7617 (N_7617,N_305,N_4165);
nor U7618 (N_7618,N_463,N_5185);
nor U7619 (N_7619,N_5630,N_2159);
or U7620 (N_7620,N_4835,N_5205);
nand U7621 (N_7621,N_2653,N_1050);
nor U7622 (N_7622,N_4768,N_2943);
xnor U7623 (N_7623,N_1172,N_271);
or U7624 (N_7624,N_4861,N_1937);
xnor U7625 (N_7625,N_1931,N_5682);
nand U7626 (N_7626,N_4829,N_71);
nand U7627 (N_7627,N_1349,N_4240);
or U7628 (N_7628,N_5895,N_3717);
and U7629 (N_7629,N_2216,N_146);
and U7630 (N_7630,N_1819,N_191);
or U7631 (N_7631,N_1009,N_3192);
or U7632 (N_7632,N_4627,N_2274);
nor U7633 (N_7633,N_1427,N_683);
nand U7634 (N_7634,N_1314,N_4341);
nand U7635 (N_7635,N_1021,N_1557);
nand U7636 (N_7636,N_3586,N_2038);
or U7637 (N_7637,N_2017,N_2601);
or U7638 (N_7638,N_3952,N_1479);
and U7639 (N_7639,N_4,N_1694);
or U7640 (N_7640,N_946,N_4063);
xor U7641 (N_7641,N_5071,N_5168);
nor U7642 (N_7642,N_4632,N_5894);
and U7643 (N_7643,N_723,N_30);
xor U7644 (N_7644,N_643,N_2985);
nor U7645 (N_7645,N_1361,N_4593);
nand U7646 (N_7646,N_3710,N_5216);
xor U7647 (N_7647,N_844,N_2584);
xnor U7648 (N_7648,N_5789,N_1637);
and U7649 (N_7649,N_3957,N_3898);
nand U7650 (N_7650,N_1359,N_1963);
and U7651 (N_7651,N_4102,N_5297);
and U7652 (N_7652,N_397,N_5495);
xnor U7653 (N_7653,N_2565,N_1738);
or U7654 (N_7654,N_3525,N_4212);
xor U7655 (N_7655,N_3566,N_2648);
nand U7656 (N_7656,N_4228,N_1754);
xor U7657 (N_7657,N_1914,N_3826);
and U7658 (N_7658,N_2608,N_4222);
and U7659 (N_7659,N_3040,N_1982);
or U7660 (N_7660,N_5072,N_5420);
nand U7661 (N_7661,N_2498,N_2590);
and U7662 (N_7662,N_3835,N_3083);
nand U7663 (N_7663,N_266,N_3985);
xnor U7664 (N_7664,N_359,N_3007);
xnor U7665 (N_7665,N_2477,N_3018);
nor U7666 (N_7666,N_4028,N_5350);
nand U7667 (N_7667,N_3702,N_2117);
nor U7668 (N_7668,N_4410,N_2534);
nor U7669 (N_7669,N_5192,N_5539);
nand U7670 (N_7670,N_2319,N_4891);
nor U7671 (N_7671,N_2756,N_695);
xnor U7672 (N_7672,N_4146,N_1730);
or U7673 (N_7673,N_5114,N_2958);
or U7674 (N_7674,N_5505,N_2807);
nand U7675 (N_7675,N_1821,N_3550);
or U7676 (N_7676,N_2075,N_4823);
or U7677 (N_7677,N_5847,N_3242);
nand U7678 (N_7678,N_5944,N_2686);
nor U7679 (N_7679,N_891,N_1806);
and U7680 (N_7680,N_2631,N_840);
xnor U7681 (N_7681,N_2229,N_2299);
and U7682 (N_7682,N_3641,N_896);
nand U7683 (N_7683,N_2142,N_2954);
nor U7684 (N_7684,N_1533,N_531);
xnor U7685 (N_7685,N_690,N_2440);
and U7686 (N_7686,N_2520,N_67);
and U7687 (N_7687,N_2994,N_4166);
nand U7688 (N_7688,N_1997,N_3867);
or U7689 (N_7689,N_5960,N_5315);
nor U7690 (N_7690,N_5151,N_1451);
or U7691 (N_7691,N_2674,N_2717);
or U7692 (N_7692,N_4266,N_36);
nand U7693 (N_7693,N_1547,N_1890);
or U7694 (N_7694,N_5258,N_3346);
nand U7695 (N_7695,N_1369,N_4517);
nand U7696 (N_7696,N_4121,N_1702);
and U7697 (N_7697,N_1281,N_1004);
xor U7698 (N_7698,N_5075,N_2261);
xnor U7699 (N_7699,N_3854,N_1595);
or U7700 (N_7700,N_5211,N_5478);
nor U7701 (N_7701,N_2172,N_3049);
or U7702 (N_7702,N_5144,N_1841);
xor U7703 (N_7703,N_1345,N_3430);
nor U7704 (N_7704,N_5474,N_5757);
or U7705 (N_7705,N_2927,N_1950);
or U7706 (N_7706,N_3745,N_5231);
or U7707 (N_7707,N_4623,N_1154);
nand U7708 (N_7708,N_5651,N_4827);
or U7709 (N_7709,N_2431,N_1222);
or U7710 (N_7710,N_2782,N_2788);
nor U7711 (N_7711,N_2221,N_5978);
and U7712 (N_7712,N_3248,N_3435);
nand U7713 (N_7713,N_4059,N_5054);
and U7714 (N_7714,N_5943,N_4230);
or U7715 (N_7715,N_906,N_5115);
nand U7716 (N_7716,N_403,N_1659);
or U7717 (N_7717,N_5698,N_4482);
and U7718 (N_7718,N_1286,N_1910);
nand U7719 (N_7719,N_3935,N_5667);
and U7720 (N_7720,N_2970,N_3474);
or U7721 (N_7721,N_3762,N_4428);
and U7722 (N_7722,N_3570,N_5340);
nor U7723 (N_7723,N_1840,N_1522);
and U7724 (N_7724,N_4029,N_3188);
xnor U7725 (N_7725,N_2112,N_2195);
nor U7726 (N_7726,N_2311,N_417);
nor U7727 (N_7727,N_1463,N_2571);
xnor U7728 (N_7728,N_4718,N_2890);
nand U7729 (N_7729,N_1208,N_1985);
xor U7730 (N_7730,N_2924,N_1662);
xnor U7731 (N_7731,N_1512,N_4513);
and U7732 (N_7732,N_2508,N_3503);
xor U7733 (N_7733,N_3978,N_5687);
or U7734 (N_7734,N_4057,N_618);
nor U7735 (N_7735,N_748,N_4564);
xor U7736 (N_7736,N_3591,N_2658);
xor U7737 (N_7737,N_4630,N_5277);
or U7738 (N_7738,N_5335,N_5629);
and U7739 (N_7739,N_3066,N_3497);
and U7740 (N_7740,N_708,N_5917);
nand U7741 (N_7741,N_4177,N_539);
nor U7742 (N_7742,N_487,N_4486);
nand U7743 (N_7743,N_5537,N_2079);
nor U7744 (N_7744,N_1348,N_5620);
nand U7745 (N_7745,N_573,N_5844);
xnor U7746 (N_7746,N_4585,N_127);
and U7747 (N_7747,N_3845,N_3751);
nand U7748 (N_7748,N_2516,N_3876);
xnor U7749 (N_7749,N_2712,N_5814);
nor U7750 (N_7750,N_4273,N_2973);
nor U7751 (N_7751,N_5512,N_446);
nand U7752 (N_7752,N_2836,N_4606);
or U7753 (N_7753,N_5903,N_2087);
nand U7754 (N_7754,N_2945,N_4663);
nor U7755 (N_7755,N_2841,N_1104);
or U7756 (N_7756,N_5897,N_5318);
xor U7757 (N_7757,N_3560,N_4904);
nor U7758 (N_7758,N_4863,N_4832);
nand U7759 (N_7759,N_5289,N_5355);
nor U7760 (N_7760,N_4002,N_2547);
nor U7761 (N_7761,N_230,N_5705);
nor U7762 (N_7762,N_3130,N_1772);
nor U7763 (N_7763,N_647,N_5173);
xnor U7764 (N_7764,N_3979,N_3394);
and U7765 (N_7765,N_1396,N_3584);
and U7766 (N_7766,N_5177,N_4285);
or U7767 (N_7767,N_990,N_4036);
nand U7768 (N_7768,N_1497,N_1942);
nor U7769 (N_7769,N_3572,N_2113);
and U7770 (N_7770,N_5799,N_2705);
nand U7771 (N_7771,N_5400,N_3070);
xnor U7772 (N_7772,N_4426,N_4852);
xnor U7773 (N_7773,N_1715,N_4109);
or U7774 (N_7774,N_3298,N_2808);
nor U7775 (N_7775,N_3307,N_5022);
nor U7776 (N_7776,N_5560,N_2202);
xor U7777 (N_7777,N_641,N_5023);
and U7778 (N_7778,N_1928,N_1904);
and U7779 (N_7779,N_2735,N_179);
xor U7780 (N_7780,N_3455,N_5927);
and U7781 (N_7781,N_1080,N_453);
nand U7782 (N_7782,N_4569,N_3665);
nor U7783 (N_7783,N_2626,N_5919);
nand U7784 (N_7784,N_4619,N_3575);
nand U7785 (N_7785,N_1379,N_3673);
nand U7786 (N_7786,N_1632,N_3618);
nand U7787 (N_7787,N_2536,N_3567);
nand U7788 (N_7788,N_5748,N_1571);
nand U7789 (N_7789,N_1979,N_380);
and U7790 (N_7790,N_832,N_3191);
or U7791 (N_7791,N_4545,N_5820);
nor U7792 (N_7792,N_2439,N_4670);
and U7793 (N_7793,N_1649,N_3186);
xnor U7794 (N_7794,N_2799,N_4162);
and U7795 (N_7795,N_2395,N_3056);
nand U7796 (N_7796,N_5492,N_3182);
and U7797 (N_7797,N_3743,N_2497);
and U7798 (N_7798,N_1466,N_2346);
and U7799 (N_7799,N_1368,N_4226);
xnor U7800 (N_7800,N_5811,N_5973);
or U7801 (N_7801,N_3805,N_3674);
nor U7802 (N_7802,N_5033,N_5499);
or U7803 (N_7803,N_614,N_1518);
and U7804 (N_7804,N_4377,N_4525);
xnor U7805 (N_7805,N_1282,N_374);
or U7806 (N_7806,N_2264,N_2235);
xnor U7807 (N_7807,N_1229,N_3421);
nand U7808 (N_7808,N_2406,N_1506);
or U7809 (N_7809,N_3224,N_5447);
and U7810 (N_7810,N_3206,N_4648);
xor U7811 (N_7811,N_4703,N_412);
and U7812 (N_7812,N_1998,N_4813);
nor U7813 (N_7813,N_5065,N_3646);
or U7814 (N_7814,N_442,N_4782);
xor U7815 (N_7815,N_4317,N_3027);
xnor U7816 (N_7816,N_2517,N_4945);
or U7817 (N_7817,N_2147,N_25);
xor U7818 (N_7818,N_5886,N_1645);
nand U7819 (N_7819,N_5833,N_1041);
and U7820 (N_7820,N_1491,N_3059);
or U7821 (N_7821,N_1727,N_5097);
nor U7822 (N_7822,N_5992,N_1889);
and U7823 (N_7823,N_3398,N_5690);
xnor U7824 (N_7824,N_926,N_4587);
nor U7825 (N_7825,N_930,N_4620);
nor U7826 (N_7826,N_3982,N_4476);
xor U7827 (N_7827,N_501,N_3468);
xor U7828 (N_7828,N_1114,N_3922);
nand U7829 (N_7829,N_5966,N_5365);
nand U7830 (N_7830,N_1544,N_5304);
and U7831 (N_7831,N_264,N_4911);
xor U7832 (N_7832,N_3326,N_665);
and U7833 (N_7833,N_3713,N_4636);
or U7834 (N_7834,N_2518,N_5535);
and U7835 (N_7835,N_1603,N_5403);
nand U7836 (N_7836,N_5699,N_1030);
and U7837 (N_7837,N_1969,N_5538);
nand U7838 (N_7838,N_3597,N_1432);
nand U7839 (N_7839,N_43,N_5079);
xnor U7840 (N_7840,N_1878,N_4292);
or U7841 (N_7841,N_538,N_4331);
xor U7842 (N_7842,N_3869,N_1067);
nand U7843 (N_7843,N_4390,N_5016);
or U7844 (N_7844,N_3987,N_3603);
or U7845 (N_7845,N_4274,N_48);
nand U7846 (N_7846,N_1072,N_2472);
and U7847 (N_7847,N_70,N_1453);
and U7848 (N_7848,N_3312,N_5300);
and U7849 (N_7849,N_3962,N_3727);
xnor U7850 (N_7850,N_650,N_2313);
and U7851 (N_7851,N_2645,N_1845);
or U7852 (N_7852,N_3255,N_2630);
xor U7853 (N_7853,N_4320,N_238);
nor U7854 (N_7854,N_5371,N_3470);
and U7855 (N_7855,N_1323,N_5968);
or U7856 (N_7856,N_4715,N_2545);
or U7857 (N_7857,N_3974,N_4198);
xnor U7858 (N_7858,N_3050,N_4046);
or U7859 (N_7859,N_534,N_3719);
nand U7860 (N_7860,N_5850,N_3020);
nand U7861 (N_7861,N_4806,N_5772);
and U7862 (N_7862,N_3943,N_5794);
and U7863 (N_7863,N_5476,N_5262);
or U7864 (N_7864,N_5634,N_481);
xnor U7865 (N_7865,N_5421,N_330);
xnor U7866 (N_7866,N_1882,N_5892);
nor U7867 (N_7867,N_3264,N_5942);
nor U7868 (N_7868,N_4357,N_3115);
or U7869 (N_7869,N_4406,N_1716);
and U7870 (N_7870,N_3376,N_1018);
nor U7871 (N_7871,N_1748,N_5666);
nand U7872 (N_7872,N_4031,N_5119);
or U7873 (N_7873,N_1742,N_2895);
and U7874 (N_7874,N_4710,N_1446);
nor U7875 (N_7875,N_4524,N_2411);
and U7876 (N_7876,N_4196,N_2208);
nor U7877 (N_7877,N_334,N_1570);
or U7878 (N_7878,N_3128,N_592);
or U7879 (N_7879,N_5645,N_941);
or U7880 (N_7880,N_5937,N_820);
or U7881 (N_7881,N_2408,N_441);
and U7882 (N_7882,N_3812,N_5728);
or U7883 (N_7883,N_5465,N_141);
nor U7884 (N_7884,N_4115,N_77);
nor U7885 (N_7885,N_969,N_897);
nor U7886 (N_7886,N_3545,N_1852);
or U7887 (N_7887,N_5302,N_2050);
or U7888 (N_7888,N_3883,N_2223);
or U7889 (N_7889,N_1697,N_4311);
nor U7890 (N_7890,N_2704,N_440);
or U7891 (N_7891,N_1029,N_4756);
nand U7892 (N_7892,N_5175,N_303);
or U7893 (N_7893,N_2512,N_4130);
xnor U7894 (N_7894,N_944,N_5838);
nor U7895 (N_7895,N_702,N_1163);
nor U7896 (N_7896,N_2531,N_4042);
nor U7897 (N_7897,N_2906,N_1917);
xor U7898 (N_7898,N_613,N_1426);
and U7899 (N_7899,N_5133,N_5274);
xor U7900 (N_7900,N_3650,N_751);
and U7901 (N_7901,N_5321,N_3262);
nand U7902 (N_7902,N_4882,N_4752);
xor U7903 (N_7903,N_1496,N_631);
nand U7904 (N_7904,N_1555,N_5988);
and U7905 (N_7905,N_4797,N_5491);
and U7906 (N_7906,N_5343,N_2981);
xor U7907 (N_7907,N_2088,N_5590);
xor U7908 (N_7908,N_5004,N_864);
and U7909 (N_7909,N_4248,N_2677);
and U7910 (N_7910,N_5542,N_2170);
xor U7911 (N_7911,N_1617,N_3327);
or U7912 (N_7912,N_105,N_5143);
xnor U7913 (N_7913,N_5719,N_358);
nand U7914 (N_7914,N_3073,N_3498);
or U7915 (N_7915,N_1084,N_1153);
xor U7916 (N_7916,N_5725,N_4018);
or U7917 (N_7917,N_2263,N_2751);
xor U7918 (N_7918,N_1304,N_2260);
xnor U7919 (N_7919,N_547,N_4454);
nor U7920 (N_7920,N_1467,N_3240);
xnor U7921 (N_7921,N_3931,N_1503);
and U7922 (N_7922,N_4416,N_2784);
xor U7923 (N_7923,N_5553,N_2992);
and U7924 (N_7924,N_1461,N_5171);
or U7925 (N_7925,N_3063,N_606);
nand U7926 (N_7926,N_1674,N_3817);
xnor U7927 (N_7927,N_4246,N_4842);
and U7928 (N_7928,N_3153,N_824);
xnor U7929 (N_7929,N_4661,N_5278);
xor U7930 (N_7930,N_2874,N_3094);
nand U7931 (N_7931,N_211,N_364);
nor U7932 (N_7932,N_3017,N_4175);
nor U7933 (N_7933,N_4217,N_2582);
and U7934 (N_7934,N_701,N_3024);
and U7935 (N_7935,N_1217,N_3938);
or U7936 (N_7936,N_5713,N_4667);
nor U7937 (N_7937,N_4455,N_1384);
xor U7938 (N_7938,N_4690,N_776);
and U7939 (N_7939,N_5762,N_5876);
xnor U7940 (N_7940,N_4848,N_5890);
or U7941 (N_7941,N_2780,N_3678);
or U7942 (N_7942,N_533,N_1449);
nand U7943 (N_7943,N_1127,N_1633);
nand U7944 (N_7944,N_11,N_5637);
or U7945 (N_7945,N_1585,N_1546);
xnor U7946 (N_7946,N_1151,N_2514);
nand U7947 (N_7947,N_574,N_3290);
nand U7948 (N_7948,N_1783,N_2326);
xnor U7949 (N_7949,N_1341,N_4298);
or U7950 (N_7950,N_3373,N_850);
xnor U7951 (N_7951,N_4973,N_593);
and U7952 (N_7952,N_2198,N_1955);
xnor U7953 (N_7953,N_4097,N_2706);
and U7954 (N_7954,N_3667,N_4456);
and U7955 (N_7955,N_2340,N_194);
nor U7956 (N_7956,N_3846,N_5427);
xor U7957 (N_7957,N_3038,N_932);
nor U7958 (N_7958,N_4883,N_5224);
or U7959 (N_7959,N_5448,N_935);
nand U7960 (N_7960,N_4976,N_1769);
nand U7961 (N_7961,N_480,N_4597);
and U7962 (N_7962,N_5873,N_693);
xor U7963 (N_7963,N_2911,N_3748);
nand U7964 (N_7964,N_532,N_5796);
or U7965 (N_7965,N_121,N_3377);
or U7966 (N_7966,N_649,N_1793);
or U7967 (N_7967,N_3078,N_4280);
nor U7968 (N_7968,N_4264,N_2347);
nor U7969 (N_7969,N_205,N_3273);
and U7970 (N_7970,N_862,N_1476);
or U7971 (N_7971,N_1513,N_1092);
nor U7972 (N_7972,N_2802,N_3277);
nor U7973 (N_7973,N_485,N_386);
xnor U7974 (N_7974,N_5675,N_5445);
nor U7975 (N_7975,N_3203,N_5298);
or U7976 (N_7976,N_3352,N_5947);
or U7977 (N_7977,N_2785,N_2627);
xnor U7978 (N_7978,N_5697,N_3261);
xor U7979 (N_7979,N_4951,N_4795);
and U7980 (N_7980,N_172,N_1370);
nor U7981 (N_7981,N_2446,N_5183);
and U7982 (N_7982,N_4030,N_3330);
and U7983 (N_7983,N_3081,N_3740);
or U7984 (N_7984,N_5354,N_5616);
nor U7985 (N_7985,N_775,N_5922);
or U7986 (N_7986,N_1717,N_4282);
or U7987 (N_7987,N_959,N_62);
nor U7988 (N_7988,N_217,N_5152);
xnor U7989 (N_7989,N_5011,N_4348);
nor U7990 (N_7990,N_3834,N_1248);
nand U7991 (N_7991,N_5801,N_536);
xnor U7992 (N_7992,N_1316,N_4190);
xnor U7993 (N_7993,N_4496,N_3489);
or U7994 (N_7994,N_4490,N_3723);
or U7995 (N_7995,N_2870,N_1666);
xnor U7996 (N_7996,N_2047,N_5490);
nor U7997 (N_7997,N_3781,N_3686);
nor U7998 (N_7998,N_5755,N_3031);
nor U7999 (N_7999,N_2572,N_365);
nand U8000 (N_8000,N_4022,N_5866);
and U8001 (N_8001,N_3291,N_2764);
xor U8002 (N_8002,N_2963,N_5444);
xor U8003 (N_8003,N_13,N_5859);
xnor U8004 (N_8004,N_2470,N_5459);
nor U8005 (N_8005,N_3639,N_1071);
nand U8006 (N_8006,N_4714,N_2310);
nand U8007 (N_8007,N_557,N_3345);
nor U8008 (N_8008,N_3016,N_306);
nand U8009 (N_8009,N_1308,N_2620);
and U8010 (N_8010,N_620,N_2877);
nor U8011 (N_8011,N_5411,N_2104);
nor U8012 (N_8012,N_4479,N_3055);
and U8013 (N_8013,N_4149,N_2126);
and U8014 (N_8014,N_1062,N_108);
and U8015 (N_8015,N_4780,N_1125);
nand U8016 (N_8016,N_449,N_4615);
xnor U8017 (N_8017,N_357,N_1835);
and U8018 (N_8018,N_798,N_5109);
or U8019 (N_8019,N_4985,N_144);
and U8020 (N_8020,N_484,N_2450);
nor U8021 (N_8021,N_4446,N_4394);
xnor U8022 (N_8022,N_2359,N_1693);
xnor U8023 (N_8023,N_739,N_1757);
or U8024 (N_8024,N_5822,N_2430);
nand U8025 (N_8025,N_5853,N_2120);
and U8026 (N_8026,N_4433,N_4692);
nor U8027 (N_8027,N_5920,N_145);
and U8028 (N_8028,N_1808,N_1048);
or U8029 (N_8029,N_3389,N_5052);
or U8030 (N_8030,N_2929,N_4318);
or U8031 (N_8031,N_5426,N_296);
nand U8032 (N_8032,N_3113,N_1223);
or U8033 (N_8033,N_3878,N_5683);
or U8034 (N_8034,N_4996,N_2925);
nor U8035 (N_8035,N_3303,N_651);
nor U8036 (N_8036,N_5453,N_3101);
xnor U8037 (N_8037,N_1117,N_561);
and U8038 (N_8038,N_4783,N_581);
and U8039 (N_8039,N_5415,N_4561);
and U8040 (N_8040,N_874,N_4591);
nand U8041 (N_8041,N_3823,N_3029);
nor U8042 (N_8042,N_5117,N_5134);
nand U8043 (N_8043,N_4450,N_1532);
or U8044 (N_8044,N_540,N_5000);
xor U8045 (N_8045,N_4251,N_5702);
nor U8046 (N_8046,N_4551,N_4785);
xor U8047 (N_8047,N_5271,N_1584);
and U8048 (N_8048,N_1441,N_603);
nand U8049 (N_8049,N_3162,N_2676);
xor U8050 (N_8050,N_5061,N_2306);
nand U8051 (N_8051,N_5069,N_66);
or U8052 (N_8052,N_5209,N_119);
nand U8053 (N_8053,N_4992,N_1832);
or U8054 (N_8054,N_309,N_5502);
xnor U8055 (N_8055,N_4010,N_856);
nor U8056 (N_8056,N_1177,N_1954);
xnor U8057 (N_8057,N_2102,N_2510);
nand U8058 (N_8058,N_1421,N_2796);
or U8059 (N_8059,N_805,N_3028);
and U8060 (N_8060,N_4484,N_2850);
nor U8061 (N_8061,N_3602,N_3501);
and U8062 (N_8062,N_3392,N_1536);
or U8063 (N_8063,N_3393,N_5513);
nand U8064 (N_8064,N_3025,N_4896);
xnor U8065 (N_8065,N_4395,N_171);
nand U8066 (N_8066,N_5057,N_4844);
and U8067 (N_8067,N_526,N_2094);
xnor U8068 (N_8068,N_3691,N_3622);
or U8069 (N_8069,N_2696,N_3134);
or U8070 (N_8070,N_5095,N_722);
nand U8071 (N_8071,N_2763,N_5222);
xor U8072 (N_8072,N_5194,N_4260);
nor U8073 (N_8073,N_4338,N_2946);
xor U8074 (N_8074,N_2466,N_5613);
and U8075 (N_8075,N_4981,N_5129);
and U8076 (N_8076,N_44,N_2399);
nand U8077 (N_8077,N_3733,N_3833);
nand U8078 (N_8078,N_5918,N_2853);
nor U8079 (N_8079,N_838,N_3281);
nand U8080 (N_8080,N_3630,N_4645);
or U8081 (N_8081,N_2922,N_5410);
nor U8082 (N_8082,N_3151,N_135);
nand U8083 (N_8083,N_4761,N_3405);
nand U8084 (N_8084,N_2482,N_3438);
or U8085 (N_8085,N_4660,N_568);
and U8086 (N_8086,N_4319,N_231);
or U8087 (N_8087,N_4430,N_1342);
and U8088 (N_8088,N_918,N_2484);
xor U8089 (N_8089,N_2819,N_5549);
nand U8090 (N_8090,N_1065,N_5830);
xor U8091 (N_8091,N_2055,N_1778);
nand U8092 (N_8092,N_4003,N_3479);
and U8093 (N_8093,N_3295,N_5904);
and U8094 (N_8094,N_5339,N_5584);
nor U8095 (N_8095,N_624,N_3642);
or U8096 (N_8096,N_5208,N_4598);
xor U8097 (N_8097,N_792,N_3267);
and U8098 (N_8098,N_4909,N_1527);
and U8099 (N_8099,N_2641,N_2760);
xnor U8100 (N_8100,N_1941,N_773);
and U8101 (N_8101,N_4011,N_3087);
or U8102 (N_8102,N_552,N_2755);
and U8103 (N_8103,N_5149,N_4754);
or U8104 (N_8104,N_5078,N_49);
nor U8105 (N_8105,N_5203,N_4510);
or U8106 (N_8106,N_1126,N_4448);
xnor U8107 (N_8107,N_3516,N_1034);
and U8108 (N_8108,N_5252,N_5206);
xnor U8109 (N_8109,N_4127,N_596);
and U8110 (N_8110,N_4227,N_3968);
xnor U8111 (N_8111,N_2412,N_625);
xor U8112 (N_8112,N_4971,N_1075);
and U8113 (N_8113,N_5841,N_4968);
xor U8114 (N_8114,N_4947,N_1591);
and U8115 (N_8115,N_1465,N_1871);
and U8116 (N_8116,N_3133,N_2275);
nand U8117 (N_8117,N_3942,N_384);
and U8118 (N_8118,N_3882,N_4726);
or U8119 (N_8119,N_4769,N_550);
nor U8120 (N_8120,N_2111,N_2614);
nand U8121 (N_8121,N_2175,N_710);
and U8122 (N_8122,N_479,N_3936);
and U8123 (N_8123,N_709,N_2242);
nand U8124 (N_8124,N_1753,N_166);
or U8125 (N_8125,N_3390,N_5454);
xor U8126 (N_8126,N_4650,N_5191);
nor U8127 (N_8127,N_5487,N_5314);
or U8128 (N_8128,N_1372,N_3351);
or U8129 (N_8129,N_2273,N_4156);
xnor U8130 (N_8130,N_513,N_5360);
and U8131 (N_8131,N_3712,N_3578);
nor U8132 (N_8132,N_2618,N_1805);
nand U8133 (N_8133,N_1433,N_3061);
nor U8134 (N_8134,N_257,N_514);
nor U8135 (N_8135,N_118,N_5092);
nand U8136 (N_8136,N_5819,N_678);
xor U8137 (N_8137,N_4239,N_5405);
or U8138 (N_8138,N_3154,N_2639);
or U8139 (N_8139,N_2160,N_3784);
and U8140 (N_8140,N_3353,N_3416);
and U8141 (N_8141,N_1181,N_2600);
or U8142 (N_8142,N_5688,N_3414);
nor U8143 (N_8143,N_1383,N_3917);
or U8144 (N_8144,N_3365,N_3688);
and U8145 (N_8145,N_5931,N_2296);
nor U8146 (N_8146,N_1844,N_3929);
nor U8147 (N_8147,N_1053,N_2370);
or U8148 (N_8148,N_5963,N_5053);
nor U8149 (N_8149,N_2091,N_3534);
nor U8150 (N_8150,N_3388,N_638);
and U8151 (N_8151,N_1775,N_3820);
or U8152 (N_8152,N_1896,N_2697);
and U8153 (N_8153,N_911,N_5275);
nor U8154 (N_8154,N_1762,N_3491);
or U8155 (N_8155,N_3951,N_2800);
and U8156 (N_8156,N_2285,N_5658);
and U8157 (N_8157,N_4027,N_662);
nand U8158 (N_8158,N_3679,N_1161);
nor U8159 (N_8159,N_5900,N_2036);
nand U8160 (N_8160,N_154,N_2679);
nand U8161 (N_8161,N_2131,N_1873);
nor U8162 (N_8162,N_3822,N_2014);
xnor U8163 (N_8163,N_1731,N_1055);
nor U8164 (N_8164,N_1305,N_1101);
xor U8165 (N_8165,N_878,N_4800);
nand U8166 (N_8166,N_203,N_1490);
nor U8167 (N_8167,N_301,N_4862);
nand U8168 (N_8168,N_3011,N_4310);
nand U8169 (N_8169,N_1724,N_3568);
and U8170 (N_8170,N_5882,N_2448);
xor U8171 (N_8171,N_3382,N_5509);
nand U8172 (N_8172,N_4540,N_4384);
nand U8173 (N_8173,N_1639,N_1083);
xor U8174 (N_8174,N_5181,N_333);
and U8175 (N_8175,N_178,N_2360);
and U8176 (N_8176,N_1480,N_4457);
and U8177 (N_8177,N_5852,N_5770);
nor U8178 (N_8178,N_5800,N_5598);
xnor U8179 (N_8179,N_4817,N_1507);
xor U8180 (N_8180,N_837,N_5089);
and U8181 (N_8181,N_5249,N_4745);
nor U8182 (N_8182,N_530,N_1107);
xnor U8183 (N_8183,N_1130,N_2543);
or U8184 (N_8184,N_458,N_1660);
xnor U8185 (N_8185,N_226,N_4374);
nor U8186 (N_8186,N_5774,N_61);
or U8187 (N_8187,N_2532,N_5048);
nor U8188 (N_8188,N_5955,N_2682);
and U8189 (N_8189,N_4034,N_2791);
and U8190 (N_8190,N_5735,N_4441);
xnor U8191 (N_8191,N_4089,N_2767);
and U8192 (N_8192,N_5723,N_1797);
xor U8193 (N_8193,N_1244,N_5738);
and U8194 (N_8194,N_1876,N_2775);
or U8195 (N_8195,N_2952,N_1087);
xnor U8196 (N_8196,N_3339,N_1469);
and U8197 (N_8197,N_1880,N_3190);
or U8198 (N_8198,N_2743,N_4792);
and U8199 (N_8199,N_4617,N_447);
nor U8200 (N_8200,N_5164,N_1144);
and U8201 (N_8201,N_4836,N_3853);
nand U8202 (N_8202,N_4182,N_55);
nor U8203 (N_8203,N_3829,N_652);
nand U8204 (N_8204,N_880,N_2062);
xnor U8205 (N_8205,N_2386,N_4138);
nor U8206 (N_8206,N_2950,N_1085);
or U8207 (N_8207,N_5170,N_704);
or U8208 (N_8208,N_1292,N_3995);
or U8209 (N_8209,N_4628,N_227);
nor U8210 (N_8210,N_3064,N_644);
nor U8211 (N_8211,N_3476,N_529);
and U8212 (N_8212,N_3253,N_3372);
and U8213 (N_8213,N_2820,N_1169);
xor U8214 (N_8214,N_5261,N_2816);
xor U8215 (N_8215,N_399,N_4025);
and U8216 (N_8216,N_4278,N_586);
and U8217 (N_8217,N_2255,N_998);
or U8218 (N_8218,N_152,N_109);
nor U8219 (N_8219,N_2410,N_4128);
xor U8220 (N_8220,N_2397,N_4706);
xnor U8221 (N_8221,N_1899,N_3615);
and U8222 (N_8222,N_3627,N_318);
or U8223 (N_8223,N_993,N_1091);
or U8224 (N_8224,N_336,N_5142);
nor U8225 (N_8225,N_985,N_5752);
or U8226 (N_8226,N_3102,N_5325);
xnor U8227 (N_8227,N_1628,N_2246);
or U8228 (N_8228,N_5609,N_4914);
and U8229 (N_8229,N_128,N_4654);
xnor U8230 (N_8230,N_5607,N_2632);
or U8231 (N_8231,N_5884,N_3543);
or U8232 (N_8232,N_3759,N_1824);
nand U8233 (N_8233,N_3100,N_3201);
and U8234 (N_8234,N_294,N_1962);
nand U8235 (N_8235,N_3739,N_884);
and U8236 (N_8236,N_4532,N_1274);
or U8237 (N_8237,N_2268,N_360);
nor U8238 (N_8238,N_4686,N_2831);
xor U8239 (N_8239,N_1764,N_842);
nor U8240 (N_8240,N_3431,N_1839);
xor U8241 (N_8241,N_1990,N_5898);
xor U8242 (N_8242,N_4079,N_3428);
or U8243 (N_8243,N_5467,N_2429);
nor U8244 (N_8244,N_1792,N_1363);
and U8245 (N_8245,N_2392,N_2896);
and U8246 (N_8246,N_1266,N_3980);
xor U8247 (N_8247,N_5040,N_585);
nand U8248 (N_8248,N_3636,N_3229);
nand U8249 (N_8249,N_2342,N_7);
nand U8250 (N_8250,N_5681,N_657);
xnor U8251 (N_8251,N_2928,N_12);
nand U8252 (N_8252,N_1182,N_5506);
xor U8253 (N_8253,N_5572,N_4418);
and U8254 (N_8254,N_2522,N_2983);
or U8255 (N_8255,N_4224,N_2662);
or U8256 (N_8256,N_2333,N_5508);
xnor U8257 (N_8257,N_5754,N_4900);
xor U8258 (N_8258,N_1658,N_1265);
nor U8259 (N_8259,N_4750,N_1944);
nand U8260 (N_8260,N_349,N_1921);
nand U8261 (N_8261,N_1149,N_2099);
nand U8262 (N_8262,N_5425,N_5373);
xor U8263 (N_8263,N_1023,N_3370);
xnor U8264 (N_8264,N_4841,N_987);
and U8265 (N_8265,N_4618,N_999);
or U8266 (N_8266,N_2180,N_1563);
nor U8267 (N_8267,N_1110,N_4075);
or U8268 (N_8268,N_5521,N_2982);
nor U8269 (N_8269,N_3170,N_2490);
and U8270 (N_8270,N_429,N_5514);
nor U8271 (N_8271,N_2300,N_5517);
nor U8272 (N_8272,N_260,N_712);
and U8273 (N_8273,N_4124,N_835);
or U8274 (N_8274,N_3559,N_5088);
and U8275 (N_8275,N_2607,N_1462);
xor U8276 (N_8276,N_4940,N_304);
xor U8277 (N_8277,N_736,N_133);
and U8278 (N_8278,N_809,N_2437);
nand U8279 (N_8279,N_3596,N_3816);
xnor U8280 (N_8280,N_5891,N_1297);
nand U8281 (N_8281,N_438,N_5786);
or U8282 (N_8282,N_3546,N_2750);
xor U8283 (N_8283,N_4193,N_3967);
nand U8284 (N_8284,N_3776,N_2733);
and U8285 (N_8285,N_3728,N_1995);
nand U8286 (N_8286,N_546,N_4676);
nor U8287 (N_8287,N_668,N_5997);
or U8288 (N_8288,N_1200,N_288);
nand U8289 (N_8289,N_4516,N_3051);
xnor U8290 (N_8290,N_3555,N_4500);
and U8291 (N_8291,N_3285,N_115);
xor U8292 (N_8292,N_786,N_4526);
nand U8293 (N_8293,N_1243,N_2663);
and U8294 (N_8294,N_5272,N_1502);
or U8295 (N_8295,N_3708,N_5996);
xnor U8296 (N_8296,N_4735,N_3251);
and U8297 (N_8297,N_4401,N_4219);
and U8298 (N_8298,N_1587,N_4241);
nor U8299 (N_8299,N_1284,N_2737);
and U8300 (N_8300,N_5399,N_21);
or U8301 (N_8301,N_5369,N_3387);
xnor U8302 (N_8302,N_5676,N_936);
xnor U8303 (N_8303,N_3091,N_4372);
xnor U8304 (N_8304,N_5533,N_4180);
xnor U8305 (N_8305,N_339,N_2889);
nor U8306 (N_8306,N_4468,N_5633);
nor U8307 (N_8307,N_4809,N_5123);
nand U8308 (N_8308,N_3539,N_2291);
or U8309 (N_8309,N_4803,N_2034);
nand U8310 (N_8310,N_2989,N_956);
and U8311 (N_8311,N_4301,N_1064);
nand U8312 (N_8312,N_5557,N_1750);
nand U8313 (N_8313,N_494,N_5046);
nand U8314 (N_8314,N_2418,N_3797);
nand U8315 (N_8315,N_3971,N_4181);
xor U8316 (N_8316,N_2135,N_1171);
nor U8317 (N_8317,N_3689,N_3768);
nand U8318 (N_8318,N_1024,N_4250);
nor U8319 (N_8319,N_4901,N_679);
or U8320 (N_8320,N_2580,N_1366);
xnor U8321 (N_8321,N_4422,N_3480);
xnor U8322 (N_8322,N_2832,N_1299);
xnor U8323 (N_8323,N_315,N_3522);
nand U8324 (N_8324,N_1678,N_952);
or U8325 (N_8325,N_3009,N_5083);
xor U8326 (N_8326,N_865,N_1389);
nand U8327 (N_8327,N_5768,N_3547);
nor U8328 (N_8328,N_5437,N_5070);
nor U8329 (N_8329,N_2867,N_470);
xor U8330 (N_8330,N_968,N_5750);
or U8331 (N_8331,N_1344,N_3996);
xnor U8332 (N_8332,N_2834,N_5585);
nand U8333 (N_8333,N_4299,N_4838);
and U8334 (N_8334,N_3406,N_1115);
xor U8335 (N_8335,N_5443,N_4412);
nor U8336 (N_8336,N_1193,N_1861);
xor U8337 (N_8337,N_4440,N_2804);
xor U8338 (N_8338,N_3207,N_1814);
nor U8339 (N_8339,N_3057,N_2975);
and U8340 (N_8340,N_4699,N_2462);
and U8341 (N_8341,N_4512,N_1240);
nand U8342 (N_8342,N_2564,N_4185);
and U8343 (N_8343,N_1386,N_281);
nor U8344 (N_8344,N_1106,N_774);
and U8345 (N_8345,N_4684,N_858);
nand U8346 (N_8346,N_4733,N_3628);
xnor U8347 (N_8347,N_4649,N_2837);
xnor U8348 (N_8348,N_1099,N_2043);
nor U8349 (N_8349,N_5268,N_2315);
or U8350 (N_8350,N_1495,N_2158);
nor U8351 (N_8351,N_1559,N_5210);
and U8352 (N_8352,N_4143,N_2668);
nand U8353 (N_8353,N_5471,N_3998);
nor U8354 (N_8354,N_1703,N_4665);
or U8355 (N_8355,N_831,N_4570);
nor U8356 (N_8356,N_819,N_5761);
nor U8357 (N_8357,N_5902,N_3737);
or U8358 (N_8358,N_4380,N_4154);
and U8359 (N_8359,N_3623,N_1482);
and U8360 (N_8360,N_3735,N_2269);
nand U8361 (N_8361,N_4421,N_2678);
xnor U8362 (N_8362,N_5763,N_5999);
and U8363 (N_8363,N_3344,N_622);
xnor U8364 (N_8364,N_2718,N_3810);
xnor U8365 (N_8365,N_3225,N_5032);
nand U8366 (N_8366,N_2644,N_5665);
nand U8367 (N_8367,N_2656,N_3770);
nor U8368 (N_8368,N_2803,N_2787);
xor U8369 (N_8369,N_791,N_63);
nor U8370 (N_8370,N_1150,N_504);
or U8371 (N_8371,N_2276,N_5783);
xor U8372 (N_8372,N_3788,N_738);
and U8373 (N_8373,N_3518,N_3420);
and U8374 (N_8374,N_4837,N_3450);
or U8375 (N_8375,N_1972,N_5500);
xor U8376 (N_8376,N_2443,N_2053);
xnor U8377 (N_8377,N_5469,N_148);
or U8378 (N_8378,N_3039,N_633);
nand U8379 (N_8379,N_3313,N_5802);
nand U8380 (N_8380,N_1936,N_4725);
and U8381 (N_8381,N_4954,N_3449);
nor U8382 (N_8382,N_3873,N_3306);
xnor U8383 (N_8383,N_4807,N_2976);
or U8384 (N_8384,N_4839,N_197);
or U8385 (N_8385,N_1443,N_3150);
nor U8386 (N_8386,N_18,N_4601);
or U8387 (N_8387,N_1688,N_3300);
nand U8388 (N_8388,N_2184,N_2197);
or U8389 (N_8389,N_4831,N_5328);
and U8390 (N_8390,N_3505,N_2684);
xor U8391 (N_8391,N_5952,N_2193);
and U8392 (N_8392,N_4675,N_5631);
nor U8393 (N_8393,N_988,N_3540);
or U8394 (N_8394,N_2936,N_1309);
or U8395 (N_8395,N_1394,N_2944);
nor U8396 (N_8396,N_1301,N_4987);
xnor U8397 (N_8397,N_2821,N_839);
or U8398 (N_8398,N_1993,N_718);
nor U8399 (N_8399,N_3909,N_35);
nand U8400 (N_8400,N_777,N_1930);
or U8401 (N_8401,N_3961,N_2655);
nor U8402 (N_8402,N_626,N_284);
or U8403 (N_8403,N_1833,N_2416);
xnor U8404 (N_8404,N_894,N_4824);
and U8405 (N_8405,N_4546,N_4393);
and U8406 (N_8406,N_3417,N_1196);
nor U8407 (N_8407,N_2494,N_3095);
xor U8408 (N_8408,N_4092,N_3911);
nor U8409 (N_8409,N_4163,N_3249);
nand U8410 (N_8410,N_3587,N_2010);
and U8411 (N_8411,N_282,N_2894);
or U8412 (N_8412,N_4503,N_4908);
nand U8413 (N_8413,N_157,N_4600);
nor U8414 (N_8414,N_126,N_5874);
and U8415 (N_8415,N_4218,N_525);
or U8416 (N_8416,N_3620,N_3441);
nor U8417 (N_8417,N_5595,N_4055);
or U8418 (N_8418,N_5744,N_2073);
xor U8419 (N_8419,N_2149,N_3945);
or U8420 (N_8420,N_2109,N_5863);
or U8421 (N_8421,N_5606,N_2955);
and U8422 (N_8422,N_88,N_5950);
and U8423 (N_8423,N_1378,N_3842);
xor U8424 (N_8424,N_2330,N_222);
and U8425 (N_8425,N_3317,N_1650);
nand U8426 (N_8426,N_5363,N_285);
nor U8427 (N_8427,N_915,N_2022);
xor U8428 (N_8428,N_3811,N_715);
nor U8429 (N_8429,N_2863,N_4171);
or U8430 (N_8430,N_5857,N_5971);
nor U8431 (N_8431,N_1922,N_462);
nand U8432 (N_8432,N_1704,N_4090);
nand U8433 (N_8433,N_2986,N_1932);
nand U8434 (N_8434,N_1528,N_5504);
and U8435 (N_8435,N_885,N_1672);
nor U8436 (N_8436,N_1020,N_2203);
nand U8437 (N_8437,N_1994,N_3527);
xnor U8438 (N_8438,N_2907,N_3507);
nand U8439 (N_8439,N_1484,N_2045);
nor U8440 (N_8440,N_1886,N_3315);
or U8441 (N_8441,N_1675,N_2917);
or U8442 (N_8442,N_5240,N_297);
or U8443 (N_8443,N_2483,N_402);
or U8444 (N_8444,N_5734,N_3160);
nand U8445 (N_8445,N_3404,N_5670);
xnor U8446 (N_8446,N_5501,N_4961);
and U8447 (N_8447,N_512,N_3458);
and U8448 (N_8448,N_4487,N_1187);
and U8449 (N_8449,N_3396,N_795);
nor U8450 (N_8450,N_781,N_5652);
and U8451 (N_8451,N_749,N_5460);
and U8452 (N_8452,N_3580,N_5266);
nor U8453 (N_8453,N_1391,N_221);
nor U8454 (N_8454,N_731,N_5503);
and U8455 (N_8455,N_869,N_2393);
xnor U8456 (N_8456,N_3117,N_1313);
and U8457 (N_8457,N_5385,N_1364);
and U8458 (N_8458,N_5721,N_2003);
nand U8459 (N_8459,N_1920,N_4186);
and U8460 (N_8460,N_4242,N_4647);
nor U8461 (N_8461,N_287,N_4801);
and U8462 (N_8462,N_892,N_1412);
or U8463 (N_8463,N_3684,N_4291);
nor U8464 (N_8464,N_5248,N_1450);
nand U8465 (N_8465,N_1837,N_2815);
and U8466 (N_8466,N_1445,N_1537);
nand U8467 (N_8467,N_5461,N_2847);
xnor U8468 (N_8468,N_2042,N_2728);
and U8469 (N_8469,N_1073,N_653);
and U8470 (N_8470,N_2708,N_1964);
xor U8471 (N_8471,N_4673,N_628);
nand U8472 (N_8472,N_490,N_3949);
nor U8473 (N_8473,N_943,N_5438);
xnor U8474 (N_8474,N_3227,N_2636);
and U8475 (N_8475,N_4637,N_2378);
nor U8476 (N_8476,N_2377,N_2240);
and U8477 (N_8477,N_4279,N_1531);
nor U8478 (N_8478,N_326,N_4543);
and U8479 (N_8479,N_545,N_2736);
nand U8480 (N_8480,N_5346,N_277);
or U8481 (N_8481,N_1278,N_0);
and U8482 (N_8482,N_5540,N_5871);
and U8483 (N_8483,N_1929,N_543);
or U8484 (N_8484,N_1358,N_740);
and U8485 (N_8485,N_2969,N_2583);
or U8486 (N_8486,N_4187,N_4353);
xor U8487 (N_8487,N_5840,N_1616);
nor U8488 (N_8488,N_3511,N_3670);
nand U8489 (N_8489,N_1111,N_5485);
xnor U8490 (N_8490,N_3499,N_905);
nand U8491 (N_8491,N_3576,N_1242);
xor U8492 (N_8492,N_2090,N_2635);
xor U8493 (N_8493,N_5122,N_3509);
and U8494 (N_8494,N_4856,N_1211);
and U8495 (N_8495,N_698,N_2427);
xnor U8496 (N_8496,N_972,N_659);
and U8497 (N_8497,N_4965,N_4614);
and U8498 (N_8498,N_5276,N_1137);
nor U8499 (N_8499,N_3395,N_1599);
nor U8500 (N_8500,N_2396,N_5578);
nand U8501 (N_8501,N_5977,N_1046);
and U8502 (N_8502,N_4984,N_2125);
xor U8503 (N_8503,N_4161,N_4452);
or U8504 (N_8504,N_3215,N_2247);
and U8505 (N_8505,N_854,N_921);
xor U8506 (N_8506,N_1088,N_261);
xnor U8507 (N_8507,N_2971,N_4975);
nor U8508 (N_8508,N_350,N_4403);
and U8509 (N_8509,N_4247,N_1118);
and U8510 (N_8510,N_4960,N_1739);
nand U8511 (N_8511,N_1414,N_5311);
nor U8512 (N_8512,N_3001,N_5908);
xor U8513 (N_8513,N_4511,N_610);
xor U8514 (N_8514,N_1551,N_2560);
or U8515 (N_8515,N_594,N_4415);
nand U8516 (N_8516,N_737,N_815);
and U8517 (N_8517,N_852,N_1796);
xor U8518 (N_8518,N_4238,N_939);
xor U8519 (N_8519,N_1545,N_3877);
xnor U8520 (N_8520,N_1902,N_1203);
nand U8521 (N_8521,N_4866,N_4694);
xnor U8522 (N_8522,N_5494,N_4967);
nand U8523 (N_8523,N_2537,N_3897);
nor U8524 (N_8524,N_5291,N_1489);
or U8525 (N_8525,N_1540,N_3118);
nor U8526 (N_8526,N_4643,N_5155);
nand U8527 (N_8527,N_5545,N_2828);
xnor U8528 (N_8528,N_2,N_1474);
and U8529 (N_8529,N_997,N_3875);
nor U8530 (N_8530,N_3609,N_5525);
nand U8531 (N_8531,N_5044,N_4069);
nand U8532 (N_8532,N_3700,N_4577);
and U8533 (N_8533,N_3086,N_4766);
xnor U8534 (N_8534,N_3105,N_1646);
nor U8535 (N_8535,N_3358,N_4588);
nand U8536 (N_8536,N_4781,N_5803);
nor U8537 (N_8537,N_5716,N_5765);
xnor U8538 (N_8538,N_4413,N_2237);
nand U8539 (N_8539,N_1564,N_3612);
xnor U8540 (N_8540,N_5924,N_4691);
nand U8541 (N_8541,N_3637,N_4905);
and U8542 (N_8542,N_45,N_660);
nor U8543 (N_8543,N_5711,N_4595);
nand U8544 (N_8544,N_4657,N_646);
and U8545 (N_8545,N_457,N_3690);
nand U8546 (N_8546,N_4677,N_5737);
nand U8547 (N_8547,N_5202,N_1049);
nand U8548 (N_8548,N_2481,N_1052);
nor U8549 (N_8549,N_2405,N_5536);
or U8550 (N_8550,N_2324,N_4131);
xor U8551 (N_8551,N_5523,N_1424);
or U8552 (N_8552,N_681,N_3481);
xor U8553 (N_8553,N_5746,N_445);
or U8554 (N_8554,N_1843,N_236);
nand U8555 (N_8555,N_4902,N_5520);
or U8556 (N_8556,N_2205,N_4872);
xor U8557 (N_8557,N_2525,N_1656);
xor U8558 (N_8558,N_3321,N_1398);
xor U8559 (N_8559,N_579,N_2417);
and U8560 (N_8560,N_2842,N_5017);
or U8561 (N_8561,N_3131,N_3085);
nor U8562 (N_8562,N_899,N_3517);
xnor U8563 (N_8563,N_2949,N_1377);
and U8564 (N_8564,N_2893,N_1239);
nand U8565 (N_8565,N_1010,N_4885);
nand U8566 (N_8566,N_207,N_3924);
nor U8567 (N_8567,N_2422,N_3019);
nand U8568 (N_8568,N_2074,N_908);
and U8569 (N_8569,N_5470,N_2972);
and U8570 (N_8570,N_4494,N_5096);
and U8571 (N_8571,N_3407,N_5647);
or U8572 (N_8572,N_2781,N_3183);
or U8573 (N_8573,N_2478,N_5479);
nand U8574 (N_8574,N_1168,N_4492);
and U8575 (N_8575,N_1059,N_2049);
or U8576 (N_8576,N_1781,N_3199);
and U8577 (N_8577,N_5279,N_4958);
xor U8578 (N_8578,N_3158,N_630);
and U8579 (N_8579,N_1976,N_2244);
xnor U8580 (N_8580,N_5440,N_5991);
nor U8581 (N_8581,N_1784,N_3535);
nand U8582 (N_8582,N_101,N_3254);
and U8583 (N_8583,N_168,N_465);
xnor U8584 (N_8584,N_5094,N_4429);
xnor U8585 (N_8585,N_4799,N_4879);
nor U8586 (N_8586,N_134,N_4191);
nand U8587 (N_8587,N_814,N_3703);
xor U8588 (N_8588,N_1492,N_416);
and U8589 (N_8589,N_1577,N_1156);
xnor U8590 (N_8590,N_5653,N_3173);
nor U8591 (N_8591,N_4775,N_883);
and U8592 (N_8592,N_4737,N_2278);
nor U8593 (N_8593,N_1874,N_747);
nor U8594 (N_8594,N_3459,N_4347);
nor U8595 (N_8595,N_4679,N_2339);
nor U8596 (N_8596,N_2226,N_2023);
xor U8597 (N_8597,N_2961,N_1916);
and U8598 (N_8598,N_2432,N_4927);
or U8599 (N_8599,N_3510,N_2912);
nor U8600 (N_8600,N_5451,N_2671);
and U8601 (N_8601,N_1343,N_979);
and U8602 (N_8602,N_3472,N_4262);
or U8603 (N_8603,N_4325,N_567);
and U8604 (N_8604,N_1303,N_4738);
and U8605 (N_8605,N_553,N_53);
and U8606 (N_8606,N_1113,N_299);
and U8607 (N_8607,N_2813,N_2384);
xnor U8608 (N_8608,N_3782,N_2316);
xnor U8609 (N_8609,N_1787,N_1339);
and U8610 (N_8610,N_5824,N_5480);
or U8611 (N_8611,N_2634,N_4938);
xor U8612 (N_8612,N_1285,N_1967);
xor U8613 (N_8613,N_3858,N_1027);
nand U8614 (N_8614,N_3933,N_4349);
xnor U8615 (N_8615,N_1096,N_5576);
or U8616 (N_8616,N_5566,N_398);
or U8617 (N_8617,N_807,N_3161);
nor U8618 (N_8618,N_4499,N_4978);
nand U8619 (N_8619,N_4033,N_448);
nand U8620 (N_8620,N_4431,N_3645);
xor U8621 (N_8621,N_2616,N_4950);
nor U8622 (N_8622,N_2228,N_570);
or U8623 (N_8623,N_5511,N_1608);
and U8624 (N_8624,N_202,N_4148);
nand U8625 (N_8625,N_3320,N_5102);
nand U8626 (N_8626,N_3880,N_2366);
xnor U8627 (N_8627,N_272,N_5082);
or U8628 (N_8628,N_4948,N_233);
xnor U8629 (N_8629,N_1827,N_1592);
nor U8630 (N_8630,N_2019,N_346);
and U8631 (N_8631,N_1556,N_3259);
or U8632 (N_8632,N_933,N_4825);
or U8633 (N_8633,N_3453,N_3973);
nor U8634 (N_8634,N_3079,N_5309);
nand U8635 (N_8635,N_4989,N_142);
nand U8636 (N_8636,N_5257,N_5259);
nand U8637 (N_8637,N_2165,N_1425);
or U8638 (N_8638,N_2089,N_3981);
and U8639 (N_8639,N_1300,N_2891);
xor U8640 (N_8640,N_1045,N_2719);
and U8641 (N_8641,N_1418,N_5428);
nor U8642 (N_8642,N_2037,N_143);
or U8643 (N_8643,N_3720,N_4123);
and U8644 (N_8644,N_10,N_673);
nor U8645 (N_8645,N_1799,N_259);
or U8646 (N_8646,N_3332,N_2795);
or U8647 (N_8647,N_4674,N_2860);
xor U8648 (N_8648,N_794,N_1749);
nor U8649 (N_8649,N_2487,N_3716);
nor U8650 (N_8650,N_4153,N_1082);
or U8651 (N_8651,N_1077,N_3760);
xor U8652 (N_8652,N_65,N_3208);
nand U8653 (N_8653,N_2007,N_796);
or U8654 (N_8654,N_2559,N_5145);
or U8655 (N_8655,N_2549,N_1891);
nor U8656 (N_8656,N_4579,N_4402);
nor U8657 (N_8657,N_4739,N_4626);
nor U8658 (N_8658,N_196,N_1051);
or U8659 (N_8659,N_3246,N_1776);
nor U8660 (N_8660,N_5732,N_4602);
nor U8661 (N_8661,N_5778,N_5139);
or U8662 (N_8662,N_1330,N_2380);
xnor U8663 (N_8663,N_3366,N_829);
nand U8664 (N_8664,N_5724,N_2769);
nor U8665 (N_8665,N_5299,N_3104);
xor U8666 (N_8666,N_87,N_1375);
nor U8667 (N_8667,N_1076,N_482);
or U8668 (N_8668,N_4592,N_1224);
and U8669 (N_8669,N_4449,N_3336);
nor U8670 (N_8670,N_1801,N_4095);
and U8671 (N_8671,N_5941,N_4970);
xnor U8672 (N_8672,N_970,N_1903);
nand U8673 (N_8673,N_1975,N_4346);
nand U8674 (N_8674,N_4195,N_3044);
nor U8675 (N_8675,N_3872,N_1420);
and U8676 (N_8676,N_3483,N_1626);
nor U8677 (N_8677,N_2869,N_1351);
nand U8678 (N_8678,N_2167,N_3905);
xor U8679 (N_8679,N_2848,N_520);
nor U8680 (N_8680,N_4167,N_876);
nor U8681 (N_8681,N_5090,N_3323);
nor U8682 (N_8682,N_2479,N_3928);
and U8683 (N_8683,N_4722,N_1017);
and U8684 (N_8684,N_198,N_2369);
nand U8685 (N_8685,N_1464,N_116);
nor U8686 (N_8686,N_4656,N_3231);
or U8687 (N_8687,N_2555,N_2628);
or U8688 (N_8688,N_1235,N_4916);
and U8689 (N_8689,N_1191,N_5825);
xor U8690 (N_8690,N_5329,N_861);
or U8691 (N_8691,N_1560,N_4963);
and U8692 (N_8692,N_1452,N_600);
nor U8693 (N_8693,N_5995,N_617);
xor U8694 (N_8694,N_3184,N_4746);
or U8695 (N_8695,N_477,N_2190);
and U8696 (N_8696,N_3753,N_4096);
nand U8697 (N_8697,N_4035,N_5693);
and U8698 (N_8698,N_2554,N_5617);
nor U8699 (N_8699,N_2419,N_5009);
xnor U8700 (N_8700,N_5059,N_1185);
nor U8701 (N_8701,N_1121,N_1575);
nand U8702 (N_8702,N_503,N_2685);
nor U8703 (N_8703,N_4157,N_576);
nor U8704 (N_8704,N_1214,N_1510);
or U8705 (N_8705,N_4140,N_1676);
and U8706 (N_8706,N_5103,N_3813);
nand U8707 (N_8707,N_5982,N_895);
or U8708 (N_8708,N_566,N_4991);
xor U8709 (N_8709,N_1516,N_4478);
nand U8710 (N_8710,N_4873,N_1178);
and U8711 (N_8711,N_5180,N_3613);
and U8712 (N_8712,N_1586,N_5058);
nand U8713 (N_8713,N_2997,N_1160);
nand U8714 (N_8714,N_4398,N_2154);
or U8715 (N_8715,N_1388,N_1019);
nand U8716 (N_8716,N_3340,N_3319);
or U8717 (N_8717,N_1943,N_241);
or U8718 (N_8718,N_5140,N_4103);
xor U8719 (N_8719,N_3411,N_4220);
xor U8720 (N_8720,N_2591,N_472);
or U8721 (N_8721,N_1604,N_456);
nand U8722 (N_8722,N_5986,N_4999);
nand U8723 (N_8723,N_5233,N_2888);
xnor U8724 (N_8724,N_4741,N_2002);
nor U8725 (N_8725,N_5779,N_716);
nand U8726 (N_8726,N_38,N_1365);
nand U8727 (N_8727,N_1254,N_4133);
or U8728 (N_8728,N_3899,N_3970);
and U8729 (N_8729,N_3993,N_4868);
or U8730 (N_8730,N_1012,N_4086);
or U8731 (N_8731,N_564,N_3901);
xor U8732 (N_8732,N_5984,N_5628);
nand U8733 (N_8733,N_4172,N_496);
nor U8734 (N_8734,N_587,N_616);
xnor U8735 (N_8735,N_3721,N_5358);
xnor U8736 (N_8736,N_2103,N_5791);
xor U8737 (N_8737,N_4072,N_3687);
nand U8738 (N_8738,N_2449,N_4669);
and U8739 (N_8739,N_789,N_4716);
or U8740 (N_8740,N_5338,N_3934);
or U8741 (N_8741,N_4688,N_4764);
nand U8742 (N_8742,N_4576,N_1454);
nand U8743 (N_8743,N_951,N_2578);
xor U8744 (N_8744,N_1040,N_3923);
nand U8745 (N_8745,N_5243,N_5618);
xor U8746 (N_8746,N_635,N_5751);
and U8747 (N_8747,N_3245,N_2209);
and U8748 (N_8748,N_4356,N_4553);
xnor U8749 (N_8749,N_4581,N_3958);
xnor U8750 (N_8750,N_4286,N_5482);
and U8751 (N_8751,N_4826,N_3328);
xor U8752 (N_8752,N_3551,N_2594);
nor U8753 (N_8753,N_608,N_3166);
nand U8754 (N_8754,N_4405,N_218);
nor U8755 (N_8755,N_4616,N_2852);
xor U8756 (N_8756,N_4608,N_1360);
or U8757 (N_8757,N_199,N_2861);
xor U8758 (N_8758,N_3741,N_5510);
or U8759 (N_8759,N_4388,N_369);
xor U8760 (N_8760,N_1868,N_1250);
nand U8761 (N_8761,N_1996,N_5326);
nor U8762 (N_8762,N_3847,N_2754);
xnor U8763 (N_8763,N_3288,N_19);
or U8764 (N_8764,N_4723,N_4604);
and U8765 (N_8765,N_3058,N_2093);
and U8766 (N_8766,N_1390,N_489);
xor U8767 (N_8767,N_1794,N_4160);
nor U8768 (N_8768,N_4436,N_817);
nand U8769 (N_8769,N_3523,N_4922);
xor U8770 (N_8770,N_3821,N_1459);
or U8771 (N_8771,N_1249,N_4112);
nor U8772 (N_8772,N_4276,N_5452);
nand U8773 (N_8773,N_3792,N_4414);
xor U8774 (N_8774,N_5221,N_2675);
or U8775 (N_8775,N_4770,N_5677);
nand U8776 (N_8776,N_4521,N_2114);
or U8777 (N_8777,N_875,N_242);
or U8778 (N_8778,N_1514,N_5345);
and U8779 (N_8779,N_4223,N_1439);
xnor U8780 (N_8780,N_4993,N_2941);
or U8781 (N_8781,N_4923,N_4720);
nand U8782 (N_8782,N_1006,N_2281);
nand U8783 (N_8783,N_1951,N_5524);
nor U8784 (N_8784,N_430,N_2515);
xor U8785 (N_8785,N_3178,N_3077);
or U8786 (N_8786,N_2964,N_4284);
or U8787 (N_8787,N_1141,N_2130);
nor U8788 (N_8788,N_2424,N_3766);
nor U8789 (N_8789,N_5586,N_1869);
and U8790 (N_8790,N_2509,N_5881);
or U8791 (N_8791,N_4355,N_1686);
and U8792 (N_8792,N_4442,N_2505);
or U8793 (N_8793,N_4082,N_5270);
nand U8794 (N_8794,N_4767,N_3860);
xnor U8795 (N_8795,N_4888,N_4944);
nor U8796 (N_8796,N_395,N_4322);
nor U8797 (N_8797,N_571,N_506);
xor U8798 (N_8798,N_806,N_3633);
nand U8799 (N_8799,N_5189,N_4438);
or U8800 (N_8800,N_2078,N_3354);
xor U8801 (N_8801,N_1593,N_5660);
nand U8802 (N_8802,N_2222,N_1279);
xor U8803 (N_8803,N_117,N_3172);
nand U8804 (N_8804,N_4070,N_483);
nor U8805 (N_8805,N_2900,N_1335);
nor U8806 (N_8806,N_5981,N_4408);
or U8807 (N_8807,N_2806,N_1139);
nor U8808 (N_8808,N_4237,N_4194);
nand U8809 (N_8809,N_5280,N_5597);
nand U8810 (N_8810,N_5013,N_518);
nor U8811 (N_8811,N_4382,N_4536);
and U8812 (N_8812,N_3619,N_898);
and U8813 (N_8813,N_3764,N_5580);
xnor U8814 (N_8814,N_92,N_2077);
or U8815 (N_8815,N_2939,N_4309);
and U8816 (N_8816,N_3232,N_2592);
or U8817 (N_8817,N_2279,N_169);
xor U8818 (N_8818,N_52,N_1621);
and U8819 (N_8819,N_2402,N_5910);
xnor U8820 (N_8820,N_2826,N_1236);
nor U8821 (N_8821,N_5316,N_3976);
nor U8822 (N_8822,N_4880,N_2790);
nand U8823 (N_8823,N_2192,N_1385);
nor U8824 (N_8824,N_3986,N_1562);
xnor U8825 (N_8825,N_3662,N_1458);
xnor U8826 (N_8826,N_2008,N_2933);
or U8827 (N_8827,N_3542,N_5696);
or U8828 (N_8828,N_1820,N_3144);
nor U8829 (N_8829,N_2916,N_3730);
xnor U8830 (N_8830,N_2409,N_3487);
or U8831 (N_8831,N_3269,N_1047);
xnor U8832 (N_8832,N_2962,N_2855);
or U8833 (N_8833,N_3278,N_4687);
nand U8834 (N_8834,N_1346,N_5472);
nor U8835 (N_8835,N_1501,N_4997);
xor U8836 (N_8836,N_1016,N_68);
xnor U8837 (N_8837,N_114,N_2302);
and U8838 (N_8838,N_4458,N_2713);
xnor U8839 (N_8839,N_3067,N_4270);
xnor U8840 (N_8840,N_5929,N_4612);
and U8841 (N_8841,N_4045,N_411);
and U8842 (N_8842,N_5541,N_2987);
xnor U8843 (N_8843,N_5228,N_4471);
and U8844 (N_8844,N_3964,N_235);
xnor U8845 (N_8845,N_3021,N_4407);
or U8846 (N_8846,N_1044,N_4708);
nand U8847 (N_8847,N_2098,N_5130);
nor U8848 (N_8848,N_3080,N_389);
xnor U8849 (N_8849,N_1371,N_902);
nor U8850 (N_8850,N_4653,N_5507);
and U8851 (N_8851,N_2447,N_3274);
nand U8852 (N_8852,N_2391,N_2566);
nand U8853 (N_8853,N_4556,N_3562);
or U8854 (N_8854,N_1237,N_4437);
xor U8855 (N_8855,N_714,N_5594);
or U8856 (N_8856,N_2458,N_2722);
or U8857 (N_8857,N_3135,N_2491);
xor U8858 (N_8858,N_4890,N_4539);
or U8859 (N_8859,N_6,N_3969);
nand U8860 (N_8860,N_1572,N_59);
or U8861 (N_8861,N_4423,N_5650);
nor U8862 (N_8862,N_713,N_5644);
xor U8863 (N_8863,N_1340,N_5450);
or U8864 (N_8864,N_1655,N_1219);
nand U8865 (N_8865,N_1317,N_5643);
xor U8866 (N_8866,N_20,N_5899);
and U8867 (N_8867,N_3034,N_5341);
or U8868 (N_8868,N_3789,N_3963);
nand U8869 (N_8869,N_1430,N_2624);
nor U8870 (N_8870,N_3143,N_3892);
nor U8871 (N_8871,N_1590,N_407);
or U8872 (N_8872,N_4255,N_79);
nand U8873 (N_8873,N_2459,N_5828);
or U8874 (N_8874,N_4101,N_3652);
xor U8875 (N_8875,N_180,N_2864);
nor U8876 (N_8876,N_1136,N_4549);
or U8877 (N_8877,N_5353,N_4533);
nor U8878 (N_8878,N_1822,N_420);
or U8879 (N_8879,N_1734,N_5409);
nor U8880 (N_8880,N_1402,N_2000);
nand U8881 (N_8881,N_3756,N_5137);
xnor U8882 (N_8882,N_753,N_4590);
and U8883 (N_8883,N_387,N_4137);
nand U8884 (N_8884,N_4933,N_2072);
xnor U8885 (N_8885,N_2548,N_4136);
and U8886 (N_8886,N_4910,N_595);
or U8887 (N_8887,N_3536,N_508);
nor U8888 (N_8888,N_766,N_1504);
and U8889 (N_8889,N_5957,N_5455);
nor U8890 (N_8890,N_3289,N_4522);
or U8891 (N_8891,N_293,N_5466);
or U8892 (N_8892,N_461,N_5442);
nand U8893 (N_8893,N_240,N_2504);
nand U8894 (N_8894,N_5288,N_5349);
nor U8895 (N_8895,N_541,N_368);
nor U8896 (N_8896,N_2503,N_5220);
or U8897 (N_8897,N_1863,N_5695);
xnor U8898 (N_8898,N_3329,N_4678);
nand U8899 (N_8899,N_572,N_497);
nor U8900 (N_8900,N_4283,N_1758);
nor U8901 (N_8901,N_1705,N_3910);
xnor U8902 (N_8902,N_1687,N_954);
xnor U8903 (N_8903,N_3955,N_2729);
nor U8904 (N_8904,N_1042,N_707);
nor U8905 (N_8905,N_2139,N_4535);
or U8906 (N_8906,N_3383,N_5132);
nor U8907 (N_8907,N_2155,N_721);
xnor U8908 (N_8908,N_1307,N_2814);
and U8909 (N_8909,N_4445,N_5244);
nor U8910 (N_8910,N_661,N_577);
nand U8911 (N_8911,N_3640,N_4383);
nand U8912 (N_8912,N_4253,N_1325);
or U8913 (N_8913,N_4020,N_4078);
and U8914 (N_8914,N_3500,N_3412);
and U8915 (N_8915,N_367,N_1726);
and U8916 (N_8916,N_2332,N_5933);
and U8917 (N_8917,N_1779,N_4586);
and U8918 (N_8918,N_5394,N_639);
nor U8919 (N_8919,N_2297,N_4465);
xor U8920 (N_8920,N_4043,N_3868);
or U8921 (N_8921,N_2734,N_2500);
xnor U8922 (N_8922,N_2926,N_2076);
nor U8923 (N_8923,N_5282,N_720);
xnor U8924 (N_8924,N_2883,N_4307);
nor U8925 (N_8925,N_1627,N_5529);
nand U8926 (N_8926,N_2404,N_967);
xnor U8927 (N_8927,N_4875,N_5729);
and U8928 (N_8928,N_782,N_192);
nand U8929 (N_8929,N_5227,N_4509);
nor U8930 (N_8930,N_5296,N_3088);
or U8931 (N_8931,N_1885,N_183);
or U8932 (N_8932,N_3308,N_5970);
nand U8933 (N_8933,N_1606,N_1907);
and U8934 (N_8934,N_2615,N_1270);
nor U8935 (N_8935,N_1992,N_2097);
nand U8936 (N_8936,N_2334,N_2873);
nor U8937 (N_8937,N_5845,N_699);
or U8938 (N_8938,N_2157,N_1022);
xor U8939 (N_8939,N_4913,N_2001);
and U8940 (N_8940,N_5118,N_5381);
nor U8941 (N_8941,N_4350,N_3036);
nor U8942 (N_8942,N_1619,N_29);
or U8943 (N_8943,N_5722,N_4071);
xor U8944 (N_8944,N_5006,N_1725);
or U8945 (N_8945,N_4466,N_4376);
or U8946 (N_8946,N_4854,N_378);
nor U8947 (N_8947,N_3552,N_5432);
xnor U8948 (N_8948,N_3682,N_3806);
nor U8949 (N_8949,N_1828,N_4790);
nor U8950 (N_8950,N_1074,N_3391);
or U8951 (N_8951,N_5295,N_863);
nor U8952 (N_8952,N_4052,N_4263);
and U8953 (N_8953,N_3502,N_5030);
or U8954 (N_8954,N_1691,N_1422);
or U8955 (N_8955,N_2381,N_5441);
nor U8956 (N_8956,N_2455,N_1089);
nand U8957 (N_8957,N_729,N_2885);
or U8958 (N_8958,N_1192,N_5486);
nand U8959 (N_8959,N_425,N_3241);
and U8960 (N_8960,N_1525,N_2445);
or U8961 (N_8961,N_2513,N_3338);
xnor U8962 (N_8962,N_900,N_1706);
and U8963 (N_8963,N_5717,N_408);
nand U8964 (N_8964,N_756,N_1913);
xnor U8965 (N_8965,N_3097,N_5165);
nand U8966 (N_8966,N_2930,N_1607);
or U8967 (N_8967,N_4693,N_1241);
or U8968 (N_8968,N_4969,N_4515);
or U8969 (N_8969,N_4534,N_5179);
or U8970 (N_8970,N_5386,N_1355);
nand U8971 (N_8971,N_1416,N_5273);
nand U8972 (N_8972,N_4776,N_4387);
or U8973 (N_8973,N_3276,N_2887);
nand U8974 (N_8974,N_691,N_760);
nand U8975 (N_8975,N_2129,N_983);
nand U8976 (N_8976,N_2105,N_4711);
nor U8977 (N_8977,N_5215,N_4192);
xnor U8978 (N_8978,N_3729,N_4352);
nand U8979 (N_8979,N_2637,N_2680);
and U8980 (N_8980,N_1774,N_1673);
nor U8981 (N_8981,N_3857,N_404);
or U8982 (N_8982,N_423,N_4234);
nor U8983 (N_8983,N_5603,N_5657);
nand U8984 (N_8984,N_2664,N_5308);
xnor U8985 (N_8985,N_5334,N_3189);
nor U8986 (N_8986,N_5916,N_254);
xor U8987 (N_8987,N_2934,N_4574);
and U8988 (N_8988,N_4758,N_3156);
xnor U8989 (N_8989,N_3219,N_2033);
nand U8990 (N_8990,N_2373,N_4696);
and U8991 (N_8991,N_4921,N_1926);
or U8992 (N_8992,N_311,N_4351);
or U8993 (N_8993,N_3574,N_14);
nor U8994 (N_8994,N_2904,N_2650);
or U8995 (N_8995,N_4537,N_3643);
nor U8996 (N_8996,N_3163,N_4189);
or U8997 (N_8997,N_3198,N_1695);
or U8998 (N_8998,N_4834,N_2323);
nand U8999 (N_8999,N_3504,N_4313);
or U9000 (N_9000,N_2429,N_483);
nor U9001 (N_9001,N_3383,N_5553);
nand U9002 (N_9002,N_4973,N_4624);
xnor U9003 (N_9003,N_4670,N_2198);
xor U9004 (N_9004,N_4426,N_5355);
nand U9005 (N_9005,N_3327,N_4448);
and U9006 (N_9006,N_4113,N_2271);
and U9007 (N_9007,N_5879,N_2759);
and U9008 (N_9008,N_5521,N_2378);
xor U9009 (N_9009,N_968,N_2587);
xnor U9010 (N_9010,N_210,N_2668);
or U9011 (N_9011,N_1728,N_3306);
nor U9012 (N_9012,N_4757,N_5395);
nand U9013 (N_9013,N_3970,N_4966);
or U9014 (N_9014,N_28,N_1130);
or U9015 (N_9015,N_1142,N_5185);
or U9016 (N_9016,N_1176,N_1145);
and U9017 (N_9017,N_1908,N_1926);
nand U9018 (N_9018,N_1986,N_1120);
and U9019 (N_9019,N_688,N_2056);
and U9020 (N_9020,N_523,N_5976);
and U9021 (N_9021,N_1831,N_5025);
xnor U9022 (N_9022,N_1010,N_794);
nand U9023 (N_9023,N_39,N_362);
and U9024 (N_9024,N_5498,N_1983);
xor U9025 (N_9025,N_135,N_980);
and U9026 (N_9026,N_3585,N_5724);
nand U9027 (N_9027,N_5678,N_3482);
and U9028 (N_9028,N_3305,N_1820);
nand U9029 (N_9029,N_587,N_1903);
and U9030 (N_9030,N_2867,N_3157);
nand U9031 (N_9031,N_3035,N_4604);
xnor U9032 (N_9032,N_3825,N_385);
or U9033 (N_9033,N_5073,N_798);
or U9034 (N_9034,N_3867,N_187);
xor U9035 (N_9035,N_1112,N_5386);
nand U9036 (N_9036,N_217,N_3377);
xor U9037 (N_9037,N_2979,N_1050);
or U9038 (N_9038,N_4210,N_4752);
nand U9039 (N_9039,N_3323,N_4524);
or U9040 (N_9040,N_554,N_3130);
nand U9041 (N_9041,N_1746,N_2415);
nand U9042 (N_9042,N_4528,N_5735);
nor U9043 (N_9043,N_2647,N_2867);
nand U9044 (N_9044,N_3807,N_739);
and U9045 (N_9045,N_4298,N_2515);
or U9046 (N_9046,N_3710,N_3535);
nand U9047 (N_9047,N_5092,N_3897);
nand U9048 (N_9048,N_716,N_2147);
xor U9049 (N_9049,N_2063,N_3623);
or U9050 (N_9050,N_5241,N_4866);
and U9051 (N_9051,N_4142,N_2012);
and U9052 (N_9052,N_1031,N_2257);
nand U9053 (N_9053,N_2800,N_4082);
or U9054 (N_9054,N_3294,N_1045);
or U9055 (N_9055,N_1432,N_1761);
nor U9056 (N_9056,N_4594,N_398);
or U9057 (N_9057,N_3736,N_1265);
and U9058 (N_9058,N_5719,N_1339);
nor U9059 (N_9059,N_5613,N_2024);
and U9060 (N_9060,N_2548,N_2964);
or U9061 (N_9061,N_4274,N_5415);
nand U9062 (N_9062,N_1791,N_5042);
or U9063 (N_9063,N_4328,N_3836);
and U9064 (N_9064,N_889,N_5468);
xnor U9065 (N_9065,N_3260,N_4373);
nand U9066 (N_9066,N_4051,N_5486);
xnor U9067 (N_9067,N_987,N_2715);
or U9068 (N_9068,N_4058,N_4508);
nand U9069 (N_9069,N_697,N_746);
xnor U9070 (N_9070,N_1382,N_2418);
nand U9071 (N_9071,N_1461,N_2923);
nand U9072 (N_9072,N_4676,N_3419);
nand U9073 (N_9073,N_5103,N_457);
xnor U9074 (N_9074,N_5479,N_1765);
nand U9075 (N_9075,N_812,N_3627);
nor U9076 (N_9076,N_678,N_279);
nand U9077 (N_9077,N_5738,N_2646);
nand U9078 (N_9078,N_740,N_3492);
or U9079 (N_9079,N_4625,N_5751);
nor U9080 (N_9080,N_1042,N_3080);
nor U9081 (N_9081,N_4760,N_4378);
and U9082 (N_9082,N_2417,N_2482);
nor U9083 (N_9083,N_2472,N_1116);
xor U9084 (N_9084,N_838,N_2880);
xnor U9085 (N_9085,N_4370,N_872);
xnor U9086 (N_9086,N_5382,N_4032);
xor U9087 (N_9087,N_4155,N_5313);
nand U9088 (N_9088,N_4335,N_461);
nor U9089 (N_9089,N_166,N_4526);
xor U9090 (N_9090,N_2773,N_2650);
nand U9091 (N_9091,N_512,N_4617);
and U9092 (N_9092,N_2547,N_2657);
nand U9093 (N_9093,N_1667,N_3883);
nor U9094 (N_9094,N_5351,N_234);
xnor U9095 (N_9095,N_4290,N_5886);
xor U9096 (N_9096,N_5448,N_4378);
nor U9097 (N_9097,N_3897,N_5615);
or U9098 (N_9098,N_3877,N_5304);
and U9099 (N_9099,N_4394,N_1770);
nor U9100 (N_9100,N_3576,N_2733);
xnor U9101 (N_9101,N_2521,N_2613);
and U9102 (N_9102,N_3389,N_729);
nor U9103 (N_9103,N_1117,N_861);
nor U9104 (N_9104,N_595,N_4387);
or U9105 (N_9105,N_2653,N_3378);
and U9106 (N_9106,N_95,N_5652);
xnor U9107 (N_9107,N_3868,N_2728);
nand U9108 (N_9108,N_4368,N_4355);
and U9109 (N_9109,N_2534,N_907);
nand U9110 (N_9110,N_3471,N_2394);
xnor U9111 (N_9111,N_3487,N_1706);
nand U9112 (N_9112,N_5973,N_3684);
nor U9113 (N_9113,N_5802,N_3608);
or U9114 (N_9114,N_3484,N_5374);
xor U9115 (N_9115,N_4340,N_2387);
nor U9116 (N_9116,N_4352,N_3284);
nor U9117 (N_9117,N_3215,N_2757);
nor U9118 (N_9118,N_2249,N_5962);
xnor U9119 (N_9119,N_2046,N_1059);
xor U9120 (N_9120,N_4018,N_1467);
nand U9121 (N_9121,N_5260,N_2247);
xor U9122 (N_9122,N_5201,N_2344);
nand U9123 (N_9123,N_4945,N_3277);
nor U9124 (N_9124,N_707,N_3566);
xor U9125 (N_9125,N_1774,N_143);
nor U9126 (N_9126,N_2632,N_3037);
or U9127 (N_9127,N_5436,N_5438);
or U9128 (N_9128,N_4777,N_5155);
or U9129 (N_9129,N_3301,N_3032);
nand U9130 (N_9130,N_2956,N_3729);
nand U9131 (N_9131,N_1975,N_5231);
or U9132 (N_9132,N_228,N_3841);
and U9133 (N_9133,N_5379,N_1429);
nor U9134 (N_9134,N_5445,N_7);
xor U9135 (N_9135,N_5761,N_5510);
xor U9136 (N_9136,N_1012,N_4763);
xor U9137 (N_9137,N_3911,N_442);
or U9138 (N_9138,N_5271,N_1305);
nand U9139 (N_9139,N_3480,N_4079);
or U9140 (N_9140,N_5086,N_1051);
nand U9141 (N_9141,N_3492,N_139);
and U9142 (N_9142,N_4901,N_3825);
or U9143 (N_9143,N_3490,N_5605);
nor U9144 (N_9144,N_5883,N_4807);
nand U9145 (N_9145,N_4925,N_2713);
nor U9146 (N_9146,N_3644,N_5434);
xor U9147 (N_9147,N_3736,N_2630);
nor U9148 (N_9148,N_4332,N_2634);
nor U9149 (N_9149,N_319,N_2380);
and U9150 (N_9150,N_2974,N_1239);
xor U9151 (N_9151,N_602,N_1876);
nand U9152 (N_9152,N_4121,N_5094);
xnor U9153 (N_9153,N_4476,N_3215);
xnor U9154 (N_9154,N_3565,N_4493);
or U9155 (N_9155,N_3695,N_4508);
xor U9156 (N_9156,N_2931,N_496);
xnor U9157 (N_9157,N_2899,N_3833);
nand U9158 (N_9158,N_4941,N_4848);
nor U9159 (N_9159,N_5444,N_1620);
nor U9160 (N_9160,N_2004,N_3932);
xor U9161 (N_9161,N_5235,N_2744);
xor U9162 (N_9162,N_2456,N_670);
xor U9163 (N_9163,N_1919,N_294);
or U9164 (N_9164,N_1540,N_1049);
nand U9165 (N_9165,N_1846,N_5334);
nand U9166 (N_9166,N_5720,N_89);
and U9167 (N_9167,N_4342,N_1390);
and U9168 (N_9168,N_4274,N_1516);
xor U9169 (N_9169,N_4313,N_1513);
nand U9170 (N_9170,N_1036,N_980);
xor U9171 (N_9171,N_3630,N_4727);
nand U9172 (N_9172,N_23,N_3071);
nor U9173 (N_9173,N_1431,N_1905);
xor U9174 (N_9174,N_1719,N_5374);
and U9175 (N_9175,N_3750,N_2342);
xnor U9176 (N_9176,N_1840,N_5058);
xor U9177 (N_9177,N_1770,N_4805);
nand U9178 (N_9178,N_1865,N_2259);
or U9179 (N_9179,N_4344,N_781);
nor U9180 (N_9180,N_5613,N_2606);
xnor U9181 (N_9181,N_4192,N_5042);
and U9182 (N_9182,N_5355,N_1801);
nor U9183 (N_9183,N_5589,N_4534);
and U9184 (N_9184,N_5105,N_1630);
nor U9185 (N_9185,N_290,N_3869);
or U9186 (N_9186,N_5974,N_2772);
nor U9187 (N_9187,N_4138,N_1376);
and U9188 (N_9188,N_1679,N_3146);
nand U9189 (N_9189,N_3162,N_4600);
or U9190 (N_9190,N_5907,N_3146);
nor U9191 (N_9191,N_5206,N_2045);
or U9192 (N_9192,N_3307,N_2280);
xor U9193 (N_9193,N_1458,N_95);
or U9194 (N_9194,N_861,N_486);
and U9195 (N_9195,N_5998,N_4603);
nor U9196 (N_9196,N_5494,N_3058);
nand U9197 (N_9197,N_801,N_5894);
or U9198 (N_9198,N_1601,N_4741);
or U9199 (N_9199,N_4859,N_5870);
nor U9200 (N_9200,N_3834,N_3224);
xor U9201 (N_9201,N_2982,N_5399);
and U9202 (N_9202,N_3941,N_2476);
and U9203 (N_9203,N_1726,N_1105);
nand U9204 (N_9204,N_4841,N_1629);
nor U9205 (N_9205,N_2501,N_5786);
or U9206 (N_9206,N_1829,N_954);
nor U9207 (N_9207,N_3545,N_1263);
or U9208 (N_9208,N_498,N_4070);
and U9209 (N_9209,N_3394,N_2623);
nor U9210 (N_9210,N_510,N_744);
or U9211 (N_9211,N_4784,N_5579);
or U9212 (N_9212,N_2323,N_2681);
nand U9213 (N_9213,N_4690,N_2799);
xnor U9214 (N_9214,N_54,N_2179);
nor U9215 (N_9215,N_5882,N_4886);
xor U9216 (N_9216,N_4599,N_1737);
xor U9217 (N_9217,N_4735,N_3583);
or U9218 (N_9218,N_1709,N_5629);
or U9219 (N_9219,N_5212,N_4042);
nand U9220 (N_9220,N_233,N_3358);
and U9221 (N_9221,N_1352,N_3746);
nand U9222 (N_9222,N_4261,N_1991);
or U9223 (N_9223,N_3907,N_4476);
and U9224 (N_9224,N_1240,N_4645);
xor U9225 (N_9225,N_855,N_135);
xnor U9226 (N_9226,N_1019,N_4795);
nor U9227 (N_9227,N_1653,N_1735);
nand U9228 (N_9228,N_2502,N_3011);
or U9229 (N_9229,N_2734,N_5083);
or U9230 (N_9230,N_2330,N_2092);
xnor U9231 (N_9231,N_4000,N_4520);
or U9232 (N_9232,N_1219,N_479);
xor U9233 (N_9233,N_164,N_235);
or U9234 (N_9234,N_4419,N_4440);
xnor U9235 (N_9235,N_2392,N_165);
nand U9236 (N_9236,N_5255,N_1932);
or U9237 (N_9237,N_5005,N_3884);
nor U9238 (N_9238,N_1662,N_1913);
nor U9239 (N_9239,N_558,N_4954);
nor U9240 (N_9240,N_3561,N_2357);
nor U9241 (N_9241,N_5118,N_4781);
nand U9242 (N_9242,N_2762,N_2219);
nor U9243 (N_9243,N_1168,N_4637);
and U9244 (N_9244,N_3454,N_5089);
nor U9245 (N_9245,N_446,N_1166);
xor U9246 (N_9246,N_5390,N_4441);
nor U9247 (N_9247,N_121,N_672);
or U9248 (N_9248,N_232,N_2147);
or U9249 (N_9249,N_1330,N_683);
xor U9250 (N_9250,N_4357,N_2242);
and U9251 (N_9251,N_517,N_2436);
nand U9252 (N_9252,N_4125,N_4280);
and U9253 (N_9253,N_2595,N_1725);
and U9254 (N_9254,N_3885,N_2482);
nand U9255 (N_9255,N_367,N_1609);
xor U9256 (N_9256,N_2152,N_4902);
nand U9257 (N_9257,N_4030,N_229);
nand U9258 (N_9258,N_1607,N_485);
xor U9259 (N_9259,N_4781,N_5514);
xnor U9260 (N_9260,N_5182,N_90);
and U9261 (N_9261,N_2191,N_5442);
nor U9262 (N_9262,N_5197,N_4460);
xor U9263 (N_9263,N_5312,N_2058);
and U9264 (N_9264,N_5353,N_5509);
or U9265 (N_9265,N_2519,N_675);
and U9266 (N_9266,N_3225,N_1590);
xnor U9267 (N_9267,N_2387,N_2788);
and U9268 (N_9268,N_3149,N_2061);
and U9269 (N_9269,N_5448,N_2149);
or U9270 (N_9270,N_1775,N_2301);
and U9271 (N_9271,N_1498,N_2263);
and U9272 (N_9272,N_69,N_2287);
nor U9273 (N_9273,N_1807,N_130);
and U9274 (N_9274,N_5488,N_5941);
and U9275 (N_9275,N_634,N_3975);
nor U9276 (N_9276,N_4114,N_819);
and U9277 (N_9277,N_3042,N_2736);
nand U9278 (N_9278,N_3005,N_3667);
nand U9279 (N_9279,N_4776,N_5719);
xor U9280 (N_9280,N_3843,N_4927);
nand U9281 (N_9281,N_2363,N_565);
nand U9282 (N_9282,N_3915,N_1481);
nor U9283 (N_9283,N_4260,N_1686);
xnor U9284 (N_9284,N_3759,N_4304);
nand U9285 (N_9285,N_5225,N_5419);
nor U9286 (N_9286,N_4095,N_2612);
and U9287 (N_9287,N_2002,N_2166);
nand U9288 (N_9288,N_5636,N_2490);
and U9289 (N_9289,N_2109,N_215);
and U9290 (N_9290,N_3679,N_5960);
or U9291 (N_9291,N_5436,N_1845);
nor U9292 (N_9292,N_4576,N_3231);
nand U9293 (N_9293,N_5606,N_4117);
nor U9294 (N_9294,N_3663,N_3430);
nor U9295 (N_9295,N_1598,N_5925);
or U9296 (N_9296,N_2846,N_1802);
nand U9297 (N_9297,N_2475,N_3659);
nand U9298 (N_9298,N_5562,N_3799);
nand U9299 (N_9299,N_2145,N_2754);
xor U9300 (N_9300,N_5242,N_4121);
nor U9301 (N_9301,N_1602,N_1673);
nor U9302 (N_9302,N_5772,N_1444);
and U9303 (N_9303,N_2803,N_1429);
nor U9304 (N_9304,N_2800,N_27);
or U9305 (N_9305,N_295,N_4258);
nor U9306 (N_9306,N_3002,N_604);
nor U9307 (N_9307,N_4977,N_2556);
or U9308 (N_9308,N_773,N_2074);
nor U9309 (N_9309,N_3760,N_2617);
nor U9310 (N_9310,N_1560,N_123);
or U9311 (N_9311,N_5390,N_3145);
nor U9312 (N_9312,N_5266,N_4883);
nand U9313 (N_9313,N_3533,N_1406);
xnor U9314 (N_9314,N_1113,N_3968);
and U9315 (N_9315,N_1878,N_5650);
nor U9316 (N_9316,N_1341,N_3360);
or U9317 (N_9317,N_3443,N_5314);
or U9318 (N_9318,N_1610,N_1810);
or U9319 (N_9319,N_4840,N_4462);
xnor U9320 (N_9320,N_1858,N_1553);
or U9321 (N_9321,N_5745,N_2083);
and U9322 (N_9322,N_1323,N_1898);
xnor U9323 (N_9323,N_1201,N_3612);
nor U9324 (N_9324,N_1474,N_4242);
nand U9325 (N_9325,N_3904,N_5896);
xnor U9326 (N_9326,N_3950,N_2972);
xnor U9327 (N_9327,N_1197,N_4130);
nand U9328 (N_9328,N_4046,N_2590);
and U9329 (N_9329,N_4265,N_3526);
nand U9330 (N_9330,N_1950,N_5511);
nor U9331 (N_9331,N_934,N_151);
and U9332 (N_9332,N_2085,N_3049);
xor U9333 (N_9333,N_4379,N_3354);
nor U9334 (N_9334,N_5920,N_5912);
nor U9335 (N_9335,N_5255,N_3220);
nor U9336 (N_9336,N_1295,N_959);
nor U9337 (N_9337,N_3764,N_1994);
nand U9338 (N_9338,N_89,N_3692);
or U9339 (N_9339,N_1972,N_3983);
and U9340 (N_9340,N_460,N_5740);
and U9341 (N_9341,N_3167,N_1600);
or U9342 (N_9342,N_3977,N_2531);
or U9343 (N_9343,N_4938,N_5976);
nand U9344 (N_9344,N_3486,N_4873);
or U9345 (N_9345,N_5272,N_3267);
nor U9346 (N_9346,N_1559,N_3986);
and U9347 (N_9347,N_555,N_4371);
and U9348 (N_9348,N_3023,N_3430);
nor U9349 (N_9349,N_1707,N_3735);
or U9350 (N_9350,N_137,N_3347);
or U9351 (N_9351,N_1366,N_2498);
nor U9352 (N_9352,N_1982,N_2349);
nor U9353 (N_9353,N_3048,N_1862);
nand U9354 (N_9354,N_1001,N_905);
xor U9355 (N_9355,N_4471,N_2730);
nor U9356 (N_9356,N_3528,N_4735);
or U9357 (N_9357,N_3114,N_5944);
or U9358 (N_9358,N_3682,N_843);
and U9359 (N_9359,N_1010,N_52);
xor U9360 (N_9360,N_397,N_4120);
xnor U9361 (N_9361,N_3295,N_3820);
xnor U9362 (N_9362,N_3948,N_2913);
nand U9363 (N_9363,N_5259,N_2864);
and U9364 (N_9364,N_4745,N_2681);
xnor U9365 (N_9365,N_5506,N_430);
xnor U9366 (N_9366,N_776,N_537);
and U9367 (N_9367,N_5700,N_3416);
nand U9368 (N_9368,N_1654,N_3472);
or U9369 (N_9369,N_1093,N_1060);
nor U9370 (N_9370,N_218,N_2479);
or U9371 (N_9371,N_4877,N_5317);
or U9372 (N_9372,N_3974,N_4108);
and U9373 (N_9373,N_1489,N_445);
nand U9374 (N_9374,N_4278,N_3350);
xnor U9375 (N_9375,N_142,N_3892);
nand U9376 (N_9376,N_348,N_5133);
or U9377 (N_9377,N_3273,N_5785);
or U9378 (N_9378,N_5144,N_5272);
or U9379 (N_9379,N_573,N_5185);
nand U9380 (N_9380,N_1415,N_4727);
or U9381 (N_9381,N_4438,N_4649);
nand U9382 (N_9382,N_309,N_3812);
xor U9383 (N_9383,N_5423,N_979);
nand U9384 (N_9384,N_1070,N_1448);
or U9385 (N_9385,N_1983,N_126);
or U9386 (N_9386,N_621,N_1076);
and U9387 (N_9387,N_1711,N_3335);
nand U9388 (N_9388,N_4421,N_4349);
or U9389 (N_9389,N_4626,N_4253);
and U9390 (N_9390,N_5036,N_5782);
xnor U9391 (N_9391,N_2207,N_1109);
and U9392 (N_9392,N_1584,N_664);
or U9393 (N_9393,N_3755,N_842);
nor U9394 (N_9394,N_2776,N_4408);
nand U9395 (N_9395,N_4771,N_2016);
or U9396 (N_9396,N_5696,N_4640);
and U9397 (N_9397,N_3132,N_2334);
nand U9398 (N_9398,N_1069,N_1283);
xnor U9399 (N_9399,N_2455,N_4175);
nand U9400 (N_9400,N_5120,N_4917);
xnor U9401 (N_9401,N_3732,N_2055);
xor U9402 (N_9402,N_1377,N_2422);
or U9403 (N_9403,N_3125,N_3373);
nand U9404 (N_9404,N_802,N_4933);
nand U9405 (N_9405,N_2966,N_3565);
xnor U9406 (N_9406,N_691,N_3877);
or U9407 (N_9407,N_1091,N_1370);
or U9408 (N_9408,N_4088,N_1659);
and U9409 (N_9409,N_4827,N_2269);
and U9410 (N_9410,N_1223,N_2242);
or U9411 (N_9411,N_5987,N_801);
nor U9412 (N_9412,N_5877,N_2505);
nand U9413 (N_9413,N_5166,N_1637);
xor U9414 (N_9414,N_1955,N_5878);
and U9415 (N_9415,N_3317,N_503);
and U9416 (N_9416,N_4816,N_391);
nand U9417 (N_9417,N_2956,N_4423);
nand U9418 (N_9418,N_4763,N_2819);
xor U9419 (N_9419,N_1375,N_329);
or U9420 (N_9420,N_1713,N_1404);
or U9421 (N_9421,N_1821,N_4453);
or U9422 (N_9422,N_1758,N_5652);
or U9423 (N_9423,N_2712,N_4540);
nor U9424 (N_9424,N_297,N_1764);
nand U9425 (N_9425,N_4658,N_2096);
and U9426 (N_9426,N_1797,N_1038);
or U9427 (N_9427,N_3747,N_4145);
nor U9428 (N_9428,N_3685,N_4373);
xor U9429 (N_9429,N_4190,N_1016);
and U9430 (N_9430,N_5342,N_1173);
and U9431 (N_9431,N_3859,N_672);
nor U9432 (N_9432,N_632,N_3944);
nand U9433 (N_9433,N_3164,N_4060);
xnor U9434 (N_9434,N_4751,N_1706);
xor U9435 (N_9435,N_1570,N_573);
xor U9436 (N_9436,N_3079,N_2822);
xor U9437 (N_9437,N_2654,N_4414);
nand U9438 (N_9438,N_5377,N_4188);
nor U9439 (N_9439,N_1919,N_1645);
xor U9440 (N_9440,N_5539,N_647);
or U9441 (N_9441,N_2186,N_2032);
or U9442 (N_9442,N_317,N_1149);
and U9443 (N_9443,N_4022,N_274);
and U9444 (N_9444,N_3100,N_3797);
nand U9445 (N_9445,N_3102,N_4330);
nor U9446 (N_9446,N_2984,N_4440);
nor U9447 (N_9447,N_783,N_1159);
nand U9448 (N_9448,N_1970,N_182);
and U9449 (N_9449,N_5856,N_5251);
or U9450 (N_9450,N_2157,N_4750);
and U9451 (N_9451,N_2860,N_1913);
or U9452 (N_9452,N_3610,N_5096);
nand U9453 (N_9453,N_1043,N_4128);
xnor U9454 (N_9454,N_4904,N_1217);
nand U9455 (N_9455,N_2884,N_104);
or U9456 (N_9456,N_2412,N_4230);
or U9457 (N_9457,N_5215,N_1894);
xnor U9458 (N_9458,N_117,N_1632);
and U9459 (N_9459,N_867,N_1115);
and U9460 (N_9460,N_5327,N_5646);
nor U9461 (N_9461,N_4821,N_1991);
nand U9462 (N_9462,N_986,N_1363);
or U9463 (N_9463,N_3941,N_1930);
and U9464 (N_9464,N_5523,N_4781);
nand U9465 (N_9465,N_3724,N_689);
or U9466 (N_9466,N_5769,N_2999);
nor U9467 (N_9467,N_3478,N_5434);
or U9468 (N_9468,N_4683,N_2564);
or U9469 (N_9469,N_367,N_4520);
xnor U9470 (N_9470,N_5095,N_2935);
nor U9471 (N_9471,N_2359,N_3180);
nand U9472 (N_9472,N_4223,N_5860);
and U9473 (N_9473,N_1138,N_1432);
nor U9474 (N_9474,N_5530,N_870);
and U9475 (N_9475,N_369,N_4836);
or U9476 (N_9476,N_302,N_2395);
and U9477 (N_9477,N_5975,N_2559);
nor U9478 (N_9478,N_4715,N_1785);
xor U9479 (N_9479,N_2032,N_1619);
nor U9480 (N_9480,N_3815,N_4143);
xor U9481 (N_9481,N_3575,N_4168);
nor U9482 (N_9482,N_5411,N_5555);
or U9483 (N_9483,N_5035,N_2003);
nor U9484 (N_9484,N_3191,N_1869);
or U9485 (N_9485,N_3305,N_1790);
xor U9486 (N_9486,N_1440,N_4823);
xnor U9487 (N_9487,N_553,N_1388);
xor U9488 (N_9488,N_5693,N_5264);
or U9489 (N_9489,N_5341,N_152);
or U9490 (N_9490,N_950,N_398);
or U9491 (N_9491,N_2743,N_383);
xor U9492 (N_9492,N_3535,N_1009);
or U9493 (N_9493,N_1429,N_3713);
nand U9494 (N_9494,N_5214,N_3036);
nand U9495 (N_9495,N_5376,N_5318);
xnor U9496 (N_9496,N_2124,N_2238);
or U9497 (N_9497,N_3099,N_5769);
nand U9498 (N_9498,N_2551,N_2142);
nor U9499 (N_9499,N_900,N_4848);
and U9500 (N_9500,N_4563,N_176);
and U9501 (N_9501,N_939,N_675);
and U9502 (N_9502,N_3350,N_5600);
xnor U9503 (N_9503,N_4030,N_13);
and U9504 (N_9504,N_1799,N_3904);
nand U9505 (N_9505,N_4568,N_5347);
nand U9506 (N_9506,N_4375,N_2745);
xor U9507 (N_9507,N_2319,N_4929);
and U9508 (N_9508,N_4876,N_3436);
nor U9509 (N_9509,N_1676,N_5627);
nor U9510 (N_9510,N_920,N_4911);
xnor U9511 (N_9511,N_4153,N_336);
or U9512 (N_9512,N_4518,N_2486);
nor U9513 (N_9513,N_4453,N_4940);
or U9514 (N_9514,N_4171,N_3367);
xnor U9515 (N_9515,N_5558,N_2423);
nor U9516 (N_9516,N_670,N_5366);
nand U9517 (N_9517,N_2528,N_83);
and U9518 (N_9518,N_5910,N_50);
nand U9519 (N_9519,N_4016,N_3593);
and U9520 (N_9520,N_4425,N_4611);
xor U9521 (N_9521,N_2027,N_4039);
nor U9522 (N_9522,N_1072,N_364);
nand U9523 (N_9523,N_2938,N_5015);
nor U9524 (N_9524,N_2672,N_2379);
xor U9525 (N_9525,N_671,N_3743);
nand U9526 (N_9526,N_3916,N_2804);
nand U9527 (N_9527,N_5384,N_2596);
nor U9528 (N_9528,N_1957,N_2694);
and U9529 (N_9529,N_5829,N_2674);
nand U9530 (N_9530,N_1074,N_4199);
or U9531 (N_9531,N_2335,N_2306);
nor U9532 (N_9532,N_3802,N_187);
nor U9533 (N_9533,N_2150,N_2797);
and U9534 (N_9534,N_3708,N_754);
or U9535 (N_9535,N_842,N_4759);
nand U9536 (N_9536,N_2975,N_4923);
nand U9537 (N_9537,N_5021,N_1390);
nand U9538 (N_9538,N_247,N_5235);
and U9539 (N_9539,N_1922,N_1968);
xnor U9540 (N_9540,N_3084,N_2814);
nand U9541 (N_9541,N_5984,N_1139);
nor U9542 (N_9542,N_3738,N_152);
xor U9543 (N_9543,N_3464,N_4758);
nor U9544 (N_9544,N_3687,N_2507);
nor U9545 (N_9545,N_61,N_5115);
or U9546 (N_9546,N_2400,N_291);
nand U9547 (N_9547,N_424,N_5261);
xnor U9548 (N_9548,N_5196,N_4542);
xnor U9549 (N_9549,N_2959,N_678);
nor U9550 (N_9550,N_3058,N_873);
nor U9551 (N_9551,N_5679,N_2633);
xor U9552 (N_9552,N_2492,N_2721);
nor U9553 (N_9553,N_4303,N_3335);
nand U9554 (N_9554,N_1881,N_4870);
or U9555 (N_9555,N_3427,N_4514);
nand U9556 (N_9556,N_608,N_5172);
nand U9557 (N_9557,N_5229,N_934);
xnor U9558 (N_9558,N_3446,N_5723);
or U9559 (N_9559,N_5091,N_2037);
nand U9560 (N_9560,N_4277,N_1598);
nand U9561 (N_9561,N_1413,N_2122);
nand U9562 (N_9562,N_3957,N_2273);
and U9563 (N_9563,N_2396,N_3865);
or U9564 (N_9564,N_1740,N_1247);
nor U9565 (N_9565,N_1617,N_2441);
xnor U9566 (N_9566,N_5584,N_2227);
nor U9567 (N_9567,N_5491,N_631);
nand U9568 (N_9568,N_3959,N_2563);
or U9569 (N_9569,N_563,N_4882);
xnor U9570 (N_9570,N_5479,N_5836);
or U9571 (N_9571,N_1599,N_269);
nand U9572 (N_9572,N_1626,N_5120);
nand U9573 (N_9573,N_3857,N_1008);
and U9574 (N_9574,N_668,N_5319);
or U9575 (N_9575,N_2827,N_574);
xnor U9576 (N_9576,N_2126,N_1653);
nand U9577 (N_9577,N_3542,N_5924);
xnor U9578 (N_9578,N_4595,N_123);
nand U9579 (N_9579,N_5500,N_3117);
nor U9580 (N_9580,N_2646,N_5735);
xor U9581 (N_9581,N_2410,N_175);
nor U9582 (N_9582,N_4051,N_5393);
xor U9583 (N_9583,N_4314,N_246);
and U9584 (N_9584,N_526,N_1885);
nand U9585 (N_9585,N_2196,N_333);
and U9586 (N_9586,N_129,N_2061);
and U9587 (N_9587,N_3568,N_575);
xnor U9588 (N_9588,N_4514,N_2865);
xor U9589 (N_9589,N_968,N_1223);
xnor U9590 (N_9590,N_4194,N_2067);
xnor U9591 (N_9591,N_1252,N_149);
nor U9592 (N_9592,N_3020,N_1565);
or U9593 (N_9593,N_3063,N_1395);
xor U9594 (N_9594,N_2538,N_4373);
or U9595 (N_9595,N_836,N_3855);
xor U9596 (N_9596,N_2719,N_104);
or U9597 (N_9597,N_1704,N_929);
nand U9598 (N_9598,N_849,N_2078);
nand U9599 (N_9599,N_4218,N_4313);
or U9600 (N_9600,N_3929,N_5455);
xor U9601 (N_9601,N_3894,N_1493);
xnor U9602 (N_9602,N_4051,N_58);
nand U9603 (N_9603,N_3865,N_873);
nor U9604 (N_9604,N_2972,N_1214);
nand U9605 (N_9605,N_4165,N_2348);
nor U9606 (N_9606,N_5383,N_1785);
nand U9607 (N_9607,N_3269,N_824);
and U9608 (N_9608,N_1983,N_3940);
nor U9609 (N_9609,N_4943,N_653);
nor U9610 (N_9610,N_5978,N_2955);
nand U9611 (N_9611,N_3697,N_3417);
or U9612 (N_9612,N_3228,N_3725);
and U9613 (N_9613,N_4256,N_920);
and U9614 (N_9614,N_5974,N_255);
or U9615 (N_9615,N_1544,N_5777);
or U9616 (N_9616,N_5532,N_4779);
nand U9617 (N_9617,N_1329,N_3698);
and U9618 (N_9618,N_376,N_82);
nand U9619 (N_9619,N_2555,N_4480);
xnor U9620 (N_9620,N_3896,N_3105);
or U9621 (N_9621,N_1687,N_630);
and U9622 (N_9622,N_844,N_5869);
or U9623 (N_9623,N_5663,N_2050);
or U9624 (N_9624,N_2924,N_1705);
and U9625 (N_9625,N_592,N_3829);
or U9626 (N_9626,N_412,N_136);
nor U9627 (N_9627,N_276,N_4044);
or U9628 (N_9628,N_5003,N_1220);
xnor U9629 (N_9629,N_2101,N_2350);
nand U9630 (N_9630,N_4573,N_4095);
and U9631 (N_9631,N_1696,N_3102);
nand U9632 (N_9632,N_5131,N_2581);
nand U9633 (N_9633,N_1710,N_485);
and U9634 (N_9634,N_3147,N_1282);
or U9635 (N_9635,N_2223,N_1074);
nand U9636 (N_9636,N_3504,N_607);
or U9637 (N_9637,N_2758,N_3363);
and U9638 (N_9638,N_5811,N_3954);
or U9639 (N_9639,N_169,N_833);
or U9640 (N_9640,N_3910,N_556);
and U9641 (N_9641,N_2238,N_5010);
nand U9642 (N_9642,N_3946,N_5862);
or U9643 (N_9643,N_4154,N_4839);
nand U9644 (N_9644,N_4141,N_4502);
nor U9645 (N_9645,N_2917,N_1015);
or U9646 (N_9646,N_1745,N_2273);
or U9647 (N_9647,N_3188,N_2177);
or U9648 (N_9648,N_3986,N_4437);
or U9649 (N_9649,N_4449,N_5383);
nor U9650 (N_9650,N_2019,N_1333);
xor U9651 (N_9651,N_5680,N_1231);
nor U9652 (N_9652,N_745,N_2524);
xnor U9653 (N_9653,N_1319,N_2684);
and U9654 (N_9654,N_5044,N_5158);
xor U9655 (N_9655,N_5525,N_5283);
nor U9656 (N_9656,N_1055,N_1411);
xor U9657 (N_9657,N_3101,N_567);
and U9658 (N_9658,N_5816,N_3853);
nand U9659 (N_9659,N_5012,N_2371);
or U9660 (N_9660,N_1985,N_2736);
and U9661 (N_9661,N_11,N_1059);
nor U9662 (N_9662,N_272,N_3423);
or U9663 (N_9663,N_1312,N_3656);
nand U9664 (N_9664,N_3057,N_2807);
nor U9665 (N_9665,N_127,N_5053);
nand U9666 (N_9666,N_747,N_425);
and U9667 (N_9667,N_3315,N_2096);
nor U9668 (N_9668,N_2601,N_3984);
nor U9669 (N_9669,N_5515,N_1213);
xnor U9670 (N_9670,N_4366,N_291);
nand U9671 (N_9671,N_93,N_2182);
nand U9672 (N_9672,N_4379,N_1480);
nor U9673 (N_9673,N_3101,N_1753);
and U9674 (N_9674,N_2332,N_791);
nand U9675 (N_9675,N_5447,N_1878);
or U9676 (N_9676,N_142,N_5100);
and U9677 (N_9677,N_3300,N_353);
xor U9678 (N_9678,N_1064,N_2840);
nor U9679 (N_9679,N_5445,N_4155);
xnor U9680 (N_9680,N_1808,N_479);
xnor U9681 (N_9681,N_481,N_2705);
and U9682 (N_9682,N_4972,N_1935);
xnor U9683 (N_9683,N_397,N_1627);
nand U9684 (N_9684,N_4152,N_3400);
or U9685 (N_9685,N_1850,N_730);
or U9686 (N_9686,N_2280,N_438);
and U9687 (N_9687,N_2022,N_4477);
nor U9688 (N_9688,N_624,N_5151);
nor U9689 (N_9689,N_2248,N_362);
or U9690 (N_9690,N_1525,N_263);
and U9691 (N_9691,N_5185,N_5611);
nor U9692 (N_9692,N_3603,N_5145);
nand U9693 (N_9693,N_3295,N_3144);
nor U9694 (N_9694,N_3295,N_1975);
and U9695 (N_9695,N_5512,N_1589);
or U9696 (N_9696,N_3419,N_1768);
and U9697 (N_9697,N_4236,N_779);
and U9698 (N_9698,N_3608,N_2807);
nand U9699 (N_9699,N_2903,N_2322);
nand U9700 (N_9700,N_4301,N_2920);
xnor U9701 (N_9701,N_345,N_680);
or U9702 (N_9702,N_1817,N_16);
nor U9703 (N_9703,N_4518,N_5286);
xor U9704 (N_9704,N_5096,N_1531);
or U9705 (N_9705,N_5627,N_1431);
and U9706 (N_9706,N_3414,N_5692);
and U9707 (N_9707,N_2708,N_2353);
xor U9708 (N_9708,N_1161,N_1584);
xnor U9709 (N_9709,N_5707,N_2128);
nor U9710 (N_9710,N_2580,N_1988);
or U9711 (N_9711,N_4624,N_5329);
nand U9712 (N_9712,N_2179,N_5159);
and U9713 (N_9713,N_3712,N_5513);
and U9714 (N_9714,N_1104,N_4463);
and U9715 (N_9715,N_3362,N_4023);
and U9716 (N_9716,N_4927,N_1374);
nor U9717 (N_9717,N_4593,N_2643);
and U9718 (N_9718,N_2335,N_4225);
nand U9719 (N_9719,N_2838,N_4558);
or U9720 (N_9720,N_2392,N_2115);
nand U9721 (N_9721,N_3824,N_3187);
nor U9722 (N_9722,N_5806,N_5171);
and U9723 (N_9723,N_3669,N_2430);
nor U9724 (N_9724,N_845,N_3744);
xnor U9725 (N_9725,N_2975,N_268);
or U9726 (N_9726,N_3258,N_187);
xor U9727 (N_9727,N_5600,N_4017);
and U9728 (N_9728,N_104,N_831);
nor U9729 (N_9729,N_5097,N_266);
and U9730 (N_9730,N_5947,N_1117);
nor U9731 (N_9731,N_4956,N_2746);
nor U9732 (N_9732,N_376,N_5374);
xnor U9733 (N_9733,N_4429,N_2152);
and U9734 (N_9734,N_1858,N_1269);
nand U9735 (N_9735,N_2983,N_3332);
or U9736 (N_9736,N_3008,N_2883);
and U9737 (N_9737,N_1126,N_1235);
or U9738 (N_9738,N_1484,N_329);
nor U9739 (N_9739,N_1083,N_3616);
and U9740 (N_9740,N_4414,N_4387);
xnor U9741 (N_9741,N_4883,N_2109);
nand U9742 (N_9742,N_4565,N_4709);
and U9743 (N_9743,N_3423,N_1217);
or U9744 (N_9744,N_1679,N_2858);
nor U9745 (N_9745,N_3554,N_5996);
and U9746 (N_9746,N_3070,N_3782);
nor U9747 (N_9747,N_2166,N_4550);
xor U9748 (N_9748,N_1785,N_5061);
or U9749 (N_9749,N_4894,N_3600);
xor U9750 (N_9750,N_5946,N_2114);
xnor U9751 (N_9751,N_2831,N_3516);
and U9752 (N_9752,N_5036,N_5500);
nor U9753 (N_9753,N_2548,N_4709);
nand U9754 (N_9754,N_4239,N_653);
xnor U9755 (N_9755,N_4095,N_1644);
and U9756 (N_9756,N_1498,N_1794);
xnor U9757 (N_9757,N_29,N_4169);
or U9758 (N_9758,N_2440,N_949);
and U9759 (N_9759,N_4662,N_1911);
or U9760 (N_9760,N_5980,N_3442);
xnor U9761 (N_9761,N_5835,N_4215);
nand U9762 (N_9762,N_2957,N_92);
nand U9763 (N_9763,N_4922,N_1396);
or U9764 (N_9764,N_2590,N_4341);
xor U9765 (N_9765,N_4509,N_4255);
or U9766 (N_9766,N_2201,N_498);
nand U9767 (N_9767,N_782,N_4187);
and U9768 (N_9768,N_2782,N_4622);
nor U9769 (N_9769,N_4213,N_4951);
xor U9770 (N_9770,N_2330,N_4302);
nand U9771 (N_9771,N_4302,N_4863);
or U9772 (N_9772,N_2049,N_2320);
or U9773 (N_9773,N_5161,N_4692);
nand U9774 (N_9774,N_2122,N_3170);
nor U9775 (N_9775,N_2439,N_5294);
xor U9776 (N_9776,N_1259,N_934);
and U9777 (N_9777,N_660,N_5849);
or U9778 (N_9778,N_4982,N_2793);
xnor U9779 (N_9779,N_4861,N_1229);
or U9780 (N_9780,N_508,N_2161);
nor U9781 (N_9781,N_5806,N_510);
nand U9782 (N_9782,N_1030,N_5471);
and U9783 (N_9783,N_4724,N_3288);
nand U9784 (N_9784,N_281,N_3294);
and U9785 (N_9785,N_4302,N_1244);
nand U9786 (N_9786,N_1449,N_226);
nand U9787 (N_9787,N_159,N_3321);
or U9788 (N_9788,N_3205,N_4199);
nor U9789 (N_9789,N_31,N_187);
nand U9790 (N_9790,N_1559,N_2446);
and U9791 (N_9791,N_120,N_1344);
or U9792 (N_9792,N_3292,N_2725);
and U9793 (N_9793,N_2184,N_5559);
nor U9794 (N_9794,N_2087,N_4328);
xnor U9795 (N_9795,N_4177,N_1422);
nor U9796 (N_9796,N_4677,N_1363);
xor U9797 (N_9797,N_4161,N_1003);
nand U9798 (N_9798,N_3023,N_3440);
nand U9799 (N_9799,N_4010,N_3470);
or U9800 (N_9800,N_280,N_5841);
nand U9801 (N_9801,N_4681,N_1999);
and U9802 (N_9802,N_5499,N_1098);
xnor U9803 (N_9803,N_3836,N_1082);
xor U9804 (N_9804,N_1866,N_4118);
nand U9805 (N_9805,N_1272,N_5734);
nor U9806 (N_9806,N_3751,N_1669);
nor U9807 (N_9807,N_4820,N_2798);
xor U9808 (N_9808,N_1815,N_422);
nor U9809 (N_9809,N_3651,N_2198);
nand U9810 (N_9810,N_5592,N_5013);
xnor U9811 (N_9811,N_5951,N_2301);
xnor U9812 (N_9812,N_4444,N_5744);
nand U9813 (N_9813,N_2465,N_1624);
or U9814 (N_9814,N_3133,N_181);
xnor U9815 (N_9815,N_4999,N_3570);
or U9816 (N_9816,N_4121,N_3044);
nor U9817 (N_9817,N_2661,N_2485);
nor U9818 (N_9818,N_399,N_5984);
xnor U9819 (N_9819,N_153,N_2839);
xor U9820 (N_9820,N_934,N_152);
xor U9821 (N_9821,N_130,N_5301);
and U9822 (N_9822,N_559,N_96);
and U9823 (N_9823,N_2009,N_4299);
nor U9824 (N_9824,N_4768,N_1995);
nand U9825 (N_9825,N_2475,N_3056);
nor U9826 (N_9826,N_3625,N_1137);
nand U9827 (N_9827,N_248,N_5030);
xor U9828 (N_9828,N_1711,N_5639);
and U9829 (N_9829,N_3039,N_1361);
nor U9830 (N_9830,N_5302,N_5797);
and U9831 (N_9831,N_1800,N_1729);
or U9832 (N_9832,N_4324,N_1012);
and U9833 (N_9833,N_1604,N_3430);
nand U9834 (N_9834,N_4362,N_1977);
nor U9835 (N_9835,N_2059,N_4603);
or U9836 (N_9836,N_978,N_2342);
nand U9837 (N_9837,N_668,N_948);
or U9838 (N_9838,N_5187,N_14);
nand U9839 (N_9839,N_4791,N_1471);
or U9840 (N_9840,N_4949,N_3610);
or U9841 (N_9841,N_5614,N_3327);
nor U9842 (N_9842,N_5202,N_5);
and U9843 (N_9843,N_4082,N_3832);
or U9844 (N_9844,N_3462,N_919);
or U9845 (N_9845,N_5711,N_4351);
or U9846 (N_9846,N_3286,N_5629);
or U9847 (N_9847,N_4012,N_27);
nand U9848 (N_9848,N_60,N_4519);
nand U9849 (N_9849,N_3508,N_2656);
or U9850 (N_9850,N_1902,N_1282);
or U9851 (N_9851,N_2726,N_2184);
or U9852 (N_9852,N_2557,N_1879);
or U9853 (N_9853,N_5037,N_4181);
xor U9854 (N_9854,N_3893,N_976);
and U9855 (N_9855,N_3856,N_3522);
or U9856 (N_9856,N_502,N_1816);
nand U9857 (N_9857,N_3228,N_4672);
and U9858 (N_9858,N_3679,N_678);
or U9859 (N_9859,N_747,N_4154);
or U9860 (N_9860,N_2553,N_1323);
or U9861 (N_9861,N_733,N_5600);
xor U9862 (N_9862,N_2205,N_3565);
xor U9863 (N_9863,N_978,N_4133);
nor U9864 (N_9864,N_5803,N_1661);
xnor U9865 (N_9865,N_585,N_5131);
xor U9866 (N_9866,N_5616,N_2253);
or U9867 (N_9867,N_3677,N_1548);
and U9868 (N_9868,N_419,N_5931);
or U9869 (N_9869,N_436,N_2207);
nor U9870 (N_9870,N_1966,N_1675);
nand U9871 (N_9871,N_590,N_544);
nor U9872 (N_9872,N_830,N_608);
xnor U9873 (N_9873,N_1884,N_5515);
nor U9874 (N_9874,N_5162,N_2130);
or U9875 (N_9875,N_4720,N_596);
nor U9876 (N_9876,N_82,N_5666);
nor U9877 (N_9877,N_3415,N_581);
and U9878 (N_9878,N_2102,N_5278);
or U9879 (N_9879,N_3963,N_1485);
nor U9880 (N_9880,N_1450,N_5105);
or U9881 (N_9881,N_5545,N_797);
xnor U9882 (N_9882,N_3169,N_5249);
and U9883 (N_9883,N_37,N_3702);
and U9884 (N_9884,N_2542,N_2652);
and U9885 (N_9885,N_5308,N_5169);
and U9886 (N_9886,N_4610,N_2676);
xnor U9887 (N_9887,N_1455,N_5199);
nor U9888 (N_9888,N_1347,N_428);
and U9889 (N_9889,N_4651,N_2615);
nand U9890 (N_9890,N_4331,N_903);
and U9891 (N_9891,N_4091,N_4411);
nor U9892 (N_9892,N_3167,N_761);
and U9893 (N_9893,N_1215,N_4856);
or U9894 (N_9894,N_2226,N_5511);
nor U9895 (N_9895,N_103,N_5805);
or U9896 (N_9896,N_1305,N_1217);
or U9897 (N_9897,N_1472,N_403);
nor U9898 (N_9898,N_1567,N_3097);
or U9899 (N_9899,N_5563,N_5406);
or U9900 (N_9900,N_3931,N_1993);
or U9901 (N_9901,N_2839,N_3704);
or U9902 (N_9902,N_4777,N_740);
or U9903 (N_9903,N_1005,N_1097);
nor U9904 (N_9904,N_3114,N_2881);
nand U9905 (N_9905,N_3258,N_674);
nor U9906 (N_9906,N_1637,N_916);
nor U9907 (N_9907,N_5077,N_3978);
xor U9908 (N_9908,N_2497,N_1726);
nor U9909 (N_9909,N_43,N_768);
nand U9910 (N_9910,N_5897,N_2786);
or U9911 (N_9911,N_4640,N_5882);
nor U9912 (N_9912,N_4156,N_3193);
xor U9913 (N_9913,N_442,N_5828);
nand U9914 (N_9914,N_1599,N_2531);
nand U9915 (N_9915,N_3452,N_3138);
nor U9916 (N_9916,N_1070,N_1348);
or U9917 (N_9917,N_4169,N_2429);
xnor U9918 (N_9918,N_1512,N_1015);
and U9919 (N_9919,N_5845,N_2227);
nor U9920 (N_9920,N_1440,N_5744);
xor U9921 (N_9921,N_2996,N_5289);
nand U9922 (N_9922,N_796,N_2759);
xnor U9923 (N_9923,N_2947,N_365);
or U9924 (N_9924,N_2457,N_3917);
and U9925 (N_9925,N_2549,N_2383);
xor U9926 (N_9926,N_2227,N_2552);
nand U9927 (N_9927,N_5509,N_2359);
nor U9928 (N_9928,N_5894,N_5955);
xor U9929 (N_9929,N_2216,N_1586);
or U9930 (N_9930,N_4126,N_5203);
xor U9931 (N_9931,N_5359,N_5797);
nor U9932 (N_9932,N_2676,N_4428);
or U9933 (N_9933,N_1513,N_3963);
nor U9934 (N_9934,N_5220,N_5707);
or U9935 (N_9935,N_1819,N_1716);
nor U9936 (N_9936,N_1873,N_1534);
or U9937 (N_9937,N_4669,N_1813);
or U9938 (N_9938,N_1213,N_3691);
nor U9939 (N_9939,N_1596,N_1819);
or U9940 (N_9940,N_4734,N_4996);
and U9941 (N_9941,N_3526,N_3744);
nor U9942 (N_9942,N_1142,N_4357);
xnor U9943 (N_9943,N_895,N_4250);
and U9944 (N_9944,N_5243,N_195);
nor U9945 (N_9945,N_5307,N_3170);
nand U9946 (N_9946,N_4610,N_4593);
nor U9947 (N_9947,N_4804,N_937);
nand U9948 (N_9948,N_1938,N_1520);
and U9949 (N_9949,N_5742,N_627);
and U9950 (N_9950,N_1335,N_4936);
xor U9951 (N_9951,N_4593,N_5074);
xor U9952 (N_9952,N_5918,N_2046);
or U9953 (N_9953,N_2980,N_3685);
and U9954 (N_9954,N_5318,N_1511);
or U9955 (N_9955,N_3236,N_3329);
or U9956 (N_9956,N_2386,N_4225);
nand U9957 (N_9957,N_5909,N_1729);
nand U9958 (N_9958,N_5993,N_717);
and U9959 (N_9959,N_3881,N_2200);
and U9960 (N_9960,N_4272,N_1069);
xor U9961 (N_9961,N_3958,N_1594);
or U9962 (N_9962,N_5507,N_1172);
xnor U9963 (N_9963,N_2067,N_5170);
xnor U9964 (N_9964,N_3891,N_378);
nor U9965 (N_9965,N_3606,N_138);
xor U9966 (N_9966,N_5803,N_4485);
xor U9967 (N_9967,N_4388,N_4694);
xnor U9968 (N_9968,N_3324,N_5766);
and U9969 (N_9969,N_1189,N_5082);
xnor U9970 (N_9970,N_3388,N_692);
or U9971 (N_9971,N_609,N_1594);
or U9972 (N_9972,N_4371,N_1770);
nand U9973 (N_9973,N_3737,N_2270);
nand U9974 (N_9974,N_4504,N_5569);
or U9975 (N_9975,N_4932,N_2352);
nor U9976 (N_9976,N_4663,N_1698);
or U9977 (N_9977,N_5567,N_2788);
nand U9978 (N_9978,N_244,N_5867);
nand U9979 (N_9979,N_2315,N_3968);
and U9980 (N_9980,N_1552,N_3579);
and U9981 (N_9981,N_1020,N_5916);
nor U9982 (N_9982,N_2243,N_3244);
xor U9983 (N_9983,N_4487,N_5437);
nor U9984 (N_9984,N_454,N_1576);
and U9985 (N_9985,N_4970,N_4586);
or U9986 (N_9986,N_3346,N_5392);
or U9987 (N_9987,N_344,N_5721);
xor U9988 (N_9988,N_1333,N_2948);
or U9989 (N_9989,N_4332,N_2526);
or U9990 (N_9990,N_1168,N_5574);
nor U9991 (N_9991,N_5566,N_606);
nand U9992 (N_9992,N_4171,N_2366);
nand U9993 (N_9993,N_4365,N_5473);
nor U9994 (N_9994,N_4172,N_268);
nand U9995 (N_9995,N_637,N_235);
and U9996 (N_9996,N_1470,N_2452);
nor U9997 (N_9997,N_5585,N_3972);
nand U9998 (N_9998,N_1385,N_1653);
nand U9999 (N_9999,N_5194,N_4372);
nor U10000 (N_10000,N_5540,N_4369);
or U10001 (N_10001,N_2504,N_5666);
or U10002 (N_10002,N_4893,N_1434);
nand U10003 (N_10003,N_2986,N_5177);
nor U10004 (N_10004,N_5932,N_2379);
nor U10005 (N_10005,N_5606,N_3814);
nor U10006 (N_10006,N_3523,N_5040);
nor U10007 (N_10007,N_5999,N_1020);
xnor U10008 (N_10008,N_5270,N_1877);
nor U10009 (N_10009,N_988,N_3040);
and U10010 (N_10010,N_2544,N_4252);
nand U10011 (N_10011,N_126,N_470);
xnor U10012 (N_10012,N_471,N_3401);
nor U10013 (N_10013,N_5135,N_4428);
or U10014 (N_10014,N_803,N_4912);
xor U10015 (N_10015,N_5061,N_2513);
nand U10016 (N_10016,N_696,N_2236);
nand U10017 (N_10017,N_2759,N_5772);
xor U10018 (N_10018,N_125,N_4662);
nor U10019 (N_10019,N_5603,N_2016);
and U10020 (N_10020,N_4421,N_275);
xor U10021 (N_10021,N_2281,N_721);
nand U10022 (N_10022,N_4416,N_5287);
or U10023 (N_10023,N_147,N_4533);
and U10024 (N_10024,N_3400,N_5084);
nor U10025 (N_10025,N_3503,N_685);
or U10026 (N_10026,N_91,N_5743);
xnor U10027 (N_10027,N_2448,N_2425);
xor U10028 (N_10028,N_305,N_3517);
nor U10029 (N_10029,N_2702,N_3122);
nand U10030 (N_10030,N_2797,N_769);
nor U10031 (N_10031,N_3162,N_1872);
nor U10032 (N_10032,N_3605,N_5489);
nand U10033 (N_10033,N_5482,N_2101);
and U10034 (N_10034,N_946,N_1591);
nor U10035 (N_10035,N_4408,N_27);
xor U10036 (N_10036,N_366,N_4086);
or U10037 (N_10037,N_713,N_3637);
nand U10038 (N_10038,N_1709,N_565);
or U10039 (N_10039,N_1173,N_1566);
nor U10040 (N_10040,N_2649,N_3389);
nor U10041 (N_10041,N_4533,N_3458);
xor U10042 (N_10042,N_919,N_5513);
or U10043 (N_10043,N_2255,N_3272);
and U10044 (N_10044,N_5249,N_5936);
or U10045 (N_10045,N_4244,N_948);
xor U10046 (N_10046,N_3121,N_3613);
xor U10047 (N_10047,N_4762,N_4356);
nor U10048 (N_10048,N_3883,N_5939);
and U10049 (N_10049,N_503,N_2225);
xor U10050 (N_10050,N_2883,N_2912);
xnor U10051 (N_10051,N_1664,N_866);
nor U10052 (N_10052,N_959,N_3833);
nor U10053 (N_10053,N_4348,N_5736);
and U10054 (N_10054,N_728,N_2934);
and U10055 (N_10055,N_3387,N_568);
xor U10056 (N_10056,N_3879,N_2262);
nor U10057 (N_10057,N_4870,N_67);
nand U10058 (N_10058,N_1081,N_2069);
nor U10059 (N_10059,N_1402,N_3334);
nand U10060 (N_10060,N_3745,N_4087);
nor U10061 (N_10061,N_3506,N_2553);
or U10062 (N_10062,N_5929,N_5381);
and U10063 (N_10063,N_1303,N_56);
or U10064 (N_10064,N_1071,N_2016);
and U10065 (N_10065,N_4630,N_2600);
nor U10066 (N_10066,N_2839,N_1457);
and U10067 (N_10067,N_4313,N_2221);
nor U10068 (N_10068,N_1840,N_3150);
nand U10069 (N_10069,N_5672,N_47);
or U10070 (N_10070,N_5325,N_4165);
nand U10071 (N_10071,N_4401,N_5650);
xor U10072 (N_10072,N_2350,N_5475);
nor U10073 (N_10073,N_3442,N_3175);
or U10074 (N_10074,N_5215,N_1058);
or U10075 (N_10075,N_4090,N_3886);
or U10076 (N_10076,N_3881,N_2179);
nand U10077 (N_10077,N_4600,N_4009);
nand U10078 (N_10078,N_1827,N_3362);
and U10079 (N_10079,N_49,N_5408);
nand U10080 (N_10080,N_4342,N_2814);
nor U10081 (N_10081,N_2260,N_5151);
and U10082 (N_10082,N_2041,N_1492);
xor U10083 (N_10083,N_3312,N_2141);
nand U10084 (N_10084,N_4783,N_3723);
nor U10085 (N_10085,N_5902,N_3200);
and U10086 (N_10086,N_415,N_5602);
and U10087 (N_10087,N_102,N_2433);
nor U10088 (N_10088,N_2783,N_3153);
xor U10089 (N_10089,N_3426,N_2622);
nor U10090 (N_10090,N_3458,N_1717);
xor U10091 (N_10091,N_3375,N_2283);
xor U10092 (N_10092,N_3164,N_5336);
and U10093 (N_10093,N_850,N_4137);
xnor U10094 (N_10094,N_2723,N_2884);
or U10095 (N_10095,N_4450,N_4668);
and U10096 (N_10096,N_5985,N_5130);
xnor U10097 (N_10097,N_1006,N_1595);
xnor U10098 (N_10098,N_643,N_3704);
nor U10099 (N_10099,N_3791,N_4212);
nand U10100 (N_10100,N_103,N_4920);
xnor U10101 (N_10101,N_296,N_1276);
and U10102 (N_10102,N_4109,N_3536);
or U10103 (N_10103,N_3765,N_3134);
xnor U10104 (N_10104,N_3550,N_4831);
nor U10105 (N_10105,N_4675,N_1631);
and U10106 (N_10106,N_4533,N_42);
xor U10107 (N_10107,N_5164,N_568);
and U10108 (N_10108,N_1912,N_1519);
nand U10109 (N_10109,N_1568,N_3215);
or U10110 (N_10110,N_2139,N_5738);
xor U10111 (N_10111,N_2659,N_3628);
or U10112 (N_10112,N_117,N_3475);
nor U10113 (N_10113,N_2989,N_4977);
nor U10114 (N_10114,N_2014,N_4123);
xnor U10115 (N_10115,N_3860,N_4902);
or U10116 (N_10116,N_97,N_681);
xor U10117 (N_10117,N_3588,N_4543);
nand U10118 (N_10118,N_946,N_4844);
or U10119 (N_10119,N_2584,N_1528);
and U10120 (N_10120,N_1673,N_3186);
or U10121 (N_10121,N_5744,N_2469);
nor U10122 (N_10122,N_1034,N_1926);
nand U10123 (N_10123,N_1517,N_2670);
nand U10124 (N_10124,N_1331,N_4082);
and U10125 (N_10125,N_5989,N_1294);
and U10126 (N_10126,N_3933,N_5900);
nand U10127 (N_10127,N_3027,N_4486);
nor U10128 (N_10128,N_1139,N_3480);
or U10129 (N_10129,N_1820,N_2604);
xor U10130 (N_10130,N_5830,N_2842);
or U10131 (N_10131,N_2493,N_1320);
xor U10132 (N_10132,N_3507,N_1231);
xnor U10133 (N_10133,N_1545,N_8);
nand U10134 (N_10134,N_839,N_3465);
or U10135 (N_10135,N_3321,N_429);
or U10136 (N_10136,N_4086,N_2184);
nand U10137 (N_10137,N_310,N_4746);
and U10138 (N_10138,N_4772,N_3128);
nand U10139 (N_10139,N_182,N_3316);
nand U10140 (N_10140,N_2061,N_3446);
nor U10141 (N_10141,N_3575,N_212);
and U10142 (N_10142,N_713,N_5311);
and U10143 (N_10143,N_3645,N_470);
nand U10144 (N_10144,N_5191,N_5465);
nand U10145 (N_10145,N_4599,N_5263);
xnor U10146 (N_10146,N_1851,N_1294);
xor U10147 (N_10147,N_1723,N_4576);
xnor U10148 (N_10148,N_4741,N_5262);
or U10149 (N_10149,N_2976,N_1307);
or U10150 (N_10150,N_1558,N_4493);
xnor U10151 (N_10151,N_5709,N_2841);
and U10152 (N_10152,N_2076,N_42);
nor U10153 (N_10153,N_1897,N_496);
nor U10154 (N_10154,N_3033,N_2242);
nor U10155 (N_10155,N_2607,N_2523);
or U10156 (N_10156,N_412,N_774);
and U10157 (N_10157,N_5652,N_1978);
nor U10158 (N_10158,N_2288,N_573);
xnor U10159 (N_10159,N_5489,N_5491);
xor U10160 (N_10160,N_1063,N_493);
nor U10161 (N_10161,N_3839,N_2677);
or U10162 (N_10162,N_650,N_3756);
nor U10163 (N_10163,N_2804,N_2698);
and U10164 (N_10164,N_64,N_4535);
and U10165 (N_10165,N_3774,N_5699);
or U10166 (N_10166,N_658,N_3945);
and U10167 (N_10167,N_1582,N_362);
xnor U10168 (N_10168,N_1246,N_582);
or U10169 (N_10169,N_2333,N_2802);
nand U10170 (N_10170,N_99,N_1414);
and U10171 (N_10171,N_5479,N_2216);
nor U10172 (N_10172,N_198,N_5246);
or U10173 (N_10173,N_5332,N_4436);
nor U10174 (N_10174,N_194,N_5910);
nand U10175 (N_10175,N_5968,N_2743);
and U10176 (N_10176,N_1456,N_438);
xor U10177 (N_10177,N_3359,N_1828);
nand U10178 (N_10178,N_1303,N_203);
or U10179 (N_10179,N_3600,N_3544);
xor U10180 (N_10180,N_3721,N_2475);
or U10181 (N_10181,N_19,N_5071);
and U10182 (N_10182,N_3539,N_3181);
xor U10183 (N_10183,N_4596,N_1992);
nand U10184 (N_10184,N_168,N_397);
nand U10185 (N_10185,N_5531,N_1478);
xor U10186 (N_10186,N_1899,N_5864);
nor U10187 (N_10187,N_1729,N_2764);
or U10188 (N_10188,N_5884,N_941);
xor U10189 (N_10189,N_5339,N_1008);
nor U10190 (N_10190,N_4566,N_1918);
nand U10191 (N_10191,N_34,N_4288);
or U10192 (N_10192,N_4952,N_2108);
and U10193 (N_10193,N_3601,N_864);
and U10194 (N_10194,N_1101,N_480);
nor U10195 (N_10195,N_3898,N_330);
nand U10196 (N_10196,N_3115,N_1011);
or U10197 (N_10197,N_3541,N_4496);
nand U10198 (N_10198,N_2723,N_339);
xor U10199 (N_10199,N_2269,N_3880);
or U10200 (N_10200,N_3385,N_4040);
or U10201 (N_10201,N_1104,N_3916);
and U10202 (N_10202,N_3852,N_728);
and U10203 (N_10203,N_3182,N_4488);
xnor U10204 (N_10204,N_4931,N_4156);
xnor U10205 (N_10205,N_968,N_5243);
nand U10206 (N_10206,N_1140,N_3486);
and U10207 (N_10207,N_2744,N_3059);
xnor U10208 (N_10208,N_3206,N_3360);
or U10209 (N_10209,N_5557,N_3424);
nand U10210 (N_10210,N_642,N_4843);
nand U10211 (N_10211,N_1115,N_19);
and U10212 (N_10212,N_5576,N_5653);
nand U10213 (N_10213,N_2418,N_5002);
nor U10214 (N_10214,N_277,N_2105);
and U10215 (N_10215,N_2371,N_1527);
or U10216 (N_10216,N_2371,N_3454);
nor U10217 (N_10217,N_3666,N_2368);
nand U10218 (N_10218,N_4710,N_3866);
nand U10219 (N_10219,N_4146,N_93);
nor U10220 (N_10220,N_399,N_2808);
xor U10221 (N_10221,N_1419,N_5253);
or U10222 (N_10222,N_573,N_5484);
xnor U10223 (N_10223,N_3503,N_4124);
nor U10224 (N_10224,N_2015,N_5667);
or U10225 (N_10225,N_4811,N_2390);
or U10226 (N_10226,N_4267,N_3168);
nor U10227 (N_10227,N_5205,N_2178);
nand U10228 (N_10228,N_1838,N_587);
nor U10229 (N_10229,N_3975,N_3147);
xnor U10230 (N_10230,N_3188,N_1462);
xor U10231 (N_10231,N_3227,N_4114);
nand U10232 (N_10232,N_2604,N_5501);
nor U10233 (N_10233,N_1954,N_663);
nand U10234 (N_10234,N_206,N_5426);
xnor U10235 (N_10235,N_3587,N_2928);
nand U10236 (N_10236,N_748,N_2293);
nor U10237 (N_10237,N_5066,N_1181);
or U10238 (N_10238,N_2070,N_522);
nand U10239 (N_10239,N_3333,N_3643);
nand U10240 (N_10240,N_3668,N_5149);
nand U10241 (N_10241,N_5398,N_3329);
and U10242 (N_10242,N_1082,N_2483);
nand U10243 (N_10243,N_1096,N_5829);
and U10244 (N_10244,N_221,N_5313);
and U10245 (N_10245,N_671,N_4644);
or U10246 (N_10246,N_4750,N_4888);
nand U10247 (N_10247,N_1901,N_1969);
nand U10248 (N_10248,N_3938,N_5462);
and U10249 (N_10249,N_2261,N_4638);
xor U10250 (N_10250,N_5606,N_3656);
nand U10251 (N_10251,N_5153,N_5775);
or U10252 (N_10252,N_3563,N_5240);
nor U10253 (N_10253,N_1228,N_914);
and U10254 (N_10254,N_2851,N_4144);
nand U10255 (N_10255,N_2938,N_2731);
nor U10256 (N_10256,N_5254,N_5947);
xor U10257 (N_10257,N_5416,N_50);
nand U10258 (N_10258,N_3594,N_5139);
or U10259 (N_10259,N_4652,N_4549);
and U10260 (N_10260,N_2648,N_4978);
or U10261 (N_10261,N_4812,N_4658);
xnor U10262 (N_10262,N_3646,N_1393);
or U10263 (N_10263,N_3660,N_2921);
nor U10264 (N_10264,N_3144,N_2805);
or U10265 (N_10265,N_5723,N_4401);
and U10266 (N_10266,N_973,N_2575);
nand U10267 (N_10267,N_1520,N_1624);
nor U10268 (N_10268,N_873,N_687);
nand U10269 (N_10269,N_1662,N_4881);
nor U10270 (N_10270,N_5999,N_3932);
nor U10271 (N_10271,N_1506,N_2244);
and U10272 (N_10272,N_961,N_4711);
xor U10273 (N_10273,N_3186,N_3532);
and U10274 (N_10274,N_2900,N_4003);
xor U10275 (N_10275,N_3787,N_2614);
xnor U10276 (N_10276,N_1871,N_2170);
or U10277 (N_10277,N_3696,N_2467);
xnor U10278 (N_10278,N_3409,N_1542);
nand U10279 (N_10279,N_3149,N_3634);
nand U10280 (N_10280,N_3752,N_3519);
nor U10281 (N_10281,N_5954,N_2576);
nand U10282 (N_10282,N_5672,N_5155);
nand U10283 (N_10283,N_2513,N_2759);
xor U10284 (N_10284,N_578,N_3695);
and U10285 (N_10285,N_1383,N_1656);
xor U10286 (N_10286,N_3712,N_619);
nand U10287 (N_10287,N_2598,N_2145);
and U10288 (N_10288,N_5843,N_0);
nor U10289 (N_10289,N_3353,N_5552);
and U10290 (N_10290,N_2964,N_453);
and U10291 (N_10291,N_3852,N_3947);
nor U10292 (N_10292,N_656,N_430);
or U10293 (N_10293,N_1286,N_2080);
and U10294 (N_10294,N_3755,N_3625);
nand U10295 (N_10295,N_3537,N_5758);
or U10296 (N_10296,N_2510,N_120);
nand U10297 (N_10297,N_629,N_1159);
nand U10298 (N_10298,N_1809,N_1656);
nor U10299 (N_10299,N_5104,N_826);
nand U10300 (N_10300,N_1557,N_5303);
nor U10301 (N_10301,N_3294,N_438);
and U10302 (N_10302,N_2504,N_4792);
and U10303 (N_10303,N_5183,N_5154);
nor U10304 (N_10304,N_4748,N_1586);
and U10305 (N_10305,N_3330,N_5461);
xor U10306 (N_10306,N_5282,N_3444);
xnor U10307 (N_10307,N_2127,N_2632);
or U10308 (N_10308,N_5739,N_408);
nor U10309 (N_10309,N_2608,N_3404);
xnor U10310 (N_10310,N_3896,N_3145);
xnor U10311 (N_10311,N_349,N_3512);
xor U10312 (N_10312,N_3253,N_1787);
nand U10313 (N_10313,N_4079,N_1212);
nor U10314 (N_10314,N_2087,N_5444);
nand U10315 (N_10315,N_1162,N_5439);
or U10316 (N_10316,N_4392,N_3418);
xor U10317 (N_10317,N_2501,N_2991);
nand U10318 (N_10318,N_4909,N_3706);
nand U10319 (N_10319,N_1147,N_3376);
and U10320 (N_10320,N_942,N_3356);
or U10321 (N_10321,N_2371,N_3944);
and U10322 (N_10322,N_4494,N_3629);
and U10323 (N_10323,N_1029,N_3166);
and U10324 (N_10324,N_5366,N_3797);
and U10325 (N_10325,N_3294,N_5663);
and U10326 (N_10326,N_1808,N_5156);
and U10327 (N_10327,N_3033,N_5156);
xor U10328 (N_10328,N_1437,N_2352);
nor U10329 (N_10329,N_5441,N_2552);
and U10330 (N_10330,N_1071,N_2408);
nand U10331 (N_10331,N_2493,N_1196);
and U10332 (N_10332,N_349,N_944);
and U10333 (N_10333,N_2653,N_310);
nand U10334 (N_10334,N_1873,N_1822);
xnor U10335 (N_10335,N_2282,N_1016);
nand U10336 (N_10336,N_829,N_5354);
nor U10337 (N_10337,N_4807,N_3601);
xor U10338 (N_10338,N_5063,N_4338);
or U10339 (N_10339,N_96,N_2851);
xor U10340 (N_10340,N_3799,N_28);
and U10341 (N_10341,N_1975,N_5148);
nand U10342 (N_10342,N_1914,N_5378);
xor U10343 (N_10343,N_5166,N_819);
nand U10344 (N_10344,N_4615,N_4795);
nor U10345 (N_10345,N_4610,N_4769);
or U10346 (N_10346,N_2285,N_4165);
or U10347 (N_10347,N_3429,N_1011);
xor U10348 (N_10348,N_4138,N_4913);
and U10349 (N_10349,N_4951,N_4574);
or U10350 (N_10350,N_5472,N_2557);
xor U10351 (N_10351,N_911,N_2156);
and U10352 (N_10352,N_797,N_3481);
nor U10353 (N_10353,N_2701,N_5710);
xnor U10354 (N_10354,N_1300,N_3477);
nor U10355 (N_10355,N_983,N_197);
or U10356 (N_10356,N_3086,N_307);
or U10357 (N_10357,N_3292,N_2497);
or U10358 (N_10358,N_4659,N_2413);
and U10359 (N_10359,N_5776,N_3401);
xor U10360 (N_10360,N_932,N_5239);
or U10361 (N_10361,N_2243,N_3792);
and U10362 (N_10362,N_3549,N_3470);
nor U10363 (N_10363,N_136,N_5505);
nor U10364 (N_10364,N_3521,N_1850);
nand U10365 (N_10365,N_2314,N_4761);
and U10366 (N_10366,N_2482,N_4187);
nor U10367 (N_10367,N_5271,N_3559);
and U10368 (N_10368,N_1626,N_5363);
nor U10369 (N_10369,N_5326,N_2840);
nand U10370 (N_10370,N_436,N_2916);
or U10371 (N_10371,N_3309,N_1750);
nand U10372 (N_10372,N_1718,N_4704);
or U10373 (N_10373,N_4982,N_3490);
xnor U10374 (N_10374,N_2676,N_5469);
nor U10375 (N_10375,N_4222,N_5372);
and U10376 (N_10376,N_1374,N_2947);
nand U10377 (N_10377,N_2545,N_2005);
and U10378 (N_10378,N_2346,N_1898);
and U10379 (N_10379,N_3848,N_4703);
or U10380 (N_10380,N_55,N_1801);
nor U10381 (N_10381,N_3496,N_3034);
and U10382 (N_10382,N_3898,N_900);
nand U10383 (N_10383,N_3741,N_1870);
nor U10384 (N_10384,N_2965,N_1222);
nand U10385 (N_10385,N_5288,N_2409);
xor U10386 (N_10386,N_4257,N_3966);
nor U10387 (N_10387,N_894,N_2184);
and U10388 (N_10388,N_3784,N_4831);
xnor U10389 (N_10389,N_4249,N_3091);
or U10390 (N_10390,N_4245,N_1109);
or U10391 (N_10391,N_5471,N_3272);
nor U10392 (N_10392,N_5256,N_5257);
nand U10393 (N_10393,N_5179,N_4657);
nor U10394 (N_10394,N_2579,N_1544);
xnor U10395 (N_10395,N_2667,N_204);
and U10396 (N_10396,N_5667,N_3904);
and U10397 (N_10397,N_1784,N_1033);
and U10398 (N_10398,N_3914,N_367);
and U10399 (N_10399,N_2296,N_3374);
xnor U10400 (N_10400,N_4529,N_4673);
nand U10401 (N_10401,N_620,N_5954);
nor U10402 (N_10402,N_5719,N_5821);
or U10403 (N_10403,N_821,N_2870);
nor U10404 (N_10404,N_5116,N_494);
nor U10405 (N_10405,N_3858,N_1989);
and U10406 (N_10406,N_1627,N_3810);
nor U10407 (N_10407,N_2921,N_3655);
nor U10408 (N_10408,N_4265,N_5301);
and U10409 (N_10409,N_1559,N_1801);
or U10410 (N_10410,N_1722,N_4000);
and U10411 (N_10411,N_1804,N_945);
xnor U10412 (N_10412,N_4048,N_3721);
nand U10413 (N_10413,N_1865,N_2034);
and U10414 (N_10414,N_3112,N_583);
nor U10415 (N_10415,N_5139,N_2415);
xnor U10416 (N_10416,N_257,N_4394);
nor U10417 (N_10417,N_2358,N_469);
nand U10418 (N_10418,N_1832,N_689);
nand U10419 (N_10419,N_3459,N_2560);
or U10420 (N_10420,N_1150,N_5278);
or U10421 (N_10421,N_650,N_1063);
or U10422 (N_10422,N_2936,N_198);
or U10423 (N_10423,N_2392,N_479);
and U10424 (N_10424,N_3160,N_4317);
xor U10425 (N_10425,N_5909,N_4730);
or U10426 (N_10426,N_1717,N_3173);
xor U10427 (N_10427,N_547,N_5037);
or U10428 (N_10428,N_5808,N_3328);
xnor U10429 (N_10429,N_2995,N_490);
and U10430 (N_10430,N_1740,N_3747);
nand U10431 (N_10431,N_2091,N_3104);
nor U10432 (N_10432,N_3676,N_4149);
and U10433 (N_10433,N_2678,N_2061);
xnor U10434 (N_10434,N_5702,N_4899);
nor U10435 (N_10435,N_59,N_931);
or U10436 (N_10436,N_4057,N_3123);
and U10437 (N_10437,N_174,N_1922);
or U10438 (N_10438,N_2163,N_5435);
nor U10439 (N_10439,N_2830,N_2036);
nand U10440 (N_10440,N_2304,N_4073);
and U10441 (N_10441,N_4328,N_118);
xnor U10442 (N_10442,N_289,N_3318);
or U10443 (N_10443,N_3882,N_2435);
xnor U10444 (N_10444,N_3389,N_5407);
nor U10445 (N_10445,N_4308,N_5867);
and U10446 (N_10446,N_1915,N_3961);
xor U10447 (N_10447,N_5357,N_5943);
or U10448 (N_10448,N_415,N_5698);
or U10449 (N_10449,N_2855,N_932);
and U10450 (N_10450,N_568,N_254);
xnor U10451 (N_10451,N_3689,N_4856);
or U10452 (N_10452,N_3513,N_1779);
or U10453 (N_10453,N_4009,N_2113);
or U10454 (N_10454,N_5297,N_5619);
nand U10455 (N_10455,N_3107,N_5101);
and U10456 (N_10456,N_4881,N_4455);
and U10457 (N_10457,N_5893,N_4123);
nand U10458 (N_10458,N_4475,N_4433);
and U10459 (N_10459,N_3012,N_3809);
nor U10460 (N_10460,N_1461,N_1981);
xor U10461 (N_10461,N_1558,N_761);
xnor U10462 (N_10462,N_2517,N_5241);
xnor U10463 (N_10463,N_2795,N_196);
and U10464 (N_10464,N_606,N_2594);
nor U10465 (N_10465,N_4805,N_2881);
nor U10466 (N_10466,N_1892,N_468);
or U10467 (N_10467,N_5989,N_2216);
or U10468 (N_10468,N_4645,N_4962);
nand U10469 (N_10469,N_3428,N_4124);
xor U10470 (N_10470,N_965,N_1603);
or U10471 (N_10471,N_168,N_2973);
nor U10472 (N_10472,N_949,N_3573);
or U10473 (N_10473,N_2401,N_3582);
nor U10474 (N_10474,N_4183,N_3987);
xnor U10475 (N_10475,N_5535,N_827);
or U10476 (N_10476,N_1286,N_3236);
xnor U10477 (N_10477,N_1923,N_5810);
xor U10478 (N_10478,N_426,N_2382);
xnor U10479 (N_10479,N_4415,N_4219);
nor U10480 (N_10480,N_1167,N_671);
xnor U10481 (N_10481,N_5555,N_5597);
xnor U10482 (N_10482,N_3046,N_1808);
nor U10483 (N_10483,N_1521,N_2455);
xor U10484 (N_10484,N_1164,N_3415);
nand U10485 (N_10485,N_113,N_5243);
and U10486 (N_10486,N_5139,N_2663);
or U10487 (N_10487,N_409,N_1278);
or U10488 (N_10488,N_5241,N_1885);
nand U10489 (N_10489,N_1848,N_4492);
and U10490 (N_10490,N_333,N_1146);
xor U10491 (N_10491,N_5386,N_2110);
nor U10492 (N_10492,N_575,N_736);
nand U10493 (N_10493,N_802,N_5116);
nor U10494 (N_10494,N_748,N_2674);
xnor U10495 (N_10495,N_4959,N_1203);
or U10496 (N_10496,N_5477,N_1323);
or U10497 (N_10497,N_3404,N_2273);
nor U10498 (N_10498,N_1174,N_4150);
or U10499 (N_10499,N_5417,N_3249);
xnor U10500 (N_10500,N_66,N_2720);
and U10501 (N_10501,N_4951,N_5650);
or U10502 (N_10502,N_2712,N_5316);
nand U10503 (N_10503,N_2630,N_3924);
or U10504 (N_10504,N_5518,N_5885);
nor U10505 (N_10505,N_3748,N_813);
nand U10506 (N_10506,N_3535,N_2462);
nand U10507 (N_10507,N_4808,N_5455);
nor U10508 (N_10508,N_1360,N_1485);
and U10509 (N_10509,N_2892,N_5156);
or U10510 (N_10510,N_2482,N_4245);
nor U10511 (N_10511,N_3459,N_2979);
xor U10512 (N_10512,N_4500,N_1736);
xor U10513 (N_10513,N_657,N_1752);
xnor U10514 (N_10514,N_2792,N_5129);
nor U10515 (N_10515,N_1746,N_922);
nand U10516 (N_10516,N_1194,N_4941);
nor U10517 (N_10517,N_3836,N_3842);
nor U10518 (N_10518,N_1316,N_1551);
and U10519 (N_10519,N_3074,N_4140);
xnor U10520 (N_10520,N_5919,N_5769);
nor U10521 (N_10521,N_407,N_929);
or U10522 (N_10522,N_3273,N_3633);
and U10523 (N_10523,N_567,N_1537);
or U10524 (N_10524,N_5825,N_206);
or U10525 (N_10525,N_4561,N_927);
and U10526 (N_10526,N_5319,N_1235);
or U10527 (N_10527,N_5103,N_4959);
xnor U10528 (N_10528,N_5281,N_5136);
and U10529 (N_10529,N_2053,N_3446);
nand U10530 (N_10530,N_4960,N_3574);
and U10531 (N_10531,N_5253,N_4833);
and U10532 (N_10532,N_1064,N_2065);
or U10533 (N_10533,N_1313,N_4717);
or U10534 (N_10534,N_5657,N_764);
xor U10535 (N_10535,N_2106,N_2349);
nor U10536 (N_10536,N_3168,N_517);
nor U10537 (N_10537,N_2187,N_2746);
xor U10538 (N_10538,N_5843,N_5113);
nand U10539 (N_10539,N_2341,N_3146);
nand U10540 (N_10540,N_1379,N_5951);
or U10541 (N_10541,N_1928,N_2930);
and U10542 (N_10542,N_2376,N_4730);
nand U10543 (N_10543,N_5299,N_5698);
nand U10544 (N_10544,N_4998,N_1475);
nor U10545 (N_10545,N_3175,N_206);
xor U10546 (N_10546,N_5647,N_2576);
or U10547 (N_10547,N_307,N_496);
nor U10548 (N_10548,N_834,N_5347);
nand U10549 (N_10549,N_1267,N_2877);
nor U10550 (N_10550,N_5559,N_3010);
nor U10551 (N_10551,N_3469,N_34);
or U10552 (N_10552,N_5634,N_4942);
and U10553 (N_10553,N_2658,N_669);
xor U10554 (N_10554,N_4815,N_4682);
or U10555 (N_10555,N_3407,N_254);
xnor U10556 (N_10556,N_252,N_2911);
nor U10557 (N_10557,N_1898,N_2811);
nand U10558 (N_10558,N_3757,N_913);
nor U10559 (N_10559,N_794,N_508);
nand U10560 (N_10560,N_2501,N_4981);
nor U10561 (N_10561,N_5181,N_4163);
xnor U10562 (N_10562,N_548,N_4069);
xnor U10563 (N_10563,N_2464,N_1764);
xnor U10564 (N_10564,N_3487,N_3585);
xnor U10565 (N_10565,N_5918,N_910);
and U10566 (N_10566,N_5339,N_5022);
nand U10567 (N_10567,N_5314,N_2622);
and U10568 (N_10568,N_1747,N_3442);
or U10569 (N_10569,N_1485,N_2572);
nor U10570 (N_10570,N_853,N_3106);
nor U10571 (N_10571,N_2699,N_189);
xor U10572 (N_10572,N_4920,N_1539);
nor U10573 (N_10573,N_1307,N_888);
nand U10574 (N_10574,N_5021,N_4487);
or U10575 (N_10575,N_1139,N_5540);
xor U10576 (N_10576,N_3492,N_3342);
or U10577 (N_10577,N_2672,N_5655);
and U10578 (N_10578,N_3148,N_3739);
or U10579 (N_10579,N_4373,N_3523);
nand U10580 (N_10580,N_3636,N_5939);
and U10581 (N_10581,N_4654,N_3103);
and U10582 (N_10582,N_3700,N_4251);
and U10583 (N_10583,N_44,N_1129);
xnor U10584 (N_10584,N_1730,N_5802);
and U10585 (N_10585,N_3396,N_1547);
or U10586 (N_10586,N_3799,N_556);
or U10587 (N_10587,N_622,N_3062);
and U10588 (N_10588,N_5035,N_890);
and U10589 (N_10589,N_1479,N_5842);
xnor U10590 (N_10590,N_2022,N_5850);
nand U10591 (N_10591,N_3726,N_1047);
or U10592 (N_10592,N_2423,N_1394);
and U10593 (N_10593,N_1936,N_5264);
xnor U10594 (N_10594,N_5622,N_129);
xor U10595 (N_10595,N_5945,N_2173);
and U10596 (N_10596,N_1639,N_5153);
nor U10597 (N_10597,N_5146,N_2406);
xor U10598 (N_10598,N_3482,N_21);
xor U10599 (N_10599,N_1987,N_2105);
and U10600 (N_10600,N_1257,N_437);
nand U10601 (N_10601,N_4933,N_1053);
nor U10602 (N_10602,N_3056,N_1173);
or U10603 (N_10603,N_2363,N_1992);
xnor U10604 (N_10604,N_4004,N_4980);
nor U10605 (N_10605,N_5907,N_941);
and U10606 (N_10606,N_3266,N_3636);
xnor U10607 (N_10607,N_4024,N_1337);
and U10608 (N_10608,N_5681,N_1531);
and U10609 (N_10609,N_3705,N_4021);
or U10610 (N_10610,N_3968,N_178);
or U10611 (N_10611,N_5820,N_3049);
nand U10612 (N_10612,N_5891,N_4550);
nor U10613 (N_10613,N_5703,N_3413);
or U10614 (N_10614,N_5907,N_4935);
or U10615 (N_10615,N_5348,N_824);
nand U10616 (N_10616,N_2116,N_2112);
and U10617 (N_10617,N_4008,N_3869);
or U10618 (N_10618,N_3021,N_4728);
or U10619 (N_10619,N_5610,N_2176);
nand U10620 (N_10620,N_2860,N_4094);
nand U10621 (N_10621,N_2550,N_5072);
and U10622 (N_10622,N_4220,N_2552);
or U10623 (N_10623,N_3967,N_2877);
and U10624 (N_10624,N_2265,N_5045);
or U10625 (N_10625,N_2700,N_1830);
or U10626 (N_10626,N_5345,N_914);
or U10627 (N_10627,N_3213,N_2041);
and U10628 (N_10628,N_5634,N_5692);
xnor U10629 (N_10629,N_4964,N_2774);
xor U10630 (N_10630,N_2656,N_5578);
nor U10631 (N_10631,N_3741,N_5707);
nor U10632 (N_10632,N_2813,N_2704);
nor U10633 (N_10633,N_3293,N_4472);
nand U10634 (N_10634,N_3756,N_3898);
xnor U10635 (N_10635,N_4972,N_4306);
xnor U10636 (N_10636,N_345,N_1376);
or U10637 (N_10637,N_4240,N_3547);
or U10638 (N_10638,N_2626,N_1760);
and U10639 (N_10639,N_1739,N_945);
nand U10640 (N_10640,N_4748,N_1483);
nor U10641 (N_10641,N_123,N_99);
xor U10642 (N_10642,N_3376,N_3859);
xnor U10643 (N_10643,N_2983,N_3799);
nand U10644 (N_10644,N_4980,N_5974);
or U10645 (N_10645,N_1547,N_1097);
xor U10646 (N_10646,N_2347,N_3218);
or U10647 (N_10647,N_3088,N_1912);
or U10648 (N_10648,N_681,N_1008);
nor U10649 (N_10649,N_4123,N_5863);
nand U10650 (N_10650,N_4876,N_1709);
nand U10651 (N_10651,N_2787,N_3264);
or U10652 (N_10652,N_1632,N_5899);
or U10653 (N_10653,N_3755,N_2443);
nand U10654 (N_10654,N_4947,N_887);
nand U10655 (N_10655,N_3044,N_5652);
nand U10656 (N_10656,N_640,N_4999);
nand U10657 (N_10657,N_2807,N_2131);
or U10658 (N_10658,N_3863,N_566);
and U10659 (N_10659,N_737,N_3584);
nand U10660 (N_10660,N_5734,N_1228);
and U10661 (N_10661,N_5789,N_3241);
nor U10662 (N_10662,N_5313,N_502);
xnor U10663 (N_10663,N_3984,N_5784);
and U10664 (N_10664,N_3929,N_4782);
and U10665 (N_10665,N_2329,N_4860);
and U10666 (N_10666,N_5364,N_1014);
and U10667 (N_10667,N_318,N_1859);
xnor U10668 (N_10668,N_3185,N_5253);
xor U10669 (N_10669,N_3099,N_3502);
or U10670 (N_10670,N_2261,N_3279);
nand U10671 (N_10671,N_3139,N_531);
xor U10672 (N_10672,N_2544,N_2075);
nand U10673 (N_10673,N_2402,N_4495);
or U10674 (N_10674,N_1736,N_2887);
nor U10675 (N_10675,N_562,N_1057);
nand U10676 (N_10676,N_2486,N_2556);
or U10677 (N_10677,N_5074,N_3930);
nand U10678 (N_10678,N_4962,N_5576);
or U10679 (N_10679,N_4655,N_3277);
xor U10680 (N_10680,N_4525,N_3295);
nor U10681 (N_10681,N_4004,N_169);
and U10682 (N_10682,N_840,N_2975);
and U10683 (N_10683,N_4372,N_5832);
or U10684 (N_10684,N_4768,N_2303);
xor U10685 (N_10685,N_632,N_4175);
or U10686 (N_10686,N_4061,N_5773);
or U10687 (N_10687,N_2023,N_2213);
or U10688 (N_10688,N_4557,N_8);
nand U10689 (N_10689,N_4746,N_1345);
nor U10690 (N_10690,N_4223,N_5475);
nand U10691 (N_10691,N_119,N_5080);
nor U10692 (N_10692,N_1906,N_5251);
or U10693 (N_10693,N_5935,N_4990);
nand U10694 (N_10694,N_2125,N_2611);
nand U10695 (N_10695,N_762,N_3808);
nor U10696 (N_10696,N_4474,N_4302);
nand U10697 (N_10697,N_5362,N_3090);
nor U10698 (N_10698,N_1092,N_5044);
nand U10699 (N_10699,N_5144,N_3927);
and U10700 (N_10700,N_167,N_2400);
nand U10701 (N_10701,N_3120,N_856);
and U10702 (N_10702,N_861,N_704);
xor U10703 (N_10703,N_778,N_4114);
nand U10704 (N_10704,N_1805,N_870);
or U10705 (N_10705,N_3144,N_1663);
and U10706 (N_10706,N_1214,N_820);
nor U10707 (N_10707,N_3662,N_126);
and U10708 (N_10708,N_1066,N_2148);
nor U10709 (N_10709,N_4360,N_4236);
nor U10710 (N_10710,N_4590,N_3598);
xor U10711 (N_10711,N_1138,N_2345);
or U10712 (N_10712,N_3475,N_948);
xnor U10713 (N_10713,N_5410,N_4883);
nor U10714 (N_10714,N_5246,N_1886);
xor U10715 (N_10715,N_505,N_2893);
xor U10716 (N_10716,N_2015,N_3950);
and U10717 (N_10717,N_103,N_1795);
nand U10718 (N_10718,N_3217,N_5426);
nor U10719 (N_10719,N_1078,N_557);
or U10720 (N_10720,N_2890,N_74);
or U10721 (N_10721,N_5777,N_2352);
and U10722 (N_10722,N_1343,N_5138);
nor U10723 (N_10723,N_4203,N_878);
or U10724 (N_10724,N_1928,N_2302);
and U10725 (N_10725,N_5953,N_4766);
and U10726 (N_10726,N_4001,N_3976);
xor U10727 (N_10727,N_4145,N_28);
and U10728 (N_10728,N_2748,N_86);
nand U10729 (N_10729,N_3934,N_4513);
and U10730 (N_10730,N_3883,N_3566);
xnor U10731 (N_10731,N_2498,N_5089);
nor U10732 (N_10732,N_5123,N_5975);
and U10733 (N_10733,N_2800,N_3108);
nand U10734 (N_10734,N_708,N_492);
nor U10735 (N_10735,N_5872,N_2791);
or U10736 (N_10736,N_1255,N_2922);
nor U10737 (N_10737,N_1425,N_1149);
and U10738 (N_10738,N_5094,N_5068);
xnor U10739 (N_10739,N_567,N_3861);
nand U10740 (N_10740,N_3832,N_1755);
nand U10741 (N_10741,N_4616,N_5870);
xor U10742 (N_10742,N_3161,N_821);
or U10743 (N_10743,N_2233,N_5851);
and U10744 (N_10744,N_2114,N_1530);
or U10745 (N_10745,N_4734,N_1458);
nor U10746 (N_10746,N_4755,N_2790);
xnor U10747 (N_10747,N_1212,N_1444);
xnor U10748 (N_10748,N_5969,N_123);
nor U10749 (N_10749,N_5843,N_3714);
xor U10750 (N_10750,N_464,N_1040);
nor U10751 (N_10751,N_4289,N_5166);
xnor U10752 (N_10752,N_1085,N_956);
nor U10753 (N_10753,N_3864,N_666);
nor U10754 (N_10754,N_5980,N_5712);
and U10755 (N_10755,N_445,N_2271);
nand U10756 (N_10756,N_3796,N_756);
nand U10757 (N_10757,N_4855,N_5534);
nor U10758 (N_10758,N_1024,N_3508);
nand U10759 (N_10759,N_5751,N_454);
nand U10760 (N_10760,N_5898,N_2380);
and U10761 (N_10761,N_3372,N_3333);
nor U10762 (N_10762,N_1602,N_3598);
and U10763 (N_10763,N_5198,N_5254);
and U10764 (N_10764,N_1350,N_5196);
or U10765 (N_10765,N_5720,N_90);
and U10766 (N_10766,N_2968,N_3627);
nor U10767 (N_10767,N_882,N_1947);
xor U10768 (N_10768,N_1864,N_3776);
and U10769 (N_10769,N_4444,N_3291);
xnor U10770 (N_10770,N_4266,N_2320);
xor U10771 (N_10771,N_318,N_4193);
nand U10772 (N_10772,N_4912,N_3553);
or U10773 (N_10773,N_3313,N_184);
nand U10774 (N_10774,N_4951,N_1381);
nor U10775 (N_10775,N_5531,N_3967);
xor U10776 (N_10776,N_3987,N_3400);
xnor U10777 (N_10777,N_1713,N_1199);
xor U10778 (N_10778,N_2304,N_5363);
nand U10779 (N_10779,N_1395,N_548);
and U10780 (N_10780,N_4255,N_5867);
xor U10781 (N_10781,N_3314,N_5493);
or U10782 (N_10782,N_5362,N_4863);
or U10783 (N_10783,N_351,N_5110);
nand U10784 (N_10784,N_4457,N_977);
nand U10785 (N_10785,N_2969,N_5571);
xnor U10786 (N_10786,N_3529,N_3389);
and U10787 (N_10787,N_2427,N_4365);
nand U10788 (N_10788,N_4827,N_3613);
nand U10789 (N_10789,N_5921,N_4001);
xnor U10790 (N_10790,N_5023,N_4332);
and U10791 (N_10791,N_192,N_5582);
or U10792 (N_10792,N_5992,N_1620);
nand U10793 (N_10793,N_541,N_5236);
and U10794 (N_10794,N_1318,N_5751);
or U10795 (N_10795,N_835,N_5628);
xor U10796 (N_10796,N_657,N_503);
or U10797 (N_10797,N_291,N_4721);
nor U10798 (N_10798,N_4482,N_3118);
nand U10799 (N_10799,N_4668,N_5151);
xnor U10800 (N_10800,N_1741,N_2682);
nand U10801 (N_10801,N_657,N_5075);
nand U10802 (N_10802,N_1972,N_4178);
xnor U10803 (N_10803,N_569,N_200);
nand U10804 (N_10804,N_5904,N_5743);
nand U10805 (N_10805,N_1293,N_96);
xnor U10806 (N_10806,N_5150,N_4400);
or U10807 (N_10807,N_3801,N_802);
nor U10808 (N_10808,N_216,N_2273);
nand U10809 (N_10809,N_1596,N_4083);
nand U10810 (N_10810,N_2119,N_2468);
or U10811 (N_10811,N_2638,N_1476);
nand U10812 (N_10812,N_304,N_217);
nand U10813 (N_10813,N_5194,N_4942);
xor U10814 (N_10814,N_5970,N_1799);
xnor U10815 (N_10815,N_5866,N_2738);
or U10816 (N_10816,N_2879,N_5560);
nor U10817 (N_10817,N_128,N_3152);
or U10818 (N_10818,N_162,N_2386);
nand U10819 (N_10819,N_4294,N_2545);
and U10820 (N_10820,N_876,N_3195);
and U10821 (N_10821,N_2282,N_4482);
nand U10822 (N_10822,N_3275,N_3080);
or U10823 (N_10823,N_3223,N_4438);
and U10824 (N_10824,N_5094,N_2860);
nand U10825 (N_10825,N_2539,N_5968);
or U10826 (N_10826,N_1740,N_1714);
nor U10827 (N_10827,N_2448,N_2137);
or U10828 (N_10828,N_5255,N_4534);
or U10829 (N_10829,N_396,N_5789);
and U10830 (N_10830,N_4671,N_353);
or U10831 (N_10831,N_26,N_2384);
nor U10832 (N_10832,N_4711,N_3280);
nand U10833 (N_10833,N_105,N_1295);
xnor U10834 (N_10834,N_5400,N_4699);
xnor U10835 (N_10835,N_1774,N_3766);
xnor U10836 (N_10836,N_527,N_2080);
nor U10837 (N_10837,N_5941,N_3183);
nor U10838 (N_10838,N_4317,N_5759);
nand U10839 (N_10839,N_1025,N_1038);
nor U10840 (N_10840,N_4705,N_2111);
nand U10841 (N_10841,N_3661,N_2560);
xor U10842 (N_10842,N_3869,N_3527);
nor U10843 (N_10843,N_5591,N_323);
xnor U10844 (N_10844,N_5782,N_2712);
nor U10845 (N_10845,N_4781,N_4980);
or U10846 (N_10846,N_4427,N_5382);
xor U10847 (N_10847,N_4527,N_322);
or U10848 (N_10848,N_5713,N_677);
xnor U10849 (N_10849,N_4762,N_623);
xor U10850 (N_10850,N_800,N_4468);
or U10851 (N_10851,N_5004,N_3158);
or U10852 (N_10852,N_5617,N_1900);
or U10853 (N_10853,N_5842,N_2155);
nor U10854 (N_10854,N_4483,N_2885);
nand U10855 (N_10855,N_5223,N_3473);
nor U10856 (N_10856,N_678,N_1645);
nor U10857 (N_10857,N_2965,N_2250);
xnor U10858 (N_10858,N_2403,N_4490);
xnor U10859 (N_10859,N_1350,N_4919);
nand U10860 (N_10860,N_2059,N_216);
or U10861 (N_10861,N_4384,N_5987);
xnor U10862 (N_10862,N_2103,N_794);
xnor U10863 (N_10863,N_316,N_2180);
xnor U10864 (N_10864,N_5497,N_4552);
nand U10865 (N_10865,N_3828,N_2990);
nand U10866 (N_10866,N_4428,N_5078);
or U10867 (N_10867,N_882,N_1873);
xor U10868 (N_10868,N_3568,N_3096);
nor U10869 (N_10869,N_5892,N_4564);
nor U10870 (N_10870,N_4463,N_4471);
nand U10871 (N_10871,N_3357,N_4564);
or U10872 (N_10872,N_1936,N_2776);
and U10873 (N_10873,N_5117,N_2623);
and U10874 (N_10874,N_1791,N_5928);
and U10875 (N_10875,N_142,N_1893);
or U10876 (N_10876,N_5194,N_5147);
or U10877 (N_10877,N_1469,N_1452);
xnor U10878 (N_10878,N_3222,N_502);
and U10879 (N_10879,N_5750,N_4439);
nand U10880 (N_10880,N_3726,N_230);
or U10881 (N_10881,N_3119,N_4443);
and U10882 (N_10882,N_3553,N_1231);
xor U10883 (N_10883,N_3844,N_5476);
nor U10884 (N_10884,N_866,N_5203);
xnor U10885 (N_10885,N_973,N_5497);
nand U10886 (N_10886,N_2010,N_1871);
xor U10887 (N_10887,N_4293,N_5608);
or U10888 (N_10888,N_428,N_4171);
nor U10889 (N_10889,N_4888,N_5983);
xnor U10890 (N_10890,N_2004,N_3967);
and U10891 (N_10891,N_3428,N_5948);
and U10892 (N_10892,N_4641,N_5629);
nor U10893 (N_10893,N_435,N_1075);
nand U10894 (N_10894,N_1632,N_3533);
and U10895 (N_10895,N_3676,N_136);
nor U10896 (N_10896,N_4146,N_2881);
nand U10897 (N_10897,N_5710,N_1265);
nand U10898 (N_10898,N_1901,N_541);
or U10899 (N_10899,N_5444,N_4307);
nand U10900 (N_10900,N_5734,N_4092);
nor U10901 (N_10901,N_1464,N_5410);
xnor U10902 (N_10902,N_2839,N_5678);
and U10903 (N_10903,N_5130,N_4826);
and U10904 (N_10904,N_4206,N_902);
nor U10905 (N_10905,N_814,N_1278);
xnor U10906 (N_10906,N_5765,N_2715);
or U10907 (N_10907,N_5377,N_5521);
nand U10908 (N_10908,N_4779,N_506);
nor U10909 (N_10909,N_884,N_859);
nand U10910 (N_10910,N_4284,N_3366);
nor U10911 (N_10911,N_111,N_3303);
and U10912 (N_10912,N_3428,N_662);
or U10913 (N_10913,N_1656,N_3050);
nor U10914 (N_10914,N_1433,N_3955);
and U10915 (N_10915,N_2990,N_1568);
and U10916 (N_10916,N_4719,N_3911);
xor U10917 (N_10917,N_3800,N_2492);
nand U10918 (N_10918,N_2282,N_1347);
nand U10919 (N_10919,N_142,N_5653);
and U10920 (N_10920,N_1503,N_2665);
and U10921 (N_10921,N_1857,N_2552);
xor U10922 (N_10922,N_1503,N_5346);
nor U10923 (N_10923,N_4439,N_1399);
nand U10924 (N_10924,N_4836,N_5703);
nand U10925 (N_10925,N_2649,N_5060);
nand U10926 (N_10926,N_3434,N_1560);
xnor U10927 (N_10927,N_2305,N_1140);
or U10928 (N_10928,N_3675,N_4325);
and U10929 (N_10929,N_541,N_3269);
xor U10930 (N_10930,N_2953,N_2532);
nor U10931 (N_10931,N_4669,N_5157);
xor U10932 (N_10932,N_3514,N_3750);
or U10933 (N_10933,N_450,N_1288);
xnor U10934 (N_10934,N_1268,N_752);
nor U10935 (N_10935,N_5490,N_1923);
xnor U10936 (N_10936,N_4615,N_4051);
xor U10937 (N_10937,N_4139,N_2561);
and U10938 (N_10938,N_3956,N_2086);
xnor U10939 (N_10939,N_2489,N_2640);
and U10940 (N_10940,N_794,N_5336);
xor U10941 (N_10941,N_2375,N_1910);
nor U10942 (N_10942,N_1428,N_2847);
nor U10943 (N_10943,N_4448,N_3622);
or U10944 (N_10944,N_2541,N_4653);
and U10945 (N_10945,N_2600,N_941);
and U10946 (N_10946,N_4648,N_2870);
xor U10947 (N_10947,N_1545,N_2626);
or U10948 (N_10948,N_2717,N_3394);
and U10949 (N_10949,N_4144,N_5652);
or U10950 (N_10950,N_4027,N_4906);
xor U10951 (N_10951,N_4470,N_5097);
or U10952 (N_10952,N_503,N_3666);
or U10953 (N_10953,N_1272,N_4585);
nand U10954 (N_10954,N_1090,N_460);
nor U10955 (N_10955,N_3904,N_4764);
nand U10956 (N_10956,N_5386,N_3502);
or U10957 (N_10957,N_2512,N_4581);
nor U10958 (N_10958,N_377,N_5854);
nor U10959 (N_10959,N_2417,N_1898);
nand U10960 (N_10960,N_2000,N_2708);
or U10961 (N_10961,N_3035,N_5827);
nor U10962 (N_10962,N_1604,N_643);
xnor U10963 (N_10963,N_180,N_5156);
nor U10964 (N_10964,N_2583,N_702);
xnor U10965 (N_10965,N_4291,N_3002);
or U10966 (N_10966,N_4006,N_4064);
or U10967 (N_10967,N_4701,N_5230);
or U10968 (N_10968,N_4163,N_3529);
and U10969 (N_10969,N_5543,N_1912);
nand U10970 (N_10970,N_839,N_3771);
xnor U10971 (N_10971,N_430,N_407);
nor U10972 (N_10972,N_611,N_5386);
and U10973 (N_10973,N_5722,N_5869);
and U10974 (N_10974,N_4238,N_3767);
or U10975 (N_10975,N_3469,N_2785);
nor U10976 (N_10976,N_4151,N_1428);
nand U10977 (N_10977,N_4676,N_1444);
xnor U10978 (N_10978,N_1324,N_4147);
xnor U10979 (N_10979,N_811,N_3980);
nand U10980 (N_10980,N_5838,N_2518);
and U10981 (N_10981,N_3578,N_87);
nor U10982 (N_10982,N_2585,N_1636);
nor U10983 (N_10983,N_2676,N_1291);
nand U10984 (N_10984,N_1972,N_5670);
and U10985 (N_10985,N_5602,N_860);
nor U10986 (N_10986,N_2693,N_5264);
nand U10987 (N_10987,N_1681,N_381);
or U10988 (N_10988,N_3108,N_2176);
and U10989 (N_10989,N_261,N_1811);
xnor U10990 (N_10990,N_1790,N_2312);
nor U10991 (N_10991,N_2051,N_4627);
nor U10992 (N_10992,N_1157,N_1012);
nor U10993 (N_10993,N_5134,N_1049);
nand U10994 (N_10994,N_2575,N_3697);
xnor U10995 (N_10995,N_4377,N_5717);
xor U10996 (N_10996,N_3447,N_2020);
xnor U10997 (N_10997,N_3686,N_3872);
nand U10998 (N_10998,N_1951,N_2164);
or U10999 (N_10999,N_1840,N_957);
and U11000 (N_11000,N_2993,N_4134);
or U11001 (N_11001,N_918,N_2044);
xnor U11002 (N_11002,N_5175,N_2183);
xnor U11003 (N_11003,N_5401,N_5917);
xor U11004 (N_11004,N_977,N_231);
nand U11005 (N_11005,N_539,N_3379);
xnor U11006 (N_11006,N_4140,N_3299);
xnor U11007 (N_11007,N_1585,N_5650);
or U11008 (N_11008,N_2806,N_1769);
or U11009 (N_11009,N_3023,N_2497);
nor U11010 (N_11010,N_2206,N_1298);
xor U11011 (N_11011,N_4085,N_2195);
nor U11012 (N_11012,N_1042,N_3491);
nor U11013 (N_11013,N_5921,N_774);
nand U11014 (N_11014,N_2672,N_613);
nor U11015 (N_11015,N_1299,N_1757);
xor U11016 (N_11016,N_2889,N_1242);
nor U11017 (N_11017,N_1120,N_1324);
xor U11018 (N_11018,N_3149,N_4678);
or U11019 (N_11019,N_720,N_1323);
xnor U11020 (N_11020,N_5947,N_2234);
and U11021 (N_11021,N_3786,N_2498);
or U11022 (N_11022,N_5670,N_5295);
nand U11023 (N_11023,N_924,N_2568);
xor U11024 (N_11024,N_569,N_576);
nand U11025 (N_11025,N_5556,N_3493);
and U11026 (N_11026,N_2165,N_1351);
and U11027 (N_11027,N_5304,N_2951);
nor U11028 (N_11028,N_4657,N_2853);
xor U11029 (N_11029,N_450,N_1930);
nor U11030 (N_11030,N_2285,N_5563);
and U11031 (N_11031,N_3099,N_2126);
xnor U11032 (N_11032,N_1495,N_5846);
and U11033 (N_11033,N_1928,N_4917);
and U11034 (N_11034,N_3392,N_2450);
and U11035 (N_11035,N_352,N_3287);
or U11036 (N_11036,N_1728,N_3246);
nor U11037 (N_11037,N_5075,N_4342);
nor U11038 (N_11038,N_3578,N_4636);
nor U11039 (N_11039,N_4353,N_4219);
and U11040 (N_11040,N_4277,N_3640);
or U11041 (N_11041,N_5646,N_4877);
xor U11042 (N_11042,N_2690,N_3339);
or U11043 (N_11043,N_3838,N_3540);
xor U11044 (N_11044,N_4909,N_1358);
or U11045 (N_11045,N_1394,N_4260);
nand U11046 (N_11046,N_5829,N_3);
or U11047 (N_11047,N_3115,N_2009);
or U11048 (N_11048,N_1422,N_385);
or U11049 (N_11049,N_2906,N_4449);
xnor U11050 (N_11050,N_5389,N_3839);
and U11051 (N_11051,N_2879,N_1076);
nor U11052 (N_11052,N_1663,N_1960);
nand U11053 (N_11053,N_2704,N_1808);
xor U11054 (N_11054,N_4052,N_3871);
xor U11055 (N_11055,N_599,N_5974);
nor U11056 (N_11056,N_1725,N_2093);
nor U11057 (N_11057,N_610,N_1394);
nand U11058 (N_11058,N_1086,N_2454);
or U11059 (N_11059,N_573,N_3601);
nor U11060 (N_11060,N_392,N_3812);
nor U11061 (N_11061,N_1041,N_1754);
or U11062 (N_11062,N_4909,N_3406);
xor U11063 (N_11063,N_4098,N_5968);
nor U11064 (N_11064,N_2983,N_2588);
and U11065 (N_11065,N_2439,N_4560);
nor U11066 (N_11066,N_807,N_4758);
or U11067 (N_11067,N_5086,N_2589);
or U11068 (N_11068,N_334,N_2841);
nor U11069 (N_11069,N_5987,N_5841);
nor U11070 (N_11070,N_1550,N_1639);
xor U11071 (N_11071,N_630,N_1422);
and U11072 (N_11072,N_1733,N_447);
and U11073 (N_11073,N_159,N_4264);
nor U11074 (N_11074,N_3108,N_4007);
nor U11075 (N_11075,N_4097,N_4890);
or U11076 (N_11076,N_3364,N_2526);
nand U11077 (N_11077,N_1736,N_2192);
xnor U11078 (N_11078,N_5792,N_4535);
xor U11079 (N_11079,N_2377,N_4551);
nand U11080 (N_11080,N_4646,N_5496);
and U11081 (N_11081,N_4853,N_5959);
and U11082 (N_11082,N_92,N_3895);
nor U11083 (N_11083,N_115,N_1831);
and U11084 (N_11084,N_1736,N_4063);
xor U11085 (N_11085,N_1901,N_668);
xnor U11086 (N_11086,N_4677,N_5220);
nor U11087 (N_11087,N_245,N_5688);
nor U11088 (N_11088,N_2441,N_5203);
nand U11089 (N_11089,N_318,N_5485);
or U11090 (N_11090,N_2258,N_2023);
xor U11091 (N_11091,N_4224,N_5237);
xor U11092 (N_11092,N_4478,N_2496);
or U11093 (N_11093,N_4377,N_1777);
xnor U11094 (N_11094,N_4482,N_5851);
nor U11095 (N_11095,N_3769,N_1051);
xnor U11096 (N_11096,N_2909,N_5124);
xor U11097 (N_11097,N_3986,N_2815);
xnor U11098 (N_11098,N_886,N_5050);
and U11099 (N_11099,N_992,N_5030);
nor U11100 (N_11100,N_5084,N_5510);
nand U11101 (N_11101,N_5064,N_2093);
nand U11102 (N_11102,N_3866,N_401);
xor U11103 (N_11103,N_3108,N_2761);
or U11104 (N_11104,N_5652,N_2249);
or U11105 (N_11105,N_1448,N_835);
and U11106 (N_11106,N_5404,N_5523);
or U11107 (N_11107,N_2395,N_4597);
xor U11108 (N_11108,N_2052,N_4177);
and U11109 (N_11109,N_3326,N_2798);
xnor U11110 (N_11110,N_242,N_1235);
and U11111 (N_11111,N_5484,N_1434);
nor U11112 (N_11112,N_4569,N_3512);
and U11113 (N_11113,N_1718,N_3668);
xnor U11114 (N_11114,N_4936,N_555);
and U11115 (N_11115,N_2462,N_2829);
xor U11116 (N_11116,N_3182,N_649);
or U11117 (N_11117,N_3174,N_551);
xor U11118 (N_11118,N_1807,N_4865);
nand U11119 (N_11119,N_307,N_4844);
nand U11120 (N_11120,N_1382,N_586);
nor U11121 (N_11121,N_5377,N_4538);
or U11122 (N_11122,N_4834,N_3653);
nand U11123 (N_11123,N_265,N_382);
nand U11124 (N_11124,N_2489,N_4660);
or U11125 (N_11125,N_2347,N_4571);
and U11126 (N_11126,N_1286,N_3062);
xor U11127 (N_11127,N_2352,N_5143);
nand U11128 (N_11128,N_2419,N_885);
nand U11129 (N_11129,N_3901,N_4998);
xnor U11130 (N_11130,N_4618,N_5766);
or U11131 (N_11131,N_2264,N_3921);
xnor U11132 (N_11132,N_5027,N_241);
xor U11133 (N_11133,N_4349,N_4143);
nand U11134 (N_11134,N_1486,N_2784);
or U11135 (N_11135,N_1093,N_1355);
or U11136 (N_11136,N_5478,N_1115);
or U11137 (N_11137,N_5414,N_3978);
xnor U11138 (N_11138,N_2798,N_2968);
xnor U11139 (N_11139,N_1029,N_810);
nor U11140 (N_11140,N_888,N_1502);
and U11141 (N_11141,N_4908,N_2063);
and U11142 (N_11142,N_3652,N_3747);
and U11143 (N_11143,N_2052,N_2417);
or U11144 (N_11144,N_1992,N_5216);
xor U11145 (N_11145,N_5562,N_4826);
nand U11146 (N_11146,N_5899,N_573);
nor U11147 (N_11147,N_939,N_715);
nor U11148 (N_11148,N_928,N_4498);
nand U11149 (N_11149,N_723,N_2070);
nor U11150 (N_11150,N_5651,N_2865);
nor U11151 (N_11151,N_1729,N_4925);
nor U11152 (N_11152,N_1853,N_1178);
or U11153 (N_11153,N_5846,N_4409);
xnor U11154 (N_11154,N_4763,N_2327);
or U11155 (N_11155,N_3262,N_705);
nor U11156 (N_11156,N_2667,N_4000);
and U11157 (N_11157,N_4901,N_2784);
nand U11158 (N_11158,N_4372,N_894);
nor U11159 (N_11159,N_4665,N_4655);
nand U11160 (N_11160,N_5250,N_3511);
or U11161 (N_11161,N_5417,N_5979);
nand U11162 (N_11162,N_3196,N_3135);
and U11163 (N_11163,N_2743,N_2658);
or U11164 (N_11164,N_5673,N_479);
xor U11165 (N_11165,N_4528,N_2189);
xor U11166 (N_11166,N_2799,N_539);
and U11167 (N_11167,N_5506,N_4284);
or U11168 (N_11168,N_216,N_352);
xnor U11169 (N_11169,N_1449,N_5845);
nand U11170 (N_11170,N_1175,N_5384);
xnor U11171 (N_11171,N_1267,N_2663);
nand U11172 (N_11172,N_2061,N_3669);
or U11173 (N_11173,N_1397,N_3257);
nand U11174 (N_11174,N_4518,N_4411);
nor U11175 (N_11175,N_2524,N_2172);
and U11176 (N_11176,N_5553,N_2588);
xor U11177 (N_11177,N_2224,N_3386);
and U11178 (N_11178,N_4498,N_2065);
nand U11179 (N_11179,N_3051,N_3735);
xor U11180 (N_11180,N_709,N_1815);
xor U11181 (N_11181,N_5645,N_5951);
xnor U11182 (N_11182,N_3201,N_4057);
or U11183 (N_11183,N_4020,N_5666);
nand U11184 (N_11184,N_1227,N_4769);
and U11185 (N_11185,N_247,N_5027);
nor U11186 (N_11186,N_4750,N_4495);
nand U11187 (N_11187,N_2031,N_3480);
xnor U11188 (N_11188,N_3825,N_3800);
xnor U11189 (N_11189,N_2749,N_597);
nand U11190 (N_11190,N_2067,N_4053);
and U11191 (N_11191,N_3354,N_5568);
nor U11192 (N_11192,N_79,N_2346);
nand U11193 (N_11193,N_3138,N_5554);
or U11194 (N_11194,N_2459,N_3898);
xnor U11195 (N_11195,N_1004,N_4822);
nand U11196 (N_11196,N_608,N_5673);
and U11197 (N_11197,N_5691,N_244);
xor U11198 (N_11198,N_3932,N_2876);
nor U11199 (N_11199,N_4361,N_1453);
nor U11200 (N_11200,N_5220,N_2591);
xnor U11201 (N_11201,N_1097,N_5757);
and U11202 (N_11202,N_1952,N_1478);
nor U11203 (N_11203,N_4806,N_2248);
xor U11204 (N_11204,N_5289,N_4129);
nand U11205 (N_11205,N_2170,N_2225);
nor U11206 (N_11206,N_5316,N_448);
nand U11207 (N_11207,N_2292,N_1043);
or U11208 (N_11208,N_2690,N_5074);
xor U11209 (N_11209,N_5885,N_4267);
xor U11210 (N_11210,N_1184,N_1347);
xnor U11211 (N_11211,N_884,N_5075);
and U11212 (N_11212,N_5256,N_2280);
and U11213 (N_11213,N_4720,N_2638);
xnor U11214 (N_11214,N_4260,N_3799);
xnor U11215 (N_11215,N_5284,N_2107);
or U11216 (N_11216,N_3579,N_420);
or U11217 (N_11217,N_3990,N_352);
nand U11218 (N_11218,N_1989,N_4218);
nor U11219 (N_11219,N_5295,N_2469);
or U11220 (N_11220,N_2643,N_321);
or U11221 (N_11221,N_416,N_316);
and U11222 (N_11222,N_735,N_4525);
and U11223 (N_11223,N_1088,N_374);
nand U11224 (N_11224,N_3704,N_4745);
nor U11225 (N_11225,N_5416,N_1748);
xor U11226 (N_11226,N_5742,N_4405);
and U11227 (N_11227,N_1028,N_5871);
nor U11228 (N_11228,N_4126,N_1853);
xnor U11229 (N_11229,N_5279,N_4272);
and U11230 (N_11230,N_985,N_1888);
or U11231 (N_11231,N_3946,N_240);
nor U11232 (N_11232,N_238,N_99);
nand U11233 (N_11233,N_4816,N_5026);
nand U11234 (N_11234,N_2890,N_1742);
xor U11235 (N_11235,N_3533,N_5646);
nand U11236 (N_11236,N_2791,N_4701);
nand U11237 (N_11237,N_2947,N_875);
nand U11238 (N_11238,N_2516,N_2096);
xor U11239 (N_11239,N_5831,N_3091);
nand U11240 (N_11240,N_5463,N_2019);
nor U11241 (N_11241,N_3680,N_4688);
or U11242 (N_11242,N_1562,N_2753);
nor U11243 (N_11243,N_4020,N_5006);
and U11244 (N_11244,N_1929,N_3685);
nand U11245 (N_11245,N_2250,N_1925);
or U11246 (N_11246,N_4039,N_1890);
xor U11247 (N_11247,N_5517,N_3977);
xnor U11248 (N_11248,N_2737,N_5998);
or U11249 (N_11249,N_4716,N_5328);
or U11250 (N_11250,N_703,N_5235);
nor U11251 (N_11251,N_4758,N_559);
and U11252 (N_11252,N_4107,N_1725);
xnor U11253 (N_11253,N_2309,N_1464);
xor U11254 (N_11254,N_4064,N_5156);
or U11255 (N_11255,N_4593,N_4494);
nand U11256 (N_11256,N_1493,N_2156);
nand U11257 (N_11257,N_4319,N_4830);
and U11258 (N_11258,N_1959,N_5772);
or U11259 (N_11259,N_3316,N_993);
nand U11260 (N_11260,N_2044,N_4680);
nand U11261 (N_11261,N_5058,N_4112);
or U11262 (N_11262,N_5649,N_4781);
xnor U11263 (N_11263,N_466,N_1646);
and U11264 (N_11264,N_5877,N_3056);
xnor U11265 (N_11265,N_327,N_3037);
or U11266 (N_11266,N_1617,N_5717);
nand U11267 (N_11267,N_2828,N_2482);
and U11268 (N_11268,N_727,N_5339);
nand U11269 (N_11269,N_1356,N_4328);
xor U11270 (N_11270,N_3229,N_5960);
nor U11271 (N_11271,N_5829,N_350);
and U11272 (N_11272,N_814,N_5902);
and U11273 (N_11273,N_1131,N_4659);
and U11274 (N_11274,N_5790,N_269);
nor U11275 (N_11275,N_5179,N_3431);
xnor U11276 (N_11276,N_4594,N_3587);
nor U11277 (N_11277,N_4608,N_2280);
or U11278 (N_11278,N_4599,N_227);
and U11279 (N_11279,N_5227,N_624);
nor U11280 (N_11280,N_2333,N_3085);
or U11281 (N_11281,N_92,N_4161);
or U11282 (N_11282,N_4119,N_5663);
nand U11283 (N_11283,N_3000,N_862);
nor U11284 (N_11284,N_1036,N_2754);
xor U11285 (N_11285,N_1238,N_3944);
xnor U11286 (N_11286,N_1313,N_5584);
xor U11287 (N_11287,N_3758,N_3029);
and U11288 (N_11288,N_2212,N_4646);
and U11289 (N_11289,N_5799,N_1465);
xor U11290 (N_11290,N_5627,N_4452);
xnor U11291 (N_11291,N_2069,N_1618);
xor U11292 (N_11292,N_3097,N_3527);
and U11293 (N_11293,N_256,N_4475);
xnor U11294 (N_11294,N_364,N_1465);
or U11295 (N_11295,N_1933,N_3701);
xor U11296 (N_11296,N_2500,N_2411);
nor U11297 (N_11297,N_4584,N_5961);
nand U11298 (N_11298,N_5210,N_619);
xnor U11299 (N_11299,N_5185,N_3151);
nand U11300 (N_11300,N_1929,N_1433);
nand U11301 (N_11301,N_4022,N_270);
or U11302 (N_11302,N_1780,N_4139);
and U11303 (N_11303,N_1779,N_2199);
and U11304 (N_11304,N_1622,N_3629);
xnor U11305 (N_11305,N_1303,N_2638);
and U11306 (N_11306,N_2575,N_4844);
or U11307 (N_11307,N_2282,N_3829);
xnor U11308 (N_11308,N_4578,N_28);
or U11309 (N_11309,N_2969,N_3265);
nor U11310 (N_11310,N_3475,N_89);
or U11311 (N_11311,N_1881,N_119);
and U11312 (N_11312,N_2078,N_1011);
and U11313 (N_11313,N_4677,N_4700);
and U11314 (N_11314,N_873,N_1726);
and U11315 (N_11315,N_1688,N_2384);
nand U11316 (N_11316,N_3362,N_128);
nand U11317 (N_11317,N_385,N_4099);
nand U11318 (N_11318,N_5728,N_2315);
and U11319 (N_11319,N_3592,N_3275);
or U11320 (N_11320,N_4958,N_555);
and U11321 (N_11321,N_2576,N_4727);
and U11322 (N_11322,N_3920,N_4953);
xnor U11323 (N_11323,N_725,N_4575);
or U11324 (N_11324,N_5446,N_1250);
xor U11325 (N_11325,N_1145,N_2765);
xor U11326 (N_11326,N_3130,N_4422);
and U11327 (N_11327,N_2017,N_3237);
nor U11328 (N_11328,N_4780,N_5274);
or U11329 (N_11329,N_1238,N_1134);
nand U11330 (N_11330,N_3895,N_1012);
and U11331 (N_11331,N_3100,N_4202);
and U11332 (N_11332,N_190,N_1470);
nor U11333 (N_11333,N_4244,N_3258);
xnor U11334 (N_11334,N_101,N_4011);
xor U11335 (N_11335,N_460,N_1341);
nor U11336 (N_11336,N_3406,N_241);
nor U11337 (N_11337,N_2065,N_1258);
nand U11338 (N_11338,N_2052,N_554);
nand U11339 (N_11339,N_3955,N_2118);
nand U11340 (N_11340,N_3302,N_5084);
nand U11341 (N_11341,N_2501,N_4082);
nand U11342 (N_11342,N_4616,N_1915);
or U11343 (N_11343,N_2155,N_1479);
xnor U11344 (N_11344,N_471,N_3037);
nand U11345 (N_11345,N_738,N_3674);
and U11346 (N_11346,N_5093,N_2668);
and U11347 (N_11347,N_4130,N_5798);
nor U11348 (N_11348,N_1245,N_717);
or U11349 (N_11349,N_4043,N_2110);
nor U11350 (N_11350,N_2533,N_1853);
and U11351 (N_11351,N_3806,N_4680);
xor U11352 (N_11352,N_3788,N_2545);
and U11353 (N_11353,N_4603,N_1159);
and U11354 (N_11354,N_5658,N_4482);
xor U11355 (N_11355,N_1640,N_3570);
nor U11356 (N_11356,N_5885,N_4977);
nand U11357 (N_11357,N_4514,N_3196);
xor U11358 (N_11358,N_521,N_4709);
nand U11359 (N_11359,N_1745,N_2846);
or U11360 (N_11360,N_4547,N_908);
xor U11361 (N_11361,N_5194,N_1089);
xor U11362 (N_11362,N_2464,N_2737);
nand U11363 (N_11363,N_3365,N_4241);
nor U11364 (N_11364,N_2012,N_5594);
nor U11365 (N_11365,N_3066,N_3423);
nand U11366 (N_11366,N_5897,N_1455);
nor U11367 (N_11367,N_1143,N_5056);
and U11368 (N_11368,N_1677,N_1852);
or U11369 (N_11369,N_4024,N_5272);
nor U11370 (N_11370,N_3764,N_417);
xnor U11371 (N_11371,N_5562,N_148);
xor U11372 (N_11372,N_359,N_3076);
nor U11373 (N_11373,N_4714,N_5255);
xor U11374 (N_11374,N_4116,N_893);
and U11375 (N_11375,N_5330,N_5910);
nor U11376 (N_11376,N_4886,N_4610);
and U11377 (N_11377,N_955,N_5271);
nand U11378 (N_11378,N_5291,N_1857);
or U11379 (N_11379,N_2249,N_1989);
and U11380 (N_11380,N_1110,N_4974);
or U11381 (N_11381,N_3857,N_3654);
xnor U11382 (N_11382,N_3883,N_5541);
and U11383 (N_11383,N_4928,N_2531);
or U11384 (N_11384,N_4724,N_5859);
xor U11385 (N_11385,N_1017,N_5685);
or U11386 (N_11386,N_1276,N_3883);
xor U11387 (N_11387,N_4201,N_1531);
nand U11388 (N_11388,N_884,N_5634);
and U11389 (N_11389,N_2566,N_2608);
or U11390 (N_11390,N_3087,N_1564);
xor U11391 (N_11391,N_2358,N_1028);
nor U11392 (N_11392,N_1977,N_1891);
nand U11393 (N_11393,N_4225,N_3780);
nor U11394 (N_11394,N_4005,N_4610);
and U11395 (N_11395,N_3793,N_3638);
and U11396 (N_11396,N_5466,N_932);
nor U11397 (N_11397,N_5023,N_5102);
and U11398 (N_11398,N_5045,N_4757);
and U11399 (N_11399,N_1621,N_5807);
nor U11400 (N_11400,N_1389,N_2936);
nor U11401 (N_11401,N_3197,N_3556);
or U11402 (N_11402,N_2083,N_2506);
and U11403 (N_11403,N_4060,N_36);
nand U11404 (N_11404,N_2366,N_315);
or U11405 (N_11405,N_3834,N_3401);
or U11406 (N_11406,N_789,N_3074);
and U11407 (N_11407,N_1915,N_5617);
nor U11408 (N_11408,N_4712,N_255);
xnor U11409 (N_11409,N_4329,N_5721);
or U11410 (N_11410,N_3449,N_1236);
nand U11411 (N_11411,N_4859,N_4284);
xor U11412 (N_11412,N_4467,N_3664);
and U11413 (N_11413,N_5011,N_3980);
xnor U11414 (N_11414,N_546,N_4005);
or U11415 (N_11415,N_1417,N_2304);
and U11416 (N_11416,N_898,N_333);
or U11417 (N_11417,N_5124,N_3646);
nand U11418 (N_11418,N_4690,N_829);
nor U11419 (N_11419,N_2986,N_2890);
nor U11420 (N_11420,N_5665,N_2068);
or U11421 (N_11421,N_3188,N_1574);
nand U11422 (N_11422,N_992,N_3461);
and U11423 (N_11423,N_2467,N_114);
nor U11424 (N_11424,N_2797,N_318);
xor U11425 (N_11425,N_3281,N_752);
nand U11426 (N_11426,N_3211,N_5072);
nand U11427 (N_11427,N_4217,N_5076);
or U11428 (N_11428,N_5662,N_2251);
xnor U11429 (N_11429,N_1816,N_1207);
or U11430 (N_11430,N_2938,N_4138);
or U11431 (N_11431,N_1209,N_4435);
nor U11432 (N_11432,N_2452,N_5190);
and U11433 (N_11433,N_5084,N_422);
xnor U11434 (N_11434,N_1070,N_1310);
or U11435 (N_11435,N_655,N_4846);
xnor U11436 (N_11436,N_621,N_4964);
xnor U11437 (N_11437,N_4214,N_230);
and U11438 (N_11438,N_761,N_56);
and U11439 (N_11439,N_1093,N_2809);
and U11440 (N_11440,N_5546,N_5716);
and U11441 (N_11441,N_5919,N_4082);
xor U11442 (N_11442,N_5162,N_365);
or U11443 (N_11443,N_5977,N_4674);
or U11444 (N_11444,N_1018,N_1357);
or U11445 (N_11445,N_3994,N_123);
nand U11446 (N_11446,N_606,N_287);
and U11447 (N_11447,N_2034,N_1771);
nor U11448 (N_11448,N_3911,N_4081);
xor U11449 (N_11449,N_1341,N_729);
xor U11450 (N_11450,N_2280,N_137);
nand U11451 (N_11451,N_4334,N_4986);
nor U11452 (N_11452,N_4917,N_2366);
xnor U11453 (N_11453,N_2700,N_3451);
nand U11454 (N_11454,N_2574,N_2381);
nor U11455 (N_11455,N_3578,N_645);
or U11456 (N_11456,N_4235,N_686);
nand U11457 (N_11457,N_484,N_1324);
or U11458 (N_11458,N_4459,N_3595);
nor U11459 (N_11459,N_5368,N_653);
nor U11460 (N_11460,N_1541,N_1162);
or U11461 (N_11461,N_751,N_2127);
or U11462 (N_11462,N_2816,N_1363);
or U11463 (N_11463,N_5484,N_4963);
nand U11464 (N_11464,N_2288,N_5700);
and U11465 (N_11465,N_1062,N_4626);
or U11466 (N_11466,N_5713,N_2370);
nand U11467 (N_11467,N_1294,N_5938);
or U11468 (N_11468,N_5206,N_4450);
and U11469 (N_11469,N_3884,N_5037);
nand U11470 (N_11470,N_1435,N_1894);
xnor U11471 (N_11471,N_4661,N_5647);
and U11472 (N_11472,N_5574,N_5740);
xor U11473 (N_11473,N_2846,N_3386);
or U11474 (N_11474,N_3303,N_3439);
xor U11475 (N_11475,N_5886,N_5348);
nand U11476 (N_11476,N_3267,N_2695);
xor U11477 (N_11477,N_3763,N_1748);
nand U11478 (N_11478,N_422,N_1819);
and U11479 (N_11479,N_4110,N_5995);
nand U11480 (N_11480,N_1664,N_3456);
nand U11481 (N_11481,N_1977,N_2430);
nand U11482 (N_11482,N_4470,N_2242);
nor U11483 (N_11483,N_3519,N_5399);
nor U11484 (N_11484,N_5479,N_3719);
and U11485 (N_11485,N_2410,N_1853);
or U11486 (N_11486,N_5709,N_4536);
nand U11487 (N_11487,N_442,N_3179);
nand U11488 (N_11488,N_1082,N_1247);
nand U11489 (N_11489,N_1604,N_1153);
or U11490 (N_11490,N_845,N_2871);
or U11491 (N_11491,N_4800,N_1172);
or U11492 (N_11492,N_3827,N_3772);
or U11493 (N_11493,N_5421,N_341);
and U11494 (N_11494,N_1508,N_4029);
xnor U11495 (N_11495,N_1781,N_742);
or U11496 (N_11496,N_1864,N_596);
nand U11497 (N_11497,N_3657,N_989);
xnor U11498 (N_11498,N_1302,N_3717);
and U11499 (N_11499,N_494,N_70);
xor U11500 (N_11500,N_4526,N_880);
or U11501 (N_11501,N_5296,N_478);
nor U11502 (N_11502,N_5673,N_3272);
and U11503 (N_11503,N_1077,N_3851);
and U11504 (N_11504,N_3680,N_2050);
nand U11505 (N_11505,N_4715,N_1382);
nor U11506 (N_11506,N_222,N_4572);
nand U11507 (N_11507,N_2981,N_5293);
or U11508 (N_11508,N_5379,N_3493);
and U11509 (N_11509,N_183,N_3507);
and U11510 (N_11510,N_845,N_2681);
xor U11511 (N_11511,N_4051,N_2173);
xor U11512 (N_11512,N_62,N_747);
and U11513 (N_11513,N_5680,N_5785);
or U11514 (N_11514,N_5146,N_781);
xor U11515 (N_11515,N_2789,N_3713);
or U11516 (N_11516,N_3875,N_2948);
xnor U11517 (N_11517,N_1237,N_105);
nand U11518 (N_11518,N_3768,N_237);
nor U11519 (N_11519,N_5067,N_856);
nand U11520 (N_11520,N_5298,N_4431);
and U11521 (N_11521,N_3526,N_5603);
nor U11522 (N_11522,N_4547,N_590);
and U11523 (N_11523,N_1420,N_3476);
and U11524 (N_11524,N_3946,N_551);
xnor U11525 (N_11525,N_3649,N_1941);
nor U11526 (N_11526,N_1674,N_4727);
nor U11527 (N_11527,N_4515,N_3392);
nor U11528 (N_11528,N_308,N_2113);
xnor U11529 (N_11529,N_2900,N_532);
xnor U11530 (N_11530,N_1605,N_1359);
xnor U11531 (N_11531,N_1284,N_4496);
nand U11532 (N_11532,N_497,N_5534);
or U11533 (N_11533,N_5031,N_5293);
xnor U11534 (N_11534,N_4606,N_963);
nand U11535 (N_11535,N_4096,N_3029);
or U11536 (N_11536,N_2131,N_2368);
and U11537 (N_11537,N_4370,N_2489);
nor U11538 (N_11538,N_941,N_2014);
nand U11539 (N_11539,N_3732,N_3876);
xor U11540 (N_11540,N_2085,N_3277);
nor U11541 (N_11541,N_807,N_1412);
nand U11542 (N_11542,N_4177,N_3622);
nand U11543 (N_11543,N_2256,N_4792);
nor U11544 (N_11544,N_896,N_5160);
xor U11545 (N_11545,N_4793,N_5836);
nand U11546 (N_11546,N_1854,N_2274);
xnor U11547 (N_11547,N_4270,N_5814);
xor U11548 (N_11548,N_1077,N_5401);
xor U11549 (N_11549,N_5117,N_313);
and U11550 (N_11550,N_328,N_3469);
nor U11551 (N_11551,N_1804,N_2940);
or U11552 (N_11552,N_2864,N_1244);
nand U11553 (N_11553,N_472,N_5632);
nand U11554 (N_11554,N_979,N_3033);
nand U11555 (N_11555,N_3012,N_1366);
nand U11556 (N_11556,N_5872,N_2879);
xnor U11557 (N_11557,N_975,N_1504);
and U11558 (N_11558,N_2785,N_1798);
xnor U11559 (N_11559,N_1099,N_1123);
nor U11560 (N_11560,N_3346,N_3088);
and U11561 (N_11561,N_5782,N_3701);
and U11562 (N_11562,N_3264,N_4457);
or U11563 (N_11563,N_1390,N_1447);
nor U11564 (N_11564,N_2003,N_4261);
nor U11565 (N_11565,N_5957,N_5921);
nand U11566 (N_11566,N_1265,N_810);
nand U11567 (N_11567,N_2208,N_1921);
or U11568 (N_11568,N_1967,N_5612);
or U11569 (N_11569,N_1514,N_4649);
xnor U11570 (N_11570,N_3779,N_5689);
or U11571 (N_11571,N_5923,N_1735);
nor U11572 (N_11572,N_2252,N_4784);
nor U11573 (N_11573,N_3920,N_2047);
xnor U11574 (N_11574,N_4668,N_2396);
or U11575 (N_11575,N_3128,N_3387);
xnor U11576 (N_11576,N_3783,N_1182);
and U11577 (N_11577,N_3021,N_442);
nand U11578 (N_11578,N_1199,N_5384);
nor U11579 (N_11579,N_146,N_2477);
nand U11580 (N_11580,N_2050,N_5529);
nand U11581 (N_11581,N_85,N_4814);
xnor U11582 (N_11582,N_3167,N_265);
or U11583 (N_11583,N_4377,N_2129);
xor U11584 (N_11584,N_64,N_3361);
nor U11585 (N_11585,N_3073,N_875);
xor U11586 (N_11586,N_1017,N_957);
or U11587 (N_11587,N_2184,N_2661);
and U11588 (N_11588,N_1778,N_763);
nor U11589 (N_11589,N_2733,N_1061);
nand U11590 (N_11590,N_5259,N_3845);
and U11591 (N_11591,N_2213,N_754);
nand U11592 (N_11592,N_2705,N_4058);
nor U11593 (N_11593,N_2543,N_2953);
and U11594 (N_11594,N_4452,N_4695);
nand U11595 (N_11595,N_2733,N_2398);
or U11596 (N_11596,N_5572,N_2661);
nor U11597 (N_11597,N_1645,N_5638);
nand U11598 (N_11598,N_2374,N_4387);
xor U11599 (N_11599,N_2442,N_562);
xor U11600 (N_11600,N_3847,N_3373);
nand U11601 (N_11601,N_2000,N_3265);
nor U11602 (N_11602,N_2978,N_5579);
nand U11603 (N_11603,N_1708,N_2614);
nor U11604 (N_11604,N_3807,N_570);
and U11605 (N_11605,N_3151,N_557);
nand U11606 (N_11606,N_4487,N_310);
nor U11607 (N_11607,N_4948,N_3059);
and U11608 (N_11608,N_869,N_2289);
xor U11609 (N_11609,N_2796,N_1714);
xnor U11610 (N_11610,N_4806,N_2266);
and U11611 (N_11611,N_1910,N_2236);
nor U11612 (N_11612,N_3439,N_5610);
xor U11613 (N_11613,N_1299,N_2658);
or U11614 (N_11614,N_4875,N_3188);
and U11615 (N_11615,N_4919,N_4185);
nor U11616 (N_11616,N_596,N_1070);
nor U11617 (N_11617,N_3623,N_4632);
and U11618 (N_11618,N_3017,N_4520);
nor U11619 (N_11619,N_1468,N_2155);
and U11620 (N_11620,N_3255,N_5812);
xnor U11621 (N_11621,N_4022,N_605);
xnor U11622 (N_11622,N_4098,N_3281);
nand U11623 (N_11623,N_1457,N_456);
nor U11624 (N_11624,N_203,N_1404);
or U11625 (N_11625,N_454,N_1666);
and U11626 (N_11626,N_4088,N_776);
nand U11627 (N_11627,N_5946,N_2838);
xnor U11628 (N_11628,N_1061,N_1287);
xor U11629 (N_11629,N_5069,N_250);
and U11630 (N_11630,N_3233,N_850);
nor U11631 (N_11631,N_626,N_5152);
or U11632 (N_11632,N_5365,N_2881);
and U11633 (N_11633,N_176,N_1239);
nand U11634 (N_11634,N_2103,N_3865);
nor U11635 (N_11635,N_2958,N_5658);
nor U11636 (N_11636,N_2835,N_1119);
nor U11637 (N_11637,N_5512,N_3886);
or U11638 (N_11638,N_4151,N_5955);
nand U11639 (N_11639,N_154,N_1132);
nor U11640 (N_11640,N_71,N_252);
nor U11641 (N_11641,N_1602,N_5609);
xor U11642 (N_11642,N_5578,N_566);
or U11643 (N_11643,N_2580,N_1706);
and U11644 (N_11644,N_4162,N_3371);
nor U11645 (N_11645,N_176,N_367);
nand U11646 (N_11646,N_4170,N_3539);
and U11647 (N_11647,N_4128,N_185);
nor U11648 (N_11648,N_4204,N_4935);
nor U11649 (N_11649,N_5871,N_2533);
xnor U11650 (N_11650,N_4498,N_2923);
nand U11651 (N_11651,N_4464,N_3169);
xnor U11652 (N_11652,N_1269,N_5077);
or U11653 (N_11653,N_473,N_3443);
nor U11654 (N_11654,N_268,N_5933);
or U11655 (N_11655,N_2605,N_2971);
nor U11656 (N_11656,N_2672,N_1455);
nor U11657 (N_11657,N_4059,N_3237);
and U11658 (N_11658,N_5789,N_1830);
or U11659 (N_11659,N_3935,N_5235);
xor U11660 (N_11660,N_3469,N_1349);
or U11661 (N_11661,N_2286,N_3269);
nor U11662 (N_11662,N_4808,N_5440);
and U11663 (N_11663,N_2453,N_2783);
and U11664 (N_11664,N_5859,N_5417);
nand U11665 (N_11665,N_43,N_4669);
nand U11666 (N_11666,N_5036,N_3980);
or U11667 (N_11667,N_5620,N_5320);
or U11668 (N_11668,N_2937,N_4092);
nand U11669 (N_11669,N_3996,N_4257);
nor U11670 (N_11670,N_239,N_1040);
nand U11671 (N_11671,N_5093,N_1439);
nand U11672 (N_11672,N_2733,N_3822);
nor U11673 (N_11673,N_3132,N_4047);
xor U11674 (N_11674,N_31,N_205);
or U11675 (N_11675,N_203,N_3276);
or U11676 (N_11676,N_3202,N_2143);
nand U11677 (N_11677,N_370,N_3915);
nand U11678 (N_11678,N_4371,N_2737);
and U11679 (N_11679,N_5906,N_2499);
xnor U11680 (N_11680,N_4575,N_4477);
nor U11681 (N_11681,N_2394,N_5989);
or U11682 (N_11682,N_3374,N_399);
nand U11683 (N_11683,N_1064,N_1382);
xnor U11684 (N_11684,N_3375,N_1882);
or U11685 (N_11685,N_3850,N_3288);
and U11686 (N_11686,N_304,N_4353);
xor U11687 (N_11687,N_465,N_2044);
or U11688 (N_11688,N_1499,N_1966);
and U11689 (N_11689,N_5357,N_4249);
nor U11690 (N_11690,N_2,N_4175);
and U11691 (N_11691,N_2555,N_5089);
xor U11692 (N_11692,N_125,N_4338);
nor U11693 (N_11693,N_1871,N_5402);
nor U11694 (N_11694,N_713,N_3853);
xor U11695 (N_11695,N_6,N_492);
xor U11696 (N_11696,N_3229,N_2135);
nor U11697 (N_11697,N_4976,N_933);
and U11698 (N_11698,N_3451,N_4451);
and U11699 (N_11699,N_5169,N_3434);
nor U11700 (N_11700,N_2581,N_4738);
nor U11701 (N_11701,N_4522,N_5623);
nor U11702 (N_11702,N_3711,N_983);
and U11703 (N_11703,N_440,N_2333);
nand U11704 (N_11704,N_2718,N_334);
nor U11705 (N_11705,N_3963,N_5604);
xnor U11706 (N_11706,N_4474,N_603);
nor U11707 (N_11707,N_4206,N_975);
or U11708 (N_11708,N_2355,N_628);
xor U11709 (N_11709,N_1040,N_5420);
nor U11710 (N_11710,N_1955,N_5779);
nor U11711 (N_11711,N_5328,N_3913);
nor U11712 (N_11712,N_5077,N_1949);
xor U11713 (N_11713,N_4107,N_3277);
or U11714 (N_11714,N_3488,N_5396);
or U11715 (N_11715,N_5669,N_1902);
nand U11716 (N_11716,N_2970,N_3882);
nor U11717 (N_11717,N_2898,N_3924);
and U11718 (N_11718,N_1644,N_1276);
nor U11719 (N_11719,N_4005,N_5452);
and U11720 (N_11720,N_3497,N_3769);
nand U11721 (N_11721,N_5363,N_5045);
xnor U11722 (N_11722,N_2016,N_5499);
xor U11723 (N_11723,N_4232,N_4875);
nand U11724 (N_11724,N_5881,N_1434);
nor U11725 (N_11725,N_3959,N_3671);
and U11726 (N_11726,N_1485,N_263);
xnor U11727 (N_11727,N_3160,N_5179);
xnor U11728 (N_11728,N_4522,N_2649);
xnor U11729 (N_11729,N_4033,N_2665);
nor U11730 (N_11730,N_3154,N_112);
and U11731 (N_11731,N_2398,N_2711);
nor U11732 (N_11732,N_3425,N_714);
and U11733 (N_11733,N_3143,N_796);
nor U11734 (N_11734,N_2037,N_2017);
nand U11735 (N_11735,N_2758,N_3);
and U11736 (N_11736,N_646,N_1936);
nand U11737 (N_11737,N_2921,N_3712);
xor U11738 (N_11738,N_246,N_1272);
xor U11739 (N_11739,N_768,N_5060);
or U11740 (N_11740,N_5584,N_707);
and U11741 (N_11741,N_3816,N_47);
or U11742 (N_11742,N_2590,N_67);
or U11743 (N_11743,N_2204,N_3536);
xor U11744 (N_11744,N_728,N_3128);
nand U11745 (N_11745,N_182,N_5961);
nand U11746 (N_11746,N_5560,N_242);
nand U11747 (N_11747,N_3214,N_5705);
nand U11748 (N_11748,N_4513,N_3688);
xor U11749 (N_11749,N_706,N_755);
nor U11750 (N_11750,N_5606,N_1783);
or U11751 (N_11751,N_5410,N_3647);
and U11752 (N_11752,N_294,N_3597);
nor U11753 (N_11753,N_2791,N_2560);
nand U11754 (N_11754,N_2486,N_1511);
nor U11755 (N_11755,N_1051,N_3096);
and U11756 (N_11756,N_3537,N_2627);
nand U11757 (N_11757,N_2426,N_5229);
or U11758 (N_11758,N_4935,N_3594);
or U11759 (N_11759,N_5209,N_3459);
nand U11760 (N_11760,N_3383,N_2555);
xor U11761 (N_11761,N_2044,N_3384);
or U11762 (N_11762,N_1268,N_3656);
nand U11763 (N_11763,N_3199,N_3269);
nand U11764 (N_11764,N_1735,N_2392);
xor U11765 (N_11765,N_5631,N_852);
or U11766 (N_11766,N_1124,N_3574);
and U11767 (N_11767,N_5901,N_1221);
or U11768 (N_11768,N_1750,N_2496);
or U11769 (N_11769,N_3280,N_3151);
nand U11770 (N_11770,N_5790,N_5600);
or U11771 (N_11771,N_1401,N_5779);
or U11772 (N_11772,N_4664,N_5816);
or U11773 (N_11773,N_2608,N_4952);
nand U11774 (N_11774,N_4305,N_4012);
nor U11775 (N_11775,N_1518,N_761);
nor U11776 (N_11776,N_3155,N_2243);
and U11777 (N_11777,N_2144,N_1140);
nand U11778 (N_11778,N_5542,N_1399);
and U11779 (N_11779,N_3730,N_4722);
or U11780 (N_11780,N_690,N_1153);
nor U11781 (N_11781,N_2403,N_5247);
and U11782 (N_11782,N_25,N_4761);
nor U11783 (N_11783,N_5600,N_1284);
or U11784 (N_11784,N_5242,N_5827);
nor U11785 (N_11785,N_1715,N_2003);
and U11786 (N_11786,N_2194,N_2721);
and U11787 (N_11787,N_867,N_1730);
and U11788 (N_11788,N_1221,N_5453);
nand U11789 (N_11789,N_2327,N_4591);
xor U11790 (N_11790,N_5479,N_2303);
nand U11791 (N_11791,N_4614,N_2494);
and U11792 (N_11792,N_1212,N_5932);
xor U11793 (N_11793,N_175,N_3354);
nor U11794 (N_11794,N_2219,N_5608);
and U11795 (N_11795,N_2801,N_3740);
nand U11796 (N_11796,N_1765,N_5363);
and U11797 (N_11797,N_3282,N_2973);
nor U11798 (N_11798,N_2873,N_610);
and U11799 (N_11799,N_97,N_4177);
nor U11800 (N_11800,N_1183,N_5349);
xor U11801 (N_11801,N_143,N_2659);
or U11802 (N_11802,N_3275,N_3948);
or U11803 (N_11803,N_5717,N_1748);
or U11804 (N_11804,N_3644,N_5822);
nand U11805 (N_11805,N_2865,N_1860);
nand U11806 (N_11806,N_2117,N_1602);
or U11807 (N_11807,N_788,N_1029);
xor U11808 (N_11808,N_3145,N_1641);
nand U11809 (N_11809,N_701,N_3352);
xnor U11810 (N_11810,N_3778,N_499);
or U11811 (N_11811,N_2218,N_3690);
xnor U11812 (N_11812,N_3434,N_4815);
and U11813 (N_11813,N_2894,N_1356);
nor U11814 (N_11814,N_5889,N_4265);
and U11815 (N_11815,N_5855,N_56);
and U11816 (N_11816,N_4157,N_5544);
or U11817 (N_11817,N_5062,N_4135);
nor U11818 (N_11818,N_1721,N_5194);
nor U11819 (N_11819,N_5628,N_4110);
or U11820 (N_11820,N_3377,N_1623);
or U11821 (N_11821,N_740,N_5566);
nor U11822 (N_11822,N_2850,N_2144);
xor U11823 (N_11823,N_5557,N_4623);
nor U11824 (N_11824,N_3567,N_4279);
or U11825 (N_11825,N_2636,N_374);
nand U11826 (N_11826,N_315,N_1981);
xnor U11827 (N_11827,N_4557,N_3967);
nand U11828 (N_11828,N_4754,N_3339);
xor U11829 (N_11829,N_5110,N_4790);
xnor U11830 (N_11830,N_5685,N_3633);
nand U11831 (N_11831,N_1346,N_1791);
and U11832 (N_11832,N_5364,N_4348);
or U11833 (N_11833,N_598,N_3041);
and U11834 (N_11834,N_1049,N_522);
xnor U11835 (N_11835,N_4588,N_1112);
or U11836 (N_11836,N_2050,N_4813);
xnor U11837 (N_11837,N_3850,N_1411);
nor U11838 (N_11838,N_1783,N_4426);
nand U11839 (N_11839,N_1235,N_3750);
or U11840 (N_11840,N_3607,N_4596);
nand U11841 (N_11841,N_4848,N_399);
xor U11842 (N_11842,N_3831,N_3179);
nand U11843 (N_11843,N_4021,N_3154);
or U11844 (N_11844,N_4653,N_3438);
xnor U11845 (N_11845,N_4284,N_5157);
nand U11846 (N_11846,N_3960,N_552);
or U11847 (N_11847,N_3388,N_127);
xnor U11848 (N_11848,N_1449,N_4833);
nand U11849 (N_11849,N_3513,N_3047);
or U11850 (N_11850,N_387,N_1135);
or U11851 (N_11851,N_2599,N_3371);
xor U11852 (N_11852,N_5546,N_5241);
nor U11853 (N_11853,N_823,N_4951);
nand U11854 (N_11854,N_1718,N_2030);
or U11855 (N_11855,N_1104,N_5086);
and U11856 (N_11856,N_4039,N_5071);
and U11857 (N_11857,N_1684,N_5898);
nand U11858 (N_11858,N_3327,N_2874);
nand U11859 (N_11859,N_441,N_5591);
nor U11860 (N_11860,N_3446,N_5160);
nor U11861 (N_11861,N_1743,N_1122);
nor U11862 (N_11862,N_3095,N_4027);
nor U11863 (N_11863,N_1815,N_3212);
xor U11864 (N_11864,N_4119,N_2108);
nand U11865 (N_11865,N_413,N_2082);
nor U11866 (N_11866,N_4727,N_1056);
xor U11867 (N_11867,N_5539,N_2041);
and U11868 (N_11868,N_2794,N_1099);
nor U11869 (N_11869,N_5572,N_4187);
nor U11870 (N_11870,N_1168,N_5162);
and U11871 (N_11871,N_4428,N_2243);
xor U11872 (N_11872,N_552,N_5047);
and U11873 (N_11873,N_4024,N_3118);
nand U11874 (N_11874,N_2804,N_4397);
nand U11875 (N_11875,N_5875,N_1211);
nor U11876 (N_11876,N_3911,N_5697);
xor U11877 (N_11877,N_4818,N_1190);
nor U11878 (N_11878,N_3556,N_3213);
nor U11879 (N_11879,N_2527,N_2516);
or U11880 (N_11880,N_5023,N_4526);
and U11881 (N_11881,N_4850,N_5170);
nor U11882 (N_11882,N_5806,N_2704);
nand U11883 (N_11883,N_4413,N_4493);
or U11884 (N_11884,N_5934,N_5696);
nor U11885 (N_11885,N_4303,N_3965);
xor U11886 (N_11886,N_3852,N_2474);
nor U11887 (N_11887,N_356,N_2665);
and U11888 (N_11888,N_2439,N_2272);
or U11889 (N_11889,N_4615,N_4878);
or U11890 (N_11890,N_3071,N_4967);
and U11891 (N_11891,N_1366,N_1355);
or U11892 (N_11892,N_4184,N_2210);
or U11893 (N_11893,N_2678,N_2100);
xor U11894 (N_11894,N_5255,N_1775);
or U11895 (N_11895,N_5428,N_3333);
nand U11896 (N_11896,N_1419,N_787);
or U11897 (N_11897,N_4904,N_1764);
or U11898 (N_11898,N_2550,N_5270);
nor U11899 (N_11899,N_4107,N_3333);
or U11900 (N_11900,N_3908,N_3722);
nand U11901 (N_11901,N_1895,N_4416);
nand U11902 (N_11902,N_1125,N_2919);
xor U11903 (N_11903,N_4666,N_762);
nand U11904 (N_11904,N_4285,N_1693);
xnor U11905 (N_11905,N_4873,N_5941);
nand U11906 (N_11906,N_1333,N_1216);
and U11907 (N_11907,N_4976,N_5538);
and U11908 (N_11908,N_1798,N_429);
and U11909 (N_11909,N_3659,N_2103);
and U11910 (N_11910,N_5827,N_5485);
or U11911 (N_11911,N_4641,N_920);
nor U11912 (N_11912,N_2566,N_713);
and U11913 (N_11913,N_5499,N_4414);
or U11914 (N_11914,N_2081,N_1874);
xnor U11915 (N_11915,N_5130,N_2124);
and U11916 (N_11916,N_1221,N_731);
or U11917 (N_11917,N_3939,N_4366);
nor U11918 (N_11918,N_5584,N_2972);
nor U11919 (N_11919,N_3659,N_1327);
nor U11920 (N_11920,N_2774,N_1223);
nor U11921 (N_11921,N_581,N_3367);
nor U11922 (N_11922,N_271,N_3678);
nor U11923 (N_11923,N_329,N_1292);
nor U11924 (N_11924,N_5508,N_3662);
nor U11925 (N_11925,N_3504,N_2030);
xnor U11926 (N_11926,N_2945,N_3775);
nor U11927 (N_11927,N_1445,N_3323);
nor U11928 (N_11928,N_3199,N_5873);
or U11929 (N_11929,N_1496,N_4532);
nor U11930 (N_11930,N_305,N_4291);
or U11931 (N_11931,N_1871,N_2971);
and U11932 (N_11932,N_207,N_3316);
nand U11933 (N_11933,N_5514,N_742);
xor U11934 (N_11934,N_1605,N_760);
or U11935 (N_11935,N_1566,N_2320);
xor U11936 (N_11936,N_4905,N_5158);
xor U11937 (N_11937,N_3243,N_171);
nand U11938 (N_11938,N_3254,N_3876);
nand U11939 (N_11939,N_1474,N_986);
nor U11940 (N_11940,N_5428,N_3543);
or U11941 (N_11941,N_5282,N_2139);
and U11942 (N_11942,N_3492,N_2581);
nor U11943 (N_11943,N_700,N_1548);
xnor U11944 (N_11944,N_4529,N_5556);
xor U11945 (N_11945,N_3603,N_2279);
and U11946 (N_11946,N_2521,N_4394);
nor U11947 (N_11947,N_2845,N_1356);
nor U11948 (N_11948,N_5779,N_4799);
and U11949 (N_11949,N_3447,N_2136);
nor U11950 (N_11950,N_1585,N_5019);
and U11951 (N_11951,N_4183,N_2917);
and U11952 (N_11952,N_292,N_2606);
nand U11953 (N_11953,N_2211,N_3451);
nor U11954 (N_11954,N_3081,N_2975);
nand U11955 (N_11955,N_1352,N_754);
and U11956 (N_11956,N_215,N_4008);
xor U11957 (N_11957,N_3744,N_3356);
and U11958 (N_11958,N_622,N_5433);
nand U11959 (N_11959,N_5015,N_1318);
xor U11960 (N_11960,N_1969,N_3398);
or U11961 (N_11961,N_5634,N_494);
and U11962 (N_11962,N_71,N_2564);
nand U11963 (N_11963,N_3138,N_716);
and U11964 (N_11964,N_5192,N_5343);
xnor U11965 (N_11965,N_1502,N_1999);
nor U11966 (N_11966,N_5074,N_4630);
xor U11967 (N_11967,N_2994,N_5901);
xor U11968 (N_11968,N_1261,N_3310);
and U11969 (N_11969,N_1675,N_3110);
nand U11970 (N_11970,N_829,N_4686);
nand U11971 (N_11971,N_0,N_3474);
xor U11972 (N_11972,N_3610,N_2360);
or U11973 (N_11973,N_5438,N_833);
or U11974 (N_11974,N_1556,N_2155);
and U11975 (N_11975,N_1800,N_3704);
nand U11976 (N_11976,N_5625,N_1626);
or U11977 (N_11977,N_3621,N_5234);
and U11978 (N_11978,N_2886,N_2992);
xor U11979 (N_11979,N_3796,N_2050);
xnor U11980 (N_11980,N_1802,N_4968);
xnor U11981 (N_11981,N_3564,N_5930);
and U11982 (N_11982,N_5243,N_5592);
or U11983 (N_11983,N_4935,N_3411);
nand U11984 (N_11984,N_499,N_865);
or U11985 (N_11985,N_5896,N_575);
or U11986 (N_11986,N_3002,N_5099);
xor U11987 (N_11987,N_5529,N_1772);
or U11988 (N_11988,N_2190,N_4065);
nor U11989 (N_11989,N_1251,N_983);
nor U11990 (N_11990,N_670,N_2249);
xor U11991 (N_11991,N_1655,N_348);
or U11992 (N_11992,N_996,N_806);
nand U11993 (N_11993,N_948,N_1470);
xor U11994 (N_11994,N_2395,N_3794);
xor U11995 (N_11995,N_1261,N_850);
nand U11996 (N_11996,N_5756,N_3060);
xnor U11997 (N_11997,N_203,N_4556);
and U11998 (N_11998,N_3793,N_4032);
nand U11999 (N_11999,N_2877,N_3983);
xor U12000 (N_12000,N_9309,N_6028);
or U12001 (N_12001,N_10982,N_8392);
nand U12002 (N_12002,N_6846,N_10320);
nand U12003 (N_12003,N_7470,N_8140);
xnor U12004 (N_12004,N_9322,N_10240);
or U12005 (N_12005,N_8966,N_6822);
nand U12006 (N_12006,N_7851,N_8930);
nor U12007 (N_12007,N_10416,N_10991);
xor U12008 (N_12008,N_6197,N_7323);
nor U12009 (N_12009,N_9068,N_10015);
and U12010 (N_12010,N_8288,N_10010);
or U12011 (N_12011,N_10467,N_6411);
and U12012 (N_12012,N_10619,N_9952);
nand U12013 (N_12013,N_8276,N_7254);
nand U12014 (N_12014,N_8393,N_11777);
or U12015 (N_12015,N_11075,N_6838);
and U12016 (N_12016,N_6778,N_7177);
nand U12017 (N_12017,N_10544,N_11570);
xnor U12018 (N_12018,N_6633,N_11686);
or U12019 (N_12019,N_8285,N_10279);
xor U12020 (N_12020,N_9125,N_7726);
nand U12021 (N_12021,N_11244,N_7795);
and U12022 (N_12022,N_8368,N_8274);
nor U12023 (N_12023,N_9311,N_7576);
and U12024 (N_12024,N_6693,N_11938);
nor U12025 (N_12025,N_11859,N_6119);
and U12026 (N_12026,N_11062,N_8204);
xor U12027 (N_12027,N_11980,N_9145);
nand U12028 (N_12028,N_9821,N_6319);
nand U12029 (N_12029,N_9875,N_11093);
or U12030 (N_12030,N_6163,N_9728);
xnor U12031 (N_12031,N_9743,N_8499);
or U12032 (N_12032,N_10996,N_7515);
or U12033 (N_12033,N_7644,N_11065);
xnor U12034 (N_12034,N_8672,N_6211);
or U12035 (N_12035,N_9308,N_9293);
or U12036 (N_12036,N_8637,N_11469);
or U12037 (N_12037,N_6338,N_7161);
nand U12038 (N_12038,N_7958,N_8382);
xnor U12039 (N_12039,N_7762,N_11308);
or U12040 (N_12040,N_10235,N_8987);
nand U12041 (N_12041,N_7180,N_11698);
nand U12042 (N_12042,N_7174,N_10345);
xor U12043 (N_12043,N_9557,N_9462);
xor U12044 (N_12044,N_11241,N_7780);
or U12045 (N_12045,N_7892,N_7568);
nor U12046 (N_12046,N_9953,N_7335);
or U12047 (N_12047,N_9035,N_8024);
nand U12048 (N_12048,N_6106,N_9285);
nor U12049 (N_12049,N_6614,N_8051);
nor U12050 (N_12050,N_8559,N_8686);
nor U12051 (N_12051,N_9710,N_6386);
or U12052 (N_12052,N_10084,N_8365);
nand U12053 (N_12053,N_11431,N_7261);
nand U12054 (N_12054,N_7998,N_6514);
or U12055 (N_12055,N_8826,N_8073);
nor U12056 (N_12056,N_9027,N_7328);
nor U12057 (N_12057,N_6388,N_6468);
xnor U12058 (N_12058,N_11547,N_6117);
and U12059 (N_12059,N_8876,N_6737);
nor U12060 (N_12060,N_9493,N_11406);
nand U12061 (N_12061,N_6036,N_7149);
nand U12062 (N_12062,N_6967,N_6749);
xnor U12063 (N_12063,N_7961,N_10876);
and U12064 (N_12064,N_7582,N_9836);
xor U12065 (N_12065,N_7759,N_9990);
nor U12066 (N_12066,N_11739,N_8287);
and U12067 (N_12067,N_7603,N_7252);
xnor U12068 (N_12068,N_8718,N_7210);
and U12069 (N_12069,N_11650,N_9809);
and U12070 (N_12070,N_11567,N_6894);
nand U12071 (N_12071,N_10228,N_6055);
nand U12072 (N_12072,N_11902,N_9296);
xnor U12073 (N_12073,N_10119,N_7037);
nand U12074 (N_12074,N_8237,N_10064);
nor U12075 (N_12075,N_6499,N_6453);
nor U12076 (N_12076,N_7807,N_6698);
nand U12077 (N_12077,N_7977,N_9519);
nand U12078 (N_12078,N_9238,N_8350);
or U12079 (N_12079,N_9741,N_8048);
nor U12080 (N_12080,N_7012,N_11633);
nand U12081 (N_12081,N_8451,N_8246);
or U12082 (N_12082,N_11656,N_7999);
xnor U12083 (N_12083,N_9759,N_8157);
or U12084 (N_12084,N_7855,N_7553);
xnor U12085 (N_12085,N_8896,N_8667);
or U12086 (N_12086,N_6017,N_8309);
xnor U12087 (N_12087,N_9352,N_7638);
xor U12088 (N_12088,N_11729,N_10535);
xor U12089 (N_12089,N_9856,N_10966);
and U12090 (N_12090,N_7092,N_7309);
nand U12091 (N_12091,N_10024,N_10198);
nand U12092 (N_12092,N_10040,N_10417);
nor U12093 (N_12093,N_6060,N_11235);
nor U12094 (N_12094,N_7287,N_9892);
xnor U12095 (N_12095,N_8016,N_8317);
nor U12096 (N_12096,N_8115,N_6566);
nand U12097 (N_12097,N_10212,N_10486);
nor U12098 (N_12098,N_11367,N_6362);
nor U12099 (N_12099,N_11850,N_6255);
and U12100 (N_12100,N_7134,N_6137);
xor U12101 (N_12101,N_9297,N_6734);
nor U12102 (N_12102,N_6038,N_10833);
or U12103 (N_12103,N_9294,N_6702);
or U12104 (N_12104,N_9957,N_8214);
nand U12105 (N_12105,N_9961,N_7670);
and U12106 (N_12106,N_8364,N_10887);
or U12107 (N_12107,N_11008,N_11087);
xnor U12108 (N_12108,N_10711,N_11792);
nor U12109 (N_12109,N_10348,N_11935);
nand U12110 (N_12110,N_7525,N_9969);
and U12111 (N_12111,N_10420,N_11309);
and U12112 (N_12112,N_7333,N_7268);
nor U12113 (N_12113,N_8687,N_11179);
xor U12114 (N_12114,N_11021,N_9355);
or U12115 (N_12115,N_7725,N_6023);
or U12116 (N_12116,N_7981,N_6571);
nor U12117 (N_12117,N_8770,N_10315);
nand U12118 (N_12118,N_10761,N_10894);
and U12119 (N_12119,N_6853,N_6562);
nor U12120 (N_12120,N_11694,N_8370);
or U12121 (N_12121,N_6673,N_9508);
nand U12122 (N_12122,N_11027,N_8516);
xor U12123 (N_12123,N_9200,N_11425);
xor U12124 (N_12124,N_7572,N_10495);
nand U12125 (N_12125,N_9636,N_7565);
nand U12126 (N_12126,N_6650,N_9602);
or U12127 (N_12127,N_10503,N_7659);
xor U12128 (N_12128,N_6477,N_7789);
nand U12129 (N_12129,N_11976,N_8971);
nand U12130 (N_12130,N_9552,N_10551);
nor U12131 (N_12131,N_8359,N_9419);
nor U12132 (N_12132,N_9469,N_9380);
and U12133 (N_12133,N_11899,N_8592);
nor U12134 (N_12134,N_8928,N_11505);
and U12135 (N_12135,N_6597,N_6294);
nor U12136 (N_12136,N_8063,N_11394);
xnor U12137 (N_12137,N_9737,N_6088);
nor U12138 (N_12138,N_8217,N_10190);
xnor U12139 (N_12139,N_11875,N_8720);
xor U12140 (N_12140,N_10293,N_7089);
nand U12141 (N_12141,N_11722,N_6905);
nor U12142 (N_12142,N_10915,N_11143);
xnor U12143 (N_12143,N_9154,N_9371);
and U12144 (N_12144,N_7269,N_7158);
nor U12145 (N_12145,N_6553,N_10643);
nand U12146 (N_12146,N_10984,N_11148);
nand U12147 (N_12147,N_10221,N_9719);
nand U12148 (N_12148,N_11231,N_8429);
nor U12149 (N_12149,N_7011,N_9008);
nand U12150 (N_12150,N_8877,N_11006);
nor U12151 (N_12151,N_11229,N_6156);
nor U12152 (N_12152,N_9692,N_8447);
or U12153 (N_12153,N_9024,N_10831);
nand U12154 (N_12154,N_10045,N_8746);
or U12155 (N_12155,N_7152,N_9253);
and U12156 (N_12156,N_11689,N_8735);
nor U12157 (N_12157,N_9264,N_10772);
and U12158 (N_12158,N_9686,N_11287);
nand U12159 (N_12159,N_10821,N_7802);
or U12160 (N_12160,N_10776,N_7581);
nor U12161 (N_12161,N_9687,N_11282);
or U12162 (N_12162,N_7523,N_10216);
nand U12163 (N_12163,N_11374,N_10395);
nor U12164 (N_12164,N_6596,N_9825);
nand U12165 (N_12165,N_11818,N_10004);
xnor U12166 (N_12166,N_9223,N_10926);
and U12167 (N_12167,N_11019,N_8294);
nor U12168 (N_12168,N_7772,N_11207);
xor U12169 (N_12169,N_8940,N_6665);
nand U12170 (N_12170,N_10734,N_10434);
or U12171 (N_12171,N_8553,N_8523);
nand U12172 (N_12172,N_7989,N_7562);
nand U12173 (N_12173,N_9472,N_10871);
or U12174 (N_12174,N_7103,N_6236);
nand U12175 (N_12175,N_10514,N_8467);
and U12176 (N_12176,N_10581,N_7895);
nor U12177 (N_12177,N_9029,N_10205);
nor U12178 (N_12178,N_11740,N_10444);
nand U12179 (N_12179,N_7372,N_6725);
nor U12180 (N_12180,N_7862,N_8114);
nor U12181 (N_12181,N_6136,N_7060);
nand U12182 (N_12182,N_9205,N_9249);
xor U12183 (N_12183,N_9321,N_10903);
nor U12184 (N_12184,N_10593,N_10510);
nand U12185 (N_12185,N_11795,N_7052);
xnor U12186 (N_12186,N_9639,N_10272);
or U12187 (N_12187,N_9921,N_6173);
xor U12188 (N_12188,N_6227,N_10282);
xor U12189 (N_12189,N_10671,N_8760);
nand U12190 (N_12190,N_6050,N_9604);
and U12191 (N_12191,N_9305,N_8052);
and U12192 (N_12192,N_7188,N_7779);
and U12193 (N_12193,N_10431,N_11528);
nor U12194 (N_12194,N_11154,N_9659);
or U12195 (N_12195,N_7547,N_10223);
nor U12196 (N_12196,N_10708,N_6828);
or U12197 (N_12197,N_11054,N_8040);
or U12198 (N_12198,N_7241,N_9358);
nand U12199 (N_12199,N_11058,N_9509);
or U12200 (N_12200,N_6341,N_8604);
and U12201 (N_12201,N_6416,N_10307);
nand U12202 (N_12202,N_8319,N_10407);
and U12203 (N_12203,N_8381,N_11300);
nor U12204 (N_12204,N_10238,N_6953);
nand U12205 (N_12205,N_11360,N_11415);
nor U12206 (N_12206,N_8191,N_6825);
nor U12207 (N_12207,N_6950,N_10536);
nand U12208 (N_12208,N_8064,N_9624);
nand U12209 (N_12209,N_11680,N_11713);
and U12210 (N_12210,N_9266,N_11095);
nor U12211 (N_12211,N_8195,N_9181);
and U12212 (N_12212,N_8180,N_6234);
or U12213 (N_12213,N_7633,N_11471);
nor U12214 (N_12214,N_9229,N_8417);
or U12215 (N_12215,N_11820,N_10846);
and U12216 (N_12216,N_10430,N_10249);
nand U12217 (N_12217,N_7048,N_11166);
or U12218 (N_12218,N_7681,N_10867);
or U12219 (N_12219,N_7208,N_7426);
and U12220 (N_12220,N_8894,N_7368);
nand U12221 (N_12221,N_6105,N_7081);
and U12222 (N_12222,N_10726,N_6839);
nor U12223 (N_12223,N_6307,N_7415);
and U12224 (N_12224,N_9009,N_8038);
xor U12225 (N_12225,N_7641,N_6048);
and U12226 (N_12226,N_7348,N_6576);
nand U12227 (N_12227,N_6854,N_9722);
or U12228 (N_12228,N_8128,N_7667);
xnor U12229 (N_12229,N_10397,N_11466);
nand U12230 (N_12230,N_11884,N_6422);
xnor U12231 (N_12231,N_11801,N_7956);
or U12232 (N_12232,N_7677,N_11053);
or U12233 (N_12233,N_7917,N_7247);
nand U12234 (N_12234,N_6719,N_7908);
and U12235 (N_12235,N_6146,N_9320);
xor U12236 (N_12236,N_10729,N_10563);
or U12237 (N_12237,N_8378,N_7800);
or U12238 (N_12238,N_9174,N_7545);
and U12239 (N_12239,N_6071,N_6465);
or U12240 (N_12240,N_9511,N_10875);
nor U12241 (N_12241,N_6252,N_8841);
and U12242 (N_12242,N_9863,N_7440);
or U12243 (N_12243,N_6029,N_7144);
or U12244 (N_12244,N_10693,N_11163);
or U12245 (N_12245,N_7450,N_11091);
xor U12246 (N_12246,N_6241,N_9279);
or U12247 (N_12247,N_6426,N_10384);
xor U12248 (N_12248,N_10487,N_10934);
and U12249 (N_12249,N_11504,N_11910);
nand U12250 (N_12250,N_10341,N_8278);
and U12251 (N_12251,N_7173,N_10394);
or U12252 (N_12252,N_9663,N_10418);
or U12253 (N_12253,N_8037,N_6686);
nor U12254 (N_12254,N_9789,N_6887);
and U12255 (N_12255,N_11584,N_6796);
nor U12256 (N_12256,N_11250,N_9445);
xnor U12257 (N_12257,N_8908,N_9310);
nand U12258 (N_12258,N_6581,N_11653);
nand U12259 (N_12259,N_6744,N_7820);
nand U12260 (N_12260,N_9740,N_8573);
nand U12261 (N_12261,N_6222,N_6543);
or U12262 (N_12262,N_6191,N_11866);
nand U12263 (N_12263,N_9072,N_8673);
and U12264 (N_12264,N_10425,N_7297);
nand U12265 (N_12265,N_8614,N_10808);
xnor U12266 (N_12266,N_6087,N_10891);
or U12267 (N_12267,N_6602,N_11121);
and U12268 (N_12268,N_9324,N_10807);
nor U12269 (N_12269,N_9696,N_7841);
nor U12270 (N_12270,N_8558,N_11554);
or U12271 (N_12271,N_8145,N_6647);
and U12272 (N_12272,N_10362,N_9045);
nand U12273 (N_12273,N_9712,N_6090);
and U12274 (N_12274,N_11495,N_11856);
nand U12275 (N_12275,N_9866,N_7314);
nor U12276 (N_12276,N_8797,N_8514);
xor U12277 (N_12277,N_9993,N_6446);
and U12278 (N_12278,N_8308,N_9669);
or U12279 (N_12279,N_11489,N_8167);
nor U12280 (N_12280,N_6459,N_10342);
xor U12281 (N_12281,N_9411,N_6867);
xor U12282 (N_12282,N_7135,N_10356);
xnor U12283 (N_12283,N_7122,N_6875);
or U12284 (N_12284,N_6215,N_9457);
nor U12285 (N_12285,N_8830,N_9974);
nor U12286 (N_12286,N_11872,N_7794);
and U12287 (N_12287,N_8799,N_8507);
or U12288 (N_12288,N_8983,N_10241);
nand U12289 (N_12289,N_7034,N_10940);
xnor U12290 (N_12290,N_11736,N_6144);
nand U12291 (N_12291,N_6978,N_10476);
nor U12292 (N_12292,N_9448,N_6271);
or U12293 (N_12293,N_6261,N_7773);
and U12294 (N_12294,N_8598,N_9651);
nand U12295 (N_12295,N_11886,N_7155);
xor U12296 (N_12296,N_9456,N_9428);
nand U12297 (N_12297,N_9482,N_10501);
nor U12298 (N_12298,N_9280,N_10368);
nor U12299 (N_12299,N_8622,N_6253);
nor U12300 (N_12300,N_7646,N_6367);
xor U12301 (N_12301,N_8496,N_9106);
or U12302 (N_12302,N_6250,N_9650);
or U12303 (N_12303,N_10043,N_8722);
nand U12304 (N_12304,N_9985,N_9037);
xnor U12305 (N_12305,N_6959,N_10391);
xnor U12306 (N_12306,N_6892,N_9331);
or U12307 (N_12307,N_9343,N_8560);
or U12308 (N_12308,N_9254,N_8478);
nand U12309 (N_12309,N_8252,N_6067);
nor U12310 (N_12310,N_7482,N_9250);
xor U12311 (N_12311,N_8679,N_6845);
nor U12312 (N_12312,N_6681,N_9244);
and U12313 (N_12313,N_7487,N_11369);
nand U12314 (N_12314,N_11128,N_9489);
xnor U12315 (N_12315,N_7987,N_10116);
and U12316 (N_12316,N_9893,N_11092);
and U12317 (N_12317,N_10294,N_9234);
nor U12318 (N_12318,N_8755,N_9175);
nand U12319 (N_12319,N_6640,N_8831);
nand U12320 (N_12320,N_9099,N_8694);
xnor U12321 (N_12321,N_7921,N_9948);
nand U12322 (N_12322,N_9655,N_8234);
nand U12323 (N_12323,N_8374,N_10259);
nor U12324 (N_12324,N_6970,N_10860);
and U12325 (N_12325,N_6044,N_8127);
xor U12326 (N_12326,N_7095,N_6405);
nor U12327 (N_12327,N_11966,N_7359);
or U12328 (N_12328,N_7975,N_11683);
and U12329 (N_12329,N_10186,N_7198);
xnor U12330 (N_12330,N_6954,N_6193);
or U12331 (N_12331,N_8203,N_11613);
nand U12332 (N_12332,N_6573,N_9590);
and U12333 (N_12333,N_8783,N_10965);
and U12334 (N_12334,N_7010,N_10817);
and U12335 (N_12335,N_9461,N_7853);
and U12336 (N_12336,N_7821,N_10660);
and U12337 (N_12337,N_11617,N_9078);
xor U12338 (N_12338,N_9513,N_11212);
nand U12339 (N_12339,N_10373,N_6040);
xor U12340 (N_12340,N_10976,N_7175);
nand U12341 (N_12341,N_8091,N_10106);
xnor U12342 (N_12342,N_11518,N_10463);
nand U12343 (N_12343,N_10367,N_8898);
nor U12344 (N_12344,N_6366,N_6893);
and U12345 (N_12345,N_8583,N_8386);
nor U12346 (N_12346,N_6728,N_7716);
xor U12347 (N_12347,N_9494,N_9715);
nor U12348 (N_12348,N_10421,N_11100);
nor U12349 (N_12349,N_11751,N_8913);
nand U12350 (N_12350,N_9323,N_6885);
nand U12351 (N_12351,N_8438,N_8771);
or U12352 (N_12352,N_10077,N_7737);
or U12353 (N_12353,N_7317,N_11553);
and U12354 (N_12354,N_8247,N_8501);
and U12355 (N_12355,N_8432,N_6783);
nor U12356 (N_12356,N_8231,N_8973);
nor U12357 (N_12357,N_10958,N_11261);
or U12358 (N_12358,N_7930,N_10554);
xnor U12359 (N_12359,N_11373,N_9017);
nand U12360 (N_12360,N_10771,N_8676);
nor U12361 (N_12361,N_6052,N_11214);
or U12362 (N_12362,N_9882,N_9680);
nor U12363 (N_12363,N_7086,N_10280);
nor U12364 (N_12364,N_11029,N_10677);
or U12365 (N_12365,N_7191,N_10100);
nand U12366 (N_12366,N_6258,N_7085);
or U12367 (N_12367,N_9334,N_6575);
or U12368 (N_12368,N_10225,N_8187);
nand U12369 (N_12369,N_7731,N_10099);
and U12370 (N_12370,N_7625,N_6302);
xnor U12371 (N_12371,N_11182,N_11947);
xnor U12372 (N_12372,N_10881,N_7993);
or U12373 (N_12373,N_10764,N_6946);
xnor U12374 (N_12374,N_6630,N_7850);
or U12375 (N_12375,N_11001,N_9353);
nor U12376 (N_12376,N_10931,N_7898);
nor U12377 (N_12377,N_7684,N_9114);
and U12378 (N_12378,N_8147,N_7929);
nor U12379 (N_12379,N_9299,N_7925);
or U12380 (N_12380,N_8304,N_11486);
nor U12381 (N_12381,N_7439,N_10402);
or U12382 (N_12382,N_8372,N_6788);
or U12383 (N_12383,N_6075,N_7378);
nand U12384 (N_12384,N_8638,N_7982);
xor U12385 (N_12385,N_8915,N_8521);
nor U12386 (N_12386,N_9661,N_7114);
nand U12387 (N_12387,N_10720,N_9278);
nor U12388 (N_12388,N_7270,N_9191);
or U12389 (N_12389,N_6122,N_7612);
nand U12390 (N_12390,N_11814,N_10977);
nor U12391 (N_12391,N_8549,N_10189);
or U12392 (N_12392,N_10951,N_9441);
xnor U12393 (N_12393,N_11366,N_11441);
or U12394 (N_12394,N_6006,N_10067);
xnor U12395 (N_12395,N_6827,N_9386);
or U12396 (N_12396,N_9622,N_8408);
xnor U12397 (N_12397,N_8716,N_7004);
or U12398 (N_12398,N_6579,N_8112);
nor U12399 (N_12399,N_10678,N_10159);
xor U12400 (N_12400,N_9032,N_9613);
or U12401 (N_12401,N_7020,N_7082);
and U12402 (N_12402,N_7922,N_8097);
and U12403 (N_12403,N_9806,N_11601);
nor U12404 (N_12404,N_10478,N_7009);
and U12405 (N_12405,N_11098,N_7057);
or U12406 (N_12406,N_7986,N_8003);
xor U12407 (N_12407,N_9935,N_7810);
or U12408 (N_12408,N_8271,N_7703);
or U12409 (N_12409,N_9786,N_7137);
xor U12410 (N_12410,N_7017,N_10797);
xnor U12411 (N_12411,N_10366,N_11968);
xor U12412 (N_12412,N_8544,N_11672);
nor U12413 (N_12413,N_11152,N_9992);
nor U12414 (N_12414,N_7952,N_6540);
and U12415 (N_12415,N_6490,N_10393);
xor U12416 (N_12416,N_9677,N_7374);
nand U12417 (N_12417,N_8596,N_8852);
or U12418 (N_12418,N_6143,N_11208);
and U12419 (N_12419,N_6114,N_9330);
or U12420 (N_12420,N_11311,N_7529);
nor U12421 (N_12421,N_11833,N_11663);
and U12422 (N_12422,N_9865,N_9698);
nor U12423 (N_12423,N_9130,N_9906);
nand U12424 (N_12424,N_7157,N_11280);
and U12425 (N_12425,N_8343,N_8919);
nor U12426 (N_12426,N_10215,N_10071);
or U12427 (N_12427,N_11749,N_6103);
nor U12428 (N_12428,N_6570,N_7027);
nor U12429 (N_12429,N_11527,N_10630);
nand U12430 (N_12430,N_6132,N_11578);
nand U12431 (N_12431,N_6772,N_11537);
nor U12432 (N_12432,N_7826,N_11953);
nand U12433 (N_12433,N_8658,N_11251);
nor U12434 (N_12434,N_6836,N_10182);
and U12435 (N_12435,N_10781,N_10335);
and U12436 (N_12436,N_6523,N_11009);
nand U12437 (N_12437,N_11523,N_11336);
nand U12438 (N_12438,N_11327,N_9938);
xnor U12439 (N_12439,N_8473,N_10167);
nand U12440 (N_12440,N_7707,N_10684);
xnor U12441 (N_12441,N_7338,N_6634);
nand U12442 (N_12442,N_9733,N_9501);
and U12443 (N_12443,N_11482,N_9559);
or U12444 (N_12444,N_10139,N_9975);
nand U12445 (N_12445,N_11540,N_9173);
nand U12446 (N_12446,N_9435,N_7859);
nor U12447 (N_12447,N_9328,N_6646);
nand U12448 (N_12448,N_6043,N_10308);
xnor U12449 (N_12449,N_7566,N_11370);
xor U12450 (N_12450,N_7894,N_10460);
xnor U12451 (N_12451,N_11422,N_11341);
xor U12452 (N_12452,N_7279,N_6568);
or U12453 (N_12453,N_7920,N_10559);
or U12454 (N_12454,N_9828,N_8741);
xnor U12455 (N_12455,N_11778,N_11183);
or U12456 (N_12456,N_9523,N_11348);
and U12457 (N_12457,N_9372,N_8701);
or U12458 (N_12458,N_8586,N_9256);
xor U12459 (N_12459,N_10137,N_6852);
nand U12460 (N_12460,N_8084,N_8227);
or U12461 (N_12461,N_6181,N_9678);
or U12462 (N_12462,N_10509,N_7281);
xor U12463 (N_12463,N_7615,N_11240);
nand U12464 (N_12464,N_7560,N_10757);
xnor U12465 (N_12465,N_7899,N_8249);
or U12466 (N_12466,N_9220,N_9911);
and U12467 (N_12467,N_6763,N_9030);
and U12468 (N_12468,N_6287,N_8182);
xnor U12469 (N_12469,N_9033,N_8474);
and U12470 (N_12470,N_11108,N_11949);
xor U12471 (N_12471,N_8680,N_11810);
xor U12472 (N_12472,N_8028,N_9754);
and U12473 (N_12473,N_6083,N_7066);
or U12474 (N_12474,N_8787,N_6395);
and U12475 (N_12475,N_11176,N_8179);
nand U12476 (N_12476,N_6432,N_9402);
nor U12477 (N_12477,N_10888,N_8832);
nand U12478 (N_12478,N_7693,N_7331);
or U12479 (N_12479,N_9695,N_8570);
xor U12480 (N_12480,N_8540,N_9356);
and U12481 (N_12481,N_10621,N_8981);
nand U12482 (N_12482,N_8357,N_6175);
or U12483 (N_12483,N_9383,N_6486);
nor U12484 (N_12484,N_9226,N_9413);
nand U12485 (N_12485,N_6670,N_7407);
nor U12486 (N_12486,N_7217,N_7651);
nand U12487 (N_12487,N_6342,N_10230);
nand U12488 (N_12488,N_7361,N_7226);
nand U12489 (N_12489,N_9385,N_7003);
nor U12490 (N_12490,N_8094,N_11526);
and U12491 (N_12491,N_9292,N_11566);
nor U12492 (N_12492,N_10911,N_7029);
xnor U12493 (N_12493,N_7105,N_10747);
xnor U12494 (N_12494,N_9189,N_7221);
xnor U12495 (N_12495,N_10906,N_7765);
nand U12496 (N_12496,N_6424,N_9901);
and U12497 (N_12497,N_10316,N_9079);
or U12498 (N_12498,N_10532,N_7481);
or U12499 (N_12499,N_6168,N_8412);
nand U12500 (N_12500,N_6606,N_9587);
xor U12501 (N_12501,N_7708,N_11799);
or U12502 (N_12502,N_10290,N_7113);
or U12503 (N_12503,N_6935,N_11755);
nor U12504 (N_12504,N_11118,N_11284);
and U12505 (N_12505,N_6390,N_11123);
and U12506 (N_12506,N_10002,N_7065);
or U12507 (N_12507,N_6934,N_6922);
nand U12508 (N_12508,N_11784,N_11853);
and U12509 (N_12509,N_6720,N_7329);
nor U12510 (N_12510,N_6368,N_7369);
or U12511 (N_12511,N_6672,N_6519);
or U12512 (N_12512,N_9543,N_8058);
xnor U12513 (N_12513,N_7750,N_8792);
or U12514 (N_12514,N_9196,N_6653);
xor U12515 (N_12515,N_10375,N_6290);
nor U12516 (N_12516,N_7970,N_6676);
xnor U12517 (N_12517,N_11016,N_9943);
nand U12518 (N_12518,N_11964,N_7377);
nand U12519 (N_12519,N_8230,N_6124);
nor U12520 (N_12520,N_11127,N_10283);
and U12521 (N_12521,N_10331,N_7249);
nor U12522 (N_12522,N_7164,N_9083);
nand U12523 (N_12523,N_9046,N_6986);
xor U12524 (N_12524,N_11496,N_10562);
or U12525 (N_12525,N_9271,N_8520);
xor U12526 (N_12526,N_10739,N_8015);
xor U12527 (N_12527,N_7013,N_7885);
nand U12528 (N_12528,N_7460,N_10859);
or U12529 (N_12529,N_9671,N_9536);
or U12530 (N_12530,N_6102,N_7963);
nor U12531 (N_12531,N_8156,N_9939);
nor U12532 (N_12532,N_9818,N_11948);
nand U12533 (N_12533,N_11137,N_11470);
or U12534 (N_12534,N_7146,N_6108);
and U12535 (N_12535,N_11582,N_7733);
nor U12536 (N_12536,N_7580,N_7237);
nor U12537 (N_12537,N_10448,N_8975);
and U12538 (N_12538,N_11703,N_6595);
and U12539 (N_12539,N_7093,N_6332);
nor U12540 (N_12540,N_6058,N_7123);
or U12541 (N_12541,N_10415,N_6812);
or U12542 (N_12542,N_11660,N_6393);
and U12543 (N_12543,N_6370,N_8618);
or U12544 (N_12544,N_7650,N_10396);
and U12545 (N_12545,N_6675,N_11797);
nor U12546 (N_12546,N_10126,N_6382);
nand U12547 (N_12547,N_8340,N_10768);
nor U12548 (N_12548,N_10756,N_8401);
and U12549 (N_12549,N_8254,N_6092);
nor U12550 (N_12550,N_7245,N_11077);
or U12551 (N_12551,N_9965,N_6361);
and U12552 (N_12552,N_8067,N_9488);
nand U12553 (N_12553,N_10093,N_11864);
nand U12554 (N_12554,N_8910,N_9274);
or U12555 (N_12555,N_10023,N_6207);
and U12556 (N_12556,N_10650,N_8630);
or U12557 (N_12557,N_6564,N_7948);
nand U12558 (N_12558,N_6112,N_6363);
xnor U12559 (N_12559,N_11117,N_11069);
nand U12560 (N_12560,N_10491,N_9013);
xor U12561 (N_12561,N_8212,N_6760);
and U12562 (N_12562,N_10047,N_9764);
or U12563 (N_12563,N_10154,N_6683);
nor U12564 (N_12564,N_11852,N_6260);
nand U12565 (N_12565,N_11565,N_7528);
and U12566 (N_12566,N_6993,N_6968);
or U12567 (N_12567,N_7604,N_6730);
nand U12568 (N_12568,N_6345,N_7818);
and U12569 (N_12569,N_10213,N_9426);
xor U12570 (N_12570,N_10305,N_11293);
nand U12571 (N_12571,N_6466,N_8697);
nor U12572 (N_12572,N_9542,N_11385);
xor U12573 (N_12573,N_10254,N_8517);
nand U12574 (N_12574,N_10200,N_9805);
or U12575 (N_12575,N_9787,N_11222);
nor U12576 (N_12576,N_9634,N_6841);
and U12577 (N_12577,N_8824,N_8996);
nor U12578 (N_12578,N_10850,N_6492);
xnor U12579 (N_12579,N_10380,N_6380);
xnor U12580 (N_12580,N_9088,N_6226);
nor U12581 (N_12581,N_6830,N_9178);
xnor U12582 (N_12582,N_11969,N_11030);
xor U12583 (N_12583,N_6014,N_11078);
xnor U12584 (N_12584,N_8057,N_8921);
or U12585 (N_12585,N_10032,N_7542);
xnor U12586 (N_12586,N_9885,N_11187);
nand U12587 (N_12587,N_7819,N_7502);
or U12588 (N_12588,N_9123,N_7583);
or U12589 (N_12589,N_10890,N_11560);
nand U12590 (N_12590,N_7064,N_10705);
or U12591 (N_12591,N_6820,N_9623);
and U12592 (N_12592,N_6298,N_8161);
nand U12593 (N_12593,N_6781,N_8873);
or U12594 (N_12594,N_8361,N_8396);
or U12595 (N_12595,N_9345,N_10017);
and U12596 (N_12596,N_10037,N_6869);
nand U12597 (N_12597,N_8154,N_9949);
and U12598 (N_12598,N_9111,N_11045);
xor U12599 (N_12599,N_10451,N_7743);
and U12600 (N_12600,N_11982,N_8899);
xnor U12601 (N_12601,N_11579,N_10779);
or U12602 (N_12602,N_9982,N_7021);
and U12603 (N_12603,N_10295,N_11681);
nor U12604 (N_12604,N_6358,N_9694);
or U12605 (N_12605,N_11220,N_8482);
xnor U12606 (N_12606,N_11842,N_6800);
nor U12607 (N_12607,N_6406,N_9766);
or U12608 (N_12608,N_9791,N_11592);
and U12609 (N_12609,N_10950,N_7763);
and U12610 (N_12610,N_6165,N_7107);
nand U12611 (N_12611,N_11272,N_8582);
and U12612 (N_12612,N_11894,N_9074);
nand U12613 (N_12613,N_6931,N_8174);
or U12614 (N_12614,N_10515,N_6666);
nand U12615 (N_12615,N_10534,N_7264);
nor U12616 (N_12616,N_11455,N_6901);
or U12617 (N_12617,N_9926,N_9515);
and U12618 (N_12618,N_8840,N_6205);
or U12619 (N_12619,N_6086,N_8461);
xor U12620 (N_12620,N_9206,N_11851);
and U12621 (N_12621,N_11180,N_6313);
nor U12622 (N_12622,N_7046,N_6498);
and U12623 (N_12623,N_11746,N_6186);
nand U12624 (N_12624,N_11215,N_7068);
nand U12625 (N_12625,N_6700,N_6503);
and U12626 (N_12626,N_7875,N_10450);
and U12627 (N_12627,N_7194,N_6199);
nor U12628 (N_12628,N_10895,N_10031);
nor U12629 (N_12629,N_10685,N_8148);
nand U12630 (N_12630,N_10400,N_10274);
xor U12631 (N_12631,N_10147,N_7480);
xnor U12632 (N_12632,N_11322,N_10819);
or U12633 (N_12633,N_11227,N_8101);
xor U12634 (N_12634,N_6328,N_11785);
nor U12635 (N_12635,N_6927,N_10907);
nor U12636 (N_12636,N_10647,N_11924);
or U12637 (N_12637,N_7401,N_11667);
nand U12638 (N_12638,N_9931,N_7058);
nand U12639 (N_12639,N_6346,N_10056);
nor U12640 (N_12640,N_6409,N_10718);
xnor U12641 (N_12641,N_6420,N_11467);
and U12642 (N_12642,N_11529,N_8326);
nand U12643 (N_12643,N_6069,N_7275);
nor U12644 (N_12644,N_8643,N_10622);
or U12645 (N_12645,N_9466,N_11643);
nand U12646 (N_12646,N_11013,N_11392);
nor U12647 (N_12647,N_8606,N_11252);
nand U12648 (N_12648,N_8151,N_10683);
nand U12649 (N_12649,N_8732,N_10474);
or U12650 (N_12650,N_11915,N_10209);
or U12651 (N_12651,N_11003,N_11141);
xnor U12652 (N_12652,N_8995,N_11766);
nor U12653 (N_12653,N_8842,N_11612);
or U12654 (N_12654,N_9567,N_11985);
nor U12655 (N_12655,N_7087,N_8020);
nor U12656 (N_12656,N_7983,N_8961);
xnor U12657 (N_12657,N_8510,N_8798);
nor U12658 (N_12658,N_7741,N_6289);
xor U12659 (N_12659,N_6138,N_6096);
xnor U12660 (N_12660,N_7610,N_6507);
and U12661 (N_12661,N_8768,N_10456);
or U12662 (N_12662,N_9364,N_6643);
or U12663 (N_12663,N_10680,N_7642);
and U12664 (N_12664,N_9006,N_6303);
or U12665 (N_12665,N_11545,N_10742);
nor U12666 (N_12666,N_6306,N_7490);
and U12667 (N_12667,N_9631,N_6376);
or U12668 (N_12668,N_7436,N_11821);
and U12669 (N_12669,N_9858,N_8713);
or U12670 (N_12670,N_8010,N_9578);
nor U12671 (N_12671,N_6975,N_7136);
nor U12672 (N_12672,N_7655,N_11641);
or U12673 (N_12673,N_10933,N_10424);
or U12674 (N_12674,N_11007,N_9082);
nor U12675 (N_12675,N_6973,N_10313);
nand U12676 (N_12676,N_9683,N_9001);
xor U12677 (N_12677,N_10443,N_8759);
nand U12678 (N_12678,N_9653,N_7654);
nor U12679 (N_12679,N_10731,N_11124);
xor U12680 (N_12680,N_9218,N_11319);
or U12681 (N_12681,N_7022,N_7947);
nor U12682 (N_12682,N_6805,N_9738);
and U12683 (N_12683,N_11279,N_9988);
nand U12684 (N_12684,N_6158,N_11424);
and U12685 (N_12685,N_8023,N_8152);
nor U12686 (N_12686,N_6526,N_9149);
or U12687 (N_12687,N_7616,N_6863);
and U12688 (N_12688,N_9153,N_9711);
nand U12689 (N_12689,N_6807,N_9550);
nor U12690 (N_12690,N_6831,N_11738);
nor U12691 (N_12691,N_9158,N_11342);
or U12692 (N_12692,N_9512,N_6774);
nand U12693 (N_12693,N_8870,N_8962);
nand U12694 (N_12694,N_8998,N_10521);
or U12695 (N_12695,N_7451,N_9562);
or U12696 (N_12696,N_10357,N_9474);
or U12697 (N_12697,N_11780,N_7721);
nand U12698 (N_12698,N_9702,N_7869);
and U12699 (N_12699,N_10462,N_9652);
xnor U12700 (N_12700,N_7283,N_7623);
and U12701 (N_12701,N_7039,N_6918);
xnor U12702 (N_12702,N_9427,N_11925);
or U12703 (N_12703,N_8576,N_10321);
xor U12704 (N_12704,N_9465,N_11926);
xnor U12705 (N_12705,N_11520,N_6379);
nand U12706 (N_12706,N_6671,N_11255);
nand U12707 (N_12707,N_10575,N_7621);
or U12708 (N_12708,N_11399,N_10763);
xor U12709 (N_12709,N_10262,N_7371);
xnor U12710 (N_12710,N_8947,N_8209);
and U12711 (N_12711,N_9752,N_8734);
and U12712 (N_12712,N_9835,N_7559);
or U12713 (N_12713,N_11916,N_6689);
nand U12714 (N_12714,N_7301,N_6256);
nor U12715 (N_12715,N_7443,N_6872);
nand U12716 (N_12716,N_11031,N_9151);
and U12717 (N_12717,N_10113,N_11408);
or U12718 (N_12718,N_7224,N_6969);
nor U12719 (N_12719,N_9422,N_7888);
nand U12720 (N_12720,N_11485,N_7475);
nand U12721 (N_12721,N_6865,N_11888);
nor U12722 (N_12722,N_9739,N_6463);
or U12723 (N_12723,N_11677,N_9487);
xnor U12724 (N_12724,N_9140,N_6004);
and U12725 (N_12725,N_10157,N_6947);
xnor U12726 (N_12726,N_10008,N_9963);
or U12727 (N_12727,N_10775,N_7661);
nor U12728 (N_12728,N_10824,N_6525);
nand U12729 (N_12729,N_11202,N_11132);
nand U12730 (N_12730,N_8483,N_6718);
xnor U12731 (N_12731,N_11357,N_7185);
and U12732 (N_12732,N_8825,N_6546);
nor U12733 (N_12733,N_11388,N_6815);
nand U12734 (N_12734,N_9528,N_6180);
and U12735 (N_12735,N_6908,N_8337);
nand U12736 (N_12736,N_10916,N_6360);
or U12737 (N_12737,N_8806,N_6484);
nand U12738 (N_12738,N_7438,N_10565);
xor U12739 (N_12739,N_10009,N_7602);
nand U12740 (N_12740,N_6440,N_9312);
nand U12741 (N_12741,N_11816,N_10095);
and U12742 (N_12742,N_11494,N_8661);
nand U12743 (N_12743,N_8351,N_8539);
and U12744 (N_12744,N_10083,N_11175);
and U12745 (N_12745,N_10029,N_6944);
and U12746 (N_12746,N_10237,N_8820);
or U12747 (N_12747,N_7445,N_7932);
and U12748 (N_12748,N_11930,N_6316);
or U12749 (N_12749,N_10264,N_6736);
or U12750 (N_12750,N_6157,N_9193);
and U12751 (N_12751,N_8920,N_6031);
nor U12752 (N_12752,N_6600,N_8267);
nand U12753 (N_12753,N_11177,N_8508);
nand U12754 (N_12754,N_9797,N_11057);
nand U12755 (N_12755,N_6835,N_6126);
and U12756 (N_12756,N_6899,N_7606);
xnor U12757 (N_12757,N_8512,N_8407);
nand U12758 (N_12758,N_10007,N_7749);
or U12759 (N_12759,N_6428,N_11574);
xor U12760 (N_12760,N_8751,N_11701);
nor U12761 (N_12761,N_10204,N_9327);
nor U12762 (N_12762,N_7539,N_8617);
nand U12763 (N_12763,N_9569,N_10155);
xor U12764 (N_12764,N_7230,N_6943);
or U12765 (N_12765,N_10136,N_7635);
nor U12766 (N_12766,N_10404,N_10207);
and U12767 (N_12767,N_6247,N_10278);
nand U12768 (N_12768,N_11479,N_6609);
nand U12769 (N_12769,N_6701,N_10108);
nand U12770 (N_12770,N_11213,N_6537);
or U12771 (N_12771,N_8767,N_10074);
nor U12772 (N_12772,N_8011,N_7832);
nor U12773 (N_12773,N_7519,N_11301);
xor U12774 (N_12774,N_11524,N_11539);
and U12775 (N_12775,N_9817,N_11534);
or U12776 (N_12776,N_7365,N_7220);
nor U12777 (N_12777,N_6979,N_7870);
xnor U12778 (N_12778,N_11502,N_7255);
nand U12779 (N_12779,N_11906,N_10707);
and U12780 (N_12780,N_7461,N_6588);
or U12781 (N_12781,N_6868,N_8550);
nor U12782 (N_12782,N_6072,N_7643);
nor U12783 (N_12783,N_6619,N_9036);
and U12784 (N_12784,N_6333,N_6073);
nand U12785 (N_12785,N_10800,N_8314);
and U12786 (N_12786,N_7246,N_7265);
nand U12787 (N_12787,N_8012,N_10667);
or U12788 (N_12788,N_8163,N_11956);
nor U12789 (N_12789,N_8413,N_9284);
and U12790 (N_12790,N_7494,N_8207);
and U12791 (N_12791,N_10442,N_9785);
nor U12792 (N_12792,N_10461,N_10972);
nand U12793 (N_12793,N_10612,N_6933);
nand U12794 (N_12794,N_11532,N_6206);
xnor U12795 (N_12795,N_9115,N_9213);
nand U12796 (N_12796,N_8444,N_9703);
nor U12797 (N_12797,N_6099,N_8153);
nand U12798 (N_12798,N_11702,N_11023);
or U12799 (N_12799,N_10413,N_6995);
xor U12800 (N_12800,N_9611,N_10242);
xor U12801 (N_12801,N_11450,N_8956);
nand U12802 (N_12802,N_8013,N_11055);
and U12803 (N_12803,N_6584,N_6135);
or U12804 (N_12804,N_9643,N_10553);
or U12805 (N_12805,N_9096,N_9831);
or U12806 (N_12806,N_7376,N_9262);
xor U12807 (N_12807,N_11822,N_10250);
or U12808 (N_12808,N_9340,N_6223);
nand U12809 (N_12809,N_7814,N_10094);
and U12810 (N_12810,N_10942,N_8730);
or U12811 (N_12811,N_8387,N_9709);
and U12812 (N_12812,N_7345,N_6876);
xor U12813 (N_12813,N_9932,N_7942);
xnor U12814 (N_12814,N_9958,N_6259);
nor U12815 (N_12815,N_7139,N_11236);
xnor U12816 (N_12816,N_9524,N_10805);
and U12817 (N_12817,N_6817,N_10560);
xor U12818 (N_12818,N_11922,N_10615);
nand U12819 (N_12819,N_6451,N_7110);
nor U12820 (N_12820,N_11162,N_11783);
or U12821 (N_12821,N_8183,N_6842);
xor U12822 (N_12822,N_8158,N_10998);
xor U12823 (N_12823,N_11892,N_6018);
nand U12824 (N_12824,N_6494,N_6452);
nand U12825 (N_12825,N_10614,N_11558);
and U12826 (N_12826,N_10656,N_9148);
nor U12827 (N_12827,N_9582,N_8323);
nand U12828 (N_12828,N_6161,N_10864);
nand U12829 (N_12829,N_7724,N_11400);
nor U12830 (N_12830,N_9049,N_11955);
nand U12831 (N_12831,N_11260,N_6678);
xnor U12832 (N_12832,N_10234,N_9908);
nand U12833 (N_12833,N_7063,N_11503);
nor U12834 (N_12834,N_11129,N_10423);
xnor U12835 (N_12835,N_10504,N_6178);
nor U12836 (N_12836,N_10746,N_7504);
or U12837 (N_12837,N_8803,N_9773);
nor U12838 (N_12838,N_8785,N_10835);
or U12839 (N_12839,N_8120,N_7098);
nand U12840 (N_12840,N_9925,N_7536);
or U12841 (N_12841,N_6989,N_9920);
xor U12842 (N_12842,N_7784,N_6263);
xor U12843 (N_12843,N_8186,N_8626);
or U12844 (N_12844,N_9910,N_8864);
nand U12845 (N_12845,N_11587,N_8437);
nor U12846 (N_12846,N_10956,N_9217);
or U12847 (N_12847,N_10825,N_7120);
or U12848 (N_12848,N_11254,N_7388);
and U12849 (N_12849,N_10379,N_8758);
and U12850 (N_12850,N_11082,N_10610);
and U12851 (N_12851,N_11530,N_7215);
nand U12852 (N_12852,N_10277,N_8061);
and U12853 (N_12853,N_8390,N_11459);
xor U12854 (N_12854,N_10929,N_8243);
nor U12855 (N_12855,N_10437,N_10105);
nor U12856 (N_12856,N_10725,N_10566);
nand U12857 (N_12857,N_9554,N_9568);
or U12858 (N_12858,N_7385,N_8989);
and U12859 (N_12859,N_11345,N_7002);
or U12860 (N_12860,N_9896,N_8450);
nand U12861 (N_12861,N_7400,N_10827);
nor U12862 (N_12862,N_7083,N_11682);
xnor U12863 (N_12863,N_7596,N_8609);
nor U12864 (N_12864,N_7231,N_9332);
xor U12865 (N_12865,N_10088,N_8053);
or U12866 (N_12866,N_9608,N_9854);
nand U12867 (N_12867,N_9923,N_11015);
xor U12868 (N_12868,N_6743,N_6123);
nand U12869 (N_12869,N_10796,N_6164);
nand U12870 (N_12870,N_11882,N_10744);
nor U12871 (N_12871,N_11996,N_10629);
xnor U12872 (N_12872,N_8788,N_9936);
xor U12873 (N_12873,N_6231,N_7940);
nor U12874 (N_12874,N_8355,N_8595);
xor U12875 (N_12875,N_9518,N_11340);
and U12876 (N_12876,N_10531,N_11131);
xnor U12877 (N_12877,N_8623,N_9406);
and U12878 (N_12878,N_7805,N_7410);
and U12879 (N_12879,N_10847,N_10922);
or U12880 (N_12880,N_11324,N_11232);
or U12881 (N_12881,N_6629,N_10855);
xor U12882 (N_12882,N_8068,N_10597);
xor U12883 (N_12883,N_7351,N_6798);
nand U12884 (N_12884,N_10889,N_8420);
xor U12885 (N_12885,N_6254,N_6620);
nor U12886 (N_12886,N_6097,N_8427);
or U12887 (N_12887,N_8575,N_9615);
and U12888 (N_12888,N_10142,N_8879);
or U12889 (N_12889,N_9198,N_8312);
or U12890 (N_12890,N_6152,N_9138);
nand U12891 (N_12891,N_6806,N_11146);
and U12892 (N_12892,N_9468,N_10928);
or U12893 (N_12893,N_10810,N_6204);
and U12894 (N_12894,N_8059,N_11610);
and U12895 (N_12895,N_8356,N_8656);
xnor U12896 (N_12896,N_9837,N_10378);
nand U12897 (N_12897,N_11988,N_10171);
nor U12898 (N_12898,N_6202,N_9022);
xor U12899 (N_12899,N_11804,N_9664);
nand U12900 (N_12900,N_9783,N_9849);
nor U12901 (N_12901,N_6660,N_10103);
and U12902 (N_12902,N_6981,N_6296);
nor U12903 (N_12903,N_11824,N_9525);
nor U12904 (N_12904,N_8903,N_10721);
or U12905 (N_12905,N_9104,N_11245);
or U12906 (N_12906,N_6403,N_6281);
nand U12907 (N_12907,N_9913,N_9420);
or U12908 (N_12908,N_9136,N_7406);
nor U12909 (N_12909,N_7984,N_11854);
xnor U12910 (N_12910,N_8834,N_9481);
nand U12911 (N_12911,N_9097,N_8717);
or U12912 (N_12912,N_8752,N_8225);
nand U12913 (N_12913,N_9230,N_9265);
nand U12914 (N_12914,N_8584,N_10627);
nor U12915 (N_12915,N_6621,N_8082);
nor U12916 (N_12916,N_9510,N_10102);
xor U12917 (N_12917,N_10381,N_7179);
nor U12918 (N_12918,N_6091,N_9396);
or U12919 (N_12919,N_10638,N_11234);
xnor U12920 (N_12920,N_7042,N_8190);
and U12921 (N_12921,N_11378,N_9918);
nand U12922 (N_12922,N_8944,N_11147);
nand U12923 (N_12923,N_9020,N_7244);
and U12924 (N_12924,N_11538,N_7740);
or U12925 (N_12925,N_7591,N_8132);
xor U12926 (N_12926,N_8535,N_10625);
and U12927 (N_12927,N_11730,N_8997);
xnor U12928 (N_12928,N_8639,N_7260);
or U12929 (N_12929,N_11246,N_10968);
xor U12930 (N_12930,N_10036,N_10848);
xnor U12931 (N_12931,N_11267,N_6732);
and U12932 (N_12932,N_7682,N_8580);
nand U12933 (N_12933,N_10701,N_11767);
nor U12934 (N_12934,N_6269,N_11052);
and U12935 (N_12935,N_10591,N_7829);
nor U12936 (N_12936,N_10193,N_6782);
and U12937 (N_12937,N_9586,N_9224);
and U12938 (N_12938,N_6487,N_6714);
nand U12939 (N_12939,N_6354,N_7293);
or U12940 (N_12940,N_10276,N_11817);
or U12941 (N_12941,N_6251,N_10006);
and U12942 (N_12942,N_9092,N_10432);
and U12943 (N_12943,N_8172,N_9603);
nor U12944 (N_12944,N_7112,N_9062);
or U12945 (N_12945,N_11855,N_8748);
xnor U12946 (N_12946,N_8951,N_10143);
nand U12947 (N_12947,N_11959,N_6723);
nor U12948 (N_12948,N_11063,N_6238);
or U12949 (N_12949,N_9588,N_7764);
nand U12950 (N_12950,N_10060,N_9382);
xnor U12951 (N_12951,N_9505,N_8953);
or U12952 (N_12952,N_10347,N_9930);
or U12953 (N_12953,N_11998,N_7758);
or U12954 (N_12954,N_6212,N_11439);
xnor U12955 (N_12955,N_9169,N_6347);
xnor U12956 (N_12956,N_9736,N_11978);
or U12957 (N_12957,N_8866,N_7469);
xnor U12958 (N_12958,N_8469,N_6475);
or U12959 (N_12959,N_7023,N_10626);
nand U12960 (N_12960,N_8479,N_10390);
nor U12961 (N_12961,N_6855,N_6589);
or U12962 (N_12962,N_6886,N_6170);
or U12963 (N_12963,N_9662,N_8126);
nor U12964 (N_12964,N_9318,N_6690);
xor U12965 (N_12965,N_11709,N_9187);
nand U12966 (N_12966,N_10013,N_11081);
or U12967 (N_12967,N_8663,N_6377);
nor U12968 (N_12968,N_11954,N_6680);
nand U12969 (N_12969,N_8160,N_9869);
nor U12970 (N_12970,N_11631,N_8056);
xnor U12971 (N_12971,N_8931,N_7196);
xnor U12972 (N_12972,N_6598,N_9618);
nor U12973 (N_12973,N_8802,N_7657);
nand U12974 (N_12974,N_7878,N_7793);
xor U12975 (N_12975,N_7059,N_7108);
and U12976 (N_12976,N_7695,N_6623);
nor U12977 (N_12977,N_8591,N_9589);
and U12978 (N_12978,N_10765,N_7834);
and U12979 (N_12979,N_8858,N_6994);
and U12980 (N_12980,N_8744,N_7510);
or U12981 (N_12981,N_8279,N_7518);
nor U12982 (N_12982,N_10266,N_7690);
and U12983 (N_12983,N_9338,N_10736);
or U12984 (N_12984,N_11887,N_6301);
nand U12985 (N_12985,N_6283,N_11898);
xor U12986 (N_12986,N_9147,N_6914);
and U12987 (N_12987,N_8887,N_9648);
nor U12988 (N_12988,N_8597,N_8196);
nand U12989 (N_12989,N_10226,N_7165);
xor U12990 (N_12990,N_8146,N_6282);
or U12991 (N_12991,N_10051,N_7953);
and U12992 (N_12992,N_10220,N_10961);
or U12993 (N_12993,N_10983,N_11868);
or U12994 (N_12994,N_7915,N_9467);
or U12995 (N_12995,N_11506,N_7026);
nor U12996 (N_12996,N_8955,N_9551);
and U12997 (N_12997,N_7036,N_7844);
nand U12998 (N_12998,N_8976,N_9793);
nor U12999 (N_12999,N_8932,N_8344);
or U13000 (N_13000,N_8108,N_11943);
or U13001 (N_13001,N_10330,N_10635);
nor U13002 (N_13002,N_9028,N_10427);
or U13003 (N_13003,N_8552,N_10947);
or U13004 (N_13004,N_7811,N_7286);
nor U13005 (N_13005,N_8371,N_11602);
or U13006 (N_13006,N_10385,N_8509);
or U13007 (N_13007,N_8327,N_8737);
nand U13008 (N_13008,N_7912,N_8769);
nor U13009 (N_13009,N_8515,N_8863);
and U13010 (N_13010,N_7968,N_9841);
xnor U13011 (N_13011,N_8524,N_6450);
nor U13012 (N_13012,N_10943,N_10523);
or U13013 (N_13013,N_10642,N_7197);
nor U13014 (N_13014,N_6433,N_11590);
nor U13015 (N_13015,N_7072,N_7393);
and U13016 (N_13016,N_6814,N_10034);
nand U13017 (N_13017,N_10464,N_10936);
or U13018 (N_13018,N_6309,N_7570);
or U13019 (N_13019,N_6167,N_11036);
nor U13020 (N_13020,N_11664,N_10080);
nand U13021 (N_13021,N_6461,N_9479);
or U13022 (N_13022,N_6115,N_7900);
nor U13023 (N_13023,N_8162,N_8796);
xor U13024 (N_13024,N_6216,N_7990);
xnor U13025 (N_13025,N_7910,N_7363);
or U13026 (N_13026,N_10208,N_11661);
nor U13027 (N_13027,N_6489,N_10360);
xor U13028 (N_13028,N_8664,N_7272);
nand U13029 (N_13029,N_8418,N_7597);
and U13030 (N_13030,N_8696,N_10986);
nand U13031 (N_13031,N_6218,N_11453);
and U13032 (N_13032,N_9635,N_9973);
nand U13033 (N_13033,N_6378,N_10913);
nand U13034 (N_13034,N_6515,N_6509);
or U13035 (N_13035,N_10937,N_7088);
nand U13036 (N_13036,N_10446,N_11094);
nor U13037 (N_13037,N_10962,N_8036);
nor U13038 (N_13038,N_6462,N_11652);
or U13039 (N_13039,N_6125,N_10382);
or U13040 (N_13040,N_11478,N_10706);
and U13041 (N_13041,N_11414,N_6171);
xnor U13042 (N_13042,N_6471,N_10700);
and U13043 (N_13043,N_8511,N_6449);
or U13044 (N_13044,N_6397,N_10654);
nand U13045 (N_13045,N_11742,N_11383);
nand U13046 (N_13046,N_8045,N_11210);
xnor U13047 (N_13047,N_6305,N_8793);
nand U13048 (N_13048,N_7337,N_10303);
nor U13049 (N_13049,N_6583,N_11627);
nand U13050 (N_13050,N_6813,N_9747);
xnor U13051 (N_13051,N_8845,N_9546);
nor U13052 (N_13052,N_11659,N_7299);
nand U13053 (N_13053,N_11691,N_7672);
xor U13054 (N_13054,N_10628,N_8611);
and U13055 (N_13055,N_6521,N_8979);
nor U13056 (N_13056,N_11937,N_8642);
nor U13057 (N_13057,N_8811,N_9561);
nor U13058 (N_13058,N_10743,N_8025);
nor U13059 (N_13059,N_9861,N_10543);
or U13060 (N_13060,N_6010,N_11628);
xor U13061 (N_13061,N_11741,N_8223);
nor U13062 (N_13062,N_11247,N_11572);
xnor U13063 (N_13063,N_7028,N_6958);
and U13064 (N_13064,N_11786,N_8589);
or U13065 (N_13065,N_6960,N_8690);
nor U13066 (N_13066,N_10253,N_8131);
and U13067 (N_13067,N_6179,N_9597);
or U13068 (N_13068,N_7362,N_7273);
nor U13069 (N_13069,N_11830,N_6321);
or U13070 (N_13070,N_10158,N_8235);
and U13071 (N_13071,N_10251,N_11986);
or U13072 (N_13072,N_6552,N_9834);
and U13073 (N_13073,N_9842,N_7373);
xor U13074 (N_13074,N_9478,N_10287);
xor U13075 (N_13075,N_6948,N_10732);
or U13076 (N_13076,N_8993,N_10927);
or U13077 (N_13077,N_9319,N_8849);
and U13078 (N_13078,N_6398,N_8200);
nor U13079 (N_13079,N_10180,N_9646);
nand U13080 (N_13080,N_11939,N_7474);
and U13081 (N_13081,N_7316,N_6056);
and U13082 (N_13082,N_6911,N_9895);
nand U13083 (N_13083,N_8765,N_8710);
nor U13084 (N_13084,N_9423,N_7903);
nor U13085 (N_13085,N_9753,N_11543);
nand U13086 (N_13086,N_11056,N_6065);
nand U13087 (N_13087,N_8405,N_10041);
nand U13088 (N_13088,N_6062,N_11706);
and U13089 (N_13089,N_8897,N_6984);
xnor U13090 (N_13090,N_6504,N_9565);
and U13091 (N_13091,N_9186,N_6063);
or U13092 (N_13092,N_11668,N_6217);
and U13093 (N_13093,N_7557,N_6615);
or U13094 (N_13094,N_10291,N_11364);
or U13095 (N_13095,N_11109,N_6860);
nor U13096 (N_13096,N_9183,N_7423);
or U13097 (N_13097,N_7151,N_11688);
nand U13098 (N_13098,N_7118,N_7396);
nor U13099 (N_13099,N_9091,N_9820);
nor U13100 (N_13100,N_6326,N_11189);
xor U13101 (N_13101,N_10533,N_8640);
nor U13102 (N_13102,N_11107,N_10479);
xor U13103 (N_13103,N_7590,N_9705);
nor U13104 (N_13104,N_6524,N_10211);
or U13105 (N_13105,N_9204,N_7813);
or U13106 (N_13106,N_7995,N_7429);
nand U13107 (N_13107,N_11990,N_9171);
or U13108 (N_13108,N_11070,N_10584);
and U13109 (N_13109,N_10281,N_9259);
or U13110 (N_13110,N_7076,N_6704);
or U13111 (N_13111,N_10109,N_6479);
or U13112 (N_13112,N_7183,N_11278);
or U13113 (N_13113,N_8660,N_8006);
and U13114 (N_13114,N_7825,N_10263);
or U13115 (N_13115,N_7148,N_11705);
or U13116 (N_13116,N_7608,N_6741);
xnor U13117 (N_13117,N_7073,N_8685);
xnor U13118 (N_13118,N_10538,N_11630);
nand U13119 (N_13119,N_7563,N_9681);
nand U13120 (N_13120,N_7347,N_8491);
nor U13121 (N_13121,N_8843,N_7311);
or U13122 (N_13122,N_11576,N_6547);
and U13123 (N_13123,N_6558,N_8236);
nor U13124 (N_13124,N_8404,N_9303);
or U13125 (N_13125,N_7162,N_6826);
nand U13126 (N_13126,N_8590,N_10069);
nor U13127 (N_13127,N_10311,N_7222);
nand U13128 (N_13128,N_11878,N_7383);
or U13129 (N_13129,N_6160,N_6717);
or U13130 (N_13130,N_7954,N_11238);
or U13131 (N_13131,N_10144,N_11867);
nor U13132 (N_13132,N_11310,N_9141);
and U13133 (N_13133,N_8952,N_8318);
or U13134 (N_13134,N_7609,N_10788);
and U13135 (N_13135,N_8454,N_10399);
nand U13136 (N_13136,N_6225,N_10063);
xor U13137 (N_13137,N_8808,N_9166);
or U13138 (N_13138,N_9346,N_6295);
and U13139 (N_13139,N_6473,N_11462);
xor U13140 (N_13140,N_10419,N_8281);
xnor U13141 (N_13141,N_10414,N_6789);
and U13142 (N_13142,N_9976,N_9379);
xnor U13143 (N_13143,N_9251,N_9026);
or U13144 (N_13144,N_6418,N_10830);
or U13145 (N_13145,N_7453,N_11909);
nand U13146 (N_13146,N_11774,N_11338);
nand U13147 (N_13147,N_6284,N_6153);
xor U13148 (N_13148,N_8711,N_10401);
nor U13149 (N_13149,N_9784,N_11900);
nor U13150 (N_13150,N_9491,N_10737);
and U13151 (N_13151,N_9053,N_11233);
and U13152 (N_13152,N_7402,N_7313);
or U13153 (N_13153,N_9347,N_11807);
nor U13154 (N_13154,N_6603,N_7116);
and U13155 (N_13155,N_10406,N_6616);
nor U13156 (N_13156,N_11256,N_11395);
nor U13157 (N_13157,N_8774,N_9649);
nand U13158 (N_13158,N_6792,N_6001);
nand U13159 (N_13159,N_8800,N_7574);
xor U13160 (N_13160,N_6923,N_7619);
xnor U13161 (N_13161,N_9214,N_9940);
xnor U13162 (N_13162,N_7882,N_10949);
and U13163 (N_13163,N_8215,N_8232);
and U13164 (N_13164,N_7387,N_7495);
and U13165 (N_13165,N_9418,N_9211);
and U13166 (N_13166,N_10669,N_7324);
xnor U13167 (N_13167,N_6569,N_6864);
nor U13168 (N_13168,N_11398,N_6275);
nor U13169 (N_13169,N_10351,N_9291);
or U13170 (N_13170,N_11809,N_10151);
nor U13171 (N_13171,N_9534,N_6429);
nand U13172 (N_13172,N_6881,N_8043);
or U13173 (N_13173,N_7697,N_9063);
and U13174 (N_13174,N_11461,N_9120);
and U13175 (N_13175,N_7302,N_10269);
and U13176 (N_13176,N_7848,N_10866);
nand U13177 (N_13177,N_10618,N_10048);
xor U13178 (N_13178,N_11734,N_7125);
or U13179 (N_13179,N_8869,N_7239);
nand U13180 (N_13180,N_9691,N_8937);
xor U13181 (N_13181,N_8321,N_10592);
nand U13182 (N_13182,N_8708,N_7535);
and U13183 (N_13183,N_11475,N_11981);
nor U13184 (N_13184,N_8850,N_10028);
xor U13185 (N_13185,N_7883,N_7195);
nand U13186 (N_13186,N_9222,N_9994);
or U13187 (N_13187,N_10588,N_6410);
xnor U13188 (N_13188,N_6085,N_10517);
nor U13189 (N_13189,N_8747,N_6765);
xor U13190 (N_13190,N_11402,N_7933);
and U13191 (N_13191,N_8719,N_7524);
xnor U13192 (N_13192,N_7617,N_8113);
or U13193 (N_13193,N_9398,N_10374);
nand U13194 (N_13194,N_6336,N_11316);
nand U13195 (N_13195,N_11829,N_9802);
or U13196 (N_13196,N_11412,N_6474);
nand U13197 (N_13197,N_11989,N_9397);
and U13198 (N_13198,N_9108,N_9778);
and U13199 (N_13199,N_7153,N_6926);
or U13200 (N_13200,N_9780,N_11771);
nand U13201 (N_13201,N_11193,N_10296);
nand U13202 (N_13202,N_10520,N_7096);
or U13203 (N_13203,N_10327,N_6373);
or U13204 (N_13204,N_10288,N_10439);
nand U13205 (N_13205,N_9116,N_10604);
nor U13206 (N_13206,N_6966,N_7432);
and U13207 (N_13207,N_9555,N_11907);
xor U13208 (N_13208,N_10993,N_8070);
and U13209 (N_13209,N_8969,N_8610);
nor U13210 (N_13210,N_7078,N_10405);
xor U13211 (N_13211,N_7828,N_9307);
xnor U13212 (N_13212,N_7816,N_11699);
nor U13213 (N_13213,N_10676,N_8414);
xnor U13214 (N_13214,N_8809,N_6592);
nand U13215 (N_13215,N_11393,N_11671);
and U13216 (N_13216,N_8780,N_9760);
xor U13217 (N_13217,N_8241,N_7278);
nor U13218 (N_13218,N_6987,N_7837);
xor U13219 (N_13219,N_7435,N_8917);
or U13220 (N_13220,N_11836,N_11992);
or U13221 (N_13221,N_7949,N_8166);
and U13222 (N_13222,N_10449,N_7491);
or U13223 (N_13223,N_11845,N_8328);
or U13224 (N_13224,N_7960,N_9055);
or U13225 (N_13225,N_8257,N_9061);
nand U13226 (N_13226,N_8542,N_10502);
or U13227 (N_13227,N_6528,N_11184);
and U13228 (N_13228,N_9878,N_10318);
nor U13229 (N_13229,N_10490,N_7192);
xnor U13230 (N_13230,N_11433,N_10754);
nor U13231 (N_13231,N_9884,N_8353);
and U13232 (N_13232,N_6897,N_8726);
and U13233 (N_13233,N_11675,N_8692);
or U13234 (N_13234,N_6677,N_10975);
and U13235 (N_13235,N_8612,N_10440);
or U13236 (N_13236,N_7150,N_6520);
nand U13237 (N_13237,N_9924,N_10722);
nand U13238 (N_13238,N_7127,N_10117);
and U13239 (N_13239,N_6964,N_11290);
and U13240 (N_13240,N_10168,N_6648);
xnor U13241 (N_13241,N_11940,N_11253);
xor U13242 (N_13242,N_10239,N_9363);
and U13243 (N_13243,N_8742,N_6532);
nand U13244 (N_13244,N_6134,N_10428);
and U13245 (N_13245,N_6563,N_10232);
nand U13246 (N_13246,N_8125,N_6556);
nand U13247 (N_13247,N_11942,N_10904);
nand U13248 (N_13248,N_6626,N_7966);
nand U13249 (N_13249,N_10516,N_6026);
xnor U13250 (N_13250,N_10326,N_8603);
and U13251 (N_13251,N_9094,N_7307);
nand U13252 (N_13252,N_10500,N_6710);
or U13253 (N_13253,N_11285,N_9235);
nand U13254 (N_13254,N_11768,N_7658);
xor U13255 (N_13255,N_11438,N_11908);
or U13256 (N_13256,N_10346,N_7355);
nand U13257 (N_13257,N_7304,N_9326);
and U13258 (N_13258,N_10657,N_9570);
nand U13259 (N_13259,N_9928,N_10148);
nor U13260 (N_13260,N_10388,N_8226);
xnor U13261 (N_13261,N_6322,N_7133);
xnor U13262 (N_13262,N_11032,N_6636);
nand U13263 (N_13263,N_9270,N_6184);
nor U13264 (N_13264,N_7000,N_8942);
nor U13265 (N_13265,N_11088,N_8035);
nand U13266 (N_13266,N_10525,N_10054);
xnor U13267 (N_13267,N_8001,N_7614);
and U13268 (N_13268,N_9549,N_6627);
and U13269 (N_13269,N_7852,N_11843);
nor U13270 (N_13270,N_7018,N_11271);
xor U13271 (N_13271,N_6318,N_11941);
or U13272 (N_13272,N_8463,N_8141);
nor U13273 (N_13273,N_6591,N_7945);
or U13274 (N_13274,N_9756,N_6904);
and U13275 (N_13275,N_7671,N_9399);
nor U13276 (N_13276,N_11102,N_8757);
xnor U13277 (N_13277,N_11423,N_9616);
nor U13278 (N_13278,N_8216,N_8706);
and U13279 (N_13279,N_10422,N_7343);
nand U13280 (N_13280,N_10170,N_10528);
nand U13281 (N_13281,N_11191,N_11420);
xnor U13282 (N_13282,N_8348,N_6768);
nor U13283 (N_13283,N_9596,N_7130);
or U13284 (N_13284,N_7736,N_11962);
or U13285 (N_13285,N_11561,N_7985);
and U13286 (N_13286,N_10997,N_10472);
xnor U13287 (N_13287,N_8307,N_8691);
nor U13288 (N_13288,N_7579,N_11315);
or U13289 (N_13289,N_9188,N_11860);
nand U13290 (N_13290,N_7492,N_11837);
xor U13291 (N_13291,N_7257,N_9209);
nor U13292 (N_13292,N_6985,N_6833);
and U13293 (N_13293,N_7514,N_8066);
nor U13294 (N_13294,N_7729,N_6408);
nor U13295 (N_13295,N_10118,N_11403);
or U13296 (N_13296,N_10376,N_9241);
nor U13297 (N_13297,N_6300,N_10897);
and U13298 (N_13298,N_8918,N_6277);
or U13299 (N_13299,N_10179,N_6713);
nor U13300 (N_13300,N_8332,N_7024);
nor U13301 (N_13301,N_7785,N_6613);
xnor U13302 (N_13302,N_11476,N_10651);
nor U13303 (N_13303,N_11103,N_6998);
nor U13304 (N_13304,N_8122,N_8439);
or U13305 (N_13305,N_6803,N_11802);
nor U13306 (N_13306,N_10173,N_7778);
nor U13307 (N_13307,N_10120,N_10663);
nor U13308 (N_13308,N_7032,N_10339);
nor U13309 (N_13309,N_9929,N_7971);
xor U13310 (N_13310,N_6155,N_8914);
xor U13311 (N_13311,N_8277,N_10369);
nand U13312 (N_13312,N_9998,N_10552);
and U13313 (N_13313,N_8533,N_9155);
nor U13314 (N_13314,N_10636,N_6011);
and U13315 (N_13315,N_9157,N_11397);
nand U13316 (N_13316,N_7312,N_8859);
or U13317 (N_13317,N_11064,N_9748);
nor U13318 (N_13318,N_9799,N_9927);
nor U13319 (N_13319,N_9808,N_6469);
xnor U13320 (N_13320,N_11831,N_10648);
or U13321 (N_13321,N_8634,N_6034);
xnor U13322 (N_13322,N_9996,N_10994);
xnor U13323 (N_13323,N_6930,N_9197);
nand U13324 (N_13324,N_6467,N_8265);
nor U13325 (N_13325,N_8428,N_6434);
nor U13326 (N_13326,N_10987,N_11626);
nor U13327 (N_13327,N_8683,N_11119);
or U13328 (N_13328,N_6724,N_7680);
xnor U13329 (N_13329,N_9883,N_7584);
or U13330 (N_13330,N_9593,N_8736);
xor U13331 (N_13331,N_9601,N_6020);
or U13332 (N_13332,N_6696,N_10632);
or U13333 (N_13333,N_7902,N_11314);
and U13334 (N_13334,N_8062,N_6230);
xnor U13335 (N_13335,N_10695,N_6310);
xor U13336 (N_13336,N_6189,N_10498);
and U13337 (N_13337,N_10793,N_10177);
xor U13338 (N_13338,N_6631,N_11018);
nor U13339 (N_13339,N_10049,N_6012);
nand U13340 (N_13340,N_11066,N_11983);
and U13341 (N_13341,N_9404,N_10248);
nand U13342 (N_13342,N_9548,N_10697);
xor U13343 (N_13343,N_8194,N_11715);
and U13344 (N_13344,N_8477,N_10481);
nor U13345 (N_13345,N_6856,N_6095);
and U13346 (N_13346,N_6239,N_6682);
nand U13347 (N_13347,N_6081,N_6688);
xor U13348 (N_13348,N_8949,N_11472);
nand U13349 (N_13349,N_8116,N_10338);
nand U13350 (N_13350,N_6002,N_9011);
nor U13351 (N_13351,N_7728,N_8324);
xnor U13352 (N_13352,N_7168,N_8219);
nor U13353 (N_13353,N_10870,N_7117);
nor U13354 (N_13354,N_9242,N_9598);
xnor U13355 (N_13355,N_11581,N_10019);
and U13356 (N_13356,N_7905,N_9228);
and U13357 (N_13357,N_8369,N_6299);
or U13358 (N_13358,N_10471,N_11413);
nor U13359 (N_13359,N_6565,N_9070);
xnor U13360 (N_13360,N_8315,N_10079);
xnor U13361 (N_13361,N_10828,N_11432);
and U13362 (N_13362,N_7586,N_7589);
nand U13363 (N_13363,N_10816,N_6608);
or U13364 (N_13364,N_7056,N_9031);
or U13365 (N_13365,N_7100,N_7186);
xor U13366 (N_13366,N_9575,N_7864);
nand U13367 (N_13367,N_9150,N_11295);
xnor U13368 (N_13368,N_10286,N_10340);
xor U13369 (N_13369,N_11020,N_10637);
nand U13370 (N_13370,N_8284,N_8173);
or U13371 (N_13371,N_9124,N_8657);
xor U13372 (N_13372,N_9388,N_7517);
nor U13373 (N_13373,N_7124,N_9771);
nor U13374 (N_13374,N_9005,N_10849);
xnor U13375 (N_13375,N_8065,N_11890);
and U13376 (N_13376,N_9433,N_11139);
or U13377 (N_13377,N_11376,N_8970);
nand U13378 (N_13378,N_9075,N_8904);
or U13379 (N_13379,N_6739,N_10901);
and U13380 (N_13380,N_8650,N_11606);
or U13381 (N_13381,N_7380,N_7449);
and U13382 (N_13382,N_8615,N_10574);
nand U13383 (N_13383,N_6910,N_7458);
or U13384 (N_13384,N_6712,N_7973);
nor U13385 (N_13385,N_8275,N_8087);
nor U13386 (N_13386,N_11085,N_11651);
xnor U13387 (N_13387,N_7868,N_6787);
nand U13388 (N_13388,N_11775,N_6924);
or U13389 (N_13389,N_7891,N_8616);
nor U13390 (N_13390,N_7771,N_10633);
nor U13391 (N_13391,N_9281,N_6077);
xor U13392 (N_13392,N_9763,N_9215);
xnor U13393 (N_13393,N_11381,N_6240);
or U13394 (N_13394,N_10999,N_11034);
nand U13395 (N_13395,N_8492,N_11457);
nor U13396 (N_13396,N_11156,N_10946);
and U13397 (N_13397,N_10769,N_10244);
nand U13398 (N_13398,N_11555,N_10484);
nor U13399 (N_13399,N_9438,N_6279);
xnor U13400 (N_13400,N_11546,N_9430);
nand U13401 (N_13401,N_7262,N_9060);
and U13402 (N_13402,N_9751,N_7531);
and U13403 (N_13403,N_10869,N_8409);
nor U13404 (N_13404,N_9888,N_9745);
and U13405 (N_13405,N_11639,N_6510);
nor U13406 (N_13406,N_7648,N_6891);
and U13407 (N_13407,N_6442,N_8847);
nand U13408 (N_13408,N_8829,N_8659);
nand U13409 (N_13409,N_9981,N_9010);
or U13410 (N_13410,N_7881,N_7370);
nor U13411 (N_13411,N_6974,N_11963);
or U13412 (N_13412,N_9946,N_8761);
and U13413 (N_13413,N_10884,N_8456);
xnor U13414 (N_13414,N_10655,N_9682);
nor U13415 (N_13415,N_9410,N_6051);
xor U13416 (N_13416,N_9002,N_11387);
nor U13417 (N_13417,N_6832,N_9131);
nand U13418 (N_13418,N_9167,N_6746);
or U13419 (N_13419,N_9859,N_8709);
xor U13420 (N_13420,N_6047,N_8865);
and U13421 (N_13421,N_11291,N_10350);
and U13422 (N_13422,N_8135,N_8916);
or U13423 (N_13423,N_10755,N_9637);
or U13424 (N_13424,N_9349,N_6767);
nand U13425 (N_13425,N_10854,N_10020);
and U13426 (N_13426,N_6762,N_9746);
nor U13427 (N_13427,N_8139,N_7496);
and U13428 (N_13428,N_11500,N_8280);
or U13429 (N_13429,N_6430,N_10760);
nor U13430 (N_13430,N_9619,N_7203);
or U13431 (N_13431,N_7755,N_10518);
or U13432 (N_13432,N_6323,N_9381);
xor U13433 (N_13433,N_8354,N_10955);
nand U13434 (N_13434,N_10511,N_8927);
nand U13435 (N_13435,N_7756,N_7465);
nand U13436 (N_13436,N_6457,N_8922);
nand U13437 (N_13437,N_7872,N_6200);
nand U13438 (N_13438,N_9881,N_10587);
xor U13439 (N_13439,N_11720,N_9109);
or U13440 (N_13440,N_8519,N_11654);
and U13441 (N_13441,N_10156,N_8588);
and U13442 (N_13442,N_6053,N_9162);
and U13443 (N_13443,N_8675,N_9656);
or U13444 (N_13444,N_10548,N_10826);
or U13445 (N_13445,N_8472,N_8791);
nor U13446 (N_13446,N_11437,N_11328);
xor U13447 (N_13447,N_9803,N_10057);
nor U13448 (N_13448,N_7774,N_9118);
nand U13449 (N_13449,N_11449,N_7962);
xor U13450 (N_13450,N_8210,N_6740);
nor U13451 (N_13451,N_9127,N_11838);
xnor U13452 (N_13452,N_6417,N_7974);
or U13453 (N_13453,N_7204,N_10196);
xnor U13454 (N_13454,N_10475,N_7403);
xor U13455 (N_13455,N_9315,N_6726);
or U13456 (N_13456,N_8460,N_10813);
nor U13457 (N_13457,N_9179,N_8188);
and U13458 (N_13458,N_11321,N_6951);
nand U13459 (N_13459,N_8410,N_9792);
or U13460 (N_13460,N_10606,N_9195);
nor U13461 (N_13461,N_7391,N_11318);
xor U13462 (N_13462,N_7830,N_6423);
nor U13463 (N_13463,N_11274,N_9514);
and U13464 (N_13464,N_6942,N_6909);
xor U13465 (N_13465,N_11089,N_7734);
nand U13466 (N_13466,N_8954,N_6495);
or U13467 (N_13467,N_10840,N_8817);
nand U13468 (N_13468,N_7994,N_11173);
nand U13469 (N_13469,N_8844,N_11551);
nor U13470 (N_13470,N_11559,N_8960);
nand U13471 (N_13471,N_11000,N_9857);
and U13472 (N_13472,N_11808,N_8862);
nor U13473 (N_13473,N_7472,N_8110);
xnor U13474 (N_13474,N_8890,N_11993);
nor U13475 (N_13475,N_7640,N_10312);
nor U13476 (N_13476,N_11934,N_10336);
xor U13477 (N_13477,N_7718,N_9247);
nand U13478 (N_13478,N_6593,N_11923);
nor U13479 (N_13479,N_10353,N_6196);
nand U13480 (N_13480,N_6066,N_10181);
nand U13481 (N_13481,N_8926,N_8292);
nor U13482 (N_13482,N_10141,N_7705);
nand U13483 (N_13483,N_7488,N_10564);
xnor U13484 (N_13484,N_8338,N_6177);
and U13485 (N_13485,N_11719,N_10787);
or U13486 (N_13486,N_8270,N_7476);
nand U13487 (N_13487,N_11268,N_8888);
xnor U13488 (N_13488,N_9317,N_10741);
or U13489 (N_13489,N_7720,N_8988);
nand U13490 (N_13490,N_9477,N_8504);
and U13491 (N_13491,N_10459,N_8201);
xnor U13492 (N_13492,N_10952,N_10539);
or U13493 (N_13493,N_8551,N_6375);
nand U13494 (N_13494,N_8165,N_6249);
nand U13495 (N_13495,N_7411,N_6977);
or U13496 (N_13496,N_9978,N_8306);
or U13497 (N_13497,N_8681,N_11511);
and U13498 (N_13498,N_11928,N_8117);
and U13499 (N_13499,N_7757,N_9533);
xor U13500 (N_13500,N_11552,N_11644);
xor U13501 (N_13501,N_8300,N_11557);
xnor U13502 (N_13502,N_8923,N_9142);
xnor U13503 (N_13503,N_9941,N_8169);
xnor U13504 (N_13504,N_11312,N_10016);
nand U13505 (N_13505,N_10979,N_7934);
nand U13506 (N_13506,N_10445,N_11716);
or U13507 (N_13507,N_7512,N_10917);
nand U13508 (N_13508,N_6916,N_10507);
xor U13509 (N_13509,N_10659,N_9983);
nor U13510 (N_13510,N_9781,N_9727);
nor U13511 (N_13511,N_7321,N_8310);
and U13512 (N_13512,N_10133,N_9947);
nor U13513 (N_13513,N_10832,N_10033);
or U13514 (N_13514,N_7205,N_9432);
nand U13515 (N_13515,N_7234,N_8525);
nor U13516 (N_13516,N_10594,N_7632);
xor U13517 (N_13517,N_11731,N_10497);
xor U13518 (N_13518,N_8571,N_11779);
xor U13519 (N_13519,N_8238,N_11292);
or U13520 (N_13520,N_6541,N_7656);
nor U13521 (N_13521,N_7722,N_11707);
nand U13522 (N_13522,N_11885,N_10302);
xor U13523 (N_13523,N_11620,N_8362);
xnor U13524 (N_13524,N_8298,N_7447);
or U13525 (N_13525,N_8777,N_11743);
and U13526 (N_13526,N_10567,N_11632);
or U13527 (N_13527,N_6557,N_9600);
nand U13528 (N_13528,N_8705,N_7075);
nand U13529 (N_13529,N_11325,N_10101);
nand U13530 (N_13530,N_9360,N_8426);
xnor U13531 (N_13531,N_11283,N_9424);
and U13532 (N_13532,N_9210,N_8004);
nand U13533 (N_13533,N_9716,N_11396);
and U13534 (N_13534,N_10363,N_8251);
or U13535 (N_13535,N_7928,N_9933);
xor U13536 (N_13536,N_10762,N_10868);
and U13537 (N_13537,N_6517,N_8794);
or U13538 (N_13538,N_9665,N_11490);
xnor U13539 (N_13539,N_8422,N_9245);
and U13540 (N_13540,N_6709,N_11178);
nand U13541 (N_13541,N_11995,N_9476);
or U13542 (N_13542,N_6365,N_11116);
nor U13543 (N_13543,N_7630,N_8621);
or U13544 (N_13544,N_10670,N_10912);
nand U13545 (N_13545,N_11136,N_8729);
nor U13546 (N_13546,N_6601,N_6412);
xnor U13547 (N_13547,N_11444,N_8096);
or U13548 (N_13548,N_8629,N_11718);
nand U13549 (N_13549,N_10602,N_11447);
nand U13550 (N_13550,N_6445,N_7880);
xnor U13551 (N_13551,N_10723,N_6560);
xor U13552 (N_13552,N_8704,N_7006);
nor U13553 (N_13553,N_9039,N_6685);
nand U13554 (N_13554,N_6425,N_7187);
and U13555 (N_13555,N_7979,N_10026);
nand U13556 (N_13556,N_8652,N_11841);
and U13557 (N_13557,N_11920,N_8105);
xnor U13558 (N_13558,N_11221,N_7896);
or U13559 (N_13559,N_10571,N_10704);
nor U13560 (N_13560,N_10337,N_11051);
xor U13561 (N_13561,N_10963,N_11390);
xor U13562 (N_13562,N_11350,N_6344);
nand U13563 (N_13563,N_6169,N_10715);
nand U13564 (N_13564,N_6224,N_10310);
nand U13565 (N_13565,N_7745,N_6003);
nor U13566 (N_13566,N_9336,N_8303);
or U13567 (N_13567,N_9579,N_6703);
nor U13568 (N_13568,N_6007,N_9470);
or U13569 (N_13569,N_8039,N_8986);
or U13570 (N_13570,N_10753,N_9498);
and U13571 (N_13571,N_9794,N_9333);
nand U13572 (N_13572,N_10658,N_6990);
or U13573 (N_13573,N_10784,N_7294);
nand U13574 (N_13574,N_6401,N_9693);
xnor U13575 (N_13575,N_7936,N_11586);
nor U13576 (N_13576,N_8872,N_8366);
and U13577 (N_13577,N_6847,N_6176);
nand U13578 (N_13578,N_9202,N_6938);
or U13579 (N_13579,N_6534,N_9298);
and U13580 (N_13580,N_9720,N_10898);
and U13581 (N_13581,N_7428,N_8466);
nand U13582 (N_13582,N_7831,N_7001);
xor U13583 (N_13583,N_8402,N_8273);
xor U13584 (N_13584,N_7441,N_6349);
xor U13585 (N_13585,N_11759,N_7552);
nand U13586 (N_13586,N_6501,N_8602);
and U13587 (N_13587,N_6921,N_7258);
and U13588 (N_13588,N_8233,N_9095);
nor U13589 (N_13589,N_6402,N_10333);
nor U13590 (N_13590,N_11670,N_10130);
and U13591 (N_13591,N_10892,N_6522);
and U13592 (N_13592,N_7767,N_8250);
xor U13593 (N_13593,N_9377,N_7532);
or U13594 (N_13594,N_8727,N_10795);
nor U13595 (N_13595,N_10780,N_8297);
or U13596 (N_13596,N_10985,N_11289);
and U13597 (N_13597,N_7503,N_6870);
nor U13598 (N_13598,N_10596,N_9675);
nor U13599 (N_13599,N_7846,N_7620);
nor U13600 (N_13600,N_7629,N_6687);
or U13601 (N_13601,N_6956,N_8042);
xor U13602 (N_13602,N_9302,N_9076);
and U13603 (N_13603,N_11913,N_11435);
nor U13604 (N_13604,N_10134,N_6142);
and U13605 (N_13605,N_11679,N_7061);
nor U13606 (N_13606,N_8118,N_6413);
or U13607 (N_13607,N_10545,N_10883);
nor U13608 (N_13608,N_9090,N_7931);
nand U13609 (N_13609,N_6786,N_11434);
nand U13610 (N_13610,N_9034,N_10477);
and U13611 (N_13611,N_6483,N_9699);
or U13612 (N_13612,N_10568,N_10107);
nor U13613 (N_13613,N_10210,N_8302);
nand U13614 (N_13614,N_9048,N_10131);
and U13615 (N_13615,N_6185,N_9626);
nand U13616 (N_13616,N_9666,N_10802);
xor U13617 (N_13617,N_8578,N_8929);
nand U13618 (N_13618,N_11080,N_8855);
xor U13619 (N_13619,N_9056,N_9919);
xnor U13620 (N_13620,N_11781,N_9535);
and U13621 (N_13621,N_10355,N_11763);
xnor U13622 (N_13622,N_9944,N_10909);
and U13623 (N_13623,N_10065,N_10389);
nor U13624 (N_13624,N_9583,N_7838);
or U13625 (N_13625,N_8159,N_6233);
nor U13626 (N_13626,N_7573,N_11275);
nand U13627 (N_13627,N_7669,N_10217);
or U13628 (N_13628,N_6773,N_8124);
nand U13629 (N_13629,N_7142,N_6308);
xnor U13630 (N_13630,N_6061,N_6793);
nand U13631 (N_13631,N_9354,N_6369);
xnor U13632 (N_13632,N_11819,N_8342);
xnor U13633 (N_13633,N_10257,N_11436);
or U13634 (N_13634,N_9384,N_8425);
nor U13635 (N_13635,N_10127,N_9374);
nand U13636 (N_13636,N_6551,N_7871);
or U13637 (N_13637,N_11160,N_10988);
nor U13638 (N_13638,N_9207,N_7225);
and U13639 (N_13639,N_10505,N_8055);
nand U13640 (N_13640,N_11918,N_7109);
xor U13641 (N_13641,N_7520,N_8049);
nor U13642 (N_13642,N_11655,N_8021);
and U13643 (N_13643,N_6188,N_9128);
or U13644 (N_13644,N_11377,N_11897);
or U13645 (N_13645,N_11113,N_7701);
and U13646 (N_13646,N_11216,N_8502);
or U13647 (N_13647,N_7689,N_11004);
or U13648 (N_13648,N_10408,N_11832);
xnor U13649 (N_13649,N_7111,N_8644);
or U13650 (N_13650,N_8083,N_9051);
nand U13651 (N_13651,N_7340,N_6480);
and U13652 (N_13652,N_9860,N_8419);
xor U13653 (N_13653,N_7322,N_9807);
xnor U13654 (N_13654,N_6912,N_6183);
or U13655 (N_13655,N_8244,N_8054);
nor U13656 (N_13656,N_8177,N_6356);
nor U13657 (N_13657,N_11977,N_10447);
nor U13658 (N_13658,N_8218,N_11673);
nand U13659 (N_13659,N_7754,N_8645);
and U13660 (N_13660,N_9295,N_6610);
and U13661 (N_13661,N_6818,N_8076);
nor U13662 (N_13662,N_10488,N_7500);
or U13663 (N_13663,N_10905,N_6902);
and U13664 (N_13664,N_8095,N_8613);
or U13665 (N_13665,N_8725,N_7685);
nand U13666 (N_13666,N_7746,N_8784);
xor U13667 (N_13667,N_11714,N_9237);
xnor U13668 (N_13668,N_11515,N_7735);
or U13669 (N_13669,N_10872,N_9537);
or U13670 (N_13670,N_10823,N_11042);
or U13671 (N_13671,N_11912,N_7732);
nand U13672 (N_13672,N_8363,N_7719);
or U13673 (N_13673,N_9540,N_10359);
nor U13674 (N_13674,N_11407,N_7660);
xnor U13675 (N_13675,N_6895,N_11149);
nand U13676 (N_13676,N_6617,N_8984);
and U13677 (N_13677,N_6607,N_6655);
nor U13678 (N_13678,N_9980,N_11521);
or U13679 (N_13679,N_7575,N_8258);
or U13680 (N_13680,N_9301,N_10834);
nand U13681 (N_13681,N_10694,N_6021);
nand U13682 (N_13682,N_9689,N_8261);
nand U13683 (N_13683,N_8878,N_9394);
xor U13684 (N_13684,N_9146,N_6731);
nor U13685 (N_13685,N_10050,N_7466);
and U13686 (N_13686,N_7706,N_8384);
or U13687 (N_13687,N_10918,N_9553);
and U13688 (N_13688,N_8047,N_9770);
and U13689 (N_13689,N_9337,N_11421);
and U13690 (N_13690,N_11865,N_6738);
xor U13691 (N_13691,N_11970,N_9772);
xor U13692 (N_13692,N_8818,N_6811);
and U13693 (N_13693,N_7444,N_7172);
nor U13694 (N_13694,N_10623,N_8431);
nor U13695 (N_13695,N_9717,N_8810);
or U13696 (N_13696,N_9914,N_7131);
or U13697 (N_13697,N_9368,N_6766);
or U13698 (N_13698,N_10561,N_6387);
or U13699 (N_13699,N_9701,N_8823);
or U13700 (N_13700,N_11599,N_6757);
or U13701 (N_13701,N_7431,N_6111);
and U13702 (N_13702,N_8620,N_9844);
xor U13703 (N_13703,N_8391,N_8339);
nand U13704 (N_13704,N_10666,N_10227);
and U13705 (N_13705,N_9726,N_10383);
nand U13706 (N_13706,N_7904,N_11984);
nand U13707 (N_13707,N_7315,N_7889);
nand U13708 (N_13708,N_11770,N_11060);
xnor U13709 (N_13709,N_10246,N_11758);
and U13710 (N_13710,N_11228,N_6320);
or U13711 (N_13711,N_6359,N_6371);
nand U13712 (N_13712,N_9177,N_9135);
xor U13713 (N_13713,N_10690,N_9782);
nand U13714 (N_13714,N_10954,N_9762);
nor U13715 (N_13715,N_7143,N_11195);
nor U13716 (N_13716,N_6851,N_9886);
nand U13717 (N_13717,N_6751,N_9164);
nand U13718 (N_13718,N_10896,N_9485);
or U13719 (N_13719,N_6915,N_6555);
nor U13720 (N_13720,N_6384,N_7527);
and U13721 (N_13721,N_7384,N_8441);
and U13722 (N_13722,N_8838,N_9584);
nand U13723 (N_13723,N_7446,N_11491);
or U13724 (N_13724,N_7276,N_10783);
or U13725 (N_13725,N_9731,N_6094);
nor U13726 (N_13726,N_7893,N_7427);
nor U13727 (N_13727,N_8239,N_6756);
xor U13728 (N_13728,N_10298,N_8446);
xnor U13729 (N_13729,N_6976,N_10689);
nand U13730 (N_13730,N_8574,N_9018);
xor U13731 (N_13731,N_8564,N_6383);
nor U13732 (N_13732,N_10146,N_9366);
or U13733 (N_13733,N_8269,N_10682);
nand U13734 (N_13734,N_8349,N_9232);
nand U13735 (N_13735,N_7879,N_6025);
nor U13736 (N_13736,N_9089,N_10372);
nor U13737 (N_13737,N_11302,N_9697);
and U13738 (N_13738,N_10605,N_8682);
xor U13739 (N_13739,N_6642,N_11451);
nand U13740 (N_13740,N_8851,N_9393);
xnor U13741 (N_13741,N_9453,N_7248);
or U13742 (N_13742,N_8938,N_6649);
xor U13743 (N_13743,N_8702,N_11563);
xnor U13744 (N_13744,N_8092,N_6862);
and U13745 (N_13745,N_8272,N_6022);
or U13746 (N_13746,N_7473,N_10344);
and U13747 (N_13747,N_7167,N_11067);
xor U13748 (N_13748,N_11155,N_8301);
nor U13749 (N_13749,N_6431,N_11769);
nand U13750 (N_13750,N_10124,N_10455);
nor U13751 (N_13751,N_6753,N_10192);
or U13752 (N_13752,N_11999,N_11826);
xor U13753 (N_13753,N_11354,N_11375);
xor U13754 (N_13754,N_8935,N_9401);
and U13755 (N_13755,N_8957,N_11508);
and U13756 (N_13756,N_6663,N_6874);
nor U13757 (N_13757,N_7710,N_11517);
or U13758 (N_13758,N_9431,N_11086);
xor U13759 (N_13759,N_9585,N_9667);
and U13760 (N_13760,N_10457,N_10686);
nor U13761 (N_13761,N_9014,N_6582);
and U13762 (N_13762,N_9599,N_7342);
xnor U13763 (N_13763,N_11676,N_11813);
or U13764 (N_13764,N_7683,N_9163);
and U13765 (N_13765,N_11440,N_6030);
nor U13766 (N_13766,N_11904,N_10749);
nor U13767 (N_13767,N_9275,N_8005);
nor U13768 (N_13768,N_11704,N_10091);
or U13769 (N_13769,N_9239,N_9572);
and U13770 (N_13770,N_6033,N_6622);
xor U13771 (N_13771,N_6444,N_6438);
xor U13772 (N_13772,N_6235,N_7907);
nand U13773 (N_13773,N_7291,N_8959);
xnor U13774 (N_13774,N_10085,N_8871);
nand U13775 (N_13775,N_10885,N_10317);
xnor U13776 (N_13776,N_7967,N_8260);
xnor U13777 (N_13777,N_10229,N_7259);
or U13778 (N_13778,N_11834,N_11794);
or U13779 (N_13779,N_8100,N_6545);
and U13780 (N_13780,N_10645,N_7747);
nand U13781 (N_13781,N_9440,N_11199);
nor U13782 (N_13782,N_6045,N_11497);
nor U13783 (N_13783,N_9843,N_9566);
nand U13784 (N_13784,N_8857,N_8388);
xnor U13785 (N_13785,N_10537,N_6339);
nand U13786 (N_13786,N_9233,N_9630);
and U13787 (N_13787,N_10978,N_8367);
nor U13788 (N_13788,N_11353,N_9304);
xor U13789 (N_13789,N_11662,N_10675);
or U13790 (N_13790,N_9227,N_8019);
and U13791 (N_13791,N_6550,N_11728);
nor U13792 (N_13792,N_10777,N_6882);
and U13793 (N_13793,N_11806,N_7627);
nor U13794 (N_13794,N_7219,N_7511);
or U13795 (N_13795,N_9066,N_10098);
and U13796 (N_13796,N_6244,N_7823);
xor U13797 (N_13797,N_6889,N_7865);
or U13798 (N_13798,N_10164,N_7964);
or U13799 (N_13799,N_9043,N_11194);
or U13800 (N_13800,N_9350,N_7126);
xor U13801 (N_13801,N_10836,N_7211);
or U13802 (N_13802,N_10590,N_10970);
xnor U13803 (N_13803,N_10012,N_11535);
nand U13804 (N_13804,N_7538,N_9098);
nor U13805 (N_13805,N_10522,N_6482);
or U13806 (N_13806,N_9870,N_10222);
and U13807 (N_13807,N_10585,N_10206);
nor U13808 (N_13808,N_9412,N_10187);
nand U13809 (N_13809,N_11591,N_7997);
nor U13810 (N_13810,N_9872,N_9755);
nand U13811 (N_13811,N_7455,N_6580);
or U13812 (N_13812,N_10325,N_10392);
nand U13813 (N_13813,N_10188,N_8819);
nor U13814 (N_13814,N_6599,N_10820);
xor U13815 (N_13815,N_10039,N_9443);
or U13816 (N_13816,N_9054,N_11605);
xnor U13817 (N_13817,N_6190,N_8750);
and U13818 (N_13818,N_8885,N_10526);
xnor U13819 (N_13819,N_8171,N_10508);
or U13820 (N_13820,N_6759,N_6802);
nor U13821 (N_13821,N_10598,N_7040);
xor U13822 (N_13822,N_11787,N_10243);
or U13823 (N_13823,N_11288,N_11076);
and U13824 (N_13824,N_8856,N_9964);
xnor U13825 (N_13825,N_6529,N_10038);
and U13826 (N_13826,N_7308,N_7354);
nand U13827 (N_13827,N_7739,N_8481);
xor U13828 (N_13828,N_11595,N_9067);
or U13829 (N_13829,N_7422,N_6844);
nand U13830 (N_13830,N_8434,N_11442);
nor U13831 (N_13831,N_8939,N_9915);
nand U13832 (N_13832,N_6039,N_6654);
and U13833 (N_13833,N_9522,N_8605);
xor U13834 (N_13834,N_8335,N_9073);
or U13835 (N_13835,N_9087,N_11693);
nand U13836 (N_13836,N_9042,N_6162);
or U13837 (N_13837,N_11823,N_7618);
nand U13838 (N_13838,N_9847,N_11750);
nor U13839 (N_13839,N_8079,N_7332);
nor U13840 (N_13840,N_9362,N_6536);
and U13841 (N_13841,N_8442,N_8654);
or U13842 (N_13842,N_8311,N_10829);
or U13843 (N_13843,N_6437,N_7325);
nand U13844 (N_13844,N_11046,N_10161);
or U13845 (N_13845,N_8150,N_11429);
and U13846 (N_13846,N_6530,N_9376);
nand U13847 (N_13847,N_7803,N_11987);
xor U13848 (N_13848,N_6439,N_9289);
and U13849 (N_13849,N_9081,N_8175);
nand U13850 (N_13850,N_11531,N_7777);
nor U13851 (N_13851,N_8475,N_11391);
or U13852 (N_13852,N_10492,N_8666);
nand U13853 (N_13853,N_9496,N_7941);
nor U13854 (N_13854,N_10255,N_9706);
and U13855 (N_13855,N_10662,N_7886);
and U13856 (N_13856,N_9216,N_10639);
xor U13857 (N_13857,N_6561,N_7071);
and U13858 (N_13858,N_10714,N_10468);
or U13859 (N_13859,N_7744,N_11840);
nand U13860 (N_13860,N_11548,N_10184);
or U13861 (N_13861,N_6458,N_6419);
nor U13862 (N_13862,N_11789,N_11756);
or U13863 (N_13863,N_10166,N_8046);
xnor U13864 (N_13864,N_10470,N_7901);
nand U13865 (N_13865,N_7349,N_6035);
or U13866 (N_13866,N_11203,N_6267);
or U13867 (N_13867,N_8077,N_9673);
nand U13868 (N_13868,N_7783,N_7781);
nand U13869 (N_13869,N_7897,N_7310);
and U13870 (N_13870,N_9904,N_11700);
or U13871 (N_13871,N_9676,N_10550);
nor U13872 (N_13872,N_10858,N_7555);
nand U13873 (N_13873,N_9788,N_10735);
or U13874 (N_13874,N_8346,N_7115);
and U13875 (N_13875,N_10653,N_6849);
nor U13876 (N_13876,N_10640,N_8423);
nand U13877 (N_13877,N_9526,N_8911);
and U13878 (N_13878,N_11330,N_6544);
or U13879 (N_13879,N_8513,N_11126);
nand U13880 (N_13880,N_7678,N_9962);
xnor U13881 (N_13881,N_8399,N_7696);
xor U13882 (N_13882,N_7533,N_6594);
nor U13883 (N_13883,N_11598,N_10055);
and U13884 (N_13884,N_9934,N_9812);
nand U13885 (N_13885,N_9823,N_9516);
xnor U13886 (N_13886,N_10052,N_10301);
nor U13887 (N_13887,N_6957,N_7860);
and U13888 (N_13888,N_8268,N_7477);
xnor U13889 (N_13889,N_9750,N_7499);
nor U13890 (N_13890,N_9225,N_6652);
and U13891 (N_13891,N_7256,N_11764);
nand U13892 (N_13892,N_8641,N_10466);
or U13893 (N_13893,N_7005,N_6089);
and U13894 (N_13894,N_7815,N_7101);
or U13895 (N_13895,N_11944,N_8565);
nand U13896 (N_13896,N_8345,N_9447);
and U13897 (N_13897,N_7381,N_7336);
nand U13898 (N_13898,N_11024,N_6314);
and U13899 (N_13899,N_9556,N_6187);
nand U13900 (N_13900,N_11171,N_9172);
or U13901 (N_13901,N_9833,N_10162);
nand U13902 (N_13902,N_11281,N_10129);
nor U13903 (N_13903,N_6799,N_8532);
or U13904 (N_13904,N_7216,N_10767);
nor U13905 (N_13905,N_8936,N_10195);
or U13906 (N_13906,N_8636,N_7652);
and U13907 (N_13907,N_9641,N_10132);
xor U13908 (N_13908,N_11480,N_8074);
xnor U13909 (N_13909,N_11172,N_7884);
nand U13910 (N_13910,N_8912,N_10110);
and U13911 (N_13911,N_11477,N_9133);
nand U13912 (N_13912,N_11638,N_7084);
or U13913 (N_13913,N_9093,N_7497);
nor U13914 (N_13914,N_7416,N_8740);
nor U13915 (N_13915,N_11028,N_7969);
and U13916 (N_13916,N_7016,N_10546);
nor U13917 (N_13917,N_6297,N_9894);
nor U13918 (N_13918,N_11997,N_11733);
nor U13919 (N_13919,N_11083,N_8228);
nor U13920 (N_13920,N_7567,N_9000);
or U13921 (N_13921,N_9129,N_6334);
and U13922 (N_13922,N_11637,N_6651);
nand U13923 (N_13923,N_7456,N_6116);
nor U13924 (N_13924,N_11573,N_10712);
xor U13925 (N_13925,N_9779,N_10631);
or U13926 (N_13926,N_9392,N_7817);
xor U13927 (N_13927,N_7647,N_8385);
or U13928 (N_13928,N_8107,N_6415);
and U13929 (N_13929,N_6708,N_11263);
xnor U13930 (N_13930,N_11488,N_7692);
nand U13931 (N_13931,N_11957,N_9822);
nor U13932 (N_13932,N_6919,N_7770);
nor U13933 (N_13933,N_11744,N_7530);
nor U13934 (N_13934,N_9194,N_6932);
nor U13935 (N_13935,N_8334,N_11286);
or U13936 (N_13936,N_7704,N_8568);
xnor U13937 (N_13937,N_8977,N_11965);
or U13938 (N_13938,N_8436,N_11975);
and U13939 (N_13939,N_7711,N_7768);
or U13940 (N_13940,N_10297,N_8199);
nor U13941 (N_13941,N_9152,N_11636);
nand U13942 (N_13942,N_11174,N_6791);
and U13943 (N_13943,N_9258,N_11352);
xnor U13944 (N_13944,N_9047,N_7193);
nor U13945 (N_13945,N_8892,N_6407);
and U13946 (N_13946,N_11674,N_10880);
or U13947 (N_13947,N_11747,N_9868);
or U13948 (N_13948,N_7202,N_11416);
xnor U13949 (N_13949,N_8883,N_7292);
nor U13950 (N_13950,N_9989,N_8111);
nand U13951 (N_13951,N_10169,N_6079);
nand U13952 (N_13952,N_6100,N_6965);
xnor U13953 (N_13953,N_8902,N_8489);
or U13954 (N_13954,N_6273,N_6129);
and U13955 (N_13955,N_11600,N_7091);
and U13956 (N_13956,N_7699,N_9351);
or U13957 (N_13957,N_10469,N_7534);
and U13958 (N_13958,N_9660,N_8480);
nor U13959 (N_13959,N_11273,N_11507);
xnor U13960 (N_13960,N_8193,N_11401);
and U13961 (N_13961,N_9015,N_8906);
and U13962 (N_13962,N_11604,N_11165);
and U13963 (N_13963,N_8594,N_8142);
xnor U13964 (N_13964,N_11418,N_10324);
and U13965 (N_13965,N_7988,N_7776);
nor U13966 (N_13966,N_7176,N_7051);
or U13967 (N_13967,N_6705,N_9917);
and U13968 (N_13968,N_6518,N_11106);
and U13969 (N_13969,N_7169,N_6272);
or U13970 (N_13970,N_11658,N_10441);
nand U13971 (N_13971,N_6819,N_10454);
xnor U13972 (N_13972,N_8259,N_8206);
or U13973 (N_13973,N_6232,N_8290);
nor U13974 (N_13974,N_9395,N_7104);
nand U13975 (N_13975,N_8445,N_9815);
nand U13976 (N_13976,N_7926,N_7459);
nor U13977 (N_13977,N_9951,N_9966);
and U13978 (N_13978,N_9845,N_6008);
nor U13979 (N_13979,N_8488,N_7356);
and U13980 (N_13980,N_11157,N_7070);
nor U13981 (N_13981,N_6980,N_7468);
xor U13982 (N_13982,N_6632,N_10398);
and U13983 (N_13983,N_9679,N_8494);
xor U13984 (N_13984,N_9484,N_8178);
nor U13985 (N_13985,N_9286,N_8316);
and U13986 (N_13986,N_6292,N_7430);
or U13987 (N_13987,N_11243,N_7698);
or U13988 (N_13988,N_11010,N_10062);
xor U13989 (N_13989,N_10925,N_7074);
or U13990 (N_13990,N_6906,N_6454);
xnor U13991 (N_13991,N_8555,N_8543);
nand U13992 (N_13992,N_9879,N_8069);
xnor U13993 (N_13993,N_9810,N_8352);
nor U13994 (N_13994,N_10070,N_8072);
xor U13995 (N_13995,N_6745,N_6809);
or U13996 (N_13996,N_6488,N_10910);
and U13997 (N_13997,N_10149,N_8990);
nand U13998 (N_13998,N_6027,N_10914);
nand U13999 (N_13999,N_6879,N_11815);
or U14000 (N_14000,N_6472,N_7766);
nand U14001 (N_14001,N_11994,N_10900);
and U14002 (N_14002,N_10719,N_8529);
xor U14003 (N_14003,N_8985,N_9970);
or U14004 (N_14004,N_10794,N_11125);
and U14005 (N_14005,N_9458,N_8189);
nor U14006 (N_14006,N_6213,N_11607);
or U14007 (N_14007,N_6210,N_8088);
xnor U14008 (N_14008,N_9203,N_7664);
and U14009 (N_14009,N_11047,N_7319);
and U14010 (N_14010,N_8470,N_8089);
nor U14011 (N_14011,N_6151,N_8255);
and U14012 (N_14012,N_8607,N_8835);
and U14013 (N_14013,N_8440,N_11169);
xnor U14014 (N_14014,N_10343,N_7206);
xor U14015 (N_14015,N_6742,N_10178);
and U14016 (N_14016,N_8703,N_8772);
xor U14017 (N_14017,N_7274,N_7457);
and U14018 (N_14018,N_11464,N_7955);
and U14019 (N_14019,N_8506,N_9184);
nand U14020 (N_14020,N_9370,N_11355);
or U14021 (N_14021,N_8398,N_8014);
and U14022 (N_14022,N_6470,N_11917);
or U14023 (N_14023,N_10601,N_7079);
and U14024 (N_14024,N_7723,N_7663);
nor U14025 (N_14025,N_8331,N_8816);
xnor U14026 (N_14026,N_7845,N_8464);
nor U14027 (N_14027,N_8029,N_9408);
or U14028 (N_14028,N_6577,N_7424);
and U14029 (N_14029,N_9816,N_8262);
and U14030 (N_14030,N_6824,N_6715);
and U14031 (N_14031,N_11448,N_8176);
nor U14032 (N_14032,N_11259,N_6447);
nand U14033 (N_14033,N_7913,N_10578);
nor U14034 (N_14034,N_8377,N_7132);
nand U14035 (N_14035,N_9544,N_10214);
nor U14036 (N_14036,N_10512,N_11846);
and U14037 (N_14037,N_9460,N_8376);
and U14038 (N_14038,N_10513,N_11869);
nor U14039 (N_14039,N_7353,N_9916);
xor U14040 (N_14040,N_9813,N_9984);
and U14041 (N_14041,N_9607,N_11487);
or U14042 (N_14042,N_11973,N_10838);
xor U14043 (N_14043,N_10292,N_10944);
nand U14044 (N_14044,N_9571,N_7673);
xor U14045 (N_14045,N_8443,N_9378);
nor U14046 (N_14046,N_10582,N_10862);
and U14047 (N_14047,N_10018,N_10845);
nor U14048 (N_14048,N_6535,N_11458);
xor U14049 (N_14049,N_8536,N_7145);
nand U14050 (N_14050,N_8941,N_7140);
nor U14051 (N_14051,N_7306,N_10969);
nor U14052 (N_14052,N_10370,N_10811);
or U14053 (N_14053,N_8781,N_7507);
and U14054 (N_14054,N_10403,N_9898);
or U14055 (N_14055,N_11861,N_9713);
nand U14056 (N_14056,N_8406,N_11501);
or U14057 (N_14057,N_10493,N_10314);
xnor U14058 (N_14058,N_11206,N_10527);
or U14059 (N_14059,N_7873,N_9730);
nor U14060 (N_14060,N_10613,N_10620);
nor U14061 (N_14061,N_7761,N_9800);
nor U14062 (N_14062,N_7366,N_11839);
nor U14063 (N_14063,N_11880,N_11430);
xor U14064 (N_14064,N_7413,N_9267);
and U14065 (N_14065,N_7522,N_9132);
nand U14066 (N_14066,N_6229,N_7201);
or U14067 (N_14067,N_9421,N_11796);
or U14068 (N_14068,N_10104,N_9903);
nand U14069 (N_14069,N_11847,N_9846);
nand U14070 (N_14070,N_11509,N_8721);
or U14071 (N_14071,N_8635,N_10557);
xor U14072 (N_14072,N_11201,N_10163);
and U14073 (N_14073,N_11188,N_9606);
nor U14074 (N_14074,N_6848,N_9897);
and U14075 (N_14075,N_9084,N_6770);
nand U14076 (N_14076,N_10709,N_11276);
or U14077 (N_14077,N_10409,N_6343);
and U14078 (N_14078,N_9658,N_6748);
or U14079 (N_14079,N_11863,N_6280);
nand U14080 (N_14080,N_9627,N_8833);
nand U14081 (N_14081,N_9415,N_7769);
xor U14082 (N_14082,N_8041,N_7866);
xnor U14083 (N_14083,N_8050,N_10971);
and U14084 (N_14084,N_10589,N_7611);
and U14085 (N_14085,N_8449,N_10774);
or U14086 (N_14086,N_11618,N_8775);
nor U14087 (N_14087,N_11483,N_6331);
and U14088 (N_14088,N_7782,N_11428);
nand U14089 (N_14089,N_11580,N_7543);
nand U14090 (N_14090,N_6794,N_11541);
nand U14091 (N_14091,N_11005,N_9777);
nor U14092 (N_14092,N_7972,N_8684);
xnor U14093 (N_14093,N_6355,N_7014);
xor U14094 (N_14094,N_6755,N_7836);
nor U14095 (N_14095,N_8528,N_7080);
nor U14096 (N_14096,N_8994,N_7327);
xnor U14097 (N_14097,N_11265,N_11329);
nor U14098 (N_14098,N_10806,N_11625);
xor U14099 (N_14099,N_7804,N_8283);
or U14100 (N_14100,N_6317,N_6291);
or U14101 (N_14101,N_6476,N_7587);
or U14102 (N_14102,N_7634,N_6441);
nor U14103 (N_14103,N_6148,N_6635);
xor U14104 (N_14104,N_10935,N_11306);
xor U14105 (N_14105,N_8670,N_6776);
nor U14106 (N_14106,N_11317,N_10853);
xnor U14107 (N_14107,N_11629,N_6624);
xor U14108 (N_14108,N_11761,N_11090);
nand U14109 (N_14109,N_10773,N_11474);
xor U14110 (N_14110,N_11585,N_6511);
xor U14111 (N_14111,N_10203,N_9819);
or U14112 (N_14112,N_6348,N_9019);
nand U14113 (N_14113,N_7015,N_6436);
xnor U14114 (N_14114,N_10702,N_11550);
xnor U14115 (N_14115,N_11405,N_8168);
nand U14116 (N_14116,N_8631,N_11493);
or U14117 (N_14117,N_6078,N_9853);
or U14118 (N_14118,N_7209,N_9725);
or U14119 (N_14119,N_9576,N_6508);
xnor U14120 (N_14120,N_9165,N_7709);
nor U14121 (N_14121,N_10473,N_10691);
xnor U14122 (N_14122,N_10583,N_11164);
nor U14123 (N_14123,N_6758,N_10586);
xor U14124 (N_14124,N_10194,N_8373);
nand U14125 (N_14125,N_7493,N_11140);
and U14126 (N_14126,N_8197,N_10923);
or U14127 (N_14127,N_10258,N_6350);
xnor U14128 (N_14128,N_10485,N_7790);
or U14129 (N_14129,N_11386,N_10687);
and U14130 (N_14130,N_6639,N_8889);
nor U14131 (N_14131,N_9517,N_10785);
and U14132 (N_14132,N_9880,N_7791);
nand U14133 (N_14133,N_9855,N_7119);
xor U14134 (N_14134,N_11079,N_7876);
and U14135 (N_14135,N_10138,N_10261);
and U14136 (N_14136,N_6962,N_8782);
xor U14137 (N_14137,N_7049,N_9848);
nand U14138 (N_14138,N_9531,N_7182);
nor U14139 (N_14139,N_7326,N_11512);
nor U14140 (N_14140,N_11379,N_7951);
or U14141 (N_14141,N_10236,N_10078);
nand U14142 (N_14142,N_8495,N_7350);
and U14143 (N_14143,N_8790,N_7801);
nand U14144 (N_14144,N_9101,N_9107);
xnor U14145 (N_14145,N_7106,N_9899);
nor U14146 (N_14146,N_9168,N_6829);
or U14147 (N_14147,N_8144,N_10433);
nand U14148 (N_14148,N_11114,N_8421);
and U14149 (N_14149,N_10941,N_11936);
xor U14150 (N_14150,N_8891,N_10082);
or U14151 (N_14151,N_6101,N_10529);
xnor U14152 (N_14152,N_11097,N_7121);
nand U14153 (N_14153,N_10160,N_10121);
nand U14154 (N_14154,N_11646,N_10759);
or U14155 (N_14155,N_7919,N_9839);
nor U14156 (N_14156,N_10358,N_6548);
or U14157 (N_14157,N_6107,N_8240);
and U14158 (N_14158,N_8527,N_7645);
xor U14159 (N_14159,N_6512,N_9668);
xor U14160 (N_14160,N_9306,N_8330);
xnor U14161 (N_14161,N_11167,N_11788);
or U14162 (N_14162,N_7943,N_11445);
nor U14163 (N_14163,N_8119,N_10247);
or U14164 (N_14164,N_7950,N_9004);
xor U14165 (N_14165,N_6925,N_8868);
or U14166 (N_14166,N_8032,N_9798);
xnor U14167 (N_14167,N_8925,N_10843);
or U14168 (N_14168,N_11726,N_10086);
nand U14169 (N_14169,N_11460,N_10270);
nor U14170 (N_14170,N_8839,N_11735);
nand U14171 (N_14171,N_11158,N_7008);
xnor U14172 (N_14172,N_10688,N_6941);
and U14173 (N_14173,N_11270,N_9862);
xnor U14174 (N_14174,N_11014,N_8485);
and U14175 (N_14175,N_9968,N_11952);
nor U14176 (N_14176,N_8459,N_10728);
nor U14177 (N_14177,N_6764,N_11933);
nor U14178 (N_14178,N_11762,N_6000);
nand U14179 (N_14179,N_9642,N_10371);
nand U14180 (N_14180,N_8884,N_10044);
nor U14181 (N_14181,N_8026,N_8143);
nand U14182 (N_14182,N_7007,N_7792);
nand U14183 (N_14183,N_6587,N_8886);
and U14184 (N_14184,N_11564,N_9450);
xnor U14185 (N_14185,N_6669,N_10145);
nor U14186 (N_14186,N_7578,N_11835);
or U14187 (N_14187,N_9945,N_6877);
xnor U14188 (N_14188,N_8893,N_8075);
or U14189 (N_14189,N_10030,N_8448);
xor U14190 (N_14190,N_6883,N_7094);
xor U14191 (N_14191,N_6542,N_9538);
xor U14192 (N_14192,N_9257,N_6667);
or U14193 (N_14193,N_7717,N_11269);
and U14194 (N_14194,N_10661,N_6775);
and U14195 (N_14195,N_11896,N_7382);
nand U14196 (N_14196,N_9463,N_6506);
nand U14197 (N_14197,N_11134,N_8022);
xnor U14198 (N_14198,N_7486,N_7053);
nand U14199 (N_14199,N_11122,N_6840);
or U14200 (N_14200,N_9339,N_11120);
or U14201 (N_14201,N_8017,N_11657);
or U14202 (N_14202,N_7425,N_11339);
and U14203 (N_14203,N_11041,N_11516);
or U14204 (N_14204,N_8557,N_9390);
nand U14205 (N_14205,N_9012,N_7448);
and U14206 (N_14206,N_11230,N_10494);
nand U14207 (N_14207,N_9612,N_7251);
nor U14208 (N_14208,N_7271,N_6754);
or U14209 (N_14209,N_11857,N_10135);
nor U14210 (N_14210,N_8587,N_10782);
or U14211 (N_14211,N_10603,N_11443);
or U14212 (N_14212,N_11049,N_10068);
xor U14213 (N_14213,N_10202,N_8895);
or U14214 (N_14214,N_10219,N_6878);
or U14215 (N_14215,N_10980,N_11929);
nor U14216 (N_14216,N_11044,N_8106);
xnor U14217 (N_14217,N_6009,N_10879);
xor U14218 (N_14218,N_9486,N_11562);
and U14219 (N_14219,N_9640,N_8531);
nand U14220 (N_14220,N_10231,N_6784);
xor U14221 (N_14221,N_7787,N_6042);
xnor U14222 (N_14222,N_9344,N_8430);
and U14223 (N_14223,N_10059,N_10924);
xor U14224 (N_14224,N_11313,N_7516);
or U14225 (N_14225,N_6131,N_11333);
or U14226 (N_14226,N_7334,N_11549);
nand U14227 (N_14227,N_7593,N_11979);
or U14228 (N_14228,N_10197,N_9922);
nor U14229 (N_14229,N_7375,N_9732);
and U14230 (N_14230,N_10021,N_6917);
xnor U14231 (N_14231,N_10758,N_10300);
nand U14232 (N_14232,N_11384,N_9221);
nor U14233 (N_14233,N_8537,N_7637);
or U14234 (N_14234,N_11827,N_7019);
nand U14235 (N_14235,N_6140,N_6460);
and U14236 (N_14236,N_7298,N_7288);
xor U14237 (N_14237,N_6549,N_6154);
or U14238 (N_14238,N_6093,N_10990);
or U14239 (N_14239,N_7390,N_8435);
nand U14240 (N_14240,N_8086,N_11622);
nor U14241 (N_14241,N_11525,N_8360);
or U14242 (N_14242,N_7569,N_10125);
nor U14243 (N_14243,N_11181,N_7405);
xnor U14244 (N_14244,N_10649,N_7691);
and U14245 (N_14245,N_11492,N_9023);
nor U14246 (N_14246,N_10172,N_8293);
xnor U14247 (N_14247,N_10865,N_9182);
nand U14248 (N_14248,N_9497,N_11363);
or U14249 (N_14249,N_10081,N_8325);
and U14250 (N_14250,N_9595,N_10863);
and U14251 (N_14251,N_8712,N_11760);
or U14252 (N_14252,N_10429,N_10699);
or U14253 (N_14253,N_9313,N_11678);
or U14254 (N_14254,N_6896,N_11358);
and U14255 (N_14255,N_7229,N_8538);
nor U14256 (N_14256,N_11239,N_10436);
and U14257 (N_14257,N_10092,N_10981);
xnor U14258 (N_14258,N_7289,N_11615);
nor U14259 (N_14259,N_9288,N_11513);
or U14260 (N_14260,N_11343,N_9180);
nor U14261 (N_14261,N_8655,N_8572);
xor U14262 (N_14262,N_9359,N_6733);
nor U14263 (N_14263,N_9907,N_10664);
nor U14264 (N_14264,N_9560,N_6590);
and U14265 (N_14265,N_6695,N_11334);
xor U14266 (N_14266,N_6991,N_11196);
or U14267 (N_14267,N_11266,N_6396);
or U14268 (N_14268,N_7033,N_10973);
and U14269 (N_14269,N_6888,N_8534);
or U14270 (N_14270,N_10046,N_6936);
xor U14271 (N_14271,N_8213,N_7433);
xor U14272 (N_14272,N_6304,N_9564);
or U14273 (N_14273,N_11692,N_10809);
and U14274 (N_14274,N_8044,N_9581);
nand U14275 (N_14275,N_7485,N_6785);
nor U14276 (N_14276,N_6691,N_9357);
or U14277 (N_14277,N_6527,N_10260);
nor U14278 (N_14278,N_8085,N_7452);
nand U14279 (N_14279,N_11603,N_6752);
and U14280 (N_14280,N_9545,N_9628);
nor U14281 (N_14281,N_11753,N_9300);
or U14282 (N_14282,N_11456,N_7595);
or U14283 (N_14283,N_9464,N_6999);
xor U14284 (N_14284,N_8256,N_8999);
nand U14285 (N_14285,N_7282,N_9707);
and U14286 (N_14286,N_6972,N_6399);
or U14287 (N_14287,N_11011,N_7067);
or U14288 (N_14288,N_11905,N_11144);
and U14289 (N_14289,N_6795,N_9342);
nor U14290 (N_14290,N_9830,N_7564);
and U14291 (N_14291,N_11623,N_11879);
xor U14292 (N_14292,N_10611,N_11197);
or U14293 (N_14293,N_11696,N_6381);
or U14294 (N_14294,N_11217,N_9059);
xor U14295 (N_14295,N_10577,N_7163);
nand U14296 (N_14296,N_7822,N_8530);
nor U14297 (N_14297,N_9316,N_10352);
and U14298 (N_14298,N_7840,N_9900);
nor U14299 (N_14299,N_10349,N_11135);
and U14300 (N_14300,N_6245,N_7159);
nor U14301 (N_14301,N_10822,N_8403);
and U14302 (N_14302,N_10967,N_9219);
xor U14303 (N_14303,N_9086,N_10111);
nor U14304 (N_14304,N_7404,N_8699);
nand U14305 (N_14305,N_8715,N_11257);
or U14306 (N_14306,N_7714,N_7386);
xnor U14307 (N_14307,N_10268,N_7238);
and U14308 (N_14308,N_8958,N_11946);
and U14309 (N_14309,N_9407,N_10097);
nor U14310 (N_14310,N_7626,N_10089);
or U14311 (N_14311,N_6414,N_7506);
xor U14312 (N_14312,N_8901,N_11298);
or U14313 (N_14313,N_10027,N_11634);
and U14314 (N_14314,N_6531,N_11361);
xnor U14315 (N_14315,N_8133,N_8497);
nand U14316 (N_14316,N_6641,N_10851);
xor U14317 (N_14317,N_10580,N_10919);
or U14318 (N_14318,N_11895,N_10233);
nand U14319 (N_14319,N_11454,N_10703);
nand U14320 (N_14320,N_8731,N_6076);
nor U14321 (N_14321,N_9688,N_10185);
nand U14322 (N_14322,N_6810,N_8668);
nand U14323 (N_14323,N_9403,N_10673);
xnor U14324 (N_14324,N_7128,N_7147);
and U14325 (N_14325,N_7668,N_8992);
xnor U14326 (N_14326,N_8827,N_7760);
nor U14327 (N_14327,N_11368,N_6220);
nor U14328 (N_14328,N_7228,N_9277);
xor U14329 (N_14329,N_11748,N_10964);
or U14330 (N_14330,N_9684,N_7594);
xor U14331 (N_14331,N_11026,N_7266);
nand U14332 (N_14332,N_7280,N_7675);
nor U14333 (N_14333,N_10480,N_10153);
nand U14334 (N_14334,N_10679,N_11754);
nor U14335 (N_14335,N_7484,N_11404);
nand U14336 (N_14336,N_9255,N_11359);
and U14337 (N_14337,N_7674,N_6939);
nor U14338 (N_14338,N_7284,N_11446);
xor U14339 (N_14339,N_6070,N_9231);
or U14340 (N_14340,N_11690,N_10218);
or U14341 (N_14341,N_6074,N_9714);
nor U14342 (N_14342,N_10713,N_10275);
nand U14343 (N_14343,N_11237,N_6963);
nand U14344 (N_14344,N_6080,N_11723);
xnor U14345 (N_14345,N_8647,N_9804);
nand U14346 (N_14346,N_9521,N_10932);
xor U14347 (N_14347,N_7540,N_11153);
nand U14348 (N_14348,N_8222,N_9829);
nand U14349 (N_14349,N_9591,N_11927);
and U14350 (N_14350,N_6790,N_9137);
or U14351 (N_14351,N_6493,N_10801);
nor U14352 (N_14352,N_9644,N_6992);
nand U14353 (N_14353,N_9176,N_11685);
xnor U14354 (N_14354,N_11111,N_6166);
nand U14355 (N_14355,N_6656,N_7521);
xor U14356 (N_14356,N_7799,N_11320);
and U14357 (N_14357,N_10183,N_11130);
xor U14358 (N_14358,N_10815,N_11209);
and U14359 (N_14359,N_9112,N_10599);
and U14360 (N_14360,N_9071,N_9025);
nor U14361 (N_14361,N_10140,N_8546);
xor U14362 (N_14362,N_9937,N_10072);
or U14363 (N_14363,N_11039,N_7843);
xor U14364 (N_14364,N_7653,N_10727);
xnor U14365 (N_14365,N_8263,N_10738);
nand U14366 (N_14366,N_9790,N_7236);
nand U14367 (N_14367,N_8104,N_9506);
nor U14368 (N_14368,N_9672,N_10750);
and U14369 (N_14369,N_7571,N_8134);
nand U14370 (N_14370,N_8671,N_11870);
or U14371 (N_14371,N_11640,N_8170);
or U14372 (N_14372,N_7129,N_7965);
xor U14373 (N_14373,N_9690,N_11427);
nand U14374 (N_14374,N_8753,N_8295);
nand U14375 (N_14375,N_9159,N_6645);
or U14376 (N_14376,N_6064,N_6421);
or U14377 (N_14377,N_9252,N_9960);
xor U14378 (N_14378,N_8963,N_6195);
nor U14379 (N_14379,N_7867,N_7160);
or U14380 (N_14380,N_7592,N_10123);
and U14381 (N_14381,N_11765,N_7916);
and U14382 (N_14382,N_10792,N_6722);
nor U14383 (N_14383,N_8242,N_10953);
and U14384 (N_14384,N_10061,N_10365);
nor U14385 (N_14385,N_11151,N_11649);
nand U14386 (N_14386,N_10745,N_8313);
or U14387 (N_14387,N_11382,N_8745);
and U14388 (N_14388,N_7200,N_6516);
and U14389 (N_14389,N_11862,N_10176);
xnor U14390 (N_14390,N_7483,N_9080);
nand U14391 (N_14391,N_11642,N_11971);
nand U14392 (N_14392,N_7199,N_6638);
nand U14393 (N_14393,N_9986,N_7223);
nor U14394 (N_14394,N_11593,N_11468);
xnor U14395 (N_14395,N_11037,N_6821);
and U14396 (N_14396,N_10025,N_7686);
xor U14397 (N_14397,N_10766,N_9113);
nand U14398 (N_14398,N_7054,N_6228);
xor U14399 (N_14399,N_8948,N_11510);
nand U14400 (N_14400,N_11035,N_11708);
and U14401 (N_14401,N_11921,N_7227);
nand U14402 (N_14402,N_8007,N_11881);
or U14403 (N_14403,N_6961,N_9439);
or U14404 (N_14404,N_6637,N_8164);
nor U14405 (N_14405,N_9761,N_7250);
nor U14406 (N_14406,N_11017,N_6857);
or U14407 (N_14407,N_11346,N_8389);
or U14408 (N_14408,N_10652,N_6539);
nor U14409 (N_14409,N_7418,N_6780);
nor U14410 (N_14410,N_6113,N_11211);
xor U14411 (N_14411,N_10452,N_11038);
xor U14412 (N_14412,N_7550,N_11347);
nor U14413 (N_14413,N_7809,N_7976);
xnor U14414 (N_14414,N_10410,N_10549);
nand U14415 (N_14415,N_11577,N_6658);
nor U14416 (N_14416,N_8674,N_10698);
nand U14417 (N_14417,N_8109,N_8950);
and U14418 (N_14418,N_7213,N_11757);
and U14419 (N_14419,N_8633,N_6448);
nor U14420 (N_14420,N_6145,N_11264);
xnor U14421 (N_14421,N_7914,N_7978);
and U14422 (N_14422,N_6374,N_7171);
and U14423 (N_14423,N_9105,N_9902);
nand U14424 (N_14424,N_10644,N_11745);
and U14425 (N_14425,N_11609,N_6502);
xor U14426 (N_14426,N_9473,N_7412);
xor U14427 (N_14427,N_11695,N_7437);
or U14428 (N_14428,N_7045,N_8754);
nand U14429 (N_14429,N_7827,N_7937);
xnor U14430 (N_14430,N_8738,N_9348);
nand U14431 (N_14431,N_7857,N_6871);
nand U14432 (N_14432,N_8299,N_6834);
nor U14433 (N_14433,N_9455,N_10939);
xor U14434 (N_14434,N_7395,N_7318);
xnor U14435 (N_14435,N_8123,N_8593);
or U14436 (N_14436,N_7996,N_11145);
and U14437 (N_14437,N_10364,N_9102);
or U14438 (N_14438,N_6049,N_10616);
or U14439 (N_14439,N_8837,N_11594);
nand U14440 (N_14440,N_10465,N_10435);
and U14441 (N_14441,N_10899,N_10634);
and U14442 (N_14442,N_10844,N_6201);
nor U14443 (N_14443,N_6329,N_9276);
nand U14444 (N_14444,N_8289,N_10558);
nand U14445 (N_14445,N_6578,N_10191);
xnor U14446 (N_14446,N_11258,N_8358);
nor U14447 (N_14447,N_9795,N_7509);
and U14448 (N_14448,N_7044,N_6394);
and U14449 (N_14449,N_9838,N_9504);
xor U14450 (N_14450,N_10572,N_8476);
nand U14451 (N_14451,N_7812,N_10804);
or U14452 (N_14452,N_6351,N_6873);
and U14453 (N_14453,N_6559,N_9287);
nor U14454 (N_14454,N_7806,N_9369);
or U14455 (N_14455,N_9547,N_7537);
or U14456 (N_14456,N_7099,N_6315);
xor U14457 (N_14457,N_11410,N_9647);
xnor U14458 (N_14458,N_10412,N_6801);
or U14459 (N_14459,N_8749,N_9283);
nand U14460 (N_14460,N_9625,N_11611);
nor U14461 (N_14461,N_11043,N_10224);
or U14462 (N_14462,N_7713,N_10786);
or U14463 (N_14463,N_9767,N_7421);
nor U14464 (N_14464,N_7856,N_10555);
nand U14465 (N_14465,N_7959,N_11498);
nand U14466 (N_14466,N_8874,N_11307);
xor U14467 (N_14467,N_9050,N_9532);
nand U14468 (N_14468,N_7541,N_6149);
xor U14469 (N_14469,N_6352,N_7212);
and U14470 (N_14470,N_7600,N_10001);
xnor U14471 (N_14471,N_7835,N_9871);
nor U14472 (N_14472,N_6288,N_6837);
and U14473 (N_14473,N_11665,N_9991);
and U14474 (N_14474,N_10908,N_9459);
and U14475 (N_14475,N_8848,N_6133);
nand U14476 (N_14476,N_10814,N_9876);
nor U14477 (N_14477,N_9955,N_9874);
nand U14478 (N_14478,N_8695,N_8964);
nor U14479 (N_14479,N_7178,N_11871);
and U14480 (N_14480,N_8646,N_6843);
nor U14481 (N_14481,N_7992,N_11931);
xor U14482 (N_14482,N_6032,N_9121);
and U14483 (N_14483,N_7320,N_9801);
and U14484 (N_14484,N_9100,N_7050);
xnor U14485 (N_14485,N_7944,N_9290);
nor U14486 (N_14486,N_8541,N_9452);
and U14487 (N_14487,N_9475,N_9103);
nor U14488 (N_14488,N_9979,N_11891);
or U14489 (N_14489,N_9248,N_10073);
or U14490 (N_14490,N_7420,N_6997);
and U14491 (N_14491,N_10267,N_6357);
xnor U14492 (N_14492,N_8689,N_9573);
nand U14493 (N_14493,N_7156,N_6392);
and U14494 (N_14494,N_11919,N_6128);
or U14495 (N_14495,N_7808,N_9890);
or U14496 (N_14496,N_6372,N_9160);
xnor U14497 (N_14497,N_10112,N_6264);
xor U14498 (N_14498,N_8846,N_11648);
and U14499 (N_14499,N_7730,N_9085);
xnor U14500 (N_14500,N_6139,N_9314);
nand U14501 (N_14501,N_9558,N_7170);
nand U14502 (N_14502,N_11499,N_6729);
nor U14503 (N_14503,N_9246,N_9503);
or U14504 (N_14504,N_7102,N_6262);
and U14505 (N_14505,N_11568,N_7624);
and U14506 (N_14506,N_8400,N_10499);
nand U14507 (N_14507,N_6159,N_11335);
nand U14508 (N_14508,N_10309,N_10607);
or U14509 (N_14509,N_8484,N_7858);
nand U14510 (N_14510,N_8500,N_7874);
nor U14511 (N_14511,N_7442,N_7399);
or U14512 (N_14512,N_8619,N_8688);
nor U14513 (N_14513,N_7636,N_7357);
nand U14514 (N_14514,N_6694,N_9405);
nand U14515 (N_14515,N_9449,N_9950);
or U14516 (N_14516,N_11072,N_8579);
and U14517 (N_14517,N_9058,N_7489);
nand U14518 (N_14518,N_7561,N_8341);
xnor U14519 (N_14519,N_9832,N_9110);
xnor U14520 (N_14520,N_7389,N_10856);
or U14521 (N_14521,N_6706,N_9044);
nor U14522 (N_14522,N_7379,N_10256);
or U14523 (N_14523,N_8411,N_6041);
xor U14524 (N_14524,N_7207,N_11185);
xor U14525 (N_14525,N_8563,N_10930);
nand U14526 (N_14526,N_8462,N_6456);
xor U14527 (N_14527,N_6928,N_8208);
nor U14528 (N_14528,N_8522,N_10878);
and U14529 (N_14529,N_9776,N_10005);
xnor U14530 (N_14530,N_6054,N_8554);
nand U14531 (N_14531,N_8562,N_6098);
or U14532 (N_14532,N_8599,N_8677);
xor U14533 (N_14533,N_9490,N_7939);
nand U14534 (N_14534,N_11773,N_10995);
and U14535 (N_14535,N_11803,N_6585);
and U14536 (N_14536,N_8743,N_8333);
nor U14537 (N_14537,N_7752,N_7909);
xnor U14538 (N_14538,N_6257,N_6659);
xor U14539 (N_14539,N_7392,N_10798);
nor U14540 (N_14540,N_9400,N_8291);
xnor U14541 (N_14541,N_10090,N_9827);
nand U14542 (N_14542,N_6777,N_9633);
or U14543 (N_14543,N_11104,N_11294);
nand U14544 (N_14544,N_10920,N_6497);
xor U14545 (N_14545,N_7055,N_8380);
nor U14546 (N_14546,N_7786,N_11426);
nor U14547 (N_14547,N_7031,N_9341);
and U14548 (N_14548,N_10717,N_8807);
nand U14549 (N_14549,N_8526,N_8875);
or U14550 (N_14550,N_8103,N_11805);
nor U14551 (N_14551,N_9236,N_10011);
nand U14552 (N_14552,N_6327,N_6612);
nor U14553 (N_14553,N_9480,N_11669);
or U14554 (N_14554,N_11050,N_10882);
nand U14555 (N_14555,N_10778,N_11793);
xor U14556 (N_14556,N_8653,N_6605);
and U14557 (N_14557,N_7341,N_8924);
nor U14558 (N_14558,N_11811,N_9768);
nand U14559 (N_14559,N_7957,N_7043);
nor U14560 (N_14560,N_11465,N_7253);
nand U14561 (N_14561,N_9995,N_6808);
nor U14562 (N_14562,N_6664,N_8625);
or U14563 (N_14563,N_9117,N_9126);
nand U14564 (N_14564,N_9563,N_6644);
and U14565 (N_14565,N_9052,N_7346);
nand U14566 (N_14566,N_9442,N_9263);
nor U14567 (N_14567,N_6110,N_8600);
nor U14568 (N_14568,N_7665,N_6268);
and U14569 (N_14569,N_6567,N_9877);
nor U14570 (N_14570,N_8880,N_10873);
xor U14571 (N_14571,N_9272,N_6141);
or U14572 (N_14572,N_6400,N_8078);
nand U14573 (N_14573,N_7367,N_11849);
or U14574 (N_14574,N_9997,N_10354);
or U14575 (N_14575,N_9594,N_6505);
and U14576 (N_14576,N_8503,N_10386);
or U14577 (N_14577,N_11967,N_9852);
nand U14578 (N_14578,N_11218,N_8248);
nor U14579 (N_14579,N_11974,N_10096);
nand U14580 (N_14580,N_6391,N_9580);
and U14581 (N_14581,N_8253,N_7797);
nand U14582 (N_14582,N_6192,N_9003);
or U14583 (N_14583,N_8822,N_9657);
nand U14584 (N_14584,N_8202,N_11514);
nor U14585 (N_14585,N_10087,N_7558);
nand U14586 (N_14586,N_9529,N_10569);
nand U14587 (N_14587,N_8487,N_6861);
xnor U14588 (N_14588,N_11371,N_6586);
nand U14589 (N_14589,N_8394,N_9954);
or U14590 (N_14590,N_9851,N_9500);
nor U14591 (N_14591,N_6082,N_8099);
xnor U14592 (N_14592,N_11356,N_7861);
and U14593 (N_14593,N_6312,N_6761);
xnor U14594 (N_14594,N_8649,N_8773);
and U14595 (N_14595,N_7154,N_7471);
or U14596 (N_14596,N_10641,N_8724);
xor U14597 (N_14597,N_8739,N_11304);
xor U14598 (N_14598,N_10668,N_11621);
nor U14599 (N_14599,N_7330,N_10482);
nand U14600 (N_14600,N_6127,N_6015);
nand U14601 (N_14601,N_8060,N_8548);
or U14602 (N_14602,N_11033,N_9199);
or U14603 (N_14603,N_6929,N_7702);
or U14604 (N_14604,N_8693,N_10003);
and U14605 (N_14605,N_8155,N_6037);
nand U14606 (N_14606,N_11790,N_7030);
or U14607 (N_14607,N_8968,N_9436);
nand U14608 (N_14608,N_7991,N_7605);
nor U14609 (N_14609,N_7360,N_7842);
or U14610 (N_14610,N_11725,N_7601);
nor U14611 (N_14611,N_7508,N_10334);
and U14612 (N_14612,N_11071,N_7277);
and U14613 (N_14613,N_11192,N_8490);
or U14614 (N_14614,N_10874,N_11883);
nand U14615 (N_14615,N_9734,N_6019);
or U14616 (N_14616,N_7918,N_11168);
nand U14617 (N_14617,N_9909,N_6265);
nand U14618 (N_14618,N_11798,N_10547);
nand U14619 (N_14619,N_8651,N_9365);
xor U14620 (N_14620,N_7077,N_9161);
or U14621 (N_14621,N_6243,N_8185);
or U14622 (N_14622,N_8465,N_6485);
nand U14623 (N_14623,N_6246,N_8397);
or U14624 (N_14624,N_11138,N_11542);
xnor U14625 (N_14625,N_8776,N_8561);
xor U14626 (N_14626,N_11084,N_11958);
and U14627 (N_14627,N_9621,N_7824);
and U14628 (N_14628,N_10595,N_10299);
or U14629 (N_14629,N_9520,N_6850);
nand U14630 (N_14630,N_9329,N_7788);
nor U14631 (N_14631,N_8433,N_6574);
xnor U14632 (N_14632,N_11473,N_9620);
nor U14633 (N_14633,N_9335,N_7798);
nand U14634 (N_14634,N_6735,N_10438);
or U14635 (N_14635,N_9240,N_7181);
nand U14636 (N_14636,N_10285,N_7295);
nand U14637 (N_14637,N_9361,N_6203);
or U14638 (N_14638,N_7417,N_6628);
or U14639 (N_14639,N_6955,N_8669);
nor U14640 (N_14640,N_7662,N_8137);
or U14641 (N_14641,N_11115,N_6455);
nand U14642 (N_14642,N_9201,N_9729);
nand U14643 (N_14643,N_7863,N_11186);
xnor U14644 (N_14644,N_9987,N_8700);
nand U14645 (N_14645,N_9574,N_8264);
and U14646 (N_14646,N_10122,N_8395);
xor U14647 (N_14647,N_6237,N_8577);
nand U14648 (N_14648,N_9826,N_9999);
nand U14649 (N_14649,N_9700,N_11727);
xnor U14650 (N_14650,N_10458,N_6945);
and U14651 (N_14651,N_6771,N_7339);
xnor U14652 (N_14652,N_7069,N_8821);
nor U14653 (N_14653,N_11721,N_8205);
nand U14654 (N_14654,N_11710,N_10790);
and U14655 (N_14655,N_7694,N_9814);
xnor U14656 (N_14656,N_8909,N_10273);
and U14657 (N_14657,N_9389,N_8662);
or U14658 (N_14658,N_6172,N_8861);
or U14659 (N_14659,N_7141,N_11889);
nand U14660 (N_14660,N_7887,N_11040);
nand U14661 (N_14661,N_11893,N_9539);
nand U14662 (N_14662,N_11991,N_11277);
xor U14663 (N_14663,N_10075,N_6940);
and U14664 (N_14664,N_8608,N_6707);
nor U14665 (N_14665,N_6121,N_10886);
or U14666 (N_14666,N_10818,N_7924);
xor U14667 (N_14667,N_8034,N_7877);
or U14668 (N_14668,N_11059,N_7688);
xnor U14669 (N_14669,N_7409,N_7166);
xor U14670 (N_14670,N_9499,N_10646);
and U14671 (N_14671,N_6385,N_11452);
and U14672 (N_14672,N_8678,N_10377);
or U14673 (N_14673,N_10751,N_6618);
nor U14674 (N_14674,N_10608,N_8698);
xor U14675 (N_14675,N_7676,N_8198);
xor U14676 (N_14676,N_11877,N_10304);
xnor U14677 (N_14677,N_7305,N_11074);
xnor U14678 (N_14678,N_10893,N_9192);
nand U14679 (N_14679,N_8943,N_8980);
nand U14680 (N_14680,N_11687,N_7463);
xnor U14681 (N_14681,N_9185,N_8789);
nor U14682 (N_14682,N_8305,N_9016);
or U14683 (N_14683,N_10992,N_9824);
or U14684 (N_14684,N_10066,N_10265);
xnor U14685 (N_14685,N_11825,N_11571);
nor U14686 (N_14686,N_9065,N_11556);
nor U14687 (N_14687,N_8416,N_11932);
and U14688 (N_14688,N_9437,N_10938);
nor U14689 (N_14689,N_11614,N_11961);
and U14690 (N_14690,N_9905,N_8779);
xor U14691 (N_14691,N_9867,N_9414);
nand U14692 (N_14692,N_9190,N_11684);
or U14693 (N_14693,N_6427,N_6554);
nor U14694 (N_14694,N_11800,N_7300);
xor U14695 (N_14695,N_10710,N_7505);
or U14696 (N_14696,N_6884,N_9873);
nand U14697 (N_14697,N_9708,N_11068);
nor U14698 (N_14698,N_11874,N_10152);
and U14699 (N_14699,N_9609,N_7599);
nor U14700 (N_14700,N_11226,N_8329);
nor U14701 (N_14701,N_11389,N_8468);
or U14702 (N_14702,N_10319,N_10861);
or U14703 (N_14703,N_7394,N_7548);
nor U14704 (N_14704,N_6147,N_8632);
xnor U14705 (N_14705,N_7296,N_6697);
or U14706 (N_14706,N_11876,N_11873);
nor U14707 (N_14707,N_9721,N_8601);
and U14708 (N_14708,N_9577,N_11616);
and U14709 (N_14709,N_7454,N_10076);
nand U14710 (N_14710,N_9077,N_10542);
nand U14711 (N_14711,N_11903,N_7546);
or U14712 (N_14712,N_9007,N_6311);
and U14713 (N_14713,N_10042,N_8452);
nand U14714 (N_14714,N_10730,N_11575);
and U14715 (N_14715,N_8627,N_9040);
or U14716 (N_14716,N_6858,N_11481);
and U14717 (N_14717,N_8778,N_10332);
nand U14718 (N_14718,N_7434,N_10842);
nor U14719 (N_14719,N_6716,N_6130);
nor U14720 (N_14720,N_6903,N_7414);
xnor U14721 (N_14721,N_10600,N_10284);
nor U14722 (N_14722,N_9942,N_7549);
nor U14723 (N_14723,N_7753,N_8945);
or U14724 (N_14724,N_10483,N_7712);
and U14725 (N_14725,N_7232,N_8033);
or U14726 (N_14726,N_6024,N_7501);
nor U14727 (N_14727,N_6150,N_11142);
nand U14728 (N_14728,N_8860,N_6662);
xnor U14729 (N_14729,N_11025,N_6804);
and U14730 (N_14730,N_10540,N_9592);
nand U14731 (N_14731,N_6364,N_7464);
nand U14732 (N_14732,N_6699,N_8336);
and U14733 (N_14733,N_10837,N_10245);
xnor U14734 (N_14734,N_6988,N_7927);
xor U14735 (N_14735,N_8967,N_11791);
nor U14736 (N_14736,N_9502,N_6330);
and U14737 (N_14737,N_8665,N_11951);
xnor U14738 (N_14738,N_10201,N_7243);
nor U14739 (N_14739,N_8900,N_8556);
or U14740 (N_14740,N_8286,N_9811);
nand U14741 (N_14741,N_11419,N_10252);
or U14742 (N_14742,N_10803,N_6182);
or U14743 (N_14743,N_11048,N_8714);
xor U14744 (N_14744,N_8093,N_6059);
and U14745 (N_14745,N_7748,N_6604);
nor U14746 (N_14746,N_7242,N_7666);
nor U14747 (N_14747,N_6747,N_10165);
or U14748 (N_14748,N_7235,N_8486);
or U14749 (N_14749,N_8795,N_8296);
nand U14750 (N_14750,N_11297,N_6880);
or U14751 (N_14751,N_6013,N_7738);
and U14752 (N_14752,N_10174,N_8723);
or U14753 (N_14753,N_6611,N_9425);
and U14754 (N_14754,N_8211,N_11161);
or U14755 (N_14755,N_10576,N_10812);
and U14756 (N_14756,N_11411,N_7090);
and U14757 (N_14757,N_6657,N_9541);
xnor U14758 (N_14758,N_6274,N_6572);
nand U14759 (N_14759,N_11597,N_6221);
and U14760 (N_14760,N_6513,N_8815);
xor U14761 (N_14761,N_10579,N_6890);
nor U14762 (N_14762,N_8415,N_6533);
or U14763 (N_14763,N_8457,N_6679);
or U14764 (N_14764,N_8018,N_11223);
xor U14765 (N_14765,N_9723,N_9429);
and U14766 (N_14766,N_6711,N_9367);
and U14767 (N_14767,N_7946,N_8804);
nor U14768 (N_14768,N_11219,N_7544);
or U14769 (N_14769,N_7911,N_9122);
or U14770 (N_14770,N_11326,N_11647);
nor U14771 (N_14771,N_6898,N_10115);
and U14772 (N_14772,N_7906,N_7267);
and U14773 (N_14773,N_9758,N_8946);
xor U14774 (N_14774,N_11198,N_7478);
nand U14775 (N_14775,N_11262,N_9208);
nor U14776 (N_14776,N_6057,N_11588);
and U14777 (N_14777,N_6491,N_9956);
xnor U14778 (N_14778,N_11544,N_10959);
xnor U14779 (N_14779,N_10957,N_8581);
nor U14780 (N_14780,N_10035,N_6949);
nand U14781 (N_14781,N_11732,N_6661);
and U14782 (N_14782,N_11409,N_8982);
and U14783 (N_14783,N_6208,N_6900);
nand U14784 (N_14784,N_9850,N_11299);
nand U14785 (N_14785,N_7923,N_7190);
nor U14786 (N_14786,N_9391,N_11380);
nor U14787 (N_14787,N_9864,N_11844);
xor U14788 (N_14788,N_6214,N_11099);
xor U14789 (N_14789,N_9260,N_10665);
nor U14790 (N_14790,N_6797,N_7462);
nor U14791 (N_14791,N_9212,N_6005);
and U14792 (N_14792,N_7138,N_10748);
nor U14793 (N_14793,N_10948,N_8453);
xnor U14794 (N_14794,N_8383,N_7551);
or U14795 (N_14795,N_7639,N_10617);
nor U14796 (N_14796,N_9654,N_11022);
nand U14797 (N_14797,N_8648,N_11752);
nand U14798 (N_14798,N_7285,N_8762);
and U14799 (N_14799,N_11200,N_6120);
xnor U14800 (N_14800,N_7189,N_6983);
xnor U14801 (N_14801,N_10609,N_6866);
or U14802 (N_14802,N_8224,N_8907);
xnor U14803 (N_14803,N_7854,N_9765);
nand U14804 (N_14804,N_8184,N_11724);
xnor U14805 (N_14805,N_8009,N_9387);
and U14806 (N_14806,N_10740,N_9638);
or U14807 (N_14807,N_11204,N_8624);
nand U14808 (N_14808,N_10672,N_9527);
nand U14809 (N_14809,N_6046,N_8229);
and U14810 (N_14810,N_8471,N_9483);
nor U14811 (N_14811,N_11776,N_6353);
or U14812 (N_14812,N_8991,N_6285);
nand U14813 (N_14813,N_7622,N_7263);
nand U14814 (N_14814,N_11224,N_11365);
nor U14815 (N_14815,N_6435,N_8545);
nand U14816 (N_14816,N_10323,N_7775);
xnor U14817 (N_14817,N_9273,N_6816);
and U14818 (N_14818,N_7240,N_8375);
xnor U14819 (N_14819,N_7849,N_6684);
xnor U14820 (N_14820,N_11349,N_9724);
nor U14821 (N_14821,N_8766,N_9769);
and U14822 (N_14822,N_8080,N_9038);
nor U14823 (N_14823,N_11096,N_6293);
nand U14824 (N_14824,N_7479,N_8130);
xnor U14825 (N_14825,N_9268,N_9492);
or U14826 (N_14826,N_11463,N_9325);
nor U14827 (N_14827,N_6625,N_6481);
nand U14828 (N_14828,N_9451,N_6118);
nor U14829 (N_14829,N_10674,N_8881);
and U14830 (N_14830,N_7498,N_9605);
or U14831 (N_14831,N_7344,N_8245);
nand U14832 (N_14832,N_11012,N_7097);
and U14833 (N_14833,N_11858,N_6174);
and U14834 (N_14834,N_7679,N_11772);
nand U14835 (N_14835,N_10791,N_8320);
xnor U14836 (N_14836,N_10175,N_10329);
nand U14837 (N_14837,N_11362,N_8974);
xnor U14838 (N_14838,N_11945,N_9744);
xnor U14839 (N_14839,N_10974,N_8812);
and U14840 (N_14840,N_9796,N_9495);
xor U14841 (N_14841,N_10945,N_10411);
nand U14842 (N_14842,N_10799,N_10556);
or U14843 (N_14843,N_6996,N_11225);
nor U14844 (N_14844,N_11712,N_8569);
nor U14845 (N_14845,N_9645,N_7742);
and U14846 (N_14846,N_6248,N_6325);
xor U14847 (N_14847,N_6496,N_8322);
xnor U14848 (N_14848,N_9261,N_8547);
xnor U14849 (N_14849,N_8081,N_7184);
nand U14850 (N_14850,N_6242,N_8102);
nor U14851 (N_14851,N_11666,N_10328);
and U14852 (N_14852,N_11323,N_9632);
and U14853 (N_14853,N_9507,N_10573);
nor U14854 (N_14854,N_8192,N_10453);
xnor U14855 (N_14855,N_7397,N_8221);
nor U14856 (N_14856,N_11950,N_11002);
nor U14857 (N_14857,N_10960,N_10128);
nor U14858 (N_14858,N_11635,N_10839);
nor U14859 (N_14859,N_8805,N_8814);
or U14860 (N_14860,N_9629,N_10570);
nor U14861 (N_14861,N_11372,N_7419);
nor U14862 (N_14862,N_9670,N_9774);
nand U14863 (N_14863,N_8828,N_9446);
nand U14864 (N_14864,N_9471,N_6692);
or U14865 (N_14865,N_8027,N_8498);
nor U14866 (N_14866,N_11112,N_11484);
and U14867 (N_14867,N_11828,N_8090);
nand U14868 (N_14868,N_10058,N_6219);
xnor U14869 (N_14869,N_6982,N_7352);
or U14870 (N_14870,N_11305,N_7839);
or U14871 (N_14871,N_9409,N_11417);
xor U14872 (N_14872,N_6109,N_10681);
nand U14873 (N_14873,N_10271,N_6538);
or U14874 (N_14874,N_6209,N_8505);
xnor U14875 (N_14875,N_11170,N_8282);
nor U14876 (N_14876,N_8764,N_8934);
nor U14877 (N_14877,N_8853,N_7556);
and U14878 (N_14878,N_6920,N_6769);
xnor U14879 (N_14879,N_7467,N_9454);
and U14880 (N_14880,N_10530,N_10921);
xor U14881 (N_14881,N_6389,N_9143);
or U14882 (N_14882,N_8136,N_8763);
xnor U14883 (N_14883,N_8493,N_10752);
or U14884 (N_14884,N_6278,N_7796);
xor U14885 (N_14885,N_6443,N_9718);
xor U14886 (N_14886,N_8733,N_11337);
nand U14887 (N_14887,N_6674,N_9610);
or U14888 (N_14888,N_7038,N_7513);
nand U14889 (N_14889,N_7047,N_6266);
or U14890 (N_14890,N_11351,N_6198);
nand U14891 (N_14891,N_10541,N_10789);
or U14892 (N_14892,N_11242,N_8138);
and U14893 (N_14893,N_10199,N_11914);
nor U14894 (N_14894,N_9840,N_7935);
nor U14895 (N_14895,N_6478,N_7890);
nand U14896 (N_14896,N_9912,N_7364);
xnor U14897 (N_14897,N_7613,N_10022);
xor U14898 (N_14898,N_9972,N_8707);
or U14899 (N_14899,N_8867,N_8786);
nor U14900 (N_14900,N_9139,N_8071);
and U14901 (N_14901,N_11110,N_8379);
nand U14902 (N_14902,N_9887,N_11344);
or U14903 (N_14903,N_10770,N_9735);
nor U14904 (N_14904,N_11619,N_8854);
or U14905 (N_14905,N_7938,N_8585);
or U14906 (N_14906,N_8121,N_11533);
xnor U14907 (N_14907,N_6340,N_6337);
or U14908 (N_14908,N_8978,N_7358);
nor U14909 (N_14909,N_7607,N_11159);
nor U14910 (N_14910,N_8181,N_7980);
or U14911 (N_14911,N_9069,N_9373);
xnor U14912 (N_14912,N_11569,N_11190);
and U14913 (N_14913,N_11150,N_7526);
nor U14914 (N_14914,N_11519,N_10150);
nor U14915 (N_14915,N_10506,N_11105);
and U14916 (N_14916,N_11522,N_9444);
and U14917 (N_14917,N_9434,N_11645);
nor U14918 (N_14918,N_6286,N_7041);
or U14919 (N_14919,N_11205,N_11248);
or U14920 (N_14920,N_6952,N_10426);
or U14921 (N_14921,N_7218,N_8882);
nand U14922 (N_14922,N_7847,N_9685);
nand U14923 (N_14923,N_6464,N_11589);
nor U14924 (N_14924,N_9775,N_9375);
nor U14925 (N_14925,N_8098,N_10696);
nor U14926 (N_14926,N_11972,N_6270);
nor U14927 (N_14927,N_11073,N_11717);
or U14928 (N_14928,N_10902,N_8756);
and U14929 (N_14929,N_7062,N_6913);
xor U14930 (N_14930,N_8567,N_10053);
nor U14931 (N_14931,N_11596,N_10114);
nand U14932 (N_14932,N_8030,N_6068);
xnor U14933 (N_14933,N_10289,N_9614);
nand U14934 (N_14934,N_9959,N_6937);
nor U14935 (N_14935,N_7631,N_9977);
and U14936 (N_14936,N_8905,N_8518);
and U14937 (N_14937,N_9530,N_6276);
nand U14938 (N_14938,N_9041,N_8813);
nor U14939 (N_14939,N_10852,N_7833);
nand U14940 (N_14940,N_9156,N_9742);
xor U14941 (N_14941,N_9889,N_9749);
xor U14942 (N_14942,N_7700,N_11697);
nor U14943 (N_14943,N_11583,N_8424);
and U14944 (N_14944,N_10857,N_7727);
or U14945 (N_14945,N_9269,N_7035);
or U14946 (N_14946,N_8801,N_6750);
and U14947 (N_14947,N_11848,N_6721);
and U14948 (N_14948,N_10692,N_7398);
nor U14949 (N_14949,N_9757,N_8000);
xor U14950 (N_14950,N_8008,N_6404);
xor U14951 (N_14951,N_6084,N_9891);
nand U14952 (N_14952,N_9134,N_11608);
nor U14953 (N_14953,N_11332,N_8566);
and U14954 (N_14954,N_6907,N_7214);
nor U14955 (N_14955,N_11133,N_6324);
and U14956 (N_14956,N_6859,N_7303);
xnor U14957 (N_14957,N_7408,N_11737);
nand U14958 (N_14958,N_7687,N_9282);
xor U14959 (N_14959,N_9057,N_6500);
nand U14960 (N_14960,N_10989,N_9674);
xnor U14961 (N_14961,N_9416,N_8347);
and U14962 (N_14962,N_10519,N_7577);
nand U14963 (N_14963,N_11061,N_10014);
and U14964 (N_14964,N_10000,N_7628);
nand U14965 (N_14965,N_10489,N_7751);
or U14966 (N_14966,N_8002,N_6104);
xnor U14967 (N_14967,N_8628,N_10841);
nand U14968 (N_14968,N_11911,N_9119);
nor U14969 (N_14969,N_11331,N_6727);
xnor U14970 (N_14970,N_8728,N_9417);
nor U14971 (N_14971,N_9064,N_9021);
nand U14972 (N_14972,N_7554,N_7588);
nor U14973 (N_14973,N_8129,N_8149);
and U14974 (N_14974,N_11901,N_9144);
nand U14975 (N_14975,N_10524,N_10387);
and U14976 (N_14976,N_6668,N_8972);
or U14977 (N_14977,N_9170,N_8220);
and U14978 (N_14978,N_10306,N_10361);
nor U14979 (N_14979,N_11812,N_10716);
or U14980 (N_14980,N_7585,N_9971);
xor U14981 (N_14981,N_10724,N_9967);
and U14982 (N_14982,N_11101,N_11711);
and U14983 (N_14983,N_8266,N_8458);
or U14984 (N_14984,N_11960,N_6194);
nor U14985 (N_14985,N_10322,N_10877);
nor U14986 (N_14986,N_10733,N_8836);
nor U14987 (N_14987,N_7715,N_7025);
nor U14988 (N_14988,N_8965,N_11296);
nand U14989 (N_14989,N_7290,N_7649);
and U14990 (N_14990,N_9704,N_11249);
nor U14991 (N_14991,N_10496,N_9243);
nand U14992 (N_14992,N_11303,N_6823);
and U14993 (N_14993,N_6779,N_6971);
nor U14994 (N_14994,N_7598,N_6016);
or U14995 (N_14995,N_10624,N_11782);
nor U14996 (N_14996,N_7233,N_8031);
nor U14997 (N_14997,N_11536,N_9617);
and U14998 (N_14998,N_11624,N_6335);
xnor U14999 (N_14999,N_8455,N_8933);
or U15000 (N_15000,N_9971,N_7271);
or U15001 (N_15001,N_11071,N_10262);
nor U15002 (N_15002,N_10113,N_8762);
nand U15003 (N_15003,N_10213,N_8923);
nand U15004 (N_15004,N_9134,N_7201);
and U15005 (N_15005,N_6352,N_6412);
nor U15006 (N_15006,N_10092,N_6931);
or U15007 (N_15007,N_9775,N_11167);
nor U15008 (N_15008,N_9381,N_8837);
nor U15009 (N_15009,N_7869,N_8682);
nand U15010 (N_15010,N_10184,N_10645);
xnor U15011 (N_15011,N_10614,N_9372);
nor U15012 (N_15012,N_8159,N_7950);
nor U15013 (N_15013,N_9837,N_8163);
or U15014 (N_15014,N_9228,N_7484);
nor U15015 (N_15015,N_9354,N_9918);
or U15016 (N_15016,N_8646,N_7949);
and U15017 (N_15017,N_9507,N_6120);
nand U15018 (N_15018,N_10518,N_6066);
nor U15019 (N_15019,N_6876,N_10567);
and U15020 (N_15020,N_8863,N_9896);
nand U15021 (N_15021,N_11395,N_11589);
xnor U15022 (N_15022,N_8277,N_9069);
nor U15023 (N_15023,N_10564,N_6408);
and U15024 (N_15024,N_9240,N_9816);
xnor U15025 (N_15025,N_6241,N_6199);
xnor U15026 (N_15026,N_9517,N_11021);
nor U15027 (N_15027,N_9742,N_10490);
nor U15028 (N_15028,N_11820,N_8439);
xor U15029 (N_15029,N_8292,N_9603);
xnor U15030 (N_15030,N_8876,N_9054);
or U15031 (N_15031,N_10171,N_6392);
nand U15032 (N_15032,N_11354,N_10780);
or U15033 (N_15033,N_11550,N_7104);
xor U15034 (N_15034,N_6206,N_8664);
xnor U15035 (N_15035,N_11667,N_11854);
or U15036 (N_15036,N_6114,N_7423);
nand U15037 (N_15037,N_10411,N_10610);
and U15038 (N_15038,N_7415,N_10206);
nand U15039 (N_15039,N_6070,N_6807);
xor U15040 (N_15040,N_8687,N_10352);
and U15041 (N_15041,N_8857,N_11194);
and U15042 (N_15042,N_11635,N_9844);
or U15043 (N_15043,N_10719,N_9170);
and U15044 (N_15044,N_7078,N_6581);
and U15045 (N_15045,N_10935,N_10287);
or U15046 (N_15046,N_8270,N_9998);
and U15047 (N_15047,N_7138,N_8498);
nor U15048 (N_15048,N_7588,N_11833);
or U15049 (N_15049,N_10434,N_11759);
or U15050 (N_15050,N_8670,N_8578);
nor U15051 (N_15051,N_6291,N_6450);
nand U15052 (N_15052,N_8284,N_7647);
and U15053 (N_15053,N_10167,N_11268);
nand U15054 (N_15054,N_7657,N_7849);
nand U15055 (N_15055,N_10950,N_11734);
nand U15056 (N_15056,N_8345,N_11812);
xnor U15057 (N_15057,N_7708,N_6666);
nand U15058 (N_15058,N_8713,N_11256);
xor U15059 (N_15059,N_7937,N_8403);
nor U15060 (N_15060,N_11689,N_7169);
or U15061 (N_15061,N_6100,N_8359);
nand U15062 (N_15062,N_6788,N_8331);
nand U15063 (N_15063,N_8707,N_6668);
nor U15064 (N_15064,N_7171,N_8630);
xnor U15065 (N_15065,N_9122,N_7306);
xor U15066 (N_15066,N_8645,N_8431);
xor U15067 (N_15067,N_10543,N_8953);
nor U15068 (N_15068,N_9508,N_8184);
nand U15069 (N_15069,N_10927,N_6807);
nor U15070 (N_15070,N_9824,N_7084);
xor U15071 (N_15071,N_6559,N_11000);
xor U15072 (N_15072,N_7650,N_10932);
or U15073 (N_15073,N_8715,N_9051);
and U15074 (N_15074,N_9207,N_11781);
or U15075 (N_15075,N_6291,N_8901);
or U15076 (N_15076,N_9985,N_7679);
xor U15077 (N_15077,N_10664,N_7518);
and U15078 (N_15078,N_9621,N_9195);
nor U15079 (N_15079,N_8873,N_8364);
nand U15080 (N_15080,N_9862,N_9301);
and U15081 (N_15081,N_8922,N_8841);
or U15082 (N_15082,N_8179,N_6941);
nor U15083 (N_15083,N_9767,N_10896);
xnor U15084 (N_15084,N_8781,N_6709);
or U15085 (N_15085,N_6237,N_9654);
nand U15086 (N_15086,N_11437,N_10845);
nand U15087 (N_15087,N_6144,N_6946);
xor U15088 (N_15088,N_11392,N_8214);
and U15089 (N_15089,N_6288,N_6488);
and U15090 (N_15090,N_9224,N_9131);
or U15091 (N_15091,N_10335,N_8741);
xnor U15092 (N_15092,N_10031,N_10766);
or U15093 (N_15093,N_9155,N_10590);
nor U15094 (N_15094,N_11786,N_6657);
nor U15095 (N_15095,N_7929,N_7518);
and U15096 (N_15096,N_9020,N_11542);
xnor U15097 (N_15097,N_9724,N_7653);
and U15098 (N_15098,N_7241,N_8254);
xor U15099 (N_15099,N_6314,N_9972);
and U15100 (N_15100,N_6414,N_7230);
nand U15101 (N_15101,N_8289,N_10369);
or U15102 (N_15102,N_6815,N_8293);
nand U15103 (N_15103,N_8914,N_10678);
and U15104 (N_15104,N_6689,N_11125);
xor U15105 (N_15105,N_11736,N_9626);
nand U15106 (N_15106,N_7809,N_7643);
nor U15107 (N_15107,N_6111,N_6108);
nand U15108 (N_15108,N_8096,N_9586);
and U15109 (N_15109,N_6521,N_7224);
nor U15110 (N_15110,N_9747,N_6747);
and U15111 (N_15111,N_7109,N_9295);
and U15112 (N_15112,N_6509,N_8423);
or U15113 (N_15113,N_11671,N_8333);
nor U15114 (N_15114,N_11297,N_11124);
nand U15115 (N_15115,N_7439,N_6603);
or U15116 (N_15116,N_9743,N_11161);
or U15117 (N_15117,N_9979,N_9657);
or U15118 (N_15118,N_7911,N_9676);
xnor U15119 (N_15119,N_11491,N_9003);
nand U15120 (N_15120,N_7973,N_7490);
and U15121 (N_15121,N_6688,N_6941);
or U15122 (N_15122,N_8374,N_9023);
xnor U15123 (N_15123,N_6321,N_8513);
and U15124 (N_15124,N_11792,N_10121);
nor U15125 (N_15125,N_10388,N_11885);
or U15126 (N_15126,N_6703,N_7360);
or U15127 (N_15127,N_8573,N_6183);
or U15128 (N_15128,N_8861,N_9691);
xnor U15129 (N_15129,N_8449,N_9907);
nand U15130 (N_15130,N_10529,N_9068);
and U15131 (N_15131,N_8723,N_6589);
nand U15132 (N_15132,N_10796,N_7556);
xor U15133 (N_15133,N_10910,N_8435);
and U15134 (N_15134,N_6559,N_8325);
or U15135 (N_15135,N_9417,N_6752);
nand U15136 (N_15136,N_11038,N_10088);
nor U15137 (N_15137,N_7726,N_6507);
nand U15138 (N_15138,N_8322,N_10654);
nand U15139 (N_15139,N_7227,N_6914);
nor U15140 (N_15140,N_6135,N_6940);
nand U15141 (N_15141,N_8377,N_9452);
or U15142 (N_15142,N_7320,N_10227);
xor U15143 (N_15143,N_9228,N_10160);
nor U15144 (N_15144,N_9931,N_11629);
and U15145 (N_15145,N_6571,N_9665);
or U15146 (N_15146,N_7799,N_6715);
nor U15147 (N_15147,N_6755,N_7002);
nor U15148 (N_15148,N_11861,N_9469);
and U15149 (N_15149,N_6332,N_7972);
nor U15150 (N_15150,N_9263,N_10776);
nand U15151 (N_15151,N_9466,N_7377);
nand U15152 (N_15152,N_9940,N_11760);
nor U15153 (N_15153,N_11566,N_7607);
nand U15154 (N_15154,N_7053,N_10929);
nand U15155 (N_15155,N_9566,N_7245);
nand U15156 (N_15156,N_7760,N_9369);
nor U15157 (N_15157,N_7549,N_7428);
xnor U15158 (N_15158,N_7057,N_9957);
or U15159 (N_15159,N_7150,N_9613);
and U15160 (N_15160,N_10571,N_9262);
xor U15161 (N_15161,N_7319,N_7529);
xnor U15162 (N_15162,N_7341,N_7918);
and U15163 (N_15163,N_10367,N_11844);
xor U15164 (N_15164,N_8204,N_11975);
or U15165 (N_15165,N_10253,N_7046);
xor U15166 (N_15166,N_9196,N_9274);
nor U15167 (N_15167,N_9601,N_11445);
or U15168 (N_15168,N_8640,N_7267);
xor U15169 (N_15169,N_8732,N_11411);
nand U15170 (N_15170,N_7177,N_11117);
nor U15171 (N_15171,N_9948,N_10822);
or U15172 (N_15172,N_9676,N_10516);
nand U15173 (N_15173,N_9701,N_10369);
nand U15174 (N_15174,N_11489,N_11895);
nand U15175 (N_15175,N_10840,N_11597);
nand U15176 (N_15176,N_6647,N_6344);
nand U15177 (N_15177,N_8760,N_6722);
and U15178 (N_15178,N_6840,N_10178);
nand U15179 (N_15179,N_8736,N_7258);
and U15180 (N_15180,N_8081,N_6550);
and U15181 (N_15181,N_8176,N_10848);
nor U15182 (N_15182,N_10720,N_8161);
and U15183 (N_15183,N_9905,N_6529);
xor U15184 (N_15184,N_6076,N_10665);
or U15185 (N_15185,N_8914,N_7573);
and U15186 (N_15186,N_8835,N_11338);
xor U15187 (N_15187,N_6794,N_7865);
nand U15188 (N_15188,N_9002,N_8256);
and U15189 (N_15189,N_7407,N_11631);
and U15190 (N_15190,N_6078,N_10007);
nor U15191 (N_15191,N_7686,N_11278);
nor U15192 (N_15192,N_11152,N_6246);
and U15193 (N_15193,N_11659,N_9184);
xor U15194 (N_15194,N_6942,N_8934);
nor U15195 (N_15195,N_6156,N_10923);
nand U15196 (N_15196,N_6776,N_6462);
nand U15197 (N_15197,N_8636,N_9092);
or U15198 (N_15198,N_11761,N_9509);
or U15199 (N_15199,N_10268,N_7035);
and U15200 (N_15200,N_6112,N_9714);
nor U15201 (N_15201,N_6053,N_11963);
nand U15202 (N_15202,N_10473,N_11838);
xnor U15203 (N_15203,N_8916,N_8004);
and U15204 (N_15204,N_8085,N_6650);
nand U15205 (N_15205,N_8208,N_8326);
xor U15206 (N_15206,N_6024,N_7681);
or U15207 (N_15207,N_7689,N_8676);
or U15208 (N_15208,N_9432,N_8191);
nor U15209 (N_15209,N_8097,N_6408);
and U15210 (N_15210,N_9344,N_9561);
nand U15211 (N_15211,N_8462,N_6099);
nor U15212 (N_15212,N_7513,N_9448);
or U15213 (N_15213,N_10869,N_11474);
xnor U15214 (N_15214,N_11869,N_6740);
and U15215 (N_15215,N_7661,N_6047);
nand U15216 (N_15216,N_10621,N_7660);
and U15217 (N_15217,N_8651,N_11531);
nor U15218 (N_15218,N_7149,N_6238);
xor U15219 (N_15219,N_8211,N_9725);
and U15220 (N_15220,N_10780,N_6030);
nor U15221 (N_15221,N_7990,N_11836);
and U15222 (N_15222,N_8515,N_10827);
and U15223 (N_15223,N_10744,N_7515);
xnor U15224 (N_15224,N_9842,N_7303);
xnor U15225 (N_15225,N_7116,N_7060);
nor U15226 (N_15226,N_9208,N_7439);
nand U15227 (N_15227,N_9727,N_6347);
xnor U15228 (N_15228,N_6282,N_6576);
and U15229 (N_15229,N_6952,N_11172);
nand U15230 (N_15230,N_8472,N_8017);
nor U15231 (N_15231,N_8791,N_9334);
nand U15232 (N_15232,N_11742,N_6383);
and U15233 (N_15233,N_8078,N_11529);
and U15234 (N_15234,N_9465,N_8611);
nand U15235 (N_15235,N_8818,N_8873);
xor U15236 (N_15236,N_6188,N_6242);
nand U15237 (N_15237,N_9134,N_7395);
xor U15238 (N_15238,N_11061,N_9811);
nand U15239 (N_15239,N_9612,N_6680);
or U15240 (N_15240,N_7826,N_6291);
or U15241 (N_15241,N_6199,N_6776);
xor U15242 (N_15242,N_8137,N_9505);
xnor U15243 (N_15243,N_11477,N_11913);
nor U15244 (N_15244,N_11029,N_8977);
nand U15245 (N_15245,N_6671,N_7672);
nand U15246 (N_15246,N_7512,N_10689);
or U15247 (N_15247,N_10203,N_7918);
or U15248 (N_15248,N_9609,N_11606);
nor U15249 (N_15249,N_9884,N_11859);
and U15250 (N_15250,N_6926,N_11750);
and U15251 (N_15251,N_8749,N_7328);
or U15252 (N_15252,N_6744,N_7482);
xor U15253 (N_15253,N_10066,N_9423);
or U15254 (N_15254,N_7450,N_11500);
or U15255 (N_15255,N_6618,N_7912);
nand U15256 (N_15256,N_10068,N_6607);
or U15257 (N_15257,N_11324,N_9313);
nor U15258 (N_15258,N_6739,N_6949);
or U15259 (N_15259,N_8710,N_11148);
nor U15260 (N_15260,N_6358,N_10006);
or U15261 (N_15261,N_7536,N_11185);
nand U15262 (N_15262,N_9599,N_6374);
nor U15263 (N_15263,N_11180,N_8515);
nor U15264 (N_15264,N_9350,N_11538);
nand U15265 (N_15265,N_7705,N_9236);
or U15266 (N_15266,N_11093,N_7519);
nand U15267 (N_15267,N_7859,N_9520);
xor U15268 (N_15268,N_8620,N_11859);
xor U15269 (N_15269,N_6166,N_8253);
and U15270 (N_15270,N_9639,N_6340);
xnor U15271 (N_15271,N_8910,N_9362);
or U15272 (N_15272,N_9908,N_7972);
xnor U15273 (N_15273,N_9482,N_7864);
nor U15274 (N_15274,N_7565,N_6822);
or U15275 (N_15275,N_8301,N_10658);
nand U15276 (N_15276,N_10364,N_9457);
or U15277 (N_15277,N_8745,N_10902);
nand U15278 (N_15278,N_8402,N_6717);
and U15279 (N_15279,N_7736,N_8050);
xnor U15280 (N_15280,N_9040,N_11089);
or U15281 (N_15281,N_9123,N_8833);
nand U15282 (N_15282,N_8093,N_6624);
and U15283 (N_15283,N_10489,N_6747);
or U15284 (N_15284,N_8688,N_11440);
or U15285 (N_15285,N_10003,N_10131);
nand U15286 (N_15286,N_9417,N_10171);
or U15287 (N_15287,N_11198,N_6113);
and U15288 (N_15288,N_8454,N_7942);
or U15289 (N_15289,N_11953,N_9576);
and U15290 (N_15290,N_11397,N_9369);
xnor U15291 (N_15291,N_8652,N_8758);
and U15292 (N_15292,N_11861,N_6526);
nor U15293 (N_15293,N_8900,N_6669);
nor U15294 (N_15294,N_7942,N_10444);
xnor U15295 (N_15295,N_6673,N_7605);
nand U15296 (N_15296,N_6006,N_8283);
nand U15297 (N_15297,N_6541,N_7904);
and U15298 (N_15298,N_10378,N_8654);
xor U15299 (N_15299,N_11966,N_6535);
xnor U15300 (N_15300,N_10755,N_6404);
xor U15301 (N_15301,N_6755,N_6350);
or U15302 (N_15302,N_8449,N_11518);
or U15303 (N_15303,N_9272,N_6457);
nand U15304 (N_15304,N_11359,N_9362);
and U15305 (N_15305,N_9953,N_10933);
xnor U15306 (N_15306,N_11605,N_7926);
nand U15307 (N_15307,N_6381,N_11061);
nor U15308 (N_15308,N_11718,N_6139);
and U15309 (N_15309,N_10621,N_8468);
xnor U15310 (N_15310,N_9208,N_9377);
and U15311 (N_15311,N_10083,N_7620);
or U15312 (N_15312,N_7500,N_6479);
nand U15313 (N_15313,N_8285,N_7583);
nand U15314 (N_15314,N_7479,N_10191);
nor U15315 (N_15315,N_8386,N_6865);
and U15316 (N_15316,N_8216,N_8426);
and U15317 (N_15317,N_8033,N_10963);
and U15318 (N_15318,N_10461,N_9127);
nor U15319 (N_15319,N_11051,N_6371);
and U15320 (N_15320,N_9047,N_10835);
xor U15321 (N_15321,N_11057,N_11633);
nor U15322 (N_15322,N_9366,N_7268);
or U15323 (N_15323,N_10258,N_7098);
nand U15324 (N_15324,N_7665,N_9057);
nor U15325 (N_15325,N_7886,N_8750);
nor U15326 (N_15326,N_11464,N_9718);
xnor U15327 (N_15327,N_7624,N_6883);
nor U15328 (N_15328,N_6475,N_8852);
xnor U15329 (N_15329,N_8867,N_11502);
or U15330 (N_15330,N_8443,N_7049);
nor U15331 (N_15331,N_11116,N_10935);
nand U15332 (N_15332,N_6908,N_11075);
nor U15333 (N_15333,N_7659,N_10985);
or U15334 (N_15334,N_11282,N_8710);
nor U15335 (N_15335,N_10571,N_6254);
xnor U15336 (N_15336,N_7989,N_10660);
xor U15337 (N_15337,N_10411,N_9269);
and U15338 (N_15338,N_10617,N_11289);
and U15339 (N_15339,N_6878,N_11004);
nor U15340 (N_15340,N_6357,N_9687);
and U15341 (N_15341,N_8439,N_11937);
nand U15342 (N_15342,N_10800,N_11326);
or U15343 (N_15343,N_8703,N_7796);
or U15344 (N_15344,N_9781,N_6493);
nor U15345 (N_15345,N_11457,N_11106);
nand U15346 (N_15346,N_10876,N_9371);
and U15347 (N_15347,N_8376,N_9800);
nor U15348 (N_15348,N_9948,N_8431);
and U15349 (N_15349,N_6039,N_7422);
xor U15350 (N_15350,N_7642,N_9303);
nor U15351 (N_15351,N_11521,N_8306);
xor U15352 (N_15352,N_10573,N_9222);
or U15353 (N_15353,N_8313,N_11271);
or U15354 (N_15354,N_10337,N_11421);
nand U15355 (N_15355,N_6786,N_8957);
and U15356 (N_15356,N_7969,N_10679);
nor U15357 (N_15357,N_6851,N_9652);
nand U15358 (N_15358,N_7489,N_7346);
nor U15359 (N_15359,N_9401,N_7066);
or U15360 (N_15360,N_8444,N_6338);
and U15361 (N_15361,N_6179,N_10953);
or U15362 (N_15362,N_11916,N_7253);
nor U15363 (N_15363,N_10577,N_6184);
nor U15364 (N_15364,N_7895,N_8377);
nand U15365 (N_15365,N_8871,N_9397);
xnor U15366 (N_15366,N_7940,N_10132);
or U15367 (N_15367,N_6176,N_6338);
nor U15368 (N_15368,N_8222,N_8988);
and U15369 (N_15369,N_8534,N_6936);
or U15370 (N_15370,N_7520,N_6631);
and U15371 (N_15371,N_8045,N_10151);
xor U15372 (N_15372,N_9658,N_7419);
or U15373 (N_15373,N_6811,N_10756);
and U15374 (N_15374,N_8736,N_7883);
nand U15375 (N_15375,N_9084,N_10084);
xor U15376 (N_15376,N_11266,N_10727);
nor U15377 (N_15377,N_7549,N_9863);
nand U15378 (N_15378,N_7527,N_11821);
and U15379 (N_15379,N_7715,N_11483);
nor U15380 (N_15380,N_6793,N_7963);
nor U15381 (N_15381,N_7995,N_7433);
nand U15382 (N_15382,N_11259,N_8284);
or U15383 (N_15383,N_7041,N_11886);
nor U15384 (N_15384,N_11020,N_9544);
xnor U15385 (N_15385,N_11082,N_9386);
xnor U15386 (N_15386,N_7891,N_9511);
or U15387 (N_15387,N_7975,N_6064);
nand U15388 (N_15388,N_6095,N_7984);
and U15389 (N_15389,N_9002,N_7507);
nand U15390 (N_15390,N_11519,N_6562);
nor U15391 (N_15391,N_10810,N_8431);
nor U15392 (N_15392,N_11618,N_10832);
xor U15393 (N_15393,N_6577,N_7474);
nand U15394 (N_15394,N_10896,N_11113);
or U15395 (N_15395,N_11393,N_10029);
nor U15396 (N_15396,N_11639,N_8732);
nor U15397 (N_15397,N_7595,N_9690);
xnor U15398 (N_15398,N_7937,N_11513);
xor U15399 (N_15399,N_11298,N_11543);
or U15400 (N_15400,N_9880,N_11747);
xnor U15401 (N_15401,N_10357,N_10286);
or U15402 (N_15402,N_11101,N_10464);
nand U15403 (N_15403,N_8299,N_6331);
nand U15404 (N_15404,N_8012,N_7068);
nor U15405 (N_15405,N_9925,N_9940);
or U15406 (N_15406,N_9034,N_10611);
nand U15407 (N_15407,N_10486,N_9964);
xnor U15408 (N_15408,N_9730,N_7632);
nor U15409 (N_15409,N_11888,N_9369);
nor U15410 (N_15410,N_11992,N_6334);
or U15411 (N_15411,N_6421,N_9980);
or U15412 (N_15412,N_6057,N_9483);
nor U15413 (N_15413,N_7001,N_11810);
nand U15414 (N_15414,N_8266,N_9242);
xor U15415 (N_15415,N_7132,N_11133);
or U15416 (N_15416,N_7435,N_8650);
nand U15417 (N_15417,N_6762,N_9495);
and U15418 (N_15418,N_11658,N_7914);
nand U15419 (N_15419,N_10015,N_6821);
and U15420 (N_15420,N_8460,N_11100);
xnor U15421 (N_15421,N_8756,N_6294);
nand U15422 (N_15422,N_8334,N_6555);
nor U15423 (N_15423,N_7081,N_8567);
and U15424 (N_15424,N_10402,N_6612);
or U15425 (N_15425,N_9294,N_10264);
xnor U15426 (N_15426,N_8537,N_6133);
or U15427 (N_15427,N_7634,N_11671);
or U15428 (N_15428,N_7049,N_9451);
or U15429 (N_15429,N_7211,N_8492);
nand U15430 (N_15430,N_7292,N_10580);
or U15431 (N_15431,N_11815,N_6206);
nor U15432 (N_15432,N_8478,N_11559);
nor U15433 (N_15433,N_8459,N_8552);
xnor U15434 (N_15434,N_11826,N_10860);
xor U15435 (N_15435,N_6786,N_10990);
and U15436 (N_15436,N_7635,N_11982);
nand U15437 (N_15437,N_9261,N_6703);
nand U15438 (N_15438,N_10187,N_6276);
nand U15439 (N_15439,N_9817,N_9385);
xor U15440 (N_15440,N_6822,N_8293);
nand U15441 (N_15441,N_11937,N_8303);
nand U15442 (N_15442,N_8459,N_7448);
or U15443 (N_15443,N_9105,N_11821);
or U15444 (N_15444,N_9281,N_8449);
and U15445 (N_15445,N_9313,N_8577);
nand U15446 (N_15446,N_8670,N_6128);
xor U15447 (N_15447,N_7385,N_10768);
xnor U15448 (N_15448,N_11924,N_9892);
nand U15449 (N_15449,N_9696,N_8099);
or U15450 (N_15450,N_6656,N_11767);
nor U15451 (N_15451,N_11690,N_8801);
and U15452 (N_15452,N_7567,N_6646);
xnor U15453 (N_15453,N_8835,N_6919);
nor U15454 (N_15454,N_8924,N_11456);
and U15455 (N_15455,N_9606,N_7075);
nand U15456 (N_15456,N_11845,N_10095);
and U15457 (N_15457,N_6689,N_8215);
nand U15458 (N_15458,N_9064,N_11647);
xor U15459 (N_15459,N_8147,N_10575);
and U15460 (N_15460,N_6277,N_9410);
nor U15461 (N_15461,N_11320,N_11979);
and U15462 (N_15462,N_7930,N_9262);
or U15463 (N_15463,N_9805,N_7807);
and U15464 (N_15464,N_7451,N_8063);
xnor U15465 (N_15465,N_7112,N_9887);
nand U15466 (N_15466,N_6711,N_7877);
and U15467 (N_15467,N_10587,N_11483);
xnor U15468 (N_15468,N_9892,N_10395);
and U15469 (N_15469,N_10624,N_8427);
and U15470 (N_15470,N_10050,N_6731);
or U15471 (N_15471,N_9084,N_11603);
nand U15472 (N_15472,N_11625,N_8816);
or U15473 (N_15473,N_7695,N_7591);
and U15474 (N_15474,N_9000,N_8800);
xor U15475 (N_15475,N_8150,N_8479);
nor U15476 (N_15476,N_9528,N_9393);
or U15477 (N_15477,N_8232,N_8390);
nor U15478 (N_15478,N_7355,N_8664);
and U15479 (N_15479,N_7039,N_9031);
nor U15480 (N_15480,N_9371,N_11412);
nor U15481 (N_15481,N_11413,N_11236);
and U15482 (N_15482,N_9993,N_6516);
or U15483 (N_15483,N_8113,N_11780);
xor U15484 (N_15484,N_11444,N_9838);
or U15485 (N_15485,N_8160,N_9892);
xor U15486 (N_15486,N_7159,N_9176);
or U15487 (N_15487,N_7508,N_7449);
xor U15488 (N_15488,N_11708,N_6241);
nand U15489 (N_15489,N_6383,N_7259);
or U15490 (N_15490,N_6655,N_7086);
or U15491 (N_15491,N_9147,N_8172);
and U15492 (N_15492,N_8564,N_9039);
nand U15493 (N_15493,N_10432,N_11137);
nand U15494 (N_15494,N_8199,N_11218);
xor U15495 (N_15495,N_6755,N_8920);
xnor U15496 (N_15496,N_10180,N_10427);
nand U15497 (N_15497,N_11782,N_10028);
and U15498 (N_15498,N_8787,N_11360);
nor U15499 (N_15499,N_10329,N_7708);
or U15500 (N_15500,N_11188,N_10687);
nor U15501 (N_15501,N_11528,N_9235);
nand U15502 (N_15502,N_9574,N_6880);
and U15503 (N_15503,N_11922,N_8051);
or U15504 (N_15504,N_11444,N_7070);
nand U15505 (N_15505,N_6106,N_9590);
nand U15506 (N_15506,N_7562,N_11371);
nor U15507 (N_15507,N_11997,N_6571);
xnor U15508 (N_15508,N_8632,N_8885);
nand U15509 (N_15509,N_8952,N_9611);
nand U15510 (N_15510,N_8668,N_7359);
xor U15511 (N_15511,N_6645,N_8870);
and U15512 (N_15512,N_11928,N_11227);
nand U15513 (N_15513,N_7626,N_10853);
and U15514 (N_15514,N_6086,N_6432);
and U15515 (N_15515,N_8766,N_9064);
nor U15516 (N_15516,N_10962,N_9335);
and U15517 (N_15517,N_9984,N_9907);
nor U15518 (N_15518,N_9082,N_11605);
xnor U15519 (N_15519,N_7237,N_11005);
or U15520 (N_15520,N_9638,N_7589);
xnor U15521 (N_15521,N_11122,N_7918);
xor U15522 (N_15522,N_8049,N_8514);
nor U15523 (N_15523,N_7174,N_7740);
nor U15524 (N_15524,N_7584,N_10840);
or U15525 (N_15525,N_8889,N_10452);
nand U15526 (N_15526,N_10046,N_8963);
and U15527 (N_15527,N_6140,N_6610);
or U15528 (N_15528,N_9336,N_7877);
nor U15529 (N_15529,N_9968,N_8779);
xor U15530 (N_15530,N_9479,N_9012);
nor U15531 (N_15531,N_10444,N_11595);
and U15532 (N_15532,N_8505,N_11588);
nand U15533 (N_15533,N_10140,N_7279);
or U15534 (N_15534,N_10254,N_6749);
nor U15535 (N_15535,N_6963,N_7252);
xnor U15536 (N_15536,N_11158,N_7027);
nor U15537 (N_15537,N_6083,N_9076);
xor U15538 (N_15538,N_10263,N_9310);
nor U15539 (N_15539,N_8473,N_9325);
xnor U15540 (N_15540,N_8703,N_11589);
or U15541 (N_15541,N_6563,N_6643);
nand U15542 (N_15542,N_9926,N_11930);
xor U15543 (N_15543,N_8817,N_7084);
and U15544 (N_15544,N_7164,N_9972);
nor U15545 (N_15545,N_11151,N_8385);
and U15546 (N_15546,N_11455,N_9977);
or U15547 (N_15547,N_8202,N_11158);
xor U15548 (N_15548,N_8820,N_6715);
or U15549 (N_15549,N_11557,N_7931);
nand U15550 (N_15550,N_9439,N_11718);
or U15551 (N_15551,N_7394,N_8618);
or U15552 (N_15552,N_7625,N_6916);
nand U15553 (N_15553,N_10354,N_9887);
xor U15554 (N_15554,N_9325,N_11112);
and U15555 (N_15555,N_7194,N_11146);
nand U15556 (N_15556,N_7810,N_11224);
nor U15557 (N_15557,N_8112,N_8963);
and U15558 (N_15558,N_9276,N_7087);
nand U15559 (N_15559,N_7411,N_6416);
nand U15560 (N_15560,N_8137,N_10686);
or U15561 (N_15561,N_9612,N_9900);
and U15562 (N_15562,N_6130,N_11381);
nand U15563 (N_15563,N_8770,N_9553);
nand U15564 (N_15564,N_11439,N_10947);
nand U15565 (N_15565,N_9411,N_6581);
xor U15566 (N_15566,N_7525,N_6219);
nand U15567 (N_15567,N_10656,N_6135);
or U15568 (N_15568,N_8317,N_6498);
or U15569 (N_15569,N_9441,N_8668);
or U15570 (N_15570,N_8938,N_6690);
nand U15571 (N_15571,N_6866,N_11435);
and U15572 (N_15572,N_8408,N_9869);
or U15573 (N_15573,N_7119,N_6620);
nor U15574 (N_15574,N_9545,N_8912);
or U15575 (N_15575,N_7877,N_10977);
nor U15576 (N_15576,N_6877,N_7799);
and U15577 (N_15577,N_10614,N_7818);
and U15578 (N_15578,N_7345,N_9172);
or U15579 (N_15579,N_7616,N_8519);
and U15580 (N_15580,N_7689,N_9798);
or U15581 (N_15581,N_9639,N_10185);
nor U15582 (N_15582,N_7828,N_10052);
nand U15583 (N_15583,N_10636,N_10047);
xor U15584 (N_15584,N_9564,N_8349);
or U15585 (N_15585,N_10077,N_6341);
nor U15586 (N_15586,N_9870,N_10238);
xor U15587 (N_15587,N_10806,N_11517);
nor U15588 (N_15588,N_8254,N_7891);
nor U15589 (N_15589,N_7882,N_7675);
nand U15590 (N_15590,N_9192,N_8862);
and U15591 (N_15591,N_6326,N_10573);
nand U15592 (N_15592,N_9868,N_8548);
nand U15593 (N_15593,N_9591,N_11500);
or U15594 (N_15594,N_10534,N_6039);
or U15595 (N_15595,N_8549,N_11327);
xnor U15596 (N_15596,N_6718,N_7951);
or U15597 (N_15597,N_8830,N_9573);
xor U15598 (N_15598,N_6418,N_10066);
and U15599 (N_15599,N_9863,N_8949);
xor U15600 (N_15600,N_10813,N_11379);
xnor U15601 (N_15601,N_9388,N_8466);
nand U15602 (N_15602,N_6835,N_9207);
nor U15603 (N_15603,N_9630,N_9169);
xor U15604 (N_15604,N_8495,N_10401);
and U15605 (N_15605,N_6680,N_10982);
nand U15606 (N_15606,N_7183,N_8576);
or U15607 (N_15607,N_8035,N_10573);
nor U15608 (N_15608,N_11228,N_7029);
xor U15609 (N_15609,N_10440,N_6871);
and U15610 (N_15610,N_8108,N_6396);
nand U15611 (N_15611,N_7077,N_8531);
and U15612 (N_15612,N_10613,N_10522);
nor U15613 (N_15613,N_6776,N_7693);
xnor U15614 (N_15614,N_11497,N_8612);
and U15615 (N_15615,N_8784,N_6904);
nor U15616 (N_15616,N_11284,N_6626);
or U15617 (N_15617,N_10521,N_10063);
nand U15618 (N_15618,N_11336,N_9082);
xor U15619 (N_15619,N_9613,N_7869);
and U15620 (N_15620,N_6561,N_9468);
and U15621 (N_15621,N_10476,N_7870);
xor U15622 (N_15622,N_8175,N_10770);
or U15623 (N_15623,N_8629,N_7955);
nor U15624 (N_15624,N_8966,N_6015);
or U15625 (N_15625,N_11832,N_7477);
nand U15626 (N_15626,N_10124,N_8959);
nand U15627 (N_15627,N_7709,N_8562);
nor U15628 (N_15628,N_6766,N_6320);
and U15629 (N_15629,N_7657,N_7300);
and U15630 (N_15630,N_10746,N_9605);
nand U15631 (N_15631,N_11755,N_10795);
or U15632 (N_15632,N_7814,N_6670);
nand U15633 (N_15633,N_8943,N_6419);
or U15634 (N_15634,N_6176,N_10809);
xnor U15635 (N_15635,N_10414,N_11468);
xor U15636 (N_15636,N_11307,N_9302);
or U15637 (N_15637,N_7613,N_7066);
xor U15638 (N_15638,N_6523,N_9909);
nand U15639 (N_15639,N_9642,N_8389);
xnor U15640 (N_15640,N_10738,N_9328);
nor U15641 (N_15641,N_11446,N_6206);
xnor U15642 (N_15642,N_10739,N_8423);
nand U15643 (N_15643,N_7501,N_7529);
and U15644 (N_15644,N_11389,N_6513);
and U15645 (N_15645,N_8786,N_10936);
nor U15646 (N_15646,N_10536,N_8114);
nor U15647 (N_15647,N_6775,N_9699);
xor U15648 (N_15648,N_8724,N_6549);
nand U15649 (N_15649,N_9771,N_10059);
and U15650 (N_15650,N_9306,N_10513);
xor U15651 (N_15651,N_9448,N_11480);
nor U15652 (N_15652,N_6698,N_9755);
or U15653 (N_15653,N_10652,N_6414);
nor U15654 (N_15654,N_7020,N_10586);
nor U15655 (N_15655,N_7815,N_9680);
or U15656 (N_15656,N_10144,N_8396);
xor U15657 (N_15657,N_8374,N_11000);
nor U15658 (N_15658,N_7564,N_11674);
nand U15659 (N_15659,N_10625,N_6059);
and U15660 (N_15660,N_10932,N_8243);
nor U15661 (N_15661,N_10156,N_6198);
nand U15662 (N_15662,N_6552,N_6762);
xnor U15663 (N_15663,N_7504,N_6929);
or U15664 (N_15664,N_10628,N_6094);
nand U15665 (N_15665,N_9665,N_10880);
nand U15666 (N_15666,N_9449,N_6405);
nor U15667 (N_15667,N_11226,N_8122);
xnor U15668 (N_15668,N_6837,N_8600);
xnor U15669 (N_15669,N_10922,N_6866);
and U15670 (N_15670,N_10803,N_6947);
or U15671 (N_15671,N_11240,N_9853);
and U15672 (N_15672,N_11720,N_7969);
or U15673 (N_15673,N_10098,N_9618);
or U15674 (N_15674,N_11371,N_9497);
nand U15675 (N_15675,N_6070,N_10376);
and U15676 (N_15676,N_9773,N_6743);
nand U15677 (N_15677,N_9518,N_6204);
or U15678 (N_15678,N_6431,N_7475);
xnor U15679 (N_15679,N_7784,N_7696);
and U15680 (N_15680,N_9975,N_9079);
or U15681 (N_15681,N_8502,N_10577);
nor U15682 (N_15682,N_8238,N_8056);
and U15683 (N_15683,N_7901,N_11131);
xnor U15684 (N_15684,N_8162,N_9900);
xnor U15685 (N_15685,N_10413,N_10683);
nand U15686 (N_15686,N_9211,N_8922);
xnor U15687 (N_15687,N_7669,N_8868);
xnor U15688 (N_15688,N_8551,N_7866);
nand U15689 (N_15689,N_8153,N_10892);
nor U15690 (N_15690,N_8065,N_9608);
nand U15691 (N_15691,N_7708,N_11408);
nand U15692 (N_15692,N_6830,N_10336);
nand U15693 (N_15693,N_9118,N_7758);
nand U15694 (N_15694,N_7211,N_8491);
nand U15695 (N_15695,N_11388,N_7905);
and U15696 (N_15696,N_11440,N_8503);
and U15697 (N_15697,N_9640,N_10952);
xor U15698 (N_15698,N_6065,N_10118);
xnor U15699 (N_15699,N_11530,N_7440);
or U15700 (N_15700,N_6612,N_7864);
nand U15701 (N_15701,N_9906,N_7219);
xor U15702 (N_15702,N_6689,N_8642);
nand U15703 (N_15703,N_7372,N_9095);
or U15704 (N_15704,N_8347,N_11653);
nand U15705 (N_15705,N_8200,N_6349);
nand U15706 (N_15706,N_10832,N_8897);
xnor U15707 (N_15707,N_6410,N_11137);
nor U15708 (N_15708,N_6337,N_7578);
and U15709 (N_15709,N_6696,N_11133);
nor U15710 (N_15710,N_8097,N_11195);
nor U15711 (N_15711,N_6758,N_6141);
and U15712 (N_15712,N_11179,N_7234);
nor U15713 (N_15713,N_9919,N_10301);
and U15714 (N_15714,N_11340,N_10425);
nor U15715 (N_15715,N_9521,N_11568);
nand U15716 (N_15716,N_9665,N_6539);
nor U15717 (N_15717,N_7890,N_11565);
or U15718 (N_15718,N_11107,N_10388);
nand U15719 (N_15719,N_7576,N_7482);
xor U15720 (N_15720,N_6628,N_8696);
nor U15721 (N_15721,N_8170,N_11440);
nor U15722 (N_15722,N_11422,N_10104);
nand U15723 (N_15723,N_7825,N_9381);
and U15724 (N_15724,N_8277,N_6825);
nand U15725 (N_15725,N_9860,N_7199);
nand U15726 (N_15726,N_10587,N_11783);
nand U15727 (N_15727,N_9569,N_7387);
xor U15728 (N_15728,N_10959,N_8016);
nand U15729 (N_15729,N_8636,N_11755);
and U15730 (N_15730,N_7786,N_9446);
nand U15731 (N_15731,N_10492,N_8828);
nand U15732 (N_15732,N_8216,N_8796);
nand U15733 (N_15733,N_9090,N_10527);
nand U15734 (N_15734,N_8839,N_7139);
nand U15735 (N_15735,N_6602,N_6113);
nor U15736 (N_15736,N_8464,N_7727);
and U15737 (N_15737,N_10611,N_9385);
or U15738 (N_15738,N_11271,N_8823);
or U15739 (N_15739,N_6420,N_8945);
nand U15740 (N_15740,N_8166,N_6271);
nor U15741 (N_15741,N_7191,N_9067);
nor U15742 (N_15742,N_6618,N_8399);
nand U15743 (N_15743,N_8461,N_10402);
and U15744 (N_15744,N_6858,N_10272);
xnor U15745 (N_15745,N_9907,N_11905);
nand U15746 (N_15746,N_6576,N_6704);
and U15747 (N_15747,N_8394,N_7446);
and U15748 (N_15748,N_10203,N_8320);
and U15749 (N_15749,N_8693,N_7559);
nor U15750 (N_15750,N_7000,N_6951);
and U15751 (N_15751,N_7971,N_11289);
nor U15752 (N_15752,N_11318,N_9257);
xor U15753 (N_15753,N_6413,N_9669);
xnor U15754 (N_15754,N_8059,N_7731);
or U15755 (N_15755,N_7527,N_9729);
or U15756 (N_15756,N_9727,N_7473);
xnor U15757 (N_15757,N_9627,N_10852);
nand U15758 (N_15758,N_11057,N_8926);
and U15759 (N_15759,N_7940,N_8476);
and U15760 (N_15760,N_9766,N_11131);
nor U15761 (N_15761,N_10261,N_8852);
nor U15762 (N_15762,N_9355,N_6887);
nand U15763 (N_15763,N_10029,N_11942);
nor U15764 (N_15764,N_10851,N_11174);
nor U15765 (N_15765,N_11232,N_8559);
nand U15766 (N_15766,N_7569,N_6332);
and U15767 (N_15767,N_11085,N_6986);
nand U15768 (N_15768,N_8651,N_11190);
nor U15769 (N_15769,N_7708,N_6712);
or U15770 (N_15770,N_6470,N_6145);
or U15771 (N_15771,N_7465,N_9067);
nor U15772 (N_15772,N_7741,N_7307);
xor U15773 (N_15773,N_7894,N_7912);
nor U15774 (N_15774,N_11184,N_10635);
nand U15775 (N_15775,N_8065,N_10724);
xor U15776 (N_15776,N_7902,N_11045);
and U15777 (N_15777,N_7889,N_9698);
nand U15778 (N_15778,N_10943,N_8276);
or U15779 (N_15779,N_11655,N_6145);
and U15780 (N_15780,N_10858,N_9242);
or U15781 (N_15781,N_9416,N_6888);
xor U15782 (N_15782,N_8754,N_9911);
and U15783 (N_15783,N_10211,N_9822);
nor U15784 (N_15784,N_8344,N_7795);
xor U15785 (N_15785,N_10434,N_8668);
and U15786 (N_15786,N_8247,N_8769);
and U15787 (N_15787,N_10295,N_8019);
and U15788 (N_15788,N_11242,N_6318);
nor U15789 (N_15789,N_11959,N_8608);
and U15790 (N_15790,N_7724,N_7981);
or U15791 (N_15791,N_8550,N_10568);
nor U15792 (N_15792,N_6281,N_7338);
or U15793 (N_15793,N_6474,N_7863);
or U15794 (N_15794,N_7626,N_11588);
xor U15795 (N_15795,N_8534,N_11290);
and U15796 (N_15796,N_9942,N_8333);
nand U15797 (N_15797,N_7406,N_10252);
and U15798 (N_15798,N_7568,N_7269);
and U15799 (N_15799,N_6362,N_10373);
xnor U15800 (N_15800,N_6380,N_8074);
or U15801 (N_15801,N_10210,N_11392);
xnor U15802 (N_15802,N_6882,N_10666);
xnor U15803 (N_15803,N_10813,N_6220);
nand U15804 (N_15804,N_11205,N_9743);
nor U15805 (N_15805,N_6543,N_8990);
and U15806 (N_15806,N_9595,N_8444);
or U15807 (N_15807,N_7847,N_6981);
nand U15808 (N_15808,N_6552,N_6538);
xnor U15809 (N_15809,N_10644,N_8466);
nor U15810 (N_15810,N_7237,N_10895);
nand U15811 (N_15811,N_11807,N_6856);
nand U15812 (N_15812,N_7768,N_11083);
xor U15813 (N_15813,N_8477,N_7660);
and U15814 (N_15814,N_8575,N_7423);
xnor U15815 (N_15815,N_6345,N_9751);
and U15816 (N_15816,N_8878,N_7547);
nand U15817 (N_15817,N_11118,N_10376);
or U15818 (N_15818,N_7688,N_8394);
and U15819 (N_15819,N_9226,N_7743);
and U15820 (N_15820,N_10898,N_9410);
xnor U15821 (N_15821,N_11891,N_10393);
nor U15822 (N_15822,N_7242,N_10323);
or U15823 (N_15823,N_6469,N_11121);
nand U15824 (N_15824,N_11580,N_8346);
nand U15825 (N_15825,N_7422,N_9027);
xnor U15826 (N_15826,N_9449,N_9093);
nor U15827 (N_15827,N_7018,N_11455);
or U15828 (N_15828,N_8791,N_9039);
nand U15829 (N_15829,N_10082,N_11112);
and U15830 (N_15830,N_8789,N_7708);
xor U15831 (N_15831,N_9821,N_6509);
xnor U15832 (N_15832,N_11734,N_8598);
and U15833 (N_15833,N_6425,N_6338);
or U15834 (N_15834,N_8134,N_11296);
nor U15835 (N_15835,N_11062,N_8848);
and U15836 (N_15836,N_11701,N_8344);
nor U15837 (N_15837,N_8890,N_9700);
or U15838 (N_15838,N_8996,N_9523);
nor U15839 (N_15839,N_11439,N_7540);
xnor U15840 (N_15840,N_7606,N_8324);
or U15841 (N_15841,N_6588,N_6479);
and U15842 (N_15842,N_8792,N_9877);
and U15843 (N_15843,N_9991,N_10580);
and U15844 (N_15844,N_6788,N_8615);
xnor U15845 (N_15845,N_10746,N_7474);
or U15846 (N_15846,N_10553,N_10955);
xnor U15847 (N_15847,N_8665,N_8866);
xor U15848 (N_15848,N_8202,N_8120);
or U15849 (N_15849,N_7171,N_9248);
xor U15850 (N_15850,N_6443,N_9332);
and U15851 (N_15851,N_9823,N_8218);
nor U15852 (N_15852,N_8148,N_11420);
nand U15853 (N_15853,N_11567,N_8861);
or U15854 (N_15854,N_10156,N_8486);
and U15855 (N_15855,N_6969,N_7976);
and U15856 (N_15856,N_8000,N_6007);
or U15857 (N_15857,N_7249,N_11786);
or U15858 (N_15858,N_6352,N_9784);
nor U15859 (N_15859,N_11498,N_8750);
xnor U15860 (N_15860,N_10575,N_9134);
nor U15861 (N_15861,N_7536,N_6459);
nor U15862 (N_15862,N_11058,N_11203);
xnor U15863 (N_15863,N_9096,N_8112);
and U15864 (N_15864,N_6860,N_8948);
xnor U15865 (N_15865,N_11608,N_9143);
xnor U15866 (N_15866,N_6457,N_6456);
nand U15867 (N_15867,N_10012,N_6522);
nor U15868 (N_15868,N_7865,N_9257);
nor U15869 (N_15869,N_6569,N_8982);
xnor U15870 (N_15870,N_10728,N_6404);
or U15871 (N_15871,N_6834,N_8529);
nor U15872 (N_15872,N_8201,N_7335);
or U15873 (N_15873,N_8216,N_7055);
nand U15874 (N_15874,N_6071,N_7023);
and U15875 (N_15875,N_9436,N_7412);
nand U15876 (N_15876,N_11543,N_7161);
and U15877 (N_15877,N_6884,N_11068);
xor U15878 (N_15878,N_11827,N_6685);
or U15879 (N_15879,N_11057,N_7295);
nor U15880 (N_15880,N_7689,N_6353);
nand U15881 (N_15881,N_8735,N_9137);
xnor U15882 (N_15882,N_7745,N_11382);
nand U15883 (N_15883,N_10330,N_6093);
nor U15884 (N_15884,N_6882,N_11429);
nand U15885 (N_15885,N_6893,N_6681);
nor U15886 (N_15886,N_10864,N_8224);
or U15887 (N_15887,N_8422,N_6712);
nand U15888 (N_15888,N_7317,N_6341);
nor U15889 (N_15889,N_9480,N_7347);
or U15890 (N_15890,N_10478,N_8422);
nor U15891 (N_15891,N_7373,N_11414);
xnor U15892 (N_15892,N_11002,N_10901);
or U15893 (N_15893,N_10024,N_9866);
and U15894 (N_15894,N_7154,N_11420);
xnor U15895 (N_15895,N_9452,N_8492);
xnor U15896 (N_15896,N_9855,N_6845);
nand U15897 (N_15897,N_10079,N_9837);
or U15898 (N_15898,N_8614,N_11085);
or U15899 (N_15899,N_11222,N_6940);
nand U15900 (N_15900,N_11946,N_8078);
xor U15901 (N_15901,N_10518,N_11732);
xor U15902 (N_15902,N_10738,N_8593);
and U15903 (N_15903,N_8115,N_7458);
xnor U15904 (N_15904,N_6096,N_11560);
and U15905 (N_15905,N_8531,N_6994);
nor U15906 (N_15906,N_10272,N_11370);
and U15907 (N_15907,N_11933,N_6911);
xnor U15908 (N_15908,N_11997,N_7856);
nand U15909 (N_15909,N_9028,N_9074);
nor U15910 (N_15910,N_11957,N_8355);
nor U15911 (N_15911,N_9798,N_7405);
nor U15912 (N_15912,N_8854,N_8243);
nor U15913 (N_15913,N_9473,N_7030);
and U15914 (N_15914,N_8261,N_7890);
nor U15915 (N_15915,N_10169,N_11241);
nand U15916 (N_15916,N_8532,N_9712);
nand U15917 (N_15917,N_8131,N_9334);
or U15918 (N_15918,N_9276,N_6422);
nor U15919 (N_15919,N_6720,N_10747);
nand U15920 (N_15920,N_6480,N_11636);
and U15921 (N_15921,N_6971,N_11044);
nand U15922 (N_15922,N_10359,N_7162);
xor U15923 (N_15923,N_9491,N_6508);
and U15924 (N_15924,N_10663,N_6424);
nor U15925 (N_15925,N_9062,N_11018);
and U15926 (N_15926,N_7904,N_7104);
nand U15927 (N_15927,N_6027,N_9020);
nand U15928 (N_15928,N_10864,N_9452);
nor U15929 (N_15929,N_11647,N_6712);
or U15930 (N_15930,N_11385,N_6541);
nor U15931 (N_15931,N_7431,N_11624);
nand U15932 (N_15932,N_11999,N_10010);
or U15933 (N_15933,N_11538,N_10382);
and U15934 (N_15934,N_8004,N_10463);
nand U15935 (N_15935,N_10538,N_7485);
nand U15936 (N_15936,N_10745,N_6639);
xor U15937 (N_15937,N_8089,N_6083);
xnor U15938 (N_15938,N_10745,N_6335);
nor U15939 (N_15939,N_8484,N_11927);
xor U15940 (N_15940,N_10030,N_11925);
xor U15941 (N_15941,N_8998,N_11956);
nand U15942 (N_15942,N_7139,N_10925);
or U15943 (N_15943,N_8627,N_8275);
or U15944 (N_15944,N_9615,N_7477);
nand U15945 (N_15945,N_8359,N_11612);
nand U15946 (N_15946,N_10718,N_10619);
and U15947 (N_15947,N_10980,N_10999);
nand U15948 (N_15948,N_6007,N_6524);
xor U15949 (N_15949,N_11129,N_7998);
nor U15950 (N_15950,N_7020,N_11847);
or U15951 (N_15951,N_9195,N_9289);
nand U15952 (N_15952,N_11322,N_7087);
and U15953 (N_15953,N_10933,N_6436);
and U15954 (N_15954,N_6058,N_11795);
or U15955 (N_15955,N_10811,N_11223);
and U15956 (N_15956,N_8034,N_9366);
nor U15957 (N_15957,N_10209,N_11693);
and U15958 (N_15958,N_7904,N_6768);
nand U15959 (N_15959,N_7636,N_7935);
and U15960 (N_15960,N_6391,N_11439);
and U15961 (N_15961,N_8294,N_11081);
nor U15962 (N_15962,N_9487,N_9473);
or U15963 (N_15963,N_10596,N_9557);
nor U15964 (N_15964,N_8969,N_7817);
xnor U15965 (N_15965,N_8764,N_7405);
or U15966 (N_15966,N_8643,N_11596);
and U15967 (N_15967,N_6688,N_6658);
nor U15968 (N_15968,N_10075,N_7556);
or U15969 (N_15969,N_10212,N_11175);
nor U15970 (N_15970,N_8164,N_11366);
xnor U15971 (N_15971,N_8057,N_11223);
xor U15972 (N_15972,N_9036,N_8806);
and U15973 (N_15973,N_6313,N_10690);
nor U15974 (N_15974,N_8544,N_7844);
nand U15975 (N_15975,N_8064,N_8020);
nor U15976 (N_15976,N_11104,N_6872);
nand U15977 (N_15977,N_7273,N_6467);
and U15978 (N_15978,N_11897,N_8012);
nor U15979 (N_15979,N_9495,N_10168);
nand U15980 (N_15980,N_9873,N_8150);
xor U15981 (N_15981,N_9776,N_11093);
nor U15982 (N_15982,N_10558,N_6328);
nand U15983 (N_15983,N_10800,N_8472);
or U15984 (N_15984,N_11379,N_11277);
nor U15985 (N_15985,N_11568,N_11515);
nor U15986 (N_15986,N_9897,N_11420);
or U15987 (N_15987,N_7346,N_10941);
or U15988 (N_15988,N_11038,N_7819);
and U15989 (N_15989,N_8369,N_7657);
nand U15990 (N_15990,N_6905,N_9017);
nand U15991 (N_15991,N_6095,N_7172);
or U15992 (N_15992,N_10513,N_11895);
nand U15993 (N_15993,N_9204,N_6393);
xor U15994 (N_15994,N_11057,N_10986);
and U15995 (N_15995,N_6003,N_7307);
and U15996 (N_15996,N_6007,N_7686);
nand U15997 (N_15997,N_6772,N_9726);
nand U15998 (N_15998,N_10860,N_11757);
and U15999 (N_15999,N_7909,N_10198);
nand U16000 (N_16000,N_9064,N_10726);
nand U16001 (N_16001,N_9169,N_8226);
nor U16002 (N_16002,N_9864,N_11976);
or U16003 (N_16003,N_6285,N_10752);
xor U16004 (N_16004,N_7449,N_11885);
xnor U16005 (N_16005,N_8743,N_7476);
xor U16006 (N_16006,N_6495,N_11038);
nor U16007 (N_16007,N_6090,N_7795);
nand U16008 (N_16008,N_9732,N_9729);
xnor U16009 (N_16009,N_7689,N_6334);
nor U16010 (N_16010,N_10455,N_6437);
xnor U16011 (N_16011,N_8990,N_8101);
nor U16012 (N_16012,N_11207,N_9488);
nand U16013 (N_16013,N_8289,N_11084);
xor U16014 (N_16014,N_11868,N_10442);
nand U16015 (N_16015,N_10697,N_10124);
nor U16016 (N_16016,N_6762,N_7268);
and U16017 (N_16017,N_9179,N_10404);
xnor U16018 (N_16018,N_6249,N_11584);
nand U16019 (N_16019,N_7127,N_6429);
xor U16020 (N_16020,N_10678,N_10374);
nor U16021 (N_16021,N_9743,N_7351);
nand U16022 (N_16022,N_10945,N_11654);
or U16023 (N_16023,N_9083,N_11507);
nand U16024 (N_16024,N_8333,N_9094);
xor U16025 (N_16025,N_7570,N_9948);
and U16026 (N_16026,N_11428,N_11119);
nand U16027 (N_16027,N_10226,N_9160);
nor U16028 (N_16028,N_7355,N_11733);
nor U16029 (N_16029,N_9737,N_6096);
xor U16030 (N_16030,N_9741,N_10659);
nor U16031 (N_16031,N_6640,N_11525);
and U16032 (N_16032,N_10255,N_11829);
xnor U16033 (N_16033,N_7579,N_10917);
and U16034 (N_16034,N_10774,N_8412);
and U16035 (N_16035,N_6461,N_10073);
or U16036 (N_16036,N_11853,N_6643);
nand U16037 (N_16037,N_10709,N_10153);
xor U16038 (N_16038,N_9286,N_11232);
nand U16039 (N_16039,N_11638,N_6809);
nand U16040 (N_16040,N_10447,N_10763);
or U16041 (N_16041,N_9166,N_7535);
xor U16042 (N_16042,N_11910,N_9515);
nand U16043 (N_16043,N_10157,N_9053);
nand U16044 (N_16044,N_8492,N_10228);
nor U16045 (N_16045,N_10728,N_8842);
or U16046 (N_16046,N_8514,N_11576);
nor U16047 (N_16047,N_6374,N_8319);
nor U16048 (N_16048,N_9030,N_8849);
nor U16049 (N_16049,N_6532,N_11467);
xnor U16050 (N_16050,N_9243,N_11718);
nand U16051 (N_16051,N_9277,N_11532);
or U16052 (N_16052,N_9489,N_7871);
and U16053 (N_16053,N_6296,N_10789);
and U16054 (N_16054,N_10132,N_8900);
nor U16055 (N_16055,N_11670,N_6824);
xnor U16056 (N_16056,N_10540,N_7623);
nand U16057 (N_16057,N_7280,N_9080);
nor U16058 (N_16058,N_8816,N_8705);
or U16059 (N_16059,N_8378,N_10108);
nor U16060 (N_16060,N_11120,N_6650);
and U16061 (N_16061,N_8910,N_7384);
nor U16062 (N_16062,N_7875,N_11386);
nand U16063 (N_16063,N_9209,N_8533);
and U16064 (N_16064,N_7241,N_6050);
xor U16065 (N_16065,N_11846,N_6331);
nand U16066 (N_16066,N_7705,N_10413);
or U16067 (N_16067,N_7470,N_7221);
or U16068 (N_16068,N_10756,N_11657);
or U16069 (N_16069,N_10912,N_8462);
and U16070 (N_16070,N_7046,N_11422);
nand U16071 (N_16071,N_8062,N_6287);
or U16072 (N_16072,N_9271,N_8449);
nor U16073 (N_16073,N_9843,N_10420);
xnor U16074 (N_16074,N_10944,N_6568);
xnor U16075 (N_16075,N_9307,N_10659);
or U16076 (N_16076,N_8909,N_10468);
nor U16077 (N_16077,N_7085,N_11134);
or U16078 (N_16078,N_11334,N_7132);
and U16079 (N_16079,N_7111,N_6412);
or U16080 (N_16080,N_8410,N_8152);
or U16081 (N_16081,N_9935,N_11177);
and U16082 (N_16082,N_11335,N_7050);
xor U16083 (N_16083,N_11395,N_11125);
nand U16084 (N_16084,N_8251,N_10186);
and U16085 (N_16085,N_11198,N_6961);
or U16086 (N_16086,N_10098,N_8345);
nand U16087 (N_16087,N_6577,N_7564);
nor U16088 (N_16088,N_10125,N_8385);
xnor U16089 (N_16089,N_6311,N_9521);
or U16090 (N_16090,N_10307,N_9594);
nor U16091 (N_16091,N_8694,N_6130);
nor U16092 (N_16092,N_9352,N_8489);
xnor U16093 (N_16093,N_11757,N_8427);
xor U16094 (N_16094,N_6671,N_11763);
or U16095 (N_16095,N_9436,N_6064);
and U16096 (N_16096,N_7561,N_8942);
nand U16097 (N_16097,N_11028,N_9850);
nor U16098 (N_16098,N_11459,N_11774);
xor U16099 (N_16099,N_9434,N_6992);
and U16100 (N_16100,N_9462,N_7176);
nand U16101 (N_16101,N_10289,N_8724);
nand U16102 (N_16102,N_9422,N_11615);
or U16103 (N_16103,N_6259,N_10754);
xnor U16104 (N_16104,N_7728,N_11101);
or U16105 (N_16105,N_11949,N_6104);
xor U16106 (N_16106,N_6348,N_8203);
nor U16107 (N_16107,N_6644,N_7492);
nand U16108 (N_16108,N_8205,N_6122);
nor U16109 (N_16109,N_11691,N_9116);
nand U16110 (N_16110,N_9458,N_11171);
xor U16111 (N_16111,N_6184,N_6953);
or U16112 (N_16112,N_9548,N_9611);
or U16113 (N_16113,N_11244,N_7709);
xor U16114 (N_16114,N_9972,N_10678);
xnor U16115 (N_16115,N_7260,N_8828);
xnor U16116 (N_16116,N_10881,N_10042);
nor U16117 (N_16117,N_10260,N_7692);
nand U16118 (N_16118,N_9319,N_9422);
or U16119 (N_16119,N_11649,N_6449);
nor U16120 (N_16120,N_10834,N_9626);
nor U16121 (N_16121,N_10264,N_11495);
or U16122 (N_16122,N_6855,N_10619);
or U16123 (N_16123,N_11330,N_8158);
nor U16124 (N_16124,N_8037,N_10043);
and U16125 (N_16125,N_7255,N_11198);
and U16126 (N_16126,N_7730,N_9151);
xnor U16127 (N_16127,N_6868,N_6554);
and U16128 (N_16128,N_8360,N_6821);
xor U16129 (N_16129,N_10911,N_11484);
and U16130 (N_16130,N_9135,N_6173);
nor U16131 (N_16131,N_7096,N_10057);
and U16132 (N_16132,N_6145,N_9161);
and U16133 (N_16133,N_11121,N_7281);
nor U16134 (N_16134,N_6324,N_7070);
and U16135 (N_16135,N_7148,N_10569);
nand U16136 (N_16136,N_7625,N_7994);
or U16137 (N_16137,N_9857,N_10587);
and U16138 (N_16138,N_7998,N_10520);
and U16139 (N_16139,N_8752,N_11495);
or U16140 (N_16140,N_7829,N_7526);
or U16141 (N_16141,N_6096,N_7628);
nand U16142 (N_16142,N_7086,N_11569);
and U16143 (N_16143,N_7824,N_7900);
nor U16144 (N_16144,N_6605,N_10358);
nand U16145 (N_16145,N_9308,N_7330);
or U16146 (N_16146,N_10938,N_8724);
nand U16147 (N_16147,N_8303,N_10657);
xnor U16148 (N_16148,N_8450,N_11970);
nor U16149 (N_16149,N_11356,N_7924);
and U16150 (N_16150,N_11864,N_6371);
xnor U16151 (N_16151,N_7879,N_9033);
xnor U16152 (N_16152,N_9706,N_6841);
nand U16153 (N_16153,N_11204,N_10615);
nor U16154 (N_16154,N_9565,N_10057);
nand U16155 (N_16155,N_9731,N_7527);
and U16156 (N_16156,N_9027,N_8884);
nor U16157 (N_16157,N_8470,N_8350);
xnor U16158 (N_16158,N_11666,N_9119);
nand U16159 (N_16159,N_9410,N_9125);
and U16160 (N_16160,N_8635,N_7577);
or U16161 (N_16161,N_7561,N_7424);
or U16162 (N_16162,N_11769,N_7083);
nor U16163 (N_16163,N_6940,N_9791);
or U16164 (N_16164,N_9873,N_10069);
and U16165 (N_16165,N_6724,N_8846);
nor U16166 (N_16166,N_7643,N_11214);
or U16167 (N_16167,N_8993,N_7479);
nand U16168 (N_16168,N_9064,N_11005);
or U16169 (N_16169,N_9566,N_10363);
or U16170 (N_16170,N_9380,N_8661);
xor U16171 (N_16171,N_6315,N_10010);
nand U16172 (N_16172,N_10478,N_8752);
xor U16173 (N_16173,N_6842,N_8147);
and U16174 (N_16174,N_7704,N_8417);
xor U16175 (N_16175,N_11094,N_8645);
and U16176 (N_16176,N_11266,N_10455);
nor U16177 (N_16177,N_7069,N_6325);
nor U16178 (N_16178,N_9637,N_11279);
xor U16179 (N_16179,N_8605,N_6423);
nor U16180 (N_16180,N_6267,N_11643);
xnor U16181 (N_16181,N_7809,N_8061);
or U16182 (N_16182,N_10687,N_6791);
nor U16183 (N_16183,N_7312,N_8235);
nand U16184 (N_16184,N_8190,N_9157);
and U16185 (N_16185,N_10527,N_10364);
xnor U16186 (N_16186,N_7294,N_7037);
or U16187 (N_16187,N_7957,N_7233);
xnor U16188 (N_16188,N_7121,N_8439);
or U16189 (N_16189,N_9035,N_8867);
xnor U16190 (N_16190,N_11988,N_10336);
and U16191 (N_16191,N_9796,N_6370);
nor U16192 (N_16192,N_9924,N_6460);
or U16193 (N_16193,N_8626,N_8645);
xor U16194 (N_16194,N_10209,N_6733);
nand U16195 (N_16195,N_9607,N_11803);
xnor U16196 (N_16196,N_10302,N_9662);
or U16197 (N_16197,N_6032,N_8621);
and U16198 (N_16198,N_10016,N_6193);
nor U16199 (N_16199,N_6187,N_9663);
nand U16200 (N_16200,N_11459,N_6343);
nand U16201 (N_16201,N_10078,N_8592);
nor U16202 (N_16202,N_7136,N_8442);
nor U16203 (N_16203,N_11250,N_9504);
and U16204 (N_16204,N_7441,N_8853);
nand U16205 (N_16205,N_9158,N_10066);
and U16206 (N_16206,N_9735,N_7257);
xor U16207 (N_16207,N_10460,N_6015);
or U16208 (N_16208,N_6069,N_7367);
xor U16209 (N_16209,N_10848,N_7862);
xnor U16210 (N_16210,N_9925,N_6513);
nor U16211 (N_16211,N_8851,N_6554);
nand U16212 (N_16212,N_11074,N_7025);
nor U16213 (N_16213,N_7238,N_9256);
nand U16214 (N_16214,N_7653,N_7434);
nor U16215 (N_16215,N_6978,N_10661);
xnor U16216 (N_16216,N_6944,N_11967);
nor U16217 (N_16217,N_7653,N_7477);
and U16218 (N_16218,N_6401,N_10721);
xor U16219 (N_16219,N_6590,N_6880);
or U16220 (N_16220,N_11168,N_9789);
or U16221 (N_16221,N_9008,N_9453);
xnor U16222 (N_16222,N_10117,N_6179);
xor U16223 (N_16223,N_10042,N_9391);
nand U16224 (N_16224,N_9160,N_9755);
or U16225 (N_16225,N_9000,N_11352);
and U16226 (N_16226,N_10024,N_11028);
nor U16227 (N_16227,N_11837,N_7561);
nor U16228 (N_16228,N_6624,N_9902);
nand U16229 (N_16229,N_6149,N_11743);
nand U16230 (N_16230,N_10402,N_9505);
nor U16231 (N_16231,N_9533,N_10327);
or U16232 (N_16232,N_9789,N_11647);
and U16233 (N_16233,N_9109,N_11515);
nor U16234 (N_16234,N_8480,N_7523);
nand U16235 (N_16235,N_9717,N_8032);
xor U16236 (N_16236,N_8488,N_6470);
nand U16237 (N_16237,N_10364,N_9498);
nor U16238 (N_16238,N_7869,N_11020);
and U16239 (N_16239,N_10049,N_9962);
and U16240 (N_16240,N_6604,N_11379);
or U16241 (N_16241,N_6452,N_6103);
or U16242 (N_16242,N_7204,N_11146);
nor U16243 (N_16243,N_8113,N_10486);
xnor U16244 (N_16244,N_8735,N_8172);
nor U16245 (N_16245,N_9993,N_6622);
nand U16246 (N_16246,N_9087,N_6184);
xor U16247 (N_16247,N_11190,N_7506);
nand U16248 (N_16248,N_8349,N_11360);
nand U16249 (N_16249,N_6372,N_10997);
or U16250 (N_16250,N_11918,N_6341);
xnor U16251 (N_16251,N_7092,N_11245);
nor U16252 (N_16252,N_6944,N_9838);
xnor U16253 (N_16253,N_6385,N_8279);
or U16254 (N_16254,N_10955,N_10089);
xnor U16255 (N_16255,N_11919,N_9585);
nor U16256 (N_16256,N_6310,N_7120);
nand U16257 (N_16257,N_6728,N_11722);
nor U16258 (N_16258,N_9652,N_7702);
or U16259 (N_16259,N_10480,N_7009);
and U16260 (N_16260,N_10804,N_6076);
nand U16261 (N_16261,N_8790,N_6146);
or U16262 (N_16262,N_7087,N_7595);
nor U16263 (N_16263,N_8046,N_6517);
and U16264 (N_16264,N_9086,N_8307);
xnor U16265 (N_16265,N_6236,N_6101);
or U16266 (N_16266,N_8283,N_10936);
xnor U16267 (N_16267,N_11678,N_6921);
or U16268 (N_16268,N_6035,N_7885);
nand U16269 (N_16269,N_7675,N_9128);
xnor U16270 (N_16270,N_7839,N_6613);
nand U16271 (N_16271,N_11620,N_6307);
xnor U16272 (N_16272,N_6336,N_6473);
nor U16273 (N_16273,N_11930,N_9537);
or U16274 (N_16274,N_9875,N_9146);
and U16275 (N_16275,N_7674,N_10383);
nand U16276 (N_16276,N_7812,N_7021);
nand U16277 (N_16277,N_11756,N_11784);
and U16278 (N_16278,N_7579,N_10174);
or U16279 (N_16279,N_10072,N_11999);
nor U16280 (N_16280,N_9287,N_7956);
or U16281 (N_16281,N_8128,N_10687);
xor U16282 (N_16282,N_9714,N_11372);
nand U16283 (N_16283,N_11813,N_7970);
xnor U16284 (N_16284,N_10940,N_8135);
and U16285 (N_16285,N_11605,N_10447);
and U16286 (N_16286,N_7389,N_8967);
nor U16287 (N_16287,N_11301,N_7269);
or U16288 (N_16288,N_10436,N_7502);
and U16289 (N_16289,N_7117,N_11574);
and U16290 (N_16290,N_10472,N_9032);
xor U16291 (N_16291,N_7239,N_7551);
and U16292 (N_16292,N_10861,N_8309);
nand U16293 (N_16293,N_8301,N_9958);
nand U16294 (N_16294,N_10402,N_6567);
or U16295 (N_16295,N_7065,N_6404);
nor U16296 (N_16296,N_8720,N_11178);
xor U16297 (N_16297,N_11807,N_9767);
and U16298 (N_16298,N_10725,N_11995);
or U16299 (N_16299,N_6824,N_6246);
and U16300 (N_16300,N_9079,N_8698);
and U16301 (N_16301,N_11423,N_10430);
or U16302 (N_16302,N_9167,N_6254);
xor U16303 (N_16303,N_11141,N_7726);
nand U16304 (N_16304,N_6126,N_7053);
nand U16305 (N_16305,N_6093,N_8186);
and U16306 (N_16306,N_11043,N_8020);
xor U16307 (N_16307,N_7809,N_6394);
or U16308 (N_16308,N_11567,N_7890);
and U16309 (N_16309,N_8011,N_7935);
or U16310 (N_16310,N_9479,N_7260);
nor U16311 (N_16311,N_9526,N_9605);
nor U16312 (N_16312,N_6105,N_7657);
nand U16313 (N_16313,N_11414,N_6983);
nor U16314 (N_16314,N_9897,N_6547);
or U16315 (N_16315,N_10206,N_9474);
xnor U16316 (N_16316,N_10706,N_11818);
nand U16317 (N_16317,N_6022,N_10762);
nand U16318 (N_16318,N_6469,N_10293);
or U16319 (N_16319,N_6829,N_8662);
xor U16320 (N_16320,N_9209,N_7762);
nand U16321 (N_16321,N_8059,N_11234);
nand U16322 (N_16322,N_7536,N_11495);
xor U16323 (N_16323,N_8070,N_9072);
xnor U16324 (N_16324,N_10382,N_8725);
and U16325 (N_16325,N_10373,N_10751);
xnor U16326 (N_16326,N_8197,N_9953);
nand U16327 (N_16327,N_9773,N_10993);
or U16328 (N_16328,N_7811,N_7612);
nand U16329 (N_16329,N_9663,N_11252);
or U16330 (N_16330,N_9871,N_10523);
and U16331 (N_16331,N_9052,N_11548);
and U16332 (N_16332,N_9204,N_9401);
and U16333 (N_16333,N_11897,N_9391);
nand U16334 (N_16334,N_10030,N_8273);
xor U16335 (N_16335,N_9649,N_11765);
xnor U16336 (N_16336,N_10775,N_9419);
xor U16337 (N_16337,N_7341,N_7935);
nor U16338 (N_16338,N_9285,N_10474);
and U16339 (N_16339,N_8915,N_8939);
xnor U16340 (N_16340,N_10863,N_10004);
nand U16341 (N_16341,N_8781,N_6432);
nor U16342 (N_16342,N_10378,N_7440);
xnor U16343 (N_16343,N_11006,N_8229);
nand U16344 (N_16344,N_11313,N_8109);
xnor U16345 (N_16345,N_10670,N_9617);
nor U16346 (N_16346,N_10782,N_9323);
xor U16347 (N_16347,N_9712,N_6297);
and U16348 (N_16348,N_11446,N_6563);
xor U16349 (N_16349,N_11261,N_9575);
nor U16350 (N_16350,N_9816,N_11541);
nand U16351 (N_16351,N_11006,N_8983);
and U16352 (N_16352,N_7019,N_10659);
xnor U16353 (N_16353,N_10329,N_9051);
nand U16354 (N_16354,N_10088,N_6912);
or U16355 (N_16355,N_6071,N_10755);
or U16356 (N_16356,N_11147,N_10187);
or U16357 (N_16357,N_10863,N_8655);
or U16358 (N_16358,N_7766,N_11547);
or U16359 (N_16359,N_7405,N_11702);
nand U16360 (N_16360,N_11797,N_10260);
or U16361 (N_16361,N_10984,N_7637);
nand U16362 (N_16362,N_8065,N_9718);
and U16363 (N_16363,N_9833,N_10664);
xor U16364 (N_16364,N_10526,N_11606);
nor U16365 (N_16365,N_11014,N_6925);
and U16366 (N_16366,N_10654,N_11191);
nor U16367 (N_16367,N_10145,N_10723);
xor U16368 (N_16368,N_10878,N_7185);
or U16369 (N_16369,N_9182,N_7322);
nor U16370 (N_16370,N_6520,N_9585);
nand U16371 (N_16371,N_9565,N_8626);
or U16372 (N_16372,N_7220,N_11147);
nor U16373 (N_16373,N_11061,N_9784);
and U16374 (N_16374,N_9985,N_10542);
xor U16375 (N_16375,N_10739,N_6576);
xor U16376 (N_16376,N_6154,N_6341);
nor U16377 (N_16377,N_8675,N_10894);
xnor U16378 (N_16378,N_11775,N_7903);
nor U16379 (N_16379,N_7994,N_11893);
and U16380 (N_16380,N_9990,N_8184);
and U16381 (N_16381,N_10063,N_7464);
xor U16382 (N_16382,N_11384,N_10386);
xor U16383 (N_16383,N_10586,N_8705);
or U16384 (N_16384,N_9922,N_10804);
nor U16385 (N_16385,N_7085,N_7271);
nor U16386 (N_16386,N_7073,N_9542);
and U16387 (N_16387,N_6776,N_6655);
and U16388 (N_16388,N_7669,N_9482);
xor U16389 (N_16389,N_8077,N_7673);
and U16390 (N_16390,N_11531,N_9773);
and U16391 (N_16391,N_6517,N_11429);
nand U16392 (N_16392,N_6466,N_10504);
xor U16393 (N_16393,N_8348,N_11263);
or U16394 (N_16394,N_10040,N_7088);
xnor U16395 (N_16395,N_10960,N_9553);
and U16396 (N_16396,N_8411,N_6444);
nand U16397 (N_16397,N_6577,N_7116);
and U16398 (N_16398,N_7837,N_8043);
and U16399 (N_16399,N_10213,N_8814);
and U16400 (N_16400,N_9309,N_6915);
or U16401 (N_16401,N_10401,N_9499);
xor U16402 (N_16402,N_11201,N_8262);
nand U16403 (N_16403,N_10885,N_10456);
xor U16404 (N_16404,N_9021,N_7363);
nor U16405 (N_16405,N_10474,N_6603);
nand U16406 (N_16406,N_6662,N_9564);
nor U16407 (N_16407,N_8812,N_7644);
or U16408 (N_16408,N_8833,N_11399);
and U16409 (N_16409,N_7087,N_11872);
or U16410 (N_16410,N_8504,N_10853);
or U16411 (N_16411,N_10538,N_10040);
xnor U16412 (N_16412,N_8327,N_7307);
nand U16413 (N_16413,N_10442,N_10139);
nor U16414 (N_16414,N_11665,N_11754);
nand U16415 (N_16415,N_10553,N_11669);
xnor U16416 (N_16416,N_6352,N_10347);
nand U16417 (N_16417,N_7156,N_7793);
nand U16418 (N_16418,N_8265,N_11355);
or U16419 (N_16419,N_8854,N_6662);
and U16420 (N_16420,N_8398,N_8534);
nor U16421 (N_16421,N_6047,N_8611);
nand U16422 (N_16422,N_7490,N_8337);
nand U16423 (N_16423,N_10169,N_9311);
nand U16424 (N_16424,N_8282,N_7232);
and U16425 (N_16425,N_10008,N_8602);
or U16426 (N_16426,N_8909,N_9100);
or U16427 (N_16427,N_10097,N_6927);
nor U16428 (N_16428,N_9969,N_10858);
nor U16429 (N_16429,N_8062,N_10167);
nor U16430 (N_16430,N_10388,N_7004);
and U16431 (N_16431,N_9522,N_11944);
nand U16432 (N_16432,N_8672,N_11599);
nand U16433 (N_16433,N_11896,N_7855);
and U16434 (N_16434,N_9619,N_7515);
xor U16435 (N_16435,N_11314,N_7107);
nand U16436 (N_16436,N_7540,N_7115);
xor U16437 (N_16437,N_7275,N_6291);
nor U16438 (N_16438,N_9111,N_10582);
or U16439 (N_16439,N_9979,N_9636);
and U16440 (N_16440,N_10875,N_10025);
xor U16441 (N_16441,N_9909,N_9767);
nand U16442 (N_16442,N_9061,N_11035);
nor U16443 (N_16443,N_7783,N_6392);
xor U16444 (N_16444,N_9698,N_10948);
and U16445 (N_16445,N_6799,N_7035);
and U16446 (N_16446,N_7953,N_6176);
xor U16447 (N_16447,N_11436,N_9087);
nor U16448 (N_16448,N_10583,N_8853);
nor U16449 (N_16449,N_11297,N_6933);
or U16450 (N_16450,N_7619,N_7365);
xor U16451 (N_16451,N_8404,N_11015);
or U16452 (N_16452,N_8594,N_8527);
and U16453 (N_16453,N_9868,N_11005);
nand U16454 (N_16454,N_11351,N_11955);
and U16455 (N_16455,N_9881,N_7392);
xor U16456 (N_16456,N_6818,N_10694);
and U16457 (N_16457,N_8791,N_9176);
nand U16458 (N_16458,N_8071,N_6439);
nand U16459 (N_16459,N_6741,N_6797);
and U16460 (N_16460,N_11497,N_11803);
xor U16461 (N_16461,N_11176,N_9885);
nor U16462 (N_16462,N_8632,N_10113);
nor U16463 (N_16463,N_11919,N_8694);
and U16464 (N_16464,N_10760,N_9598);
xor U16465 (N_16465,N_11624,N_10737);
nor U16466 (N_16466,N_9542,N_11190);
nor U16467 (N_16467,N_10378,N_10285);
nand U16468 (N_16468,N_6127,N_10922);
and U16469 (N_16469,N_7165,N_11937);
nor U16470 (N_16470,N_8379,N_9446);
xnor U16471 (N_16471,N_8684,N_10146);
xor U16472 (N_16472,N_11667,N_7508);
nand U16473 (N_16473,N_8703,N_9044);
and U16474 (N_16474,N_7468,N_9200);
and U16475 (N_16475,N_9764,N_7630);
and U16476 (N_16476,N_7875,N_7289);
nor U16477 (N_16477,N_7980,N_10490);
and U16478 (N_16478,N_8877,N_9747);
xor U16479 (N_16479,N_9020,N_11399);
and U16480 (N_16480,N_9987,N_10146);
nand U16481 (N_16481,N_7338,N_9141);
or U16482 (N_16482,N_11917,N_6427);
and U16483 (N_16483,N_10009,N_7692);
and U16484 (N_16484,N_8795,N_11482);
nand U16485 (N_16485,N_8269,N_7139);
or U16486 (N_16486,N_6742,N_8902);
xnor U16487 (N_16487,N_7475,N_11547);
nand U16488 (N_16488,N_10623,N_8530);
and U16489 (N_16489,N_9718,N_6942);
and U16490 (N_16490,N_10192,N_7692);
and U16491 (N_16491,N_8882,N_9224);
or U16492 (N_16492,N_11815,N_7427);
and U16493 (N_16493,N_9346,N_9143);
xor U16494 (N_16494,N_8682,N_9609);
and U16495 (N_16495,N_6917,N_8632);
or U16496 (N_16496,N_6891,N_8252);
nor U16497 (N_16497,N_7529,N_11080);
nand U16498 (N_16498,N_7918,N_9401);
or U16499 (N_16499,N_10614,N_8690);
nand U16500 (N_16500,N_9861,N_6721);
nand U16501 (N_16501,N_8764,N_6773);
and U16502 (N_16502,N_9110,N_6528);
or U16503 (N_16503,N_11826,N_6451);
nand U16504 (N_16504,N_6593,N_8236);
nor U16505 (N_16505,N_11280,N_8115);
nand U16506 (N_16506,N_8931,N_7708);
or U16507 (N_16507,N_8949,N_8602);
xor U16508 (N_16508,N_10097,N_7510);
xnor U16509 (N_16509,N_6520,N_8911);
nand U16510 (N_16510,N_11136,N_11251);
and U16511 (N_16511,N_11755,N_9602);
or U16512 (N_16512,N_9647,N_7927);
xor U16513 (N_16513,N_6450,N_8139);
nor U16514 (N_16514,N_11344,N_6975);
nor U16515 (N_16515,N_11670,N_10369);
and U16516 (N_16516,N_7110,N_6328);
and U16517 (N_16517,N_10530,N_9160);
and U16518 (N_16518,N_11263,N_7348);
xnor U16519 (N_16519,N_6871,N_9776);
xor U16520 (N_16520,N_7384,N_6478);
nor U16521 (N_16521,N_6443,N_6920);
nor U16522 (N_16522,N_8752,N_6400);
xor U16523 (N_16523,N_7406,N_6947);
nand U16524 (N_16524,N_7795,N_6292);
nand U16525 (N_16525,N_11506,N_8443);
or U16526 (N_16526,N_11798,N_6469);
nor U16527 (N_16527,N_7055,N_7474);
xnor U16528 (N_16528,N_8322,N_8106);
xnor U16529 (N_16529,N_8149,N_6072);
nor U16530 (N_16530,N_9157,N_7514);
xnor U16531 (N_16531,N_10570,N_10154);
nor U16532 (N_16532,N_9806,N_8708);
and U16533 (N_16533,N_6124,N_11641);
nand U16534 (N_16534,N_9552,N_6551);
and U16535 (N_16535,N_8550,N_8311);
nor U16536 (N_16536,N_8884,N_8487);
or U16537 (N_16537,N_9985,N_9540);
or U16538 (N_16538,N_8806,N_7849);
nand U16539 (N_16539,N_10740,N_9183);
or U16540 (N_16540,N_7227,N_8535);
or U16541 (N_16541,N_6463,N_6699);
xnor U16542 (N_16542,N_10733,N_6245);
xnor U16543 (N_16543,N_11597,N_10632);
nor U16544 (N_16544,N_6379,N_9220);
and U16545 (N_16545,N_11366,N_11625);
nor U16546 (N_16546,N_7328,N_8738);
nand U16547 (N_16547,N_9301,N_7546);
xor U16548 (N_16548,N_6858,N_6196);
nor U16549 (N_16549,N_10834,N_7905);
nor U16550 (N_16550,N_11588,N_7038);
nor U16551 (N_16551,N_10574,N_8274);
nor U16552 (N_16552,N_10824,N_6196);
or U16553 (N_16553,N_11528,N_11793);
and U16554 (N_16554,N_7538,N_11153);
or U16555 (N_16555,N_6725,N_10918);
nand U16556 (N_16556,N_9627,N_11501);
nor U16557 (N_16557,N_6772,N_9893);
xor U16558 (N_16558,N_7771,N_9389);
and U16559 (N_16559,N_6307,N_7840);
or U16560 (N_16560,N_7278,N_9858);
nand U16561 (N_16561,N_8443,N_7647);
and U16562 (N_16562,N_11955,N_6084);
nand U16563 (N_16563,N_10361,N_9348);
and U16564 (N_16564,N_11711,N_10575);
and U16565 (N_16565,N_7698,N_9634);
and U16566 (N_16566,N_8486,N_7935);
and U16567 (N_16567,N_7563,N_7513);
nand U16568 (N_16568,N_11433,N_11667);
nand U16569 (N_16569,N_9175,N_8507);
nand U16570 (N_16570,N_6696,N_10325);
nand U16571 (N_16571,N_8820,N_7196);
nor U16572 (N_16572,N_11883,N_7603);
and U16573 (N_16573,N_6906,N_10476);
nand U16574 (N_16574,N_8525,N_6422);
nor U16575 (N_16575,N_6741,N_11593);
nand U16576 (N_16576,N_10768,N_9572);
or U16577 (N_16577,N_10159,N_6992);
nor U16578 (N_16578,N_7236,N_11384);
nand U16579 (N_16579,N_9902,N_11893);
nand U16580 (N_16580,N_8948,N_6568);
nor U16581 (N_16581,N_10723,N_10878);
and U16582 (N_16582,N_10533,N_10151);
nand U16583 (N_16583,N_7512,N_7551);
nor U16584 (N_16584,N_10679,N_11345);
nand U16585 (N_16585,N_8639,N_9974);
and U16586 (N_16586,N_11365,N_8272);
and U16587 (N_16587,N_7566,N_8490);
or U16588 (N_16588,N_10960,N_8681);
or U16589 (N_16589,N_6810,N_10494);
and U16590 (N_16590,N_8819,N_10644);
and U16591 (N_16591,N_6959,N_7017);
nor U16592 (N_16592,N_6603,N_6012);
nor U16593 (N_16593,N_6971,N_9582);
xor U16594 (N_16594,N_7883,N_6504);
nor U16595 (N_16595,N_8745,N_9958);
xnor U16596 (N_16596,N_7718,N_9970);
nand U16597 (N_16597,N_7607,N_7133);
nand U16598 (N_16598,N_11536,N_9559);
and U16599 (N_16599,N_9376,N_10857);
nand U16600 (N_16600,N_8410,N_11938);
nor U16601 (N_16601,N_9581,N_6580);
and U16602 (N_16602,N_11040,N_9904);
nor U16603 (N_16603,N_9484,N_10263);
and U16604 (N_16604,N_8779,N_7508);
nor U16605 (N_16605,N_11982,N_6182);
xor U16606 (N_16606,N_9622,N_9940);
or U16607 (N_16607,N_8576,N_11969);
nand U16608 (N_16608,N_7043,N_8589);
xor U16609 (N_16609,N_11683,N_7790);
or U16610 (N_16610,N_7721,N_11271);
or U16611 (N_16611,N_8454,N_10120);
xor U16612 (N_16612,N_9919,N_9696);
xor U16613 (N_16613,N_7557,N_7099);
nand U16614 (N_16614,N_6805,N_9148);
and U16615 (N_16615,N_11776,N_7293);
nand U16616 (N_16616,N_7596,N_8391);
xnor U16617 (N_16617,N_11716,N_10012);
and U16618 (N_16618,N_10042,N_10261);
nor U16619 (N_16619,N_10664,N_9882);
and U16620 (N_16620,N_11812,N_10024);
nand U16621 (N_16621,N_10520,N_8873);
or U16622 (N_16622,N_8815,N_10192);
or U16623 (N_16623,N_8085,N_7922);
or U16624 (N_16624,N_7863,N_9094);
nor U16625 (N_16625,N_6210,N_6614);
xor U16626 (N_16626,N_7950,N_7743);
nor U16627 (N_16627,N_7278,N_7753);
nor U16628 (N_16628,N_9005,N_11276);
nand U16629 (N_16629,N_9584,N_9567);
and U16630 (N_16630,N_8829,N_6693);
or U16631 (N_16631,N_10858,N_6511);
xor U16632 (N_16632,N_7016,N_11270);
and U16633 (N_16633,N_6215,N_10121);
xnor U16634 (N_16634,N_6428,N_7232);
or U16635 (N_16635,N_6723,N_11369);
nand U16636 (N_16636,N_8124,N_8224);
nor U16637 (N_16637,N_6466,N_9004);
nand U16638 (N_16638,N_6941,N_6823);
xor U16639 (N_16639,N_6388,N_7463);
xnor U16640 (N_16640,N_9843,N_7893);
and U16641 (N_16641,N_11889,N_8360);
nor U16642 (N_16642,N_9949,N_11964);
and U16643 (N_16643,N_7369,N_10842);
nor U16644 (N_16644,N_9592,N_10145);
or U16645 (N_16645,N_8125,N_8635);
nand U16646 (N_16646,N_8650,N_11611);
xnor U16647 (N_16647,N_11682,N_6044);
xnor U16648 (N_16648,N_8324,N_7730);
or U16649 (N_16649,N_9186,N_9054);
nor U16650 (N_16650,N_11817,N_6975);
xor U16651 (N_16651,N_9448,N_9889);
nand U16652 (N_16652,N_7488,N_11026);
nor U16653 (N_16653,N_6393,N_10220);
xnor U16654 (N_16654,N_7633,N_7194);
nor U16655 (N_16655,N_9817,N_11461);
nand U16656 (N_16656,N_8266,N_11599);
nor U16657 (N_16657,N_8506,N_9831);
nand U16658 (N_16658,N_7566,N_6397);
nor U16659 (N_16659,N_6210,N_9678);
xnor U16660 (N_16660,N_7249,N_7246);
xnor U16661 (N_16661,N_6252,N_9026);
nand U16662 (N_16662,N_8007,N_9291);
nand U16663 (N_16663,N_10781,N_7769);
or U16664 (N_16664,N_9286,N_8611);
nand U16665 (N_16665,N_6817,N_9878);
or U16666 (N_16666,N_8861,N_7587);
and U16667 (N_16667,N_10987,N_9528);
xor U16668 (N_16668,N_8521,N_10146);
xor U16669 (N_16669,N_6771,N_7347);
xor U16670 (N_16670,N_8791,N_6262);
and U16671 (N_16671,N_11128,N_9512);
and U16672 (N_16672,N_11174,N_7995);
and U16673 (N_16673,N_7843,N_7160);
and U16674 (N_16674,N_7701,N_11577);
and U16675 (N_16675,N_8181,N_7781);
nand U16676 (N_16676,N_9672,N_7893);
and U16677 (N_16677,N_11542,N_6981);
or U16678 (N_16678,N_11825,N_11860);
nand U16679 (N_16679,N_9995,N_8338);
or U16680 (N_16680,N_8814,N_6517);
xnor U16681 (N_16681,N_10012,N_11756);
nand U16682 (N_16682,N_9820,N_10003);
xnor U16683 (N_16683,N_8361,N_11437);
xor U16684 (N_16684,N_10526,N_11598);
nor U16685 (N_16685,N_8174,N_6928);
xor U16686 (N_16686,N_10361,N_9422);
xnor U16687 (N_16687,N_7633,N_11250);
and U16688 (N_16688,N_6079,N_10945);
or U16689 (N_16689,N_6177,N_7528);
and U16690 (N_16690,N_8750,N_10398);
or U16691 (N_16691,N_9830,N_10510);
nand U16692 (N_16692,N_11778,N_9317);
and U16693 (N_16693,N_9380,N_10468);
and U16694 (N_16694,N_6261,N_8656);
xor U16695 (N_16695,N_7032,N_9256);
or U16696 (N_16696,N_10331,N_6433);
and U16697 (N_16697,N_10295,N_8245);
xnor U16698 (N_16698,N_6070,N_11880);
or U16699 (N_16699,N_10966,N_11349);
and U16700 (N_16700,N_8044,N_7834);
nand U16701 (N_16701,N_6436,N_7552);
nand U16702 (N_16702,N_6638,N_10999);
xor U16703 (N_16703,N_11802,N_6285);
nand U16704 (N_16704,N_6708,N_6961);
or U16705 (N_16705,N_7300,N_8004);
and U16706 (N_16706,N_8415,N_10469);
nor U16707 (N_16707,N_11426,N_8348);
and U16708 (N_16708,N_11046,N_7118);
and U16709 (N_16709,N_6879,N_6481);
xnor U16710 (N_16710,N_8296,N_10071);
xor U16711 (N_16711,N_6939,N_6695);
nor U16712 (N_16712,N_7203,N_8989);
and U16713 (N_16713,N_6136,N_6444);
nand U16714 (N_16714,N_8512,N_11575);
or U16715 (N_16715,N_9909,N_10928);
and U16716 (N_16716,N_10334,N_10426);
nor U16717 (N_16717,N_6791,N_8269);
nand U16718 (N_16718,N_9752,N_10294);
xor U16719 (N_16719,N_9531,N_8826);
xor U16720 (N_16720,N_11770,N_8215);
nand U16721 (N_16721,N_11830,N_8536);
nand U16722 (N_16722,N_11556,N_11758);
xnor U16723 (N_16723,N_10609,N_6728);
nand U16724 (N_16724,N_8638,N_9337);
and U16725 (N_16725,N_11509,N_6666);
and U16726 (N_16726,N_10462,N_10907);
xnor U16727 (N_16727,N_11004,N_8168);
nand U16728 (N_16728,N_7399,N_8008);
xnor U16729 (N_16729,N_7653,N_9148);
xor U16730 (N_16730,N_7415,N_8310);
xnor U16731 (N_16731,N_11497,N_9976);
or U16732 (N_16732,N_6551,N_11633);
nor U16733 (N_16733,N_6668,N_9734);
and U16734 (N_16734,N_8935,N_8295);
and U16735 (N_16735,N_9000,N_11597);
nand U16736 (N_16736,N_9204,N_11491);
xnor U16737 (N_16737,N_8331,N_8988);
xor U16738 (N_16738,N_11604,N_9960);
nand U16739 (N_16739,N_9409,N_6873);
or U16740 (N_16740,N_7483,N_11350);
or U16741 (N_16741,N_11942,N_10911);
and U16742 (N_16742,N_7928,N_11395);
xnor U16743 (N_16743,N_11239,N_10602);
xor U16744 (N_16744,N_7563,N_11692);
xor U16745 (N_16745,N_9933,N_9561);
nand U16746 (N_16746,N_11045,N_6799);
nand U16747 (N_16747,N_10005,N_6378);
xor U16748 (N_16748,N_10356,N_7481);
nor U16749 (N_16749,N_10823,N_6592);
nand U16750 (N_16750,N_8863,N_10980);
xor U16751 (N_16751,N_7964,N_7561);
nand U16752 (N_16752,N_7093,N_7148);
or U16753 (N_16753,N_7375,N_7492);
nand U16754 (N_16754,N_10673,N_9372);
xnor U16755 (N_16755,N_6104,N_10988);
and U16756 (N_16756,N_11887,N_8786);
xnor U16757 (N_16757,N_8534,N_11401);
xor U16758 (N_16758,N_9420,N_7390);
nand U16759 (N_16759,N_6699,N_11121);
nand U16760 (N_16760,N_6029,N_7197);
or U16761 (N_16761,N_8275,N_9411);
nor U16762 (N_16762,N_7523,N_9061);
and U16763 (N_16763,N_7678,N_8046);
nor U16764 (N_16764,N_7423,N_6180);
xor U16765 (N_16765,N_8832,N_10039);
xor U16766 (N_16766,N_10239,N_11301);
nor U16767 (N_16767,N_9644,N_7792);
nor U16768 (N_16768,N_11992,N_11095);
xor U16769 (N_16769,N_11665,N_8954);
and U16770 (N_16770,N_11863,N_8530);
and U16771 (N_16771,N_9534,N_11417);
nor U16772 (N_16772,N_7533,N_11789);
nand U16773 (N_16773,N_6569,N_11681);
and U16774 (N_16774,N_7910,N_6318);
and U16775 (N_16775,N_7653,N_6294);
and U16776 (N_16776,N_8537,N_11484);
xor U16777 (N_16777,N_6251,N_10509);
nand U16778 (N_16778,N_8148,N_6451);
and U16779 (N_16779,N_11264,N_7454);
xnor U16780 (N_16780,N_6978,N_8066);
and U16781 (N_16781,N_6430,N_11561);
nand U16782 (N_16782,N_7503,N_9961);
or U16783 (N_16783,N_11010,N_8356);
nor U16784 (N_16784,N_7085,N_10092);
nand U16785 (N_16785,N_7900,N_7514);
or U16786 (N_16786,N_8128,N_7036);
xnor U16787 (N_16787,N_9731,N_8913);
and U16788 (N_16788,N_9125,N_6542);
nor U16789 (N_16789,N_10300,N_6849);
nor U16790 (N_16790,N_9859,N_6783);
xnor U16791 (N_16791,N_7218,N_11001);
nand U16792 (N_16792,N_9800,N_6166);
nor U16793 (N_16793,N_9551,N_9887);
nand U16794 (N_16794,N_9042,N_6379);
nor U16795 (N_16795,N_9112,N_6817);
or U16796 (N_16796,N_10411,N_8576);
nor U16797 (N_16797,N_8388,N_6397);
nand U16798 (N_16798,N_8107,N_6746);
nor U16799 (N_16799,N_8467,N_9347);
and U16800 (N_16800,N_8230,N_10158);
or U16801 (N_16801,N_8209,N_10028);
xor U16802 (N_16802,N_6431,N_10304);
nor U16803 (N_16803,N_10198,N_6455);
and U16804 (N_16804,N_7027,N_6293);
xor U16805 (N_16805,N_11156,N_11977);
or U16806 (N_16806,N_7469,N_10038);
xnor U16807 (N_16807,N_7001,N_7556);
nand U16808 (N_16808,N_11042,N_11901);
and U16809 (N_16809,N_9968,N_10779);
xnor U16810 (N_16810,N_7687,N_6996);
nor U16811 (N_16811,N_6789,N_10777);
nand U16812 (N_16812,N_9098,N_9833);
nor U16813 (N_16813,N_7262,N_10409);
or U16814 (N_16814,N_9388,N_10442);
nor U16815 (N_16815,N_7622,N_9194);
nor U16816 (N_16816,N_6839,N_6598);
xor U16817 (N_16817,N_10979,N_7049);
xnor U16818 (N_16818,N_6212,N_7121);
and U16819 (N_16819,N_10353,N_10943);
nor U16820 (N_16820,N_10757,N_6567);
and U16821 (N_16821,N_6406,N_6679);
xnor U16822 (N_16822,N_10100,N_9142);
nor U16823 (N_16823,N_10721,N_9685);
nor U16824 (N_16824,N_11777,N_9734);
and U16825 (N_16825,N_9516,N_8440);
nand U16826 (N_16826,N_7740,N_8876);
or U16827 (N_16827,N_7146,N_6189);
nor U16828 (N_16828,N_10071,N_6993);
nor U16829 (N_16829,N_11213,N_8000);
or U16830 (N_16830,N_8390,N_9144);
xnor U16831 (N_16831,N_10750,N_8260);
or U16832 (N_16832,N_8815,N_8072);
or U16833 (N_16833,N_11287,N_10319);
xnor U16834 (N_16834,N_7174,N_11172);
nor U16835 (N_16835,N_10641,N_6007);
nor U16836 (N_16836,N_7352,N_7644);
and U16837 (N_16837,N_10991,N_9786);
xor U16838 (N_16838,N_7895,N_7712);
nor U16839 (N_16839,N_9057,N_6629);
or U16840 (N_16840,N_11918,N_9650);
and U16841 (N_16841,N_10523,N_10014);
nor U16842 (N_16842,N_8347,N_9483);
xor U16843 (N_16843,N_9600,N_8579);
or U16844 (N_16844,N_9734,N_11487);
nand U16845 (N_16845,N_11167,N_6180);
xor U16846 (N_16846,N_7224,N_6661);
or U16847 (N_16847,N_10709,N_6712);
or U16848 (N_16848,N_10205,N_8412);
nor U16849 (N_16849,N_6145,N_8272);
or U16850 (N_16850,N_8376,N_11313);
or U16851 (N_16851,N_10653,N_11154);
and U16852 (N_16852,N_6327,N_8788);
xor U16853 (N_16853,N_6044,N_7399);
and U16854 (N_16854,N_6966,N_10709);
xnor U16855 (N_16855,N_8319,N_11338);
or U16856 (N_16856,N_6626,N_8259);
nand U16857 (N_16857,N_10168,N_11611);
nand U16858 (N_16858,N_8602,N_11378);
xor U16859 (N_16859,N_10418,N_7708);
xnor U16860 (N_16860,N_11789,N_11491);
xor U16861 (N_16861,N_10595,N_7702);
nor U16862 (N_16862,N_11626,N_11006);
nor U16863 (N_16863,N_6139,N_9416);
nand U16864 (N_16864,N_10852,N_6769);
nor U16865 (N_16865,N_11309,N_10658);
xor U16866 (N_16866,N_8148,N_8609);
nand U16867 (N_16867,N_8597,N_9356);
nor U16868 (N_16868,N_6195,N_9835);
nor U16869 (N_16869,N_8131,N_10935);
nor U16870 (N_16870,N_11968,N_8338);
or U16871 (N_16871,N_9219,N_6294);
nand U16872 (N_16872,N_11656,N_8044);
xnor U16873 (N_16873,N_10209,N_8071);
or U16874 (N_16874,N_7658,N_6061);
xnor U16875 (N_16875,N_7913,N_11183);
or U16876 (N_16876,N_6997,N_10895);
nor U16877 (N_16877,N_7584,N_7219);
xor U16878 (N_16878,N_6298,N_10226);
or U16879 (N_16879,N_8926,N_10892);
xor U16880 (N_16880,N_9011,N_6810);
nor U16881 (N_16881,N_9917,N_7713);
or U16882 (N_16882,N_11594,N_9796);
or U16883 (N_16883,N_8085,N_10268);
nand U16884 (N_16884,N_6385,N_11008);
xnor U16885 (N_16885,N_9108,N_8261);
nand U16886 (N_16886,N_6775,N_6741);
nor U16887 (N_16887,N_6490,N_11849);
nand U16888 (N_16888,N_11349,N_10812);
nor U16889 (N_16889,N_11581,N_9314);
nor U16890 (N_16890,N_6272,N_11667);
or U16891 (N_16891,N_7034,N_7202);
nor U16892 (N_16892,N_9478,N_9991);
or U16893 (N_16893,N_9014,N_8791);
or U16894 (N_16894,N_10508,N_11952);
or U16895 (N_16895,N_11809,N_7574);
and U16896 (N_16896,N_8342,N_7758);
and U16897 (N_16897,N_7963,N_9571);
and U16898 (N_16898,N_10126,N_9395);
or U16899 (N_16899,N_6287,N_9278);
or U16900 (N_16900,N_9451,N_7853);
nand U16901 (N_16901,N_6198,N_9289);
nor U16902 (N_16902,N_11777,N_6411);
xnor U16903 (N_16903,N_8073,N_6195);
or U16904 (N_16904,N_8603,N_7635);
and U16905 (N_16905,N_11398,N_8354);
or U16906 (N_16906,N_11426,N_10802);
nand U16907 (N_16907,N_11690,N_10528);
xor U16908 (N_16908,N_11875,N_10994);
nand U16909 (N_16909,N_11545,N_8725);
and U16910 (N_16910,N_7135,N_10437);
or U16911 (N_16911,N_10823,N_8399);
nand U16912 (N_16912,N_10242,N_8616);
nor U16913 (N_16913,N_8330,N_7642);
nor U16914 (N_16914,N_10470,N_6907);
xor U16915 (N_16915,N_7269,N_7013);
xor U16916 (N_16916,N_11163,N_8250);
nand U16917 (N_16917,N_7289,N_6782);
nor U16918 (N_16918,N_11613,N_10739);
xnor U16919 (N_16919,N_8897,N_8599);
nand U16920 (N_16920,N_8463,N_8603);
xor U16921 (N_16921,N_10455,N_10310);
or U16922 (N_16922,N_7390,N_7010);
nand U16923 (N_16923,N_11940,N_7887);
and U16924 (N_16924,N_10849,N_8253);
or U16925 (N_16925,N_10217,N_7174);
nor U16926 (N_16926,N_9539,N_7316);
or U16927 (N_16927,N_7461,N_10106);
and U16928 (N_16928,N_6838,N_6254);
nand U16929 (N_16929,N_6922,N_10501);
or U16930 (N_16930,N_7076,N_7987);
nand U16931 (N_16931,N_11376,N_7950);
nand U16932 (N_16932,N_10162,N_10224);
or U16933 (N_16933,N_11617,N_7372);
xor U16934 (N_16934,N_7174,N_6600);
and U16935 (N_16935,N_6959,N_8890);
and U16936 (N_16936,N_8951,N_8870);
nand U16937 (N_16937,N_10223,N_9544);
nand U16938 (N_16938,N_8876,N_10152);
nand U16939 (N_16939,N_8115,N_7292);
nor U16940 (N_16940,N_11818,N_11299);
xnor U16941 (N_16941,N_7949,N_7551);
nand U16942 (N_16942,N_11639,N_10865);
or U16943 (N_16943,N_6691,N_11751);
or U16944 (N_16944,N_10763,N_9884);
or U16945 (N_16945,N_7708,N_8023);
or U16946 (N_16946,N_8738,N_11089);
xor U16947 (N_16947,N_8036,N_11611);
nor U16948 (N_16948,N_11170,N_6452);
nor U16949 (N_16949,N_9419,N_11410);
or U16950 (N_16950,N_11386,N_9697);
or U16951 (N_16951,N_6658,N_7059);
or U16952 (N_16952,N_10994,N_11229);
or U16953 (N_16953,N_7412,N_6100);
and U16954 (N_16954,N_9321,N_10850);
or U16955 (N_16955,N_6224,N_10833);
nand U16956 (N_16956,N_9831,N_9122);
xor U16957 (N_16957,N_7380,N_8868);
nor U16958 (N_16958,N_9130,N_6517);
and U16959 (N_16959,N_8844,N_11403);
or U16960 (N_16960,N_8294,N_7781);
nor U16961 (N_16961,N_7323,N_6815);
nand U16962 (N_16962,N_6765,N_6181);
and U16963 (N_16963,N_10391,N_8568);
or U16964 (N_16964,N_9605,N_11837);
nand U16965 (N_16965,N_9528,N_6258);
xnor U16966 (N_16966,N_9099,N_7628);
nand U16967 (N_16967,N_9907,N_10177);
or U16968 (N_16968,N_9884,N_11197);
or U16969 (N_16969,N_10624,N_7570);
nor U16970 (N_16970,N_10391,N_7515);
nand U16971 (N_16971,N_6597,N_10860);
nor U16972 (N_16972,N_8613,N_10537);
nand U16973 (N_16973,N_8726,N_10801);
nor U16974 (N_16974,N_9707,N_8464);
and U16975 (N_16975,N_8223,N_7456);
xnor U16976 (N_16976,N_9109,N_6185);
and U16977 (N_16977,N_6213,N_10837);
and U16978 (N_16978,N_7702,N_8537);
nor U16979 (N_16979,N_11096,N_9155);
xor U16980 (N_16980,N_9354,N_8771);
or U16981 (N_16981,N_6634,N_9029);
nand U16982 (N_16982,N_11696,N_6417);
nand U16983 (N_16983,N_10661,N_10383);
nor U16984 (N_16984,N_11476,N_6110);
or U16985 (N_16985,N_7184,N_7226);
nor U16986 (N_16986,N_6483,N_10072);
nor U16987 (N_16987,N_6318,N_9159);
nor U16988 (N_16988,N_6772,N_11449);
nor U16989 (N_16989,N_8832,N_7098);
nand U16990 (N_16990,N_8243,N_8713);
xnor U16991 (N_16991,N_8412,N_7014);
or U16992 (N_16992,N_10946,N_10649);
and U16993 (N_16993,N_8552,N_6708);
nor U16994 (N_16994,N_11341,N_9332);
xor U16995 (N_16995,N_8275,N_9303);
or U16996 (N_16996,N_10194,N_8799);
xor U16997 (N_16997,N_10782,N_11642);
xor U16998 (N_16998,N_9359,N_10189);
and U16999 (N_16999,N_7973,N_8006);
or U17000 (N_17000,N_7265,N_9521);
nor U17001 (N_17001,N_8620,N_10435);
nor U17002 (N_17002,N_6906,N_10390);
nand U17003 (N_17003,N_7377,N_10633);
and U17004 (N_17004,N_11334,N_7342);
and U17005 (N_17005,N_9657,N_8587);
nand U17006 (N_17006,N_8723,N_11113);
or U17007 (N_17007,N_8261,N_10981);
and U17008 (N_17008,N_11881,N_6876);
and U17009 (N_17009,N_8271,N_9145);
xor U17010 (N_17010,N_10809,N_8016);
xnor U17011 (N_17011,N_7604,N_6212);
nor U17012 (N_17012,N_6287,N_8974);
xor U17013 (N_17013,N_11029,N_6073);
and U17014 (N_17014,N_11193,N_7444);
and U17015 (N_17015,N_7889,N_7895);
xor U17016 (N_17016,N_11039,N_10182);
or U17017 (N_17017,N_7031,N_10483);
nor U17018 (N_17018,N_9828,N_9887);
xor U17019 (N_17019,N_9141,N_7994);
and U17020 (N_17020,N_9574,N_11596);
xor U17021 (N_17021,N_9478,N_6921);
or U17022 (N_17022,N_9991,N_11285);
and U17023 (N_17023,N_6090,N_8797);
nor U17024 (N_17024,N_7591,N_9114);
and U17025 (N_17025,N_8795,N_11210);
nor U17026 (N_17026,N_11526,N_10738);
and U17027 (N_17027,N_10268,N_8921);
or U17028 (N_17028,N_9827,N_7046);
or U17029 (N_17029,N_10554,N_8897);
xor U17030 (N_17030,N_10426,N_10773);
xnor U17031 (N_17031,N_10374,N_10755);
nand U17032 (N_17032,N_6508,N_11774);
or U17033 (N_17033,N_6611,N_10428);
and U17034 (N_17034,N_10487,N_9825);
and U17035 (N_17035,N_8673,N_10081);
or U17036 (N_17036,N_7115,N_11564);
nand U17037 (N_17037,N_10925,N_8017);
or U17038 (N_17038,N_6446,N_8251);
xnor U17039 (N_17039,N_6344,N_10004);
or U17040 (N_17040,N_7291,N_11150);
nand U17041 (N_17041,N_8594,N_9792);
nand U17042 (N_17042,N_11630,N_8233);
nor U17043 (N_17043,N_8432,N_11201);
or U17044 (N_17044,N_6743,N_10802);
nand U17045 (N_17045,N_8975,N_11386);
or U17046 (N_17046,N_7963,N_11144);
or U17047 (N_17047,N_10031,N_8014);
or U17048 (N_17048,N_9129,N_8771);
nor U17049 (N_17049,N_8723,N_10212);
or U17050 (N_17050,N_9281,N_11685);
and U17051 (N_17051,N_11976,N_7256);
nand U17052 (N_17052,N_6570,N_9315);
nand U17053 (N_17053,N_8455,N_6436);
nand U17054 (N_17054,N_7009,N_6935);
nand U17055 (N_17055,N_11174,N_6161);
or U17056 (N_17056,N_6859,N_11640);
nor U17057 (N_17057,N_8768,N_6489);
nand U17058 (N_17058,N_9913,N_7161);
nor U17059 (N_17059,N_8859,N_11092);
xor U17060 (N_17060,N_11290,N_10823);
or U17061 (N_17061,N_8960,N_10175);
nor U17062 (N_17062,N_10534,N_6621);
nand U17063 (N_17063,N_7175,N_8468);
xor U17064 (N_17064,N_7262,N_10289);
nor U17065 (N_17065,N_11609,N_9074);
nor U17066 (N_17066,N_7940,N_6368);
or U17067 (N_17067,N_6334,N_9473);
and U17068 (N_17068,N_6895,N_6782);
and U17069 (N_17069,N_6569,N_9706);
nor U17070 (N_17070,N_8665,N_7817);
xor U17071 (N_17071,N_10550,N_11834);
xnor U17072 (N_17072,N_9308,N_9365);
and U17073 (N_17073,N_8796,N_11428);
xor U17074 (N_17074,N_8906,N_7442);
nand U17075 (N_17075,N_6911,N_6488);
and U17076 (N_17076,N_8031,N_8835);
or U17077 (N_17077,N_8059,N_9771);
xnor U17078 (N_17078,N_10155,N_8633);
or U17079 (N_17079,N_7592,N_8071);
nand U17080 (N_17080,N_8987,N_11692);
and U17081 (N_17081,N_9512,N_8845);
and U17082 (N_17082,N_9038,N_6581);
nor U17083 (N_17083,N_11323,N_9219);
nor U17084 (N_17084,N_10909,N_8914);
nor U17085 (N_17085,N_10720,N_7439);
nand U17086 (N_17086,N_8043,N_11446);
or U17087 (N_17087,N_7044,N_9258);
and U17088 (N_17088,N_6580,N_10523);
and U17089 (N_17089,N_10110,N_8252);
xnor U17090 (N_17090,N_6305,N_6647);
and U17091 (N_17091,N_9990,N_8416);
and U17092 (N_17092,N_11303,N_7009);
xnor U17093 (N_17093,N_10666,N_10920);
or U17094 (N_17094,N_10004,N_8207);
xor U17095 (N_17095,N_7834,N_11420);
nand U17096 (N_17096,N_8181,N_7923);
xnor U17097 (N_17097,N_7309,N_9526);
nand U17098 (N_17098,N_9569,N_6233);
nor U17099 (N_17099,N_6590,N_8577);
nor U17100 (N_17100,N_10499,N_9421);
nor U17101 (N_17101,N_8679,N_9719);
nand U17102 (N_17102,N_9152,N_11665);
xor U17103 (N_17103,N_9250,N_8783);
or U17104 (N_17104,N_6822,N_11114);
and U17105 (N_17105,N_10135,N_8624);
nor U17106 (N_17106,N_11024,N_8025);
nor U17107 (N_17107,N_10035,N_7095);
xor U17108 (N_17108,N_11078,N_9758);
or U17109 (N_17109,N_10369,N_6617);
and U17110 (N_17110,N_8177,N_6628);
xor U17111 (N_17111,N_6902,N_10977);
and U17112 (N_17112,N_10309,N_6657);
nor U17113 (N_17113,N_9728,N_10647);
and U17114 (N_17114,N_9584,N_6921);
nor U17115 (N_17115,N_7256,N_9897);
or U17116 (N_17116,N_11706,N_9803);
nor U17117 (N_17117,N_9534,N_11531);
or U17118 (N_17118,N_9320,N_9406);
xor U17119 (N_17119,N_11481,N_6353);
nand U17120 (N_17120,N_6758,N_7153);
nor U17121 (N_17121,N_8500,N_8714);
xor U17122 (N_17122,N_6309,N_6156);
xnor U17123 (N_17123,N_8160,N_10088);
xor U17124 (N_17124,N_9592,N_9566);
nor U17125 (N_17125,N_9452,N_7841);
or U17126 (N_17126,N_10644,N_10084);
xor U17127 (N_17127,N_8263,N_8433);
xor U17128 (N_17128,N_9838,N_6429);
nand U17129 (N_17129,N_6582,N_10204);
xor U17130 (N_17130,N_10721,N_9207);
and U17131 (N_17131,N_10271,N_8889);
xor U17132 (N_17132,N_10096,N_10807);
or U17133 (N_17133,N_7483,N_6723);
and U17134 (N_17134,N_8186,N_9449);
or U17135 (N_17135,N_9103,N_6232);
nand U17136 (N_17136,N_10001,N_11270);
nor U17137 (N_17137,N_7290,N_9455);
or U17138 (N_17138,N_6627,N_10567);
nor U17139 (N_17139,N_10212,N_6850);
and U17140 (N_17140,N_8524,N_11885);
and U17141 (N_17141,N_8113,N_9778);
nand U17142 (N_17142,N_6532,N_11538);
nor U17143 (N_17143,N_10212,N_11987);
xnor U17144 (N_17144,N_6116,N_7497);
xor U17145 (N_17145,N_6020,N_9985);
nor U17146 (N_17146,N_11315,N_9957);
nand U17147 (N_17147,N_8521,N_11209);
nand U17148 (N_17148,N_6394,N_8667);
xor U17149 (N_17149,N_10441,N_6605);
nand U17150 (N_17150,N_10525,N_7588);
nor U17151 (N_17151,N_9752,N_7374);
and U17152 (N_17152,N_11657,N_11299);
or U17153 (N_17153,N_11316,N_11321);
xor U17154 (N_17154,N_7372,N_7152);
nand U17155 (N_17155,N_7280,N_10985);
nand U17156 (N_17156,N_11505,N_10939);
nand U17157 (N_17157,N_6268,N_7357);
nand U17158 (N_17158,N_8729,N_9620);
or U17159 (N_17159,N_11622,N_11212);
or U17160 (N_17160,N_11798,N_7610);
and U17161 (N_17161,N_8734,N_8706);
xnor U17162 (N_17162,N_11018,N_10167);
and U17163 (N_17163,N_7552,N_11667);
nor U17164 (N_17164,N_6634,N_6798);
or U17165 (N_17165,N_10992,N_11308);
or U17166 (N_17166,N_9437,N_7600);
xnor U17167 (N_17167,N_8855,N_6078);
xnor U17168 (N_17168,N_8346,N_11211);
nor U17169 (N_17169,N_11610,N_11788);
or U17170 (N_17170,N_10061,N_7499);
nand U17171 (N_17171,N_8036,N_7106);
xor U17172 (N_17172,N_11622,N_7966);
xor U17173 (N_17173,N_10822,N_10219);
xor U17174 (N_17174,N_10898,N_6465);
nor U17175 (N_17175,N_7051,N_10580);
nor U17176 (N_17176,N_8277,N_8012);
and U17177 (N_17177,N_7047,N_8302);
nor U17178 (N_17178,N_11411,N_11188);
xnor U17179 (N_17179,N_10321,N_11341);
and U17180 (N_17180,N_8216,N_9444);
nand U17181 (N_17181,N_10752,N_10862);
or U17182 (N_17182,N_11415,N_8281);
and U17183 (N_17183,N_6886,N_9981);
nor U17184 (N_17184,N_9343,N_11925);
nor U17185 (N_17185,N_10793,N_11275);
or U17186 (N_17186,N_10812,N_8304);
nand U17187 (N_17187,N_11114,N_6743);
xor U17188 (N_17188,N_6769,N_8887);
and U17189 (N_17189,N_8105,N_8113);
xnor U17190 (N_17190,N_8767,N_8834);
or U17191 (N_17191,N_8970,N_11084);
or U17192 (N_17192,N_11787,N_10951);
nor U17193 (N_17193,N_8467,N_7938);
or U17194 (N_17194,N_9603,N_9127);
and U17195 (N_17195,N_10367,N_9797);
xor U17196 (N_17196,N_11713,N_9802);
nor U17197 (N_17197,N_10336,N_10405);
nor U17198 (N_17198,N_11341,N_10032);
or U17199 (N_17199,N_6867,N_11973);
or U17200 (N_17200,N_11085,N_8344);
nor U17201 (N_17201,N_11404,N_9819);
and U17202 (N_17202,N_8953,N_9805);
xor U17203 (N_17203,N_10198,N_8078);
nand U17204 (N_17204,N_10626,N_11815);
xor U17205 (N_17205,N_10803,N_6058);
xnor U17206 (N_17206,N_6697,N_10562);
nand U17207 (N_17207,N_6860,N_9125);
nor U17208 (N_17208,N_8174,N_7398);
nand U17209 (N_17209,N_7500,N_7959);
xor U17210 (N_17210,N_8428,N_7649);
nor U17211 (N_17211,N_9524,N_11707);
nand U17212 (N_17212,N_9504,N_6615);
xor U17213 (N_17213,N_10925,N_8520);
nand U17214 (N_17214,N_6104,N_11885);
nand U17215 (N_17215,N_7207,N_10673);
and U17216 (N_17216,N_11191,N_11151);
nor U17217 (N_17217,N_11318,N_9496);
nor U17218 (N_17218,N_9750,N_8442);
nor U17219 (N_17219,N_8532,N_10183);
nor U17220 (N_17220,N_6806,N_9864);
nor U17221 (N_17221,N_11409,N_11638);
nor U17222 (N_17222,N_11793,N_6314);
xor U17223 (N_17223,N_10002,N_9442);
nor U17224 (N_17224,N_9575,N_9096);
and U17225 (N_17225,N_8353,N_8291);
nand U17226 (N_17226,N_9431,N_6706);
xor U17227 (N_17227,N_9444,N_9113);
and U17228 (N_17228,N_6743,N_10740);
or U17229 (N_17229,N_8512,N_10381);
or U17230 (N_17230,N_8111,N_9869);
and U17231 (N_17231,N_10073,N_8073);
xnor U17232 (N_17232,N_8645,N_9445);
and U17233 (N_17233,N_10740,N_8250);
nor U17234 (N_17234,N_7234,N_6133);
xnor U17235 (N_17235,N_8242,N_7426);
and U17236 (N_17236,N_9268,N_7217);
nor U17237 (N_17237,N_7560,N_10965);
nand U17238 (N_17238,N_11192,N_9607);
or U17239 (N_17239,N_6814,N_8773);
nand U17240 (N_17240,N_9216,N_8922);
or U17241 (N_17241,N_9217,N_6529);
nand U17242 (N_17242,N_6160,N_11185);
nor U17243 (N_17243,N_11128,N_11069);
nor U17244 (N_17244,N_10923,N_6251);
or U17245 (N_17245,N_6129,N_7047);
nand U17246 (N_17246,N_10216,N_9221);
nand U17247 (N_17247,N_7159,N_8214);
and U17248 (N_17248,N_10468,N_10383);
or U17249 (N_17249,N_8690,N_7947);
and U17250 (N_17250,N_8283,N_10968);
nor U17251 (N_17251,N_11581,N_10724);
and U17252 (N_17252,N_7149,N_7477);
nor U17253 (N_17253,N_6864,N_9708);
nand U17254 (N_17254,N_7914,N_8650);
or U17255 (N_17255,N_6004,N_9595);
nand U17256 (N_17256,N_11454,N_6296);
nand U17257 (N_17257,N_7904,N_7091);
nand U17258 (N_17258,N_10453,N_8843);
nor U17259 (N_17259,N_9804,N_11683);
or U17260 (N_17260,N_11376,N_11262);
or U17261 (N_17261,N_9676,N_8814);
nor U17262 (N_17262,N_8934,N_8332);
nor U17263 (N_17263,N_10017,N_6887);
or U17264 (N_17264,N_11296,N_7493);
or U17265 (N_17265,N_8865,N_6350);
nor U17266 (N_17266,N_11085,N_6102);
or U17267 (N_17267,N_8148,N_11907);
and U17268 (N_17268,N_11741,N_8791);
nand U17269 (N_17269,N_8539,N_10114);
xnor U17270 (N_17270,N_8702,N_9234);
or U17271 (N_17271,N_6068,N_7596);
and U17272 (N_17272,N_10231,N_10236);
and U17273 (N_17273,N_8778,N_10973);
xor U17274 (N_17274,N_11543,N_7938);
nor U17275 (N_17275,N_6422,N_6462);
nand U17276 (N_17276,N_11379,N_7276);
or U17277 (N_17277,N_10441,N_7668);
xnor U17278 (N_17278,N_6339,N_8537);
nand U17279 (N_17279,N_10655,N_10918);
xor U17280 (N_17280,N_8740,N_11173);
xnor U17281 (N_17281,N_11667,N_11905);
or U17282 (N_17282,N_9206,N_8227);
and U17283 (N_17283,N_11511,N_7213);
xor U17284 (N_17284,N_7996,N_10991);
or U17285 (N_17285,N_8580,N_7268);
and U17286 (N_17286,N_6729,N_9494);
nand U17287 (N_17287,N_11313,N_8825);
or U17288 (N_17288,N_6297,N_11071);
xnor U17289 (N_17289,N_9941,N_7066);
nor U17290 (N_17290,N_11122,N_11356);
xor U17291 (N_17291,N_7480,N_10240);
nand U17292 (N_17292,N_7340,N_6105);
xor U17293 (N_17293,N_8742,N_7713);
xor U17294 (N_17294,N_8793,N_10820);
nand U17295 (N_17295,N_7453,N_9782);
or U17296 (N_17296,N_9063,N_10373);
nand U17297 (N_17297,N_7709,N_8740);
xnor U17298 (N_17298,N_9693,N_8290);
or U17299 (N_17299,N_11939,N_9254);
or U17300 (N_17300,N_8409,N_6228);
and U17301 (N_17301,N_8503,N_11136);
and U17302 (N_17302,N_10005,N_8517);
xor U17303 (N_17303,N_8403,N_9606);
xor U17304 (N_17304,N_7225,N_10456);
or U17305 (N_17305,N_10408,N_11399);
nand U17306 (N_17306,N_10623,N_11282);
xnor U17307 (N_17307,N_8431,N_8960);
or U17308 (N_17308,N_9843,N_8067);
and U17309 (N_17309,N_9515,N_6986);
xnor U17310 (N_17310,N_11512,N_8083);
nand U17311 (N_17311,N_11993,N_11831);
xnor U17312 (N_17312,N_11153,N_8447);
xor U17313 (N_17313,N_11310,N_6833);
or U17314 (N_17314,N_8252,N_10629);
and U17315 (N_17315,N_9550,N_8626);
nand U17316 (N_17316,N_8278,N_9780);
nand U17317 (N_17317,N_8661,N_8721);
xnor U17318 (N_17318,N_7300,N_7265);
nand U17319 (N_17319,N_11996,N_6977);
xnor U17320 (N_17320,N_11212,N_7347);
and U17321 (N_17321,N_6270,N_7982);
xnor U17322 (N_17322,N_9448,N_8701);
or U17323 (N_17323,N_10917,N_9190);
nand U17324 (N_17324,N_6543,N_8473);
xnor U17325 (N_17325,N_6306,N_8624);
nand U17326 (N_17326,N_10387,N_10231);
nor U17327 (N_17327,N_11413,N_8979);
xor U17328 (N_17328,N_9718,N_6804);
nor U17329 (N_17329,N_10909,N_11252);
or U17330 (N_17330,N_9179,N_9918);
nor U17331 (N_17331,N_7910,N_9909);
and U17332 (N_17332,N_7117,N_11618);
or U17333 (N_17333,N_9582,N_11061);
and U17334 (N_17334,N_11351,N_6100);
or U17335 (N_17335,N_6515,N_6300);
and U17336 (N_17336,N_6627,N_10458);
and U17337 (N_17337,N_6360,N_6473);
or U17338 (N_17338,N_9877,N_6372);
nand U17339 (N_17339,N_9181,N_8301);
or U17340 (N_17340,N_8795,N_6619);
or U17341 (N_17341,N_8624,N_9148);
nand U17342 (N_17342,N_7542,N_9021);
xor U17343 (N_17343,N_11390,N_9000);
nand U17344 (N_17344,N_6009,N_7096);
or U17345 (N_17345,N_10442,N_9119);
and U17346 (N_17346,N_8553,N_11176);
xor U17347 (N_17347,N_11233,N_11479);
xor U17348 (N_17348,N_11331,N_8287);
nand U17349 (N_17349,N_6379,N_10909);
nand U17350 (N_17350,N_6333,N_6143);
and U17351 (N_17351,N_9327,N_9844);
nor U17352 (N_17352,N_10159,N_9280);
nor U17353 (N_17353,N_11923,N_9742);
nor U17354 (N_17354,N_6136,N_8592);
nand U17355 (N_17355,N_9616,N_7782);
nor U17356 (N_17356,N_10494,N_8092);
and U17357 (N_17357,N_9850,N_8909);
xnor U17358 (N_17358,N_11728,N_9119);
nand U17359 (N_17359,N_7178,N_10115);
or U17360 (N_17360,N_11499,N_6462);
or U17361 (N_17361,N_9335,N_6653);
or U17362 (N_17362,N_6322,N_8029);
and U17363 (N_17363,N_9481,N_7455);
nor U17364 (N_17364,N_7435,N_9741);
xor U17365 (N_17365,N_9814,N_11906);
and U17366 (N_17366,N_8775,N_6483);
xor U17367 (N_17367,N_11796,N_6851);
and U17368 (N_17368,N_8468,N_7052);
nor U17369 (N_17369,N_6125,N_10997);
or U17370 (N_17370,N_8082,N_10016);
and U17371 (N_17371,N_7368,N_6079);
or U17372 (N_17372,N_9285,N_11358);
and U17373 (N_17373,N_11471,N_7259);
and U17374 (N_17374,N_10804,N_10581);
nor U17375 (N_17375,N_10324,N_10191);
nand U17376 (N_17376,N_10491,N_11411);
xor U17377 (N_17377,N_11845,N_11846);
nor U17378 (N_17378,N_7913,N_11218);
xnor U17379 (N_17379,N_7274,N_7633);
and U17380 (N_17380,N_8832,N_6856);
nor U17381 (N_17381,N_9765,N_9182);
nand U17382 (N_17382,N_9216,N_8463);
nor U17383 (N_17383,N_7904,N_11128);
nor U17384 (N_17384,N_8674,N_7566);
nand U17385 (N_17385,N_8608,N_7825);
nand U17386 (N_17386,N_8594,N_8112);
xor U17387 (N_17387,N_8604,N_9098);
and U17388 (N_17388,N_9051,N_6213);
nor U17389 (N_17389,N_11577,N_10633);
nand U17390 (N_17390,N_10667,N_10845);
nand U17391 (N_17391,N_8869,N_8139);
nor U17392 (N_17392,N_10824,N_6446);
nor U17393 (N_17393,N_11426,N_7559);
nand U17394 (N_17394,N_9814,N_6009);
xnor U17395 (N_17395,N_6103,N_8841);
nor U17396 (N_17396,N_10760,N_8200);
or U17397 (N_17397,N_10377,N_6830);
and U17398 (N_17398,N_8891,N_9418);
xor U17399 (N_17399,N_8316,N_10696);
nor U17400 (N_17400,N_8653,N_6248);
xor U17401 (N_17401,N_10341,N_11511);
and U17402 (N_17402,N_8630,N_7077);
and U17403 (N_17403,N_9747,N_7005);
nand U17404 (N_17404,N_7150,N_11360);
nor U17405 (N_17405,N_11466,N_10497);
xnor U17406 (N_17406,N_10294,N_7189);
nand U17407 (N_17407,N_6322,N_7351);
nand U17408 (N_17408,N_11242,N_11554);
nor U17409 (N_17409,N_11618,N_7755);
nor U17410 (N_17410,N_9029,N_6653);
nor U17411 (N_17411,N_9012,N_6234);
nor U17412 (N_17412,N_9264,N_7487);
or U17413 (N_17413,N_10520,N_9699);
nor U17414 (N_17414,N_8642,N_7962);
or U17415 (N_17415,N_11569,N_6607);
or U17416 (N_17416,N_11727,N_10483);
or U17417 (N_17417,N_9646,N_7916);
xnor U17418 (N_17418,N_9964,N_6757);
xor U17419 (N_17419,N_9307,N_8367);
and U17420 (N_17420,N_7268,N_8701);
or U17421 (N_17421,N_7847,N_8664);
nor U17422 (N_17422,N_10524,N_11475);
nor U17423 (N_17423,N_7943,N_10190);
or U17424 (N_17424,N_8355,N_6524);
and U17425 (N_17425,N_8148,N_7662);
nand U17426 (N_17426,N_10744,N_6609);
nand U17427 (N_17427,N_10972,N_9596);
nor U17428 (N_17428,N_8314,N_7520);
nor U17429 (N_17429,N_8632,N_8490);
nand U17430 (N_17430,N_6981,N_11307);
xor U17431 (N_17431,N_11909,N_9276);
nand U17432 (N_17432,N_9262,N_7762);
or U17433 (N_17433,N_6467,N_11270);
nor U17434 (N_17434,N_7734,N_8005);
xnor U17435 (N_17435,N_10933,N_9544);
nand U17436 (N_17436,N_9318,N_7147);
or U17437 (N_17437,N_10622,N_10959);
and U17438 (N_17438,N_6939,N_11151);
nand U17439 (N_17439,N_11254,N_11658);
or U17440 (N_17440,N_6953,N_11785);
nor U17441 (N_17441,N_8149,N_9978);
xor U17442 (N_17442,N_6637,N_8408);
nand U17443 (N_17443,N_7354,N_10690);
nand U17444 (N_17444,N_7835,N_7651);
or U17445 (N_17445,N_6608,N_10474);
and U17446 (N_17446,N_7580,N_6239);
nand U17447 (N_17447,N_6991,N_8004);
xnor U17448 (N_17448,N_9078,N_8062);
and U17449 (N_17449,N_7496,N_8390);
xor U17450 (N_17450,N_11834,N_8874);
nor U17451 (N_17451,N_6335,N_6445);
nand U17452 (N_17452,N_9842,N_8893);
and U17453 (N_17453,N_8559,N_8940);
xnor U17454 (N_17454,N_7361,N_11279);
nor U17455 (N_17455,N_6524,N_6400);
nand U17456 (N_17456,N_8904,N_11213);
or U17457 (N_17457,N_7459,N_6886);
and U17458 (N_17458,N_6757,N_10750);
and U17459 (N_17459,N_8578,N_9989);
xor U17460 (N_17460,N_7046,N_8757);
nand U17461 (N_17461,N_10058,N_6761);
xnor U17462 (N_17462,N_6394,N_11736);
xnor U17463 (N_17463,N_11807,N_9629);
nand U17464 (N_17464,N_9811,N_9055);
nor U17465 (N_17465,N_11954,N_8016);
xnor U17466 (N_17466,N_6136,N_8366);
nand U17467 (N_17467,N_10408,N_8343);
nand U17468 (N_17468,N_10620,N_8183);
nand U17469 (N_17469,N_11457,N_9425);
and U17470 (N_17470,N_6529,N_6369);
nor U17471 (N_17471,N_7316,N_6408);
nor U17472 (N_17472,N_8773,N_10601);
xnor U17473 (N_17473,N_6683,N_10126);
nor U17474 (N_17474,N_9689,N_8514);
nor U17475 (N_17475,N_6667,N_9655);
xor U17476 (N_17476,N_10016,N_9321);
xnor U17477 (N_17477,N_7977,N_10833);
and U17478 (N_17478,N_11214,N_6086);
nor U17479 (N_17479,N_10628,N_7834);
nor U17480 (N_17480,N_9449,N_8076);
and U17481 (N_17481,N_11423,N_7933);
and U17482 (N_17482,N_8758,N_7162);
nand U17483 (N_17483,N_7643,N_7854);
nor U17484 (N_17484,N_8392,N_7175);
and U17485 (N_17485,N_9409,N_11338);
or U17486 (N_17486,N_8687,N_8002);
nor U17487 (N_17487,N_6350,N_6420);
nor U17488 (N_17488,N_9037,N_11600);
and U17489 (N_17489,N_11438,N_6908);
nor U17490 (N_17490,N_7664,N_9791);
xnor U17491 (N_17491,N_10838,N_9463);
nand U17492 (N_17492,N_6742,N_9652);
and U17493 (N_17493,N_9566,N_10214);
and U17494 (N_17494,N_10431,N_9086);
or U17495 (N_17495,N_7671,N_10699);
nor U17496 (N_17496,N_10643,N_8376);
or U17497 (N_17497,N_10015,N_9246);
and U17498 (N_17498,N_6153,N_11224);
nand U17499 (N_17499,N_9069,N_9306);
or U17500 (N_17500,N_10762,N_8074);
xor U17501 (N_17501,N_10636,N_11357);
xor U17502 (N_17502,N_10084,N_7368);
xor U17503 (N_17503,N_7108,N_10099);
nor U17504 (N_17504,N_7631,N_11440);
nand U17505 (N_17505,N_7321,N_8536);
nand U17506 (N_17506,N_7899,N_7749);
nor U17507 (N_17507,N_10180,N_10898);
nand U17508 (N_17508,N_9287,N_8227);
nor U17509 (N_17509,N_10968,N_6163);
xor U17510 (N_17510,N_11704,N_7812);
nor U17511 (N_17511,N_6320,N_8781);
nand U17512 (N_17512,N_11775,N_10987);
xnor U17513 (N_17513,N_9882,N_7426);
xor U17514 (N_17514,N_9961,N_10059);
nand U17515 (N_17515,N_6848,N_8981);
and U17516 (N_17516,N_6209,N_10580);
nor U17517 (N_17517,N_7693,N_10516);
or U17518 (N_17518,N_7345,N_10743);
xnor U17519 (N_17519,N_8009,N_11918);
or U17520 (N_17520,N_6599,N_7488);
nor U17521 (N_17521,N_10342,N_10925);
nand U17522 (N_17522,N_10768,N_6620);
nor U17523 (N_17523,N_9082,N_9442);
nand U17524 (N_17524,N_8218,N_6791);
xnor U17525 (N_17525,N_9656,N_11742);
and U17526 (N_17526,N_7129,N_6623);
and U17527 (N_17527,N_8291,N_11772);
nor U17528 (N_17528,N_9380,N_10672);
nand U17529 (N_17529,N_10101,N_6861);
nand U17530 (N_17530,N_11070,N_10860);
nand U17531 (N_17531,N_10505,N_9945);
nor U17532 (N_17532,N_8057,N_6874);
xor U17533 (N_17533,N_10268,N_6021);
nor U17534 (N_17534,N_9540,N_6842);
or U17535 (N_17535,N_6201,N_11661);
or U17536 (N_17536,N_7677,N_6497);
nor U17537 (N_17537,N_11381,N_8874);
nand U17538 (N_17538,N_8202,N_6093);
or U17539 (N_17539,N_11233,N_7071);
nor U17540 (N_17540,N_6147,N_10675);
or U17541 (N_17541,N_6076,N_7208);
nor U17542 (N_17542,N_7301,N_9998);
xnor U17543 (N_17543,N_8031,N_11854);
or U17544 (N_17544,N_6038,N_9671);
nor U17545 (N_17545,N_7581,N_9668);
nand U17546 (N_17546,N_10678,N_7857);
or U17547 (N_17547,N_8036,N_8185);
nor U17548 (N_17548,N_8050,N_9988);
xor U17549 (N_17549,N_8653,N_7358);
or U17550 (N_17550,N_8753,N_8935);
and U17551 (N_17551,N_9414,N_9164);
xor U17552 (N_17552,N_9179,N_11299);
or U17553 (N_17553,N_10952,N_6378);
nand U17554 (N_17554,N_6470,N_11466);
nor U17555 (N_17555,N_8453,N_9441);
nor U17556 (N_17556,N_9940,N_9057);
nor U17557 (N_17557,N_7352,N_10647);
and U17558 (N_17558,N_10047,N_8157);
nor U17559 (N_17559,N_10888,N_6169);
nor U17560 (N_17560,N_9700,N_6577);
and U17561 (N_17561,N_11188,N_7469);
or U17562 (N_17562,N_7571,N_6550);
nand U17563 (N_17563,N_6988,N_8095);
xor U17564 (N_17564,N_9219,N_10770);
nor U17565 (N_17565,N_11382,N_6498);
nand U17566 (N_17566,N_7498,N_11766);
xor U17567 (N_17567,N_10922,N_9363);
and U17568 (N_17568,N_11552,N_8126);
or U17569 (N_17569,N_10358,N_9731);
xor U17570 (N_17570,N_6890,N_11577);
nor U17571 (N_17571,N_7030,N_7994);
nor U17572 (N_17572,N_11491,N_6430);
and U17573 (N_17573,N_6325,N_7609);
and U17574 (N_17574,N_8121,N_8612);
or U17575 (N_17575,N_7582,N_8253);
and U17576 (N_17576,N_7829,N_9397);
nor U17577 (N_17577,N_8679,N_8975);
nor U17578 (N_17578,N_11526,N_10369);
nor U17579 (N_17579,N_11749,N_7833);
and U17580 (N_17580,N_6126,N_6461);
xnor U17581 (N_17581,N_7879,N_11024);
or U17582 (N_17582,N_8924,N_10504);
nor U17583 (N_17583,N_10082,N_10227);
nand U17584 (N_17584,N_6972,N_10624);
nand U17585 (N_17585,N_11857,N_10248);
nand U17586 (N_17586,N_9261,N_6237);
xnor U17587 (N_17587,N_7669,N_10478);
xor U17588 (N_17588,N_9315,N_11890);
and U17589 (N_17589,N_10446,N_8348);
nor U17590 (N_17590,N_10918,N_10164);
xnor U17591 (N_17591,N_7404,N_7826);
xnor U17592 (N_17592,N_10534,N_7009);
xnor U17593 (N_17593,N_6218,N_11964);
xor U17594 (N_17594,N_10718,N_8575);
or U17595 (N_17595,N_10350,N_6312);
nor U17596 (N_17596,N_11977,N_6064);
xnor U17597 (N_17597,N_11073,N_9805);
nor U17598 (N_17598,N_11031,N_8091);
and U17599 (N_17599,N_9872,N_9250);
and U17600 (N_17600,N_9608,N_6842);
and U17601 (N_17601,N_8094,N_8564);
xor U17602 (N_17602,N_10552,N_9246);
and U17603 (N_17603,N_7311,N_7654);
xnor U17604 (N_17604,N_10987,N_7815);
xor U17605 (N_17605,N_8164,N_8813);
nand U17606 (N_17606,N_9609,N_10085);
and U17607 (N_17607,N_10460,N_11049);
xor U17608 (N_17608,N_10073,N_8212);
or U17609 (N_17609,N_9850,N_6302);
or U17610 (N_17610,N_7268,N_9271);
nand U17611 (N_17611,N_10203,N_11322);
xor U17612 (N_17612,N_9686,N_6730);
nor U17613 (N_17613,N_8217,N_8078);
nand U17614 (N_17614,N_8070,N_9568);
nor U17615 (N_17615,N_11206,N_7671);
nor U17616 (N_17616,N_10832,N_10933);
and U17617 (N_17617,N_6315,N_7844);
xor U17618 (N_17618,N_7998,N_9153);
xnor U17619 (N_17619,N_8980,N_8081);
or U17620 (N_17620,N_6517,N_6739);
and U17621 (N_17621,N_7437,N_11557);
nor U17622 (N_17622,N_8319,N_11196);
nor U17623 (N_17623,N_9009,N_10637);
nand U17624 (N_17624,N_6982,N_8403);
xor U17625 (N_17625,N_6892,N_11742);
xor U17626 (N_17626,N_10036,N_9365);
nand U17627 (N_17627,N_11252,N_8326);
or U17628 (N_17628,N_11612,N_8259);
and U17629 (N_17629,N_9127,N_11138);
and U17630 (N_17630,N_8882,N_11733);
nand U17631 (N_17631,N_8119,N_6270);
and U17632 (N_17632,N_9868,N_10005);
and U17633 (N_17633,N_9535,N_9586);
nand U17634 (N_17634,N_6316,N_10029);
nand U17635 (N_17635,N_8922,N_11149);
and U17636 (N_17636,N_7271,N_8067);
xnor U17637 (N_17637,N_9774,N_8607);
or U17638 (N_17638,N_7671,N_11065);
xnor U17639 (N_17639,N_7405,N_9270);
and U17640 (N_17640,N_6430,N_10658);
and U17641 (N_17641,N_10589,N_11545);
and U17642 (N_17642,N_10673,N_9994);
nor U17643 (N_17643,N_7834,N_7816);
nand U17644 (N_17644,N_6434,N_6878);
and U17645 (N_17645,N_11471,N_11488);
xnor U17646 (N_17646,N_8133,N_10968);
and U17647 (N_17647,N_11053,N_7576);
xor U17648 (N_17648,N_9150,N_8831);
and U17649 (N_17649,N_7996,N_9868);
and U17650 (N_17650,N_10244,N_6108);
nor U17651 (N_17651,N_8686,N_8712);
xor U17652 (N_17652,N_6710,N_11903);
xnor U17653 (N_17653,N_6516,N_6159);
nand U17654 (N_17654,N_10932,N_9640);
or U17655 (N_17655,N_11258,N_10644);
and U17656 (N_17656,N_10415,N_7824);
xnor U17657 (N_17657,N_10058,N_6570);
nor U17658 (N_17658,N_10145,N_11203);
and U17659 (N_17659,N_7385,N_9510);
or U17660 (N_17660,N_8155,N_11993);
or U17661 (N_17661,N_9856,N_8704);
or U17662 (N_17662,N_9965,N_9816);
or U17663 (N_17663,N_7877,N_6179);
or U17664 (N_17664,N_10137,N_6866);
nor U17665 (N_17665,N_8908,N_10100);
xnor U17666 (N_17666,N_11616,N_11938);
nor U17667 (N_17667,N_6620,N_7919);
nand U17668 (N_17668,N_6442,N_7736);
nor U17669 (N_17669,N_6992,N_6784);
nand U17670 (N_17670,N_8567,N_7182);
or U17671 (N_17671,N_7705,N_10960);
or U17672 (N_17672,N_7049,N_6435);
and U17673 (N_17673,N_11490,N_10683);
or U17674 (N_17674,N_8146,N_6533);
nand U17675 (N_17675,N_9163,N_11629);
xnor U17676 (N_17676,N_7235,N_7422);
nand U17677 (N_17677,N_9717,N_7826);
or U17678 (N_17678,N_6229,N_8464);
and U17679 (N_17679,N_8529,N_11366);
nor U17680 (N_17680,N_10303,N_11223);
or U17681 (N_17681,N_8790,N_11668);
or U17682 (N_17682,N_6589,N_6822);
nor U17683 (N_17683,N_9218,N_6783);
and U17684 (N_17684,N_10656,N_11317);
and U17685 (N_17685,N_8367,N_8396);
nand U17686 (N_17686,N_10843,N_11393);
and U17687 (N_17687,N_11714,N_10124);
nand U17688 (N_17688,N_6913,N_11948);
xor U17689 (N_17689,N_9335,N_8899);
nand U17690 (N_17690,N_11277,N_8194);
nor U17691 (N_17691,N_11763,N_7724);
nand U17692 (N_17692,N_11494,N_10902);
or U17693 (N_17693,N_8223,N_9997);
nor U17694 (N_17694,N_6451,N_10764);
nor U17695 (N_17695,N_10441,N_11374);
or U17696 (N_17696,N_10137,N_9453);
xnor U17697 (N_17697,N_8250,N_10926);
nand U17698 (N_17698,N_7446,N_9722);
xor U17699 (N_17699,N_11286,N_6426);
or U17700 (N_17700,N_11570,N_9436);
nor U17701 (N_17701,N_7865,N_9971);
or U17702 (N_17702,N_7099,N_11656);
xor U17703 (N_17703,N_6192,N_6758);
xnor U17704 (N_17704,N_10412,N_11476);
or U17705 (N_17705,N_11325,N_7077);
and U17706 (N_17706,N_9826,N_8562);
or U17707 (N_17707,N_10285,N_8878);
nor U17708 (N_17708,N_8610,N_10299);
or U17709 (N_17709,N_9961,N_6990);
nor U17710 (N_17710,N_8174,N_8673);
nor U17711 (N_17711,N_9285,N_7242);
nand U17712 (N_17712,N_11199,N_6469);
or U17713 (N_17713,N_9102,N_10142);
or U17714 (N_17714,N_11005,N_8122);
nor U17715 (N_17715,N_9159,N_11832);
nor U17716 (N_17716,N_11792,N_8088);
or U17717 (N_17717,N_7098,N_9596);
nand U17718 (N_17718,N_11942,N_7753);
and U17719 (N_17719,N_9921,N_8489);
and U17720 (N_17720,N_7011,N_7141);
or U17721 (N_17721,N_6580,N_7364);
or U17722 (N_17722,N_10551,N_10394);
xnor U17723 (N_17723,N_11636,N_10708);
or U17724 (N_17724,N_10915,N_10094);
xor U17725 (N_17725,N_6445,N_9420);
or U17726 (N_17726,N_7012,N_11131);
nand U17727 (N_17727,N_8604,N_9970);
nor U17728 (N_17728,N_7421,N_6569);
xor U17729 (N_17729,N_11448,N_7659);
nand U17730 (N_17730,N_9255,N_7804);
and U17731 (N_17731,N_6012,N_9470);
or U17732 (N_17732,N_7770,N_6355);
xnor U17733 (N_17733,N_6057,N_11782);
or U17734 (N_17734,N_9641,N_9850);
nor U17735 (N_17735,N_8130,N_11631);
and U17736 (N_17736,N_9312,N_11131);
or U17737 (N_17737,N_11166,N_6243);
xnor U17738 (N_17738,N_6149,N_9432);
nor U17739 (N_17739,N_11886,N_11050);
xnor U17740 (N_17740,N_9100,N_7804);
nor U17741 (N_17741,N_6319,N_11398);
or U17742 (N_17742,N_11505,N_9451);
and U17743 (N_17743,N_8690,N_10585);
and U17744 (N_17744,N_11423,N_7818);
xor U17745 (N_17745,N_8352,N_11144);
nor U17746 (N_17746,N_7144,N_10560);
nor U17747 (N_17747,N_6151,N_10205);
nand U17748 (N_17748,N_11028,N_6167);
nor U17749 (N_17749,N_9516,N_8911);
and U17750 (N_17750,N_11929,N_11173);
xor U17751 (N_17751,N_7756,N_7248);
nand U17752 (N_17752,N_6696,N_7967);
xnor U17753 (N_17753,N_10634,N_7947);
nor U17754 (N_17754,N_6193,N_8648);
and U17755 (N_17755,N_10008,N_7003);
and U17756 (N_17756,N_9821,N_11115);
and U17757 (N_17757,N_9381,N_11385);
nor U17758 (N_17758,N_10767,N_6377);
nor U17759 (N_17759,N_10663,N_8956);
and U17760 (N_17760,N_10767,N_9644);
xor U17761 (N_17761,N_7749,N_6057);
or U17762 (N_17762,N_11967,N_10998);
xnor U17763 (N_17763,N_6760,N_11583);
or U17764 (N_17764,N_11671,N_8233);
nor U17765 (N_17765,N_10753,N_11403);
or U17766 (N_17766,N_10686,N_11147);
and U17767 (N_17767,N_7898,N_10479);
nand U17768 (N_17768,N_7166,N_8928);
nand U17769 (N_17769,N_9892,N_8510);
nand U17770 (N_17770,N_10031,N_7974);
nand U17771 (N_17771,N_7138,N_10925);
or U17772 (N_17772,N_9987,N_7941);
or U17773 (N_17773,N_6128,N_9855);
or U17774 (N_17774,N_9636,N_6654);
nor U17775 (N_17775,N_10603,N_8735);
or U17776 (N_17776,N_10552,N_9723);
nor U17777 (N_17777,N_8708,N_7611);
nand U17778 (N_17778,N_9578,N_9689);
or U17779 (N_17779,N_10708,N_6303);
and U17780 (N_17780,N_9941,N_6562);
nor U17781 (N_17781,N_10403,N_8786);
xor U17782 (N_17782,N_7458,N_11066);
and U17783 (N_17783,N_10894,N_7320);
or U17784 (N_17784,N_6996,N_7191);
xor U17785 (N_17785,N_7255,N_6938);
or U17786 (N_17786,N_10470,N_8035);
nand U17787 (N_17787,N_7520,N_10261);
nor U17788 (N_17788,N_9329,N_6432);
or U17789 (N_17789,N_8701,N_11244);
and U17790 (N_17790,N_9307,N_11002);
nand U17791 (N_17791,N_9366,N_8298);
xor U17792 (N_17792,N_11599,N_8007);
xnor U17793 (N_17793,N_8436,N_8629);
nor U17794 (N_17794,N_11623,N_6231);
nand U17795 (N_17795,N_10412,N_9089);
xnor U17796 (N_17796,N_6443,N_10863);
nor U17797 (N_17797,N_7393,N_11427);
nand U17798 (N_17798,N_9694,N_6628);
nor U17799 (N_17799,N_9046,N_10271);
or U17800 (N_17800,N_9119,N_7703);
and U17801 (N_17801,N_7883,N_8523);
or U17802 (N_17802,N_11493,N_10764);
and U17803 (N_17803,N_9445,N_8514);
nand U17804 (N_17804,N_11742,N_6374);
and U17805 (N_17805,N_6860,N_9255);
xnor U17806 (N_17806,N_9582,N_9824);
and U17807 (N_17807,N_10780,N_9126);
xor U17808 (N_17808,N_6003,N_6144);
nand U17809 (N_17809,N_10463,N_10731);
or U17810 (N_17810,N_7168,N_9531);
nand U17811 (N_17811,N_9380,N_8309);
or U17812 (N_17812,N_11202,N_10408);
xor U17813 (N_17813,N_7356,N_9092);
nor U17814 (N_17814,N_9915,N_8635);
nand U17815 (N_17815,N_6223,N_7277);
or U17816 (N_17816,N_8429,N_11020);
xnor U17817 (N_17817,N_9818,N_10082);
xnor U17818 (N_17818,N_8032,N_9333);
xnor U17819 (N_17819,N_10405,N_10632);
and U17820 (N_17820,N_8134,N_8044);
or U17821 (N_17821,N_6292,N_6755);
nand U17822 (N_17822,N_10554,N_7215);
nand U17823 (N_17823,N_11638,N_11501);
or U17824 (N_17824,N_6919,N_6951);
nor U17825 (N_17825,N_8226,N_8147);
nand U17826 (N_17826,N_11020,N_9826);
nand U17827 (N_17827,N_8934,N_6405);
nand U17828 (N_17828,N_7995,N_6965);
and U17829 (N_17829,N_9572,N_9633);
or U17830 (N_17830,N_6097,N_11088);
nor U17831 (N_17831,N_8766,N_6851);
nand U17832 (N_17832,N_6400,N_11243);
or U17833 (N_17833,N_11274,N_6628);
xor U17834 (N_17834,N_9220,N_9775);
or U17835 (N_17835,N_11544,N_10052);
nand U17836 (N_17836,N_9686,N_9045);
and U17837 (N_17837,N_11985,N_9873);
nor U17838 (N_17838,N_7586,N_7850);
or U17839 (N_17839,N_7379,N_9483);
nor U17840 (N_17840,N_10477,N_9625);
and U17841 (N_17841,N_6917,N_9836);
nor U17842 (N_17842,N_8616,N_6017);
or U17843 (N_17843,N_7300,N_11401);
xor U17844 (N_17844,N_6479,N_9442);
or U17845 (N_17845,N_10561,N_6229);
or U17846 (N_17846,N_8140,N_11415);
or U17847 (N_17847,N_6705,N_6664);
nor U17848 (N_17848,N_6080,N_10835);
nand U17849 (N_17849,N_9251,N_7668);
or U17850 (N_17850,N_8018,N_8758);
nor U17851 (N_17851,N_8539,N_11228);
or U17852 (N_17852,N_10288,N_9133);
nand U17853 (N_17853,N_6321,N_11636);
nor U17854 (N_17854,N_7389,N_9715);
nor U17855 (N_17855,N_9608,N_8519);
or U17856 (N_17856,N_11737,N_10355);
nand U17857 (N_17857,N_10154,N_9236);
nand U17858 (N_17858,N_7237,N_6159);
nor U17859 (N_17859,N_11248,N_10043);
nor U17860 (N_17860,N_11696,N_11280);
xnor U17861 (N_17861,N_6568,N_7529);
nand U17862 (N_17862,N_11089,N_6228);
or U17863 (N_17863,N_6310,N_9286);
xor U17864 (N_17864,N_11566,N_9190);
xor U17865 (N_17865,N_11670,N_9164);
and U17866 (N_17866,N_10271,N_6349);
nor U17867 (N_17867,N_9550,N_10338);
nand U17868 (N_17868,N_11571,N_6779);
and U17869 (N_17869,N_11645,N_6959);
xnor U17870 (N_17870,N_6561,N_6127);
nor U17871 (N_17871,N_11239,N_8381);
xnor U17872 (N_17872,N_11523,N_8089);
and U17873 (N_17873,N_9867,N_6287);
and U17874 (N_17874,N_9505,N_10460);
nand U17875 (N_17875,N_9851,N_9465);
xnor U17876 (N_17876,N_10228,N_11240);
and U17877 (N_17877,N_10142,N_6591);
or U17878 (N_17878,N_9917,N_8087);
or U17879 (N_17879,N_7338,N_11248);
nand U17880 (N_17880,N_10306,N_11709);
xor U17881 (N_17881,N_8751,N_6642);
nor U17882 (N_17882,N_11334,N_11631);
and U17883 (N_17883,N_11949,N_8842);
nor U17884 (N_17884,N_10310,N_6638);
or U17885 (N_17885,N_11518,N_10801);
xnor U17886 (N_17886,N_10847,N_8650);
nor U17887 (N_17887,N_6943,N_9412);
nor U17888 (N_17888,N_7459,N_8160);
or U17889 (N_17889,N_6783,N_7946);
or U17890 (N_17890,N_8178,N_7277);
or U17891 (N_17891,N_11774,N_8001);
nor U17892 (N_17892,N_8174,N_6816);
or U17893 (N_17893,N_10304,N_9342);
nand U17894 (N_17894,N_6317,N_7436);
nor U17895 (N_17895,N_10738,N_8050);
or U17896 (N_17896,N_9235,N_10187);
or U17897 (N_17897,N_6477,N_9369);
nor U17898 (N_17898,N_8264,N_9706);
and U17899 (N_17899,N_8415,N_11719);
and U17900 (N_17900,N_6506,N_7992);
and U17901 (N_17901,N_7570,N_7094);
or U17902 (N_17902,N_6675,N_7819);
and U17903 (N_17903,N_10514,N_6451);
and U17904 (N_17904,N_6574,N_9764);
nor U17905 (N_17905,N_8677,N_6193);
nor U17906 (N_17906,N_10766,N_9147);
xor U17907 (N_17907,N_10411,N_6646);
or U17908 (N_17908,N_6527,N_7246);
nor U17909 (N_17909,N_11805,N_8818);
and U17910 (N_17910,N_7199,N_6635);
xnor U17911 (N_17911,N_11858,N_11779);
and U17912 (N_17912,N_9517,N_7195);
or U17913 (N_17913,N_8167,N_9619);
xnor U17914 (N_17914,N_7884,N_11204);
nor U17915 (N_17915,N_9160,N_8330);
or U17916 (N_17916,N_11133,N_9073);
nor U17917 (N_17917,N_9986,N_6963);
nand U17918 (N_17918,N_11803,N_8923);
xnor U17919 (N_17919,N_6928,N_9538);
xnor U17920 (N_17920,N_8780,N_7161);
xnor U17921 (N_17921,N_11441,N_8974);
nor U17922 (N_17922,N_10715,N_9615);
and U17923 (N_17923,N_9654,N_6349);
nor U17924 (N_17924,N_6877,N_10941);
or U17925 (N_17925,N_11388,N_7195);
nor U17926 (N_17926,N_6728,N_8100);
or U17927 (N_17927,N_10120,N_7002);
nor U17928 (N_17928,N_8988,N_10427);
or U17929 (N_17929,N_11387,N_6038);
and U17930 (N_17930,N_6429,N_9169);
or U17931 (N_17931,N_10891,N_7357);
xnor U17932 (N_17932,N_8690,N_6495);
nor U17933 (N_17933,N_11833,N_10790);
and U17934 (N_17934,N_8514,N_6615);
nand U17935 (N_17935,N_7538,N_8819);
nor U17936 (N_17936,N_8391,N_8940);
nand U17937 (N_17937,N_8404,N_9663);
and U17938 (N_17938,N_9067,N_7085);
and U17939 (N_17939,N_11716,N_8548);
xnor U17940 (N_17940,N_9805,N_9318);
nand U17941 (N_17941,N_10137,N_9845);
nand U17942 (N_17942,N_9406,N_10426);
and U17943 (N_17943,N_10259,N_9883);
and U17944 (N_17944,N_9148,N_10006);
or U17945 (N_17945,N_8517,N_9377);
nand U17946 (N_17946,N_7511,N_6991);
nand U17947 (N_17947,N_6417,N_9774);
nand U17948 (N_17948,N_6669,N_11178);
nor U17949 (N_17949,N_10611,N_6238);
nor U17950 (N_17950,N_9104,N_8160);
and U17951 (N_17951,N_11763,N_6237);
or U17952 (N_17952,N_8867,N_10567);
nor U17953 (N_17953,N_9293,N_11458);
and U17954 (N_17954,N_10232,N_7021);
or U17955 (N_17955,N_8921,N_8422);
nor U17956 (N_17956,N_8837,N_9595);
nor U17957 (N_17957,N_11414,N_10505);
or U17958 (N_17958,N_10457,N_11951);
nand U17959 (N_17959,N_10773,N_8521);
or U17960 (N_17960,N_8186,N_7031);
xor U17961 (N_17961,N_10855,N_9738);
or U17962 (N_17962,N_7402,N_7954);
xor U17963 (N_17963,N_10432,N_11837);
nand U17964 (N_17964,N_11115,N_9675);
and U17965 (N_17965,N_6705,N_9404);
or U17966 (N_17966,N_8915,N_7717);
or U17967 (N_17967,N_6075,N_11303);
nand U17968 (N_17968,N_6700,N_6931);
xor U17969 (N_17969,N_7584,N_9772);
nor U17970 (N_17970,N_8798,N_6407);
nor U17971 (N_17971,N_9213,N_6279);
or U17972 (N_17972,N_10549,N_7298);
xnor U17973 (N_17973,N_11856,N_10261);
nand U17974 (N_17974,N_8912,N_7590);
nor U17975 (N_17975,N_6964,N_6750);
or U17976 (N_17976,N_7250,N_10023);
nand U17977 (N_17977,N_8950,N_9487);
xnor U17978 (N_17978,N_9900,N_7257);
xnor U17979 (N_17979,N_11346,N_9060);
or U17980 (N_17980,N_9160,N_6513);
nor U17981 (N_17981,N_11024,N_11741);
or U17982 (N_17982,N_8242,N_10353);
nand U17983 (N_17983,N_11229,N_6716);
nand U17984 (N_17984,N_8300,N_11307);
xnor U17985 (N_17985,N_10002,N_9073);
xnor U17986 (N_17986,N_8145,N_10659);
xor U17987 (N_17987,N_10125,N_6093);
or U17988 (N_17988,N_9863,N_8939);
xnor U17989 (N_17989,N_6982,N_7136);
xor U17990 (N_17990,N_10454,N_11003);
nand U17991 (N_17991,N_9790,N_8272);
and U17992 (N_17992,N_8574,N_6490);
and U17993 (N_17993,N_8959,N_7772);
xnor U17994 (N_17994,N_10518,N_11172);
and U17995 (N_17995,N_10039,N_7141);
or U17996 (N_17996,N_6113,N_10303);
xnor U17997 (N_17997,N_6135,N_6551);
nand U17998 (N_17998,N_9109,N_10020);
and U17999 (N_17999,N_6409,N_6718);
or U18000 (N_18000,N_14640,N_13698);
or U18001 (N_18001,N_13560,N_14930);
xor U18002 (N_18002,N_16591,N_12846);
nand U18003 (N_18003,N_15394,N_13623);
xor U18004 (N_18004,N_14012,N_15479);
and U18005 (N_18005,N_16727,N_12312);
or U18006 (N_18006,N_12109,N_14550);
and U18007 (N_18007,N_16376,N_12696);
and U18008 (N_18008,N_15119,N_13512);
or U18009 (N_18009,N_17622,N_12406);
or U18010 (N_18010,N_16031,N_16078);
or U18011 (N_18011,N_12530,N_13946);
xor U18012 (N_18012,N_12172,N_15336);
xor U18013 (N_18013,N_13876,N_17774);
nor U18014 (N_18014,N_17023,N_15967);
nor U18015 (N_18015,N_14295,N_14228);
or U18016 (N_18016,N_16751,N_17334);
and U18017 (N_18017,N_16250,N_15720);
or U18018 (N_18018,N_12650,N_17255);
xor U18019 (N_18019,N_16420,N_17997);
and U18020 (N_18020,N_16425,N_17800);
nor U18021 (N_18021,N_17271,N_14394);
nand U18022 (N_18022,N_16045,N_13828);
or U18023 (N_18023,N_17596,N_13167);
and U18024 (N_18024,N_17985,N_14419);
and U18025 (N_18025,N_13227,N_17559);
nor U18026 (N_18026,N_13031,N_12408);
or U18027 (N_18027,N_15292,N_13399);
xor U18028 (N_18028,N_15484,N_17682);
and U18029 (N_18029,N_15994,N_13354);
nor U18030 (N_18030,N_12361,N_15126);
xor U18031 (N_18031,N_14893,N_16408);
nand U18032 (N_18032,N_13845,N_14351);
or U18033 (N_18033,N_15669,N_15014);
nand U18034 (N_18034,N_17427,N_12049);
nor U18035 (N_18035,N_14598,N_17109);
nand U18036 (N_18036,N_15900,N_16547);
or U18037 (N_18037,N_13786,N_15189);
xnor U18038 (N_18038,N_13100,N_15745);
nor U18039 (N_18039,N_13886,N_16556);
nor U18040 (N_18040,N_12558,N_14060);
xnor U18041 (N_18041,N_17553,N_13517);
or U18042 (N_18042,N_15478,N_13674);
nor U18043 (N_18043,N_14954,N_13937);
nand U18044 (N_18044,N_13120,N_15671);
and U18045 (N_18045,N_15579,N_14609);
and U18046 (N_18046,N_12646,N_17328);
nand U18047 (N_18047,N_17524,N_13864);
or U18048 (N_18048,N_15784,N_13222);
and U18049 (N_18049,N_17148,N_16961);
nand U18050 (N_18050,N_13065,N_17108);
and U18051 (N_18051,N_14159,N_13596);
or U18052 (N_18052,N_15053,N_12034);
or U18053 (N_18053,N_13478,N_12201);
and U18054 (N_18054,N_12750,N_16357);
nor U18055 (N_18055,N_13720,N_13440);
nor U18056 (N_18056,N_17058,N_12197);
or U18057 (N_18057,N_16388,N_15064);
and U18058 (N_18058,N_16351,N_16415);
xnor U18059 (N_18059,N_15698,N_16356);
nand U18060 (N_18060,N_12166,N_15420);
nand U18061 (N_18061,N_12340,N_13418);
xnor U18062 (N_18062,N_14076,N_12680);
xor U18063 (N_18063,N_12392,N_15772);
and U18064 (N_18064,N_15695,N_13826);
nand U18065 (N_18065,N_17024,N_15067);
nor U18066 (N_18066,N_16043,N_16720);
nand U18067 (N_18067,N_12501,N_14339);
or U18068 (N_18068,N_16283,N_13693);
and U18069 (N_18069,N_13882,N_17638);
xor U18070 (N_18070,N_17820,N_12565);
xnor U18071 (N_18071,N_16678,N_14164);
nor U18072 (N_18072,N_14755,N_15454);
nand U18073 (N_18073,N_17726,N_12857);
and U18074 (N_18074,N_15604,N_16249);
and U18075 (N_18075,N_14660,N_13525);
and U18076 (N_18076,N_14858,N_13490);
and U18077 (N_18077,N_17277,N_17176);
nor U18078 (N_18078,N_17137,N_13842);
nor U18079 (N_18079,N_17920,N_12967);
and U18080 (N_18080,N_16321,N_14008);
and U18081 (N_18081,N_16381,N_16701);
nor U18082 (N_18082,N_14585,N_12099);
nor U18083 (N_18083,N_13138,N_12313);
and U18084 (N_18084,N_15356,N_14980);
nor U18085 (N_18085,N_14089,N_15260);
nand U18086 (N_18086,N_15875,N_15502);
xor U18087 (N_18087,N_13562,N_15208);
or U18088 (N_18088,N_13157,N_17078);
nand U18089 (N_18089,N_17215,N_16465);
or U18090 (N_18090,N_12947,N_12956);
or U18091 (N_18091,N_15930,N_17057);
xnor U18092 (N_18092,N_16979,N_13898);
nand U18093 (N_18093,N_12207,N_12798);
and U18094 (N_18094,N_13821,N_15061);
and U18095 (N_18095,N_13630,N_14125);
or U18096 (N_18096,N_13203,N_13284);
or U18097 (N_18097,N_12998,N_17380);
nor U18098 (N_18098,N_14627,N_14850);
or U18099 (N_18099,N_16307,N_14939);
or U18100 (N_18100,N_17847,N_16478);
nor U18101 (N_18101,N_15021,N_17092);
xnor U18102 (N_18102,N_17205,N_14170);
nand U18103 (N_18103,N_14617,N_14018);
nor U18104 (N_18104,N_16118,N_17438);
nand U18105 (N_18105,N_15599,N_13285);
nand U18106 (N_18106,N_15643,N_15752);
nor U18107 (N_18107,N_13906,N_16772);
and U18108 (N_18108,N_15924,N_17956);
and U18109 (N_18109,N_17305,N_15607);
and U18110 (N_18110,N_12054,N_14263);
nand U18111 (N_18111,N_17494,N_17294);
xor U18112 (N_18112,N_16875,N_17100);
or U18113 (N_18113,N_17029,N_17744);
or U18114 (N_18114,N_13761,N_12215);
xnor U18115 (N_18115,N_16059,N_16286);
xor U18116 (N_18116,N_12676,N_16771);
nand U18117 (N_18117,N_14487,N_16521);
and U18118 (N_18118,N_15595,N_15330);
or U18119 (N_18119,N_17165,N_16574);
xnor U18120 (N_18120,N_16306,N_13461);
nor U18121 (N_18121,N_14815,N_12435);
nand U18122 (N_18122,N_16567,N_15042);
xnor U18123 (N_18123,N_15613,N_13738);
or U18124 (N_18124,N_14092,N_17031);
xnor U18125 (N_18125,N_14162,N_12569);
or U18126 (N_18126,N_13335,N_12059);
nand U18127 (N_18127,N_13978,N_14541);
nand U18128 (N_18128,N_13178,N_16021);
or U18129 (N_18129,N_14239,N_17374);
nand U18130 (N_18130,N_16393,N_13330);
and U18131 (N_18131,N_13088,N_14686);
xor U18132 (N_18132,N_14182,N_15633);
nor U18133 (N_18133,N_15080,N_17127);
xnor U18134 (N_18134,N_13292,N_14624);
or U18135 (N_18135,N_16717,N_17437);
nor U18136 (N_18136,N_14603,N_13627);
and U18137 (N_18137,N_15906,N_13732);
nand U18138 (N_18138,N_13366,N_13348);
nor U18139 (N_18139,N_12048,N_14253);
nand U18140 (N_18140,N_16016,N_14774);
or U18141 (N_18141,N_15419,N_12179);
nand U18142 (N_18142,N_15111,N_17829);
and U18143 (N_18143,N_15960,N_15760);
and U18144 (N_18144,N_17190,N_16217);
or U18145 (N_18145,N_13391,N_14035);
and U18146 (N_18146,N_15827,N_15040);
nor U18147 (N_18147,N_12670,N_15023);
or U18148 (N_18148,N_12892,N_15546);
and U18149 (N_18149,N_13448,N_15674);
nor U18150 (N_18150,N_13777,N_16175);
and U18151 (N_18151,N_17219,N_16134);
xnor U18152 (N_18152,N_16238,N_14479);
nor U18153 (N_18153,N_16819,N_17584);
or U18154 (N_18154,N_14636,N_13244);
and U18155 (N_18155,N_15904,N_13671);
xor U18156 (N_18156,N_14269,N_13874);
and U18157 (N_18157,N_14410,N_13406);
nand U18158 (N_18158,N_12330,N_14115);
xnor U18159 (N_18159,N_17362,N_12071);
xor U18160 (N_18160,N_15059,N_17548);
xor U18161 (N_18161,N_17513,N_14177);
nor U18162 (N_18162,N_15953,N_12092);
xor U18163 (N_18163,N_14973,N_15622);
nor U18164 (N_18164,N_16589,N_14129);
and U18165 (N_18165,N_15136,N_15476);
nor U18166 (N_18166,N_17655,N_12479);
nand U18167 (N_18167,N_17320,N_17620);
nand U18168 (N_18168,N_12613,N_13832);
nor U18169 (N_18169,N_17865,N_16966);
nor U18170 (N_18170,N_17636,N_13730);
nor U18171 (N_18171,N_17687,N_16988);
nand U18172 (N_18172,N_17248,N_15085);
xnor U18173 (N_18173,N_12877,N_15615);
nor U18174 (N_18174,N_15097,N_17943);
and U18175 (N_18175,N_14390,N_16504);
nand U18176 (N_18176,N_16329,N_16121);
nand U18177 (N_18177,N_14097,N_17476);
xnor U18178 (N_18178,N_12326,N_13942);
or U18179 (N_18179,N_13545,N_14465);
xor U18180 (N_18180,N_17010,N_17204);
nor U18181 (N_18181,N_13111,N_16784);
or U18182 (N_18182,N_17265,N_13806);
nand U18183 (N_18183,N_15333,N_14155);
and U18184 (N_18184,N_17173,N_13612);
nand U18185 (N_18185,N_13689,N_14167);
nor U18186 (N_18186,N_13997,N_12553);
nand U18187 (N_18187,N_16492,N_13704);
or U18188 (N_18188,N_13305,N_12057);
nand U18189 (N_18189,N_15029,N_12536);
xnor U18190 (N_18190,N_13661,N_12873);
and U18191 (N_18191,N_13588,N_16170);
nand U18192 (N_18192,N_12181,N_16494);
or U18193 (N_18193,N_13282,N_14629);
and U18194 (N_18194,N_15503,N_17583);
nand U18195 (N_18195,N_15340,N_12683);
or U18196 (N_18196,N_12955,N_17144);
nand U18197 (N_18197,N_17314,N_14392);
or U18198 (N_18198,N_16682,N_17626);
nand U18199 (N_18199,N_15367,N_12617);
nand U18200 (N_18200,N_12209,N_13712);
and U18201 (N_18201,N_16490,N_16934);
xnor U18202 (N_18202,N_12285,N_17512);
nand U18203 (N_18203,N_13395,N_12411);
and U18204 (N_18204,N_14433,N_13579);
or U18205 (N_18205,N_12428,N_16167);
nor U18206 (N_18206,N_13012,N_15481);
and U18207 (N_18207,N_15654,N_15285);
or U18208 (N_18208,N_16877,N_16578);
nand U18209 (N_18209,N_13384,N_17135);
xor U18210 (N_18210,N_14538,N_14327);
or U18211 (N_18211,N_17295,N_14929);
nand U18212 (N_18212,N_14564,N_14428);
or U18213 (N_18213,N_14287,N_16073);
nand U18214 (N_18214,N_16011,N_13411);
and U18215 (N_18215,N_16534,N_12451);
or U18216 (N_18216,N_14025,N_13115);
nand U18217 (N_18217,N_13185,N_14854);
and U18218 (N_18218,N_14848,N_15282);
nand U18219 (N_18219,N_14693,N_13850);
xor U18220 (N_18220,N_16263,N_13913);
or U18221 (N_18221,N_17492,N_13270);
or U18222 (N_18222,N_17214,N_15177);
xnor U18223 (N_18223,N_13615,N_17593);
or U18224 (N_18224,N_12318,N_15482);
xor U18225 (N_18225,N_14211,N_15157);
and U18226 (N_18226,N_16199,N_14223);
xnor U18227 (N_18227,N_14168,N_16613);
xnor U18228 (N_18228,N_12114,N_12611);
or U18229 (N_18229,N_15466,N_17142);
xnor U18230 (N_18230,N_17821,N_17832);
and U18231 (N_18231,N_15699,N_13307);
or U18232 (N_18232,N_16565,N_15103);
xnor U18233 (N_18233,N_12818,N_13625);
or U18234 (N_18234,N_16990,N_12102);
or U18235 (N_18235,N_15555,N_12307);
nand U18236 (N_18236,N_15648,N_14944);
nand U18237 (N_18237,N_16790,N_14749);
and U18238 (N_18238,N_12813,N_17973);
xnor U18239 (N_18239,N_16974,N_13094);
or U18240 (N_18240,N_14937,N_16821);
or U18241 (N_18241,N_13553,N_12015);
xor U18242 (N_18242,N_14404,N_17016);
xnor U18243 (N_18243,N_17924,N_17202);
and U18244 (N_18244,N_17530,N_13133);
or U18245 (N_18245,N_17796,N_14837);
nor U18246 (N_18246,N_16582,N_15563);
nor U18247 (N_18247,N_12586,N_14555);
nor U18248 (N_18248,N_15318,N_16846);
or U18249 (N_18249,N_12189,N_16583);
or U18250 (N_18250,N_17318,N_14391);
nand U18251 (N_18251,N_17151,N_16312);
xor U18252 (N_18252,N_14865,N_13408);
nand U18253 (N_18253,N_13509,N_13707);
and U18254 (N_18254,N_15694,N_17431);
nor U18255 (N_18255,N_17471,N_13278);
nor U18256 (N_18256,N_12602,N_15378);
and U18257 (N_18257,N_16100,N_15066);
nand U18258 (N_18258,N_17749,N_12856);
nor U18259 (N_18259,N_13890,N_14007);
or U18260 (N_18260,N_12573,N_15984);
nor U18261 (N_18261,N_16781,N_15594);
or U18262 (N_18262,N_12767,N_16479);
xor U18263 (N_18263,N_17837,N_17845);
or U18264 (N_18264,N_14792,N_12665);
nand U18265 (N_18265,N_13437,N_16538);
or U18266 (N_18266,N_15676,N_15940);
nor U18267 (N_18267,N_17025,N_12694);
and U18268 (N_18268,N_16467,N_12921);
and U18269 (N_18269,N_13021,N_15848);
and U18270 (N_18270,N_14030,N_14374);
nor U18271 (N_18271,N_12011,N_13682);
nand U18272 (N_18272,N_17805,N_17627);
nand U18273 (N_18273,N_16335,N_16262);
or U18274 (N_18274,N_13762,N_13257);
xnor U18275 (N_18275,N_13843,N_13158);
and U18276 (N_18276,N_12023,N_15450);
or U18277 (N_18277,N_17790,N_12702);
or U18278 (N_18278,N_15187,N_13286);
and U18279 (N_18279,N_12876,N_13793);
and U18280 (N_18280,N_14703,N_16115);
nor U18281 (N_18281,N_13804,N_15740);
nor U18282 (N_18282,N_17946,N_12780);
and U18283 (N_18283,N_12283,N_16274);
or U18284 (N_18284,N_12546,N_12792);
nor U18285 (N_18285,N_14868,N_12174);
nor U18286 (N_18286,N_15712,N_16624);
or U18287 (N_18287,N_17383,N_15518);
or U18288 (N_18288,N_14688,N_17140);
or U18289 (N_18289,N_13599,N_12708);
nand U18290 (N_18290,N_15448,N_17143);
nor U18291 (N_18291,N_13811,N_14108);
nor U18292 (N_18292,N_16296,N_14153);
and U18293 (N_18293,N_15000,N_13518);
nor U18294 (N_18294,N_15320,N_15039);
xor U18295 (N_18295,N_14742,N_16850);
or U18296 (N_18296,N_14107,N_13802);
and U18297 (N_18297,N_15362,N_14024);
nand U18298 (N_18298,N_16663,N_17649);
nand U18299 (N_18299,N_12465,N_16174);
xor U18300 (N_18300,N_17098,N_15507);
xor U18301 (N_18301,N_16012,N_13260);
nand U18302 (N_18302,N_13870,N_17218);
or U18303 (N_18303,N_16339,N_14981);
xnor U18304 (N_18304,N_12137,N_12452);
nand U18305 (N_18305,N_17485,N_15554);
nand U18306 (N_18306,N_13197,N_17003);
nor U18307 (N_18307,N_16868,N_15220);
nand U18308 (N_18308,N_12888,N_14475);
nand U18309 (N_18309,N_16019,N_13442);
or U18310 (N_18310,N_12365,N_13912);
xnor U18311 (N_18311,N_13940,N_17657);
and U18312 (N_18312,N_17911,N_13367);
xnor U18313 (N_18313,N_14208,N_16382);
and U18314 (N_18314,N_14446,N_12150);
nor U18315 (N_18315,N_17772,N_12551);
or U18316 (N_18316,N_17838,N_15808);
or U18317 (N_18317,N_14521,N_13232);
or U18318 (N_18318,N_13077,N_13679);
nor U18319 (N_18319,N_16438,N_12934);
xor U18320 (N_18320,N_14161,N_16168);
nand U18321 (N_18321,N_14847,N_14418);
nor U18322 (N_18322,N_13023,N_13556);
xor U18323 (N_18323,N_15128,N_14885);
and U18324 (N_18324,N_12806,N_14867);
nor U18325 (N_18325,N_15880,N_13321);
nor U18326 (N_18326,N_13951,N_17076);
xor U18327 (N_18327,N_14041,N_13034);
xnor U18328 (N_18328,N_17203,N_14569);
nand U18329 (N_18329,N_16499,N_15972);
nor U18330 (N_18330,N_15195,N_13008);
or U18331 (N_18331,N_14065,N_14481);
nand U18332 (N_18332,N_15660,N_15913);
nor U18333 (N_18333,N_12117,N_17562);
nor U18334 (N_18334,N_14591,N_17775);
xnor U18335 (N_18335,N_13691,N_17718);
and U18336 (N_18336,N_16914,N_16927);
nor U18337 (N_18337,N_15332,N_17987);
nand U18338 (N_18338,N_13746,N_16700);
xnor U18339 (N_18339,N_12458,N_14921);
nand U18340 (N_18340,N_17952,N_15001);
and U18341 (N_18341,N_14158,N_17711);
and U18342 (N_18342,N_13606,N_17680);
and U18343 (N_18343,N_15713,N_17576);
and U18344 (N_18344,N_17310,N_12072);
or U18345 (N_18345,N_12191,N_14179);
and U18346 (N_18346,N_14554,N_16691);
nor U18347 (N_18347,N_12265,N_17433);
nand U18348 (N_18348,N_13935,N_16667);
nor U18349 (N_18349,N_17830,N_16553);
and U18350 (N_18350,N_17698,N_15603);
nor U18351 (N_18351,N_12468,N_16096);
and U18352 (N_18352,N_16715,N_14903);
xor U18353 (N_18353,N_16967,N_14956);
xnor U18354 (N_18354,N_16977,N_15211);
nand U18355 (N_18355,N_12014,N_13421);
or U18356 (N_18356,N_15504,N_12502);
nand U18357 (N_18357,N_14950,N_13371);
xor U18358 (N_18358,N_13372,N_13540);
xnor U18359 (N_18359,N_13955,N_13767);
or U18360 (N_18360,N_15487,N_16512);
nor U18361 (N_18361,N_17477,N_13680);
and U18362 (N_18362,N_12804,N_12075);
or U18363 (N_18363,N_14307,N_12599);
xnor U18364 (N_18364,N_16234,N_17560);
and U18365 (N_18365,N_15771,N_14063);
nor U18366 (N_18366,N_12902,N_17416);
and U18367 (N_18367,N_13485,N_12887);
and U18368 (N_18368,N_17895,N_13353);
nand U18369 (N_18369,N_14265,N_16284);
nor U18370 (N_18370,N_16281,N_15212);
and U18371 (N_18371,N_15756,N_17856);
nor U18372 (N_18372,N_15982,N_17609);
nand U18373 (N_18373,N_16742,N_13010);
xor U18374 (N_18374,N_12381,N_14005);
nand U18375 (N_18375,N_15846,N_17557);
nor U18376 (N_18376,N_16859,N_16370);
nor U18377 (N_18377,N_12860,N_15765);
xnor U18378 (N_18378,N_17551,N_14246);
nand U18379 (N_18379,N_12649,N_15248);
nand U18380 (N_18380,N_16780,N_13592);
nor U18381 (N_18381,N_13175,N_14335);
or U18382 (N_18382,N_17146,N_13424);
nor U18383 (N_18383,N_15156,N_16147);
xnor U18384 (N_18384,N_17330,N_14117);
nor U18385 (N_18385,N_16664,N_17113);
nand U18386 (N_18386,N_15832,N_13780);
nand U18387 (N_18387,N_15526,N_12672);
xnor U18388 (N_18388,N_15255,N_15072);
nand U18389 (N_18389,N_15662,N_14254);
or U18390 (N_18390,N_13091,N_14764);
nor U18391 (N_18391,N_15922,N_16256);
xor U18392 (N_18392,N_16493,N_14836);
nand U18393 (N_18393,N_16159,N_15191);
xnor U18394 (N_18394,N_12513,N_12834);
nor U18395 (N_18395,N_17942,N_14765);
xor U18396 (N_18396,N_15363,N_17402);
xnor U18397 (N_18397,N_15343,N_14189);
nor U18398 (N_18398,N_17145,N_12699);
xnor U18399 (N_18399,N_17611,N_15531);
or U18400 (N_18400,N_15709,N_14979);
xnor U18401 (N_18401,N_13847,N_17222);
and U18402 (N_18402,N_13871,N_15583);
or U18403 (N_18403,N_17722,N_12076);
or U18404 (N_18404,N_13194,N_13127);
and U18405 (N_18405,N_12450,N_16833);
xnor U18406 (N_18406,N_14985,N_13651);
nand U18407 (N_18407,N_17356,N_14845);
and U18408 (N_18408,N_14841,N_13719);
xnor U18409 (N_18409,N_13998,N_15584);
nand U18410 (N_18410,N_15124,N_13563);
nor U18411 (N_18411,N_13668,N_12367);
nand U18412 (N_18412,N_12751,N_17065);
xor U18413 (N_18413,N_14319,N_16911);
and U18414 (N_18414,N_14578,N_16188);
nor U18415 (N_18415,N_17090,N_15327);
nor U18416 (N_18416,N_16303,N_17914);
or U18417 (N_18417,N_13963,N_14875);
xnor U18418 (N_18418,N_12145,N_15895);
nand U18419 (N_18419,N_16050,N_13574);
or U18420 (N_18420,N_13894,N_15152);
xor U18421 (N_18421,N_16783,N_14236);
nand U18422 (N_18422,N_15426,N_17293);
and U18423 (N_18423,N_17990,N_12871);
xor U18424 (N_18424,N_12488,N_13984);
and U18425 (N_18425,N_15317,N_15371);
or U18426 (N_18426,N_15655,N_14644);
xnor U18427 (N_18427,N_16947,N_15711);
and U18428 (N_18428,N_15125,N_13479);
nor U18429 (N_18429,N_16738,N_15821);
nor U18430 (N_18430,N_15705,N_17502);
nor U18431 (N_18431,N_13609,N_17464);
nand U18432 (N_18432,N_16787,N_15102);
xnor U18433 (N_18433,N_14347,N_13188);
nor U18434 (N_18434,N_12142,N_15130);
xor U18435 (N_18435,N_16861,N_12690);
and U18436 (N_18436,N_16520,N_12969);
nor U18437 (N_18437,N_17554,N_13794);
nor U18438 (N_18438,N_16855,N_14006);
or U18439 (N_18439,N_17770,N_13357);
nor U18440 (N_18440,N_13007,N_17333);
nor U18441 (N_18441,N_12541,N_15743);
nand U18442 (N_18442,N_12907,N_17795);
and U18443 (N_18443,N_13328,N_13944);
nand U18444 (N_18444,N_13900,N_13466);
nor U18445 (N_18445,N_16802,N_13125);
nor U18446 (N_18446,N_14322,N_12080);
xor U18447 (N_18447,N_14403,N_17996);
nor U18448 (N_18448,N_13660,N_17834);
or U18449 (N_18449,N_17189,N_13058);
nor U18450 (N_18450,N_17967,N_13267);
and U18451 (N_18451,N_12854,N_17186);
and U18452 (N_18452,N_14238,N_14360);
nand U18453 (N_18453,N_16056,N_14892);
nor U18454 (N_18454,N_16090,N_16254);
or U18455 (N_18455,N_12688,N_17587);
nand U18456 (N_18456,N_13241,N_12590);
nand U18457 (N_18457,N_17629,N_16754);
nor U18458 (N_18458,N_13672,N_15068);
nand U18459 (N_18459,N_12821,N_12772);
and U18460 (N_18460,N_12130,N_17979);
nand U18461 (N_18461,N_17699,N_16987);
nand U18462 (N_18462,N_17094,N_16758);
and U18463 (N_18463,N_12227,N_15893);
nand U18464 (N_18464,N_14436,N_12753);
nand U18465 (N_18465,N_13758,N_13015);
nor U18466 (N_18466,N_13699,N_14061);
xnor U18467 (N_18467,N_17342,N_12002);
nand U18468 (N_18468,N_14338,N_15473);
or U18469 (N_18469,N_14308,N_15204);
xor U18470 (N_18470,N_13510,N_14028);
and U18471 (N_18471,N_12111,N_12833);
xor U18472 (N_18472,N_15580,N_16311);
xnor U18473 (N_18473,N_15192,N_13867);
xor U18474 (N_18474,N_13796,N_12448);
nand U18475 (N_18475,N_15364,N_15673);
nand U18476 (N_18476,N_17287,N_12837);
nor U18477 (N_18477,N_12814,N_17216);
nand U18478 (N_18478,N_17085,N_16362);
and U18479 (N_18479,N_14626,N_14518);
or U18480 (N_18480,N_12636,N_14361);
nor U18481 (N_18481,N_16554,N_15852);
or U18482 (N_18482,N_15529,N_17961);
nor U18483 (N_18483,N_15155,N_16642);
or U18484 (N_18484,N_17463,N_12006);
nand U18485 (N_18485,N_12924,N_13373);
or U18486 (N_18486,N_15480,N_12441);
nand U18487 (N_18487,N_13716,N_14466);
nor U18488 (N_18488,N_13452,N_16404);
and U18489 (N_18489,N_13962,N_14655);
nor U18490 (N_18490,N_16464,N_17175);
or U18491 (N_18491,N_17958,N_15618);
xor U18492 (N_18492,N_12718,N_15471);
and U18493 (N_18493,N_12198,N_17086);
xor U18494 (N_18494,N_17007,N_13050);
nand U18495 (N_18495,N_12195,N_14922);
nand U18496 (N_18496,N_14400,N_15379);
and U18497 (N_18497,N_14207,N_16455);
and U18498 (N_18498,N_14496,N_12495);
and U18499 (N_18499,N_13848,N_13684);
xor U18500 (N_18500,N_13763,N_12762);
xnor U18501 (N_18501,N_16635,N_13187);
nand U18502 (N_18502,N_13533,N_14318);
nand U18503 (N_18503,N_16940,N_12494);
xor U18504 (N_18504,N_17254,N_13745);
nor U18505 (N_18505,N_12661,N_15091);
xor U18506 (N_18506,N_17909,N_12754);
xor U18507 (N_18507,N_12894,N_12788);
xor U18508 (N_18508,N_17927,N_13255);
nand U18509 (N_18509,N_13096,N_12154);
and U18510 (N_18510,N_17074,N_17678);
and U18511 (N_18511,N_12525,N_17809);
and U18512 (N_18512,N_17051,N_12524);
or U18513 (N_18513,N_16346,N_13742);
xnor U18514 (N_18514,N_15276,N_15810);
xor U18515 (N_18515,N_13457,N_12604);
nor U18516 (N_18516,N_16973,N_12261);
nor U18517 (N_18517,N_16536,N_14553);
nand U18518 (N_18518,N_13280,N_14923);
nor U18519 (N_18519,N_14622,N_17603);
or U18520 (N_18520,N_16571,N_13364);
nor U18521 (N_18521,N_12695,N_17739);
nand U18522 (N_18522,N_15755,N_17659);
xor U18523 (N_18523,N_16178,N_12052);
nor U18524 (N_18524,N_13797,N_16579);
or U18525 (N_18525,N_14454,N_14099);
nor U18526 (N_18526,N_16835,N_12795);
nor U18527 (N_18527,N_15235,N_12404);
xor U18528 (N_18528,N_15751,N_12129);
or U18529 (N_18529,N_15012,N_14671);
xnor U18530 (N_18530,N_15744,N_12592);
xor U18531 (N_18531,N_13580,N_17831);
xnor U18532 (N_18532,N_12564,N_14567);
and U18533 (N_18533,N_17843,N_16689);
and U18534 (N_18534,N_17097,N_12187);
xor U18535 (N_18535,N_16766,N_17632);
or U18536 (N_18536,N_14291,N_15849);
nor U18537 (N_18537,N_13456,N_15890);
nand U18538 (N_18538,N_14781,N_17537);
xor U18539 (N_18539,N_16009,N_13902);
and U18540 (N_18540,N_13272,N_16913);
or U18541 (N_18541,N_12156,N_17241);
nand U18542 (N_18542,N_12230,N_13729);
xnor U18543 (N_18543,N_12440,N_14013);
and U18544 (N_18544,N_17220,N_14494);
xor U18545 (N_18545,N_12042,N_17999);
or U18546 (N_18546,N_13887,N_13250);
nand U18547 (N_18547,N_15207,N_14397);
and U18548 (N_18548,N_15147,N_14513);
nor U18549 (N_18549,N_13905,N_14286);
and U18550 (N_18550,N_15108,N_17634);
or U18551 (N_18551,N_16373,N_13739);
or U18552 (N_18552,N_16709,N_14719);
nor U18553 (N_18553,N_14314,N_13991);
xor U18554 (N_18554,N_17459,N_17177);
or U18555 (N_18555,N_14812,N_17890);
xnor U18556 (N_18556,N_12143,N_17578);
and U18557 (N_18557,N_12044,N_13980);
xnor U18558 (N_18558,N_15035,N_12779);
nand U18559 (N_18559,N_16300,N_15350);
or U18560 (N_18560,N_14673,N_13165);
xor U18561 (N_18561,N_17458,N_16450);
or U18562 (N_18562,N_16825,N_17107);
nand U18563 (N_18563,N_16858,N_17604);
or U18564 (N_18564,N_16153,N_16525);
nand U18565 (N_18565,N_15288,N_14098);
nor U18566 (N_18566,N_17676,N_13202);
nand U18567 (N_18567,N_15884,N_14422);
nand U18568 (N_18568,N_14209,N_16395);
xnor U18569 (N_18569,N_15310,N_14925);
nor U18570 (N_18570,N_13494,N_14299);
or U18571 (N_18571,N_13493,N_15169);
or U18572 (N_18572,N_13646,N_15174);
xnor U18573 (N_18573,N_13514,N_16791);
nand U18574 (N_18574,N_17325,N_13032);
nor U18575 (N_18575,N_15561,N_17719);
or U18576 (N_18576,N_12509,N_14434);
and U18577 (N_18577,N_12697,N_12959);
xnor U18578 (N_18578,N_17251,N_12936);
nor U18579 (N_18579,N_12686,N_15831);
or U18580 (N_18580,N_13378,N_16082);
xor U18581 (N_18581,N_15414,N_14916);
xnor U18582 (N_18582,N_17577,N_13888);
or U18583 (N_18583,N_12855,N_17612);
nand U18584 (N_18584,N_16081,N_15725);
xnor U18585 (N_18585,N_13818,N_14345);
and U18586 (N_18586,N_13976,N_17658);
nand U18587 (N_18587,N_17470,N_15016);
or U18588 (N_18588,N_12413,N_17417);
xor U18589 (N_18589,N_16734,N_16810);
nor U18590 (N_18590,N_13869,N_13289);
xnor U18591 (N_18591,N_16005,N_12355);
nor U18592 (N_18592,N_13474,N_16968);
xnor U18593 (N_18593,N_14819,N_14342);
xnor U18594 (N_18594,N_14429,N_17129);
nand U18595 (N_18595,N_17637,N_13329);
or U18596 (N_18596,N_14232,N_15565);
nor U18597 (N_18597,N_12065,N_16461);
nand U18598 (N_18598,N_16721,N_17316);
or U18599 (N_18599,N_16265,N_17889);
xnor U18600 (N_18600,N_17907,N_14779);
nor U18601 (N_18601,N_14376,N_13619);
nor U18602 (N_18602,N_14300,N_14643);
or U18603 (N_18603,N_13643,N_12040);
or U18604 (N_18604,N_12489,N_14290);
nor U18605 (N_18605,N_14831,N_13859);
or U18606 (N_18606,N_14399,N_14027);
or U18607 (N_18607,N_17787,N_15228);
or U18608 (N_18608,N_13423,N_13341);
nand U18609 (N_18609,N_13337,N_16864);
or U18610 (N_18610,N_15786,N_13141);
xor U18611 (N_18611,N_17880,N_13799);
or U18612 (N_18612,N_13361,N_15860);
xnor U18613 (N_18613,N_17691,N_17257);
nand U18614 (N_18614,N_12983,N_16120);
or U18615 (N_18615,N_15537,N_15256);
nor U18616 (N_18616,N_14011,N_15154);
nand U18617 (N_18617,N_17336,N_16474);
xor U18618 (N_18618,N_15954,N_15724);
nand U18619 (N_18619,N_14407,N_16716);
xor U18620 (N_18620,N_15467,N_14563);
nor U18621 (N_18621,N_15365,N_17963);
and U18622 (N_18622,N_14420,N_15366);
and U18623 (N_18623,N_12865,N_17565);
nor U18624 (N_18624,N_12678,N_16289);
xor U18625 (N_18625,N_14090,N_13727);
nand U18626 (N_18626,N_14709,N_13801);
nor U18627 (N_18627,N_15305,N_16023);
or U18628 (N_18628,N_17601,N_13349);
xnor U18629 (N_18629,N_14252,N_14015);
and U18630 (N_18630,N_12240,N_15238);
xnor U18631 (N_18631,N_17839,N_14692);
or U18632 (N_18632,N_16441,N_13820);
xnor U18633 (N_18633,N_16419,N_17340);
xor U18634 (N_18634,N_16837,N_12485);
nor U18635 (N_18635,N_15098,N_14572);
or U18636 (N_18636,N_12389,N_14458);
nand U18637 (N_18637,N_15115,N_15224);
or U18638 (N_18638,N_16181,N_17894);
nand U18639 (N_18639,N_17976,N_15523);
nand U18640 (N_18640,N_12578,N_16743);
xnor U18641 (N_18641,N_15817,N_17684);
nor U18642 (N_18642,N_17588,N_14156);
and U18643 (N_18643,N_13183,N_12321);
nand U18644 (N_18644,N_12991,N_14844);
or U18645 (N_18645,N_15055,N_14963);
nand U18646 (N_18646,N_15451,N_14143);
and U18647 (N_18647,N_13476,N_17182);
or U18648 (N_18648,N_17027,N_14512);
nand U18649 (N_18649,N_15240,N_14835);
nand U18650 (N_18650,N_15179,N_14310);
xor U18651 (N_18651,N_15289,N_16714);
nor U18652 (N_18652,N_15283,N_14224);
or U18653 (N_18653,N_15800,N_16332);
nor U18654 (N_18654,N_17389,N_13539);
and U18655 (N_18655,N_13340,N_12802);
xnor U18656 (N_18656,N_12825,N_13929);
nor U18657 (N_18657,N_15881,N_12790);
and U18658 (N_18658,N_17993,N_16744);
nand U18659 (N_18659,N_16224,N_15286);
or U18660 (N_18660,N_17918,N_13294);
or U18661 (N_18661,N_12009,N_13046);
nor U18662 (N_18662,N_14717,N_16920);
nor U18663 (N_18663,N_14186,N_13863);
or U18664 (N_18664,N_16029,N_12214);
xor U18665 (N_18665,N_17589,N_12518);
nor U18666 (N_18666,N_12831,N_12184);
and U18667 (N_18667,N_13705,N_12671);
nor U18668 (N_18668,N_13404,N_17931);
or U18669 (N_18669,N_17422,N_12260);
nor U18670 (N_18670,N_14192,N_15767);
or U18671 (N_18671,N_16187,N_17018);
nor U18672 (N_18672,N_14771,N_17447);
nand U18673 (N_18673,N_14105,N_12226);
and U18674 (N_18674,N_16200,N_16301);
or U18675 (N_18675,N_17628,N_16259);
or U18676 (N_18676,N_12133,N_12358);
or U18677 (N_18677,N_15358,N_15623);
or U18678 (N_18678,N_15346,N_15008);
nand U18679 (N_18679,N_14811,N_14796);
or U18680 (N_18680,N_16692,N_17111);
nor U18681 (N_18681,N_17908,N_14745);
and U18682 (N_18682,N_17073,N_16114);
and U18683 (N_18683,N_13465,N_15242);
and U18684 (N_18684,N_16902,N_12897);
nor U18685 (N_18685,N_14009,N_12722);
nand U18686 (N_18686,N_13338,N_13104);
or U18687 (N_18687,N_12108,N_16051);
or U18688 (N_18688,N_14853,N_13189);
xor U18689 (N_18689,N_16818,N_16632);
or U18690 (N_18690,N_17697,N_13313);
nand U18691 (N_18691,N_12012,N_14017);
nor U18692 (N_18692,N_17398,N_14411);
and U18693 (N_18693,N_17666,N_15046);
nor U18694 (N_18694,N_13788,N_12120);
and U18695 (N_18695,N_13965,N_15637);
and U18696 (N_18696,N_14722,N_17338);
nand U18697 (N_18697,N_12374,N_16385);
nor U18698 (N_18698,N_16518,N_16496);
nand U18699 (N_18699,N_15640,N_15413);
and U18700 (N_18700,N_13246,N_17905);
xor U18701 (N_18701,N_14780,N_17102);
nand U18702 (N_18702,N_13392,N_12923);
nand U18703 (N_18703,N_12740,N_13151);
and U18704 (N_18704,N_16577,N_13445);
or U18705 (N_18705,N_15197,N_13491);
xnor U18706 (N_18706,N_16996,N_15566);
and U18707 (N_18707,N_12761,N_15418);
nor U18708 (N_18708,N_17012,N_13939);
or U18709 (N_18709,N_14653,N_16733);
nand U18710 (N_18710,N_17217,N_17779);
nand U18711 (N_18711,N_15412,N_13638);
nor U18712 (N_18712,N_14071,N_15069);
nor U18713 (N_18713,N_17806,N_12679);
nor U18714 (N_18714,N_15178,N_12760);
xnor U18715 (N_18715,N_14714,N_17081);
or U18716 (N_18716,N_15337,N_16360);
xnor U18717 (N_18717,N_15807,N_15748);
or U18718 (N_18718,N_15287,N_17299);
xor U18719 (N_18719,N_13640,N_15051);
xor U18720 (N_18720,N_17555,N_17474);
or U18721 (N_18721,N_15963,N_12832);
nor U18722 (N_18722,N_15959,N_16022);
or U18723 (N_18723,N_12669,N_13492);
xnor U18724 (N_18724,N_14121,N_14368);
and U18725 (N_18725,N_17974,N_15460);
xnor U18726 (N_18726,N_13968,N_12380);
nand U18727 (N_18727,N_15759,N_14150);
and U18728 (N_18728,N_12729,N_17740);
nand U18729 (N_18729,N_17357,N_13812);
nor U18730 (N_18730,N_15243,N_14059);
nand U18731 (N_18731,N_14602,N_12687);
nand U18732 (N_18732,N_16297,N_16466);
nor U18733 (N_18733,N_13024,N_17793);
and U18734 (N_18734,N_12382,N_14529);
nand U18735 (N_18735,N_17759,N_17645);
nand U18736 (N_18736,N_17157,N_13056);
xnor U18737 (N_18737,N_12148,N_15445);
nand U18738 (N_18738,N_14704,N_14927);
xor U18739 (N_18739,N_15057,N_16778);
nor U18740 (N_18740,N_12487,N_17878);
or U18741 (N_18741,N_12940,N_12126);
and U18742 (N_18742,N_14081,N_12375);
nor U18743 (N_18743,N_12852,N_15218);
or U18744 (N_18744,N_15020,N_13792);
or U18745 (N_18745,N_13261,N_16058);
xor U18746 (N_18746,N_14346,N_14851);
and U18747 (N_18747,N_14273,N_13374);
and U18748 (N_18748,N_13854,N_14967);
or U18749 (N_18749,N_12001,N_14309);
and U18750 (N_18750,N_15568,N_15512);
nor U18751 (N_18751,N_12799,N_16398);
and U18752 (N_18752,N_13775,N_16895);
and U18753 (N_18753,N_16434,N_17667);
nand U18754 (N_18754,N_15505,N_16405);
and U18755 (N_18755,N_17172,N_14356);
and U18756 (N_18756,N_12352,N_16854);
nand U18757 (N_18757,N_15635,N_15045);
xor U18758 (N_18758,N_13557,N_12193);
or U18759 (N_18759,N_14902,N_14943);
and U18760 (N_18760,N_15998,N_16278);
and U18761 (N_18761,N_16759,N_16728);
nand U18762 (N_18762,N_15280,N_17866);
and U18763 (N_18763,N_16696,N_16951);
or U18764 (N_18764,N_12845,N_12867);
or U18765 (N_18765,N_12152,N_15321);
or U18766 (N_18766,N_16719,N_16269);
or U18767 (N_18767,N_14301,N_17066);
nand U18768 (N_18768,N_12107,N_16909);
nand U18769 (N_18769,N_13018,N_12535);
and U18770 (N_18770,N_14216,N_13287);
nand U18771 (N_18771,N_16018,N_17317);
nor U18772 (N_18772,N_13172,N_16811);
nand U18773 (N_18773,N_13972,N_14485);
or U18774 (N_18774,N_14510,N_16559);
nand U18775 (N_18775,N_14750,N_16602);
nor U18776 (N_18776,N_17767,N_17858);
nor U18777 (N_18777,N_17377,N_13891);
xnor U18778 (N_18778,N_14801,N_16834);
and U18779 (N_18779,N_14031,N_13325);
or U18780 (N_18780,N_16817,N_13550);
nand U18781 (N_18781,N_16449,N_15862);
nand U18782 (N_18782,N_15736,N_16007);
xor U18783 (N_18783,N_15086,N_16756);
or U18784 (N_18784,N_15475,N_12891);
nor U18785 (N_18785,N_16879,N_15778);
nor U18786 (N_18786,N_13069,N_13230);
nor U18787 (N_18787,N_14570,N_13587);
nor U18788 (N_18788,N_15534,N_17867);
nor U18789 (N_18789,N_12917,N_14234);
nand U18790 (N_18790,N_17538,N_17479);
xor U18791 (N_18791,N_16748,N_15923);
xnor U18792 (N_18792,N_12878,N_16436);
nor U18793 (N_18793,N_17898,N_15681);
nand U18794 (N_18794,N_13528,N_14492);
xnor U18795 (N_18795,N_12973,N_13221);
and U18796 (N_18796,N_15575,N_13385);
nand U18797 (N_18797,N_14408,N_14083);
xnor U18798 (N_18798,N_16594,N_15170);
nor U18799 (N_18799,N_16173,N_15649);
xor U18800 (N_18800,N_15704,N_16564);
nand U18801 (N_18801,N_17225,N_14800);
nor U18802 (N_18802,N_16535,N_12393);
and U18803 (N_18803,N_17826,N_13042);
nor U18804 (N_18804,N_12801,N_14476);
xor U18805 (N_18805,N_14978,N_13928);
xnor U18806 (N_18806,N_14870,N_16661);
nor U18807 (N_18807,N_14452,N_16592);
xor U18808 (N_18808,N_14438,N_12439);
nor U18809 (N_18809,N_13590,N_15747);
and U18810 (N_18810,N_16399,N_17863);
or U18811 (N_18811,N_14472,N_16662);
nor U18812 (N_18812,N_16773,N_15347);
or U18813 (N_18813,N_14661,N_17520);
or U18814 (N_18814,N_14393,N_15768);
nand U18815 (N_18815,N_17529,N_13311);
and U18816 (N_18816,N_13195,N_17117);
xor U18817 (N_18817,N_15270,N_16223);
nand U18818 (N_18818,N_16899,N_15722);
and U18819 (N_18819,N_15840,N_12616);
nand U18820 (N_18820,N_12110,N_13598);
or U18821 (N_18821,N_16292,N_14450);
nor U18822 (N_18822,N_15483,N_12582);
or U18823 (N_18823,N_13081,N_16670);
and U18824 (N_18824,N_14227,N_12388);
or U18825 (N_18825,N_14102,N_12241);
and U18826 (N_18826,N_16057,N_17088);
xnor U18827 (N_18827,N_16085,N_17252);
xor U18828 (N_18828,N_15630,N_14961);
xor U18829 (N_18829,N_17169,N_12083);
and U18830 (N_18830,N_15521,N_15446);
and U18831 (N_18831,N_12293,N_12890);
or U18832 (N_18832,N_15430,N_12274);
nand U18833 (N_18833,N_13150,N_12398);
nor U18834 (N_18834,N_17366,N_14183);
xnor U18835 (N_18835,N_14776,N_13872);
nor U18836 (N_18836,N_13637,N_17991);
nand U18837 (N_18837,N_13584,N_13360);
nor U18838 (N_18838,N_15241,N_14205);
nor U18839 (N_18839,N_12254,N_17307);
and U18840 (N_18840,N_15329,N_16230);
nor U18841 (N_18841,N_16629,N_13487);
nor U18842 (N_18842,N_13659,N_13807);
or U18843 (N_18843,N_12259,N_14244);
nor U18844 (N_18844,N_15833,N_13060);
xor U18845 (N_18845,N_15250,N_14919);
xnor U18846 (N_18846,N_16070,N_17118);
nor U18847 (N_18847,N_17616,N_15397);
or U18848 (N_18848,N_15536,N_17712);
or U18849 (N_18849,N_13486,N_17695);
xor U18850 (N_18850,N_14969,N_12805);
or U18851 (N_18851,N_17037,N_15581);
nor U18852 (N_18852,N_17407,N_13009);
and U18853 (N_18853,N_16067,N_13570);
nor U18854 (N_18854,N_14856,N_17948);
xor U18855 (N_18855,N_17469,N_15406);
xor U18856 (N_18856,N_16586,N_16872);
xnor U18857 (N_18857,N_17761,N_14171);
and U18858 (N_18858,N_16651,N_16731);
nand U18859 (N_18859,N_12419,N_14451);
and U18860 (N_18860,N_15592,N_14064);
nor U18861 (N_18861,N_17408,N_17495);
or U18862 (N_18862,N_15107,N_12467);
xnor U18863 (N_18863,N_14638,N_17516);
nor U18864 (N_18864,N_16261,N_13142);
nor U18865 (N_18865,N_17980,N_16653);
and U18866 (N_18866,N_16129,N_17563);
nand U18867 (N_18867,N_12157,N_14491);
nand U18868 (N_18868,N_15464,N_13884);
nand U18869 (N_18869,N_15530,N_15183);
nor U18870 (N_18870,N_14424,N_14758);
and U18871 (N_18871,N_13837,N_15060);
xor U18872 (N_18872,N_14940,N_12493);
nor U18873 (N_18873,N_16650,N_16617);
nor U18874 (N_18874,N_17276,N_12963);
xor U18875 (N_18875,N_17738,N_14042);
or U18876 (N_18876,N_15639,N_14199);
and U18877 (N_18877,N_13889,N_16686);
nand U18878 (N_18878,N_14784,N_12962);
or U18879 (N_18879,N_12399,N_17701);
xnor U18880 (N_18880,N_12433,N_17835);
or U18881 (N_18881,N_15334,N_13030);
xor U18882 (N_18882,N_15750,N_13409);
xor U18883 (N_18883,N_13650,N_15210);
or U18884 (N_18884,N_16160,N_15409);
nor U18885 (N_18885,N_12540,N_17455);
xnor U18886 (N_18886,N_17008,N_16593);
nand U18887 (N_18887,N_17468,N_14384);
or U18888 (N_18888,N_12035,N_14302);
nor U18889 (N_18889,N_13342,N_15868);
or U18890 (N_18890,N_12990,N_12840);
nor U18891 (N_18891,N_12882,N_15985);
nor U18892 (N_18892,N_17497,N_17694);
nor U18893 (N_18893,N_12239,N_13473);
or U18894 (N_18894,N_16486,N_15795);
nand U18895 (N_18895,N_16161,N_14833);
xor U18896 (N_18896,N_16006,N_17877);
nand U18897 (N_18897,N_12626,N_14039);
nor U18898 (N_18898,N_13992,N_13726);
xor U18899 (N_18899,N_15634,N_13613);
nand U18900 (N_18900,N_12310,N_15938);
nand U18901 (N_18901,N_13441,N_15710);
and U18902 (N_18902,N_12903,N_14545);
and U18903 (N_18903,N_16491,N_16513);
and U18904 (N_18904,N_13607,N_12290);
nor U18905 (N_18905,N_13783,N_16840);
nor U18906 (N_18906,N_16334,N_13973);
nand U18907 (N_18907,N_17541,N_15354);
xnor U18908 (N_18908,N_17746,N_12422);
xnor U18909 (N_18909,N_15411,N_12384);
nand U18910 (N_18910,N_12203,N_13676);
nand U18911 (N_18911,N_13087,N_16392);
xor U18912 (N_18912,N_16368,N_17937);
or U18913 (N_18913,N_15325,N_15281);
nand U18914 (N_18914,N_14639,N_13920);
and U18915 (N_18915,N_12477,N_13401);
or U18916 (N_18916,N_12537,N_16896);
nand U18917 (N_18917,N_12838,N_13415);
and U18918 (N_18918,N_13315,N_16195);
and U18919 (N_18919,N_15970,N_16533);
nand U18920 (N_18920,N_12031,N_13426);
xor U18921 (N_18921,N_15058,N_15421);
xor U18922 (N_18922,N_15685,N_17064);
nor U18923 (N_18923,N_15359,N_13781);
nand U18924 (N_18924,N_17284,N_12010);
or U18925 (N_18925,N_16371,N_17644);
or U18926 (N_18926,N_15692,N_13186);
xnor U18927 (N_18927,N_14303,N_15423);
and U18928 (N_18928,N_12091,N_15261);
or U18929 (N_18929,N_15036,N_15844);
xor U18930 (N_18930,N_13673,N_14710);
xnor U18931 (N_18931,N_13468,N_17812);
xnor U18932 (N_18932,N_16888,N_14305);
nand U18933 (N_18933,N_12715,N_15990);
nand U18934 (N_18934,N_13089,N_13683);
nor U18935 (N_18935,N_14972,N_17624);
or U18936 (N_18936,N_17765,N_16828);
or U18937 (N_18937,N_12655,N_14165);
and U18938 (N_18938,N_17704,N_12577);
or U18939 (N_18939,N_15707,N_13519);
and U18940 (N_18940,N_14798,N_13283);
or U18941 (N_18941,N_13542,N_13082);
or U18942 (N_18942,N_16708,N_13713);
nand U18943 (N_18943,N_15087,N_12591);
xnor U18944 (N_18944,N_12974,N_16505);
xor U18945 (N_18945,N_13760,N_15777);
xnor U18946 (N_18946,N_16137,N_16313);
or U18947 (N_18947,N_17810,N_17180);
nor U18948 (N_18948,N_17410,N_12161);
and U18949 (N_18949,N_16805,N_16202);
nand U18950 (N_18950,N_12327,N_16131);
xor U18951 (N_18951,N_14977,N_12084);
xor U18952 (N_18952,N_17984,N_15864);
and U18953 (N_18953,N_13369,N_14565);
nand U18954 (N_18954,N_16000,N_13678);
and U18955 (N_18955,N_15018,N_13223);
and U18956 (N_18956,N_15733,N_14995);
xor U18957 (N_18957,N_14221,N_14349);
or U18958 (N_18958,N_13201,N_12159);
nor U18959 (N_18959,N_13159,N_16605);
or U18960 (N_18960,N_15686,N_16637);
nor U18961 (N_18961,N_16946,N_16367);
nand U18962 (N_18962,N_14568,N_12607);
xor U18963 (N_18963,N_15780,N_14723);
and U18964 (N_18964,N_12123,N_15749);
nand U18965 (N_18965,N_15578,N_16345);
nand U18966 (N_18966,N_14528,N_16726);
nor U18967 (N_18967,N_15117,N_15009);
nor U18968 (N_18968,N_13904,N_12733);
or U18969 (N_18969,N_14430,N_12069);
xnor U18970 (N_18970,N_16232,N_15296);
and U18971 (N_18971,N_15586,N_17283);
or U18972 (N_18972,N_12869,N_14970);
xor U18973 (N_18973,N_15146,N_14577);
nor U18974 (N_18974,N_17358,N_16075);
nand U18975 (N_18975,N_14700,N_12085);
nand U18976 (N_18976,N_13722,N_16489);
nand U18977 (N_18977,N_13743,N_12797);
nand U18978 (N_18978,N_12763,N_16792);
and U18979 (N_18979,N_13084,N_15376);
or U18980 (N_18980,N_13537,N_17188);
xnor U18981 (N_18981,N_12105,N_16816);
or U18982 (N_18982,N_12884,N_13814);
nand U18983 (N_18983,N_16444,N_16183);
or U18984 (N_18984,N_13521,N_16690);
nand U18985 (N_18985,N_17361,N_17087);
and U18986 (N_18986,N_13822,N_15026);
xor U18987 (N_18987,N_14315,N_15857);
xnor U18988 (N_18988,N_14185,N_17005);
nand U18989 (N_18989,N_17350,N_14600);
and U18990 (N_18990,N_15878,N_16767);
or U18991 (N_18991,N_13621,N_16248);
or U18992 (N_18992,N_15472,N_16965);
and U18993 (N_18993,N_12423,N_14274);
nand U18994 (N_18994,N_16725,N_13749);
nand U18995 (N_18995,N_15118,N_14000);
and U18996 (N_18996,N_13855,N_16750);
or U18997 (N_18997,N_17539,N_12574);
or U18998 (N_18998,N_17399,N_13865);
or U18999 (N_18999,N_13985,N_15730);
or U19000 (N_19000,N_16247,N_14537);
nand U19001 (N_19001,N_14124,N_16668);
nand U19002 (N_19002,N_15813,N_17501);
nand U19003 (N_19003,N_12979,N_15004);
nand U19004 (N_19004,N_16540,N_16912);
and U19005 (N_19005,N_13098,N_14739);
nor U19006 (N_19006,N_13482,N_13318);
or U19007 (N_19007,N_17448,N_13657);
or U19008 (N_19008,N_15600,N_14701);
nor U19009 (N_19009,N_12858,N_13785);
xor U19010 (N_19010,N_15935,N_16656);
nor U19011 (N_19011,N_12472,N_15799);
nand U19012 (N_19012,N_13685,N_14744);
nand U19013 (N_19013,N_17828,N_15049);
nor U19014 (N_19014,N_12853,N_16218);
nor U19015 (N_19015,N_12757,N_14684);
nand U19016 (N_19016,N_16566,N_17282);
nand U19017 (N_19017,N_12336,N_12557);
or U19018 (N_19018,N_17460,N_14058);
and U19019 (N_19019,N_15488,N_14533);
or U19020 (N_19020,N_14592,N_15232);
or U19021 (N_19021,N_13218,N_13677);
or U19022 (N_19022,N_13803,N_12430);
nor U19023 (N_19023,N_15688,N_13248);
nand U19024 (N_19024,N_15331,N_14100);
or U19025 (N_19025,N_13039,N_13264);
and U19026 (N_19026,N_16904,N_17365);
xnor U19027 (N_19027,N_12322,N_17549);
nand U19028 (N_19028,N_16881,N_13987);
and U19029 (N_19029,N_16749,N_15665);
or U19030 (N_19030,N_17147,N_12589);
or U19031 (N_19031,N_17119,N_16033);
and U19032 (N_19032,N_14272,N_13467);
and U19033 (N_19033,N_13352,N_12886);
nand U19034 (N_19034,N_14251,N_12681);
nor U19035 (N_19035,N_15415,N_15316);
and U19036 (N_19036,N_16763,N_17435);
nor U19037 (N_19037,N_13066,N_13417);
nand U19038 (N_19038,N_15932,N_12820);
and U19039 (N_19039,N_16106,N_17183);
xnor U19040 (N_19040,N_17263,N_17411);
nand U19041 (N_19041,N_15104,N_17729);
nor U19042 (N_19042,N_17857,N_16551);
nand U19043 (N_19043,N_12499,N_16685);
nor U19044 (N_19044,N_16171,N_12412);
nand U19045 (N_19045,N_17095,N_14548);
nand U19046 (N_19046,N_17970,N_17260);
or U19047 (N_19047,N_17089,N_15013);
and U19048 (N_19048,N_15015,N_16891);
or U19049 (N_19049,N_15572,N_13496);
and U19050 (N_19050,N_14282,N_12545);
xor U19051 (N_19051,N_14761,N_12220);
and U19052 (N_19052,N_17043,N_13724);
nor U19053 (N_19053,N_14195,N_13200);
nand U19054 (N_19054,N_12828,N_16755);
and U19055 (N_19055,N_14877,N_12177);
or U19056 (N_19056,N_12125,N_12675);
nor U19057 (N_19057,N_14321,N_15819);
xnor U19058 (N_19058,N_17875,N_14549);
nor U19059 (N_19059,N_14682,N_12022);
nor U19060 (N_19060,N_17423,N_15186);
nand U19061 (N_19061,N_14524,N_12575);
or U19062 (N_19062,N_15028,N_17640);
or U19063 (N_19063,N_14874,N_16004);
nand U19064 (N_19064,N_17243,N_12416);
nor U19065 (N_19065,N_14020,N_16795);
and U19066 (N_19066,N_12960,N_12462);
nand U19067 (N_19067,N_13225,N_13757);
xnor U19068 (N_19068,N_13047,N_13447);
and U19069 (N_19069,N_12032,N_16839);
and U19070 (N_19070,N_12583,N_13860);
xor U19071 (N_19071,N_17932,N_12579);
nand U19072 (N_19072,N_14516,N_17515);
or U19073 (N_19073,N_14382,N_17641);
nor U19074 (N_19074,N_14370,N_13868);
xnor U19075 (N_19075,N_16226,N_14337);
xor U19076 (N_19076,N_16258,N_14788);
xor U19077 (N_19077,N_12725,N_15313);
nand U19078 (N_19078,N_12053,N_13603);
xor U19079 (N_19079,N_12736,N_15934);
xnor U19080 (N_19080,N_14501,N_13045);
xnor U19081 (N_19081,N_15386,N_13893);
nor U19082 (N_19082,N_17904,N_14918);
xnor U19083 (N_19083,N_15929,N_15950);
xor U19084 (N_19084,N_17324,N_16597);
nand U19085 (N_19085,N_15219,N_12335);
nand U19086 (N_19086,N_13198,N_12263);
nand U19087 (N_19087,N_14072,N_12829);
or U19088 (N_19088,N_13219,N_14111);
or U19089 (N_19089,N_17126,N_15134);
nor U19090 (N_19090,N_14464,N_15562);
or U19091 (N_19091,N_14154,N_12889);
nor U19092 (N_19092,N_15943,N_16820);
nor U19093 (N_19093,N_15741,N_12601);
nor U19094 (N_19094,N_13171,N_13160);
and U19095 (N_19095,N_12713,N_14584);
xor U19096 (N_19096,N_14695,N_15239);
nor U19097 (N_19097,N_17245,N_16204);
and U19098 (N_19098,N_17929,N_14678);
or U19099 (N_19099,N_15843,N_14840);
and U19100 (N_19100,N_12663,N_16266);
or U19101 (N_19101,N_12395,N_16723);
nor U19102 (N_19102,N_12248,N_17381);
xnor U19103 (N_19103,N_16182,N_14733);
and U19104 (N_19104,N_14738,N_13048);
nand U19105 (N_19105,N_17692,N_13209);
nand U19106 (N_19106,N_14362,N_14932);
xor U19107 (N_19107,N_14279,N_16177);
nand U19108 (N_19108,N_15886,N_17951);
xnor U19109 (N_19109,N_14445,N_14604);
xnor U19110 (N_19110,N_15380,N_17955);
nor U19111 (N_19111,N_13930,N_16519);
and U19112 (N_19112,N_12953,N_15803);
or U19113 (N_19113,N_17558,N_15041);
and U19114 (N_19114,N_13931,N_17590);
or U19115 (N_19115,N_16570,N_16330);
and U19116 (N_19116,N_16054,N_13444);
nand U19117 (N_19117,N_15145,N_13829);
nand U19118 (N_19118,N_13302,N_17972);
xnor U19119 (N_19119,N_12050,N_17434);
or U19120 (N_19120,N_16826,N_16609);
nand U19121 (N_19121,N_12212,N_13927);
and U19122 (N_19122,N_15094,N_13547);
xnor U19123 (N_19123,N_17244,N_16130);
nand U19124 (N_19124,N_13595,N_14741);
nand U19125 (N_19125,N_17017,N_17352);
and U19126 (N_19126,N_14131,N_16391);
nand U19127 (N_19127,N_16095,N_17511);
nor U19128 (N_19128,N_13319,N_15809);
and U19129 (N_19129,N_17783,N_13304);
xor U19130 (N_19130,N_16856,N_12251);
nor U19131 (N_19131,N_13001,N_13568);
xnor U19132 (N_19132,N_16800,N_14401);
or U19133 (N_19133,N_13438,N_15141);
xnor U19134 (N_19134,N_12017,N_12748);
or U19135 (N_19135,N_14552,N_12511);
and U19136 (N_19136,N_17114,N_14612);
or U19137 (N_19137,N_14975,N_14677);
xnor U19138 (N_19138,N_12724,N_16848);
nor U19139 (N_19139,N_12927,N_15717);
nand U19140 (N_19140,N_13005,N_12548);
nand U19141 (N_19141,N_12952,N_13443);
or U19142 (N_19142,N_16342,N_14280);
nand U19143 (N_19143,N_15101,N_12684);
nand U19144 (N_19144,N_16769,N_16572);
nor U19145 (N_19145,N_13692,N_13370);
and U19146 (N_19146,N_16140,N_16354);
and U19147 (N_19147,N_16829,N_17070);
or U19148 (N_19148,N_12556,N_17080);
nand U19149 (N_19149,N_13453,N_16959);
xnor U19150 (N_19150,N_14797,N_14074);
xor U19151 (N_19151,N_13303,N_12486);
and U19152 (N_19152,N_15077,N_14996);
nand U19153 (N_19153,N_17959,N_14526);
nand U19154 (N_19154,N_12914,N_13633);
nor U19155 (N_19155,N_12378,N_12839);
nor U19156 (N_19156,N_17891,N_17275);
nand U19157 (N_19157,N_14908,N_17156);
xor U19158 (N_19158,N_12136,N_14910);
xnor U19159 (N_19159,N_13310,N_15268);
nand U19160 (N_19160,N_17213,N_14799);
or U19161 (N_19161,N_17015,N_15920);
or U19162 (N_19162,N_12247,N_16548);
nor U19163 (N_19163,N_13559,N_17486);
nand U19164 (N_19164,N_15582,N_17885);
xnor U19165 (N_19165,N_15689,N_14412);
and U19166 (N_19166,N_12164,N_13152);
nand U19167 (N_19167,N_14264,N_17406);
nor U19168 (N_19168,N_13475,N_16128);
nor U19169 (N_19169,N_15159,N_13134);
nor U19170 (N_19170,N_12163,N_15715);
nor U19171 (N_19171,N_12279,N_16995);
or U19172 (N_19172,N_12308,N_12905);
nor U19173 (N_19173,N_14285,N_14816);
and U19174 (N_19174,N_16430,N_15133);
and U19175 (N_19175,N_12747,N_12316);
and U19176 (N_19176,N_14862,N_13220);
xor U19177 (N_19177,N_14260,N_16397);
xor U19178 (N_19178,N_16882,N_13675);
and U19179 (N_19179,N_13498,N_17014);
xnor U19180 (N_19180,N_14707,N_16847);
xnor U19181 (N_19181,N_13787,N_14243);
or U19182 (N_19182,N_16476,N_12311);
and U19183 (N_19183,N_17050,N_15845);
nand U19184 (N_19184,N_14630,N_16950);
or U19185 (N_19185,N_12532,N_12778);
nand U19186 (N_19186,N_13697,N_15931);
nor U19187 (N_19187,N_13083,N_17605);
and U19188 (N_19188,N_17773,N_14872);
nor U19189 (N_19189,N_15903,N_15190);
xnor U19190 (N_19190,N_13497,N_15509);
or U19191 (N_19191,N_12060,N_15075);
nor U19192 (N_19192,N_13873,N_13429);
xor U19193 (N_19193,N_14775,N_12256);
nand U19194 (N_19194,N_17077,N_12712);
nand U19195 (N_19195,N_12872,N_13731);
and U19196 (N_19196,N_14455,N_17376);
nand U19197 (N_19197,N_17982,N_15424);
xor U19198 (N_19198,N_17185,N_13339);
or U19199 (N_19199,N_14365,N_17262);
xnor U19200 (N_19200,N_15114,N_12994);
nand U19201 (N_19201,N_13488,N_12250);
xnor U19202 (N_19202,N_14520,N_13414);
or U19203 (N_19203,N_16944,N_16604);
or U19204 (N_19204,N_16435,N_16677);
nor U19205 (N_19205,N_17617,N_12843);
or U19206 (N_19206,N_12144,N_14073);
nor U19207 (N_19207,N_13434,N_16952);
and U19208 (N_19208,N_14116,N_16908);
and U19209 (N_19209,N_12349,N_16276);
nand U19210 (N_19210,N_17194,N_16774);
and U19211 (N_19211,N_14945,N_16517);
xnor U19212 (N_19212,N_12173,N_16270);
nor U19213 (N_19213,N_14133,N_16179);
nor U19214 (N_19214,N_14367,N_15957);
or U19215 (N_19215,N_12062,N_14233);
nand U19216 (N_19216,N_16407,N_16762);
and U19217 (N_19217,N_15564,N_14118);
nor U19218 (N_19218,N_12498,N_16573);
or U19219 (N_19219,N_17514,N_13538);
xnor U19220 (N_19220,N_17052,N_17082);
and U19221 (N_19221,N_14915,N_15326);
xnor U19222 (N_19222,N_17208,N_16152);
or U19223 (N_19223,N_17332,N_17199);
nor U19224 (N_19224,N_12744,N_17210);
xnor U19225 (N_19225,N_15459,N_14222);
xor U19226 (N_19226,N_16630,N_14718);
and U19227 (N_19227,N_16061,N_15663);
nand U19228 (N_19228,N_15796,N_12096);
xor U19229 (N_19229,N_14645,N_14657);
nand U19230 (N_19230,N_14278,N_16132);
and U19231 (N_19231,N_16884,N_12510);
xnor U19232 (N_19232,N_13377,N_12563);
and U19233 (N_19233,N_12771,N_14457);
nor U19234 (N_19234,N_17371,N_14336);
nand U19235 (N_19235,N_12842,N_17827);
or U19236 (N_19236,N_17167,N_13143);
nand U19237 (N_19237,N_15918,N_16104);
nor U19238 (N_19238,N_15858,N_14949);
and U19239 (N_19239,N_12968,N_17011);
nand U19240 (N_19240,N_15814,N_15361);
nand U19241 (N_19241,N_17006,N_14490);
nor U19242 (N_19242,N_13608,N_15383);
nand U19243 (N_19243,N_14823,N_16347);
and U19244 (N_19244,N_15558,N_16378);
and U19245 (N_19245,N_14534,N_15797);
nor U19246 (N_19246,N_13979,N_13095);
or U19247 (N_19247,N_17508,N_17425);
and U19248 (N_19248,N_17442,N_13981);
xor U19249 (N_19249,N_15766,N_16924);
or U19250 (N_19250,N_12296,N_12314);
xnor U19251 (N_19251,N_13116,N_14822);
xor U19252 (N_19252,N_14898,N_16633);
or U19253 (N_19253,N_12738,N_15429);
nand U19254 (N_19254,N_15802,N_17531);
nand U19255 (N_19255,N_17814,N_14649);
xor U19256 (N_19256,N_17594,N_15999);
nor U19257 (N_19257,N_16528,N_17206);
and U19258 (N_19258,N_16192,N_13051);
nor U19259 (N_19259,N_17751,N_13075);
or U19260 (N_19260,N_17540,N_15165);
nor U19261 (N_19261,N_17685,N_14654);
nand U19262 (N_19262,N_16116,N_14477);
nand U19263 (N_19263,N_16348,N_14329);
nand U19264 (N_19264,N_15670,N_14702);
and U19265 (N_19265,N_17269,N_13162);
or U19266 (N_19266,N_14421,N_14289);
and U19267 (N_19267,N_15616,N_15794);
xnor U19268 (N_19268,N_13103,N_17518);
nor U19269 (N_19269,N_16530,N_16133);
or U19270 (N_19270,N_16295,N_14724);
nor U19271 (N_19271,N_17267,N_14842);
xnor U19272 (N_19272,N_17321,N_15902);
nand U19273 (N_19273,N_14958,N_17526);
or U19274 (N_19274,N_12466,N_14762);
xor U19275 (N_19275,N_14522,N_12608);
or U19276 (N_19276,N_16473,N_14378);
nand U19277 (N_19277,N_15556,N_17794);
nor U19278 (N_19278,N_15543,N_17478);
or U19279 (N_19279,N_16666,N_13136);
nor U19280 (N_19280,N_17329,N_14936);
and U19281 (N_19281,N_12656,N_14032);
and U19282 (N_19282,N_12396,N_12478);
nand U19283 (N_19283,N_16906,N_14110);
or U19284 (N_19284,N_13254,N_15293);
nor U19285 (N_19285,N_12919,N_12400);
or U19286 (N_19286,N_12138,N_16963);
xnor U19287 (N_19287,N_12056,N_17363);
and U19288 (N_19288,N_12570,N_17799);
and U19289 (N_19289,N_17735,N_16046);
or U19290 (N_19290,N_14573,N_14093);
or U19291 (N_19291,N_13546,N_12543);
xor U19292 (N_19292,N_13897,N_17566);
nor U19293 (N_19293,N_13368,N_13102);
nand U19294 (N_19294,N_12965,N_14881);
or U19295 (N_19295,N_17347,N_13413);
and U19296 (N_19296,N_16543,N_12379);
nor U19297 (N_19297,N_15801,N_15050);
nand U19298 (N_19298,N_13346,N_16049);
xnor U19299 (N_19299,N_17552,N_13741);
and U19300 (N_19300,N_17154,N_13212);
and U19301 (N_19301,N_17266,N_15398);
nor U19302 (N_19302,N_15727,N_13618);
and U19303 (N_19303,N_14964,N_15407);
and U19304 (N_19304,N_14556,N_17270);
nor U19305 (N_19305,N_13324,N_16194);
and U19306 (N_19306,N_14886,N_15861);
xnor U19307 (N_19307,N_17734,N_16417);
nor U19308 (N_19308,N_15739,N_14359);
nand U19309 (N_19309,N_13379,N_12043);
nand U19310 (N_19310,N_17258,N_16638);
or U19311 (N_19311,N_16599,N_13345);
or U19312 (N_19312,N_16801,N_12356);
or U19313 (N_19313,N_12576,N_13332);
and U19314 (N_19314,N_13856,N_12124);
xnor U19315 (N_19315,N_17933,N_17776);
xnor U19316 (N_19316,N_16641,N_17394);
nor U19317 (N_19317,N_16219,N_13184);
nor U19318 (N_19318,N_14340,N_13564);
xnor U19319 (N_19319,N_16184,N_12320);
nor U19320 (N_19320,N_14748,N_15110);
nand U19321 (N_19321,N_17833,N_16327);
nand U19322 (N_19322,N_15153,N_17125);
nand U19323 (N_19323,N_14270,N_13959);
nor U19324 (N_19324,N_13628,N_14843);
nand U19325 (N_19325,N_12692,N_12064);
xor U19326 (N_19326,N_13989,N_14261);
or U19327 (N_19327,N_16098,N_16815);
nand U19328 (N_19328,N_13617,N_17000);
nand U19329 (N_19329,N_13751,N_17373);
xor U19330 (N_19330,N_17466,N_12781);
xor U19331 (N_19331,N_14103,N_17150);
and U19332 (N_19332,N_14883,N_15638);
or U19333 (N_19333,N_14866,N_16558);
or U19334 (N_19334,N_13526,N_15109);
or U19335 (N_19335,N_12765,N_17720);
or U19336 (N_19336,N_15882,N_16210);
xnor U19337 (N_19337,N_13552,N_12640);
xnor U19338 (N_19338,N_13798,N_16437);
or U19339 (N_19339,N_17375,N_16092);
nor U19340 (N_19340,N_13054,N_16620);
or U19341 (N_19341,N_13237,N_15952);
or U19342 (N_19342,N_12000,N_12614);
and U19343 (N_19343,N_15834,N_12223);
xnor U19344 (N_19344,N_15251,N_15345);
or U19345 (N_19345,N_13561,N_16865);
and U19346 (N_19346,N_13331,N_16735);
nand U19347 (N_19347,N_16084,N_16350);
xor U19348 (N_19348,N_14839,N_17153);
nand U19349 (N_19349,N_16587,N_17912);
nand U19350 (N_19350,N_12588,N_15926);
nor U19351 (N_19351,N_17916,N_17498);
nor U19352 (N_19352,N_17110,N_12809);
nand U19353 (N_19353,N_14813,N_13735);
xnor U19354 (N_19354,N_13688,N_13299);
nor U19355 (N_19355,N_14611,N_16369);
and U19356 (N_19356,N_13534,N_15166);
and U19357 (N_19357,N_12776,N_16010);
or U19358 (N_19358,N_15435,N_14527);
or U19359 (N_19359,N_16358,N_15092);
xor U19360 (N_19360,N_17762,N_14493);
or U19361 (N_19361,N_17586,N_14001);
or U19362 (N_19362,N_14576,N_17343);
xor U19363 (N_19363,N_16511,N_15619);
xnor U19364 (N_19364,N_14810,N_17564);
and U19365 (N_19365,N_13149,N_16621);
nand U19366 (N_19366,N_15812,N_13076);
and U19367 (N_19367,N_13591,N_14968);
or U19368 (N_19368,N_12045,N_15514);
nor U19369 (N_19369,N_12824,N_15951);
nor U19370 (N_19370,N_13737,N_12603);
nand U19371 (N_19371,N_14791,N_12741);
nor U19372 (N_19372,N_15449,N_17162);
nand U19373 (N_19373,N_17160,N_15003);
nand U19374 (N_19374,N_17700,N_14593);
nand U19375 (N_19375,N_16139,N_13582);
and U19376 (N_19376,N_15590,N_12039);
xor U19377 (N_19377,N_17781,N_13956);
and U19378 (N_19378,N_14857,N_17472);
and U19379 (N_19379,N_15837,N_15073);
and U19380 (N_19380,N_14219,N_16117);
or U19381 (N_19381,N_16922,N_17032);
nor U19382 (N_19382,N_16379,N_17730);
or U19383 (N_19383,N_14230,N_15818);
nor U19384 (N_19384,N_14873,N_17059);
nand U19385 (N_19385,N_14137,N_16457);
or U19386 (N_19386,N_17780,N_17309);
nand U19387 (N_19387,N_13196,N_16089);
nand U19388 (N_19388,N_14130,N_12390);
and U19389 (N_19389,N_12094,N_17950);
xnor U19390 (N_19390,N_17001,N_12016);
nor U19391 (N_19391,N_13969,N_12176);
xnor U19392 (N_19392,N_17367,N_13101);
or U19393 (N_19393,N_17654,N_15899);
or U19394 (N_19394,N_16316,N_14887);
or U19395 (N_19395,N_15888,N_13156);
and U19396 (N_19396,N_13885,N_15941);
nand U19397 (N_19397,N_12003,N_15339);
nand U19398 (N_19398,N_15731,N_16060);
and U19399 (N_19399,N_17409,N_13527);
nand U19400 (N_19400,N_13316,N_17351);
and U19401 (N_19401,N_17349,N_14034);
xnor U19402 (N_19402,N_14960,N_17099);
nor U19403 (N_19403,N_13966,N_16706);
and U19404 (N_19404,N_13504,N_13649);
xor U19405 (N_19405,N_13129,N_13362);
or U19406 (N_19406,N_14375,N_13878);
or U19407 (N_19407,N_15877,N_13639);
nand U19408 (N_19408,N_15474,N_17071);
or U19409 (N_19409,N_12168,N_16156);
nand U19410 (N_19410,N_17851,N_15945);
xnor U19411 (N_19411,N_16193,N_17013);
xnor U19412 (N_19412,N_17242,N_16673);
nor U19413 (N_19413,N_14313,N_12520);
nor U19414 (N_19414,N_12061,N_15194);
and U19415 (N_19415,N_17364,N_15642);
and U19416 (N_19416,N_13242,N_12020);
nor U19417 (N_19417,N_13210,N_16887);
and U19418 (N_19418,N_14292,N_16893);
or U19419 (N_19419,N_14148,N_15517);
and U19420 (N_19420,N_12512,N_12077);
nor U19421 (N_19421,N_12027,N_13524);
or U19422 (N_19422,N_17964,N_12185);
xor U19423 (N_19423,N_17079,N_17298);
or U19424 (N_19424,N_14806,N_13916);
xor U19425 (N_19425,N_17412,N_16788);
nand U19426 (N_19426,N_15025,N_12796);
or U19427 (N_19427,N_13410,N_13072);
xnor U19428 (N_19428,N_13744,N_13427);
nor U19429 (N_19429,N_15458,N_15357);
xnor U19430 (N_19430,N_12323,N_13027);
nor U19431 (N_19431,N_17707,N_17803);
nor U19432 (N_19432,N_14460,N_16981);
and U19433 (N_19433,N_17568,N_15279);
nor U19434 (N_19434,N_13019,N_16785);
or U19435 (N_19435,N_12848,N_12264);
or U19436 (N_19436,N_16770,N_16867);
xnor U19437 (N_19437,N_17346,N_17750);
and U19438 (N_19438,N_17978,N_17572);
nor U19439 (N_19439,N_13097,N_16227);
xor U19440 (N_19440,N_12253,N_14160);
or U19441 (N_19441,N_17581,N_17782);
nand U19442 (N_19442,N_15065,N_15129);
nor U19443 (N_19443,N_17892,N_12647);
and U19444 (N_19444,N_15489,N_12587);
nand U19445 (N_19445,N_17849,N_16876);
xnor U19446 (N_19446,N_15770,N_17546);
xnor U19447 (N_19447,N_12980,N_14051);
nand U19448 (N_19448,N_15525,N_13140);
nor U19449 (N_19449,N_12737,N_16757);
or U19450 (N_19450,N_15519,N_14712);
nor U19451 (N_19451,N_15559,N_14675);
xnor U19452 (N_19452,N_12095,N_17115);
or U19453 (N_19453,N_17256,N_13375);
xor U19454 (N_19454,N_13841,N_13029);
or U19455 (N_19455,N_12639,N_14235);
or U19456 (N_19456,N_13899,N_16919);
nor U19457 (N_19457,N_15328,N_16874);
nor U19458 (N_19458,N_13124,N_15936);
nor U19459 (N_19459,N_16282,N_13472);
and U19460 (N_19460,N_17400,N_12633);
and U19461 (N_19461,N_16324,N_13532);
or U19462 (N_19462,N_13733,N_13224);
and U19463 (N_19463,N_13663,N_16241);
nor U19464 (N_19464,N_17665,N_14846);
xor U19465 (N_19465,N_14054,N_15782);
xor U19466 (N_19466,N_16042,N_14385);
or U19467 (N_19467,N_13213,N_15360);
xnor U19468 (N_19468,N_13957,N_16453);
nor U19469 (N_19469,N_16222,N_16976);
nor U19470 (N_19470,N_17179,N_12706);
nand U19471 (N_19471,N_17072,N_15410);
nand U19472 (N_19472,N_14906,N_13228);
xor U19473 (N_19473,N_17174,N_15463);
and U19474 (N_19474,N_14296,N_13117);
nor U19475 (N_19475,N_13243,N_15234);
or U19476 (N_19476,N_15522,N_12328);
nor U19477 (N_19477,N_12418,N_12449);
and U19478 (N_19478,N_15143,N_15874);
xnor U19479 (N_19479,N_12782,N_13269);
and U19480 (N_19480,N_13789,N_12698);
and U19481 (N_19481,N_16648,N_13240);
xor U19482 (N_19482,N_13917,N_14417);
or U19483 (N_19483,N_15245,N_16779);
and U19484 (N_19484,N_16196,N_15465);
nand U19485 (N_19485,N_16309,N_12024);
xnor U19486 (N_19486,N_16040,N_14245);
nand U19487 (N_19487,N_12562,N_16514);
nor U19488 (N_19488,N_14331,N_15158);
xnor U19489 (N_19489,N_12391,N_12070);
or U19490 (N_19490,N_16151,N_15396);
or U19491 (N_19491,N_13543,N_17860);
and U19492 (N_19492,N_17664,N_16890);
or U19493 (N_19493,N_13003,N_17771);
or U19494 (N_19494,N_17020,N_15173);
nor U19495 (N_19495,N_12811,N_14698);
or U19496 (N_19496,N_14530,N_15010);
and U19497 (N_19497,N_16304,N_14132);
nor U19498 (N_19498,N_17240,N_16760);
nor U19499 (N_19499,N_12581,N_14557);
nor U19500 (N_19500,N_14931,N_12063);
and U19501 (N_19501,N_13934,N_16026);
and U19502 (N_19502,N_14262,N_17313);
nor U19503 (N_19503,N_13333,N_12728);
nor U19504 (N_19504,N_13708,N_17510);
xnor U19505 (N_19505,N_12295,N_14631);
or U19506 (N_19506,N_13576,N_13624);
xor U19507 (N_19507,N_15230,N_16426);
and U19508 (N_19508,N_15138,N_13208);
or U19509 (N_19509,N_13105,N_16189);
nand U19510 (N_19510,N_15493,N_13723);
or U19511 (N_19511,N_15105,N_16480);
nor U19512 (N_19512,N_14193,N_16123);
or U19513 (N_19513,N_14010,N_14934);
or U19514 (N_19514,N_16338,N_12492);
nor U19515 (N_19515,N_12461,N_13002);
and U19516 (N_19516,N_12835,N_16414);
nand U19517 (N_19517,N_16411,N_13851);
nand U19518 (N_19518,N_17981,N_15167);
nand U19519 (N_19519,N_16999,N_17047);
xor U19520 (N_19520,N_12267,N_15106);
xnor U19521 (N_19521,N_15301,N_15433);
nand U19522 (N_19522,N_17672,N_17116);
nand U19523 (N_19523,N_16439,N_14459);
or U19524 (N_19524,N_15746,N_14651);
or U19525 (N_19525,N_12749,N_16674);
nor U19526 (N_19526,N_16563,N_15865);
xor U19527 (N_19527,N_14021,N_17791);
nor U19528 (N_19528,N_17819,N_15573);
xor U19529 (N_19529,N_12542,N_17921);
xnor U19530 (N_19530,N_13049,N_17004);
nand U19531 (N_19531,N_14825,N_13513);
or U19532 (N_19532,N_12674,N_13190);
or U19533 (N_19533,N_17528,N_15200);
and U19534 (N_19534,N_17138,N_14023);
xnor U19535 (N_19535,N_17936,N_15381);
xor U19536 (N_19536,N_14589,N_15646);
xnor U19537 (N_19537,N_16150,N_15520);
nand U19538 (N_19538,N_16113,N_15961);
and U19539 (N_19539,N_13655,N_17229);
nand U19540 (N_19540,N_12334,N_17850);
xor U19541 (N_19541,N_16387,N_14597);
xnor U19542 (N_19542,N_17101,N_15498);
xor U19543 (N_19543,N_13207,N_16396);
xnor U19544 (N_19544,N_13577,N_13053);
nor U19545 (N_19545,N_16044,N_16091);
xor U19546 (N_19546,N_17378,N_17450);
nor U19547 (N_19547,N_13161,N_15390);
nor U19548 (N_19548,N_15038,N_12135);
xor U19549 (N_19549,N_12621,N_17056);
nand U19550 (N_19550,N_17688,N_17723);
nor U19551 (N_19551,N_17525,N_15116);
nor U19552 (N_19552,N_17923,N_12146);
nand U19553 (N_19553,N_13507,N_14616);
nand U19554 (N_19554,N_15215,N_16889);
or U19555 (N_19555,N_12272,N_13128);
nand U19556 (N_19556,N_15551,N_12228);
nand U19557 (N_19557,N_14141,N_14992);
nand U19558 (N_19558,N_13950,N_17752);
nand U19559 (N_19559,N_12402,N_17067);
xnor U19560 (N_19560,N_12474,N_15675);
and U19561 (N_19561,N_14519,N_14139);
and U19562 (N_19562,N_17181,N_13800);
and U19563 (N_19563,N_17755,N_16314);
nor U19564 (N_19564,N_13480,N_12484);
and U19565 (N_19565,N_15995,N_15425);
xnor U19566 (N_19566,N_14989,N_12118);
or U19567 (N_19567,N_14628,N_17656);
or U19568 (N_19568,N_16665,N_15894);
xor U19569 (N_19569,N_16076,N_17965);
nor U19570 (N_19570,N_14861,N_14605);
or U19571 (N_19571,N_17989,N_14151);
nor U19572 (N_19572,N_14696,N_12457);
nor U19573 (N_19573,N_13694,N_17264);
nor U19574 (N_19574,N_14942,N_15237);
and U19575 (N_19575,N_12417,N_14507);
xnor U19576 (N_19576,N_14607,N_15277);
nor U19577 (N_19577,N_14136,N_17874);
or U19578 (N_19578,N_12844,N_13728);
nand U19579 (N_19579,N_12170,N_16694);
xnor U19580 (N_19580,N_13435,N_16416);
xor U19581 (N_19581,N_17368,N_16208);
and U19582 (N_19582,N_16552,N_15535);
or U19583 (N_19583,N_13146,N_16017);
or U19584 (N_19584,N_17945,N_12134);
xnor U19585 (N_19585,N_12768,N_14366);
or U19586 (N_19586,N_14281,N_15539);
and U19587 (N_19587,N_17390,N_12055);
or U19588 (N_19588,N_12658,N_16484);
nand U19589 (N_19589,N_15351,N_16052);
or U19590 (N_19590,N_17397,N_14869);
xor U19591 (N_19591,N_14019,N_13387);
xnor U19592 (N_19592,N_14834,N_16972);
or U19593 (N_19593,N_13062,N_15225);
nand U19594 (N_19594,N_12700,N_12629);
nor U19595 (N_19595,N_16343,N_17681);
xor U19596 (N_19596,N_13288,N_14425);
xnor U19597 (N_19597,N_16341,N_13110);
nor U19598 (N_19598,N_16843,N_12766);
nor U19599 (N_19599,N_12104,N_15434);
or U19600 (N_19600,N_13502,N_13376);
nor U19601 (N_19601,N_12362,N_12703);
nand U19602 (N_19602,N_17758,N_16730);
nor U19603 (N_19603,N_14713,N_14641);
xor U19604 (N_19604,N_16764,N_12442);
xnor U19605 (N_19605,N_16111,N_16542);
nand U19606 (N_19606,N_16149,N_13344);
nor U19607 (N_19607,N_14146,N_13589);
nand U19608 (N_19608,N_16809,N_16812);
nand U19609 (N_19609,N_13594,N_12568);
or U19610 (N_19610,N_14852,N_14191);
and U19611 (N_19611,N_14715,N_16127);
xor U19612 (N_19612,N_13610,N_14509);
or U19613 (N_19613,N_14298,N_12158);
nand U19614 (N_19614,N_14379,N_17575);
or U19615 (N_19615,N_13016,N_13701);
nor U19616 (N_19616,N_13363,N_12132);
xnor U19617 (N_19617,N_13320,N_13113);
xor U19618 (N_19618,N_16099,N_16836);
or U19619 (N_19619,N_12775,N_14163);
and U19620 (N_19620,N_13875,N_17901);
nor U19621 (N_19621,N_17742,N_14217);
or U19622 (N_19622,N_16038,N_12232);
or U19623 (N_19623,N_15258,N_16623);
nor U19624 (N_19624,N_14395,N_16507);
and U19625 (N_19625,N_16628,N_12153);
or U19626 (N_19626,N_17597,N_12935);
xor U19627 (N_19627,N_16205,N_13073);
xnor U19628 (N_19628,N_17348,N_15298);
nor U19629 (N_19629,N_16323,N_13949);
or U19630 (N_19630,N_14928,N_16639);
and U19631 (N_19631,N_13717,N_12115);
nor U19632 (N_19632,N_15416,N_13279);
nand U19633 (N_19633,N_12951,N_15557);
and U19634 (N_19634,N_12641,N_12018);
and U19635 (N_19635,N_15732,N_17505);
and U19636 (N_19636,N_14088,N_14759);
nor U19637 (N_19637,N_17084,N_13455);
nor U19638 (N_19638,N_14697,N_14571);
or U19639 (N_19639,N_13274,N_14112);
and U19640 (N_19640,N_14443,N_14055);
and U19641 (N_19641,N_13477,N_12431);
and U19642 (N_19642,N_12632,N_12631);
xnor U19643 (N_19643,N_14855,N_12127);
nor U19644 (N_19644,N_16401,N_13262);
or U19645 (N_19645,N_16203,N_14484);
nor U19646 (N_19646,N_14431,N_14084);
nor U19647 (N_19647,N_13558,N_16803);
and U19648 (N_19648,N_17053,N_14444);
or U19649 (N_19649,N_12369,N_16186);
and U19650 (N_19650,N_17674,N_16034);
or U19651 (N_19651,N_13795,N_15427);
or U19652 (N_19652,N_15149,N_14829);
and U19653 (N_19653,N_17237,N_12719);
or U19654 (N_19654,N_12029,N_13721);
or U19655 (N_19655,N_17096,N_17503);
or U19656 (N_19656,N_12387,N_12469);
or U19657 (N_19657,N_12992,N_17545);
nand U19658 (N_19658,N_14500,N_16252);
nand U19659 (N_19659,N_17727,N_15206);
nand U19660 (N_19660,N_17253,N_15297);
or U19661 (N_19661,N_15650,N_16197);
nand U19662 (N_19662,N_13092,N_14990);
nor U19663 (N_19663,N_16529,N_12268);
xnor U19664 (N_19664,N_14026,N_17855);
xnor U19665 (N_19665,N_13834,N_14646);
and U19666 (N_19666,N_12735,N_15596);
nor U19667 (N_19667,N_15876,N_15442);
xor U19668 (N_19668,N_15198,N_14668);
nor U19669 (N_19669,N_15438,N_17339);
nand U19670 (N_19670,N_15974,N_14909);
xnor U19671 (N_19671,N_12344,N_16144);
nor U19672 (N_19672,N_17887,N_15629);
xnor U19673 (N_19673,N_13988,N_15348);
nand U19674 (N_19674,N_16279,N_12421);
nand U19675 (N_19675,N_15684,N_12303);
nor U19676 (N_19676,N_13108,N_14414);
xor U19677 (N_19677,N_16141,N_16969);
xor U19678 (N_19678,N_13943,N_14743);
or U19679 (N_19679,N_15497,N_12455);
xnor U19680 (N_19680,N_14828,N_13634);
nand U19681 (N_19681,N_16544,N_16615);
and U19682 (N_19682,N_17290,N_17312);
nor U19683 (N_19683,N_14914,N_12710);
nor U19684 (N_19684,N_15404,N_14284);
xnor U19685 (N_19685,N_16169,N_13040);
nor U19686 (N_19686,N_12634,N_15184);
nand U19687 (N_19687,N_16814,N_13109);
nor U19688 (N_19688,N_14109,N_17547);
nor U19689 (N_19689,N_16483,N_15823);
and U19690 (N_19690,N_14043,N_17928);
or U19691 (N_19691,N_12555,N_16580);
xnor U19692 (N_19692,N_17766,N_14889);
or U19693 (N_19693,N_16937,N_15311);
nand U19694 (N_19694,N_14333,N_13808);
xnor U19695 (N_19695,N_14817,N_13130);
nor U19696 (N_19696,N_15408,N_14242);
or U19697 (N_19697,N_12204,N_14531);
nand U19698 (N_19698,N_13541,N_16956);
and U19699 (N_19699,N_17760,N_16119);
xnor U19700 (N_19700,N_13236,N_15043);
or U19701 (N_19701,N_14511,N_12434);
nor U19702 (N_19702,N_17614,N_13265);
and U19703 (N_19703,N_13665,N_15402);
nand U19704 (N_19704,N_12534,N_14767);
and U19705 (N_19705,N_17482,N_15549);
nor U19706 (N_19706,N_16619,N_16923);
xnor U19707 (N_19707,N_15925,N_16001);
nand U19708 (N_19708,N_12864,N_12899);
or U19709 (N_19709,N_15625,N_12183);
and U19710 (N_19710,N_15437,N_16823);
nor U19711 (N_19711,N_15323,N_17571);
xor U19712 (N_19712,N_15078,N_14878);
xor U19713 (N_19713,N_12922,N_13791);
nor U19714 (N_19714,N_15955,N_14982);
nor U19715 (N_19715,N_17585,N_15605);
xor U19716 (N_19716,N_14664,N_13114);
nand U19717 (N_19717,N_12572,N_15140);
nor U19718 (N_19718,N_16172,N_15528);
nor U19719 (N_19719,N_15641,N_15550);
or U19720 (N_19720,N_14933,N_17743);
or U19721 (N_19721,N_12995,N_14827);
xnor U19722 (N_19722,N_14448,N_13405);
nand U19723 (N_19723,N_17039,N_15664);
or U19724 (N_19724,N_15762,N_16782);
and U19725 (N_19725,N_12910,N_13881);
nor U19726 (N_19726,N_17035,N_13776);
and U19727 (N_19727,N_15290,N_13193);
nor U19728 (N_19728,N_16055,N_14249);
and U19729 (N_19729,N_12926,N_17403);
xnor U19730 (N_19730,N_13334,N_16957);
xnor U19731 (N_19731,N_15885,N_16808);
xor U19732 (N_19732,N_15652,N_17120);
nand U19733 (N_19733,N_17444,N_13239);
and U19734 (N_19734,N_16422,N_16454);
nand U19735 (N_19735,N_12597,N_17807);
nor U19736 (N_19736,N_13986,N_15668);
or U19737 (N_19737,N_13071,N_14993);
and U19738 (N_19738,N_17106,N_16938);
nand U19739 (N_19739,N_14096,N_13398);
or U19740 (N_19740,N_15306,N_17473);
nor U19741 (N_19741,N_13901,N_14432);
and U19742 (N_19742,N_14447,N_12988);
nand U19743 (N_19743,N_13947,N_17523);
nor U19744 (N_19744,N_17567,N_13226);
xor U19745 (N_19745,N_12594,N_16452);
nor U19746 (N_19746,N_13170,N_13043);
nor U19747 (N_19747,N_13838,N_14040);
xnor U19748 (N_19748,N_14355,N_12357);
or U19749 (N_19749,N_17105,N_17045);
and U19750 (N_19750,N_14138,N_12306);
nand U19751 (N_19751,N_16921,N_12819);
or U19752 (N_19752,N_12803,N_13460);
and U19753 (N_19753,N_14128,N_14049);
or U19754 (N_19754,N_12623,N_17432);
and U19755 (N_19755,N_15417,N_15392);
and U19756 (N_19756,N_16585,N_14772);
nor U19757 (N_19757,N_17164,N_15769);
or U19758 (N_19758,N_14737,N_13764);
or U19759 (N_19759,N_13217,N_12252);
or U19760 (N_19760,N_15883,N_12506);
and U19761 (N_19761,N_15956,N_13948);
xnor U19762 (N_19762,N_13394,N_12445);
nand U19763 (N_19763,N_14473,N_16697);
nand U19764 (N_19764,N_15263,N_12471);
xor U19765 (N_19765,N_14691,N_12481);
xor U19766 (N_19766,N_16699,N_17496);
or U19767 (N_19767,N_13858,N_13953);
nor U19768 (N_19768,N_15139,N_17195);
and U19769 (N_19769,N_17207,N_14632);
xnor U19770 (N_19770,N_14389,N_14561);
nor U19771 (N_19771,N_17690,N_17491);
xnor U19772 (N_19772,N_12909,N_14706);
and U19773 (N_19773,N_16273,N_12325);
nand U19774 (N_19774,N_15791,N_16233);
or U19775 (N_19775,N_16077,N_17815);
or U19776 (N_19776,N_17939,N_14659);
nand U19777 (N_19777,N_16645,N_14052);
nand U19778 (N_19778,N_16916,N_13135);
nand U19779 (N_19779,N_13508,N_12342);
nand U19780 (N_19780,N_16984,N_12977);
nor U19781 (N_19781,N_14426,N_17713);
xor U19782 (N_19782,N_17484,N_12533);
nor U19783 (N_19783,N_12727,N_15910);
and U19784 (N_19784,N_13817,N_12807);
and U19785 (N_19785,N_14753,N_16598);
nand U19786 (N_19786,N_13725,N_17128);
and U19787 (N_19787,N_15763,N_14770);
or U19788 (N_19788,N_15700,N_13347);
or U19789 (N_19789,N_17802,N_12332);
and U19790 (N_19790,N_17028,N_17938);
nand U19791 (N_19791,N_15236,N_13877);
nand U19792 (N_19792,N_16331,N_15088);
nor U19793 (N_19793,N_13174,N_12383);
nand U19794 (N_19794,N_15811,N_14144);
or U19795 (N_19795,N_14240,N_13464);
or U19796 (N_19796,N_17853,N_16502);
xnor U19797 (N_19797,N_16337,N_17158);
nor U19798 (N_19798,N_17103,N_14106);
and U19799 (N_19799,N_15644,N_16732);
xnor U19800 (N_19800,N_17869,N_15728);
or U19801 (N_19801,N_16928,N_12415);
and U19802 (N_19802,N_16145,N_12224);
nor U19803 (N_19803,N_15853,N_14683);
nand U19804 (N_19804,N_16107,N_12709);
and U19805 (N_19805,N_16244,N_13958);
and U19806 (N_19806,N_12717,N_14293);
xnor U19807 (N_19807,N_14396,N_13191);
nand U19808 (N_19808,N_13118,N_16612);
nor U19809 (N_19809,N_17285,N_14328);
and U19810 (N_19810,N_15569,N_16359);
xnor U19811 (N_19811,N_16071,N_15137);
nor U19812 (N_19812,N_15172,N_13481);
nand U19813 (N_19813,N_17428,N_13086);
xnor U19814 (N_19814,N_13471,N_12885);
and U19815 (N_19815,N_16275,N_14066);
xnor U19816 (N_19816,N_12624,N_14502);
xnor U19817 (N_19817,N_17439,N_12271);
or U19818 (N_19818,N_15829,N_16964);
nor U19819 (N_19819,N_12970,N_14948);
nor U19820 (N_19820,N_14255,N_17132);
and U19821 (N_19821,N_16355,N_16500);
xnor U19822 (N_19822,N_14383,N_13593);
and U19823 (N_19823,N_17710,N_15304);
nand U19824 (N_19824,N_12593,N_12841);
nor U19825 (N_19825,N_12815,N_12866);
nor U19826 (N_19826,N_15606,N_13861);
nand U19827 (N_19827,N_13063,N_16983);
nor U19828 (N_19828,N_15863,N_17836);
xnor U19829 (N_19829,N_17646,N_13567);
and U19830 (N_19830,N_14896,N_16786);
and U19831 (N_19831,N_16384,N_15687);
nor U19832 (N_19832,N_14803,N_14172);
xor U19833 (N_19833,N_16647,N_12305);
nor U19834 (N_19834,N_17949,N_14271);
xnor U19835 (N_19835,N_16614,N_15589);
nand U19836 (N_19836,N_14354,N_16066);
nor U19837 (N_19837,N_12281,N_15254);
or U19838 (N_19838,N_12480,N_17778);
or U19839 (N_19839,N_13211,N_17247);
and U19840 (N_19840,N_15896,N_12081);
nor U19841 (N_19841,N_16857,N_17910);
xnor U19842 (N_19842,N_17703,N_15062);
nand U19843 (N_19843,N_13205,N_12874);
nor U19844 (N_19844,N_16844,N_16497);
xor U19845 (N_19845,N_13578,N_16590);
or U19846 (N_19846,N_17480,N_12282);
nand U19847 (N_19847,N_15850,N_16948);
or U19848 (N_19848,N_13469,N_16900);
nand U19849 (N_19849,N_12302,N_12566);
nor U19850 (N_19850,N_13971,N_17902);
and U19851 (N_19851,N_13823,N_15447);
and U19852 (N_19852,N_17226,N_16272);
or U19853 (N_19853,N_12456,N_13924);
xor U19854 (N_19854,N_14381,N_13715);
nor U19855 (N_19855,N_15854,N_16707);
and U19856 (N_19856,N_15656,N_16982);
nand U19857 (N_19857,N_17768,N_12008);
or U19858 (N_19858,N_13425,N_14127);
nor U19859 (N_19859,N_17618,N_15653);
nor U19860 (N_19860,N_14663,N_14204);
or U19861 (N_19861,N_15907,N_15160);
xor U19862 (N_19862,N_14740,N_13954);
nand U19863 (N_19863,N_12243,N_12635);
nand U19864 (N_19864,N_16832,N_17689);
or U19865 (N_19865,N_16804,N_12812);
nand U19866 (N_19866,N_15836,N_17487);
nand U19867 (N_19867,N_16498,N_12221);
nor U19868 (N_19868,N_17139,N_12827);
xor U19869 (N_19869,N_17859,N_16428);
xnor U19870 (N_19870,N_14363,N_17709);
or U19871 (N_19871,N_14608,N_13298);
and U19872 (N_19872,N_17302,N_16251);
nor U19873 (N_19873,N_13711,N_14016);
or U19874 (N_19874,N_14826,N_12870);
nand U19875 (N_19875,N_15185,N_12284);
nand U19876 (N_19876,N_15542,N_13275);
and U19877 (N_19877,N_12394,N_17813);
and U19878 (N_19878,N_15735,N_17230);
nand U19879 (N_19879,N_16980,N_14924);
nand U19880 (N_19880,N_13554,N_17044);
or U19881 (N_19881,N_17415,N_16185);
nor U19882 (N_19882,N_12515,N_12742);
nor U19883 (N_19883,N_16905,N_15533);
and U19884 (N_19884,N_15672,N_14056);
nor U19885 (N_19885,N_17879,N_17651);
nand U19886 (N_19886,N_14558,N_15872);
xnor U19887 (N_19887,N_17705,N_12139);
and U19888 (N_19888,N_13107,N_16108);
and U19889 (N_19889,N_17610,N_12350);
nor U19890 (N_19890,N_15315,N_15176);
nand U19891 (N_19891,N_12716,N_15706);
nand U19892 (N_19892,N_15898,N_13600);
or U19893 (N_19893,N_15144,N_14888);
or U19894 (N_19894,N_15513,N_12192);
or U19895 (N_19895,N_17745,N_14332);
or U19896 (N_19896,N_16032,N_12759);
xnor U19897 (N_19897,N_12116,N_15122);
nand U19898 (N_19898,N_17062,N_12464);
nand U19899 (N_19899,N_14188,N_16722);
nor U19900 (N_19900,N_16068,N_16027);
and U19901 (N_19901,N_13503,N_15302);
xor U19902 (N_19902,N_15494,N_16606);
or U19903 (N_19903,N_12453,N_12554);
nor U19904 (N_19904,N_13119,N_16575);
or U19905 (N_19905,N_13622,N_17500);
xnor U19906 (N_19906,N_13535,N_15636);
nand U19907 (N_19907,N_12160,N_12999);
nor U19908 (N_19908,N_14069,N_17854);
nand U19909 (N_19909,N_13849,N_15249);
and U19910 (N_19910,N_14959,N_16539);
xnor U19911 (N_19911,N_14905,N_13483);
or U19912 (N_19912,N_14086,N_14768);
xnor U19913 (N_19913,N_14517,N_15148);
nor U19914 (N_19914,N_15349,N_16508);
nand U19915 (N_19915,N_12437,N_15199);
or U19916 (N_19916,N_14804,N_17893);
and U19917 (N_19917,N_15291,N_17733);
nor U19918 (N_19918,N_12122,N_15506);
or U19919 (N_19919,N_12620,N_16713);
or U19920 (N_19920,N_15373,N_16989);
and U19921 (N_19921,N_16315,N_13765);
and U19922 (N_19922,N_12549,N_14897);
nand U19923 (N_19923,N_16992,N_16320);
xnor U19924 (N_19924,N_12359,N_13827);
nor U19925 (N_19925,N_14966,N_16545);
or U19926 (N_19926,N_12496,N_16293);
and U19927 (N_19927,N_17331,N_15400);
nor U19928 (N_19928,N_17519,N_16901);
and U19929 (N_19929,N_14642,N_17022);
nand U19930 (N_19930,N_14725,N_15496);
nor U19931 (N_19931,N_13176,N_15355);
or U19932 (N_19932,N_12784,N_13139);
nor U19933 (N_19933,N_14259,N_15793);
and U19934 (N_19934,N_14048,N_14462);
nor U19935 (N_19935,N_14014,N_13000);
or U19936 (N_19936,N_15944,N_16506);
or U19937 (N_19937,N_17280,N_16030);
nand U19938 (N_19938,N_12560,N_12660);
nor U19939 (N_19939,N_13925,N_13572);
xor U19940 (N_19940,N_14453,N_15074);
or U19941 (N_19941,N_15196,N_12800);
nor U19942 (N_19942,N_12906,N_16394);
nor U19943 (N_19943,N_16008,N_16209);
or U19944 (N_19944,N_13343,N_15939);
and U19945 (N_19945,N_16557,N_14508);
xor U19946 (N_19946,N_14711,N_13740);
nand U19947 (N_19947,N_16561,N_12341);
nand U19948 (N_19948,N_12664,N_16326);
nand U19949 (N_19949,N_16102,N_12298);
xor U19950 (N_19950,N_16531,N_14560);
and U19951 (N_19951,N_17171,N_15781);
nor U19952 (N_19952,N_17763,N_16813);
or U19953 (N_19953,N_17871,N_12476);
nand U19954 (N_19954,N_16361,N_17002);
or U19955 (N_19955,N_15295,N_16103);
xnor U19956 (N_19956,N_16231,N_15027);
or U19957 (N_19957,N_12657,N_15716);
or U19958 (N_19958,N_15047,N_16014);
nor U19959 (N_19959,N_14311,N_13079);
or U19960 (N_19960,N_14358,N_12758);
and U19961 (N_19961,N_12373,N_15515);
and U19962 (N_19962,N_17359,N_13544);
and U19963 (N_19963,N_14237,N_15593);
nand U19964 (N_19964,N_15161,N_12943);
xor U19965 (N_19965,N_16290,N_16146);
nor U19966 (N_19966,N_16584,N_16657);
xnor U19967 (N_19967,N_16998,N_14539);
or U19968 (N_19968,N_12826,N_12351);
or U19969 (N_19969,N_13614,N_13597);
nor U19970 (N_19970,N_15738,N_13666);
or U19971 (N_19971,N_17424,N_14650);
nor U19972 (N_19972,N_14785,N_17041);
nand U19973 (N_19973,N_13300,N_15299);
xnor U19974 (N_19974,N_16595,N_17234);
nand U19975 (N_19975,N_13710,N_14917);
xnor U19976 (N_19976,N_16257,N_16777);
and U19977 (N_19977,N_13253,N_15678);
nor U19978 (N_19978,N_17784,N_13909);
nand U19979 (N_19979,N_17201,N_14595);
nor U19980 (N_19980,N_14763,N_13641);
and U19981 (N_19981,N_14140,N_13389);
or U19982 (N_19982,N_15457,N_13840);
xor U19983 (N_19983,N_16710,N_13911);
or U19984 (N_19984,N_12216,N_13439);
nor U19985 (N_19985,N_17289,N_16340);
or U19986 (N_19986,N_13709,N_13922);
nand U19987 (N_19987,N_13784,N_13815);
or U19988 (N_19988,N_14377,N_15921);
and U19989 (N_19989,N_12519,N_13181);
or U19990 (N_19990,N_14734,N_15132);
nor U19991 (N_19991,N_14206,N_15300);
and U19992 (N_19992,N_12278,N_16445);
nand U19993 (N_19993,N_15054,N_12682);
xor U19994 (N_19994,N_17130,N_12538);
xor U19995 (N_19995,N_15369,N_15142);
nor U19996 (N_19996,N_15702,N_13604);
and U19997 (N_19997,N_13995,N_13993);
nand U19998 (N_19998,N_12584,N_12794);
and U19999 (N_19999,N_15908,N_15395);
xor U20000 (N_20000,N_16447,N_14876);
or U20001 (N_20001,N_14621,N_14437);
nand U20002 (N_20002,N_12859,N_15491);
xor U20003 (N_20003,N_14574,N_15538);
nor U20004 (N_20004,N_12273,N_16409);
and U20005 (N_20005,N_17250,N_13206);
xnor U20006 (N_20006,N_17957,N_15949);
nor U20007 (N_20007,N_17499,N_17198);
xnor U20008 (N_20008,N_14618,N_13122);
nor U20009 (N_20009,N_14101,N_12883);
or U20010 (N_20010,N_17852,N_13041);
or U20011 (N_20011,N_13403,N_12409);
nor U20012 (N_20012,N_15005,N_16807);
and U20013 (N_20013,N_16488,N_16933);
or U20014 (N_20014,N_13702,N_13199);
nand U20015 (N_20015,N_12005,N_15353);
xor U20016 (N_20016,N_12734,N_17488);
xnor U20017 (N_20017,N_14614,N_14350);
nand U20018 (N_20018,N_17048,N_13400);
nor U20019 (N_20019,N_12141,N_13658);
xnor U20020 (N_20020,N_12523,N_13301);
and U20021 (N_20021,N_13919,N_13351);
or U20022 (N_20022,N_14726,N_14665);
nand U20023 (N_20023,N_13216,N_15370);
or U20024 (N_20024,N_17344,N_15084);
or U20025 (N_20025,N_14523,N_17947);
or U20026 (N_20026,N_12958,N_12237);
and U20027 (N_20027,N_16581,N_14757);
and U20028 (N_20028,N_17619,N_15374);
nand U20029 (N_20029,N_13631,N_14091);
nand U20030 (N_20030,N_17152,N_14789);
or U20031 (N_20031,N_17986,N_14787);
nor U20032 (N_20032,N_13067,N_15456);
nor U20033 (N_20033,N_12377,N_15867);
or U20034 (N_20034,N_16079,N_16333);
or U20035 (N_20035,N_16523,N_15901);
and U20036 (N_20036,N_15227,N_13131);
nand U20037 (N_20037,N_17725,N_15401);
xnor U20038 (N_20038,N_12851,N_17769);
and U20039 (N_20039,N_15734,N_16024);
xnor U20040 (N_20040,N_13251,N_15477);
and U20041 (N_20041,N_13990,N_17224);
xnor U20042 (N_20042,N_12677,N_14998);
nand U20043 (N_20043,N_12932,N_15151);
or U20044 (N_20044,N_15422,N_14427);
and U20045 (N_20045,N_13489,N_13177);
nand U20046 (N_20046,N_13495,N_12058);
or U20047 (N_20047,N_17872,N_17714);
xnor U20048 (N_20048,N_15726,N_14463);
and U20049 (N_20049,N_16878,N_17281);
xnor U20050 (N_20050,N_13994,N_14540);
and U20051 (N_20051,N_17124,N_14879);
or U20052 (N_20052,N_12030,N_14890);
xor U20053 (N_20053,N_13830,N_15452);
and U20054 (N_20054,N_14790,N_16365);
nor U20055 (N_20055,N_14147,N_14095);
xor U20056 (N_20056,N_17797,N_12089);
or U20057 (N_20057,N_14736,N_17451);
nor U20058 (N_20058,N_12188,N_12933);
or U20059 (N_20059,N_17042,N_15790);
nor U20060 (N_20060,N_15612,N_13235);
or U20061 (N_20061,N_15181,N_15830);
or U20062 (N_20062,N_17788,N_13879);
or U20063 (N_20063,N_13961,N_12246);
xor U20064 (N_20064,N_13844,N_14832);
and U20065 (N_20065,N_17969,N_15917);
or U20066 (N_20066,N_13520,N_14951);
or U20067 (N_20067,N_13999,N_17239);
nor U20068 (N_20068,N_16427,N_12167);
or U20069 (N_20069,N_16277,N_12202);
nor U20070 (N_20070,N_17209,N_12026);
and U20071 (N_20071,N_17311,N_14178);
and U20072 (N_20072,N_12986,N_14283);
nand U20073 (N_20073,N_14904,N_16799);
xor U20074 (N_20074,N_12755,N_12021);
nand U20075 (N_20075,N_12103,N_16410);
xor U20076 (N_20076,N_12255,N_12333);
nand U20077 (N_20077,N_13234,N_16910);
nor U20078 (N_20078,N_14900,N_12165);
and U20079 (N_20079,N_12033,N_13750);
and U20080 (N_20080,N_13669,N_16649);
xnor U20081 (N_20081,N_16601,N_15385);
nand U20082 (N_20082,N_16242,N_15560);
nand U20083 (N_20083,N_16469,N_17161);
xor U20084 (N_20084,N_14470,N_12401);
or U20085 (N_20085,N_14202,N_12286);
xnor U20086 (N_20086,N_14694,N_15244);
or U20087 (N_20087,N_16086,N_12025);
xnor U20088 (N_20088,N_16190,N_16915);
nor U20089 (N_20089,N_13586,N_16157);
xor U20090 (N_20090,N_16962,N_13933);
nor U20091 (N_20091,N_12438,N_14082);
nand U20092 (N_20092,N_14341,N_14075);
xnor U20093 (N_20093,N_12638,N_15099);
or U20094 (N_20094,N_14467,N_12880);
and U20095 (N_20095,N_17323,N_13926);
or U20096 (N_20096,N_15723,N_16424);
or U20097 (N_20097,N_16550,N_14080);
nand U20098 (N_20098,N_16349,N_14002);
and U20099 (N_20099,N_17315,N_16468);
nand U20100 (N_20100,N_16712,N_12275);
xnor U20101 (N_20101,N_14482,N_15510);
xnor U20102 (N_20102,N_13908,N_14708);
nor U20103 (N_20103,N_17992,N_12950);
and U20104 (N_20104,N_16596,N_12211);
nand U20105 (N_20105,N_16069,N_16562);
nand U20106 (N_20106,N_14610,N_12106);
and U20107 (N_20107,N_16072,N_16020);
or U20108 (N_20108,N_12830,N_12266);
nand U20109 (N_20109,N_13652,N_13974);
nand U20110 (N_20110,N_17136,N_12291);
or U20111 (N_20111,N_16138,N_13064);
and U20112 (N_20112,N_12370,N_16824);
or U20113 (N_20113,N_17121,N_17238);
nor U20114 (N_20114,N_15842,N_15981);
nor U20115 (N_20115,N_15859,N_14247);
xnor U20116 (N_20116,N_14323,N_15887);
or U20117 (N_20117,N_15737,N_17535);
nor U20118 (N_20118,N_14735,N_17228);
xnor U20119 (N_20119,N_14838,N_12961);
xnor U20120 (N_20120,N_12225,N_17054);
nand U20121 (N_20121,N_13748,N_14625);
or U20122 (N_20122,N_14256,N_16681);
and U20123 (N_20123,N_14070,N_14398);
nor U20124 (N_20124,N_14210,N_14173);
xor U20125 (N_20125,N_16724,N_17764);
xor U20126 (N_20126,N_15822,N_17231);
nor U20127 (N_20127,N_12213,N_17360);
nand U20128 (N_20128,N_16446,N_13099);
nor U20129 (N_20129,N_14756,N_14891);
and U20130 (N_20130,N_13297,N_17886);
xnor U20131 (N_20131,N_13436,N_15547);
nand U20132 (N_20132,N_13505,N_15757);
and U20133 (N_20133,N_12726,N_13459);
or U20134 (N_20134,N_13295,N_17388);
nand U20135 (N_20135,N_12785,N_16470);
nor U20136 (N_20136,N_15703,N_17683);
nand U20137 (N_20137,N_15532,N_13753);
xor U20138 (N_20138,N_15229,N_14807);
or U20139 (N_20139,N_17715,N_15776);
or U20140 (N_20140,N_13420,N_15691);
xor U20141 (N_20141,N_16831,N_14123);
xnor U20142 (N_20142,N_13428,N_12946);
nor U20143 (N_20143,N_12235,N_17977);
and U20144 (N_20144,N_14687,N_13790);
and U20145 (N_20145,N_12605,N_16789);
and U20146 (N_20146,N_13290,N_16124);
or U20147 (N_20147,N_15785,N_16793);
and U20148 (N_20148,N_17261,N_15701);
and U20149 (N_20149,N_16737,N_17922);
nand U20150 (N_20150,N_16176,N_12928);
nor U20151 (N_20151,N_16698,N_12304);
xor U20152 (N_20152,N_16643,N_12447);
and U20153 (N_20153,N_17149,N_16862);
xor U20154 (N_20154,N_14515,N_14306);
and U20155 (N_20155,N_17647,N_15682);
nand U20156 (N_20156,N_16287,N_16253);
nand U20157 (N_20157,N_12233,N_15889);
nor U20158 (N_20158,N_14175,N_13173);
nor U20159 (N_20159,N_12348,N_13770);
and U20160 (N_20160,N_12976,N_12731);
or U20161 (N_20161,N_13506,N_12756);
and U20162 (N_20162,N_16994,N_12787);
or U20163 (N_20163,N_16221,N_15658);
xnor U20164 (N_20164,N_13522,N_12879);
nand U20165 (N_20165,N_16993,N_16687);
nor U20166 (N_20166,N_15816,N_16930);
or U20167 (N_20167,N_16317,N_14672);
and U20168 (N_20168,N_17556,N_16122);
or U20169 (N_20169,N_16260,N_12231);
or U20170 (N_20170,N_14114,N_12850);
xnor U20171 (N_20171,N_15617,N_17630);
or U20172 (N_20172,N_12745,N_16569);
and U20173 (N_20173,N_17650,N_15620);
nand U20174 (N_20174,N_16794,N_13382);
nand U20175 (N_20175,N_15588,N_12707);
or U20176 (N_20176,N_16344,N_15131);
and U20177 (N_20177,N_17436,N_15697);
and U20178 (N_20178,N_17643,N_12073);
or U20179 (N_20179,N_17068,N_14488);
nor U20180 (N_20180,N_16495,N_14721);
xor U20181 (N_20181,N_17353,N_16932);
or U20182 (N_20182,N_15964,N_17322);
and U20183 (N_20183,N_14225,N_13006);
or U20184 (N_20184,N_12236,N_17613);
nand U20185 (N_20185,N_15677,N_17273);
nor U20186 (N_20186,N_12861,N_12339);
nor U20187 (N_20187,N_14907,N_17903);
xor U20188 (N_20188,N_15828,N_14215);
xor U20189 (N_20189,N_16683,N_12704);
or U20190 (N_20190,N_17792,N_14581);
nor U20191 (N_20191,N_13656,N_12643);
nor U20192 (N_20192,N_16640,N_12673);
nand U20193 (N_20193,N_16220,N_16375);
nor U20194 (N_20194,N_12004,N_15405);
or U20195 (N_20195,N_13277,N_12667);
or U20196 (N_20196,N_16255,N_17061);
nor U20197 (N_20197,N_16860,N_13626);
or U20198 (N_20198,N_13644,N_17822);
nand U20199 (N_20199,N_16267,N_12653);
and U20200 (N_20200,N_13895,N_12360);
nand U20201 (N_20201,N_17465,N_13805);
and U20202 (N_20202,N_13852,N_17274);
nor U20203 (N_20203,N_14920,N_16631);
or U20204 (N_20204,N_15113,N_15492);
and U20205 (N_20205,N_15403,N_13910);
and U20206 (N_20206,N_17897,N_14729);
and U20207 (N_20207,N_14895,N_14190);
or U20208 (N_20208,N_14212,N_16841);
xor U20209 (N_20209,N_16418,N_14871);
nand U20210 (N_20210,N_16776,N_14689);
xor U20211 (N_20211,N_12199,N_15826);
or U20212 (N_20212,N_13154,N_17184);
and U20213 (N_20213,N_17542,N_17490);
nand U20214 (N_20214,N_12862,N_16885);
and U20215 (N_20215,N_12299,N_17452);
nor U20216 (N_20216,N_16903,N_17884);
xnor U20217 (N_20217,N_12426,N_12131);
xor U20218 (N_20218,N_12277,N_16421);
or U20219 (N_20219,N_16931,N_17653);
nor U20220 (N_20220,N_17034,N_13771);
nor U20221 (N_20221,N_16626,N_16112);
nand U20222 (N_20222,N_13752,N_13662);
xor U20223 (N_20223,N_12893,N_15271);
nor U20224 (N_20224,N_15787,N_17301);
nand U20225 (N_20225,N_15511,N_17517);
and U20226 (N_20226,N_14461,N_16087);
xnor U20227 (N_20227,N_12913,N_12732);
or U20228 (N_20228,N_15916,N_17372);
nand U20229 (N_20229,N_17083,N_14633);
or U20230 (N_20230,N_13530,N_16588);
nand U20231 (N_20231,N_14181,N_16025);
and U20232 (N_20232,N_16936,N_14901);
xor U20233 (N_20233,N_12178,N_13565);
nand U20234 (N_20234,N_15912,N_12808);
or U20235 (N_20235,N_12301,N_14805);
or U20236 (N_20236,N_13147,N_17534);
xnor U20237 (N_20237,N_14022,N_17785);
xnor U20238 (N_20238,N_14241,N_17249);
or U20239 (N_20239,N_12964,N_14679);
xnor U20240 (N_20240,N_16524,N_14566);
or U20241 (N_20241,N_13463,N_16526);
or U20242 (N_20242,N_15661,N_12693);
nand U20243 (N_20243,N_16655,N_12847);
and U20244 (N_20244,N_15063,N_16684);
and U20245 (N_20245,N_12454,N_15037);
xnor U20246 (N_20246,N_13714,N_15983);
or U20247 (N_20247,N_16048,N_15666);
or U20248 (N_20248,N_13432,N_14087);
nor U20249 (N_20249,N_13747,N_14266);
or U20250 (N_20250,N_14596,N_15231);
and U20251 (N_20251,N_15608,N_15567);
xnor U20252 (N_20252,N_13153,N_14547);
nor U20253 (N_20253,N_12067,N_13336);
xnor U20254 (N_20254,N_16215,N_14288);
nor U20255 (N_20255,N_12528,N_17615);
nor U20256 (N_20256,N_12128,N_16768);
or U20257 (N_20257,N_16652,N_17606);
nand U20258 (N_20258,N_12093,N_14166);
xnor U20259 (N_20259,N_13022,N_13703);
nand U20260 (N_20260,N_13182,N_12875);
and U20261 (N_20261,N_14499,N_15322);
xnor U20262 (N_20262,N_17748,N_13121);
and U20263 (N_20263,N_14911,N_17063);
xor U20264 (N_20264,N_15123,N_16136);
nand U20265 (N_20265,N_15986,N_16955);
or U20266 (N_20266,N_17708,N_17233);
xor U20267 (N_20267,N_17396,N_13214);
nand U20268 (N_20268,N_17392,N_16403);
or U20269 (N_20269,N_13635,N_16003);
and U20270 (N_20270,N_17670,N_13308);
or U20271 (N_20271,N_17953,N_13231);
xor U20272 (N_20272,N_15275,N_15324);
nor U20273 (N_20273,N_15048,N_16985);
nand U20274 (N_20274,N_16537,N_16065);
or U20275 (N_20275,N_17141,N_16166);
nor U20276 (N_20276,N_16747,N_12714);
nand U20277 (N_20277,N_17662,N_14497);
nand U20278 (N_20278,N_15342,N_14648);
nor U20279 (N_20279,N_13773,N_14546);
and U20280 (N_20280,N_12353,N_16991);
or U20281 (N_20281,N_16971,N_12982);
nor U20282 (N_20282,N_14794,N_12036);
xor U20283 (N_20283,N_17917,N_14348);
nor U20284 (N_20284,N_13754,N_14435);
nand U20285 (N_20285,N_16143,N_16285);
nand U20286 (N_20286,N_12082,N_13548);
nand U20287 (N_20287,N_15384,N_14231);
and U20288 (N_20288,N_12346,N_17337);
or U20289 (N_20289,N_14119,N_16929);
and U20290 (N_20290,N_16064,N_15838);
xor U20291 (N_20291,N_12881,N_15680);
nor U20292 (N_20292,N_15079,N_17187);
and U20293 (N_20293,N_15841,N_13025);
or U20294 (N_20294,N_12645,N_12309);
or U20295 (N_20295,N_15991,N_16851);
nand U20296 (N_20296,N_14976,N_15436);
nand U20297 (N_20297,N_17716,N_13323);
or U20298 (N_20298,N_14258,N_15262);
nor U20299 (N_20299,N_13317,N_15135);
nor U20300 (N_20300,N_13923,N_13259);
nand U20301 (N_20301,N_13273,N_15485);
and U20302 (N_20302,N_14373,N_16353);
or U20303 (N_20303,N_13163,N_14504);
nor U20304 (N_20304,N_14987,N_13123);
nand U20305 (N_20305,N_16328,N_17268);
nor U20306 (N_20306,N_12078,N_16164);
and U20307 (N_20307,N_15928,N_13907);
nand U20308 (N_20308,N_15314,N_14135);
or U20309 (N_20309,N_14894,N_14325);
nor U20310 (N_20310,N_13381,N_15019);
and U20311 (N_20311,N_13772,N_17954);
nor U20312 (N_20312,N_17561,N_17532);
nor U20313 (N_20313,N_17212,N_15548);
nand U20314 (N_20314,N_12978,N_16213);
and U20315 (N_20315,N_12473,N_13070);
xor U20316 (N_20316,N_16873,N_14532);
or U20317 (N_20317,N_17570,N_14952);
nand U20318 (N_20318,N_13035,N_17580);
nor U20319 (N_20319,N_13575,N_15375);
and U20320 (N_20320,N_16695,N_16907);
or U20321 (N_20321,N_12823,N_16765);
nand U20322 (N_20322,N_14849,N_17211);
xnor U20323 (N_20323,N_14441,N_12789);
or U20324 (N_20324,N_14716,N_16047);
nand U20325 (N_20325,N_12140,N_16960);
or U20326 (N_20326,N_12270,N_15089);
xor U20327 (N_20327,N_13020,N_15987);
nor U20328 (N_20328,N_14468,N_14194);
or U20329 (N_20329,N_12619,N_15444);
or U20330 (N_20330,N_13839,N_15601);
or U20331 (N_20331,N_16827,N_16180);
or U20332 (N_20332,N_16618,N_16080);
nor U20333 (N_20333,N_13967,N_13686);
xnor U20334 (N_20334,N_16676,N_12625);
nor U20335 (N_20335,N_16863,N_15431);
or U20336 (N_20336,N_15202,N_15708);
or U20337 (N_20337,N_15246,N_14559);
nand U20338 (N_20338,N_13501,N_15033);
xnor U20339 (N_20339,N_12319,N_14669);
or U20340 (N_20340,N_13080,N_12786);
nand U20341 (N_20341,N_13892,N_16942);
nand U20342 (N_20342,N_16162,N_12628);
nand U20343 (N_20343,N_14169,N_13846);
or U20344 (N_20344,N_12206,N_12531);
or U20345 (N_20345,N_15758,N_16752);
nor U20346 (N_20346,N_15856,N_13531);
nand U20347 (N_20347,N_15259,N_16958);
and U20348 (N_20348,N_15495,N_14197);
xor U20349 (N_20349,N_13831,N_16308);
nand U20350 (N_20350,N_15667,N_12689);
xor U20351 (N_20351,N_12019,N_16458);
nand U20352 (N_20352,N_12547,N_16448);
and U20353 (N_20353,N_14731,N_15552);
and U20354 (N_20354,N_12347,N_15870);
xor U20355 (N_20355,N_12007,N_13736);
and U20356 (N_20356,N_14478,N_15387);
and U20357 (N_20357,N_12162,N_17668);
or U20358 (N_20358,N_16703,N_15815);
nand U20359 (N_20359,N_15468,N_13004);
xor U20360 (N_20360,N_13695,N_14656);
nor U20361 (N_20361,N_13551,N_15690);
or U20362 (N_20362,N_13145,N_13011);
and U20363 (N_20363,N_12925,N_15683);
nor U20364 (N_20364,N_14297,N_16206);
and U20365 (N_20365,N_15764,N_13215);
and U20366 (N_20366,N_17123,N_17308);
xnor U20367 (N_20367,N_14586,N_14613);
nand U20368 (N_20368,N_15993,N_17221);
and U20369 (N_20369,N_16871,N_12410);
nand U20370 (N_20370,N_12315,N_14200);
or U20371 (N_20371,N_16201,N_15714);
and U20372 (N_20372,N_13941,N_13412);
and U20373 (N_20373,N_15992,N_12930);
xnor U20374 (N_20374,N_13918,N_13914);
xnor U20375 (N_20375,N_15017,N_15946);
nand U20376 (N_20376,N_13960,N_17461);
and U20377 (N_20377,N_15647,N_17663);
xnor U20378 (N_20378,N_13549,N_15213);
nand U20379 (N_20379,N_14647,N_14046);
nand U20380 (N_20380,N_17808,N_13033);
xnor U20381 (N_20381,N_14085,N_15976);
nand U20382 (N_20382,N_16897,N_17178);
xnor U20383 (N_20383,N_16622,N_17930);
nor U20384 (N_20384,N_16830,N_13276);
or U20385 (N_20385,N_13038,N_14104);
or U20386 (N_20386,N_17426,N_17112);
nand U20387 (N_20387,N_17467,N_14357);
xor U20388 (N_20388,N_17754,N_17675);
nor U20389 (N_20389,N_14038,N_13416);
nor U20390 (N_20390,N_15789,N_17481);
nand U20391 (N_20391,N_12098,N_13458);
and U20392 (N_20392,N_13350,N_13536);
or U20393 (N_20393,N_17454,N_16997);
nand U20394 (N_20394,N_16485,N_12521);
and U20395 (N_20395,N_12149,N_13938);
xnor U20396 (N_20396,N_14637,N_15377);
xor U20397 (N_20397,N_15265,N_13529);
or U20398 (N_20398,N_13383,N_17881);
nand U20399 (N_20399,N_16481,N_14680);
nand U20400 (N_20400,N_14525,N_13779);
nand U20401 (N_20401,N_13074,N_15508);
nor U20402 (N_20402,N_16842,N_13014);
or U20403 (N_20403,N_12971,N_14860);
and U20404 (N_20404,N_14535,N_12218);
nor U20405 (N_20405,N_12938,N_13936);
nor U20406 (N_20406,N_12822,N_16741);
nor U20407 (N_20407,N_14635,N_14690);
nor U20408 (N_20408,N_13585,N_17841);
nand U20409 (N_20409,N_15839,N_17811);
xnor U20410 (N_20410,N_16806,N_15610);
xor U20411 (N_20411,N_12366,N_16953);
nor U20412 (N_20412,N_15214,N_12863);
and U20413 (N_20413,N_16798,N_16211);
nor U20414 (N_20414,N_17574,N_17962);
and U20415 (N_20415,N_17387,N_17196);
or U20416 (N_20416,N_17456,N_12425);
and U20417 (N_20417,N_13144,N_17652);
xor U20418 (N_20418,N_14882,N_17550);
nand U20419 (N_20419,N_17319,N_14120);
or U20420 (N_20420,N_13358,N_12343);
nor U20421 (N_20421,N_13204,N_16039);
and U20422 (N_20422,N_14988,N_14582);
nand U20423 (N_20423,N_16477,N_13862);
nor U20424 (N_20424,N_17395,N_12901);
nand U20425 (N_20425,N_17075,N_14751);
xnor U20426 (N_20426,N_15034,N_15804);
or U20427 (N_20427,N_12997,N_16866);
or U20428 (N_20428,N_12276,N_12262);
nand U20429 (N_20429,N_13386,N_17876);
or U20430 (N_20430,N_13055,N_13611);
and U20431 (N_20431,N_12013,N_15031);
nor U20432 (N_20432,N_12526,N_14991);
nor U20433 (N_20433,N_12987,N_13090);
nor U20434 (N_20434,N_13975,N_12544);
or U20435 (N_20435,N_16363,N_15968);
and U20436 (N_20436,N_12269,N_15626);
nor U20437 (N_20437,N_15969,N_14406);
and U20438 (N_20438,N_15469,N_16386);
nand U20439 (N_20439,N_13629,N_12770);
xor U20440 (N_20440,N_16753,N_14782);
or U20441 (N_20441,N_15627,N_14619);
nor U20442 (N_20442,N_16796,N_13078);
xnor U20443 (N_20443,N_14946,N_13810);
or U20444 (N_20444,N_13866,N_12836);
or U20445 (N_20445,N_17864,N_17279);
nor U20446 (N_20446,N_14536,N_17483);
and U20447 (N_20447,N_13499,N_13249);
nor U20448 (N_20448,N_12596,N_16711);
or U20449 (N_20449,N_17009,N_12491);
and U20450 (N_20450,N_17303,N_12300);
and U20451 (N_20451,N_16013,N_17868);
nand U20452 (N_20452,N_12609,N_12783);
or U20453 (N_20453,N_14415,N_14113);
xnor U20454 (N_20454,N_17862,N_17379);
and U20455 (N_20455,N_17040,N_12595);
xor U20456 (N_20456,N_15657,N_14974);
nand U20457 (N_20457,N_16739,N_14667);
nor U20458 (N_20458,N_15312,N_16680);
and U20459 (N_20459,N_14326,N_15947);
nor U20460 (N_20460,N_16239,N_12559);
nand U20461 (N_20461,N_13996,N_16364);
xnor U20462 (N_20462,N_14732,N_12711);
or U20463 (N_20463,N_14666,N_12651);
nor U20464 (N_20464,N_17060,N_15443);
nand U20465 (N_20465,N_16745,N_13945);
nor U20466 (N_20466,N_16225,N_16482);
nand U20467 (N_20467,N_13028,N_15500);
nor U20468 (N_20468,N_14786,N_14685);
xor U20469 (N_20469,N_12119,N_14126);
nand U20470 (N_20470,N_14439,N_17168);
and U20471 (N_20471,N_13903,N_14174);
nor U20472 (N_20472,N_13632,N_14824);
xor U20473 (N_20473,N_16883,N_14324);
nand U20474 (N_20474,N_16926,N_14471);
nand U20475 (N_20475,N_13645,N_14575);
nand U20476 (N_20476,N_12503,N_17840);
xor U20477 (N_20477,N_15222,N_17522);
nand U20478 (N_20478,N_12929,N_12317);
nor U20479 (N_20479,N_17846,N_12490);
nand U20480 (N_20480,N_14276,N_15168);
and U20481 (N_20481,N_12730,N_14728);
xor U20482 (N_20482,N_13449,N_15274);
nor U20483 (N_20483,N_12238,N_13667);
or U20484 (N_20484,N_15659,N_17291);
nand U20485 (N_20485,N_17926,N_17883);
and U20486 (N_20486,N_12773,N_16560);
xor U20487 (N_20487,N_17595,N_12849);
nor U20488 (N_20488,N_13268,N_12405);
nand U20489 (N_20489,N_16366,N_15914);
xnor U20490 (N_20490,N_12895,N_17983);
xor U20491 (N_20491,N_13180,N_13824);
or U20492 (N_20492,N_13642,N_13462);
nor U20493 (N_20493,N_15007,N_16627);
nand U20494 (N_20494,N_12101,N_15052);
nor U20495 (N_20495,N_13833,N_15544);
and U20496 (N_20496,N_17717,N_12470);
nor U20497 (N_20497,N_12208,N_15645);
and U20498 (N_20498,N_14498,N_17915);
or U20499 (N_20499,N_12739,N_12210);
nor U20500 (N_20500,N_15393,N_16288);
nor U20501 (N_20501,N_12097,N_16377);
nand U20502 (N_20502,N_12429,N_17069);
nand U20503 (N_20503,N_15996,N_14720);
and U20504 (N_20504,N_14676,N_12904);
nor U20505 (N_20505,N_16838,N_15997);
xnor U20506 (N_20506,N_17777,N_13037);
nand U20507 (N_20507,N_13256,N_12637);
nand U20508 (N_20508,N_17753,N_14899);
or U20509 (N_20509,N_12618,N_12386);
xnor U20510 (N_20510,N_12948,N_12483);
or U20511 (N_20511,N_16105,N_17602);
and U20512 (N_20512,N_16527,N_13245);
or U20513 (N_20513,N_12414,N_17232);
and U20514 (N_20514,N_17413,N_16237);
and U20515 (N_20515,N_17591,N_16229);
nor U20516 (N_20516,N_15721,N_17579);
nand U20517 (N_20517,N_12219,N_15775);
xnor U20518 (N_20518,N_14416,N_17419);
and U20519 (N_20519,N_16456,N_14971);
or U20520 (N_20520,N_12615,N_13670);
and U20521 (N_20521,N_14953,N_12896);
and U20522 (N_20522,N_15389,N_16374);
nand U20523 (N_20523,N_16945,N_15501);
nand U20524 (N_20524,N_17122,N_14187);
nand U20525 (N_20525,N_17728,N_17844);
nand U20526 (N_20526,N_12497,N_15879);
nand U20527 (N_20527,N_15284,N_13825);
and U20528 (N_20528,N_17706,N_13653);
nor U20529 (N_20529,N_16294,N_17457);
and U20530 (N_20530,N_16383,N_14122);
nor U20531 (N_20531,N_12630,N_12654);
nor U20532 (N_20532,N_14077,N_13921);
or U20533 (N_20533,N_14402,N_14814);
xor U20534 (N_20534,N_13696,N_12723);
nor U20535 (N_20535,N_12229,N_15391);
nor U20536 (N_20536,N_15761,N_14134);
or U20537 (N_20537,N_13271,N_14821);
xnor U20538 (N_20538,N_12746,N_14079);
nor U20539 (N_20539,N_14820,N_17648);
nor U20540 (N_20540,N_14662,N_13883);
xor U20541 (N_20541,N_15965,N_13402);
and U20542 (N_20542,N_16390,N_15609);
and U20543 (N_20543,N_14218,N_15855);
xor U20544 (N_20544,N_15773,N_12817);
and U20545 (N_20545,N_14754,N_12600);
and U20546 (N_20546,N_15209,N_17430);
nand U20547 (N_20547,N_17036,N_17677);
xnor U20548 (N_20548,N_16302,N_13013);
nand U20549 (N_20549,N_15093,N_17599);
or U20550 (N_20550,N_14606,N_16126);
nand U20551 (N_20551,N_15193,N_12337);
nand U20552 (N_20552,N_13647,N_16845);
nor U20553 (N_20553,N_17848,N_13880);
nand U20554 (N_20554,N_12996,N_13853);
and U20555 (N_20555,N_16074,N_12443);
and U20556 (N_20556,N_16636,N_12505);
or U20557 (N_20557,N_15527,N_12816);
xnor U20558 (N_20558,N_15919,N_12652);
nor U20559 (N_20559,N_13620,N_14727);
or U20560 (N_20560,N_12945,N_14773);
xnor U20561 (N_20561,N_17971,N_14203);
and U20562 (N_20562,N_17441,N_15971);
or U20563 (N_20563,N_12810,N_16740);
nand U20564 (N_20564,N_15006,N_14388);
nand U20565 (N_20565,N_13036,N_16412);
or U20566 (N_20566,N_15871,N_16522);
nand U20567 (N_20567,N_16880,N_15696);
xor U20568 (N_20568,N_15545,N_15120);
nand U20569 (N_20569,N_13690,N_12463);
or U20570 (N_20570,N_16148,N_14777);
nand U20571 (N_20571,N_17446,N_12529);
nand U20572 (N_20572,N_13085,N_12436);
xnor U20573 (N_20573,N_14440,N_15825);
xnor U20574 (N_20574,N_15335,N_15962);
nand U20575 (N_20575,N_15090,N_12606);
nand U20576 (N_20576,N_15428,N_17757);
nor U20577 (N_20577,N_13061,N_12420);
or U20578 (N_20578,N_17453,N_15806);
nor U20579 (N_20579,N_17091,N_16898);
and U20580 (N_20580,N_12939,N_12552);
or U20581 (N_20581,N_12427,N_13247);
and U20582 (N_20582,N_12984,N_12194);
nor U20583 (N_20583,N_17801,N_12200);
or U20584 (N_20584,N_15978,N_12385);
or U20585 (N_20585,N_15927,N_17533);
nor U20586 (N_20586,N_13857,N_14409);
and U20587 (N_20587,N_14830,N_16037);
nor U20588 (N_20588,N_12147,N_13816);
nand U20589 (N_20589,N_17669,N_12989);
nand U20590 (N_20590,N_17507,N_13706);
nand U20591 (N_20591,N_17988,N_12051);
nand U20592 (N_20592,N_16036,N_15044);
and U20593 (N_20593,N_13569,N_12975);
xor U20594 (N_20594,N_17335,N_13396);
nand U20595 (N_20595,N_17134,N_17882);
xor U20596 (N_20596,N_16053,N_12460);
nor U20597 (N_20597,N_12459,N_16125);
and U20598 (N_20598,N_16515,N_15892);
xnor U20599 (N_20599,N_14142,N_16634);
or U20600 (N_20600,N_15203,N_14634);
nand U20601 (N_20601,N_16406,N_13059);
xor U20602 (N_20602,N_17445,N_14965);
nand U20603 (N_20603,N_16062,N_17341);
nor U20604 (N_20604,N_17934,N_12249);
and U20605 (N_20605,N_16402,N_13093);
and U20606 (N_20606,N_17354,N_15897);
and U20607 (N_20607,N_15486,N_14003);
nor U20608 (N_20608,N_13555,N_12791);
and U20609 (N_20609,N_15267,N_14752);
nor U20610 (N_20610,N_12508,N_16607);
nand U20611 (N_20611,N_14859,N_14615);
or U20612 (N_20612,N_12364,N_17679);
or U20613 (N_20613,N_12234,N_13700);
xnor U20614 (N_20614,N_16729,N_12685);
or U20615 (N_20615,N_13390,N_14579);
nor U20616 (N_20616,N_15591,N_14769);
or U20617 (N_20617,N_12205,N_17440);
and U20618 (N_20618,N_15432,N_14864);
nand U20619 (N_20619,N_16503,N_16925);
nand U20620 (N_20620,N_15252,N_13571);
and U20621 (N_20621,N_17131,N_17197);
xnor U20622 (N_20622,N_14353,N_15264);
and U20623 (N_20623,N_15127,N_15150);
xor U20624 (N_20624,N_17741,N_12868);
xor U20625 (N_20625,N_17246,N_13293);
and U20626 (N_20626,N_16207,N_13484);
nand U20627 (N_20627,N_16892,N_16336);
nand U20628 (N_20628,N_15273,N_16644);
and U20629 (N_20629,N_12292,N_13327);
or U20630 (N_20630,N_14670,N_17049);
and U20631 (N_20631,N_15729,N_12090);
xnor U20632 (N_20632,N_14983,N_15988);
xor U20633 (N_20633,N_15388,N_14456);
nor U20634 (N_20634,N_12527,N_14380);
and U20635 (N_20635,N_12777,N_17304);
nor U20636 (N_20636,N_16214,N_14583);
xor U20637 (N_20637,N_13263,N_15182);
or U20638 (N_20638,N_13835,N_17443);
or U20639 (N_20639,N_12368,N_15597);
or U20640 (N_20640,N_15121,N_16761);
nor U20641 (N_20641,N_13322,N_14316);
xor U20642 (N_20642,N_17393,N_15217);
nand U20643 (N_20643,N_15847,N_15915);
xor U20644 (N_20644,N_13407,N_14778);
xnor U20645 (N_20645,N_14994,N_12793);
nor U20646 (N_20646,N_17300,N_13052);
xnor U20647 (N_20647,N_17170,N_13451);
xor U20648 (N_20648,N_16509,N_17418);
nand U20649 (N_20649,N_13759,N_17935);
nand U20650 (N_20650,N_14884,N_13766);
xor U20651 (N_20651,N_13281,N_15453);
nand U20652 (N_20652,N_16318,N_16475);
xnor U20653 (N_20653,N_14495,N_14795);
nand U20654 (N_20654,N_12500,N_15980);
and U20655 (N_20655,N_16372,N_17021);
nor U20656 (N_20656,N_16775,N_16097);
xor U20657 (N_20657,N_12222,N_16975);
and U20658 (N_20658,N_15082,N_17686);
and U20659 (N_20659,N_12954,N_17600);
nor U20660 (N_20660,N_13915,N_15341);
and U20661 (N_20661,N_17913,N_16440);
xnor U20662 (N_20662,N_15171,N_12662);
or U20663 (N_20663,N_12363,N_13819);
or U20664 (N_20664,N_16002,N_16568);
xnor U20665 (N_20665,N_17543,N_17582);
xnor U20666 (N_20666,N_17306,N_12898);
or U20667 (N_20667,N_16501,N_14157);
and U20668 (N_20668,N_13616,N_12949);
nor U20669 (N_20669,N_15788,N_17861);
and U20670 (N_20670,N_14248,N_12585);
nor U20671 (N_20671,N_12920,N_16083);
xnor U20672 (N_20672,N_12774,N_17296);
or U20673 (N_20673,N_15076,N_17286);
and U20674 (N_20674,N_12539,N_12180);
xor U20675 (N_20675,N_12912,N_12743);
and U20676 (N_20676,N_17133,N_15221);
and U20677 (N_20677,N_17429,N_15909);
nor U20678 (N_20678,N_16460,N_13581);
or U20679 (N_20679,N_17736,N_14352);
xnor U20680 (N_20680,N_17975,N_17941);
nand U20681 (N_20681,N_14544,N_16413);
nor U20682 (N_20682,N_12659,N_15873);
xnor U20683 (N_20683,N_14372,N_12580);
nor U20684 (N_20684,N_17223,N_17816);
or U20685 (N_20685,N_14926,N_15175);
nand U20686 (N_20686,N_13516,N_14213);
or U20687 (N_20687,N_16978,N_15180);
or U20688 (N_20688,N_16704,N_12475);
and U20689 (N_20689,N_15783,N_16616);
nand U20690 (N_20690,N_13397,N_17404);
and U20691 (N_20691,N_12701,N_17382);
nand U20692 (N_20692,N_16702,N_17527);
xnor U20693 (N_20693,N_12287,N_14505);
nand U20694 (N_20694,N_14036,N_16451);
or U20695 (N_20695,N_17747,N_12916);
nor U20696 (N_20696,N_15937,N_17896);
nand U20697 (N_20697,N_13419,N_17919);
nor U20698 (N_20698,N_15490,N_12088);
and U20699 (N_20699,N_16015,N_16541);
nand U20700 (N_20700,N_15278,N_13952);
nand U20701 (N_20701,N_17489,N_14912);
and U20702 (N_20702,N_17817,N_14267);
nand U20703 (N_20703,N_17414,N_15577);
xor U20704 (N_20704,N_14746,N_16970);
nand U20705 (N_20705,N_15966,N_13266);
nand U20706 (N_20706,N_17994,N_12345);
and U20707 (N_20707,N_13970,N_12993);
or U20708 (N_20708,N_14176,N_14793);
or U20709 (N_20709,N_14489,N_17944);
nor U20710 (N_20710,N_15628,N_16688);
nand U20711 (N_20711,N_16941,N_14955);
xnor U20712 (N_20712,N_12113,N_16935);
or U20713 (N_20713,N_13258,N_15308);
or U20714 (N_20714,N_16986,N_17191);
nor U20715 (N_20715,N_12245,N_14474);
nand U20716 (N_20716,N_12937,N_12918);
nor U20717 (N_20717,N_15798,N_16869);
or U20718 (N_20718,N_14369,N_12079);
nand U20719 (N_20719,N_13896,N_13326);
or U20720 (N_20720,N_15719,N_15201);
nand U20721 (N_20721,N_13314,N_17297);
or U20722 (N_20722,N_15774,N_12666);
nand U20723 (N_20723,N_16212,N_15163);
xnor U20724 (N_20724,N_17673,N_13681);
nand U20725 (N_20725,N_14652,N_12908);
xnor U20726 (N_20726,N_16094,N_14730);
or U20727 (N_20727,N_15948,N_12074);
nand U20728 (N_20728,N_16659,N_13734);
nand U20729 (N_20729,N_15835,N_14094);
nand U20730 (N_20730,N_15977,N_13179);
nand U20731 (N_20731,N_15570,N_12086);
or U20732 (N_20732,N_16110,N_16063);
nor U20733 (N_20733,N_15022,N_16549);
xor U20734 (N_20734,N_15611,N_16135);
and U20735 (N_20735,N_14317,N_12514);
or U20736 (N_20736,N_17789,N_16041);
or U20737 (N_20737,N_17236,N_14334);
and U20738 (N_20738,N_12915,N_17506);
xnor U20739 (N_20739,N_17824,N_13983);
or U20740 (N_20740,N_17818,N_15382);
xor U20741 (N_20741,N_12182,N_12175);
nor U20742 (N_20742,N_12432,N_17998);
and U20743 (N_20743,N_13433,N_12517);
xor U20744 (N_20744,N_17449,N_17345);
xor U20745 (N_20745,N_17384,N_15679);
xnor U20746 (N_20746,N_15030,N_17960);
and U20747 (N_20747,N_13112,N_12705);
nor U20748 (N_20748,N_13813,N_15753);
and U20749 (N_20749,N_13057,N_14145);
nand U20750 (N_20750,N_17544,N_14620);
xor U20751 (N_20751,N_15096,N_13044);
nand U20752 (N_20752,N_13566,N_14486);
and U20753 (N_20753,N_17899,N_16918);
xnor U20754 (N_20754,N_17405,N_12196);
xnor U20755 (N_20755,N_15516,N_12931);
and U20756 (N_20756,N_16271,N_17696);
xor U20757 (N_20757,N_15455,N_17193);
xor U20758 (N_20758,N_14580,N_12155);
nor U20759 (N_20759,N_16516,N_14050);
or U20760 (N_20760,N_12444,N_14935);
nor U20761 (N_20761,N_13238,N_14588);
xor U20762 (N_20762,N_15070,N_14201);
and U20763 (N_20763,N_12372,N_16433);
nor U20764 (N_20764,N_14623,N_12507);
xnor U20765 (N_20765,N_14294,N_12288);
nor U20766 (N_20766,N_13664,N_16510);
nor U20767 (N_20767,N_13312,N_16280);
nor U20768 (N_20768,N_14957,N_15975);
nor U20769 (N_20769,N_12942,N_12376);
xnor U20770 (N_20770,N_15319,N_13166);
xor U20771 (N_20771,N_14152,N_14562);
xnor U20772 (N_20772,N_14760,N_17925);
xnor U20773 (N_20773,N_13636,N_15631);
and U20774 (N_20774,N_16155,N_17631);
or U20775 (N_20775,N_17660,N_14196);
and U20776 (N_20776,N_16746,N_16870);
nand U20777 (N_20777,N_14226,N_15309);
nor U20778 (N_20778,N_13687,N_12504);
nand U20779 (N_20779,N_13932,N_12041);
nor U20780 (N_20780,N_17093,N_14442);
nand U20781 (N_20781,N_14913,N_13430);
nand U20782 (N_20782,N_14483,N_13500);
xor U20783 (N_20783,N_17639,N_15499);
or U20784 (N_20784,N_15632,N_14543);
and U20785 (N_20785,N_15011,N_14149);
nor U20786 (N_20786,N_17420,N_16028);
xnor U20787 (N_20787,N_15624,N_13977);
or U20788 (N_20788,N_17607,N_15307);
xnor U20789 (N_20789,N_14067,N_12424);
xnor U20790 (N_20790,N_15942,N_16235);
and U20791 (N_20791,N_17421,N_12407);
nand U20792 (N_20792,N_12257,N_12066);
or U20793 (N_20793,N_15216,N_15233);
xnor U20794 (N_20794,N_12217,N_16216);
nor U20795 (N_20795,N_16319,N_16852);
nor U20796 (N_20796,N_14037,N_15824);
xnor U20797 (N_20797,N_13233,N_16949);
and U20798 (N_20798,N_17166,N_17509);
nor U20799 (N_20799,N_14257,N_12900);
nor U20800 (N_20800,N_14387,N_17995);
xnor U20801 (N_20801,N_12037,N_15820);
nand U20802 (N_20802,N_13106,N_14999);
nand U20803 (N_20803,N_14250,N_13515);
xor U20804 (N_20804,N_16646,N_14078);
and U20805 (N_20805,N_17259,N_17671);
nand U20806 (N_20806,N_12627,N_17278);
nor U20807 (N_20807,N_14045,N_12482);
nand U20808 (N_20808,N_15541,N_14599);
nand U20809 (N_20809,N_17030,N_15602);
or U20810 (N_20810,N_12371,N_15693);
and U20811 (N_20811,N_15805,N_16886);
nor U20812 (N_20812,N_14180,N_14344);
nand U20813 (N_20813,N_13359,N_16093);
xnor U20814 (N_20814,N_15621,N_13422);
nand U20815 (N_20815,N_13026,N_16675);
and U20816 (N_20816,N_13511,N_13601);
and U20817 (N_20817,N_17798,N_17155);
nand U20818 (N_20818,N_15223,N_16546);
nor U20819 (N_20819,N_16431,N_16660);
or U20820 (N_20820,N_16380,N_16429);
and U20821 (N_20821,N_14029,N_16142);
nor U20822 (N_20822,N_12612,N_13388);
xnor U20823 (N_20823,N_17104,N_17288);
xnor U20824 (N_20824,N_16705,N_16462);
nand U20825 (N_20825,N_16228,N_13431);
nand U20826 (N_20826,N_15905,N_17756);
or U20827 (N_20827,N_16245,N_15587);
or U20828 (N_20828,N_14423,N_12169);
or U20829 (N_20829,N_17693,N_17968);
nor U20830 (N_20830,N_16736,N_12644);
and U20831 (N_20831,N_17504,N_16487);
xnor U20832 (N_20832,N_15368,N_15576);
nand U20833 (N_20833,N_15032,N_14514);
or U20834 (N_20834,N_17608,N_13836);
and U20835 (N_20835,N_14044,N_14304);
or U20836 (N_20836,N_17369,N_17598);
or U20837 (N_20837,N_15083,N_17635);
xnor U20838 (N_20838,N_14062,N_15095);
or U20839 (N_20839,N_16305,N_16400);
nand U20840 (N_20840,N_14275,N_14312);
or U20841 (N_20841,N_12981,N_15253);
xor U20842 (N_20842,N_12642,N_14033);
or U20843 (N_20843,N_12720,N_12354);
xnor U20844 (N_20844,N_14802,N_16088);
xnor U20845 (N_20845,N_12280,N_16243);
and U20846 (N_20846,N_15462,N_17192);
or U20847 (N_20847,N_16432,N_14277);
nor U20848 (N_20848,N_15571,N_14068);
nand U20849 (N_20849,N_14268,N_13964);
nor U20850 (N_20850,N_16654,N_15911);
or U20851 (N_20851,N_12764,N_17842);
and U20852 (N_20852,N_16298,N_17272);
or U20853 (N_20853,N_13809,N_15933);
or U20854 (N_20854,N_17573,N_14783);
or U20855 (N_20855,N_15470,N_12028);
and U20856 (N_20856,N_16672,N_15303);
nand U20857 (N_20857,N_15002,N_13774);
or U20858 (N_20858,N_12567,N_12610);
and U20859 (N_20859,N_17621,N_12516);
and U20860 (N_20860,N_15112,N_16954);
xnor U20861 (N_20861,N_12691,N_12550);
nor U20862 (N_20862,N_12769,N_16389);
nand U20863 (N_20863,N_12047,N_16658);
or U20864 (N_20864,N_14594,N_12294);
xnor U20865 (N_20865,N_14057,N_15071);
or U20866 (N_20866,N_17966,N_14214);
nor U20867 (N_20867,N_15891,N_17536);
xnor U20868 (N_20868,N_12622,N_14004);
xor U20869 (N_20869,N_16423,N_16158);
nor U20870 (N_20870,N_17786,N_14480);
or U20871 (N_20871,N_16472,N_13148);
and U20872 (N_20872,N_17825,N_13155);
or U20873 (N_20873,N_16849,N_15439);
or U20874 (N_20874,N_16352,N_14386);
and U20875 (N_20875,N_12752,N_13356);
nor U20876 (N_20876,N_13982,N_12121);
or U20877 (N_20877,N_17642,N_12329);
nand U20878 (N_20878,N_17327,N_17569);
xnor U20879 (N_20879,N_15989,N_14808);
nor U20880 (N_20880,N_15100,N_15164);
and U20881 (N_20881,N_12957,N_17163);
nor U20882 (N_20882,N_16442,N_16669);
or U20883 (N_20883,N_15272,N_15598);
xor U20884 (N_20884,N_14818,N_15056);
xnor U20885 (N_20885,N_15081,N_13252);
or U20886 (N_20886,N_16291,N_15188);
xnor U20887 (N_20887,N_15269,N_15585);
nand U20888 (N_20888,N_12324,N_15226);
nor U20889 (N_20889,N_14863,N_14986);
nand U20890 (N_20890,N_12068,N_13450);
xnor U20891 (N_20891,N_15372,N_14220);
nand U20892 (N_20892,N_15247,N_15024);
and U20893 (N_20893,N_15866,N_13756);
and U20894 (N_20894,N_17046,N_13768);
or U20895 (N_20895,N_13355,N_17737);
xor U20896 (N_20896,N_17200,N_16240);
and U20897 (N_20897,N_16610,N_16611);
nand U20898 (N_20898,N_15257,N_15344);
xnor U20899 (N_20899,N_13393,N_16310);
and U20900 (N_20900,N_13365,N_16532);
or U20901 (N_20901,N_14747,N_15338);
and U20902 (N_20902,N_17633,N_13380);
and U20903 (N_20903,N_13192,N_16198);
xor U20904 (N_20904,N_17724,N_13137);
nand U20905 (N_20905,N_14699,N_17721);
xnor U20906 (N_20906,N_13291,N_16693);
or U20907 (N_20907,N_17227,N_16625);
or U20908 (N_20908,N_12151,N_16163);
nand U20909 (N_20909,N_13583,N_14681);
xor U20910 (N_20910,N_12289,N_16299);
nand U20911 (N_20911,N_16463,N_15779);
or U20912 (N_20912,N_14542,N_14590);
or U20913 (N_20913,N_12403,N_17731);
nand U20914 (N_20914,N_14506,N_14469);
nand U20915 (N_20915,N_17462,N_12446);
or U20916 (N_20916,N_16322,N_12338);
or U20917 (N_20917,N_13168,N_14766);
and U20918 (N_20918,N_17906,N_12242);
xnor U20919 (N_20919,N_14947,N_13296);
nor U20920 (N_20920,N_17870,N_13068);
nand U20921 (N_20921,N_14405,N_14984);
xnor U20922 (N_20922,N_15792,N_14962);
xnor U20923 (N_20923,N_14047,N_16165);
nor U20924 (N_20924,N_17386,N_14674);
nor U20925 (N_20925,N_14371,N_13454);
nor U20926 (N_20926,N_12985,N_15352);
xnor U20927 (N_20927,N_15294,N_17355);
or U20928 (N_20928,N_16853,N_16101);
nand U20929 (N_20929,N_16154,N_15869);
nand U20930 (N_20930,N_13778,N_13648);
xnor U20931 (N_20931,N_16939,N_16246);
xnor U20932 (N_20932,N_12087,N_13164);
and U20933 (N_20933,N_12100,N_17823);
or U20934 (N_20934,N_13132,N_12171);
or U20935 (N_20935,N_14413,N_15574);
nor U20936 (N_20936,N_14658,N_17804);
nor U20937 (N_20937,N_16576,N_13169);
xor U20938 (N_20938,N_17661,N_15979);
nand U20939 (N_20939,N_12112,N_15399);
nor U20940 (N_20940,N_16191,N_17026);
xnor U20941 (N_20941,N_14941,N_15651);
or U20942 (N_20942,N_13523,N_12046);
or U20943 (N_20943,N_15973,N_12244);
xnor U20944 (N_20944,N_13782,N_14364);
and U20945 (N_20945,N_16109,N_15540);
and U20946 (N_20946,N_13309,N_17370);
nand U20947 (N_20947,N_13306,N_16471);
or U20948 (N_20948,N_13602,N_12561);
xnor U20949 (N_20949,N_17391,N_12522);
or U20950 (N_20950,N_14705,N_13755);
nor U20951 (N_20951,N_16671,N_17702);
nand U20952 (N_20952,N_16555,N_17292);
and U20953 (N_20953,N_17159,N_16943);
nor U20954 (N_20954,N_17401,N_17235);
nand U20955 (N_20955,N_17038,N_17732);
nand U20956 (N_20956,N_16268,N_14551);
xnor U20957 (N_20957,N_17326,N_15524);
nor U20958 (N_20958,N_17521,N_16600);
or U20959 (N_20959,N_12668,N_16035);
nand U20960 (N_20960,N_13605,N_16608);
and U20961 (N_20961,N_17625,N_14053);
xor U20962 (N_20962,N_13718,N_12944);
nor U20963 (N_20963,N_12598,N_12941);
xor U20964 (N_20964,N_15851,N_16718);
nand U20965 (N_20965,N_13573,N_15205);
nand U20966 (N_20966,N_12297,N_17475);
or U20967 (N_20967,N_16264,N_14503);
nor U20968 (N_20968,N_15266,N_17055);
nand U20969 (N_20969,N_13769,N_13470);
and U20970 (N_20970,N_17900,N_17385);
or U20971 (N_20971,N_15162,N_14198);
and U20972 (N_20972,N_14330,N_16443);
xnor U20973 (N_20973,N_16236,N_16822);
and U20974 (N_20974,N_16603,N_15440);
nor U20975 (N_20975,N_16797,N_12397);
or U20976 (N_20976,N_12911,N_13017);
and U20977 (N_20977,N_13126,N_17623);
and U20978 (N_20978,N_14184,N_17888);
nand U20979 (N_20979,N_14320,N_15614);
xnor U20980 (N_20980,N_15461,N_14880);
nor U20981 (N_20981,N_14587,N_16325);
xor U20982 (N_20982,N_16459,N_14229);
xor U20983 (N_20983,N_16917,N_12571);
or U20984 (N_20984,N_14809,N_14601);
and U20985 (N_20985,N_12331,N_12972);
nor U20986 (N_20986,N_12038,N_14343);
and U20987 (N_20987,N_15754,N_14938);
nand U20988 (N_20988,N_13654,N_12258);
nand U20989 (N_20989,N_15958,N_12186);
or U20990 (N_20990,N_13229,N_15441);
and U20991 (N_20991,N_17940,N_17493);
nand U20992 (N_20992,N_15718,N_15553);
nand U20993 (N_20993,N_17873,N_14449);
and U20994 (N_20994,N_13446,N_15742);
and U20995 (N_20995,N_12190,N_17019);
nor U20996 (N_20996,N_16679,N_14997);
nor U20997 (N_20997,N_12721,N_17592);
or U20998 (N_20998,N_16894,N_12966);
nor U20999 (N_20999,N_17033,N_12648);
or U21000 (N_21000,N_17946,N_13268);
xnor U21001 (N_21001,N_12702,N_17399);
nand U21002 (N_21002,N_12763,N_14842);
nand U21003 (N_21003,N_13217,N_16104);
and U21004 (N_21004,N_17139,N_17743);
and U21005 (N_21005,N_12641,N_13367);
nand U21006 (N_21006,N_17495,N_16157);
nor U21007 (N_21007,N_14409,N_13697);
xnor U21008 (N_21008,N_14851,N_12548);
nor U21009 (N_21009,N_14358,N_14919);
nand U21010 (N_21010,N_12289,N_12306);
xor U21011 (N_21011,N_14974,N_12911);
xor U21012 (N_21012,N_13619,N_13632);
xnor U21013 (N_21013,N_13368,N_16047);
nor U21014 (N_21014,N_17425,N_15556);
nand U21015 (N_21015,N_17241,N_17162);
nand U21016 (N_21016,N_14353,N_16014);
xnor U21017 (N_21017,N_15308,N_16133);
nand U21018 (N_21018,N_13004,N_12348);
and U21019 (N_21019,N_12537,N_17140);
or U21020 (N_21020,N_15710,N_15684);
nand U21021 (N_21021,N_14604,N_16862);
nand U21022 (N_21022,N_12322,N_15617);
nand U21023 (N_21023,N_13251,N_14669);
nor U21024 (N_21024,N_14661,N_12602);
nor U21025 (N_21025,N_17317,N_14561);
xnor U21026 (N_21026,N_12571,N_12074);
nor U21027 (N_21027,N_16917,N_17832);
nor U21028 (N_21028,N_13522,N_13472);
nand U21029 (N_21029,N_15605,N_17217);
xnor U21030 (N_21030,N_13483,N_13214);
or U21031 (N_21031,N_12953,N_15683);
nor U21032 (N_21032,N_15640,N_15528);
xnor U21033 (N_21033,N_17197,N_16391);
nor U21034 (N_21034,N_15902,N_13005);
xnor U21035 (N_21035,N_17057,N_16955);
or U21036 (N_21036,N_17271,N_16375);
xor U21037 (N_21037,N_15657,N_16078);
xor U21038 (N_21038,N_16271,N_17935);
nor U21039 (N_21039,N_15262,N_16893);
nor U21040 (N_21040,N_15800,N_13398);
nand U21041 (N_21041,N_15049,N_16057);
and U21042 (N_21042,N_15021,N_15458);
or U21043 (N_21043,N_13550,N_12493);
nor U21044 (N_21044,N_17767,N_14958);
or U21045 (N_21045,N_15165,N_12239);
nand U21046 (N_21046,N_13907,N_16273);
nor U21047 (N_21047,N_15293,N_13628);
nor U21048 (N_21048,N_16458,N_12766);
or U21049 (N_21049,N_13193,N_12058);
xnor U21050 (N_21050,N_12728,N_12035);
nand U21051 (N_21051,N_12517,N_17858);
or U21052 (N_21052,N_17051,N_15604);
nand U21053 (N_21053,N_17819,N_14394);
or U21054 (N_21054,N_12763,N_15244);
nor U21055 (N_21055,N_13165,N_16574);
or U21056 (N_21056,N_14220,N_12944);
xnor U21057 (N_21057,N_17662,N_13971);
nor U21058 (N_21058,N_12361,N_15008);
nor U21059 (N_21059,N_13160,N_12150);
nor U21060 (N_21060,N_14017,N_12118);
and U21061 (N_21061,N_15335,N_14245);
or U21062 (N_21062,N_16080,N_17583);
xor U21063 (N_21063,N_17234,N_14901);
nor U21064 (N_21064,N_12981,N_14999);
xor U21065 (N_21065,N_17854,N_12092);
and U21066 (N_21066,N_12152,N_14262);
nor U21067 (N_21067,N_15357,N_17392);
nor U21068 (N_21068,N_14469,N_17992);
xnor U21069 (N_21069,N_17078,N_17527);
nand U21070 (N_21070,N_14572,N_15279);
nor U21071 (N_21071,N_13169,N_16231);
and U21072 (N_21072,N_15723,N_15639);
nand U21073 (N_21073,N_14527,N_14366);
or U21074 (N_21074,N_13923,N_15452);
or U21075 (N_21075,N_12604,N_14689);
nand U21076 (N_21076,N_16358,N_16808);
nor U21077 (N_21077,N_17942,N_15533);
or U21078 (N_21078,N_16341,N_17737);
or U21079 (N_21079,N_14659,N_15141);
xnor U21080 (N_21080,N_17963,N_14688);
and U21081 (N_21081,N_15895,N_16916);
xor U21082 (N_21082,N_15038,N_12473);
nor U21083 (N_21083,N_16747,N_13391);
or U21084 (N_21084,N_13227,N_15521);
xor U21085 (N_21085,N_15865,N_12610);
xnor U21086 (N_21086,N_14266,N_16967);
or U21087 (N_21087,N_15987,N_13453);
and U21088 (N_21088,N_17705,N_15615);
nor U21089 (N_21089,N_15350,N_13955);
xor U21090 (N_21090,N_16970,N_15609);
xnor U21091 (N_21091,N_14640,N_15540);
nand U21092 (N_21092,N_16866,N_16327);
xor U21093 (N_21093,N_13118,N_12189);
xor U21094 (N_21094,N_14054,N_14561);
and U21095 (N_21095,N_16824,N_17957);
nand U21096 (N_21096,N_17375,N_17563);
and U21097 (N_21097,N_14343,N_12016);
xnor U21098 (N_21098,N_12821,N_13973);
and U21099 (N_21099,N_12430,N_14145);
nand U21100 (N_21100,N_12088,N_17222);
and U21101 (N_21101,N_16996,N_14140);
and U21102 (N_21102,N_17740,N_17720);
nor U21103 (N_21103,N_15223,N_14996);
and U21104 (N_21104,N_15222,N_16183);
xnor U21105 (N_21105,N_14830,N_15990);
or U21106 (N_21106,N_12464,N_17464);
nand U21107 (N_21107,N_12955,N_17358);
and U21108 (N_21108,N_13312,N_15974);
nor U21109 (N_21109,N_17404,N_16398);
nand U21110 (N_21110,N_17701,N_16627);
nand U21111 (N_21111,N_13930,N_17123);
or U21112 (N_21112,N_12005,N_12890);
nor U21113 (N_21113,N_15118,N_15505);
nand U21114 (N_21114,N_16101,N_16780);
nor U21115 (N_21115,N_17093,N_13555);
nor U21116 (N_21116,N_16951,N_17348);
nand U21117 (N_21117,N_14297,N_17619);
nor U21118 (N_21118,N_12923,N_17542);
nand U21119 (N_21119,N_16271,N_12616);
nand U21120 (N_21120,N_13340,N_17595);
nand U21121 (N_21121,N_14881,N_12329);
xor U21122 (N_21122,N_13970,N_12106);
or U21123 (N_21123,N_15468,N_17465);
and U21124 (N_21124,N_17075,N_13091);
or U21125 (N_21125,N_14374,N_15379);
xor U21126 (N_21126,N_14311,N_15946);
nand U21127 (N_21127,N_12669,N_16409);
xor U21128 (N_21128,N_13184,N_15400);
nor U21129 (N_21129,N_13447,N_16657);
and U21130 (N_21130,N_15044,N_13582);
or U21131 (N_21131,N_16457,N_15147);
nand U21132 (N_21132,N_12144,N_16820);
nor U21133 (N_21133,N_15288,N_15330);
or U21134 (N_21134,N_13879,N_15638);
nand U21135 (N_21135,N_15036,N_15300);
xor U21136 (N_21136,N_15147,N_12328);
and U21137 (N_21137,N_12961,N_16203);
nand U21138 (N_21138,N_15125,N_16421);
xnor U21139 (N_21139,N_15767,N_15772);
or U21140 (N_21140,N_16751,N_14067);
or U21141 (N_21141,N_17770,N_15927);
and U21142 (N_21142,N_13128,N_13022);
or U21143 (N_21143,N_13269,N_13447);
or U21144 (N_21144,N_13176,N_16324);
or U21145 (N_21145,N_12342,N_13505);
or U21146 (N_21146,N_16290,N_13095);
nor U21147 (N_21147,N_14711,N_14202);
or U21148 (N_21148,N_15212,N_13496);
nand U21149 (N_21149,N_12536,N_17358);
and U21150 (N_21150,N_13672,N_15717);
and U21151 (N_21151,N_16318,N_15558);
nor U21152 (N_21152,N_17071,N_16650);
or U21153 (N_21153,N_16955,N_14203);
xnor U21154 (N_21154,N_12728,N_13759);
xnor U21155 (N_21155,N_16144,N_13863);
nor U21156 (N_21156,N_13197,N_13085);
and U21157 (N_21157,N_15665,N_17848);
and U21158 (N_21158,N_13704,N_14070);
or U21159 (N_21159,N_14348,N_13887);
xor U21160 (N_21160,N_15422,N_16498);
nor U21161 (N_21161,N_15218,N_13903);
nand U21162 (N_21162,N_12845,N_15326);
or U21163 (N_21163,N_16894,N_15348);
or U21164 (N_21164,N_15051,N_16419);
xor U21165 (N_21165,N_13135,N_16066);
or U21166 (N_21166,N_12914,N_15290);
xor U21167 (N_21167,N_17096,N_13639);
nor U21168 (N_21168,N_16908,N_15390);
xor U21169 (N_21169,N_13216,N_15690);
nand U21170 (N_21170,N_14009,N_16202);
nor U21171 (N_21171,N_15490,N_16829);
or U21172 (N_21172,N_17425,N_17804);
nand U21173 (N_21173,N_17554,N_12332);
or U21174 (N_21174,N_15979,N_13700);
nor U21175 (N_21175,N_15132,N_14606);
nor U21176 (N_21176,N_16439,N_13985);
or U21177 (N_21177,N_14035,N_15515);
xnor U21178 (N_21178,N_14985,N_12239);
or U21179 (N_21179,N_17562,N_13215);
nor U21180 (N_21180,N_15380,N_13550);
nand U21181 (N_21181,N_15464,N_16467);
nor U21182 (N_21182,N_15023,N_16402);
nand U21183 (N_21183,N_16861,N_13561);
and U21184 (N_21184,N_13472,N_12039);
nand U21185 (N_21185,N_17604,N_12859);
or U21186 (N_21186,N_14408,N_17584);
or U21187 (N_21187,N_15387,N_16102);
nor U21188 (N_21188,N_17866,N_13934);
xnor U21189 (N_21189,N_12950,N_14236);
xnor U21190 (N_21190,N_14008,N_13582);
and U21191 (N_21191,N_17806,N_12384);
nand U21192 (N_21192,N_12911,N_17501);
and U21193 (N_21193,N_16644,N_15580);
and U21194 (N_21194,N_14837,N_14996);
nand U21195 (N_21195,N_15203,N_14214);
xor U21196 (N_21196,N_14364,N_14218);
or U21197 (N_21197,N_14020,N_15578);
or U21198 (N_21198,N_13573,N_14805);
nand U21199 (N_21199,N_16067,N_14545);
and U21200 (N_21200,N_14982,N_17309);
xnor U21201 (N_21201,N_12822,N_14916);
nor U21202 (N_21202,N_17751,N_14957);
xor U21203 (N_21203,N_15367,N_17399);
and U21204 (N_21204,N_14399,N_14279);
xor U21205 (N_21205,N_17581,N_17670);
xnor U21206 (N_21206,N_12778,N_15826);
and U21207 (N_21207,N_14158,N_13548);
and U21208 (N_21208,N_17821,N_17710);
or U21209 (N_21209,N_12775,N_16596);
or U21210 (N_21210,N_15091,N_15985);
or U21211 (N_21211,N_12559,N_17209);
nor U21212 (N_21212,N_16605,N_14053);
nor U21213 (N_21213,N_14061,N_16426);
xor U21214 (N_21214,N_13337,N_12311);
xnor U21215 (N_21215,N_13719,N_17299);
and U21216 (N_21216,N_13369,N_14766);
nand U21217 (N_21217,N_15588,N_17908);
nand U21218 (N_21218,N_12074,N_16062);
and U21219 (N_21219,N_16706,N_17987);
nor U21220 (N_21220,N_17286,N_13537);
xor U21221 (N_21221,N_15092,N_13833);
nand U21222 (N_21222,N_12691,N_13321);
nor U21223 (N_21223,N_16101,N_14616);
and U21224 (N_21224,N_15517,N_12319);
and U21225 (N_21225,N_16231,N_17428);
nand U21226 (N_21226,N_12198,N_17942);
and U21227 (N_21227,N_17342,N_15855);
nor U21228 (N_21228,N_14520,N_14762);
nor U21229 (N_21229,N_12650,N_17842);
or U21230 (N_21230,N_15826,N_13398);
nand U21231 (N_21231,N_16751,N_17818);
or U21232 (N_21232,N_14273,N_17904);
nor U21233 (N_21233,N_16658,N_17612);
or U21234 (N_21234,N_17150,N_14091);
nand U21235 (N_21235,N_15059,N_14145);
xnor U21236 (N_21236,N_13395,N_16360);
xor U21237 (N_21237,N_16524,N_13137);
and U21238 (N_21238,N_12098,N_15289);
or U21239 (N_21239,N_15513,N_15711);
nor U21240 (N_21240,N_14685,N_12378);
xnor U21241 (N_21241,N_15225,N_15031);
or U21242 (N_21242,N_15858,N_12340);
or U21243 (N_21243,N_13985,N_13340);
or U21244 (N_21244,N_15643,N_17699);
nand U21245 (N_21245,N_14730,N_16393);
xnor U21246 (N_21246,N_14180,N_13069);
or U21247 (N_21247,N_15776,N_12118);
nor U21248 (N_21248,N_13686,N_13320);
nor U21249 (N_21249,N_16873,N_13771);
nand U21250 (N_21250,N_15037,N_17942);
nand U21251 (N_21251,N_14363,N_17750);
nand U21252 (N_21252,N_13905,N_15123);
and U21253 (N_21253,N_15075,N_15148);
nor U21254 (N_21254,N_13059,N_16352);
and U21255 (N_21255,N_16154,N_15254);
and U21256 (N_21256,N_14238,N_13384);
or U21257 (N_21257,N_15150,N_15700);
and U21258 (N_21258,N_16092,N_16681);
nand U21259 (N_21259,N_16717,N_15180);
nand U21260 (N_21260,N_13758,N_14237);
nor U21261 (N_21261,N_12735,N_17308);
or U21262 (N_21262,N_12111,N_13028);
xnor U21263 (N_21263,N_13673,N_17654);
or U21264 (N_21264,N_14021,N_17822);
or U21265 (N_21265,N_13971,N_14636);
nand U21266 (N_21266,N_17458,N_14178);
nand U21267 (N_21267,N_14599,N_17722);
and U21268 (N_21268,N_13473,N_15138);
xnor U21269 (N_21269,N_15943,N_17830);
and U21270 (N_21270,N_16072,N_14995);
nand U21271 (N_21271,N_17136,N_14958);
nor U21272 (N_21272,N_13854,N_12633);
nor U21273 (N_21273,N_15715,N_13225);
and U21274 (N_21274,N_17430,N_13957);
or U21275 (N_21275,N_17090,N_17059);
or U21276 (N_21276,N_12726,N_12444);
or U21277 (N_21277,N_15953,N_14823);
xor U21278 (N_21278,N_12455,N_17210);
and U21279 (N_21279,N_14387,N_16309);
or U21280 (N_21280,N_17844,N_12015);
nand U21281 (N_21281,N_12437,N_14917);
nand U21282 (N_21282,N_14228,N_14887);
nand U21283 (N_21283,N_17655,N_15509);
or U21284 (N_21284,N_14757,N_15364);
nor U21285 (N_21285,N_17699,N_16001);
or U21286 (N_21286,N_13960,N_17978);
nor U21287 (N_21287,N_12559,N_16942);
nand U21288 (N_21288,N_14074,N_15525);
xor U21289 (N_21289,N_16160,N_15290);
or U21290 (N_21290,N_12226,N_17735);
xnor U21291 (N_21291,N_12589,N_12683);
nor U21292 (N_21292,N_12263,N_13012);
nand U21293 (N_21293,N_13566,N_15331);
and U21294 (N_21294,N_14495,N_16834);
and U21295 (N_21295,N_14289,N_15536);
and U21296 (N_21296,N_17070,N_14049);
nand U21297 (N_21297,N_12146,N_17915);
and U21298 (N_21298,N_15371,N_12327);
nor U21299 (N_21299,N_14833,N_15001);
or U21300 (N_21300,N_17438,N_13754);
or U21301 (N_21301,N_12116,N_13769);
or U21302 (N_21302,N_17304,N_15745);
nor U21303 (N_21303,N_17160,N_17860);
nand U21304 (N_21304,N_16154,N_16954);
nor U21305 (N_21305,N_14661,N_13225);
or U21306 (N_21306,N_12446,N_17176);
xor U21307 (N_21307,N_17985,N_15640);
nand U21308 (N_21308,N_12543,N_17312);
nand U21309 (N_21309,N_17468,N_12501);
xor U21310 (N_21310,N_14538,N_16203);
and U21311 (N_21311,N_13151,N_14082);
nand U21312 (N_21312,N_16650,N_14872);
xnor U21313 (N_21313,N_15367,N_14634);
or U21314 (N_21314,N_13397,N_15457);
or U21315 (N_21315,N_14734,N_16963);
nand U21316 (N_21316,N_15918,N_16976);
or U21317 (N_21317,N_14017,N_12860);
and U21318 (N_21318,N_13567,N_14553);
nand U21319 (N_21319,N_17202,N_15251);
and U21320 (N_21320,N_15495,N_15250);
or U21321 (N_21321,N_14778,N_12157);
or U21322 (N_21322,N_13464,N_12449);
xnor U21323 (N_21323,N_13073,N_16780);
nand U21324 (N_21324,N_17450,N_14612);
or U21325 (N_21325,N_15542,N_15457);
and U21326 (N_21326,N_14200,N_15168);
and U21327 (N_21327,N_15283,N_17125);
nor U21328 (N_21328,N_16844,N_16640);
and U21329 (N_21329,N_14742,N_16736);
nand U21330 (N_21330,N_16126,N_16835);
xnor U21331 (N_21331,N_13086,N_17255);
and U21332 (N_21332,N_16689,N_12925);
and U21333 (N_21333,N_12788,N_14746);
xor U21334 (N_21334,N_13619,N_12236);
nand U21335 (N_21335,N_17791,N_13608);
xor U21336 (N_21336,N_17030,N_16296);
nand U21337 (N_21337,N_17550,N_15159);
and U21338 (N_21338,N_17188,N_12292);
or U21339 (N_21339,N_14888,N_15599);
and U21340 (N_21340,N_16178,N_13117);
or U21341 (N_21341,N_16936,N_17225);
nand U21342 (N_21342,N_14220,N_17257);
xor U21343 (N_21343,N_13486,N_12478);
or U21344 (N_21344,N_14143,N_14696);
or U21345 (N_21345,N_17260,N_17261);
nor U21346 (N_21346,N_14376,N_16998);
or U21347 (N_21347,N_13850,N_13594);
and U21348 (N_21348,N_17881,N_13388);
or U21349 (N_21349,N_15210,N_16062);
nand U21350 (N_21350,N_17064,N_16098);
nand U21351 (N_21351,N_15228,N_12295);
or U21352 (N_21352,N_17590,N_16202);
xnor U21353 (N_21353,N_13296,N_13970);
nand U21354 (N_21354,N_15711,N_16465);
nor U21355 (N_21355,N_13229,N_17203);
xnor U21356 (N_21356,N_17141,N_14410);
xnor U21357 (N_21357,N_15162,N_13557);
nor U21358 (N_21358,N_16243,N_15758);
nor U21359 (N_21359,N_12129,N_17566);
xor U21360 (N_21360,N_13337,N_13030);
or U21361 (N_21361,N_12247,N_14962);
and U21362 (N_21362,N_17025,N_12919);
xor U21363 (N_21363,N_17392,N_17377);
nor U21364 (N_21364,N_17050,N_14240);
xnor U21365 (N_21365,N_13039,N_15933);
or U21366 (N_21366,N_13689,N_14153);
nor U21367 (N_21367,N_15293,N_12500);
nand U21368 (N_21368,N_12380,N_14097);
nor U21369 (N_21369,N_13975,N_14860);
or U21370 (N_21370,N_13975,N_15537);
nor U21371 (N_21371,N_13983,N_14760);
and U21372 (N_21372,N_17177,N_15993);
and U21373 (N_21373,N_14968,N_14048);
or U21374 (N_21374,N_12415,N_16044);
nand U21375 (N_21375,N_16509,N_16565);
and U21376 (N_21376,N_14946,N_15669);
and U21377 (N_21377,N_16213,N_16156);
and U21378 (N_21378,N_15395,N_17593);
nand U21379 (N_21379,N_12588,N_14262);
nand U21380 (N_21380,N_15805,N_15232);
and U21381 (N_21381,N_17610,N_12299);
nand U21382 (N_21382,N_17639,N_14795);
nor U21383 (N_21383,N_14620,N_14021);
and U21384 (N_21384,N_15970,N_16265);
nand U21385 (N_21385,N_12760,N_16240);
xnor U21386 (N_21386,N_14270,N_12449);
nand U21387 (N_21387,N_15107,N_15417);
and U21388 (N_21388,N_12581,N_13701);
or U21389 (N_21389,N_15898,N_12603);
and U21390 (N_21390,N_13484,N_17707);
xor U21391 (N_21391,N_16278,N_14198);
nor U21392 (N_21392,N_17433,N_16286);
xnor U21393 (N_21393,N_13562,N_16951);
or U21394 (N_21394,N_17597,N_12959);
and U21395 (N_21395,N_14797,N_14599);
nand U21396 (N_21396,N_17226,N_12616);
and U21397 (N_21397,N_15526,N_15586);
nand U21398 (N_21398,N_13401,N_17179);
xor U21399 (N_21399,N_15622,N_12456);
xnor U21400 (N_21400,N_14417,N_17880);
nand U21401 (N_21401,N_15966,N_14023);
nand U21402 (N_21402,N_12574,N_15080);
or U21403 (N_21403,N_12205,N_12395);
or U21404 (N_21404,N_16484,N_14282);
nand U21405 (N_21405,N_15924,N_14675);
or U21406 (N_21406,N_17480,N_12973);
or U21407 (N_21407,N_12396,N_17269);
and U21408 (N_21408,N_16798,N_14995);
nor U21409 (N_21409,N_17875,N_12686);
nor U21410 (N_21410,N_15854,N_14303);
nand U21411 (N_21411,N_12588,N_13733);
or U21412 (N_21412,N_17559,N_16025);
or U21413 (N_21413,N_17390,N_13493);
or U21414 (N_21414,N_12726,N_16608);
nor U21415 (N_21415,N_14085,N_15471);
xnor U21416 (N_21416,N_13693,N_15422);
nand U21417 (N_21417,N_14787,N_13999);
xor U21418 (N_21418,N_16454,N_16215);
or U21419 (N_21419,N_15738,N_12420);
nor U21420 (N_21420,N_17339,N_13240);
and U21421 (N_21421,N_17049,N_16616);
xor U21422 (N_21422,N_17737,N_14167);
and U21423 (N_21423,N_17978,N_12872);
or U21424 (N_21424,N_13266,N_15038);
xnor U21425 (N_21425,N_13413,N_14176);
nand U21426 (N_21426,N_12142,N_12143);
and U21427 (N_21427,N_13954,N_17956);
and U21428 (N_21428,N_13404,N_16760);
and U21429 (N_21429,N_14107,N_17816);
or U21430 (N_21430,N_14132,N_13239);
xnor U21431 (N_21431,N_15863,N_13077);
nor U21432 (N_21432,N_14044,N_13599);
xnor U21433 (N_21433,N_17863,N_17699);
nor U21434 (N_21434,N_12480,N_15613);
nor U21435 (N_21435,N_12788,N_17970);
and U21436 (N_21436,N_12154,N_13836);
xor U21437 (N_21437,N_12540,N_17818);
and U21438 (N_21438,N_12903,N_12771);
or U21439 (N_21439,N_16029,N_14660);
nor U21440 (N_21440,N_15389,N_14750);
or U21441 (N_21441,N_15715,N_17480);
xor U21442 (N_21442,N_12431,N_17750);
and U21443 (N_21443,N_17551,N_13836);
and U21444 (N_21444,N_12734,N_12728);
xor U21445 (N_21445,N_15511,N_16978);
nand U21446 (N_21446,N_16302,N_14840);
or U21447 (N_21447,N_17033,N_14711);
xnor U21448 (N_21448,N_17737,N_13481);
or U21449 (N_21449,N_13523,N_12942);
or U21450 (N_21450,N_14573,N_14563);
xnor U21451 (N_21451,N_16047,N_14738);
nor U21452 (N_21452,N_15360,N_12392);
nand U21453 (N_21453,N_16848,N_17939);
nand U21454 (N_21454,N_12498,N_16354);
nand U21455 (N_21455,N_16630,N_15925);
or U21456 (N_21456,N_12198,N_12361);
or U21457 (N_21457,N_12647,N_14642);
and U21458 (N_21458,N_12834,N_12523);
and U21459 (N_21459,N_12603,N_17160);
nand U21460 (N_21460,N_14682,N_15522);
nor U21461 (N_21461,N_12358,N_13313);
and U21462 (N_21462,N_14371,N_17074);
or U21463 (N_21463,N_12965,N_17135);
or U21464 (N_21464,N_15042,N_15909);
and U21465 (N_21465,N_17453,N_16908);
or U21466 (N_21466,N_17755,N_12375);
and U21467 (N_21467,N_15851,N_13646);
and U21468 (N_21468,N_15310,N_14939);
nand U21469 (N_21469,N_16452,N_13954);
nand U21470 (N_21470,N_15013,N_16405);
nand U21471 (N_21471,N_14454,N_14981);
nand U21472 (N_21472,N_13204,N_15356);
or U21473 (N_21473,N_13585,N_12476);
nor U21474 (N_21474,N_13759,N_16290);
xnor U21475 (N_21475,N_15412,N_14970);
and U21476 (N_21476,N_13139,N_15891);
or U21477 (N_21477,N_13281,N_14950);
nand U21478 (N_21478,N_13234,N_16850);
nand U21479 (N_21479,N_14845,N_17687);
nand U21480 (N_21480,N_17317,N_12768);
nor U21481 (N_21481,N_16835,N_12505);
or U21482 (N_21482,N_14720,N_17710);
nor U21483 (N_21483,N_15931,N_16778);
nor U21484 (N_21484,N_14557,N_15807);
xnor U21485 (N_21485,N_12591,N_17402);
nand U21486 (N_21486,N_13471,N_13622);
and U21487 (N_21487,N_15895,N_13013);
nand U21488 (N_21488,N_16708,N_17146);
or U21489 (N_21489,N_16661,N_12520);
and U21490 (N_21490,N_14407,N_16168);
and U21491 (N_21491,N_15024,N_12670);
nor U21492 (N_21492,N_15937,N_17904);
and U21493 (N_21493,N_12379,N_14436);
and U21494 (N_21494,N_12356,N_13634);
nand U21495 (N_21495,N_17724,N_17310);
nand U21496 (N_21496,N_17888,N_15634);
or U21497 (N_21497,N_16981,N_17175);
nand U21498 (N_21498,N_14938,N_13816);
and U21499 (N_21499,N_17695,N_14463);
or U21500 (N_21500,N_15509,N_17792);
xnor U21501 (N_21501,N_12068,N_13981);
nor U21502 (N_21502,N_13913,N_14636);
xnor U21503 (N_21503,N_16057,N_12819);
nor U21504 (N_21504,N_16285,N_16620);
or U21505 (N_21505,N_15355,N_17149);
xnor U21506 (N_21506,N_14059,N_17036);
nand U21507 (N_21507,N_12120,N_15229);
or U21508 (N_21508,N_13768,N_16363);
or U21509 (N_21509,N_16804,N_14830);
and U21510 (N_21510,N_17610,N_14507);
or U21511 (N_21511,N_14259,N_15225);
and U21512 (N_21512,N_14563,N_12042);
xor U21513 (N_21513,N_14591,N_15793);
nor U21514 (N_21514,N_14173,N_13641);
or U21515 (N_21515,N_17518,N_12649);
xnor U21516 (N_21516,N_15259,N_15942);
or U21517 (N_21517,N_12708,N_14280);
nand U21518 (N_21518,N_16516,N_16471);
nand U21519 (N_21519,N_15102,N_15034);
or U21520 (N_21520,N_14846,N_14449);
nand U21521 (N_21521,N_14932,N_17093);
xor U21522 (N_21522,N_16800,N_16872);
xnor U21523 (N_21523,N_15499,N_12609);
nand U21524 (N_21524,N_12788,N_16446);
or U21525 (N_21525,N_12122,N_14950);
nor U21526 (N_21526,N_13965,N_17224);
and U21527 (N_21527,N_16217,N_15272);
nor U21528 (N_21528,N_14475,N_15207);
nand U21529 (N_21529,N_15856,N_13784);
xor U21530 (N_21530,N_12718,N_17296);
or U21531 (N_21531,N_14966,N_12957);
and U21532 (N_21532,N_17368,N_16866);
or U21533 (N_21533,N_12569,N_13293);
or U21534 (N_21534,N_12485,N_17920);
nor U21535 (N_21535,N_17190,N_17420);
nand U21536 (N_21536,N_17400,N_15941);
xnor U21537 (N_21537,N_17097,N_17483);
nand U21538 (N_21538,N_12928,N_14038);
or U21539 (N_21539,N_13966,N_12924);
and U21540 (N_21540,N_12234,N_14309);
nand U21541 (N_21541,N_14118,N_17249);
xor U21542 (N_21542,N_16250,N_12178);
or U21543 (N_21543,N_17341,N_16955);
nor U21544 (N_21544,N_14206,N_17159);
xnor U21545 (N_21545,N_16046,N_17525);
nand U21546 (N_21546,N_15057,N_17541);
xor U21547 (N_21547,N_13850,N_14423);
nand U21548 (N_21548,N_12441,N_17321);
nor U21549 (N_21549,N_15328,N_12191);
xor U21550 (N_21550,N_14274,N_14710);
and U21551 (N_21551,N_13560,N_12184);
and U21552 (N_21552,N_12336,N_16325);
xor U21553 (N_21553,N_15587,N_12853);
xor U21554 (N_21554,N_14635,N_16336);
or U21555 (N_21555,N_17645,N_13277);
nand U21556 (N_21556,N_13027,N_13867);
or U21557 (N_21557,N_12140,N_16080);
nor U21558 (N_21558,N_16406,N_17426);
and U21559 (N_21559,N_14147,N_16161);
nor U21560 (N_21560,N_17428,N_13221);
xnor U21561 (N_21561,N_14261,N_16263);
xnor U21562 (N_21562,N_17803,N_13795);
xor U21563 (N_21563,N_13319,N_13331);
or U21564 (N_21564,N_16362,N_15206);
nand U21565 (N_21565,N_17752,N_14441);
or U21566 (N_21566,N_16591,N_16022);
or U21567 (N_21567,N_14543,N_17115);
or U21568 (N_21568,N_14574,N_17080);
xnor U21569 (N_21569,N_13529,N_16450);
nor U21570 (N_21570,N_15379,N_16109);
and U21571 (N_21571,N_14798,N_12154);
or U21572 (N_21572,N_14447,N_14673);
nand U21573 (N_21573,N_13640,N_17433);
or U21574 (N_21574,N_12377,N_15139);
nand U21575 (N_21575,N_16222,N_15882);
xnor U21576 (N_21576,N_13606,N_17529);
or U21577 (N_21577,N_16803,N_15744);
nor U21578 (N_21578,N_17515,N_12603);
or U21579 (N_21579,N_14324,N_14363);
or U21580 (N_21580,N_12236,N_15517);
nand U21581 (N_21581,N_17300,N_12713);
nor U21582 (N_21582,N_16987,N_12543);
xnor U21583 (N_21583,N_13994,N_16552);
xor U21584 (N_21584,N_13067,N_14751);
or U21585 (N_21585,N_13662,N_13162);
nor U21586 (N_21586,N_16771,N_17701);
xor U21587 (N_21587,N_14189,N_12192);
and U21588 (N_21588,N_12255,N_16865);
xor U21589 (N_21589,N_17487,N_12006);
or U21590 (N_21590,N_14873,N_17438);
nand U21591 (N_21591,N_15244,N_14029);
and U21592 (N_21592,N_13549,N_16863);
and U21593 (N_21593,N_12319,N_15083);
nand U21594 (N_21594,N_16334,N_12457);
nand U21595 (N_21595,N_13464,N_12388);
nor U21596 (N_21596,N_12626,N_15809);
and U21597 (N_21597,N_12903,N_15153);
and U21598 (N_21598,N_15919,N_17176);
or U21599 (N_21599,N_15838,N_13436);
nand U21600 (N_21600,N_14986,N_17163);
xnor U21601 (N_21601,N_14412,N_17800);
and U21602 (N_21602,N_15825,N_15353);
or U21603 (N_21603,N_16014,N_17866);
xnor U21604 (N_21604,N_13539,N_15504);
or U21605 (N_21605,N_15806,N_15631);
xnor U21606 (N_21606,N_13647,N_13033);
or U21607 (N_21607,N_16126,N_14559);
nor U21608 (N_21608,N_12884,N_15549);
xor U21609 (N_21609,N_17356,N_15350);
or U21610 (N_21610,N_13358,N_13395);
and U21611 (N_21611,N_15954,N_15743);
nor U21612 (N_21612,N_14104,N_12329);
nor U21613 (N_21613,N_15023,N_14661);
xor U21614 (N_21614,N_13466,N_15698);
and U21615 (N_21615,N_12377,N_16333);
and U21616 (N_21616,N_13792,N_12945);
and U21617 (N_21617,N_12842,N_14976);
xor U21618 (N_21618,N_13216,N_14754);
and U21619 (N_21619,N_14085,N_16191);
nor U21620 (N_21620,N_14142,N_15722);
xnor U21621 (N_21621,N_14522,N_16979);
nand U21622 (N_21622,N_13513,N_12378);
nand U21623 (N_21623,N_17633,N_13548);
nand U21624 (N_21624,N_16351,N_14829);
and U21625 (N_21625,N_17608,N_14656);
nand U21626 (N_21626,N_16234,N_12549);
or U21627 (N_21627,N_13714,N_12784);
and U21628 (N_21628,N_15803,N_12815);
and U21629 (N_21629,N_13654,N_12157);
nand U21630 (N_21630,N_15703,N_13895);
xor U21631 (N_21631,N_17803,N_12857);
or U21632 (N_21632,N_14529,N_15946);
nor U21633 (N_21633,N_16653,N_15889);
nand U21634 (N_21634,N_13407,N_13910);
or U21635 (N_21635,N_15327,N_16813);
nor U21636 (N_21636,N_15144,N_12686);
nand U21637 (N_21637,N_13462,N_13745);
nor U21638 (N_21638,N_15061,N_13052);
nand U21639 (N_21639,N_14805,N_16560);
and U21640 (N_21640,N_14613,N_13476);
nand U21641 (N_21641,N_12055,N_16769);
and U21642 (N_21642,N_16580,N_17363);
nor U21643 (N_21643,N_17205,N_12937);
nor U21644 (N_21644,N_13450,N_16997);
or U21645 (N_21645,N_12606,N_15703);
nand U21646 (N_21646,N_16510,N_15768);
nor U21647 (N_21647,N_12758,N_15145);
and U21648 (N_21648,N_12379,N_15645);
nor U21649 (N_21649,N_12623,N_14109);
nand U21650 (N_21650,N_12113,N_17000);
xnor U21651 (N_21651,N_14474,N_17801);
xor U21652 (N_21652,N_13963,N_17033);
or U21653 (N_21653,N_16189,N_16370);
xor U21654 (N_21654,N_15281,N_13290);
nor U21655 (N_21655,N_14143,N_16154);
or U21656 (N_21656,N_13353,N_14776);
nand U21657 (N_21657,N_14374,N_12207);
or U21658 (N_21658,N_12952,N_12217);
and U21659 (N_21659,N_15086,N_17504);
or U21660 (N_21660,N_12364,N_17412);
nor U21661 (N_21661,N_14444,N_12909);
nor U21662 (N_21662,N_13194,N_13211);
xor U21663 (N_21663,N_13907,N_13723);
or U21664 (N_21664,N_12821,N_12877);
nor U21665 (N_21665,N_12429,N_13760);
and U21666 (N_21666,N_13379,N_15414);
xor U21667 (N_21667,N_15190,N_16313);
xor U21668 (N_21668,N_14618,N_17677);
xnor U21669 (N_21669,N_13328,N_13253);
and U21670 (N_21670,N_15105,N_14266);
nand U21671 (N_21671,N_15101,N_16682);
xor U21672 (N_21672,N_14228,N_14928);
or U21673 (N_21673,N_15989,N_12901);
nand U21674 (N_21674,N_12104,N_17100);
nor U21675 (N_21675,N_16127,N_14292);
nand U21676 (N_21676,N_12550,N_14030);
or U21677 (N_21677,N_17951,N_14743);
and U21678 (N_21678,N_12007,N_14755);
or U21679 (N_21679,N_14020,N_15533);
or U21680 (N_21680,N_14775,N_13738);
and U21681 (N_21681,N_16114,N_16066);
nor U21682 (N_21682,N_17453,N_15027);
and U21683 (N_21683,N_15359,N_13336);
or U21684 (N_21684,N_14926,N_14843);
and U21685 (N_21685,N_17915,N_12247);
and U21686 (N_21686,N_12914,N_12409);
xor U21687 (N_21687,N_16962,N_16485);
nand U21688 (N_21688,N_14173,N_16976);
xnor U21689 (N_21689,N_14430,N_16812);
or U21690 (N_21690,N_15937,N_14761);
nor U21691 (N_21691,N_15554,N_12729);
or U21692 (N_21692,N_14563,N_15593);
or U21693 (N_21693,N_13740,N_17029);
and U21694 (N_21694,N_13564,N_13315);
nor U21695 (N_21695,N_17337,N_16153);
and U21696 (N_21696,N_16432,N_15030);
nor U21697 (N_21697,N_12361,N_14189);
or U21698 (N_21698,N_17486,N_16672);
nor U21699 (N_21699,N_15421,N_12806);
and U21700 (N_21700,N_14462,N_15643);
xnor U21701 (N_21701,N_15414,N_13685);
xnor U21702 (N_21702,N_16368,N_15309);
or U21703 (N_21703,N_13553,N_15225);
or U21704 (N_21704,N_16910,N_13038);
nand U21705 (N_21705,N_17273,N_15436);
or U21706 (N_21706,N_12424,N_14815);
nor U21707 (N_21707,N_16108,N_15692);
xor U21708 (N_21708,N_17311,N_12849);
and U21709 (N_21709,N_14738,N_12766);
xor U21710 (N_21710,N_17640,N_16499);
and U21711 (N_21711,N_14634,N_15691);
and U21712 (N_21712,N_15787,N_14096);
nor U21713 (N_21713,N_16855,N_17677);
nand U21714 (N_21714,N_13810,N_13833);
xnor U21715 (N_21715,N_13504,N_17838);
nand U21716 (N_21716,N_12180,N_14128);
xor U21717 (N_21717,N_17033,N_15139);
or U21718 (N_21718,N_15348,N_15018);
xor U21719 (N_21719,N_17110,N_17172);
xnor U21720 (N_21720,N_13409,N_15483);
and U21721 (N_21721,N_13684,N_14961);
xor U21722 (N_21722,N_14823,N_12259);
nand U21723 (N_21723,N_17534,N_14098);
nor U21724 (N_21724,N_14194,N_17333);
and U21725 (N_21725,N_14475,N_14812);
or U21726 (N_21726,N_13883,N_13942);
xnor U21727 (N_21727,N_14696,N_12812);
and U21728 (N_21728,N_12978,N_12564);
xor U21729 (N_21729,N_12360,N_12895);
and U21730 (N_21730,N_13359,N_17672);
nand U21731 (N_21731,N_14843,N_14110);
nor U21732 (N_21732,N_16599,N_17173);
nand U21733 (N_21733,N_17945,N_12449);
and U21734 (N_21734,N_16064,N_14188);
nor U21735 (N_21735,N_12852,N_15229);
nor U21736 (N_21736,N_17535,N_14185);
or U21737 (N_21737,N_14028,N_13703);
and U21738 (N_21738,N_17852,N_16456);
or U21739 (N_21739,N_16521,N_13930);
and U21740 (N_21740,N_15943,N_14279);
or U21741 (N_21741,N_12442,N_14834);
or U21742 (N_21742,N_16392,N_17268);
nor U21743 (N_21743,N_17699,N_13194);
nor U21744 (N_21744,N_13614,N_17714);
and U21745 (N_21745,N_17382,N_17212);
xnor U21746 (N_21746,N_16877,N_12994);
or U21747 (N_21747,N_16580,N_15146);
or U21748 (N_21748,N_17210,N_14220);
nor U21749 (N_21749,N_12099,N_12485);
or U21750 (N_21750,N_13655,N_12856);
nor U21751 (N_21751,N_13511,N_13115);
nor U21752 (N_21752,N_16204,N_16740);
xor U21753 (N_21753,N_13692,N_16616);
nand U21754 (N_21754,N_16970,N_15068);
nor U21755 (N_21755,N_17484,N_17078);
or U21756 (N_21756,N_13731,N_13978);
or U21757 (N_21757,N_15426,N_13143);
or U21758 (N_21758,N_13298,N_15627);
nor U21759 (N_21759,N_16460,N_12179);
nor U21760 (N_21760,N_17116,N_17496);
xor U21761 (N_21761,N_17141,N_16571);
nor U21762 (N_21762,N_12036,N_13232);
xnor U21763 (N_21763,N_16560,N_12343);
nor U21764 (N_21764,N_17421,N_16320);
nand U21765 (N_21765,N_14326,N_16841);
xnor U21766 (N_21766,N_13153,N_14682);
nor U21767 (N_21767,N_13825,N_14026);
or U21768 (N_21768,N_17805,N_15158);
and U21769 (N_21769,N_17984,N_13575);
nand U21770 (N_21770,N_15267,N_12228);
or U21771 (N_21771,N_14943,N_14463);
xnor U21772 (N_21772,N_12421,N_15906);
xnor U21773 (N_21773,N_16389,N_15265);
nor U21774 (N_21774,N_13121,N_14539);
and U21775 (N_21775,N_17641,N_15148);
nor U21776 (N_21776,N_16175,N_15446);
nor U21777 (N_21777,N_12188,N_16570);
nor U21778 (N_21778,N_15585,N_14351);
or U21779 (N_21779,N_14722,N_14500);
nor U21780 (N_21780,N_13861,N_17697);
nand U21781 (N_21781,N_12733,N_15714);
nor U21782 (N_21782,N_17690,N_13450);
and U21783 (N_21783,N_12708,N_12391);
nor U21784 (N_21784,N_12651,N_16873);
and U21785 (N_21785,N_16376,N_14708);
and U21786 (N_21786,N_16144,N_14572);
and U21787 (N_21787,N_13934,N_17666);
or U21788 (N_21788,N_12503,N_12716);
nor U21789 (N_21789,N_15897,N_15659);
xnor U21790 (N_21790,N_12734,N_16125);
nand U21791 (N_21791,N_15759,N_15127);
nor U21792 (N_21792,N_15593,N_15538);
or U21793 (N_21793,N_17297,N_14830);
xor U21794 (N_21794,N_15496,N_17742);
nor U21795 (N_21795,N_16234,N_16152);
nand U21796 (N_21796,N_15073,N_13281);
or U21797 (N_21797,N_13445,N_14389);
and U21798 (N_21798,N_16938,N_12354);
and U21799 (N_21799,N_12795,N_14426);
or U21800 (N_21800,N_13208,N_16787);
or U21801 (N_21801,N_15548,N_16718);
xnor U21802 (N_21802,N_16077,N_14629);
nand U21803 (N_21803,N_14173,N_14829);
nand U21804 (N_21804,N_12056,N_13010);
xor U21805 (N_21805,N_12874,N_12512);
and U21806 (N_21806,N_12217,N_12123);
and U21807 (N_21807,N_14400,N_12582);
nor U21808 (N_21808,N_12633,N_14689);
and U21809 (N_21809,N_13291,N_12687);
or U21810 (N_21810,N_13237,N_12455);
or U21811 (N_21811,N_16839,N_13608);
nor U21812 (N_21812,N_15606,N_16058);
or U21813 (N_21813,N_14961,N_14200);
nor U21814 (N_21814,N_15493,N_14176);
nand U21815 (N_21815,N_13291,N_17064);
nand U21816 (N_21816,N_17400,N_12568);
and U21817 (N_21817,N_12694,N_16000);
nand U21818 (N_21818,N_14122,N_15184);
or U21819 (N_21819,N_17226,N_12015);
xor U21820 (N_21820,N_13291,N_13368);
nand U21821 (N_21821,N_17144,N_16973);
or U21822 (N_21822,N_13143,N_16117);
xor U21823 (N_21823,N_16504,N_16508);
and U21824 (N_21824,N_17456,N_12996);
or U21825 (N_21825,N_14462,N_13623);
nor U21826 (N_21826,N_17167,N_14990);
nand U21827 (N_21827,N_17619,N_14849);
xnor U21828 (N_21828,N_15789,N_17283);
nand U21829 (N_21829,N_14549,N_14576);
or U21830 (N_21830,N_13322,N_16547);
nor U21831 (N_21831,N_14267,N_13884);
xor U21832 (N_21832,N_14582,N_17170);
nand U21833 (N_21833,N_16878,N_14278);
nand U21834 (N_21834,N_17025,N_12811);
xor U21835 (N_21835,N_15173,N_13375);
and U21836 (N_21836,N_14555,N_15027);
nor U21837 (N_21837,N_14882,N_15776);
xor U21838 (N_21838,N_12258,N_16878);
nor U21839 (N_21839,N_17307,N_17536);
and U21840 (N_21840,N_12404,N_15290);
nand U21841 (N_21841,N_12076,N_13692);
nand U21842 (N_21842,N_14047,N_17669);
nand U21843 (N_21843,N_16493,N_14190);
and U21844 (N_21844,N_17300,N_16017);
and U21845 (N_21845,N_16892,N_16519);
and U21846 (N_21846,N_16067,N_12270);
nor U21847 (N_21847,N_17058,N_16582);
xnor U21848 (N_21848,N_14125,N_12629);
nand U21849 (N_21849,N_15638,N_15555);
nand U21850 (N_21850,N_15919,N_12298);
and U21851 (N_21851,N_12103,N_17618);
or U21852 (N_21852,N_15504,N_14475);
nor U21853 (N_21853,N_12319,N_16322);
and U21854 (N_21854,N_15724,N_15400);
nor U21855 (N_21855,N_15061,N_14627);
and U21856 (N_21856,N_12180,N_13407);
and U21857 (N_21857,N_13366,N_14911);
nor U21858 (N_21858,N_15220,N_13503);
nor U21859 (N_21859,N_14710,N_17194);
nand U21860 (N_21860,N_16888,N_13128);
and U21861 (N_21861,N_13965,N_14288);
nor U21862 (N_21862,N_13138,N_15003);
and U21863 (N_21863,N_13528,N_13960);
or U21864 (N_21864,N_12319,N_12314);
or U21865 (N_21865,N_12417,N_13891);
xor U21866 (N_21866,N_13481,N_17127);
nor U21867 (N_21867,N_12085,N_13803);
nor U21868 (N_21868,N_12417,N_14549);
nand U21869 (N_21869,N_12272,N_16431);
or U21870 (N_21870,N_13377,N_15556);
nand U21871 (N_21871,N_17909,N_17401);
or U21872 (N_21872,N_17182,N_15220);
xnor U21873 (N_21873,N_15600,N_12127);
nor U21874 (N_21874,N_16103,N_15272);
nor U21875 (N_21875,N_15060,N_17824);
nor U21876 (N_21876,N_15013,N_15422);
and U21877 (N_21877,N_14745,N_13584);
and U21878 (N_21878,N_17052,N_16228);
xor U21879 (N_21879,N_12765,N_12301);
xor U21880 (N_21880,N_14574,N_16330);
and U21881 (N_21881,N_17004,N_14346);
nor U21882 (N_21882,N_14389,N_12881);
nor U21883 (N_21883,N_15130,N_17178);
nor U21884 (N_21884,N_16691,N_13871);
and U21885 (N_21885,N_17883,N_12025);
xor U21886 (N_21886,N_12238,N_16936);
or U21887 (N_21887,N_17892,N_16980);
nor U21888 (N_21888,N_15099,N_15200);
and U21889 (N_21889,N_12376,N_14328);
and U21890 (N_21890,N_17057,N_16883);
nand U21891 (N_21891,N_15361,N_15123);
and U21892 (N_21892,N_14514,N_13920);
nor U21893 (N_21893,N_13140,N_12197);
or U21894 (N_21894,N_16005,N_12910);
xnor U21895 (N_21895,N_13615,N_17188);
nand U21896 (N_21896,N_15277,N_15282);
nor U21897 (N_21897,N_13626,N_17729);
nor U21898 (N_21898,N_13398,N_17090);
xnor U21899 (N_21899,N_16740,N_15098);
xnor U21900 (N_21900,N_17256,N_14110);
xor U21901 (N_21901,N_14289,N_14155);
nor U21902 (N_21902,N_12183,N_12121);
nand U21903 (N_21903,N_15060,N_15998);
and U21904 (N_21904,N_16140,N_14865);
nor U21905 (N_21905,N_16835,N_14886);
and U21906 (N_21906,N_17587,N_15758);
and U21907 (N_21907,N_12943,N_12594);
nor U21908 (N_21908,N_14932,N_14282);
xnor U21909 (N_21909,N_14793,N_16620);
and U21910 (N_21910,N_14108,N_15937);
and U21911 (N_21911,N_13980,N_13053);
and U21912 (N_21912,N_14772,N_12854);
xnor U21913 (N_21913,N_17103,N_14349);
and U21914 (N_21914,N_13832,N_12342);
nand U21915 (N_21915,N_16305,N_16295);
and U21916 (N_21916,N_16451,N_13188);
and U21917 (N_21917,N_13567,N_15794);
xor U21918 (N_21918,N_16377,N_17096);
nand U21919 (N_21919,N_17775,N_17504);
and U21920 (N_21920,N_12090,N_12772);
or U21921 (N_21921,N_17737,N_12753);
xor U21922 (N_21922,N_15448,N_15678);
nand U21923 (N_21923,N_16284,N_13340);
nor U21924 (N_21924,N_17182,N_15498);
or U21925 (N_21925,N_12985,N_15485);
nand U21926 (N_21926,N_15682,N_14628);
or U21927 (N_21927,N_15950,N_16932);
nand U21928 (N_21928,N_13966,N_14228);
nand U21929 (N_21929,N_15370,N_17349);
and U21930 (N_21930,N_15043,N_15188);
xor U21931 (N_21931,N_16794,N_13271);
or U21932 (N_21932,N_13598,N_12379);
or U21933 (N_21933,N_13219,N_12659);
nor U21934 (N_21934,N_16982,N_16834);
or U21935 (N_21935,N_14461,N_12184);
xor U21936 (N_21936,N_14724,N_12185);
and U21937 (N_21937,N_14102,N_15587);
nand U21938 (N_21938,N_17360,N_14962);
and U21939 (N_21939,N_14533,N_13164);
nor U21940 (N_21940,N_12063,N_16590);
nand U21941 (N_21941,N_13739,N_12541);
nand U21942 (N_21942,N_12256,N_15045);
and U21943 (N_21943,N_17637,N_13024);
and U21944 (N_21944,N_16785,N_15471);
nor U21945 (N_21945,N_16356,N_12548);
xnor U21946 (N_21946,N_13649,N_14113);
xnor U21947 (N_21947,N_14304,N_17208);
nand U21948 (N_21948,N_14981,N_17450);
nand U21949 (N_21949,N_12571,N_13282);
nor U21950 (N_21950,N_14404,N_12586);
or U21951 (N_21951,N_12756,N_15906);
nor U21952 (N_21952,N_13313,N_16965);
nor U21953 (N_21953,N_15179,N_17719);
nand U21954 (N_21954,N_17173,N_16100);
and U21955 (N_21955,N_12922,N_12789);
nor U21956 (N_21956,N_17754,N_14379);
or U21957 (N_21957,N_15207,N_12076);
nor U21958 (N_21958,N_13595,N_16994);
xor U21959 (N_21959,N_17616,N_12805);
xnor U21960 (N_21960,N_15276,N_13180);
nor U21961 (N_21961,N_12378,N_17080);
nand U21962 (N_21962,N_14079,N_14942);
or U21963 (N_21963,N_16388,N_17401);
nor U21964 (N_21964,N_12321,N_12615);
or U21965 (N_21965,N_13409,N_13012);
xor U21966 (N_21966,N_15796,N_15383);
and U21967 (N_21967,N_13253,N_13344);
nand U21968 (N_21968,N_17838,N_14922);
or U21969 (N_21969,N_17030,N_13923);
nand U21970 (N_21970,N_16270,N_13272);
and U21971 (N_21971,N_17526,N_17008);
or U21972 (N_21972,N_15692,N_17212);
or U21973 (N_21973,N_15192,N_17075);
and U21974 (N_21974,N_17627,N_14467);
nand U21975 (N_21975,N_17613,N_15905);
nand U21976 (N_21976,N_17845,N_13838);
nand U21977 (N_21977,N_12379,N_12757);
xnor U21978 (N_21978,N_14232,N_15828);
nor U21979 (N_21979,N_16707,N_12580);
xnor U21980 (N_21980,N_12909,N_14793);
and U21981 (N_21981,N_12394,N_14027);
and U21982 (N_21982,N_13103,N_15952);
xnor U21983 (N_21983,N_13496,N_12476);
nor U21984 (N_21984,N_13499,N_13252);
nand U21985 (N_21985,N_16006,N_15256);
nand U21986 (N_21986,N_12552,N_15759);
and U21987 (N_21987,N_16668,N_16123);
nand U21988 (N_21988,N_16542,N_15702);
nor U21989 (N_21989,N_13007,N_13756);
xnor U21990 (N_21990,N_15409,N_15374);
nor U21991 (N_21991,N_14528,N_15754);
and U21992 (N_21992,N_12783,N_15264);
xor U21993 (N_21993,N_13197,N_12191);
nor U21994 (N_21994,N_12677,N_15666);
nand U21995 (N_21995,N_16420,N_14990);
nor U21996 (N_21996,N_13882,N_14964);
nand U21997 (N_21997,N_13233,N_13833);
nor U21998 (N_21998,N_12754,N_17479);
nand U21999 (N_21999,N_16766,N_17688);
xnor U22000 (N_22000,N_14070,N_14870);
xor U22001 (N_22001,N_12672,N_13414);
and U22002 (N_22002,N_15198,N_12162);
nand U22003 (N_22003,N_17595,N_16208);
or U22004 (N_22004,N_13449,N_16145);
and U22005 (N_22005,N_14426,N_17901);
or U22006 (N_22006,N_16361,N_14709);
xor U22007 (N_22007,N_14245,N_12570);
and U22008 (N_22008,N_17455,N_17021);
nand U22009 (N_22009,N_12346,N_16552);
xor U22010 (N_22010,N_15851,N_15553);
nand U22011 (N_22011,N_14890,N_17200);
xnor U22012 (N_22012,N_15381,N_16196);
xor U22013 (N_22013,N_15909,N_14284);
xnor U22014 (N_22014,N_17153,N_15800);
or U22015 (N_22015,N_12367,N_12071);
nor U22016 (N_22016,N_13354,N_17756);
nor U22017 (N_22017,N_17241,N_16878);
and U22018 (N_22018,N_17224,N_12706);
or U22019 (N_22019,N_13029,N_14525);
xor U22020 (N_22020,N_17350,N_13143);
xnor U22021 (N_22021,N_14029,N_12156);
and U22022 (N_22022,N_12867,N_13505);
nor U22023 (N_22023,N_13254,N_14227);
or U22024 (N_22024,N_17392,N_16084);
nand U22025 (N_22025,N_14405,N_17976);
and U22026 (N_22026,N_12712,N_17378);
and U22027 (N_22027,N_15875,N_14165);
xor U22028 (N_22028,N_15680,N_14558);
nor U22029 (N_22029,N_16588,N_13877);
and U22030 (N_22030,N_16895,N_15557);
nor U22031 (N_22031,N_15176,N_14294);
nor U22032 (N_22032,N_17537,N_14999);
nor U22033 (N_22033,N_15190,N_12840);
and U22034 (N_22034,N_12048,N_13649);
nor U22035 (N_22035,N_12734,N_14577);
and U22036 (N_22036,N_17387,N_15845);
nor U22037 (N_22037,N_17293,N_12701);
or U22038 (N_22038,N_16762,N_14837);
xor U22039 (N_22039,N_15920,N_15071);
xor U22040 (N_22040,N_12233,N_13144);
nor U22041 (N_22041,N_14019,N_17629);
nand U22042 (N_22042,N_13082,N_15109);
and U22043 (N_22043,N_14753,N_14736);
and U22044 (N_22044,N_17933,N_15917);
and U22045 (N_22045,N_12712,N_13364);
and U22046 (N_22046,N_12744,N_13102);
and U22047 (N_22047,N_17683,N_15200);
and U22048 (N_22048,N_16046,N_12442);
and U22049 (N_22049,N_12706,N_13054);
and U22050 (N_22050,N_16318,N_16297);
xnor U22051 (N_22051,N_14443,N_13515);
nand U22052 (N_22052,N_12957,N_17871);
xor U22053 (N_22053,N_16241,N_15301);
nand U22054 (N_22054,N_15559,N_13350);
nand U22055 (N_22055,N_17020,N_14866);
or U22056 (N_22056,N_16927,N_14071);
and U22057 (N_22057,N_14253,N_16132);
and U22058 (N_22058,N_12695,N_13660);
nor U22059 (N_22059,N_12836,N_14105);
nand U22060 (N_22060,N_12167,N_12113);
nor U22061 (N_22061,N_16085,N_16621);
nand U22062 (N_22062,N_17144,N_15944);
or U22063 (N_22063,N_13626,N_17844);
nor U22064 (N_22064,N_17736,N_14359);
xnor U22065 (N_22065,N_13704,N_14063);
and U22066 (N_22066,N_13953,N_15302);
or U22067 (N_22067,N_17018,N_14900);
and U22068 (N_22068,N_12944,N_16191);
nand U22069 (N_22069,N_13072,N_16297);
nor U22070 (N_22070,N_14969,N_17098);
or U22071 (N_22071,N_12161,N_13391);
or U22072 (N_22072,N_13746,N_12325);
xnor U22073 (N_22073,N_15837,N_16584);
xor U22074 (N_22074,N_15571,N_17763);
and U22075 (N_22075,N_13377,N_13081);
xnor U22076 (N_22076,N_12963,N_17218);
nor U22077 (N_22077,N_13130,N_12084);
nor U22078 (N_22078,N_15637,N_14502);
nand U22079 (N_22079,N_17222,N_13154);
xor U22080 (N_22080,N_12637,N_17246);
nor U22081 (N_22081,N_15614,N_13765);
and U22082 (N_22082,N_12723,N_14589);
or U22083 (N_22083,N_13676,N_14301);
nand U22084 (N_22084,N_17232,N_15068);
xor U22085 (N_22085,N_16357,N_13803);
or U22086 (N_22086,N_14628,N_13457);
xnor U22087 (N_22087,N_12926,N_14454);
nor U22088 (N_22088,N_14055,N_12187);
and U22089 (N_22089,N_14775,N_12166);
nand U22090 (N_22090,N_15138,N_13105);
nand U22091 (N_22091,N_13749,N_16218);
and U22092 (N_22092,N_12329,N_12530);
and U22093 (N_22093,N_15639,N_14909);
nor U22094 (N_22094,N_14181,N_16480);
nor U22095 (N_22095,N_17516,N_15460);
xnor U22096 (N_22096,N_14614,N_17023);
or U22097 (N_22097,N_14175,N_12544);
nand U22098 (N_22098,N_12562,N_12945);
xnor U22099 (N_22099,N_16380,N_14411);
nor U22100 (N_22100,N_15171,N_13211);
nor U22101 (N_22101,N_12669,N_16941);
nor U22102 (N_22102,N_14317,N_13133);
nor U22103 (N_22103,N_14428,N_14670);
nor U22104 (N_22104,N_16564,N_13792);
xnor U22105 (N_22105,N_13050,N_14400);
nor U22106 (N_22106,N_16750,N_16469);
and U22107 (N_22107,N_12905,N_16941);
or U22108 (N_22108,N_12462,N_17020);
and U22109 (N_22109,N_14590,N_16502);
xnor U22110 (N_22110,N_16676,N_15316);
nand U22111 (N_22111,N_12008,N_14848);
and U22112 (N_22112,N_16991,N_13706);
nor U22113 (N_22113,N_13947,N_14659);
and U22114 (N_22114,N_17747,N_16373);
xnor U22115 (N_22115,N_15718,N_17297);
or U22116 (N_22116,N_13227,N_12576);
nand U22117 (N_22117,N_17831,N_12710);
and U22118 (N_22118,N_16589,N_16291);
or U22119 (N_22119,N_17588,N_15582);
or U22120 (N_22120,N_16166,N_15711);
nand U22121 (N_22121,N_12723,N_14144);
and U22122 (N_22122,N_17335,N_13753);
nand U22123 (N_22123,N_13133,N_12017);
nor U22124 (N_22124,N_13387,N_14973);
nand U22125 (N_22125,N_17266,N_17713);
xor U22126 (N_22126,N_17701,N_12014);
nand U22127 (N_22127,N_12840,N_17486);
and U22128 (N_22128,N_14365,N_15210);
or U22129 (N_22129,N_15942,N_13321);
nand U22130 (N_22130,N_15596,N_13649);
nand U22131 (N_22131,N_12559,N_16765);
or U22132 (N_22132,N_14334,N_12476);
nor U22133 (N_22133,N_16480,N_16758);
nor U22134 (N_22134,N_17078,N_15046);
nor U22135 (N_22135,N_14632,N_12212);
and U22136 (N_22136,N_12932,N_16122);
or U22137 (N_22137,N_12899,N_17957);
and U22138 (N_22138,N_16969,N_13080);
or U22139 (N_22139,N_12249,N_13963);
or U22140 (N_22140,N_12195,N_12219);
nor U22141 (N_22141,N_16308,N_13284);
nand U22142 (N_22142,N_15760,N_14342);
or U22143 (N_22143,N_14523,N_16406);
or U22144 (N_22144,N_16396,N_15413);
xor U22145 (N_22145,N_13516,N_16767);
xnor U22146 (N_22146,N_13569,N_13040);
or U22147 (N_22147,N_13560,N_14490);
xor U22148 (N_22148,N_16243,N_15604);
and U22149 (N_22149,N_15784,N_12817);
or U22150 (N_22150,N_15984,N_13809);
nand U22151 (N_22151,N_16583,N_14085);
nor U22152 (N_22152,N_14164,N_16716);
or U22153 (N_22153,N_14900,N_12693);
or U22154 (N_22154,N_14946,N_17330);
nor U22155 (N_22155,N_15778,N_15197);
nor U22156 (N_22156,N_16813,N_17092);
and U22157 (N_22157,N_13609,N_13791);
nor U22158 (N_22158,N_14783,N_14296);
or U22159 (N_22159,N_13356,N_13364);
nor U22160 (N_22160,N_15267,N_12701);
or U22161 (N_22161,N_12653,N_15597);
nand U22162 (N_22162,N_16247,N_16923);
xnor U22163 (N_22163,N_16138,N_15691);
nor U22164 (N_22164,N_13525,N_14074);
or U22165 (N_22165,N_14372,N_14146);
or U22166 (N_22166,N_15835,N_13525);
or U22167 (N_22167,N_14209,N_17125);
nand U22168 (N_22168,N_13277,N_16165);
or U22169 (N_22169,N_17631,N_12577);
or U22170 (N_22170,N_13802,N_17944);
xor U22171 (N_22171,N_15901,N_17655);
and U22172 (N_22172,N_15746,N_14826);
xnor U22173 (N_22173,N_15559,N_12988);
and U22174 (N_22174,N_12424,N_14690);
and U22175 (N_22175,N_17397,N_16792);
xnor U22176 (N_22176,N_13388,N_12044);
xor U22177 (N_22177,N_14206,N_14344);
and U22178 (N_22178,N_12324,N_12251);
xor U22179 (N_22179,N_14490,N_13688);
and U22180 (N_22180,N_16297,N_14291);
and U22181 (N_22181,N_15270,N_14866);
nor U22182 (N_22182,N_15621,N_14885);
and U22183 (N_22183,N_15281,N_15673);
nor U22184 (N_22184,N_16776,N_13121);
nor U22185 (N_22185,N_15708,N_17450);
nand U22186 (N_22186,N_14142,N_16438);
nor U22187 (N_22187,N_16710,N_15980);
xor U22188 (N_22188,N_14228,N_15557);
xor U22189 (N_22189,N_15757,N_12731);
or U22190 (N_22190,N_17435,N_12038);
nand U22191 (N_22191,N_12388,N_15311);
nor U22192 (N_22192,N_14609,N_14405);
nor U22193 (N_22193,N_12944,N_16821);
and U22194 (N_22194,N_15272,N_14820);
or U22195 (N_22195,N_16925,N_16255);
or U22196 (N_22196,N_15914,N_14775);
or U22197 (N_22197,N_13723,N_17811);
and U22198 (N_22198,N_16142,N_13809);
xor U22199 (N_22199,N_13104,N_16272);
and U22200 (N_22200,N_17834,N_15455);
nor U22201 (N_22201,N_14086,N_17055);
nand U22202 (N_22202,N_13069,N_17940);
nand U22203 (N_22203,N_14584,N_16683);
nor U22204 (N_22204,N_12706,N_15805);
and U22205 (N_22205,N_12938,N_16078);
nor U22206 (N_22206,N_14434,N_12621);
nand U22207 (N_22207,N_12982,N_14804);
or U22208 (N_22208,N_16427,N_17042);
or U22209 (N_22209,N_17734,N_13257);
nor U22210 (N_22210,N_15231,N_17539);
nor U22211 (N_22211,N_13880,N_15304);
or U22212 (N_22212,N_17232,N_14489);
nand U22213 (N_22213,N_12793,N_16992);
xor U22214 (N_22214,N_12734,N_14415);
or U22215 (N_22215,N_14769,N_16045);
nor U22216 (N_22216,N_12481,N_17372);
and U22217 (N_22217,N_15336,N_12792);
nand U22218 (N_22218,N_15160,N_12201);
nor U22219 (N_22219,N_15800,N_17170);
or U22220 (N_22220,N_15214,N_12790);
xor U22221 (N_22221,N_14401,N_16945);
or U22222 (N_22222,N_17648,N_16879);
and U22223 (N_22223,N_17144,N_17694);
nand U22224 (N_22224,N_14887,N_17703);
xnor U22225 (N_22225,N_17825,N_15770);
xor U22226 (N_22226,N_12708,N_14474);
xor U22227 (N_22227,N_14872,N_16309);
nor U22228 (N_22228,N_16666,N_12572);
or U22229 (N_22229,N_16968,N_17455);
or U22230 (N_22230,N_14556,N_13208);
and U22231 (N_22231,N_13717,N_14845);
nand U22232 (N_22232,N_14025,N_12753);
xnor U22233 (N_22233,N_17472,N_14188);
nand U22234 (N_22234,N_13500,N_14030);
nor U22235 (N_22235,N_17813,N_12548);
nor U22236 (N_22236,N_15657,N_16149);
nand U22237 (N_22237,N_12539,N_17069);
xor U22238 (N_22238,N_16579,N_17569);
and U22239 (N_22239,N_12467,N_12760);
nand U22240 (N_22240,N_13298,N_15471);
and U22241 (N_22241,N_15592,N_14535);
and U22242 (N_22242,N_12050,N_17336);
and U22243 (N_22243,N_14859,N_16350);
or U22244 (N_22244,N_16867,N_14000);
nor U22245 (N_22245,N_12539,N_17284);
nor U22246 (N_22246,N_16028,N_13221);
or U22247 (N_22247,N_15680,N_17981);
xor U22248 (N_22248,N_15266,N_17545);
and U22249 (N_22249,N_15895,N_15412);
or U22250 (N_22250,N_14681,N_16715);
and U22251 (N_22251,N_12797,N_13847);
nor U22252 (N_22252,N_14655,N_12577);
nand U22253 (N_22253,N_14420,N_16007);
nor U22254 (N_22254,N_13848,N_13557);
and U22255 (N_22255,N_17927,N_12594);
nor U22256 (N_22256,N_17729,N_13175);
nand U22257 (N_22257,N_13869,N_15504);
nand U22258 (N_22258,N_13503,N_14466);
nand U22259 (N_22259,N_15421,N_14195);
nand U22260 (N_22260,N_13949,N_16060);
and U22261 (N_22261,N_14322,N_12603);
and U22262 (N_22262,N_12636,N_13623);
xor U22263 (N_22263,N_14120,N_16329);
and U22264 (N_22264,N_13635,N_16818);
nor U22265 (N_22265,N_12913,N_15292);
nor U22266 (N_22266,N_16313,N_16613);
and U22267 (N_22267,N_16640,N_16427);
or U22268 (N_22268,N_13208,N_13032);
or U22269 (N_22269,N_15832,N_13866);
nand U22270 (N_22270,N_14218,N_16422);
or U22271 (N_22271,N_16108,N_14597);
and U22272 (N_22272,N_15411,N_13521);
nand U22273 (N_22273,N_12383,N_13468);
and U22274 (N_22274,N_14504,N_13648);
and U22275 (N_22275,N_17124,N_12919);
or U22276 (N_22276,N_17641,N_12870);
xnor U22277 (N_22277,N_12023,N_17743);
or U22278 (N_22278,N_15386,N_16653);
nor U22279 (N_22279,N_17889,N_14750);
xor U22280 (N_22280,N_16190,N_14121);
and U22281 (N_22281,N_15065,N_13261);
nand U22282 (N_22282,N_16330,N_17641);
and U22283 (N_22283,N_13101,N_12619);
xor U22284 (N_22284,N_16738,N_15377);
nor U22285 (N_22285,N_14742,N_12320);
xnor U22286 (N_22286,N_16675,N_14494);
nand U22287 (N_22287,N_14073,N_16881);
nor U22288 (N_22288,N_17635,N_16257);
and U22289 (N_22289,N_13456,N_15064);
xnor U22290 (N_22290,N_15918,N_13969);
xnor U22291 (N_22291,N_17794,N_12558);
nand U22292 (N_22292,N_17302,N_15441);
xor U22293 (N_22293,N_16459,N_16395);
nor U22294 (N_22294,N_16325,N_17453);
nand U22295 (N_22295,N_17758,N_12528);
or U22296 (N_22296,N_15136,N_14644);
and U22297 (N_22297,N_16682,N_13540);
and U22298 (N_22298,N_12727,N_16385);
xor U22299 (N_22299,N_16038,N_15133);
nor U22300 (N_22300,N_15101,N_15700);
nand U22301 (N_22301,N_17225,N_14876);
xnor U22302 (N_22302,N_16029,N_17108);
and U22303 (N_22303,N_12819,N_13982);
nand U22304 (N_22304,N_12244,N_15010);
xor U22305 (N_22305,N_16917,N_17445);
nand U22306 (N_22306,N_13193,N_16030);
or U22307 (N_22307,N_17337,N_17744);
nand U22308 (N_22308,N_13831,N_16522);
nand U22309 (N_22309,N_12618,N_16717);
nor U22310 (N_22310,N_12505,N_15506);
nor U22311 (N_22311,N_13509,N_17024);
nand U22312 (N_22312,N_13657,N_13396);
and U22313 (N_22313,N_16932,N_15947);
nand U22314 (N_22314,N_13593,N_14902);
or U22315 (N_22315,N_12203,N_13547);
xor U22316 (N_22316,N_14947,N_15348);
or U22317 (N_22317,N_15661,N_17885);
nand U22318 (N_22318,N_12119,N_12345);
nand U22319 (N_22319,N_13342,N_12623);
nand U22320 (N_22320,N_14610,N_14470);
nor U22321 (N_22321,N_12911,N_17734);
nor U22322 (N_22322,N_16411,N_15457);
xor U22323 (N_22323,N_15533,N_14531);
xor U22324 (N_22324,N_15984,N_16980);
or U22325 (N_22325,N_12547,N_13160);
nand U22326 (N_22326,N_13494,N_12905);
or U22327 (N_22327,N_14498,N_13014);
xor U22328 (N_22328,N_17940,N_15950);
nand U22329 (N_22329,N_16936,N_14721);
xor U22330 (N_22330,N_17703,N_13624);
and U22331 (N_22331,N_12884,N_16876);
nand U22332 (N_22332,N_13683,N_16984);
xor U22333 (N_22333,N_17264,N_16181);
and U22334 (N_22334,N_12540,N_15949);
nor U22335 (N_22335,N_16147,N_14029);
nand U22336 (N_22336,N_13332,N_15257);
nand U22337 (N_22337,N_12692,N_15420);
or U22338 (N_22338,N_16384,N_15180);
nor U22339 (N_22339,N_16099,N_17442);
or U22340 (N_22340,N_14313,N_17312);
nor U22341 (N_22341,N_12262,N_17142);
xor U22342 (N_22342,N_12157,N_14098);
nor U22343 (N_22343,N_14390,N_15130);
nor U22344 (N_22344,N_13897,N_17478);
or U22345 (N_22345,N_17844,N_14243);
xor U22346 (N_22346,N_17522,N_13728);
xnor U22347 (N_22347,N_14679,N_14118);
nand U22348 (N_22348,N_16344,N_17054);
xnor U22349 (N_22349,N_17586,N_15370);
nor U22350 (N_22350,N_12476,N_12775);
xnor U22351 (N_22351,N_17331,N_15573);
xnor U22352 (N_22352,N_12358,N_12821);
nand U22353 (N_22353,N_14391,N_13465);
and U22354 (N_22354,N_15508,N_14400);
nand U22355 (N_22355,N_14652,N_14062);
and U22356 (N_22356,N_16302,N_16987);
nand U22357 (N_22357,N_16052,N_16884);
nor U22358 (N_22358,N_13301,N_13610);
nor U22359 (N_22359,N_14989,N_15003);
and U22360 (N_22360,N_13253,N_12186);
nand U22361 (N_22361,N_17008,N_13094);
xnor U22362 (N_22362,N_17227,N_14379);
and U22363 (N_22363,N_16194,N_13669);
or U22364 (N_22364,N_17212,N_12471);
or U22365 (N_22365,N_12496,N_12948);
nand U22366 (N_22366,N_13905,N_14504);
xor U22367 (N_22367,N_13253,N_15942);
nand U22368 (N_22368,N_14458,N_15123);
and U22369 (N_22369,N_16128,N_17011);
nand U22370 (N_22370,N_17536,N_15226);
or U22371 (N_22371,N_17315,N_17249);
and U22372 (N_22372,N_13844,N_16242);
nor U22373 (N_22373,N_15388,N_15135);
and U22374 (N_22374,N_12985,N_15828);
nor U22375 (N_22375,N_15503,N_12870);
xor U22376 (N_22376,N_13784,N_15883);
and U22377 (N_22377,N_16243,N_14575);
nor U22378 (N_22378,N_13975,N_16811);
or U22379 (N_22379,N_13421,N_14085);
nor U22380 (N_22380,N_17545,N_14718);
nand U22381 (N_22381,N_14483,N_16052);
nand U22382 (N_22382,N_16660,N_13089);
xnor U22383 (N_22383,N_16511,N_13243);
nand U22384 (N_22384,N_14388,N_17748);
nor U22385 (N_22385,N_17181,N_15015);
and U22386 (N_22386,N_16501,N_12691);
xnor U22387 (N_22387,N_13733,N_14334);
or U22388 (N_22388,N_15509,N_17940);
nand U22389 (N_22389,N_17744,N_17398);
xor U22390 (N_22390,N_14369,N_14289);
nand U22391 (N_22391,N_14141,N_16898);
nor U22392 (N_22392,N_15425,N_13334);
and U22393 (N_22393,N_12727,N_16128);
and U22394 (N_22394,N_12786,N_12582);
xnor U22395 (N_22395,N_13641,N_15463);
or U22396 (N_22396,N_17886,N_17852);
nor U22397 (N_22397,N_12407,N_15413);
nor U22398 (N_22398,N_13681,N_15414);
and U22399 (N_22399,N_14621,N_13450);
nand U22400 (N_22400,N_15977,N_12063);
or U22401 (N_22401,N_15507,N_16207);
nor U22402 (N_22402,N_14213,N_12305);
xnor U22403 (N_22403,N_14663,N_13846);
nor U22404 (N_22404,N_13986,N_16500);
or U22405 (N_22405,N_16239,N_14128);
nor U22406 (N_22406,N_17864,N_15152);
nor U22407 (N_22407,N_13132,N_15247);
nor U22408 (N_22408,N_17849,N_17404);
nand U22409 (N_22409,N_14219,N_13657);
or U22410 (N_22410,N_14891,N_15916);
xor U22411 (N_22411,N_12977,N_14500);
and U22412 (N_22412,N_12883,N_16940);
and U22413 (N_22413,N_17216,N_15076);
nor U22414 (N_22414,N_15038,N_14906);
or U22415 (N_22415,N_15538,N_13644);
xnor U22416 (N_22416,N_16338,N_15803);
and U22417 (N_22417,N_16854,N_16198);
xor U22418 (N_22418,N_17424,N_17028);
or U22419 (N_22419,N_14802,N_14256);
and U22420 (N_22420,N_12676,N_17873);
or U22421 (N_22421,N_14346,N_13891);
and U22422 (N_22422,N_15778,N_14410);
nand U22423 (N_22423,N_17669,N_14737);
or U22424 (N_22424,N_13761,N_13771);
nand U22425 (N_22425,N_14478,N_17048);
nor U22426 (N_22426,N_14424,N_13371);
nand U22427 (N_22427,N_13128,N_17650);
or U22428 (N_22428,N_13001,N_13740);
and U22429 (N_22429,N_17181,N_17549);
or U22430 (N_22430,N_13948,N_15260);
or U22431 (N_22431,N_16126,N_15897);
nor U22432 (N_22432,N_13514,N_12042);
or U22433 (N_22433,N_15236,N_15832);
nand U22434 (N_22434,N_12209,N_14875);
nor U22435 (N_22435,N_17887,N_12651);
nor U22436 (N_22436,N_12337,N_15143);
or U22437 (N_22437,N_13385,N_17451);
or U22438 (N_22438,N_12965,N_12475);
nor U22439 (N_22439,N_12842,N_16069);
nand U22440 (N_22440,N_16475,N_17575);
and U22441 (N_22441,N_14463,N_15547);
or U22442 (N_22442,N_16780,N_12018);
nor U22443 (N_22443,N_14617,N_17122);
nand U22444 (N_22444,N_16007,N_16563);
nand U22445 (N_22445,N_17905,N_14714);
and U22446 (N_22446,N_12719,N_13527);
nand U22447 (N_22447,N_17417,N_13871);
and U22448 (N_22448,N_12279,N_14262);
and U22449 (N_22449,N_14955,N_15870);
or U22450 (N_22450,N_14887,N_12327);
nor U22451 (N_22451,N_12159,N_16073);
xnor U22452 (N_22452,N_15352,N_14624);
nand U22453 (N_22453,N_17560,N_12124);
nor U22454 (N_22454,N_16797,N_12307);
and U22455 (N_22455,N_15702,N_13609);
nand U22456 (N_22456,N_14273,N_17397);
nor U22457 (N_22457,N_17933,N_16287);
or U22458 (N_22458,N_12222,N_15073);
nand U22459 (N_22459,N_17770,N_17729);
nor U22460 (N_22460,N_13942,N_14841);
or U22461 (N_22461,N_15903,N_12423);
or U22462 (N_22462,N_13892,N_13847);
nand U22463 (N_22463,N_12066,N_14032);
or U22464 (N_22464,N_13593,N_15540);
or U22465 (N_22465,N_12095,N_17766);
xor U22466 (N_22466,N_12927,N_15595);
and U22467 (N_22467,N_16005,N_14610);
xnor U22468 (N_22468,N_17210,N_15919);
nor U22469 (N_22469,N_14458,N_15948);
or U22470 (N_22470,N_16970,N_13712);
and U22471 (N_22471,N_17482,N_12921);
nand U22472 (N_22472,N_17450,N_14813);
xor U22473 (N_22473,N_16417,N_17639);
xnor U22474 (N_22474,N_15403,N_16704);
and U22475 (N_22475,N_15021,N_14957);
xor U22476 (N_22476,N_14088,N_15951);
xor U22477 (N_22477,N_15010,N_15734);
xnor U22478 (N_22478,N_12665,N_17207);
xor U22479 (N_22479,N_15858,N_16900);
xnor U22480 (N_22480,N_12363,N_16293);
or U22481 (N_22481,N_17799,N_17412);
and U22482 (N_22482,N_13111,N_14711);
or U22483 (N_22483,N_12545,N_15274);
nor U22484 (N_22484,N_17990,N_17702);
or U22485 (N_22485,N_12616,N_16490);
xnor U22486 (N_22486,N_15154,N_15925);
nor U22487 (N_22487,N_17120,N_13163);
xnor U22488 (N_22488,N_16464,N_17540);
nor U22489 (N_22489,N_17959,N_17733);
xor U22490 (N_22490,N_13337,N_17319);
nand U22491 (N_22491,N_15168,N_13770);
nand U22492 (N_22492,N_14071,N_17316);
nor U22493 (N_22493,N_17403,N_17840);
nand U22494 (N_22494,N_16474,N_15006);
xor U22495 (N_22495,N_15814,N_17709);
xnor U22496 (N_22496,N_12758,N_15950);
xnor U22497 (N_22497,N_16346,N_15870);
nor U22498 (N_22498,N_14834,N_17702);
or U22499 (N_22499,N_12337,N_12232);
or U22500 (N_22500,N_17436,N_14851);
or U22501 (N_22501,N_16554,N_17190);
and U22502 (N_22502,N_15760,N_15562);
xor U22503 (N_22503,N_12568,N_17144);
and U22504 (N_22504,N_15631,N_15135);
nand U22505 (N_22505,N_15450,N_15225);
nand U22506 (N_22506,N_14928,N_13147);
xnor U22507 (N_22507,N_14368,N_15436);
nor U22508 (N_22508,N_13209,N_16214);
nor U22509 (N_22509,N_12698,N_12471);
nor U22510 (N_22510,N_14117,N_14429);
nor U22511 (N_22511,N_14188,N_17985);
xnor U22512 (N_22512,N_14422,N_13771);
xor U22513 (N_22513,N_14558,N_16459);
xnor U22514 (N_22514,N_13022,N_16303);
nor U22515 (N_22515,N_13262,N_16645);
or U22516 (N_22516,N_16626,N_15023);
nor U22517 (N_22517,N_14734,N_15952);
nand U22518 (N_22518,N_14042,N_15839);
or U22519 (N_22519,N_13027,N_15226);
xnor U22520 (N_22520,N_15239,N_14551);
xor U22521 (N_22521,N_17636,N_15425);
or U22522 (N_22522,N_14535,N_14181);
nor U22523 (N_22523,N_17015,N_15588);
nand U22524 (N_22524,N_12039,N_15593);
xnor U22525 (N_22525,N_16360,N_13643);
and U22526 (N_22526,N_12796,N_14495);
nor U22527 (N_22527,N_16915,N_14808);
or U22528 (N_22528,N_17913,N_13073);
xor U22529 (N_22529,N_15985,N_17178);
and U22530 (N_22530,N_13794,N_17075);
or U22531 (N_22531,N_12756,N_17106);
nand U22532 (N_22532,N_16076,N_16389);
nand U22533 (N_22533,N_12570,N_16351);
nor U22534 (N_22534,N_13068,N_13502);
nor U22535 (N_22535,N_17494,N_15861);
nor U22536 (N_22536,N_14598,N_17418);
or U22537 (N_22537,N_14313,N_16866);
or U22538 (N_22538,N_17729,N_14518);
xor U22539 (N_22539,N_13654,N_14145);
xor U22540 (N_22540,N_15127,N_13062);
and U22541 (N_22541,N_14649,N_16067);
nor U22542 (N_22542,N_15062,N_12689);
nor U22543 (N_22543,N_15463,N_13810);
nor U22544 (N_22544,N_12115,N_14159);
nor U22545 (N_22545,N_15215,N_12641);
or U22546 (N_22546,N_13727,N_12232);
nor U22547 (N_22547,N_12218,N_13144);
and U22548 (N_22548,N_16254,N_12763);
and U22549 (N_22549,N_14140,N_15663);
nor U22550 (N_22550,N_13246,N_12490);
xnor U22551 (N_22551,N_17112,N_14308);
and U22552 (N_22552,N_17719,N_17979);
or U22553 (N_22553,N_16483,N_13615);
or U22554 (N_22554,N_13097,N_17892);
nand U22555 (N_22555,N_17531,N_14767);
nand U22556 (N_22556,N_17190,N_15844);
and U22557 (N_22557,N_12433,N_13986);
nand U22558 (N_22558,N_12402,N_13993);
xor U22559 (N_22559,N_13812,N_16978);
xor U22560 (N_22560,N_17484,N_14145);
or U22561 (N_22561,N_15492,N_13400);
and U22562 (N_22562,N_16266,N_16220);
nand U22563 (N_22563,N_12655,N_13414);
nand U22564 (N_22564,N_16056,N_13324);
xnor U22565 (N_22565,N_16545,N_12500);
nor U22566 (N_22566,N_14045,N_16326);
or U22567 (N_22567,N_15287,N_15507);
xnor U22568 (N_22568,N_15029,N_14990);
or U22569 (N_22569,N_16700,N_16905);
xor U22570 (N_22570,N_14209,N_13817);
nor U22571 (N_22571,N_12137,N_16780);
and U22572 (N_22572,N_15175,N_15708);
xnor U22573 (N_22573,N_15269,N_14289);
nor U22574 (N_22574,N_16567,N_16260);
or U22575 (N_22575,N_17801,N_15372);
and U22576 (N_22576,N_16486,N_13803);
or U22577 (N_22577,N_16678,N_13289);
or U22578 (N_22578,N_12322,N_13151);
nand U22579 (N_22579,N_12157,N_17084);
nor U22580 (N_22580,N_15579,N_17179);
xnor U22581 (N_22581,N_15515,N_17769);
xor U22582 (N_22582,N_14166,N_12917);
or U22583 (N_22583,N_15108,N_15503);
or U22584 (N_22584,N_15149,N_12624);
nand U22585 (N_22585,N_12941,N_12929);
nor U22586 (N_22586,N_16130,N_12051);
nor U22587 (N_22587,N_17055,N_15954);
nand U22588 (N_22588,N_12572,N_13032);
nor U22589 (N_22589,N_17079,N_16937);
nand U22590 (N_22590,N_14399,N_14308);
or U22591 (N_22591,N_17532,N_12443);
nor U22592 (N_22592,N_17243,N_16716);
nor U22593 (N_22593,N_12737,N_15623);
and U22594 (N_22594,N_13953,N_12848);
or U22595 (N_22595,N_17508,N_16628);
nor U22596 (N_22596,N_14827,N_17278);
nor U22597 (N_22597,N_17554,N_13213);
and U22598 (N_22598,N_17490,N_17869);
nor U22599 (N_22599,N_15652,N_17054);
xor U22600 (N_22600,N_15539,N_17520);
or U22601 (N_22601,N_13283,N_17822);
nor U22602 (N_22602,N_14139,N_16198);
nand U22603 (N_22603,N_16386,N_15206);
or U22604 (N_22604,N_13168,N_15184);
or U22605 (N_22605,N_16411,N_17813);
or U22606 (N_22606,N_12236,N_15120);
and U22607 (N_22607,N_13289,N_14659);
nand U22608 (N_22608,N_17726,N_15343);
nor U22609 (N_22609,N_12232,N_13191);
nor U22610 (N_22610,N_17584,N_17794);
or U22611 (N_22611,N_16301,N_12822);
nor U22612 (N_22612,N_15228,N_17516);
and U22613 (N_22613,N_17676,N_12737);
nor U22614 (N_22614,N_14133,N_16466);
or U22615 (N_22615,N_12923,N_15150);
and U22616 (N_22616,N_17998,N_15817);
nand U22617 (N_22617,N_16930,N_13484);
and U22618 (N_22618,N_16560,N_15268);
and U22619 (N_22619,N_17476,N_16452);
or U22620 (N_22620,N_13508,N_16146);
and U22621 (N_22621,N_13497,N_15405);
nor U22622 (N_22622,N_13842,N_16049);
and U22623 (N_22623,N_16801,N_15389);
xor U22624 (N_22624,N_15418,N_15031);
xnor U22625 (N_22625,N_14527,N_12830);
or U22626 (N_22626,N_12351,N_14647);
xnor U22627 (N_22627,N_16528,N_15618);
and U22628 (N_22628,N_12004,N_13661);
and U22629 (N_22629,N_15737,N_15480);
nor U22630 (N_22630,N_16924,N_13492);
nand U22631 (N_22631,N_12220,N_12409);
nor U22632 (N_22632,N_12236,N_14189);
xnor U22633 (N_22633,N_15371,N_14828);
and U22634 (N_22634,N_13443,N_12456);
xor U22635 (N_22635,N_16625,N_17662);
xnor U22636 (N_22636,N_13134,N_12471);
nor U22637 (N_22637,N_12697,N_17647);
and U22638 (N_22638,N_15929,N_16404);
nand U22639 (N_22639,N_15939,N_16021);
and U22640 (N_22640,N_17212,N_16826);
nand U22641 (N_22641,N_16173,N_15866);
nor U22642 (N_22642,N_14662,N_14837);
or U22643 (N_22643,N_15806,N_17967);
xor U22644 (N_22644,N_16236,N_16873);
nand U22645 (N_22645,N_16417,N_14124);
nor U22646 (N_22646,N_13493,N_15541);
or U22647 (N_22647,N_15025,N_17221);
and U22648 (N_22648,N_14215,N_13914);
nand U22649 (N_22649,N_15073,N_15962);
xnor U22650 (N_22650,N_17258,N_16429);
xor U22651 (N_22651,N_13550,N_15365);
nand U22652 (N_22652,N_12208,N_15258);
nor U22653 (N_22653,N_14462,N_16362);
or U22654 (N_22654,N_12218,N_16935);
nor U22655 (N_22655,N_14674,N_14432);
nor U22656 (N_22656,N_14038,N_13200);
and U22657 (N_22657,N_17825,N_16203);
nand U22658 (N_22658,N_12430,N_14850);
nand U22659 (N_22659,N_14759,N_17494);
nor U22660 (N_22660,N_12075,N_16291);
and U22661 (N_22661,N_13690,N_16210);
and U22662 (N_22662,N_13208,N_16423);
nor U22663 (N_22663,N_14983,N_13225);
xor U22664 (N_22664,N_14263,N_15253);
and U22665 (N_22665,N_12519,N_13700);
xnor U22666 (N_22666,N_16481,N_15815);
xor U22667 (N_22667,N_17272,N_17761);
xnor U22668 (N_22668,N_14578,N_13798);
and U22669 (N_22669,N_14976,N_15558);
xnor U22670 (N_22670,N_15835,N_16748);
nor U22671 (N_22671,N_16068,N_15169);
nand U22672 (N_22672,N_14816,N_17815);
or U22673 (N_22673,N_15442,N_12438);
nand U22674 (N_22674,N_13995,N_17430);
and U22675 (N_22675,N_13118,N_12477);
and U22676 (N_22676,N_16921,N_14705);
xor U22677 (N_22677,N_13075,N_14295);
nand U22678 (N_22678,N_13697,N_15262);
nand U22679 (N_22679,N_14931,N_17005);
and U22680 (N_22680,N_13656,N_12098);
nand U22681 (N_22681,N_14125,N_15452);
nand U22682 (N_22682,N_15109,N_17089);
nor U22683 (N_22683,N_13761,N_17638);
or U22684 (N_22684,N_13239,N_14406);
nand U22685 (N_22685,N_15027,N_16600);
or U22686 (N_22686,N_16904,N_17924);
nand U22687 (N_22687,N_13280,N_13612);
xnor U22688 (N_22688,N_14159,N_14906);
and U22689 (N_22689,N_16619,N_14550);
xnor U22690 (N_22690,N_17289,N_15632);
xnor U22691 (N_22691,N_15567,N_15520);
nor U22692 (N_22692,N_12084,N_12716);
xnor U22693 (N_22693,N_14988,N_14412);
and U22694 (N_22694,N_13843,N_14283);
nor U22695 (N_22695,N_15726,N_16444);
nand U22696 (N_22696,N_13794,N_13188);
or U22697 (N_22697,N_12226,N_16334);
nand U22698 (N_22698,N_12595,N_15810);
nor U22699 (N_22699,N_17197,N_12595);
and U22700 (N_22700,N_17933,N_16498);
xnor U22701 (N_22701,N_13398,N_15935);
or U22702 (N_22702,N_14328,N_12445);
nor U22703 (N_22703,N_12512,N_15359);
or U22704 (N_22704,N_13672,N_14526);
nand U22705 (N_22705,N_12533,N_15011);
nand U22706 (N_22706,N_12700,N_12434);
nor U22707 (N_22707,N_16172,N_17317);
xor U22708 (N_22708,N_16027,N_17868);
xnor U22709 (N_22709,N_14421,N_13429);
nor U22710 (N_22710,N_13386,N_12598);
nand U22711 (N_22711,N_15168,N_12041);
or U22712 (N_22712,N_13485,N_12542);
nand U22713 (N_22713,N_12804,N_12197);
nand U22714 (N_22714,N_14779,N_16502);
xor U22715 (N_22715,N_14054,N_14461);
nor U22716 (N_22716,N_12230,N_17448);
and U22717 (N_22717,N_16669,N_17887);
or U22718 (N_22718,N_15346,N_12825);
or U22719 (N_22719,N_14349,N_13311);
or U22720 (N_22720,N_16375,N_14823);
and U22721 (N_22721,N_14227,N_12832);
or U22722 (N_22722,N_17734,N_15390);
and U22723 (N_22723,N_17642,N_13449);
and U22724 (N_22724,N_13743,N_12762);
and U22725 (N_22725,N_13206,N_16644);
or U22726 (N_22726,N_13402,N_16551);
xor U22727 (N_22727,N_14046,N_16234);
nor U22728 (N_22728,N_15526,N_16629);
nand U22729 (N_22729,N_14366,N_12440);
xnor U22730 (N_22730,N_15031,N_16041);
xor U22731 (N_22731,N_12075,N_14632);
and U22732 (N_22732,N_15721,N_14669);
nand U22733 (N_22733,N_15475,N_17466);
and U22734 (N_22734,N_17734,N_17873);
and U22735 (N_22735,N_15118,N_12408);
nor U22736 (N_22736,N_15464,N_17447);
nor U22737 (N_22737,N_15894,N_17660);
xor U22738 (N_22738,N_15339,N_17238);
nor U22739 (N_22739,N_12446,N_17822);
xor U22740 (N_22740,N_16110,N_13688);
or U22741 (N_22741,N_16082,N_12754);
nand U22742 (N_22742,N_16712,N_16113);
and U22743 (N_22743,N_15665,N_17774);
or U22744 (N_22744,N_17623,N_13395);
nand U22745 (N_22745,N_16018,N_16821);
xnor U22746 (N_22746,N_17510,N_17174);
nand U22747 (N_22747,N_15415,N_16972);
nand U22748 (N_22748,N_14441,N_14859);
or U22749 (N_22749,N_14004,N_14811);
or U22750 (N_22750,N_14582,N_12271);
and U22751 (N_22751,N_14259,N_12272);
and U22752 (N_22752,N_17141,N_15444);
nand U22753 (N_22753,N_14807,N_12863);
or U22754 (N_22754,N_15831,N_15278);
xor U22755 (N_22755,N_15823,N_12425);
nand U22756 (N_22756,N_16638,N_17172);
nor U22757 (N_22757,N_14302,N_14238);
nand U22758 (N_22758,N_12518,N_14424);
and U22759 (N_22759,N_15270,N_12195);
xnor U22760 (N_22760,N_12071,N_17330);
nor U22761 (N_22761,N_15897,N_14589);
and U22762 (N_22762,N_16249,N_12974);
nor U22763 (N_22763,N_17497,N_15231);
nor U22764 (N_22764,N_17590,N_14607);
and U22765 (N_22765,N_14680,N_12967);
or U22766 (N_22766,N_12243,N_14759);
xnor U22767 (N_22767,N_17052,N_17130);
nand U22768 (N_22768,N_15004,N_13362);
or U22769 (N_22769,N_17009,N_14422);
nand U22770 (N_22770,N_15680,N_14048);
or U22771 (N_22771,N_12118,N_15546);
xnor U22772 (N_22772,N_15986,N_16018);
or U22773 (N_22773,N_14286,N_14212);
xor U22774 (N_22774,N_16351,N_15023);
nand U22775 (N_22775,N_14774,N_16303);
or U22776 (N_22776,N_14262,N_14927);
or U22777 (N_22777,N_14782,N_14643);
xnor U22778 (N_22778,N_15422,N_14145);
or U22779 (N_22779,N_15326,N_16910);
and U22780 (N_22780,N_14192,N_15170);
xor U22781 (N_22781,N_13338,N_17700);
nor U22782 (N_22782,N_16786,N_12014);
xor U22783 (N_22783,N_14293,N_13144);
xor U22784 (N_22784,N_12418,N_16691);
xor U22785 (N_22785,N_16349,N_15552);
nand U22786 (N_22786,N_12225,N_12733);
or U22787 (N_22787,N_16063,N_13721);
and U22788 (N_22788,N_14015,N_14128);
nand U22789 (N_22789,N_12801,N_17697);
nand U22790 (N_22790,N_16874,N_14586);
and U22791 (N_22791,N_12193,N_16167);
nand U22792 (N_22792,N_17410,N_13019);
or U22793 (N_22793,N_16676,N_15701);
xor U22794 (N_22794,N_12109,N_17862);
nor U22795 (N_22795,N_12518,N_12110);
or U22796 (N_22796,N_17300,N_14729);
nand U22797 (N_22797,N_17108,N_12112);
or U22798 (N_22798,N_15336,N_17626);
nor U22799 (N_22799,N_15344,N_16644);
or U22800 (N_22800,N_14045,N_15875);
or U22801 (N_22801,N_17183,N_15047);
nand U22802 (N_22802,N_13094,N_17248);
nand U22803 (N_22803,N_13039,N_12650);
nand U22804 (N_22804,N_17009,N_14444);
nand U22805 (N_22805,N_15225,N_17858);
nand U22806 (N_22806,N_12765,N_13977);
xor U22807 (N_22807,N_17535,N_12905);
and U22808 (N_22808,N_12667,N_12880);
xnor U22809 (N_22809,N_17105,N_16667);
xnor U22810 (N_22810,N_17111,N_14086);
or U22811 (N_22811,N_12199,N_13963);
and U22812 (N_22812,N_14565,N_16534);
xnor U22813 (N_22813,N_15429,N_12493);
and U22814 (N_22814,N_13978,N_13159);
and U22815 (N_22815,N_14617,N_14732);
or U22816 (N_22816,N_17975,N_16337);
nand U22817 (N_22817,N_13571,N_16719);
or U22818 (N_22818,N_17822,N_17759);
and U22819 (N_22819,N_12007,N_17611);
xor U22820 (N_22820,N_15391,N_14202);
and U22821 (N_22821,N_17093,N_14402);
and U22822 (N_22822,N_15666,N_14729);
nand U22823 (N_22823,N_13217,N_15788);
xor U22824 (N_22824,N_17549,N_12018);
nand U22825 (N_22825,N_14644,N_12300);
or U22826 (N_22826,N_15235,N_13148);
and U22827 (N_22827,N_16227,N_12912);
or U22828 (N_22828,N_14851,N_17659);
xor U22829 (N_22829,N_15640,N_13862);
and U22830 (N_22830,N_15002,N_16137);
nor U22831 (N_22831,N_12749,N_14953);
and U22832 (N_22832,N_16487,N_13059);
or U22833 (N_22833,N_17325,N_15170);
or U22834 (N_22834,N_14522,N_13681);
nand U22835 (N_22835,N_14882,N_17609);
xnor U22836 (N_22836,N_16863,N_17436);
nor U22837 (N_22837,N_13603,N_12374);
nand U22838 (N_22838,N_15426,N_17197);
xnor U22839 (N_22839,N_16846,N_16489);
xnor U22840 (N_22840,N_15224,N_17610);
nand U22841 (N_22841,N_12548,N_14883);
xnor U22842 (N_22842,N_17443,N_13213);
and U22843 (N_22843,N_15168,N_15635);
nor U22844 (N_22844,N_13872,N_14200);
nor U22845 (N_22845,N_13673,N_14033);
nor U22846 (N_22846,N_17643,N_13010);
nand U22847 (N_22847,N_15625,N_17871);
nand U22848 (N_22848,N_12757,N_13674);
and U22849 (N_22849,N_13954,N_16422);
and U22850 (N_22850,N_12278,N_13134);
nand U22851 (N_22851,N_16217,N_12990);
xor U22852 (N_22852,N_14426,N_16026);
and U22853 (N_22853,N_15556,N_17921);
or U22854 (N_22854,N_16834,N_16417);
nor U22855 (N_22855,N_16363,N_13899);
and U22856 (N_22856,N_12058,N_17608);
xnor U22857 (N_22857,N_15946,N_16732);
nor U22858 (N_22858,N_14371,N_14179);
and U22859 (N_22859,N_13276,N_17851);
and U22860 (N_22860,N_12906,N_16339);
or U22861 (N_22861,N_14324,N_17204);
xor U22862 (N_22862,N_13839,N_16155);
xnor U22863 (N_22863,N_13521,N_17123);
nand U22864 (N_22864,N_17549,N_15919);
nor U22865 (N_22865,N_16683,N_13103);
xor U22866 (N_22866,N_12957,N_17029);
nor U22867 (N_22867,N_14887,N_15169);
nor U22868 (N_22868,N_12769,N_13232);
and U22869 (N_22869,N_15705,N_15777);
and U22870 (N_22870,N_14528,N_13102);
nor U22871 (N_22871,N_15490,N_12230);
and U22872 (N_22872,N_15456,N_13127);
nor U22873 (N_22873,N_15713,N_16061);
xnor U22874 (N_22874,N_14508,N_15591);
and U22875 (N_22875,N_13502,N_12354);
or U22876 (N_22876,N_12264,N_13117);
and U22877 (N_22877,N_15334,N_15045);
or U22878 (N_22878,N_13838,N_14987);
nand U22879 (N_22879,N_15200,N_17375);
nand U22880 (N_22880,N_13983,N_12217);
xor U22881 (N_22881,N_13687,N_14834);
nand U22882 (N_22882,N_16736,N_15202);
nor U22883 (N_22883,N_12858,N_12317);
nand U22884 (N_22884,N_16094,N_14625);
xnor U22885 (N_22885,N_17188,N_13066);
nor U22886 (N_22886,N_17311,N_16165);
xnor U22887 (N_22887,N_17194,N_15714);
nor U22888 (N_22888,N_17994,N_17268);
or U22889 (N_22889,N_14291,N_17344);
xor U22890 (N_22890,N_16048,N_14272);
nor U22891 (N_22891,N_17500,N_14110);
or U22892 (N_22892,N_12831,N_17500);
xor U22893 (N_22893,N_15275,N_17891);
nand U22894 (N_22894,N_14171,N_13774);
xnor U22895 (N_22895,N_13732,N_12766);
xnor U22896 (N_22896,N_16694,N_13776);
xnor U22897 (N_22897,N_16841,N_13925);
or U22898 (N_22898,N_17605,N_16838);
or U22899 (N_22899,N_13433,N_13137);
nor U22900 (N_22900,N_12018,N_12213);
xnor U22901 (N_22901,N_13835,N_13218);
and U22902 (N_22902,N_13793,N_17561);
and U22903 (N_22903,N_16255,N_15885);
or U22904 (N_22904,N_17027,N_12411);
nor U22905 (N_22905,N_13199,N_14092);
and U22906 (N_22906,N_14462,N_12741);
nand U22907 (N_22907,N_12713,N_15441);
or U22908 (N_22908,N_13069,N_13195);
xnor U22909 (N_22909,N_16612,N_15205);
nor U22910 (N_22910,N_15971,N_17595);
nand U22911 (N_22911,N_16907,N_12253);
nor U22912 (N_22912,N_13282,N_16128);
xnor U22913 (N_22913,N_14372,N_13115);
and U22914 (N_22914,N_14693,N_15315);
nand U22915 (N_22915,N_14814,N_14900);
xnor U22916 (N_22916,N_13687,N_15042);
or U22917 (N_22917,N_12016,N_14372);
and U22918 (N_22918,N_14419,N_13714);
nor U22919 (N_22919,N_12257,N_14519);
and U22920 (N_22920,N_14289,N_15246);
nand U22921 (N_22921,N_16347,N_12632);
or U22922 (N_22922,N_14066,N_15843);
nor U22923 (N_22923,N_15650,N_15585);
nand U22924 (N_22924,N_14867,N_16305);
or U22925 (N_22925,N_12182,N_14270);
nand U22926 (N_22926,N_16960,N_12626);
xor U22927 (N_22927,N_17397,N_16230);
xor U22928 (N_22928,N_13783,N_13816);
nand U22929 (N_22929,N_14699,N_16072);
xnor U22930 (N_22930,N_15757,N_16220);
or U22931 (N_22931,N_13738,N_12058);
nand U22932 (N_22932,N_12077,N_14985);
and U22933 (N_22933,N_16636,N_14540);
or U22934 (N_22934,N_13734,N_15294);
nand U22935 (N_22935,N_15235,N_16357);
or U22936 (N_22936,N_15512,N_14785);
or U22937 (N_22937,N_16958,N_14061);
and U22938 (N_22938,N_15682,N_16671);
xor U22939 (N_22939,N_17448,N_14438);
nor U22940 (N_22940,N_13789,N_17408);
xnor U22941 (N_22941,N_15533,N_14836);
nor U22942 (N_22942,N_14338,N_17448);
xnor U22943 (N_22943,N_14916,N_15403);
or U22944 (N_22944,N_13893,N_15696);
or U22945 (N_22945,N_16003,N_17557);
xor U22946 (N_22946,N_16830,N_17186);
and U22947 (N_22947,N_13369,N_12505);
or U22948 (N_22948,N_14241,N_13326);
or U22949 (N_22949,N_17387,N_17627);
nor U22950 (N_22950,N_17420,N_13773);
and U22951 (N_22951,N_12194,N_17674);
xor U22952 (N_22952,N_12220,N_14545);
and U22953 (N_22953,N_16536,N_17530);
xnor U22954 (N_22954,N_17739,N_16120);
nor U22955 (N_22955,N_13155,N_17066);
and U22956 (N_22956,N_15088,N_13312);
xor U22957 (N_22957,N_17318,N_13246);
nor U22958 (N_22958,N_15613,N_13782);
nand U22959 (N_22959,N_14969,N_12023);
and U22960 (N_22960,N_15165,N_13522);
xnor U22961 (N_22961,N_15083,N_12597);
and U22962 (N_22962,N_12483,N_14763);
nand U22963 (N_22963,N_16760,N_12808);
and U22964 (N_22964,N_12221,N_14997);
nor U22965 (N_22965,N_13250,N_15867);
and U22966 (N_22966,N_17372,N_14160);
and U22967 (N_22967,N_14954,N_12979);
nand U22968 (N_22968,N_17528,N_15995);
and U22969 (N_22969,N_16494,N_12526);
nand U22970 (N_22970,N_17243,N_15168);
and U22971 (N_22971,N_17519,N_16923);
xor U22972 (N_22972,N_13139,N_13628);
or U22973 (N_22973,N_13664,N_17169);
nor U22974 (N_22974,N_13089,N_12836);
xor U22975 (N_22975,N_15677,N_15306);
xnor U22976 (N_22976,N_15384,N_17742);
nand U22977 (N_22977,N_12068,N_14554);
nand U22978 (N_22978,N_16899,N_17120);
nand U22979 (N_22979,N_17954,N_14184);
xnor U22980 (N_22980,N_15377,N_12628);
nor U22981 (N_22981,N_17355,N_15174);
and U22982 (N_22982,N_15535,N_17607);
nand U22983 (N_22983,N_15268,N_17751);
or U22984 (N_22984,N_15038,N_12341);
and U22985 (N_22985,N_16600,N_14015);
and U22986 (N_22986,N_17900,N_13222);
nor U22987 (N_22987,N_15550,N_13828);
nor U22988 (N_22988,N_16072,N_12489);
nor U22989 (N_22989,N_15794,N_17799);
nor U22990 (N_22990,N_13644,N_15891);
or U22991 (N_22991,N_15950,N_17085);
nor U22992 (N_22992,N_15995,N_12878);
nand U22993 (N_22993,N_13980,N_13323);
xor U22994 (N_22994,N_12535,N_16107);
and U22995 (N_22995,N_16371,N_13374);
xnor U22996 (N_22996,N_14940,N_13997);
nand U22997 (N_22997,N_17472,N_13136);
xor U22998 (N_22998,N_14540,N_14529);
nor U22999 (N_22999,N_13904,N_13105);
nand U23000 (N_23000,N_14018,N_17334);
xor U23001 (N_23001,N_15729,N_14114);
or U23002 (N_23002,N_17875,N_17207);
nand U23003 (N_23003,N_12033,N_14102);
nand U23004 (N_23004,N_17008,N_16514);
and U23005 (N_23005,N_17407,N_15941);
nand U23006 (N_23006,N_16225,N_14147);
xnor U23007 (N_23007,N_14838,N_17963);
nor U23008 (N_23008,N_13988,N_13380);
or U23009 (N_23009,N_17658,N_12936);
or U23010 (N_23010,N_12036,N_12882);
nor U23011 (N_23011,N_13478,N_15990);
and U23012 (N_23012,N_17021,N_16841);
xnor U23013 (N_23013,N_13433,N_16282);
and U23014 (N_23014,N_12274,N_15585);
nand U23015 (N_23015,N_12352,N_13353);
or U23016 (N_23016,N_12584,N_14422);
xnor U23017 (N_23017,N_17486,N_13535);
nand U23018 (N_23018,N_16541,N_17874);
nor U23019 (N_23019,N_17766,N_12367);
xnor U23020 (N_23020,N_16379,N_14454);
nand U23021 (N_23021,N_15811,N_12588);
nor U23022 (N_23022,N_17864,N_16216);
xnor U23023 (N_23023,N_13129,N_14845);
or U23024 (N_23024,N_16768,N_14113);
nand U23025 (N_23025,N_13665,N_12811);
and U23026 (N_23026,N_14420,N_12409);
nand U23027 (N_23027,N_17098,N_16925);
nor U23028 (N_23028,N_16315,N_17935);
nand U23029 (N_23029,N_17757,N_14962);
nor U23030 (N_23030,N_12067,N_14926);
and U23031 (N_23031,N_16284,N_14472);
nand U23032 (N_23032,N_13870,N_14989);
nand U23033 (N_23033,N_17615,N_13713);
xor U23034 (N_23034,N_13604,N_13792);
or U23035 (N_23035,N_12599,N_17998);
or U23036 (N_23036,N_12365,N_13653);
and U23037 (N_23037,N_15635,N_13583);
nand U23038 (N_23038,N_13234,N_12914);
nor U23039 (N_23039,N_12296,N_14844);
nor U23040 (N_23040,N_14934,N_13220);
nor U23041 (N_23041,N_14210,N_17076);
and U23042 (N_23042,N_13653,N_14536);
or U23043 (N_23043,N_14736,N_14273);
xnor U23044 (N_23044,N_14640,N_15346);
nand U23045 (N_23045,N_15918,N_15823);
nor U23046 (N_23046,N_13958,N_17166);
nor U23047 (N_23047,N_17131,N_13693);
nor U23048 (N_23048,N_16441,N_15452);
nor U23049 (N_23049,N_13572,N_14767);
nand U23050 (N_23050,N_15613,N_17130);
xnor U23051 (N_23051,N_15991,N_17195);
or U23052 (N_23052,N_14543,N_16901);
xnor U23053 (N_23053,N_15090,N_17440);
and U23054 (N_23054,N_13852,N_15314);
and U23055 (N_23055,N_13013,N_17715);
or U23056 (N_23056,N_15070,N_17842);
xnor U23057 (N_23057,N_13113,N_16119);
xnor U23058 (N_23058,N_17814,N_14146);
or U23059 (N_23059,N_15208,N_14992);
nand U23060 (N_23060,N_13692,N_15721);
and U23061 (N_23061,N_15900,N_13134);
xnor U23062 (N_23062,N_14852,N_17376);
nand U23063 (N_23063,N_15764,N_14149);
nor U23064 (N_23064,N_15563,N_17426);
nand U23065 (N_23065,N_15265,N_15684);
nor U23066 (N_23066,N_14603,N_15503);
or U23067 (N_23067,N_12103,N_15093);
and U23068 (N_23068,N_16006,N_13628);
and U23069 (N_23069,N_14092,N_16942);
nor U23070 (N_23070,N_13239,N_16635);
nand U23071 (N_23071,N_14941,N_13465);
nand U23072 (N_23072,N_16116,N_17696);
or U23073 (N_23073,N_17552,N_13623);
or U23074 (N_23074,N_15600,N_13223);
xnor U23075 (N_23075,N_15102,N_14479);
xor U23076 (N_23076,N_13156,N_17116);
and U23077 (N_23077,N_15349,N_14922);
xnor U23078 (N_23078,N_17311,N_14685);
nor U23079 (N_23079,N_15681,N_13279);
or U23080 (N_23080,N_12331,N_16677);
xor U23081 (N_23081,N_13874,N_15695);
nand U23082 (N_23082,N_17544,N_14538);
or U23083 (N_23083,N_14733,N_12125);
and U23084 (N_23084,N_13645,N_16595);
and U23085 (N_23085,N_16200,N_12536);
or U23086 (N_23086,N_13782,N_12943);
nand U23087 (N_23087,N_16107,N_12261);
and U23088 (N_23088,N_13824,N_15888);
nor U23089 (N_23089,N_15050,N_16298);
xor U23090 (N_23090,N_15765,N_12711);
xor U23091 (N_23091,N_14734,N_13121);
nand U23092 (N_23092,N_13359,N_17500);
nor U23093 (N_23093,N_16626,N_16081);
nor U23094 (N_23094,N_17540,N_12018);
nor U23095 (N_23095,N_14575,N_14139);
nor U23096 (N_23096,N_12895,N_12606);
nor U23097 (N_23097,N_15271,N_14699);
nand U23098 (N_23098,N_15001,N_13141);
xor U23099 (N_23099,N_17061,N_14085);
or U23100 (N_23100,N_14117,N_15649);
nand U23101 (N_23101,N_12405,N_14061);
nor U23102 (N_23102,N_16697,N_13706);
xnor U23103 (N_23103,N_12425,N_16687);
and U23104 (N_23104,N_15822,N_15890);
nand U23105 (N_23105,N_17007,N_12698);
and U23106 (N_23106,N_17682,N_17620);
nand U23107 (N_23107,N_15998,N_14814);
xor U23108 (N_23108,N_16070,N_14055);
nor U23109 (N_23109,N_17110,N_16633);
nor U23110 (N_23110,N_12404,N_15320);
or U23111 (N_23111,N_13792,N_15301);
xor U23112 (N_23112,N_14736,N_16319);
or U23113 (N_23113,N_14850,N_12598);
nor U23114 (N_23114,N_16152,N_13853);
nand U23115 (N_23115,N_16753,N_17783);
nand U23116 (N_23116,N_17179,N_14411);
xor U23117 (N_23117,N_15563,N_17289);
xnor U23118 (N_23118,N_15048,N_15818);
xnor U23119 (N_23119,N_16304,N_14631);
nor U23120 (N_23120,N_15056,N_16526);
nand U23121 (N_23121,N_12907,N_15089);
and U23122 (N_23122,N_16101,N_13994);
nand U23123 (N_23123,N_14270,N_17452);
nand U23124 (N_23124,N_16797,N_12609);
and U23125 (N_23125,N_14097,N_14425);
nor U23126 (N_23126,N_12695,N_15315);
xnor U23127 (N_23127,N_17648,N_12476);
nand U23128 (N_23128,N_14703,N_15798);
nand U23129 (N_23129,N_14692,N_16294);
or U23130 (N_23130,N_17804,N_16286);
nor U23131 (N_23131,N_12769,N_15600);
and U23132 (N_23132,N_17904,N_14193);
nand U23133 (N_23133,N_13132,N_15431);
and U23134 (N_23134,N_12665,N_14032);
and U23135 (N_23135,N_15193,N_15595);
or U23136 (N_23136,N_13591,N_14288);
nand U23137 (N_23137,N_15941,N_16565);
and U23138 (N_23138,N_12408,N_16507);
nor U23139 (N_23139,N_12709,N_16549);
and U23140 (N_23140,N_16169,N_12161);
nor U23141 (N_23141,N_17832,N_14895);
or U23142 (N_23142,N_14461,N_17888);
or U23143 (N_23143,N_15350,N_12300);
xor U23144 (N_23144,N_17056,N_13084);
nand U23145 (N_23145,N_17137,N_13034);
nor U23146 (N_23146,N_16923,N_17526);
nor U23147 (N_23147,N_16390,N_14555);
and U23148 (N_23148,N_14564,N_15749);
and U23149 (N_23149,N_14236,N_16620);
xor U23150 (N_23150,N_17173,N_14814);
and U23151 (N_23151,N_16609,N_16645);
nor U23152 (N_23152,N_14656,N_13197);
or U23153 (N_23153,N_17957,N_16091);
or U23154 (N_23154,N_14181,N_12125);
nand U23155 (N_23155,N_17970,N_16602);
xnor U23156 (N_23156,N_12489,N_16334);
nand U23157 (N_23157,N_13372,N_15727);
nand U23158 (N_23158,N_16690,N_17242);
nor U23159 (N_23159,N_15909,N_13624);
nand U23160 (N_23160,N_15691,N_16093);
nand U23161 (N_23161,N_13112,N_14602);
nand U23162 (N_23162,N_12806,N_17698);
or U23163 (N_23163,N_16862,N_15696);
nor U23164 (N_23164,N_17847,N_12897);
nand U23165 (N_23165,N_14269,N_17538);
xnor U23166 (N_23166,N_13768,N_14090);
xnor U23167 (N_23167,N_16797,N_17927);
and U23168 (N_23168,N_14580,N_13769);
xnor U23169 (N_23169,N_16479,N_17625);
or U23170 (N_23170,N_14918,N_13269);
nor U23171 (N_23171,N_16121,N_16639);
and U23172 (N_23172,N_15598,N_12240);
nand U23173 (N_23173,N_17720,N_14675);
or U23174 (N_23174,N_16751,N_13449);
or U23175 (N_23175,N_16189,N_12492);
nor U23176 (N_23176,N_14375,N_15583);
and U23177 (N_23177,N_13982,N_12902);
nor U23178 (N_23178,N_14667,N_17450);
nand U23179 (N_23179,N_17975,N_13592);
and U23180 (N_23180,N_13530,N_14539);
nor U23181 (N_23181,N_15326,N_14383);
or U23182 (N_23182,N_13030,N_13607);
or U23183 (N_23183,N_12582,N_17783);
or U23184 (N_23184,N_17860,N_13391);
or U23185 (N_23185,N_15344,N_13760);
or U23186 (N_23186,N_13737,N_17461);
nand U23187 (N_23187,N_15596,N_17673);
nor U23188 (N_23188,N_15533,N_13237);
and U23189 (N_23189,N_13892,N_13681);
or U23190 (N_23190,N_13655,N_17106);
or U23191 (N_23191,N_15340,N_14031);
xor U23192 (N_23192,N_16372,N_12065);
nand U23193 (N_23193,N_17553,N_16560);
or U23194 (N_23194,N_14033,N_14656);
nand U23195 (N_23195,N_16581,N_14794);
nand U23196 (N_23196,N_14019,N_14732);
and U23197 (N_23197,N_16538,N_16239);
and U23198 (N_23198,N_13996,N_12377);
and U23199 (N_23199,N_14021,N_16491);
and U23200 (N_23200,N_12952,N_15408);
nor U23201 (N_23201,N_16574,N_15247);
nor U23202 (N_23202,N_16316,N_16787);
and U23203 (N_23203,N_13647,N_15924);
nor U23204 (N_23204,N_12928,N_15052);
or U23205 (N_23205,N_16264,N_13759);
and U23206 (N_23206,N_14905,N_14652);
or U23207 (N_23207,N_12144,N_15632);
or U23208 (N_23208,N_17864,N_13765);
or U23209 (N_23209,N_15703,N_13829);
xor U23210 (N_23210,N_13917,N_13636);
or U23211 (N_23211,N_13955,N_17670);
nand U23212 (N_23212,N_14691,N_12671);
and U23213 (N_23213,N_15709,N_14315);
and U23214 (N_23214,N_16997,N_14673);
nor U23215 (N_23215,N_17110,N_12441);
xor U23216 (N_23216,N_17761,N_13350);
nor U23217 (N_23217,N_14915,N_13251);
xnor U23218 (N_23218,N_13267,N_16487);
xnor U23219 (N_23219,N_12756,N_13418);
or U23220 (N_23220,N_15277,N_17107);
nand U23221 (N_23221,N_13207,N_14028);
or U23222 (N_23222,N_12824,N_17677);
nor U23223 (N_23223,N_12780,N_16040);
nor U23224 (N_23224,N_12528,N_17599);
nand U23225 (N_23225,N_15094,N_17791);
xnor U23226 (N_23226,N_13649,N_14188);
xor U23227 (N_23227,N_15593,N_16991);
xor U23228 (N_23228,N_17033,N_17079);
xnor U23229 (N_23229,N_13365,N_13924);
nand U23230 (N_23230,N_12018,N_13750);
or U23231 (N_23231,N_16150,N_14259);
xnor U23232 (N_23232,N_15413,N_12229);
xnor U23233 (N_23233,N_13585,N_13329);
or U23234 (N_23234,N_13776,N_13029);
nor U23235 (N_23235,N_15205,N_15820);
or U23236 (N_23236,N_17787,N_13064);
and U23237 (N_23237,N_14784,N_13571);
xnor U23238 (N_23238,N_17824,N_15772);
nand U23239 (N_23239,N_15631,N_12208);
or U23240 (N_23240,N_15295,N_13776);
xnor U23241 (N_23241,N_12533,N_15806);
xnor U23242 (N_23242,N_12437,N_12931);
xnor U23243 (N_23243,N_14464,N_17403);
nor U23244 (N_23244,N_14029,N_15064);
or U23245 (N_23245,N_16165,N_14339);
xor U23246 (N_23246,N_15143,N_14435);
or U23247 (N_23247,N_17322,N_14461);
nor U23248 (N_23248,N_12384,N_16185);
nand U23249 (N_23249,N_16505,N_13416);
nand U23250 (N_23250,N_13024,N_17302);
nand U23251 (N_23251,N_14224,N_14199);
or U23252 (N_23252,N_15528,N_12877);
xnor U23253 (N_23253,N_13933,N_13590);
xor U23254 (N_23254,N_13463,N_12352);
or U23255 (N_23255,N_16534,N_13477);
xor U23256 (N_23256,N_16913,N_17165);
xor U23257 (N_23257,N_16853,N_13226);
or U23258 (N_23258,N_16418,N_16842);
or U23259 (N_23259,N_15278,N_15836);
nand U23260 (N_23260,N_12268,N_12311);
and U23261 (N_23261,N_15411,N_17123);
nand U23262 (N_23262,N_13981,N_13439);
and U23263 (N_23263,N_12970,N_17984);
nand U23264 (N_23264,N_14311,N_16905);
or U23265 (N_23265,N_15722,N_17417);
xnor U23266 (N_23266,N_17314,N_17996);
nand U23267 (N_23267,N_16346,N_16004);
nor U23268 (N_23268,N_17769,N_15723);
nand U23269 (N_23269,N_16538,N_17967);
nor U23270 (N_23270,N_17592,N_15262);
nand U23271 (N_23271,N_12543,N_13068);
and U23272 (N_23272,N_12595,N_16886);
xnor U23273 (N_23273,N_12853,N_16120);
nand U23274 (N_23274,N_13426,N_12286);
nand U23275 (N_23275,N_12584,N_15315);
and U23276 (N_23276,N_12269,N_16350);
nor U23277 (N_23277,N_13672,N_17777);
xor U23278 (N_23278,N_17262,N_16873);
nand U23279 (N_23279,N_14305,N_17080);
xnor U23280 (N_23280,N_17975,N_16800);
xnor U23281 (N_23281,N_15898,N_13434);
and U23282 (N_23282,N_12034,N_12015);
and U23283 (N_23283,N_14856,N_16107);
nor U23284 (N_23284,N_16960,N_14669);
and U23285 (N_23285,N_12624,N_16310);
and U23286 (N_23286,N_13439,N_14330);
or U23287 (N_23287,N_14946,N_14405);
and U23288 (N_23288,N_17375,N_17823);
or U23289 (N_23289,N_16172,N_16651);
xnor U23290 (N_23290,N_17853,N_13928);
nand U23291 (N_23291,N_16865,N_12180);
or U23292 (N_23292,N_13116,N_12822);
and U23293 (N_23293,N_14877,N_12413);
and U23294 (N_23294,N_13930,N_14764);
and U23295 (N_23295,N_17320,N_17861);
nand U23296 (N_23296,N_17659,N_15297);
and U23297 (N_23297,N_13778,N_16526);
and U23298 (N_23298,N_14581,N_16340);
or U23299 (N_23299,N_13902,N_15251);
nor U23300 (N_23300,N_14124,N_12136);
and U23301 (N_23301,N_15639,N_12870);
and U23302 (N_23302,N_14971,N_12539);
and U23303 (N_23303,N_13497,N_16142);
and U23304 (N_23304,N_16958,N_15514);
or U23305 (N_23305,N_16920,N_12188);
or U23306 (N_23306,N_17030,N_14587);
nor U23307 (N_23307,N_12374,N_13891);
nand U23308 (N_23308,N_16265,N_16425);
or U23309 (N_23309,N_14190,N_15964);
xnor U23310 (N_23310,N_12055,N_14795);
xnor U23311 (N_23311,N_13877,N_17259);
nand U23312 (N_23312,N_13845,N_16643);
xor U23313 (N_23313,N_15951,N_16726);
nor U23314 (N_23314,N_12188,N_15758);
xor U23315 (N_23315,N_12197,N_15338);
nor U23316 (N_23316,N_13886,N_14942);
and U23317 (N_23317,N_12059,N_15135);
nand U23318 (N_23318,N_16567,N_13888);
or U23319 (N_23319,N_14735,N_14484);
nor U23320 (N_23320,N_13398,N_14272);
xor U23321 (N_23321,N_17973,N_16771);
nand U23322 (N_23322,N_13527,N_17531);
or U23323 (N_23323,N_13643,N_13087);
and U23324 (N_23324,N_14381,N_15417);
or U23325 (N_23325,N_12468,N_17732);
or U23326 (N_23326,N_17482,N_17764);
or U23327 (N_23327,N_16593,N_12828);
nand U23328 (N_23328,N_15446,N_13299);
nand U23329 (N_23329,N_16365,N_16742);
nand U23330 (N_23330,N_13143,N_17409);
and U23331 (N_23331,N_12370,N_16128);
and U23332 (N_23332,N_17469,N_13279);
or U23333 (N_23333,N_16105,N_14813);
and U23334 (N_23334,N_12961,N_15101);
xor U23335 (N_23335,N_15367,N_15652);
nor U23336 (N_23336,N_12363,N_14326);
nand U23337 (N_23337,N_13314,N_16891);
xor U23338 (N_23338,N_12695,N_15877);
and U23339 (N_23339,N_12329,N_16849);
xor U23340 (N_23340,N_15415,N_14337);
nor U23341 (N_23341,N_17190,N_13362);
nand U23342 (N_23342,N_14254,N_17468);
nor U23343 (N_23343,N_17381,N_13268);
nor U23344 (N_23344,N_16526,N_15905);
xor U23345 (N_23345,N_15525,N_15794);
nand U23346 (N_23346,N_12424,N_17178);
or U23347 (N_23347,N_15379,N_12108);
or U23348 (N_23348,N_14544,N_16507);
nor U23349 (N_23349,N_14260,N_16058);
xnor U23350 (N_23350,N_12803,N_12233);
or U23351 (N_23351,N_13982,N_15587);
and U23352 (N_23352,N_17042,N_17881);
and U23353 (N_23353,N_16543,N_15543);
xor U23354 (N_23354,N_15679,N_13657);
nor U23355 (N_23355,N_12285,N_17413);
nor U23356 (N_23356,N_16697,N_16768);
xnor U23357 (N_23357,N_13173,N_14863);
xnor U23358 (N_23358,N_14112,N_12325);
or U23359 (N_23359,N_12719,N_16911);
xor U23360 (N_23360,N_17925,N_17169);
and U23361 (N_23361,N_12387,N_14748);
and U23362 (N_23362,N_13127,N_17510);
nand U23363 (N_23363,N_15581,N_12979);
and U23364 (N_23364,N_13210,N_12724);
nand U23365 (N_23365,N_12819,N_15227);
xnor U23366 (N_23366,N_13448,N_15799);
or U23367 (N_23367,N_15096,N_12439);
nand U23368 (N_23368,N_17237,N_17318);
and U23369 (N_23369,N_16080,N_16814);
xor U23370 (N_23370,N_12166,N_13295);
and U23371 (N_23371,N_14442,N_12672);
or U23372 (N_23372,N_15970,N_14172);
or U23373 (N_23373,N_17105,N_12961);
nor U23374 (N_23374,N_14323,N_12971);
or U23375 (N_23375,N_15635,N_16868);
and U23376 (N_23376,N_14468,N_13606);
or U23377 (N_23377,N_15761,N_17652);
and U23378 (N_23378,N_16887,N_15017);
nand U23379 (N_23379,N_17557,N_16064);
nand U23380 (N_23380,N_13326,N_15494);
nor U23381 (N_23381,N_14365,N_17886);
xnor U23382 (N_23382,N_14209,N_17464);
nor U23383 (N_23383,N_14086,N_16813);
nand U23384 (N_23384,N_14335,N_13792);
and U23385 (N_23385,N_16533,N_16126);
nor U23386 (N_23386,N_17778,N_13919);
nor U23387 (N_23387,N_14849,N_17052);
nor U23388 (N_23388,N_16030,N_12912);
xor U23389 (N_23389,N_17102,N_17849);
xnor U23390 (N_23390,N_14344,N_14541);
and U23391 (N_23391,N_15027,N_15487);
nor U23392 (N_23392,N_12877,N_13469);
nor U23393 (N_23393,N_12449,N_15639);
or U23394 (N_23394,N_16030,N_13686);
nor U23395 (N_23395,N_14049,N_16986);
xnor U23396 (N_23396,N_14625,N_16642);
or U23397 (N_23397,N_14269,N_13507);
nor U23398 (N_23398,N_13982,N_13114);
nor U23399 (N_23399,N_12079,N_16327);
and U23400 (N_23400,N_12036,N_12353);
or U23401 (N_23401,N_13285,N_17016);
or U23402 (N_23402,N_17914,N_16331);
and U23403 (N_23403,N_13875,N_14173);
or U23404 (N_23404,N_16101,N_13561);
xnor U23405 (N_23405,N_13489,N_14961);
and U23406 (N_23406,N_13305,N_16895);
and U23407 (N_23407,N_17557,N_16495);
xnor U23408 (N_23408,N_12404,N_12810);
xor U23409 (N_23409,N_13807,N_12194);
nand U23410 (N_23410,N_12296,N_13131);
xor U23411 (N_23411,N_16957,N_12558);
and U23412 (N_23412,N_14456,N_17849);
xor U23413 (N_23413,N_15975,N_17822);
nor U23414 (N_23414,N_13511,N_13720);
and U23415 (N_23415,N_16707,N_12398);
xnor U23416 (N_23416,N_15503,N_12659);
xnor U23417 (N_23417,N_12538,N_16144);
xnor U23418 (N_23418,N_15097,N_13747);
xor U23419 (N_23419,N_17490,N_14742);
nor U23420 (N_23420,N_16863,N_17603);
nand U23421 (N_23421,N_17393,N_16378);
and U23422 (N_23422,N_13517,N_13091);
or U23423 (N_23423,N_16316,N_15031);
or U23424 (N_23424,N_17116,N_17336);
xnor U23425 (N_23425,N_15663,N_12819);
xor U23426 (N_23426,N_12481,N_13488);
and U23427 (N_23427,N_16884,N_12944);
nand U23428 (N_23428,N_12525,N_15514);
or U23429 (N_23429,N_13608,N_13809);
nor U23430 (N_23430,N_15501,N_13610);
or U23431 (N_23431,N_13316,N_14678);
nand U23432 (N_23432,N_12062,N_17612);
nor U23433 (N_23433,N_17742,N_14285);
xnor U23434 (N_23434,N_14339,N_12715);
or U23435 (N_23435,N_13439,N_17663);
xnor U23436 (N_23436,N_13618,N_15136);
or U23437 (N_23437,N_13902,N_14868);
or U23438 (N_23438,N_15074,N_17296);
and U23439 (N_23439,N_14055,N_14225);
nand U23440 (N_23440,N_16925,N_15722);
or U23441 (N_23441,N_13963,N_16808);
or U23442 (N_23442,N_17984,N_13062);
and U23443 (N_23443,N_14245,N_14700);
and U23444 (N_23444,N_17844,N_14437);
nand U23445 (N_23445,N_16438,N_17089);
or U23446 (N_23446,N_17345,N_15404);
xnor U23447 (N_23447,N_15970,N_17537);
nand U23448 (N_23448,N_14862,N_14437);
nand U23449 (N_23449,N_14187,N_14782);
xor U23450 (N_23450,N_14615,N_15152);
xnor U23451 (N_23451,N_14688,N_16588);
xor U23452 (N_23452,N_14825,N_17843);
and U23453 (N_23453,N_17164,N_14847);
nor U23454 (N_23454,N_15652,N_17315);
nor U23455 (N_23455,N_17389,N_13687);
xor U23456 (N_23456,N_16374,N_16005);
nand U23457 (N_23457,N_16811,N_17356);
or U23458 (N_23458,N_16554,N_15124);
xor U23459 (N_23459,N_16691,N_13131);
and U23460 (N_23460,N_12855,N_15996);
nand U23461 (N_23461,N_17046,N_12527);
nor U23462 (N_23462,N_13136,N_17695);
or U23463 (N_23463,N_12355,N_15805);
and U23464 (N_23464,N_16268,N_15469);
nand U23465 (N_23465,N_13902,N_15247);
xnor U23466 (N_23466,N_16937,N_17376);
nand U23467 (N_23467,N_14607,N_16509);
nand U23468 (N_23468,N_17222,N_15714);
and U23469 (N_23469,N_15858,N_13356);
and U23470 (N_23470,N_15969,N_14679);
nor U23471 (N_23471,N_12013,N_17869);
nor U23472 (N_23472,N_14774,N_16253);
and U23473 (N_23473,N_12254,N_15002);
or U23474 (N_23474,N_13579,N_13230);
nor U23475 (N_23475,N_12135,N_15266);
nand U23476 (N_23476,N_15465,N_13737);
and U23477 (N_23477,N_12162,N_17070);
xnor U23478 (N_23478,N_15247,N_17607);
nor U23479 (N_23479,N_17909,N_15838);
nand U23480 (N_23480,N_13817,N_13312);
nor U23481 (N_23481,N_17386,N_13141);
and U23482 (N_23482,N_12784,N_17464);
and U23483 (N_23483,N_17853,N_16778);
nand U23484 (N_23484,N_17122,N_12973);
xnor U23485 (N_23485,N_15711,N_17986);
nand U23486 (N_23486,N_13076,N_12400);
nand U23487 (N_23487,N_12816,N_14616);
nor U23488 (N_23488,N_17453,N_16838);
xor U23489 (N_23489,N_12476,N_13811);
and U23490 (N_23490,N_17504,N_16035);
nor U23491 (N_23491,N_12661,N_17024);
or U23492 (N_23492,N_14194,N_15039);
nand U23493 (N_23493,N_12596,N_13738);
or U23494 (N_23494,N_12973,N_17539);
nor U23495 (N_23495,N_15263,N_15874);
or U23496 (N_23496,N_17838,N_12223);
and U23497 (N_23497,N_16759,N_15472);
or U23498 (N_23498,N_12915,N_15820);
nor U23499 (N_23499,N_16381,N_16198);
or U23500 (N_23500,N_17936,N_12076);
and U23501 (N_23501,N_13511,N_17424);
nand U23502 (N_23502,N_16747,N_17924);
and U23503 (N_23503,N_14445,N_16956);
and U23504 (N_23504,N_15188,N_17658);
nor U23505 (N_23505,N_14859,N_13874);
xnor U23506 (N_23506,N_17717,N_16578);
or U23507 (N_23507,N_12908,N_16382);
nand U23508 (N_23508,N_15780,N_12365);
or U23509 (N_23509,N_15004,N_14271);
nand U23510 (N_23510,N_14095,N_14677);
or U23511 (N_23511,N_15174,N_13620);
xor U23512 (N_23512,N_14158,N_15838);
nand U23513 (N_23513,N_12108,N_16321);
nor U23514 (N_23514,N_14226,N_16744);
nand U23515 (N_23515,N_17863,N_17561);
or U23516 (N_23516,N_15827,N_17287);
nor U23517 (N_23517,N_15675,N_13121);
nand U23518 (N_23518,N_17555,N_16648);
xor U23519 (N_23519,N_13656,N_16192);
or U23520 (N_23520,N_17988,N_17597);
nand U23521 (N_23521,N_14553,N_13709);
xnor U23522 (N_23522,N_14180,N_12677);
nor U23523 (N_23523,N_15966,N_13213);
and U23524 (N_23524,N_12747,N_16661);
xnor U23525 (N_23525,N_14258,N_12402);
xor U23526 (N_23526,N_17599,N_14248);
nand U23527 (N_23527,N_15288,N_13851);
nor U23528 (N_23528,N_15524,N_17413);
or U23529 (N_23529,N_17688,N_17864);
and U23530 (N_23530,N_16083,N_16839);
xnor U23531 (N_23531,N_16402,N_14792);
xor U23532 (N_23532,N_12390,N_16505);
xor U23533 (N_23533,N_16884,N_17524);
and U23534 (N_23534,N_14319,N_12559);
xnor U23535 (N_23535,N_12292,N_15696);
and U23536 (N_23536,N_14513,N_17101);
or U23537 (N_23537,N_17775,N_15904);
nand U23538 (N_23538,N_14896,N_13210);
and U23539 (N_23539,N_14972,N_15176);
or U23540 (N_23540,N_16070,N_17509);
and U23541 (N_23541,N_12196,N_13288);
nor U23542 (N_23542,N_16674,N_16252);
xor U23543 (N_23543,N_13334,N_13644);
or U23544 (N_23544,N_16950,N_16570);
nand U23545 (N_23545,N_13197,N_12579);
xor U23546 (N_23546,N_15660,N_12510);
or U23547 (N_23547,N_16721,N_17766);
xor U23548 (N_23548,N_16189,N_12361);
nor U23549 (N_23549,N_12753,N_15633);
and U23550 (N_23550,N_16533,N_12492);
nor U23551 (N_23551,N_17337,N_14981);
nand U23552 (N_23552,N_16156,N_16976);
or U23553 (N_23553,N_16980,N_12318);
nand U23554 (N_23554,N_13099,N_15801);
nand U23555 (N_23555,N_16856,N_16867);
and U23556 (N_23556,N_15675,N_17116);
and U23557 (N_23557,N_15097,N_12998);
and U23558 (N_23558,N_12846,N_14827);
and U23559 (N_23559,N_12877,N_13666);
nand U23560 (N_23560,N_14155,N_17003);
or U23561 (N_23561,N_15966,N_14272);
nor U23562 (N_23562,N_13740,N_13553);
xnor U23563 (N_23563,N_16273,N_16431);
xor U23564 (N_23564,N_14750,N_15645);
nand U23565 (N_23565,N_16499,N_17844);
nand U23566 (N_23566,N_12123,N_17274);
nand U23567 (N_23567,N_14384,N_13210);
or U23568 (N_23568,N_13176,N_15335);
nand U23569 (N_23569,N_16545,N_12018);
or U23570 (N_23570,N_14947,N_14919);
nor U23571 (N_23571,N_12662,N_12031);
or U23572 (N_23572,N_14803,N_12915);
or U23573 (N_23573,N_17730,N_16928);
nor U23574 (N_23574,N_15251,N_12279);
or U23575 (N_23575,N_16056,N_13697);
or U23576 (N_23576,N_16128,N_14476);
nand U23577 (N_23577,N_15603,N_14724);
or U23578 (N_23578,N_12999,N_16154);
xor U23579 (N_23579,N_12389,N_16477);
and U23580 (N_23580,N_16184,N_13741);
xor U23581 (N_23581,N_14136,N_17714);
nor U23582 (N_23582,N_16964,N_16649);
and U23583 (N_23583,N_17306,N_17658);
and U23584 (N_23584,N_16237,N_15675);
nor U23585 (N_23585,N_14674,N_14768);
or U23586 (N_23586,N_15190,N_13618);
xnor U23587 (N_23587,N_14523,N_12094);
nand U23588 (N_23588,N_16297,N_13123);
or U23589 (N_23589,N_15874,N_17752);
nor U23590 (N_23590,N_16627,N_13117);
and U23591 (N_23591,N_14891,N_13478);
or U23592 (N_23592,N_13082,N_13432);
nor U23593 (N_23593,N_15584,N_12134);
xnor U23594 (N_23594,N_15774,N_15396);
nor U23595 (N_23595,N_16195,N_16918);
nor U23596 (N_23596,N_14108,N_17462);
nor U23597 (N_23597,N_13272,N_17035);
xnor U23598 (N_23598,N_12204,N_12517);
nand U23599 (N_23599,N_13478,N_17695);
or U23600 (N_23600,N_15332,N_13173);
or U23601 (N_23601,N_17078,N_14999);
and U23602 (N_23602,N_15794,N_16275);
nor U23603 (N_23603,N_12237,N_15987);
and U23604 (N_23604,N_14487,N_13179);
or U23605 (N_23605,N_13341,N_12961);
xnor U23606 (N_23606,N_17241,N_15380);
nand U23607 (N_23607,N_17487,N_13290);
nand U23608 (N_23608,N_12431,N_16712);
nand U23609 (N_23609,N_14108,N_16448);
xor U23610 (N_23610,N_16815,N_14736);
or U23611 (N_23611,N_14460,N_13525);
and U23612 (N_23612,N_12445,N_13943);
nand U23613 (N_23613,N_17174,N_12723);
or U23614 (N_23614,N_17018,N_14521);
xor U23615 (N_23615,N_15921,N_14828);
xnor U23616 (N_23616,N_15883,N_16487);
or U23617 (N_23617,N_16285,N_16923);
nor U23618 (N_23618,N_14149,N_13251);
nor U23619 (N_23619,N_13388,N_17976);
or U23620 (N_23620,N_17509,N_14686);
and U23621 (N_23621,N_12199,N_16839);
and U23622 (N_23622,N_17968,N_15946);
and U23623 (N_23623,N_13648,N_16525);
or U23624 (N_23624,N_12948,N_17661);
or U23625 (N_23625,N_15454,N_16821);
nor U23626 (N_23626,N_12339,N_12713);
xor U23627 (N_23627,N_17709,N_14858);
nor U23628 (N_23628,N_12292,N_16587);
nand U23629 (N_23629,N_15763,N_13694);
or U23630 (N_23630,N_13016,N_17096);
xor U23631 (N_23631,N_13293,N_12286);
xnor U23632 (N_23632,N_13053,N_12426);
xnor U23633 (N_23633,N_13298,N_16472);
nor U23634 (N_23634,N_16037,N_17975);
nand U23635 (N_23635,N_15176,N_14373);
xor U23636 (N_23636,N_14072,N_14530);
and U23637 (N_23637,N_13938,N_16095);
or U23638 (N_23638,N_14281,N_13331);
xnor U23639 (N_23639,N_17097,N_17456);
nor U23640 (N_23640,N_13619,N_14946);
nand U23641 (N_23641,N_17923,N_13246);
nor U23642 (N_23642,N_12492,N_15901);
or U23643 (N_23643,N_13531,N_12703);
nand U23644 (N_23644,N_17485,N_13079);
and U23645 (N_23645,N_15317,N_12464);
nor U23646 (N_23646,N_13401,N_14197);
nand U23647 (N_23647,N_17922,N_14288);
or U23648 (N_23648,N_14900,N_17541);
or U23649 (N_23649,N_17894,N_14446);
and U23650 (N_23650,N_13455,N_13310);
and U23651 (N_23651,N_15787,N_16157);
nand U23652 (N_23652,N_13964,N_14537);
xor U23653 (N_23653,N_15729,N_12556);
or U23654 (N_23654,N_14456,N_17693);
nand U23655 (N_23655,N_15150,N_14865);
xor U23656 (N_23656,N_16176,N_16109);
nand U23657 (N_23657,N_14962,N_17860);
or U23658 (N_23658,N_17770,N_12937);
xnor U23659 (N_23659,N_13926,N_13536);
nor U23660 (N_23660,N_13202,N_13286);
nor U23661 (N_23661,N_17072,N_13055);
or U23662 (N_23662,N_12619,N_15047);
or U23663 (N_23663,N_12677,N_16320);
or U23664 (N_23664,N_13224,N_16621);
nand U23665 (N_23665,N_12688,N_14381);
xor U23666 (N_23666,N_12758,N_13752);
and U23667 (N_23667,N_14991,N_14094);
nand U23668 (N_23668,N_12595,N_17142);
xor U23669 (N_23669,N_12887,N_16133);
nor U23670 (N_23670,N_13130,N_12924);
or U23671 (N_23671,N_12614,N_16587);
or U23672 (N_23672,N_12535,N_13405);
or U23673 (N_23673,N_16478,N_16805);
or U23674 (N_23674,N_13396,N_16202);
nor U23675 (N_23675,N_15339,N_15601);
or U23676 (N_23676,N_12524,N_12768);
xor U23677 (N_23677,N_15222,N_12626);
and U23678 (N_23678,N_14472,N_15906);
and U23679 (N_23679,N_13179,N_15144);
or U23680 (N_23680,N_16342,N_16901);
xor U23681 (N_23681,N_15170,N_13623);
nand U23682 (N_23682,N_13340,N_12569);
or U23683 (N_23683,N_13199,N_17415);
or U23684 (N_23684,N_13206,N_15758);
xnor U23685 (N_23685,N_15779,N_15794);
and U23686 (N_23686,N_14079,N_14353);
nand U23687 (N_23687,N_17664,N_14396);
nand U23688 (N_23688,N_12193,N_17620);
nand U23689 (N_23689,N_16615,N_16334);
nand U23690 (N_23690,N_13200,N_16923);
xnor U23691 (N_23691,N_12703,N_12213);
nand U23692 (N_23692,N_17822,N_17376);
and U23693 (N_23693,N_16414,N_12422);
nand U23694 (N_23694,N_14484,N_12021);
xor U23695 (N_23695,N_15130,N_12718);
nand U23696 (N_23696,N_13956,N_14798);
nand U23697 (N_23697,N_12933,N_16486);
and U23698 (N_23698,N_13518,N_12249);
xnor U23699 (N_23699,N_17473,N_13924);
and U23700 (N_23700,N_14219,N_16729);
nor U23701 (N_23701,N_15547,N_15486);
or U23702 (N_23702,N_14567,N_17523);
and U23703 (N_23703,N_13181,N_17954);
and U23704 (N_23704,N_12599,N_16469);
or U23705 (N_23705,N_15402,N_14359);
nor U23706 (N_23706,N_15527,N_13363);
xor U23707 (N_23707,N_14293,N_16015);
or U23708 (N_23708,N_17887,N_16932);
nor U23709 (N_23709,N_12313,N_17231);
or U23710 (N_23710,N_16346,N_16910);
and U23711 (N_23711,N_13530,N_15147);
or U23712 (N_23712,N_14209,N_16663);
nand U23713 (N_23713,N_16484,N_17110);
and U23714 (N_23714,N_12729,N_14918);
nand U23715 (N_23715,N_15065,N_16006);
nand U23716 (N_23716,N_12031,N_14556);
and U23717 (N_23717,N_16346,N_14793);
and U23718 (N_23718,N_14247,N_15790);
xnor U23719 (N_23719,N_13334,N_17762);
nand U23720 (N_23720,N_14423,N_13757);
nor U23721 (N_23721,N_16255,N_12564);
nand U23722 (N_23722,N_14903,N_15351);
nor U23723 (N_23723,N_12565,N_16135);
or U23724 (N_23724,N_15824,N_12386);
or U23725 (N_23725,N_13269,N_15702);
nand U23726 (N_23726,N_12815,N_13274);
nand U23727 (N_23727,N_15676,N_15155);
xor U23728 (N_23728,N_14347,N_17369);
nor U23729 (N_23729,N_15402,N_13104);
xor U23730 (N_23730,N_14707,N_12018);
nand U23731 (N_23731,N_16949,N_12949);
nand U23732 (N_23732,N_14572,N_17629);
nand U23733 (N_23733,N_12101,N_12795);
and U23734 (N_23734,N_16489,N_12219);
nand U23735 (N_23735,N_15615,N_12403);
xor U23736 (N_23736,N_17869,N_12124);
xnor U23737 (N_23737,N_16561,N_15285);
and U23738 (N_23738,N_15267,N_16887);
nand U23739 (N_23739,N_14662,N_17552);
nor U23740 (N_23740,N_17020,N_12421);
or U23741 (N_23741,N_16326,N_14391);
xor U23742 (N_23742,N_15350,N_12911);
nand U23743 (N_23743,N_14852,N_14758);
xor U23744 (N_23744,N_15061,N_15756);
nand U23745 (N_23745,N_12751,N_13371);
nand U23746 (N_23746,N_17644,N_14017);
or U23747 (N_23747,N_17532,N_14715);
and U23748 (N_23748,N_13653,N_15414);
or U23749 (N_23749,N_15547,N_13058);
nand U23750 (N_23750,N_17601,N_15325);
xor U23751 (N_23751,N_13282,N_13561);
nor U23752 (N_23752,N_12797,N_16203);
nor U23753 (N_23753,N_14822,N_15213);
xnor U23754 (N_23754,N_12496,N_14961);
nor U23755 (N_23755,N_13763,N_14860);
xnor U23756 (N_23756,N_13996,N_14157);
and U23757 (N_23757,N_17147,N_13080);
nor U23758 (N_23758,N_17204,N_16585);
nor U23759 (N_23759,N_15614,N_14102);
nor U23760 (N_23760,N_13843,N_14452);
nor U23761 (N_23761,N_16187,N_17911);
and U23762 (N_23762,N_12941,N_14706);
or U23763 (N_23763,N_13037,N_12392);
nand U23764 (N_23764,N_16454,N_13339);
or U23765 (N_23765,N_16279,N_16756);
nand U23766 (N_23766,N_16059,N_15682);
nand U23767 (N_23767,N_14811,N_12080);
nand U23768 (N_23768,N_17127,N_12751);
or U23769 (N_23769,N_12584,N_16166);
nand U23770 (N_23770,N_14025,N_16688);
nor U23771 (N_23771,N_16806,N_13205);
xnor U23772 (N_23772,N_17757,N_17793);
or U23773 (N_23773,N_14204,N_13630);
nand U23774 (N_23774,N_12916,N_17036);
nor U23775 (N_23775,N_14934,N_16761);
or U23776 (N_23776,N_14498,N_17822);
and U23777 (N_23777,N_14544,N_14862);
or U23778 (N_23778,N_13653,N_15793);
nand U23779 (N_23779,N_15066,N_14805);
nand U23780 (N_23780,N_15689,N_15986);
or U23781 (N_23781,N_12469,N_14846);
xor U23782 (N_23782,N_15286,N_13445);
and U23783 (N_23783,N_15780,N_13795);
xnor U23784 (N_23784,N_16084,N_12664);
or U23785 (N_23785,N_14671,N_16781);
nor U23786 (N_23786,N_17611,N_13222);
and U23787 (N_23787,N_17848,N_12458);
and U23788 (N_23788,N_17013,N_13449);
nor U23789 (N_23789,N_17982,N_13727);
or U23790 (N_23790,N_14437,N_12845);
and U23791 (N_23791,N_14888,N_16884);
nor U23792 (N_23792,N_13759,N_14822);
xnor U23793 (N_23793,N_13360,N_12774);
and U23794 (N_23794,N_17052,N_12102);
xor U23795 (N_23795,N_13485,N_15985);
xor U23796 (N_23796,N_14077,N_17935);
and U23797 (N_23797,N_16776,N_17423);
and U23798 (N_23798,N_16346,N_17995);
nand U23799 (N_23799,N_16703,N_13622);
or U23800 (N_23800,N_16636,N_16292);
or U23801 (N_23801,N_13894,N_12925);
xor U23802 (N_23802,N_14084,N_13088);
and U23803 (N_23803,N_13361,N_13504);
nor U23804 (N_23804,N_13262,N_15217);
or U23805 (N_23805,N_12557,N_15975);
xnor U23806 (N_23806,N_16734,N_14408);
nor U23807 (N_23807,N_14759,N_13782);
xnor U23808 (N_23808,N_17053,N_17110);
nand U23809 (N_23809,N_14428,N_13222);
nand U23810 (N_23810,N_13120,N_17465);
or U23811 (N_23811,N_16598,N_14290);
and U23812 (N_23812,N_14570,N_15193);
or U23813 (N_23813,N_16789,N_15499);
or U23814 (N_23814,N_13452,N_16399);
xor U23815 (N_23815,N_12841,N_12017);
or U23816 (N_23816,N_12142,N_12520);
and U23817 (N_23817,N_17905,N_13991);
and U23818 (N_23818,N_14774,N_14351);
or U23819 (N_23819,N_12660,N_14854);
nor U23820 (N_23820,N_13939,N_14825);
nor U23821 (N_23821,N_13116,N_16464);
and U23822 (N_23822,N_12746,N_12544);
nand U23823 (N_23823,N_13957,N_12859);
nand U23824 (N_23824,N_17009,N_14545);
nor U23825 (N_23825,N_16249,N_13280);
nand U23826 (N_23826,N_14063,N_17926);
or U23827 (N_23827,N_17071,N_14208);
or U23828 (N_23828,N_17332,N_15507);
nor U23829 (N_23829,N_16245,N_13981);
nor U23830 (N_23830,N_17768,N_12946);
nand U23831 (N_23831,N_15545,N_17079);
or U23832 (N_23832,N_17507,N_12337);
nor U23833 (N_23833,N_13625,N_12797);
nor U23834 (N_23834,N_15309,N_15813);
nand U23835 (N_23835,N_15453,N_15799);
and U23836 (N_23836,N_17256,N_16541);
nor U23837 (N_23837,N_13491,N_14172);
nand U23838 (N_23838,N_14735,N_16960);
or U23839 (N_23839,N_12274,N_16650);
nand U23840 (N_23840,N_15893,N_12799);
or U23841 (N_23841,N_12252,N_12745);
xnor U23842 (N_23842,N_15320,N_16696);
nand U23843 (N_23843,N_17881,N_17559);
or U23844 (N_23844,N_12265,N_16307);
nor U23845 (N_23845,N_14402,N_15969);
or U23846 (N_23846,N_15438,N_14083);
and U23847 (N_23847,N_17141,N_13818);
nand U23848 (N_23848,N_12844,N_14490);
or U23849 (N_23849,N_16134,N_15894);
nor U23850 (N_23850,N_15445,N_17118);
nand U23851 (N_23851,N_16329,N_17483);
or U23852 (N_23852,N_14171,N_12391);
xor U23853 (N_23853,N_16661,N_12616);
nand U23854 (N_23854,N_13926,N_17214);
xor U23855 (N_23855,N_14996,N_14032);
or U23856 (N_23856,N_14891,N_16950);
or U23857 (N_23857,N_15546,N_15176);
or U23858 (N_23858,N_14680,N_16666);
and U23859 (N_23859,N_16782,N_15720);
nor U23860 (N_23860,N_15761,N_15977);
xnor U23861 (N_23861,N_13198,N_16079);
or U23862 (N_23862,N_17459,N_14545);
xnor U23863 (N_23863,N_15550,N_14093);
or U23864 (N_23864,N_12972,N_13811);
xnor U23865 (N_23865,N_13852,N_12624);
and U23866 (N_23866,N_15896,N_13882);
nand U23867 (N_23867,N_13009,N_12707);
xnor U23868 (N_23868,N_12853,N_14614);
and U23869 (N_23869,N_16012,N_12840);
or U23870 (N_23870,N_15660,N_12556);
nor U23871 (N_23871,N_15525,N_17497);
nor U23872 (N_23872,N_14097,N_13108);
and U23873 (N_23873,N_14992,N_14537);
nand U23874 (N_23874,N_15198,N_17125);
nor U23875 (N_23875,N_17366,N_12546);
xor U23876 (N_23876,N_13593,N_14294);
nand U23877 (N_23877,N_16693,N_12796);
and U23878 (N_23878,N_12138,N_14091);
xnor U23879 (N_23879,N_15286,N_15168);
or U23880 (N_23880,N_15414,N_14273);
nor U23881 (N_23881,N_12944,N_12731);
and U23882 (N_23882,N_16451,N_16417);
nor U23883 (N_23883,N_15614,N_15075);
or U23884 (N_23884,N_13816,N_17799);
or U23885 (N_23885,N_17397,N_16647);
nor U23886 (N_23886,N_14347,N_15849);
nor U23887 (N_23887,N_12559,N_14743);
xor U23888 (N_23888,N_13391,N_14043);
xor U23889 (N_23889,N_15841,N_15461);
xor U23890 (N_23890,N_12033,N_13582);
or U23891 (N_23891,N_15977,N_15060);
and U23892 (N_23892,N_13700,N_17292);
and U23893 (N_23893,N_15664,N_15970);
xor U23894 (N_23894,N_14631,N_13672);
and U23895 (N_23895,N_15773,N_15718);
nor U23896 (N_23896,N_15246,N_13388);
and U23897 (N_23897,N_14753,N_12340);
xor U23898 (N_23898,N_16234,N_13865);
and U23899 (N_23899,N_13578,N_13874);
and U23900 (N_23900,N_12037,N_16196);
and U23901 (N_23901,N_12379,N_15030);
nand U23902 (N_23902,N_16156,N_16266);
or U23903 (N_23903,N_17349,N_17091);
and U23904 (N_23904,N_17329,N_16023);
nor U23905 (N_23905,N_12475,N_13320);
nor U23906 (N_23906,N_14200,N_15443);
or U23907 (N_23907,N_12935,N_14883);
or U23908 (N_23908,N_16977,N_14596);
or U23909 (N_23909,N_16345,N_17873);
or U23910 (N_23910,N_17406,N_15909);
and U23911 (N_23911,N_13967,N_17375);
and U23912 (N_23912,N_16257,N_12867);
and U23913 (N_23913,N_12462,N_12298);
xor U23914 (N_23914,N_15644,N_16568);
nor U23915 (N_23915,N_15815,N_17616);
or U23916 (N_23916,N_16135,N_12736);
nand U23917 (N_23917,N_15050,N_16549);
or U23918 (N_23918,N_15290,N_17626);
nor U23919 (N_23919,N_15890,N_13328);
nor U23920 (N_23920,N_16347,N_12604);
nand U23921 (N_23921,N_14564,N_17794);
or U23922 (N_23922,N_17085,N_13880);
nor U23923 (N_23923,N_16797,N_16813);
or U23924 (N_23924,N_17144,N_12379);
nor U23925 (N_23925,N_13750,N_14954);
xnor U23926 (N_23926,N_13943,N_17738);
or U23927 (N_23927,N_13402,N_17584);
or U23928 (N_23928,N_13430,N_14416);
or U23929 (N_23929,N_17160,N_13836);
or U23930 (N_23930,N_16917,N_14836);
xnor U23931 (N_23931,N_14756,N_16497);
xnor U23932 (N_23932,N_12917,N_13822);
and U23933 (N_23933,N_14785,N_13089);
and U23934 (N_23934,N_15559,N_15558);
nand U23935 (N_23935,N_12082,N_17627);
nand U23936 (N_23936,N_16588,N_14891);
nor U23937 (N_23937,N_12978,N_14325);
nand U23938 (N_23938,N_13295,N_17064);
xor U23939 (N_23939,N_16689,N_13572);
and U23940 (N_23940,N_12813,N_13306);
and U23941 (N_23941,N_12127,N_12502);
xnor U23942 (N_23942,N_15931,N_14865);
nand U23943 (N_23943,N_15097,N_17115);
or U23944 (N_23944,N_17226,N_12645);
nor U23945 (N_23945,N_15953,N_17177);
nand U23946 (N_23946,N_15012,N_15383);
xor U23947 (N_23947,N_12943,N_14625);
nor U23948 (N_23948,N_14540,N_13554);
or U23949 (N_23949,N_17696,N_15645);
or U23950 (N_23950,N_16640,N_17363);
or U23951 (N_23951,N_14871,N_17721);
and U23952 (N_23952,N_13082,N_15884);
nor U23953 (N_23953,N_16093,N_15528);
nand U23954 (N_23954,N_12717,N_15314);
or U23955 (N_23955,N_13395,N_13821);
xnor U23956 (N_23956,N_13107,N_15295);
nor U23957 (N_23957,N_13724,N_17688);
or U23958 (N_23958,N_13176,N_16635);
nor U23959 (N_23959,N_14563,N_16346);
or U23960 (N_23960,N_17297,N_16831);
or U23961 (N_23961,N_14590,N_13640);
nand U23962 (N_23962,N_13516,N_12005);
nor U23963 (N_23963,N_14650,N_16332);
or U23964 (N_23964,N_15740,N_15876);
and U23965 (N_23965,N_13588,N_17448);
nand U23966 (N_23966,N_13161,N_16405);
and U23967 (N_23967,N_13332,N_12137);
or U23968 (N_23968,N_13190,N_17909);
xor U23969 (N_23969,N_15239,N_15883);
nor U23970 (N_23970,N_16039,N_14390);
nand U23971 (N_23971,N_17266,N_16202);
xor U23972 (N_23972,N_12231,N_14250);
and U23973 (N_23973,N_12848,N_13546);
and U23974 (N_23974,N_15102,N_14526);
and U23975 (N_23975,N_12994,N_14651);
nor U23976 (N_23976,N_14400,N_15222);
xnor U23977 (N_23977,N_15069,N_14975);
and U23978 (N_23978,N_12913,N_14276);
nand U23979 (N_23979,N_13586,N_16868);
nor U23980 (N_23980,N_16339,N_17874);
and U23981 (N_23981,N_17588,N_13909);
and U23982 (N_23982,N_14362,N_13042);
nand U23983 (N_23983,N_17945,N_15781);
and U23984 (N_23984,N_14630,N_13014);
nor U23985 (N_23985,N_15042,N_16744);
or U23986 (N_23986,N_17804,N_13265);
nand U23987 (N_23987,N_17590,N_16262);
nor U23988 (N_23988,N_14730,N_17056);
or U23989 (N_23989,N_15100,N_15516);
or U23990 (N_23990,N_13179,N_12385);
nand U23991 (N_23991,N_16514,N_16569);
nand U23992 (N_23992,N_17675,N_14498);
or U23993 (N_23993,N_14673,N_16268);
xnor U23994 (N_23994,N_15982,N_13573);
or U23995 (N_23995,N_12659,N_12495);
xor U23996 (N_23996,N_13167,N_13813);
nor U23997 (N_23997,N_14989,N_14705);
nand U23998 (N_23998,N_13175,N_12490);
and U23999 (N_23999,N_17546,N_13751);
nand U24000 (N_24000,N_18706,N_22486);
and U24001 (N_24001,N_20016,N_23718);
and U24002 (N_24002,N_20900,N_20702);
or U24003 (N_24003,N_23008,N_23181);
nand U24004 (N_24004,N_19414,N_22570);
or U24005 (N_24005,N_22099,N_22635);
or U24006 (N_24006,N_22840,N_23986);
xor U24007 (N_24007,N_23442,N_19478);
nand U24008 (N_24008,N_20932,N_20278);
nand U24009 (N_24009,N_20110,N_19546);
xor U24010 (N_24010,N_23599,N_20600);
nand U24011 (N_24011,N_22980,N_19244);
and U24012 (N_24012,N_19079,N_23713);
nor U24013 (N_24013,N_18530,N_21875);
xor U24014 (N_24014,N_20248,N_21074);
nor U24015 (N_24015,N_19234,N_18463);
nor U24016 (N_24016,N_22675,N_23731);
and U24017 (N_24017,N_20700,N_19967);
nor U24018 (N_24018,N_22030,N_21424);
nand U24019 (N_24019,N_21646,N_19831);
and U24020 (N_24020,N_23628,N_20586);
or U24021 (N_24021,N_19773,N_23434);
nor U24022 (N_24022,N_23423,N_22159);
and U24023 (N_24023,N_20670,N_19516);
xnor U24024 (N_24024,N_22390,N_21033);
or U24025 (N_24025,N_20575,N_21671);
nor U24026 (N_24026,N_19371,N_23418);
or U24027 (N_24027,N_23488,N_18562);
and U24028 (N_24028,N_21075,N_19986);
or U24029 (N_24029,N_23946,N_19577);
or U24030 (N_24030,N_18435,N_18039);
nand U24031 (N_24031,N_20273,N_18479);
nand U24032 (N_24032,N_19570,N_22612);
and U24033 (N_24033,N_22291,N_21821);
or U24034 (N_24034,N_19131,N_23658);
xor U24035 (N_24035,N_21307,N_18174);
xnor U24036 (N_24036,N_20287,N_22445);
xnor U24037 (N_24037,N_20719,N_23023);
or U24038 (N_24038,N_22845,N_23825);
or U24039 (N_24039,N_20406,N_18887);
nor U24040 (N_24040,N_23426,N_23154);
and U24041 (N_24041,N_20696,N_22951);
or U24042 (N_24042,N_18468,N_19307);
xnor U24043 (N_24043,N_19521,N_23917);
nand U24044 (N_24044,N_20063,N_21803);
and U24045 (N_24045,N_18205,N_23724);
or U24046 (N_24046,N_23575,N_20377);
and U24047 (N_24047,N_22254,N_18391);
xor U24048 (N_24048,N_18017,N_18349);
and U24049 (N_24049,N_18751,N_21406);
or U24050 (N_24050,N_19606,N_23498);
nor U24051 (N_24051,N_20197,N_23045);
and U24052 (N_24052,N_20056,N_21389);
nor U24053 (N_24053,N_20324,N_19688);
nor U24054 (N_24054,N_18976,N_21077);
nor U24055 (N_24055,N_21285,N_19196);
nor U24056 (N_24056,N_19907,N_22844);
and U24057 (N_24057,N_19670,N_21594);
or U24058 (N_24058,N_21174,N_21528);
and U24059 (N_24059,N_22412,N_23531);
and U24060 (N_24060,N_18951,N_23074);
nand U24061 (N_24061,N_18116,N_21711);
xor U24062 (N_24062,N_19397,N_23119);
xnor U24063 (N_24063,N_23709,N_19737);
xor U24064 (N_24064,N_22233,N_20089);
nor U24065 (N_24065,N_21036,N_20505);
or U24066 (N_24066,N_22137,N_18258);
nor U24067 (N_24067,N_22642,N_19123);
nand U24068 (N_24068,N_19048,N_19214);
or U24069 (N_24069,N_19037,N_22732);
or U24070 (N_24070,N_19204,N_20202);
nor U24071 (N_24071,N_18268,N_20754);
xor U24072 (N_24072,N_21527,N_19050);
nor U24073 (N_24073,N_19456,N_20687);
nand U24074 (N_24074,N_19013,N_21859);
xnor U24075 (N_24075,N_18748,N_18277);
nor U24076 (N_24076,N_21502,N_21087);
nand U24077 (N_24077,N_18735,N_20163);
nand U24078 (N_24078,N_18266,N_20513);
and U24079 (N_24079,N_22878,N_19875);
nand U24080 (N_24080,N_20769,N_19353);
nor U24081 (N_24081,N_20786,N_18177);
nand U24082 (N_24082,N_18111,N_21520);
and U24083 (N_24083,N_18134,N_21691);
nor U24084 (N_24084,N_19629,N_22721);
nor U24085 (N_24085,N_20666,N_23920);
and U24086 (N_24086,N_22671,N_21190);
nor U24087 (N_24087,N_22831,N_18308);
or U24088 (N_24088,N_21352,N_20443);
or U24089 (N_24089,N_23554,N_18130);
or U24090 (N_24090,N_18305,N_20931);
or U24091 (N_24091,N_19291,N_22909);
xor U24092 (N_24092,N_20418,N_19853);
nor U24093 (N_24093,N_19847,N_21464);
nor U24094 (N_24094,N_23254,N_18097);
or U24095 (N_24095,N_23561,N_21833);
and U24096 (N_24096,N_18488,N_21119);
xor U24097 (N_24097,N_23640,N_23876);
nand U24098 (N_24098,N_19855,N_22304);
nor U24099 (N_24099,N_20721,N_23543);
and U24100 (N_24100,N_20693,N_19660);
and U24101 (N_24101,N_23886,N_19945);
xor U24102 (N_24102,N_19439,N_23056);
and U24103 (N_24103,N_20389,N_22761);
nand U24104 (N_24104,N_21591,N_18731);
nor U24105 (N_24105,N_21703,N_23742);
xnor U24106 (N_24106,N_22672,N_20662);
nor U24107 (N_24107,N_22320,N_20155);
nor U24108 (N_24108,N_18697,N_19802);
nor U24109 (N_24109,N_19457,N_18696);
or U24110 (N_24110,N_21214,N_18024);
nand U24111 (N_24111,N_23456,N_22783);
nor U24112 (N_24112,N_20676,N_19318);
nor U24113 (N_24113,N_20371,N_23809);
nand U24114 (N_24114,N_23943,N_22210);
nor U24115 (N_24115,N_18456,N_23659);
or U24116 (N_24116,N_19380,N_20745);
or U24117 (N_24117,N_23245,N_22859);
nand U24118 (N_24118,N_18596,N_18858);
or U24119 (N_24119,N_23545,N_23732);
xnor U24120 (N_24120,N_23955,N_23118);
nor U24121 (N_24121,N_21630,N_22084);
nor U24122 (N_24122,N_20374,N_23156);
or U24123 (N_24123,N_18331,N_19984);
xor U24124 (N_24124,N_23264,N_20205);
or U24125 (N_24125,N_19539,N_22925);
or U24126 (N_24126,N_23180,N_20869);
nand U24127 (N_24127,N_21079,N_18516);
nand U24128 (N_24128,N_19257,N_22299);
nor U24129 (N_24129,N_21521,N_18060);
nand U24130 (N_24130,N_22382,N_18941);
nand U24131 (N_24131,N_20706,N_19210);
xnor U24132 (N_24132,N_18050,N_18149);
nor U24133 (N_24133,N_22292,N_19655);
and U24134 (N_24134,N_20093,N_20494);
nand U24135 (N_24135,N_21861,N_19563);
or U24136 (N_24136,N_18685,N_20148);
nor U24137 (N_24137,N_18635,N_23193);
nor U24138 (N_24138,N_21633,N_23482);
nand U24139 (N_24139,N_19512,N_22873);
xor U24140 (N_24140,N_20958,N_18838);
xor U24141 (N_24141,N_21506,N_23146);
or U24142 (N_24142,N_22947,N_18671);
xor U24143 (N_24143,N_23785,N_18375);
or U24144 (N_24144,N_21608,N_19315);
or U24145 (N_24145,N_18025,N_18873);
xnor U24146 (N_24146,N_22248,N_22008);
xnor U24147 (N_24147,N_20780,N_22900);
nor U24148 (N_24148,N_20943,N_20841);
nor U24149 (N_24149,N_20495,N_23585);
nand U24150 (N_24150,N_20348,N_23263);
nor U24151 (N_24151,N_22729,N_20989);
nand U24152 (N_24152,N_19718,N_20556);
and U24153 (N_24153,N_22190,N_21136);
xor U24154 (N_24154,N_22867,N_23214);
and U24155 (N_24155,N_18726,N_23944);
xor U24156 (N_24156,N_21185,N_23484);
and U24157 (N_24157,N_20652,N_22754);
and U24158 (N_24158,N_22162,N_22046);
or U24159 (N_24159,N_20010,N_19709);
xor U24160 (N_24160,N_19236,N_23379);
nand U24161 (N_24161,N_18533,N_22067);
nor U24162 (N_24162,N_19114,N_19668);
xor U24163 (N_24163,N_22599,N_22032);
and U24164 (N_24164,N_23170,N_23136);
or U24165 (N_24165,N_18762,N_22948);
nor U24166 (N_24166,N_22243,N_20161);
xnor U24167 (N_24167,N_19129,N_20923);
or U24168 (N_24168,N_20315,N_21897);
nor U24169 (N_24169,N_22954,N_18743);
or U24170 (N_24170,N_21868,N_21088);
or U24171 (N_24171,N_19385,N_22056);
xor U24172 (N_24172,N_23516,N_23728);
xor U24173 (N_24173,N_21197,N_20435);
or U24174 (N_24174,N_21783,N_21923);
nand U24175 (N_24175,N_21975,N_18480);
or U24176 (N_24176,N_19951,N_22722);
xnor U24177 (N_24177,N_22763,N_18826);
or U24178 (N_24178,N_18422,N_18753);
xnor U24179 (N_24179,N_19506,N_23090);
xor U24180 (N_24180,N_22197,N_22713);
or U24181 (N_24181,N_22282,N_20028);
xor U24182 (N_24182,N_19806,N_21405);
or U24183 (N_24183,N_19648,N_19116);
nand U24184 (N_24184,N_21461,N_23567);
nor U24185 (N_24185,N_19029,N_18990);
or U24186 (N_24186,N_20400,N_21382);
xor U24187 (N_24187,N_19974,N_22790);
and U24188 (N_24188,N_23113,N_23149);
nor U24189 (N_24189,N_18080,N_23082);
or U24190 (N_24190,N_21613,N_18891);
nand U24191 (N_24191,N_18355,N_22189);
xor U24192 (N_24192,N_18105,N_23458);
nor U24193 (N_24193,N_22655,N_18723);
nand U24194 (N_24194,N_22780,N_18249);
xor U24195 (N_24195,N_18358,N_23541);
nand U24196 (N_24196,N_23235,N_18471);
nor U24197 (N_24197,N_20920,N_18368);
and U24198 (N_24198,N_18282,N_22420);
and U24199 (N_24199,N_22198,N_20818);
nand U24200 (N_24200,N_22235,N_23588);
xnor U24201 (N_24201,N_18169,N_20812);
nor U24202 (N_24202,N_20827,N_18011);
nor U24203 (N_24203,N_23514,N_20608);
nor U24204 (N_24204,N_20991,N_20549);
nand U24205 (N_24205,N_18522,N_19437);
nand U24206 (N_24206,N_19392,N_20762);
nand U24207 (N_24207,N_18323,N_22202);
and U24208 (N_24208,N_21243,N_20722);
and U24209 (N_24209,N_18770,N_21771);
nand U24210 (N_24210,N_22938,N_20641);
xnor U24211 (N_24211,N_22674,N_19821);
xor U24212 (N_24212,N_20902,N_21336);
nor U24213 (N_24213,N_21017,N_23021);
nor U24214 (N_24214,N_19698,N_22886);
nand U24215 (N_24215,N_23753,N_20862);
xor U24216 (N_24216,N_20551,N_22171);
nand U24217 (N_24217,N_18839,N_21732);
or U24218 (N_24218,N_22003,N_18700);
nand U24219 (N_24219,N_19369,N_22220);
xor U24220 (N_24220,N_19289,N_21616);
nand U24221 (N_24221,N_20100,N_19556);
nor U24222 (N_24222,N_19839,N_23756);
and U24223 (N_24223,N_21916,N_23397);
or U24224 (N_24224,N_22005,N_22510);
nand U24225 (N_24225,N_19733,N_18356);
xor U24226 (N_24226,N_18804,N_18380);
nor U24227 (N_24227,N_18805,N_20440);
nor U24228 (N_24228,N_18867,N_18360);
nor U24229 (N_24229,N_20948,N_23726);
nand U24230 (N_24230,N_20524,N_22592);
nand U24231 (N_24231,N_23915,N_21652);
nor U24232 (N_24232,N_22520,N_23346);
xor U24233 (N_24233,N_18737,N_19153);
nand U24234 (N_24234,N_21724,N_20635);
nand U24235 (N_24235,N_19156,N_23173);
or U24236 (N_24236,N_21702,N_21130);
nor U24237 (N_24237,N_23331,N_20013);
and U24238 (N_24238,N_21693,N_18216);
nand U24239 (N_24239,N_23020,N_23782);
nor U24240 (N_24240,N_21857,N_21663);
nor U24241 (N_24241,N_18992,N_18178);
or U24242 (N_24242,N_21941,N_22996);
nor U24243 (N_24243,N_22772,N_21626);
nand U24244 (N_24244,N_23054,N_23185);
or U24245 (N_24245,N_21765,N_19589);
nor U24246 (N_24246,N_20843,N_21120);
nand U24247 (N_24247,N_23820,N_23794);
and U24248 (N_24248,N_23924,N_22419);
xor U24249 (N_24249,N_19646,N_23835);
nor U24250 (N_24250,N_19502,N_20191);
xor U24251 (N_24251,N_19745,N_18874);
xnor U24252 (N_24252,N_18603,N_21681);
or U24253 (N_24253,N_18580,N_18864);
nand U24254 (N_24254,N_23127,N_22236);
xor U24255 (N_24255,N_22625,N_20103);
nand U24256 (N_24256,N_20265,N_22766);
and U24257 (N_24257,N_23392,N_21995);
and U24258 (N_24258,N_23240,N_20154);
and U24259 (N_24259,N_22854,N_18629);
xnor U24260 (N_24260,N_23981,N_20113);
xor U24261 (N_24261,N_23361,N_23810);
and U24262 (N_24262,N_22455,N_21426);
nand U24263 (N_24263,N_18009,N_19363);
or U24264 (N_24264,N_23050,N_18270);
nand U24265 (N_24265,N_21982,N_23819);
xnor U24266 (N_24266,N_21436,N_20636);
or U24267 (N_24267,N_18401,N_23026);
or U24268 (N_24268,N_18822,N_21296);
nand U24269 (N_24269,N_18657,N_18734);
nand U24270 (N_24270,N_20253,N_19599);
xor U24271 (N_24271,N_23988,N_19095);
xnor U24272 (N_24272,N_19561,N_19921);
and U24273 (N_24273,N_20376,N_20069);
or U24274 (N_24274,N_22490,N_21287);
or U24275 (N_24275,N_20590,N_23918);
or U24276 (N_24276,N_19404,N_19055);
nor U24277 (N_24277,N_21469,N_22629);
and U24278 (N_24278,N_21679,N_18912);
nand U24279 (N_24279,N_20227,N_22069);
and U24280 (N_24280,N_21231,N_18363);
xor U24281 (N_24281,N_20574,N_23631);
and U24282 (N_24282,N_23357,N_23879);
nor U24283 (N_24283,N_20293,N_23675);
nand U24284 (N_24284,N_18512,N_21943);
nor U24285 (N_24285,N_22566,N_18392);
and U24286 (N_24286,N_19374,N_18460);
nand U24287 (N_24287,N_18883,N_19631);
nor U24288 (N_24288,N_20898,N_21624);
and U24289 (N_24289,N_22196,N_20825);
xnor U24290 (N_24290,N_23394,N_21741);
nor U24291 (N_24291,N_18991,N_20528);
or U24292 (N_24292,N_20074,N_19477);
nor U24293 (N_24293,N_21516,N_18774);
and U24294 (N_24294,N_23586,N_18281);
nand U24295 (N_24295,N_20997,N_20472);
xor U24296 (N_24296,N_19836,N_23928);
nand U24297 (N_24297,N_18928,N_20157);
or U24298 (N_24298,N_23351,N_23603);
or U24299 (N_24299,N_20101,N_22088);
and U24300 (N_24300,N_20428,N_18683);
xnor U24301 (N_24301,N_19626,N_23171);
nand U24302 (N_24302,N_18232,N_22558);
or U24303 (N_24303,N_20115,N_22294);
nor U24304 (N_24304,N_19008,N_20726);
and U24305 (N_24305,N_23198,N_19225);
nand U24306 (N_24306,N_19043,N_22902);
xor U24307 (N_24307,N_19507,N_18535);
nor U24308 (N_24308,N_19499,N_23776);
xor U24309 (N_24309,N_23578,N_22562);
or U24310 (N_24310,N_23987,N_18336);
nor U24311 (N_24311,N_19068,N_21622);
nor U24312 (N_24312,N_19989,N_23716);
xnor U24313 (N_24313,N_22179,N_18299);
xnor U24314 (N_24314,N_19260,N_22051);
xor U24315 (N_24315,N_19928,N_23060);
nand U24316 (N_24316,N_23129,N_19316);
xnor U24317 (N_24317,N_18104,N_21704);
and U24318 (N_24318,N_21488,N_19194);
nor U24319 (N_24319,N_22230,N_21480);
or U24320 (N_24320,N_22329,N_20168);
nand U24321 (N_24321,N_22348,N_18901);
xor U24322 (N_24322,N_23938,N_23985);
or U24323 (N_24323,N_20125,N_23333);
nor U24324 (N_24324,N_18252,N_20033);
and U24325 (N_24325,N_22019,N_21498);
nand U24326 (N_24326,N_18601,N_22715);
nor U24327 (N_24327,N_22185,N_22495);
nand U24328 (N_24328,N_19440,N_21438);
and U24329 (N_24329,N_23192,N_18856);
and U24330 (N_24330,N_19940,N_22983);
xor U24331 (N_24331,N_23283,N_21987);
nor U24332 (N_24332,N_23232,N_22373);
nand U24333 (N_24333,N_22211,N_22680);
nor U24334 (N_24334,N_20462,N_22618);
xor U24335 (N_24335,N_23102,N_21717);
nor U24336 (N_24336,N_23693,N_20610);
and U24337 (N_24337,N_20170,N_20815);
or U24338 (N_24338,N_20309,N_19803);
or U24339 (N_24339,N_23803,N_23128);
nor U24340 (N_24340,N_20866,N_20468);
nand U24341 (N_24341,N_21390,N_21866);
xor U24342 (N_24342,N_21556,N_20102);
nor U24343 (N_24343,N_19579,N_18989);
nand U24344 (N_24344,N_22424,N_18439);
or U24345 (N_24345,N_21337,N_20996);
xnor U24346 (N_24346,N_18996,N_21294);
nand U24347 (N_24347,N_19387,N_18651);
nor U24348 (N_24348,N_23559,N_23654);
or U24349 (N_24349,N_19540,N_18892);
xnor U24350 (N_24350,N_19623,N_23404);
xor U24351 (N_24351,N_23857,N_19863);
nor U24352 (N_24352,N_22985,N_20381);
or U24353 (N_24353,N_21864,N_22911);
nor U24354 (N_24354,N_21614,N_19609);
nand U24355 (N_24355,N_20759,N_18402);
xnor U24356 (N_24356,N_18264,N_19366);
nor U24357 (N_24357,N_19014,N_21819);
nand U24358 (N_24358,N_20247,N_19750);
nand U24359 (N_24359,N_19751,N_22021);
and U24360 (N_24360,N_22040,N_22107);
or U24361 (N_24361,N_22444,N_23634);
nand U24362 (N_24362,N_21175,N_22508);
nor U24363 (N_24363,N_18257,N_22462);
or U24364 (N_24364,N_19526,N_21945);
nand U24365 (N_24365,N_20139,N_20334);
and U24366 (N_24366,N_22564,N_22781);
nor U24367 (N_24367,N_23501,N_21936);
xor U24368 (N_24368,N_21440,N_21199);
or U24369 (N_24369,N_19759,N_21661);
or U24370 (N_24370,N_21226,N_23900);
xnor U24371 (N_24371,N_22260,N_20336);
or U24372 (N_24372,N_19286,N_20385);
nand U24373 (N_24373,N_19616,N_19304);
and U24374 (N_24374,N_20517,N_20986);
or U24375 (N_24375,N_19358,N_19324);
or U24376 (N_24376,N_19040,N_23068);
or U24377 (N_24377,N_21582,N_21649);
xnor U24378 (N_24378,N_23160,N_20254);
or U24379 (N_24379,N_18703,N_18312);
and U24380 (N_24380,N_23353,N_21192);
or U24381 (N_24381,N_23885,N_18865);
and U24382 (N_24382,N_21940,N_22406);
or U24383 (N_24383,N_22020,N_23960);
nand U24384 (N_24384,N_22608,N_19902);
or U24385 (N_24385,N_23787,N_22333);
xnor U24386 (N_24386,N_18552,N_22026);
and U24387 (N_24387,N_23152,N_21770);
xnor U24388 (N_24388,N_18715,N_23461);
xor U24389 (N_24389,N_21718,N_22031);
and U24390 (N_24390,N_22851,N_19532);
or U24391 (N_24391,N_23682,N_23535);
nor U24392 (N_24392,N_18612,N_23937);
nor U24393 (N_24393,N_18511,N_18563);
nand U24394 (N_24394,N_19480,N_21415);
nand U24395 (N_24395,N_20893,N_18881);
or U24396 (N_24396,N_18483,N_21499);
and U24397 (N_24397,N_23676,N_18727);
nand U24398 (N_24398,N_20279,N_21368);
nand U24399 (N_24399,N_19443,N_18139);
nand U24400 (N_24400,N_23906,N_19880);
xnor U24401 (N_24401,N_22443,N_19336);
xor U24402 (N_24402,N_18524,N_18493);
xor U24403 (N_24403,N_19044,N_18879);
and U24404 (N_24404,N_22609,N_18566);
nor U24405 (N_24405,N_22789,N_22212);
xor U24406 (N_24406,N_23277,N_22002);
nor U24407 (N_24407,N_18972,N_22901);
xor U24408 (N_24408,N_22429,N_21339);
or U24409 (N_24409,N_22531,N_21056);
or U24410 (N_24410,N_20260,N_18747);
nand U24411 (N_24411,N_20886,N_20143);
nand U24412 (N_24412,N_20697,N_18558);
and U24413 (N_24413,N_22472,N_19973);
nand U24414 (N_24414,N_19819,N_18153);
nor U24415 (N_24415,N_23830,N_20582);
nand U24416 (N_24416,N_18414,N_21458);
xor U24417 (N_24417,N_23183,N_19628);
and U24418 (N_24418,N_23190,N_21090);
nor U24419 (N_24419,N_22459,N_22744);
nand U24420 (N_24420,N_21282,N_19882);
nor U24421 (N_24421,N_20741,N_23207);
nand U24422 (N_24422,N_18910,N_21909);
xor U24423 (N_24423,N_18370,N_20919);
and U24424 (N_24424,N_19031,N_20519);
or U24425 (N_24425,N_22264,N_23096);
and U24426 (N_24426,N_22506,N_18203);
or U24427 (N_24427,N_19103,N_19189);
xnor U24428 (N_24428,N_22926,N_21672);
nand U24429 (N_24429,N_21588,N_21767);
or U24430 (N_24430,N_22155,N_22118);
nor U24431 (N_24431,N_22327,N_23690);
nor U24432 (N_24432,N_20425,N_20643);
or U24433 (N_24433,N_22969,N_23393);
xor U24434 (N_24434,N_20166,N_22138);
and U24435 (N_24435,N_22071,N_23762);
nor U24436 (N_24436,N_21844,N_23580);
or U24437 (N_24437,N_20152,N_23812);
or U24438 (N_24438,N_22711,N_18669);
and U24439 (N_24439,N_21253,N_23839);
nand U24440 (N_24440,N_22317,N_19181);
xor U24441 (N_24441,N_21358,N_20094);
nor U24442 (N_24442,N_20077,N_19461);
and U24443 (N_24443,N_19442,N_23719);
xnor U24444 (N_24444,N_23976,N_23605);
and U24445 (N_24445,N_21429,N_21377);
and U24446 (N_24446,N_22613,N_21446);
or U24447 (N_24447,N_21885,N_22820);
nand U24448 (N_24448,N_23187,N_23560);
or U24449 (N_24449,N_21599,N_20508);
nand U24450 (N_24450,N_22688,N_23715);
or U24451 (N_24451,N_20908,N_20193);
nor U24452 (N_24452,N_19786,N_18262);
nor U24453 (N_24453,N_21057,N_18689);
nor U24454 (N_24454,N_21233,N_19932);
nand U24455 (N_24455,N_22270,N_20224);
nor U24456 (N_24456,N_23088,N_23743);
xor U24457 (N_24457,N_19725,N_20477);
nand U24458 (N_24458,N_19518,N_22582);
xnor U24459 (N_24459,N_20968,N_21105);
nand U24460 (N_24460,N_23382,N_21944);
or U24461 (N_24461,N_20399,N_22414);
and U24462 (N_24462,N_23657,N_18157);
nor U24463 (N_24463,N_23548,N_19898);
or U24464 (N_24464,N_22116,N_23505);
nand U24465 (N_24465,N_20024,N_19209);
and U24466 (N_24466,N_18560,N_18182);
nand U24467 (N_24467,N_18056,N_18749);
or U24468 (N_24468,N_18475,N_23048);
nor U24469 (N_24469,N_21579,N_21383);
nand U24470 (N_24470,N_23660,N_23574);
nand U24471 (N_24471,N_19983,N_22421);
nor U24472 (N_24472,N_23081,N_18223);
nor U24473 (N_24473,N_21500,N_23737);
nand U24474 (N_24474,N_19975,N_22023);
nand U24475 (N_24475,N_19262,N_21990);
nor U24476 (N_24476,N_18429,N_21523);
and U24477 (N_24477,N_23973,N_20867);
nor U24478 (N_24478,N_18317,N_19202);
nor U24479 (N_24479,N_21388,N_18746);
nor U24480 (N_24480,N_19362,N_22393);
or U24481 (N_24481,N_23705,N_18984);
nand U24482 (N_24482,N_19686,N_21935);
and U24483 (N_24483,N_18809,N_19294);
or U24484 (N_24484,N_22387,N_18244);
or U24485 (N_24485,N_21882,N_19666);
or U24486 (N_24486,N_21809,N_21788);
and U24487 (N_24487,N_23523,N_20577);
nand U24488 (N_24488,N_23789,N_21730);
nor U24489 (N_24489,N_19224,N_23865);
or U24490 (N_24490,N_23923,N_22918);
nand U24491 (N_24491,N_21238,N_19149);
xor U24492 (N_24492,N_20145,N_18474);
and U24493 (N_24493,N_21843,N_18947);
nor U24494 (N_24494,N_22979,N_22661);
nand U24495 (N_24495,N_21964,N_23869);
and U24496 (N_24496,N_20169,N_20219);
and U24497 (N_24497,N_18896,N_20097);
or U24498 (N_24498,N_18756,N_23925);
xnor U24499 (N_24499,N_20092,N_22471);
or U24500 (N_24500,N_21662,N_20391);
xor U24501 (N_24501,N_19379,N_21565);
or U24502 (N_24502,N_21725,N_19946);
and U24503 (N_24503,N_23701,N_22483);
nor U24504 (N_24504,N_23165,N_22364);
or U24505 (N_24505,N_23733,N_23860);
and U24506 (N_24506,N_19100,N_21140);
xor U24507 (N_24507,N_19144,N_19108);
nor U24508 (N_24508,N_18725,N_23914);
xnor U24509 (N_24509,N_19567,N_21554);
nor U24510 (N_24510,N_19060,N_19922);
nor U24511 (N_24511,N_21315,N_23518);
xor U24512 (N_24512,N_19419,N_20743);
nand U24513 (N_24513,N_21176,N_21660);
and U24514 (N_24514,N_18131,N_23215);
xnor U24515 (N_24515,N_21530,N_21570);
nand U24516 (N_24516,N_19382,N_22978);
xnor U24517 (N_24517,N_19656,N_19991);
and U24518 (N_24518,N_18226,N_20209);
xor U24519 (N_24519,N_20884,N_23166);
and U24520 (N_24520,N_20914,N_21733);
xnor U24521 (N_24521,N_18199,N_18457);
nor U24522 (N_24522,N_23189,N_22353);
nor U24523 (N_24523,N_19180,N_23005);
and U24524 (N_24524,N_22651,N_20804);
or U24525 (N_24525,N_21618,N_21609);
xnor U24526 (N_24526,N_20455,N_21902);
xor U24527 (N_24527,N_21158,N_21305);
nor U24528 (N_24528,N_21013,N_18803);
and U24529 (N_24529,N_22309,N_20109);
xor U24530 (N_24530,N_22541,N_22803);
or U24531 (N_24531,N_21610,N_22982);
xor U24532 (N_24532,N_23587,N_22142);
xor U24533 (N_24533,N_23700,N_19730);
nor U24534 (N_24534,N_20823,N_20890);
and U24535 (N_24535,N_22059,N_18962);
and U24536 (N_24536,N_20498,N_21380);
nand U24537 (N_24537,N_21888,N_20790);
xnor U24538 (N_24538,N_23802,N_21895);
or U24539 (N_24539,N_22677,N_22000);
and U24540 (N_24540,N_22514,N_19494);
xor U24541 (N_24541,N_19511,N_23913);
or U24542 (N_24542,N_20795,N_18890);
xnor U24543 (N_24543,N_23788,N_20714);
nor U24544 (N_24544,N_22193,N_23901);
and U24545 (N_24545,N_21103,N_21291);
xor U24546 (N_24546,N_18549,N_21467);
xor U24547 (N_24547,N_23816,N_20207);
xnor U24548 (N_24548,N_20980,N_21557);
nor U24549 (N_24549,N_18241,N_20189);
or U24550 (N_24550,N_23669,N_21481);
and U24551 (N_24551,N_22690,N_22731);
nor U24552 (N_24552,N_18255,N_22434);
nor U24553 (N_24553,N_20308,N_18383);
and U24554 (N_24554,N_23451,N_19098);
or U24555 (N_24555,N_20648,N_18759);
xor U24556 (N_24556,N_22795,N_18985);
or U24557 (N_24557,N_21970,N_20945);
nand U24558 (N_24558,N_22047,N_18889);
nand U24559 (N_24559,N_19585,N_21801);
nor U24560 (N_24560,N_20190,N_22517);
and U24561 (N_24561,N_21992,N_21543);
nand U24562 (N_24562,N_23064,N_21327);
nand U24563 (N_24563,N_21782,N_20546);
and U24564 (N_24564,N_19702,N_20793);
nor U24565 (N_24565,N_22039,N_21988);
nand U24566 (N_24566,N_18274,N_18110);
xor U24567 (N_24567,N_22726,N_22042);
and U24568 (N_24568,N_19357,N_23932);
or U24569 (N_24569,N_20460,N_21719);
nand U24570 (N_24570,N_23499,N_19647);
nor U24571 (N_24571,N_18037,N_21714);
or U24572 (N_24572,N_20680,N_21839);
or U24573 (N_24573,N_18786,N_18510);
xor U24574 (N_24574,N_23954,N_20222);
or U24575 (N_24575,N_22866,N_18300);
or U24576 (N_24576,N_21981,N_21189);
nand U24577 (N_24577,N_19465,N_21700);
xnor U24578 (N_24578,N_23570,N_23852);
or U24579 (N_24579,N_19453,N_20164);
and U24580 (N_24580,N_19490,N_18303);
and U24581 (N_24581,N_18797,N_22644);
xor U24582 (N_24582,N_22773,N_22013);
and U24583 (N_24583,N_19232,N_19901);
and U24584 (N_24584,N_21925,N_23179);
xor U24585 (N_24585,N_21360,N_20707);
nor U24586 (N_24586,N_20122,N_19947);
nor U24587 (N_24587,N_23592,N_21802);
nor U24588 (N_24588,N_23234,N_23624);
or U24589 (N_24589,N_19271,N_23695);
or U24590 (N_24590,N_21448,N_20985);
xnor U24591 (N_24591,N_20799,N_19411);
and U24592 (N_24592,N_21129,N_20963);
nand U24593 (N_24593,N_18810,N_21369);
and U24594 (N_24594,N_20817,N_23194);
nor U24595 (N_24595,N_22734,N_23793);
nor U24596 (N_24596,N_20403,N_22559);
and U24597 (N_24597,N_18246,N_20547);
nand U24598 (N_24598,N_23062,N_22561);
and U24599 (N_24599,N_18772,N_20330);
xor U24600 (N_24600,N_20310,N_21670);
nand U24601 (N_24601,N_18885,N_22590);
or U24602 (N_24602,N_18942,N_22375);
or U24603 (N_24603,N_21128,N_20014);
or U24604 (N_24604,N_19912,N_20323);
xor U24605 (N_24605,N_21146,N_22109);
and U24606 (N_24606,N_23509,N_18278);
and U24607 (N_24607,N_23431,N_21216);
nor U24608 (N_24608,N_18019,N_22952);
nand U24609 (N_24609,N_18194,N_20312);
and U24610 (N_24610,N_22676,N_23783);
xor U24611 (N_24611,N_20162,N_19734);
nand U24612 (N_24612,N_23757,N_20881);
or U24613 (N_24613,N_18489,N_22226);
and U24614 (N_24614,N_23153,N_20185);
xnor U24615 (N_24615,N_22234,N_19762);
nor U24616 (N_24616,N_21739,N_21785);
and U24617 (N_24617,N_19939,N_23284);
or U24618 (N_24618,N_19154,N_20467);
or U24619 (N_24619,N_22287,N_22526);
or U24620 (N_24620,N_18417,N_19782);
nand U24621 (N_24621,N_23542,N_23683);
and U24622 (N_24622,N_22043,N_20611);
or U24623 (N_24623,N_23590,N_21764);
or U24624 (N_24624,N_18782,N_20430);
and U24625 (N_24625,N_20704,N_22749);
nor U24626 (N_24626,N_23476,N_23650);
nand U24627 (N_24627,N_22576,N_19517);
or U24628 (N_24628,N_21221,N_23133);
nor U24629 (N_24629,N_20669,N_22385);
or U24630 (N_24630,N_20561,N_18348);
nor U24631 (N_24631,N_22546,N_18775);
or U24632 (N_24632,N_22437,N_20760);
xnor U24633 (N_24633,N_21856,N_18316);
nor U24634 (N_24634,N_20142,N_22916);
nand U24635 (N_24635,N_20675,N_20564);
nor U24636 (N_24636,N_20961,N_23201);
nand U24637 (N_24637,N_19534,N_23416);
and U24638 (N_24638,N_23995,N_21867);
nand U24639 (N_24639,N_22652,N_18636);
and U24640 (N_24640,N_21269,N_18291);
or U24641 (N_24641,N_22693,N_20683);
or U24642 (N_24642,N_22409,N_18583);
and U24643 (N_24643,N_20034,N_21536);
xor U24644 (N_24644,N_21954,N_21628);
xor U24645 (N_24645,N_20402,N_22764);
nand U24646 (N_24646,N_19824,N_20619);
and U24647 (N_24647,N_19651,N_21366);
nand U24648 (N_24648,N_22791,N_20011);
nor U24649 (N_24649,N_20274,N_19551);
xnor U24650 (N_24650,N_22993,N_23714);
nand U24651 (N_24651,N_23046,N_20550);
nand U24652 (N_24652,N_23880,N_21705);
xor U24653 (N_24653,N_19719,N_22686);
nand U24654 (N_24654,N_19780,N_23041);
nand U24655 (N_24655,N_20245,N_22206);
or U24656 (N_24656,N_20553,N_23366);
xnor U24657 (N_24657,N_20257,N_19910);
and U24658 (N_24658,N_23405,N_18869);
or U24659 (N_24659,N_18042,N_19238);
xor U24660 (N_24660,N_20108,N_18953);
xor U24661 (N_24661,N_22577,N_18144);
nor U24662 (N_24662,N_20369,N_22182);
and U24663 (N_24663,N_20781,N_18712);
and U24664 (N_24664,N_19297,N_22014);
or U24665 (N_24665,N_18376,N_21999);
xor U24666 (N_24666,N_19147,N_22906);
xor U24667 (N_24667,N_22426,N_19279);
or U24668 (N_24668,N_19092,N_21592);
or U24669 (N_24669,N_19956,N_18201);
or U24670 (N_24670,N_20794,N_22295);
nand U24671 (N_24671,N_23725,N_19229);
nor U24672 (N_24672,N_18394,N_20447);
nor U24673 (N_24673,N_19992,N_20331);
and U24674 (N_24674,N_20290,N_22267);
or U24675 (N_24675,N_23139,N_22673);
and U24676 (N_24676,N_23015,N_18967);
or U24677 (N_24677,N_20918,N_20066);
xor U24678 (N_24678,N_20858,N_20378);
nor U24679 (N_24679,N_20756,N_22836);
or U24680 (N_24680,N_23184,N_18476);
or U24681 (N_24681,N_19252,N_20390);
or U24682 (N_24682,N_23467,N_21680);
and U24683 (N_24683,N_19481,N_21977);
xnor U24684 (N_24684,N_22275,N_21386);
and U24685 (N_24685,N_23933,N_23990);
or U24686 (N_24686,N_21025,N_23890);
or U24687 (N_24687,N_19350,N_23178);
or U24688 (N_24688,N_23304,N_22743);
and U24689 (N_24689,N_22286,N_21097);
xnor U24690 (N_24690,N_19966,N_22268);
and U24691 (N_24691,N_18564,N_18592);
xor U24692 (N_24692,N_19683,N_18799);
and U24693 (N_24693,N_20850,N_20957);
xor U24694 (N_24694,N_21361,N_22025);
xnor U24695 (N_24695,N_20929,N_19074);
xor U24696 (N_24696,N_21540,N_22811);
xnor U24697 (N_24697,N_22572,N_20039);
or U24698 (N_24698,N_20239,N_19545);
nor U24699 (N_24699,N_20629,N_19876);
nand U24700 (N_24700,N_20969,N_19038);
nor U24701 (N_24701,N_18306,N_22346);
xor U24702 (N_24702,N_20196,N_22915);
or U24703 (N_24703,N_19790,N_21181);
nor U24704 (N_24704,N_23306,N_18432);
or U24705 (N_24705,N_19096,N_20276);
nor U24706 (N_24706,N_18974,N_18238);
xor U24707 (N_24707,N_21298,N_22464);
and U24708 (N_24708,N_22435,N_18343);
and U24709 (N_24709,N_19842,N_22501);
nor U24710 (N_24710,N_20184,N_21201);
nor U24711 (N_24711,N_23555,N_19157);
and U24712 (N_24712,N_19554,N_19326);
nand U24713 (N_24713,N_18664,N_22209);
nor U24714 (N_24714,N_18227,N_20394);
nand U24715 (N_24715,N_23012,N_19838);
xor U24716 (N_24716,N_19188,N_23813);
or U24717 (N_24717,N_23330,N_23579);
xnor U24718 (N_24718,N_20792,N_21252);
or U24719 (N_24719,N_20382,N_23770);
and U24720 (N_24720,N_21643,N_20798);
or U24721 (N_24721,N_22802,N_20225);
nor U24722 (N_24722,N_19987,N_23063);
and U24723 (N_24723,N_22068,N_21423);
xor U24724 (N_24724,N_23630,N_20978);
and U24725 (N_24725,N_22966,N_23758);
nor U24726 (N_24726,N_20746,N_18212);
or U24727 (N_24727,N_19845,N_20548);
xor U24728 (N_24728,N_23889,N_23596);
or U24729 (N_24729,N_18224,N_21601);
or U24730 (N_24730,N_23249,N_21441);
and U24731 (N_24731,N_23462,N_23104);
and U24732 (N_24732,N_22864,N_23343);
nor U24733 (N_24733,N_18181,N_22816);
nor U24734 (N_24734,N_21734,N_19265);
xor U24735 (N_24735,N_18800,N_23007);
xor U24736 (N_24736,N_21775,N_19749);
nand U24737 (N_24737,N_23754,N_23365);
nor U24738 (N_24738,N_18913,N_21302);
nor U24739 (N_24739,N_19109,N_20305);
nor U24740 (N_24740,N_23708,N_20606);
nand U24741 (N_24741,N_18646,N_21114);
nand U24742 (N_24742,N_21309,N_19586);
xnor U24743 (N_24743,N_19724,N_20514);
and U24744 (N_24744,N_22436,N_20776);
and U24745 (N_24745,N_19931,N_18487);
nor U24746 (N_24746,N_21378,N_22753);
xor U24747 (N_24747,N_20578,N_23058);
xnor U24748 (N_24748,N_20195,N_20764);
nand U24749 (N_24749,N_20484,N_21677);
and U24750 (N_24750,N_23172,N_23196);
nor U24751 (N_24751,N_22641,N_19615);
nand U24752 (N_24752,N_18140,N_20822);
nor U24753 (N_24753,N_23391,N_19378);
and U24754 (N_24754,N_19583,N_23864);
nand U24755 (N_24755,N_23667,N_20739);
and U24756 (N_24756,N_18490,N_18849);
nand U24757 (N_24757,N_19372,N_19543);
nand U24758 (N_24758,N_18209,N_18707);
xor U24759 (N_24759,N_22861,N_23573);
nand U24760 (N_24760,N_23419,N_21153);
nor U24761 (N_24761,N_20729,N_23326);
and U24762 (N_24762,N_19302,N_23912);
nor U24763 (N_24763,N_18903,N_21259);
or U24764 (N_24764,N_20420,N_19565);
nand U24765 (N_24765,N_18637,N_21356);
and U24766 (N_24766,N_22667,N_19247);
or U24767 (N_24767,N_21706,N_19953);
nor U24768 (N_24768,N_22771,N_21150);
xnor U24769 (N_24769,N_20834,N_18354);
nand U24770 (N_24770,N_23735,N_20870);
nor U24771 (N_24771,N_21141,N_20583);
or U24772 (N_24772,N_22144,N_21972);
and U24773 (N_24773,N_21632,N_20596);
and U24774 (N_24774,N_22133,N_23790);
or U24775 (N_24775,N_22843,N_18057);
nand U24776 (N_24776,N_23140,N_21698);
xnor U24777 (N_24777,N_22480,N_18773);
or U24778 (N_24778,N_20004,N_22416);
xor U24779 (N_24779,N_22229,N_20045);
or U24780 (N_24780,N_22890,N_23740);
nor U24781 (N_24781,N_18733,N_19944);
xor U24782 (N_24782,N_19199,N_21837);
or U24783 (N_24783,N_19635,N_22452);
nor U24784 (N_24784,N_19010,N_22044);
and U24785 (N_24785,N_21590,N_23532);
nor U24786 (N_24786,N_23292,N_22018);
and U24787 (N_24787,N_19240,N_22087);
and U24788 (N_24788,N_21071,N_21538);
and U24789 (N_24789,N_21673,N_21629);
and U24790 (N_24790,N_18143,N_23571);
and U24791 (N_24791,N_19971,N_21627);
and U24792 (N_24792,N_19455,N_20612);
nor U24793 (N_24793,N_20288,N_20452);
nand U24794 (N_24794,N_18228,N_21533);
or U24795 (N_24795,N_22876,N_21603);
nor U24796 (N_24796,N_22953,N_23847);
and U24797 (N_24797,N_19761,N_22892);
nor U24798 (N_24798,N_23850,N_18290);
nor U24799 (N_24799,N_22687,N_21452);
nor U24800 (N_24800,N_23327,N_18961);
xnor U24801 (N_24801,N_19659,N_18843);
and U24802 (N_24802,N_22316,N_23703);
or U24803 (N_24803,N_23206,N_19256);
and U24804 (N_24804,N_22737,N_21445);
nor U24805 (N_24805,N_21014,N_22156);
and U24806 (N_24806,N_22929,N_20008);
xnor U24807 (N_24807,N_20047,N_19650);
and U24808 (N_24808,N_21664,N_21760);
and U24809 (N_24809,N_19796,N_20392);
and U24810 (N_24810,N_20953,N_19663);
xnor U24811 (N_24811,N_22650,N_22240);
or U24812 (N_24812,N_23006,N_23897);
or U24813 (N_24813,N_20249,N_19717);
xnor U24814 (N_24814,N_19636,N_19864);
xnor U24815 (N_24815,N_18859,N_20509);
nand U24816 (N_24816,N_19432,N_20552);
nand U24817 (N_24817,N_21234,N_19425);
xnor U24818 (N_24818,N_18789,N_20339);
nor U24819 (N_24819,N_22485,N_22848);
and U24820 (N_24820,N_19744,N_21820);
or U24821 (N_24821,N_19337,N_18211);
nor U24822 (N_24822,N_19760,N_23468);
and U24823 (N_24823,N_19361,N_19584);
or U24824 (N_24824,N_19772,N_19830);
xor U24825 (N_24825,N_21183,N_20593);
nor U24826 (N_24826,N_20007,N_20232);
and U24827 (N_24827,N_22511,N_22922);
and U24828 (N_24828,N_21612,N_22654);
nand U24829 (N_24829,N_20458,N_18607);
nand U24830 (N_24830,N_20214,N_22507);
xnor U24831 (N_24831,N_23301,N_22895);
and U24832 (N_24832,N_22817,N_20545);
or U24833 (N_24833,N_21780,N_18128);
and U24834 (N_24834,N_19815,N_21102);
and U24835 (N_24835,N_19482,N_23681);
xor U24836 (N_24836,N_20820,N_19080);
nor U24837 (N_24837,N_22147,N_18876);
or U24838 (N_24838,N_22569,N_19416);
xor U24839 (N_24839,N_20678,N_21756);
nor U24840 (N_24840,N_20431,N_23831);
nand U24841 (N_24841,N_21484,N_20365);
xor U24842 (N_24842,N_22921,N_20126);
xor U24843 (N_24843,N_18018,N_22163);
nor U24844 (N_24844,N_18918,N_21451);
nor U24845 (N_24845,N_20557,N_23470);
or U24846 (N_24846,N_18367,N_23524);
and U24847 (N_24847,N_18074,N_21407);
or U24848 (N_24848,N_21121,N_20592);
or U24849 (N_24849,N_22967,N_20272);
or U24850 (N_24850,N_22124,N_21408);
nor U24851 (N_24851,N_19633,N_18068);
or U24852 (N_24852,N_22215,N_23004);
and U24853 (N_24853,N_23145,N_21125);
nor U24854 (N_24854,N_18204,N_21475);
nor U24855 (N_24855,N_19476,N_23300);
or U24856 (N_24856,N_19776,N_22343);
or U24857 (N_24857,N_21418,N_23257);
or U24858 (N_24858,N_23086,N_21666);
xnor U24859 (N_24859,N_18172,N_22955);
nor U24860 (N_24860,N_18240,N_19529);
or U24861 (N_24861,N_18574,N_18245);
nor U24862 (N_24862,N_18504,N_19905);
and U24863 (N_24863,N_21574,N_19275);
xor U24864 (N_24864,N_19678,N_22446);
xor U24865 (N_24865,N_22549,N_21073);
xnor U24866 (N_24866,N_20298,N_19729);
or U24867 (N_24867,N_22319,N_23115);
nand U24868 (N_24868,N_18925,N_21490);
or U24869 (N_24869,N_23256,N_21171);
and U24870 (N_24870,N_19429,N_20591);
or U24871 (N_24871,N_18778,N_22679);
and U24872 (N_24872,N_20448,N_20188);
nor U24873 (N_24873,N_21062,N_20638);
nand U24874 (N_24874,N_18661,N_23280);
or U24875 (N_24875,N_18467,N_18729);
nand U24876 (N_24876,N_20690,N_23414);
nor U24877 (N_24877,N_19450,N_21258);
nor U24878 (N_24878,N_23842,N_20748);
nor U24879 (N_24879,N_19320,N_18094);
nand U24880 (N_24880,N_22388,N_18548);
or U24881 (N_24881,N_20563,N_18922);
nor U24882 (N_24882,N_18003,N_20114);
xnor U24883 (N_24883,N_23956,N_18935);
nor U24884 (N_24884,N_19267,N_20150);
nor U24885 (N_24885,N_23838,N_20727);
nand U24886 (N_24886,N_23084,N_18096);
and U24887 (N_24887,N_18162,N_22055);
or U24888 (N_24888,N_21311,N_23823);
and U24889 (N_24889,N_23114,N_18052);
nand U24890 (N_24890,N_23436,N_21228);
or U24891 (N_24891,N_18176,N_19205);
nand U24892 (N_24892,N_19997,N_21561);
nor U24893 (N_24893,N_22888,N_18448);
or U24894 (N_24894,N_19243,N_22405);
and U24895 (N_24895,N_18667,N_20282);
nand U24896 (N_24896,N_22784,N_21286);
nand U24897 (N_24897,N_21491,N_18923);
xor U24898 (N_24898,N_22274,N_19850);
xor U24899 (N_24899,N_21310,N_23796);
and U24900 (N_24900,N_20380,N_21263);
nor U24901 (N_24901,N_20566,N_18528);
nand U24902 (N_24902,N_20464,N_20277);
xor U24903 (N_24903,N_18846,N_23372);
nand U24904 (N_24904,N_20473,N_23248);
nand U24905 (N_24905,N_23875,N_19553);
nor U24906 (N_24906,N_23291,N_18173);
nand U24907 (N_24907,N_21346,N_21419);
nor U24908 (N_24908,N_22552,N_23622);
or U24909 (N_24909,N_19661,N_21720);
and U24910 (N_24910,N_18112,N_19924);
nor U24911 (N_24911,N_23325,N_18640);
xor U24912 (N_24912,N_23453,N_22942);
nor U24913 (N_24913,N_23583,N_19693);
nand U24914 (N_24914,N_22034,N_21694);
and U24915 (N_24915,N_21918,N_21914);
and U24916 (N_24916,N_22941,N_21133);
nand U24917 (N_24917,N_18195,N_18156);
nand U24918 (N_24918,N_22752,N_22887);
nand U24919 (N_24919,N_22774,N_22639);
nor U24920 (N_24920,N_22504,N_18345);
and U24921 (N_24921,N_22322,N_21752);
xnor U24922 (N_24922,N_23625,N_20763);
or U24923 (N_24923,N_23919,N_23929);
xor U24924 (N_24924,N_21932,N_20941);
nand U24925 (N_24925,N_21316,N_20842);
and U24926 (N_24926,N_21170,N_22823);
nor U24927 (N_24927,N_21598,N_18286);
xnor U24928 (N_24928,N_19186,N_23446);
nand U24929 (N_24929,N_18981,N_23014);
nand U24930 (N_24930,N_22366,N_22580);
and U24931 (N_24931,N_21876,N_19808);
and U24932 (N_24932,N_23017,N_20751);
nand U24933 (N_24933,N_21262,N_22134);
or U24934 (N_24934,N_22932,N_20237);
and U24935 (N_24935,N_19854,N_18243);
nand U24936 (N_24936,N_20328,N_23226);
xnor U24937 (N_24937,N_23829,N_18900);
or U24938 (N_24938,N_22298,N_20303);
xor U24939 (N_24939,N_22863,N_23795);
nand U24940 (N_24940,N_20609,N_22398);
xnor U24941 (N_24941,N_20783,N_20252);
xnor U24942 (N_24942,N_20705,N_19137);
nor U24943 (N_24943,N_23904,N_22312);
nand U24944 (N_24944,N_22169,N_20589);
xnor U24945 (N_24945,N_20501,N_21048);
and U24946 (N_24946,N_21235,N_18693);
and U24947 (N_24947,N_23859,N_19305);
nand U24948 (N_24948,N_21357,N_20295);
xor U24949 (N_24949,N_21825,N_19743);
nand U24950 (N_24950,N_19012,N_22386);
nand U24951 (N_24951,N_23407,N_20785);
nand U24952 (N_24952,N_19388,N_19671);
nand U24953 (N_24953,N_18400,N_21886);
or U24954 (N_24954,N_22477,N_22702);
nand U24955 (N_24955,N_23091,N_21300);
and U24956 (N_24956,N_19283,N_21272);
nor U24957 (N_24957,N_23177,N_22244);
nor U24958 (N_24958,N_21278,N_20499);
or U24959 (N_24959,N_21938,N_20141);
nor U24960 (N_24960,N_18835,N_21620);
nand U24961 (N_24961,N_20280,N_19692);
xor U24962 (N_24962,N_18135,N_19654);
nor U24963 (N_24963,N_18430,N_20856);
nor U24964 (N_24964,N_19331,N_22422);
nand U24965 (N_24965,N_21035,N_20967);
nand U24966 (N_24966,N_21038,N_19998);
and U24967 (N_24967,N_20084,N_23386);
xnor U24968 (N_24968,N_20082,N_19783);
and U24969 (N_24969,N_18395,N_22540);
xor U24970 (N_24970,N_23098,N_19258);
and U24971 (N_24971,N_18462,N_18327);
and U24972 (N_24972,N_20438,N_21248);
and U24973 (N_24973,N_21122,N_20261);
or U24974 (N_24974,N_19877,N_18730);
and U24975 (N_24975,N_23600,N_23100);
xnor U24976 (N_24976,N_19359,N_23341);
and U24977 (N_24977,N_22733,N_18248);
xor U24978 (N_24978,N_19197,N_20401);
and U24979 (N_24979,N_18870,N_18676);
nand U24980 (N_24980,N_20570,N_20851);
and U24981 (N_24981,N_23422,N_19559);
nor U24982 (N_24982,N_19192,N_23345);
nor U24983 (N_24983,N_20536,N_20079);
and U24984 (N_24984,N_22696,N_21064);
or U24985 (N_24985,N_18148,N_18256);
or U24986 (N_24986,N_18289,N_18897);
nor U24987 (N_24987,N_22293,N_22806);
and U24988 (N_24988,N_20568,N_21755);
nor U24989 (N_24989,N_22692,N_19332);
xor U24990 (N_24990,N_22814,N_18217);
nor U24991 (N_24991,N_19611,N_19282);
nor U24992 (N_24992,N_21878,N_23390);
xnor U24993 (N_24993,N_20058,N_23251);
nand U24994 (N_24994,N_18325,N_20955);
and U24995 (N_24995,N_22659,N_23526);
nand U24996 (N_24996,N_19470,N_23899);
nand U24997 (N_24997,N_22201,N_20623);
or U24998 (N_24998,N_21118,N_21251);
and U24999 (N_24999,N_19067,N_18828);
and U25000 (N_25000,N_20387,N_20810);
or U25001 (N_25001,N_23072,N_20417);
and U25002 (N_25002,N_22093,N_23908);
xnor U25003 (N_25003,N_18572,N_18551);
xnor U25004 (N_25004,N_20833,N_18526);
xnor U25005 (N_25005,N_20144,N_22368);
nand U25006 (N_25006,N_22272,N_21351);
or U25007 (N_25007,N_18590,N_23360);
and U25008 (N_25008,N_20976,N_21708);
and U25009 (N_25009,N_19617,N_20345);
or U25010 (N_25010,N_19794,N_21161);
and U25011 (N_25011,N_18641,N_18817);
and U25012 (N_25012,N_18218,N_22203);
nor U25013 (N_25013,N_19222,N_21365);
nor U25014 (N_25014,N_22458,N_20216);
or U25015 (N_25015,N_19217,N_18072);
nor U25016 (N_25016,N_21081,N_19193);
or U25017 (N_25017,N_19393,N_21794);
and U25018 (N_25018,N_21962,N_18340);
nor U25019 (N_25019,N_22256,N_23144);
xor U25020 (N_25020,N_19233,N_21395);
xor U25021 (N_25021,N_18819,N_19007);
and U25022 (N_25022,N_20429,N_21580);
nor U25023 (N_25023,N_22581,N_19523);
nor U25024 (N_25024,N_23413,N_21726);
nand U25025 (N_25025,N_18496,N_23730);
nor U25026 (N_25026,N_23504,N_21841);
nand U25027 (N_25027,N_22102,N_18263);
and U25028 (N_25028,N_22986,N_22062);
and U25029 (N_25029,N_23018,N_23942);
and U25030 (N_25030,N_20865,N_19295);
nand U25031 (N_25031,N_20479,N_23975);
nor U25032 (N_25032,N_21342,N_20750);
nand U25033 (N_25033,N_18197,N_20829);
or U25034 (N_25034,N_23710,N_19680);
nor U25035 (N_25035,N_19814,N_18154);
nor U25036 (N_25036,N_20119,N_22296);
or U25037 (N_25037,N_19662,N_18613);
nor U25038 (N_25038,N_18279,N_22064);
or U25039 (N_25039,N_23849,N_22136);
or U25040 (N_25040,N_22542,N_20981);
nor U25041 (N_25041,N_20504,N_19400);
xor U25042 (N_25042,N_22548,N_20306);
nand U25043 (N_25043,N_18214,N_20281);
and U25044 (N_25044,N_23980,N_23959);
xnor U25045 (N_25045,N_20104,N_21638);
nor U25046 (N_25046,N_21522,N_22606);
nand U25047 (N_25047,N_19753,N_23692);
xor U25048 (N_25048,N_19102,N_23738);
nor U25049 (N_25049,N_18577,N_19462);
nor U25050 (N_25050,N_19447,N_19327);
nor U25051 (N_25051,N_20083,N_21526);
xor U25052 (N_25052,N_21364,N_22894);
xnor U25053 (N_25053,N_21871,N_22998);
nor U25054 (N_25054,N_23679,N_19917);
and U25055 (N_25055,N_21463,N_21193);
and U25056 (N_25056,N_22984,N_23022);
nor U25057 (N_25057,N_21754,N_22395);
or U25058 (N_25058,N_23261,N_19219);
nand U25059 (N_25059,N_22208,N_21318);
and U25060 (N_25060,N_21224,N_21308);
and U25061 (N_25061,N_19161,N_19832);
or U25062 (N_25062,N_22880,N_22290);
nor U25063 (N_25063,N_19968,N_18499);
or U25064 (N_25064,N_23949,N_23157);
or U25065 (N_25065,N_19001,N_21814);
or U25066 (N_25066,N_19644,N_20791);
or U25067 (N_25067,N_23244,N_21343);
nor U25068 (N_25068,N_19119,N_23241);
or U25069 (N_25069,N_19952,N_22977);
and U25070 (N_25070,N_19538,N_19564);
and U25071 (N_25071,N_21134,N_22280);
nor U25072 (N_25072,N_23781,N_23668);
nand U25073 (N_25073,N_19531,N_19996);
and U25074 (N_25074,N_18624,N_23702);
and U25075 (N_25075,N_19915,N_18066);
and U25076 (N_25076,N_20134,N_19960);
or U25077 (N_25077,N_19127,N_22796);
or U25078 (N_25078,N_23321,N_22937);
and U25079 (N_25079,N_22360,N_21835);
nand U25080 (N_25080,N_20465,N_21401);
xnor U25081 (N_25081,N_20631,N_22804);
nand U25082 (N_25082,N_21776,N_19328);
or U25083 (N_25083,N_22075,N_18320);
nor U25084 (N_25084,N_22038,N_21653);
and U25085 (N_25085,N_23337,N_18397);
and U25086 (N_25086,N_21092,N_20407);
and U25087 (N_25087,N_23111,N_20735);
or U25088 (N_25088,N_21571,N_21659);
or U25089 (N_25089,N_21743,N_22228);
and U25090 (N_25090,N_23786,N_19272);
nor U25091 (N_25091,N_19568,N_18745);
and U25092 (N_25092,N_22371,N_23840);
and U25093 (N_25093,N_23992,N_21967);
nor U25094 (N_25094,N_22470,N_20029);
nor U25095 (N_25095,N_21564,N_23473);
xor U25096 (N_25096,N_23285,N_19859);
and U25097 (N_25097,N_22266,N_22076);
or U25098 (N_25098,N_22259,N_19602);
or U25099 (N_25099,N_19207,N_22720);
xnor U25100 (N_25100,N_21723,N_18924);
xnor U25101 (N_25101,N_20990,N_20208);
and U25102 (N_25102,N_21761,N_20944);
and U25103 (N_25103,N_18332,N_22798);
or U25104 (N_25104,N_20311,N_21830);
nand U25105 (N_25105,N_23367,N_23520);
xnor U25106 (N_25106,N_21093,N_21486);
and U25107 (N_25107,N_21430,N_22015);
nor U25108 (N_25108,N_22809,N_19211);
or U25109 (N_25109,N_18532,N_22289);
nand U25110 (N_25110,N_23642,N_19590);
xor U25111 (N_25111,N_18167,N_18611);
and U25112 (N_25112,N_22184,N_20432);
nor U25113 (N_25113,N_20246,N_22621);
or U25114 (N_25114,N_19488,N_23601);
or U25115 (N_25115,N_23447,N_21169);
nor U25116 (N_25116,N_19087,N_23720);
xor U25117 (N_25117,N_22199,N_20607);
nand U25118 (N_25118,N_22376,N_20284);
or U25119 (N_25119,N_23176,N_23148);
or U25120 (N_25120,N_22740,N_22633);
nor U25121 (N_25121,N_22626,N_19542);
or U25122 (N_25122,N_20040,N_18073);
or U25123 (N_25123,N_19231,N_19312);
nor U25124 (N_25124,N_20772,N_20386);
nand U25125 (N_25125,N_22466,N_18619);
nand U25126 (N_25126,N_18053,N_18409);
and U25127 (N_25127,N_18188,N_23250);
and U25128 (N_25128,N_18694,N_23493);
xor U25129 (N_25129,N_19237,N_21028);
xnor U25130 (N_25130,N_21293,N_19804);
and U25131 (N_25131,N_18427,N_18145);
nand U25132 (N_25132,N_23478,N_19338);
and U25133 (N_25133,N_22278,N_20182);
xnor U25134 (N_25134,N_19682,N_20343);
xor U25135 (N_25135,N_22883,N_22321);
xnor U25136 (N_25136,N_23983,N_21508);
nor U25137 (N_25137,N_18081,N_21299);
and U25138 (N_25138,N_20634,N_22684);
or U25139 (N_25139,N_21002,N_22725);
or U25140 (N_25140,N_18170,N_23441);
xnor U25141 (N_25141,N_20904,N_21605);
nor U25142 (N_25142,N_18930,N_18665);
and U25143 (N_25143,N_18543,N_18117);
xor U25144 (N_25144,N_23510,N_20534);
and U25145 (N_25145,N_23662,N_20491);
nor U25146 (N_25146,N_22849,N_23200);
xor U25147 (N_25147,N_19870,N_19916);
nand U25148 (N_25148,N_19198,N_18424);
nor U25149 (N_25149,N_19402,N_23641);
nor U25150 (N_25150,N_19428,N_19084);
nand U25151 (N_25151,N_19800,N_22465);
nor U25152 (N_25152,N_20483,N_19903);
xnor U25153 (N_25153,N_23141,N_20234);
xnor U25154 (N_25154,N_19065,N_21373);
and U25155 (N_25155,N_21562,N_23359);
and U25156 (N_25156,N_23401,N_19448);
nand U25157 (N_25157,N_19547,N_20217);
or U25158 (N_25158,N_19742,N_22453);
or U25159 (N_25159,N_18521,N_18122);
or U25160 (N_25160,N_20872,N_22276);
and U25161 (N_25161,N_18501,N_22022);
and U25162 (N_25162,N_23077,N_19066);
nor U25163 (N_25163,N_19852,N_20071);
nand U25164 (N_25164,N_21091,N_23950);
nor U25165 (N_25165,N_18163,N_18779);
nor U25166 (N_25166,N_22463,N_19436);
xnor U25167 (N_25167,N_22350,N_20304);
and U25168 (N_25168,N_20717,N_20372);
nand U25169 (N_25169,N_22800,N_22449);
nor U25170 (N_25170,N_22242,N_19406);
or U25171 (N_25171,N_20035,N_21676);
nand U25172 (N_25172,N_18591,N_19451);
xnor U25173 (N_25173,N_21768,N_23475);
nand U25174 (N_25174,N_20226,N_18339);
or U25175 (N_25175,N_20845,N_18855);
xor U25176 (N_25176,N_19711,N_22824);
nand U25177 (N_25177,N_20689,N_21085);
and U25178 (N_25178,N_23972,N_19923);
or U25179 (N_25179,N_18680,N_20062);
and U25180 (N_25180,N_21177,N_19172);
nand U25181 (N_25181,N_18709,N_19057);
nand U25182 (N_25182,N_19073,N_18210);
xor U25183 (N_25183,N_23606,N_19438);
and U25184 (N_25184,N_22448,N_23075);
and U25185 (N_25185,N_21434,N_20340);
xor U25186 (N_25186,N_19857,N_21773);
and U25187 (N_25187,N_22423,N_23922);
xor U25188 (N_25188,N_18550,N_23844);
and U25189 (N_25189,N_20543,N_20362);
nor U25190 (N_25190,N_19679,N_20531);
nand U25191 (N_25191,N_21110,N_21747);
nor U25192 (N_25192,N_18911,N_21000);
and U25193 (N_25193,N_21642,N_20601);
xnor U25194 (N_25194,N_23318,N_23266);
xnor U25195 (N_25195,N_18717,N_20118);
and U25196 (N_25196,N_20615,N_20868);
and U25197 (N_25197,N_19155,N_19755);
and U25198 (N_25198,N_19770,N_20567);
xor U25199 (N_25199,N_23723,N_23883);
nand U25200 (N_25200,N_19555,N_18030);
and U25201 (N_25201,N_20604,N_18109);
or U25202 (N_25202,N_18147,N_19489);
and U25203 (N_25203,N_20470,N_19657);
and U25204 (N_25204,N_18638,N_23517);
or U25205 (N_25205,N_21946,N_20771);
xnor U25206 (N_25206,N_18741,N_20351);
or U25207 (N_25207,N_18541,N_22396);
nor U25208 (N_25208,N_21641,N_22351);
and U25209 (N_25209,N_22748,N_20879);
nor U25210 (N_25210,N_22930,N_22787);
nor U25211 (N_25211,N_18004,N_20354);
nand U25212 (N_25212,N_22315,N_22313);
and U25213 (N_25213,N_18193,N_21535);
xor U25214 (N_25214,N_20733,N_18755);
xor U25215 (N_25215,N_22092,N_23030);
nor U25216 (N_25216,N_20200,N_21492);
and U25217 (N_25217,N_23238,N_22957);
xor U25218 (N_25218,N_18569,N_18008);
nor U25219 (N_25219,N_19818,N_20379);
nor U25220 (N_25220,N_21137,N_21926);
xnor U25221 (N_25221,N_18525,N_18559);
nand U25222 (N_25222,N_21162,N_18660);
nand U25223 (N_25223,N_20667,N_18032);
or U25224 (N_25224,N_22369,N_19019);
nor U25225 (N_25225,N_21986,N_19299);
and U25226 (N_25226,N_21011,N_22086);
nand U25227 (N_25227,N_23874,N_19005);
nor U25228 (N_25228,N_23195,N_23837);
or U25229 (N_25229,N_19999,N_19027);
and U25230 (N_25230,N_20935,N_20891);
xnor U25231 (N_25231,N_20983,N_18121);
nand U25232 (N_25232,N_23328,N_21865);
or U25233 (N_25233,N_22175,N_21537);
nor U25234 (N_25234,N_20715,N_18477);
nor U25235 (N_25235,N_22610,N_19308);
and U25236 (N_25236,N_23465,N_22871);
and U25237 (N_25237,N_20533,N_23308);
nor U25238 (N_25238,N_21347,N_22944);
nand U25239 (N_25239,N_20959,N_22807);
or U25240 (N_25240,N_20826,N_19731);
or U25241 (N_25241,N_20711,N_22853);
and U25242 (N_25242,N_19170,N_22362);
nand U25243 (N_25243,N_19562,N_19817);
nor U25244 (N_25244,N_20210,N_19274);
xnor U25245 (N_25245,N_21583,N_18997);
nor U25246 (N_25246,N_19071,N_22247);
nor U25247 (N_25247,N_18691,N_18609);
or U25248 (N_25248,N_20426,N_23103);
nor U25249 (N_25249,N_21061,N_18125);
nand U25250 (N_25250,N_20043,N_19469);
and U25251 (N_25251,N_19571,N_18337);
nor U25252 (N_25252,N_23472,N_19942);
or U25253 (N_25253,N_18568,N_19047);
and U25254 (N_25254,N_18904,N_21872);
xnor U25255 (N_25255,N_20454,N_19421);
and U25256 (N_25256,N_22950,N_21225);
nor U25257 (N_25257,N_19130,N_19914);
xnor U25258 (N_25258,N_22830,N_18594);
nor U25259 (N_25259,N_19690,N_23589);
or U25260 (N_25260,N_19938,N_22401);
nand U25261 (N_25261,N_19069,N_18419);
xor U25262 (N_25262,N_21958,N_21160);
or U25263 (N_25263,N_19619,N_22279);
nand U25264 (N_25264,N_22325,N_21212);
and U25265 (N_25265,N_19449,N_21266);
or U25266 (N_25266,N_21957,N_23817);
nand U25267 (N_25267,N_22167,N_20744);
nand U25268 (N_25268,N_19174,N_21712);
nor U25269 (N_25269,N_19463,N_22105);
nor U25270 (N_25270,N_22028,N_22263);
and U25271 (N_25271,N_20414,N_21144);
xnor U25272 (N_25272,N_23409,N_20373);
and U25273 (N_25273,N_23150,N_19321);
or U25274 (N_25274,N_18531,N_21167);
nor U25275 (N_25275,N_23191,N_18547);
nor U25276 (N_25276,N_20892,N_19747);
xor U25277 (N_25277,N_23135,N_18738);
nand U25278 (N_25278,N_22328,N_19242);
and U25279 (N_25279,N_18233,N_18150);
or U25280 (N_25280,N_18051,N_23527);
or U25281 (N_25281,N_21265,N_22835);
nor U25282 (N_25282,N_19959,N_18653);
and U25283 (N_25283,N_22094,N_21501);
and U25284 (N_25284,N_19970,N_22815);
and U25285 (N_25285,N_21920,N_20896);
or U25286 (N_25286,N_20995,N_21047);
nand U25287 (N_25287,N_21211,N_18518);
or U25288 (N_25288,N_23697,N_22855);
and U25289 (N_25289,N_18708,N_20887);
nand U25290 (N_25290,N_19288,N_22330);
or U25291 (N_25291,N_23334,N_18393);
nand U25292 (N_25292,N_21059,N_20544);
xor U25293 (N_25293,N_18036,N_20921);
xor U25294 (N_25294,N_19475,N_18484);
xor U25295 (N_25295,N_23289,N_19961);
nor U25296 (N_25296,N_21381,N_21393);
xnor U25297 (N_25297,N_23673,N_20000);
and U25298 (N_25298,N_19741,N_23227);
nor U25299 (N_25299,N_18681,N_23698);
nor U25300 (N_25300,N_21959,N_21731);
nor U25301 (N_25301,N_19778,N_22638);
xor U25302 (N_25302,N_18035,N_21332);
nand U25303 (N_25303,N_21009,N_18616);
xnor U25304 (N_25304,N_20064,N_19685);
xnor U25305 (N_25305,N_22927,N_18898);
or U25306 (N_25306,N_22326,N_20121);
nand U25307 (N_25307,N_21639,N_22252);
or U25308 (N_25308,N_21922,N_18141);
xor U25309 (N_25309,N_18219,N_21392);
nor U25310 (N_25310,N_23247,N_21858);
xnor U25311 (N_25311,N_22213,N_21005);
xnor U25312 (N_25312,N_23204,N_18374);
nand U25313 (N_25313,N_19701,N_21797);
nand U25314 (N_25314,N_23001,N_20725);
and U25315 (N_25315,N_22881,N_21511);
xor U25316 (N_25316,N_19860,N_21478);
xnor U25317 (N_25317,N_20357,N_23494);
or U25318 (N_25318,N_23584,N_22427);
nand U25319 (N_25319,N_19810,N_20668);
and U25320 (N_25320,N_22344,N_18824);
nor U25321 (N_25321,N_20646,N_22173);
or U25322 (N_25322,N_21541,N_18271);
nand U25323 (N_25323,N_23161,N_20442);
nor U25324 (N_25324,N_21482,N_19089);
nand U25325 (N_25325,N_19248,N_18587);
and U25326 (N_25326,N_23246,N_20054);
or U25327 (N_25327,N_19422,N_21550);
or U25328 (N_25328,N_21551,N_19887);
or U25329 (N_25329,N_19344,N_22945);
or U25330 (N_25330,N_23533,N_21046);
xnor U25331 (N_25331,N_21039,N_23824);
and U25332 (N_25332,N_20671,N_18929);
xnor U25333 (N_25333,N_20857,N_20677);
nor U25334 (N_25334,N_19981,N_20327);
nor U25335 (N_25335,N_20716,N_20321);
xnor U25336 (N_25336,N_19634,N_21289);
or U25337 (N_25337,N_22745,N_22872);
nand U25338 (N_25338,N_22431,N_22903);
nand U25339 (N_25339,N_21152,N_22232);
xor U25340 (N_25340,N_23355,N_23038);
and U25341 (N_25341,N_19355,N_21054);
or U25342 (N_25342,N_22095,N_21873);
nor U25343 (N_25343,N_23858,N_19978);
nor U25344 (N_25344,N_18556,N_20506);
nor U25345 (N_25345,N_22367,N_20159);
and U25346 (N_25346,N_19176,N_23370);
nand U25347 (N_25347,N_18041,N_20761);
nor U25348 (N_25348,N_19011,N_20699);
nand U25349 (N_25349,N_21006,N_23395);
nor U25350 (N_25350,N_19846,N_21929);
or U25351 (N_25351,N_21145,N_20584);
or U25352 (N_25352,N_23572,N_18814);
and U25353 (N_25353,N_21060,N_18830);
or U25354 (N_25354,N_20805,N_23349);
and U25355 (N_25355,N_19062,N_22917);
or U25356 (N_25356,N_23962,N_20003);
or U25357 (N_25357,N_19165,N_21900);
nand U25358 (N_25358,N_23094,N_23704);
nand U25359 (N_25359,N_22365,N_23217);
or U25360 (N_25360,N_21427,N_20212);
nor U25361 (N_25361,N_23905,N_21433);
and U25362 (N_25362,N_20269,N_23338);
xnor U25363 (N_25363,N_21329,N_21391);
and U25364 (N_25364,N_23818,N_23564);
and U25365 (N_25365,N_22834,N_22544);
xor U25366 (N_25366,N_23688,N_19187);
nand U25367 (N_25367,N_22080,N_23282);
xor U25368 (N_25368,N_21787,N_19757);
nand U25369 (N_25369,N_20466,N_22852);
and U25370 (N_25370,N_18310,N_19957);
and U25371 (N_25371,N_23747,N_21838);
nor U25372 (N_25372,N_19649,N_19454);
nor U25373 (N_25373,N_20774,N_20091);
or U25374 (N_25374,N_22574,N_20138);
or U25375 (N_25375,N_23597,N_23556);
nand U25376 (N_25376,N_20367,N_22828);
xor U25377 (N_25377,N_19822,N_22063);
nand U25378 (N_25378,N_18048,N_18260);
or U25379 (N_25379,N_20221,N_23910);
nand U25380 (N_25380,N_21001,N_19403);
xnor U25381 (N_25381,N_18015,N_19705);
xor U25382 (N_25382,N_18390,N_21796);
nor U25383 (N_25383,N_18007,N_21517);
nand U25384 (N_25384,N_21581,N_20682);
xor U25385 (N_25385,N_20243,N_23323);
or U25386 (N_25386,N_18454,N_21560);
or U25387 (N_25387,N_19381,N_18837);
or U25388 (N_25388,N_21350,N_23258);
nand U25389 (N_25389,N_18721,N_22534);
and U25390 (N_25390,N_19833,N_18906);
nand U25391 (N_25391,N_23274,N_18287);
nand U25392 (N_25392,N_19088,N_18673);
nor U25393 (N_25393,N_23536,N_22868);
nand U25394 (N_25394,N_22205,N_20569);
nor U25395 (N_25395,N_19004,N_18410);
xnor U25396 (N_25396,N_23699,N_23273);
nor U25397 (N_25397,N_19906,N_18654);
xnor U25398 (N_25398,N_19061,N_21674);
nor U25399 (N_25399,N_18719,N_18161);
and U25400 (N_25400,N_21529,N_20581);
and U25401 (N_25401,N_20299,N_18608);
and U25402 (N_25402,N_19576,N_20427);
xor U25403 (N_25403,N_22899,N_20770);
xnor U25404 (N_25404,N_18098,N_18101);
nand U25405 (N_25405,N_19943,N_20542);
and U25406 (N_25406,N_21372,N_18465);
nand U25407 (N_25407,N_23961,N_23806);
nor U25408 (N_25408,N_18793,N_18384);
and U25409 (N_25409,N_18444,N_23761);
xor U25410 (N_25410,N_22218,N_22949);
and U25411 (N_25411,N_22097,N_22874);
xor U25412 (N_25412,N_18341,N_21034);
nor U25413 (N_25413,N_20486,N_19423);
xor U25414 (N_25414,N_18815,N_19689);
nand U25415 (N_25415,N_22122,N_19828);
xnor U25416 (N_25416,N_18398,N_19658);
and U25417 (N_25417,N_19897,N_23674);
nand U25418 (N_25418,N_23502,N_18138);
nor U25419 (N_25419,N_21991,N_18038);
or U25420 (N_25420,N_21275,N_21655);
xor U25421 (N_25421,N_19612,N_23410);
xnor U25422 (N_25422,N_19435,N_21815);
and U25423 (N_25423,N_21113,N_23836);
xor U25424 (N_25424,N_21431,N_19934);
nor U25425 (N_25425,N_18220,N_19714);
nor U25426 (N_25426,N_21037,N_20415);
and U25427 (N_25427,N_23159,N_19345);
or U25428 (N_25428,N_18237,N_19351);
xor U25429 (N_25429,N_23109,N_23678);
nand U25430 (N_25430,N_19637,N_22165);
or U25431 (N_25431,N_21016,N_23029);
or U25432 (N_25432,N_19900,N_22591);
xor U25433 (N_25433,N_20366,N_21572);
nor U25434 (N_25434,N_18118,N_23666);
nand U25435 (N_25435,N_21187,N_21354);
xnor U25436 (N_25436,N_21345,N_20538);
nand U25437 (N_25437,N_19323,N_22865);
and U25438 (N_25438,N_21688,N_20560);
and U25439 (N_25439,N_19894,N_20489);
or U25440 (N_25440,N_18155,N_22965);
and U25441 (N_25441,N_23952,N_21280);
and U25442 (N_25442,N_18634,N_20068);
xnor U25443 (N_25443,N_22587,N_20723);
nand U25444 (N_25444,N_23270,N_18295);
or U25445 (N_25445,N_23428,N_20768);
xnor U25446 (N_25446,N_19713,N_20067);
xor U25447 (N_25447,N_21104,N_18538);
nor U25448 (N_25448,N_18982,N_23108);
nand U25449 (N_25449,N_18311,N_21968);
or U25450 (N_25450,N_18453,N_23460);
xor U25451 (N_25451,N_18492,N_23239);
xor U25452 (N_25452,N_19873,N_18225);
xnor U25453 (N_25453,N_19809,N_22170);
nor U25454 (N_25454,N_21899,N_23314);
and U25455 (N_25455,N_22238,N_18168);
nand U25456 (N_25456,N_18652,N_23228);
or U25457 (N_25457,N_19296,N_23255);
nor U25458 (N_25458,N_22755,N_23911);
nand U25459 (N_25459,N_18656,N_22451);
xor U25460 (N_25460,N_21495,N_23477);
or U25461 (N_25461,N_19527,N_19150);
or U25462 (N_25462,N_18359,N_22433);
or U25463 (N_25463,N_18404,N_20368);
and U25464 (N_25464,N_22728,N_19241);
xnor U25465 (N_25465,N_18812,N_20235);
xnor U25466 (N_25466,N_22223,N_19801);
and U25467 (N_25467,N_23290,N_18326);
or U25468 (N_25468,N_22904,N_20889);
nand U25469 (N_25469,N_19250,N_20565);
and U25470 (N_25470,N_18451,N_23339);
or U25471 (N_25471,N_20128,N_20970);
nand U25472 (N_25472,N_18190,N_18567);
or U25473 (N_25473,N_21951,N_18836);
nor U25474 (N_25474,N_23644,N_19665);
nand U25475 (N_25475,N_18369,N_20174);
nor U25476 (N_25476,N_18561,N_23891);
xor U25477 (N_25477,N_22324,N_19486);
nand U25478 (N_25478,N_22225,N_18978);
xor U25479 (N_25479,N_18180,N_23613);
nand U25480 (N_25480,N_23155,N_23645);
nand U25481 (N_25481,N_19510,N_19728);
nand U25482 (N_25482,N_23188,N_23841);
nand U25483 (N_25483,N_21874,N_20412);
and U25484 (N_25484,N_19441,N_23617);
and U25485 (N_25485,N_18000,N_19572);
nor U25486 (N_25486,N_18771,N_19881);
nand U25487 (N_25487,N_19862,N_19417);
or U25488 (N_25488,N_22710,N_18166);
and U25489 (N_25489,N_20081,N_20740);
xor U25490 (N_25490,N_18861,N_20910);
xnor U25491 (N_25491,N_21753,N_18710);
nor U25492 (N_25492,N_23066,N_18850);
xnor U25493 (N_25493,N_20052,N_21924);
xor U25494 (N_25494,N_19009,N_19168);
xnor U25495 (N_25495,N_21525,N_21514);
or U25496 (N_25496,N_22216,N_22617);
xnor U25497 (N_25497,N_21784,N_20938);
nor U25498 (N_25498,N_18344,N_23224);
xor U25499 (N_25499,N_21288,N_19078);
xor U25500 (N_25500,N_20839,N_18905);
or U25501 (N_25501,N_18099,N_20861);
and U25502 (N_25502,N_22334,N_20585);
and U25503 (N_25503,N_20041,N_23611);
nor U25504 (N_25504,N_20410,N_22340);
or U25505 (N_25505,N_21004,N_23286);
and U25506 (N_25506,N_23126,N_18328);
nand U25507 (N_25507,N_18610,N_22535);
nand U25508 (N_25508,N_23412,N_18416);
nor U25509 (N_25509,N_19085,N_18043);
or U25510 (N_25510,N_21552,N_19813);
xnor U25511 (N_25511,N_23013,N_18124);
nand U25512 (N_25512,N_19848,N_19059);
nand U25513 (N_25513,N_22145,N_23777);
and U25514 (N_25514,N_22825,N_23882);
nor U25515 (N_25515,N_19020,N_23907);
nor U25516 (N_25516,N_18963,N_20076);
or U25517 (N_25517,N_23034,N_18086);
nor U25518 (N_25518,N_23593,N_20692);
xor U25519 (N_25519,N_19988,N_23500);
xnor U25520 (N_25520,N_23492,N_23798);
nand U25521 (N_25521,N_19826,N_22792);
or U25522 (N_25522,N_21051,N_22705);
or U25523 (N_25523,N_20605,N_22632);
nand U25524 (N_25524,N_20659,N_22049);
xnor U25525 (N_25525,N_20397,N_23799);
nor U25526 (N_25526,N_23417,N_21950);
xnor U25527 (N_25527,N_20873,N_18767);
nand U25528 (N_25528,N_20960,N_20813);
or U25529 (N_25529,N_21374,N_20926);
nor U25530 (N_25530,N_23684,N_20332);
nor U25531 (N_25531,N_19861,N_22877);
and U25532 (N_25532,N_20413,N_20992);
xnor U25533 (N_25533,N_18440,N_19218);
or U25534 (N_25534,N_18866,N_18378);
or U25535 (N_25535,N_21811,N_23032);
nor U25536 (N_25536,N_23398,N_23582);
xor U25537 (N_25537,N_19034,N_23260);
or U25538 (N_25538,N_21891,N_22271);
nor U25539 (N_25539,N_21032,N_20808);
nor U25540 (N_25540,N_21227,N_21795);
xnor U25541 (N_25541,N_19064,N_22553);
or U25542 (N_25542,N_21568,N_19513);
nand U25543 (N_25543,N_22380,N_20971);
nand U25544 (N_25544,N_23450,N_20198);
or U25545 (N_25545,N_22723,N_23898);
or U25546 (N_25546,N_18386,N_22649);
and U25547 (N_25547,N_18371,N_19138);
and U25548 (N_25548,N_19908,N_19466);
and U25549 (N_25549,N_21123,N_20502);
nor U25550 (N_25550,N_20844,N_18014);
or U25551 (N_25551,N_22048,N_21515);
nand U25552 (N_25552,N_18208,N_23002);
nand U25553 (N_25553,N_19918,N_22976);
xnor U25554 (N_25554,N_19032,N_20732);
xor U25555 (N_25555,N_20123,N_20500);
or U25556 (N_25556,N_19413,N_22704);
or U25557 (N_25557,N_21686,N_22461);
nor U25558 (N_25558,N_18055,N_18600);
nand U25559 (N_25559,N_20811,N_21931);
and U25560 (N_25560,N_20994,N_21683);
nor U25561 (N_25561,N_22637,N_21748);
and U25562 (N_25562,N_18365,N_21947);
and U25563 (N_25563,N_21786,N_20488);
nand U25564 (N_25564,N_20322,N_20863);
or U25565 (N_25565,N_23033,N_20049);
xnor U25566 (N_25566,N_20156,N_20433);
xor U25567 (N_25567,N_21880,N_21910);
nor U25568 (N_25568,N_18119,N_23303);
xor U25569 (N_25569,N_22265,N_21301);
or U25570 (N_25570,N_19124,N_21505);
xnor U25571 (N_25571,N_23348,N_21735);
nand U25572 (N_25572,N_23243,N_19591);
or U25573 (N_25573,N_20912,N_22914);
nand U25574 (N_25574,N_19505,N_20485);
or U25575 (N_25575,N_19962,N_19954);
or U25576 (N_25576,N_18764,N_18598);
nand U25577 (N_25577,N_22301,N_23727);
or U25578 (N_25578,N_21284,N_23252);
nor U25579 (N_25579,N_21115,N_23894);
nor U25580 (N_25580,N_18724,N_23383);
xor U25581 (N_25581,N_20286,N_19627);
or U25582 (N_25582,N_19184,N_20907);
nand U25583 (N_25583,N_19593,N_18956);
xnor U25584 (N_25584,N_18265,N_18644);
nor U25585 (N_25585,N_18346,N_23320);
xor U25586 (N_25586,N_19023,N_20847);
xor U25587 (N_25587,N_21439,N_18909);
nor U25588 (N_25588,N_19867,N_19641);
nand U25589 (N_25589,N_21063,N_20819);
or U25590 (N_25590,N_23661,N_22565);
xor U25591 (N_25591,N_22413,N_20654);
xor U25592 (N_25592,N_19458,N_22856);
nor U25593 (N_25593,N_21921,N_22140);
and U25594 (N_25594,N_18763,N_20803);
xor U25595 (N_25595,N_21042,N_22973);
nor U25596 (N_25596,N_20255,N_22594);
or U25597 (N_25597,N_18841,N_18498);
xor U25598 (N_25598,N_18969,N_23298);
and U25599 (N_25599,N_23811,N_23872);
xnor U25600 (N_25600,N_20537,N_18632);
nand U25601 (N_25601,N_21507,N_20171);
and U25602 (N_25602,N_22822,N_22146);
and U25603 (N_25603,N_23202,N_23267);
and U25604 (N_25604,N_18461,N_20213);
nand U25605 (N_25605,N_22827,N_18497);
or U25606 (N_25606,N_22288,N_23769);
and U25607 (N_25607,N_20053,N_18713);
xor U25608 (N_25608,N_21894,N_18293);
nor U25609 (N_25609,N_18674,N_19795);
xor U25610 (N_25610,N_22779,N_21400);
nand U25611 (N_25611,N_21805,N_21200);
and U25612 (N_25612,N_21058,N_20098);
or U25613 (N_25613,N_22691,N_21544);
nand U25614 (N_25614,N_18821,N_18275);
nand U25615 (N_25615,N_21772,N_18095);
xor U25616 (N_25616,N_19002,N_20338);
or U25617 (N_25617,N_20974,N_19398);
nand U25618 (N_25618,N_23037,N_22079);
nor U25619 (N_25619,N_23169,N_19091);
or U25620 (N_25620,N_20618,N_19035);
nor U25621 (N_25621,N_23691,N_23052);
or U25622 (N_25622,N_18403,N_23120);
or U25623 (N_25623,N_20882,N_21198);
xor U25624 (N_25624,N_18589,N_18089);
or U25625 (N_25625,N_18433,N_18750);
xor U25626 (N_25626,N_19972,N_21604);
and U25627 (N_25627,N_18645,N_21637);
or U25628 (N_25628,N_20444,N_21917);
nand U25629 (N_25629,N_22306,N_21460);
nand U25630 (N_25630,N_18267,N_21453);
nand U25631 (N_25631,N_21566,N_19046);
nor U25632 (N_25632,N_23941,N_22217);
and U25633 (N_25633,N_20337,N_19788);
xor U25634 (N_25634,N_19206,N_18469);
nor U25635 (N_25635,N_20951,N_22668);
or U25636 (N_25636,N_18509,N_21396);
and U25637 (N_25637,N_21829,N_22057);
nor U25638 (N_25638,N_22689,N_19926);
xnor U25639 (N_25639,N_22597,N_20355);
nand U25640 (N_25640,N_20685,N_19723);
and U25641 (N_25641,N_22885,N_19239);
nand U25642 (N_25642,N_21040,N_22224);
and U25643 (N_25643,N_21824,N_23110);
nand U25644 (N_25644,N_19774,N_21328);
or U25645 (N_25645,N_20642,N_19785);
nand U25646 (N_25646,N_20215,N_19158);
nor U25647 (N_25647,N_23751,N_20289);
nor U25648 (N_25648,N_20072,N_20353);
xor U25649 (N_25649,N_21030,N_19920);
xnor U25650 (N_25650,N_19533,N_22919);
and U25651 (N_25651,N_20395,N_20984);
nor U25652 (N_25652,N_21690,N_21519);
nor U25653 (N_25653,N_23099,N_21143);
xnor U25654 (N_25654,N_21100,N_19587);
xor U25655 (N_25655,N_19712,N_19752);
nor U25656 (N_25656,N_19816,N_23199);
or U25657 (N_25657,N_19573,N_21668);
or U25658 (N_25658,N_21949,N_22428);
nor U25659 (N_25659,N_21509,N_23854);
nand U25660 (N_25660,N_18452,N_18618);
nand U25661 (N_25661,N_23364,N_18540);
xnor U25662 (N_25662,N_22089,N_20342);
or U25663 (N_25663,N_20326,N_23851);
and U25664 (N_25664,N_23871,N_19213);
or U25665 (N_25665,N_20266,N_21607);
and U25666 (N_25666,N_23866,N_22589);
and U25667 (N_25667,N_19115,N_19837);
and U25668 (N_25668,N_21989,N_23024);
or U25669 (N_25669,N_19146,N_20023);
nand U25670 (N_25670,N_23736,N_20728);
nand U25671 (N_25671,N_18958,N_23208);
and U25672 (N_25672,N_20300,N_22370);
xor U25673 (N_25673,N_19121,N_20220);
and U25674 (N_25674,N_21050,N_18515);
and U25675 (N_25675,N_23807,N_23759);
and U25676 (N_25676,N_23095,N_21385);
nand U25677 (N_25677,N_18206,N_20718);
nand U25678 (N_25678,N_18478,N_20173);
xor U25679 (N_25679,N_23335,N_19107);
or U25680 (N_25680,N_23469,N_20075);
or U25681 (N_25681,N_20752,N_20319);
or U25682 (N_25682,N_21095,N_22241);
nand U25683 (N_25683,N_18980,N_23003);
xor U25684 (N_25684,N_22354,N_20112);
nor U25685 (N_25685,N_21665,N_20656);
nor U25686 (N_25686,N_21892,N_21281);
nand U25687 (N_25687,N_19525,N_19255);
nand U25688 (N_25688,N_18482,N_22920);
nand U25689 (N_25689,N_18852,N_22447);
or U25690 (N_25690,N_23763,N_23294);
nand U25691 (N_25691,N_18939,N_22997);
or U25692 (N_25692,N_19151,N_20526);
and U25693 (N_25693,N_18588,N_22397);
and U25694 (N_25694,N_19569,N_19675);
xnor U25695 (N_25695,N_18288,N_18269);
and U25696 (N_25696,N_19784,N_21800);
and U25697 (N_25697,N_22624,N_22331);
xor U25698 (N_25698,N_23036,N_20925);
xor U25699 (N_25699,N_18895,N_23752);
nor U25700 (N_25700,N_23106,N_18643);
and U25701 (N_25701,N_22303,N_20832);
nor U25702 (N_25702,N_18565,N_20017);
and U25703 (N_25703,N_20036,N_18539);
xnor U25704 (N_25704,N_23205,N_19139);
nor U25705 (N_25705,N_19110,N_23948);
and U25706 (N_25706,N_21147,N_22793);
and U25707 (N_25707,N_21132,N_20541);
or U25708 (N_25708,N_20576,N_19950);
nand U25709 (N_25709,N_20934,N_23540);
nor U25710 (N_25710,N_19618,N_20778);
or U25711 (N_25711,N_22336,N_22522);
xnor U25712 (N_25712,N_18085,N_19082);
nand U25713 (N_25713,N_19251,N_22181);
nand U25714 (N_25714,N_21135,N_19883);
or U25715 (N_25715,N_23373,N_22826);
or U25716 (N_25716,N_20695,N_21778);
or U25717 (N_25717,N_19904,N_18381);
and U25718 (N_25718,N_23163,N_22222);
nor U25719 (N_25719,N_22665,N_23481);
or U25720 (N_25720,N_22494,N_19278);
xor U25721 (N_25721,N_18171,N_20979);
nand U25722 (N_25722,N_22029,N_18872);
nor U25723 (N_25723,N_19016,N_18351);
nand U25724 (N_25724,N_19086,N_18780);
and U25725 (N_25725,N_19738,N_23305);
xnor U25726 (N_25726,N_21222,N_19508);
and U25727 (N_25727,N_22607,N_20238);
and U25728 (N_25728,N_20329,N_20042);
xor U25729 (N_25729,N_18952,N_21576);
nand U25730 (N_25730,N_19985,N_22527);
and U25731 (N_25731,N_21631,N_18627);
or U25732 (N_25732,N_20888,N_22939);
and U25733 (N_25733,N_21203,N_21956);
xor U25734 (N_25734,N_19550,N_20977);
or U25735 (N_25735,N_20905,N_19969);
or U25736 (N_25736,N_20523,N_19026);
xor U25737 (N_25737,N_21578,N_18933);
and U25738 (N_25738,N_23354,N_20796);
nor U25739 (N_25739,N_22438,N_18485);
xor U25740 (N_25740,N_18357,N_21744);
and U25741 (N_25741,N_18302,N_19434);
nor U25742 (N_25742,N_22718,N_20002);
nor U25743 (N_25743,N_23071,N_22337);
and U25744 (N_25744,N_19133,N_18798);
xor U25745 (N_25745,N_23568,N_20838);
or U25746 (N_25746,N_19866,N_21779);
nor U25747 (N_25747,N_19500,N_23878);
nor U25748 (N_25748,N_20684,N_22940);
and U25749 (N_25749,N_18988,N_18825);
nor U25750 (N_25750,N_20603,N_21026);
and U25751 (N_25751,N_20875,N_23242);
nor U25752 (N_25752,N_21911,N_20899);
or U25753 (N_25753,N_21548,N_23892);
nor U25754 (N_25754,N_19356,N_20837);
xor U25755 (N_25755,N_22117,N_19259);
nor U25756 (N_25756,N_23779,N_23996);
or U25757 (N_25757,N_18029,N_22399);
xor U25758 (N_25758,N_23921,N_20022);
and U25759 (N_25759,N_20496,N_22778);
xnor U25760 (N_25760,N_21425,N_19293);
nand U25761 (N_25761,N_20160,N_20436);
and U25762 (N_25762,N_22910,N_22045);
or U25763 (N_25763,N_20025,N_18207);
or U25764 (N_25764,N_22862,N_20840);
nand U25765 (N_25765,N_18688,N_20797);
nor U25766 (N_25766,N_20388,N_20701);
nand U25767 (N_25767,N_18880,N_22307);
nor U25768 (N_25768,N_21763,N_23598);
nor U25769 (N_25769,N_19191,N_22261);
nor U25770 (N_25770,N_21376,N_22052);
xnor U25771 (N_25771,N_22730,N_22669);
or U25772 (N_25772,N_23553,N_20051);
xnor U25773 (N_25773,N_21031,N_20318);
xnor U25774 (N_25774,N_21531,N_23271);
xor U25775 (N_25775,N_22481,N_19311);
xor U25776 (N_25776,N_23307,N_19528);
nor U25777 (N_25777,N_18175,N_22214);
nor U25778 (N_25778,N_23411,N_22112);
or U25779 (N_25779,N_19995,N_18284);
xor U25780 (N_25780,N_19491,N_20895);
or U25781 (N_25781,N_19113,N_22227);
nand U25782 (N_25782,N_20674,N_21842);
nor U25783 (N_25783,N_21933,N_23765);
nand U25784 (N_25784,N_21569,N_20130);
nor U25785 (N_25785,N_21634,N_20644);
nand U25786 (N_25786,N_21242,N_21976);
and U25787 (N_25787,N_20933,N_20048);
xor U25788 (N_25788,N_21593,N_21919);
and U25789 (N_25789,N_21331,N_20622);
and U25790 (N_25790,N_19185,N_23653);
xor U25791 (N_25791,N_19672,N_18418);
nor U25792 (N_25792,N_20645,N_19827);
xor U25793 (N_25793,N_19099,N_19395);
or U25794 (N_25794,N_19888,N_23513);
xor U25795 (N_25795,N_20095,N_23455);
xnor U25796 (N_25796,N_19937,N_20755);
and U25797 (N_25797,N_18436,N_19173);
xor U25798 (N_25798,N_23374,N_21029);
and U25799 (N_25799,N_23686,N_20060);
nor U25800 (N_25800,N_23296,N_18977);
nand U25801 (N_25801,N_22183,N_19166);
and U25802 (N_25802,N_19805,N_18298);
nand U25803 (N_25803,N_20046,N_22148);
xor U25804 (N_25804,N_23376,N_18185);
nand U25805 (N_25805,N_19253,N_21220);
xnor U25806 (N_25806,N_19203,N_18934);
xnor U25807 (N_25807,N_23474,N_19269);
nand U25808 (N_25808,N_21149,N_22516);
nor U25809 (N_25809,N_23025,N_22394);
nor U25810 (N_25810,N_18597,N_21094);
nor U25811 (N_25811,N_22457,N_20554);
or U25812 (N_25812,N_19597,N_21173);
xor U25813 (N_25813,N_18083,N_19024);
or U25814 (N_25814,N_20736,N_23219);
nor U25815 (N_25815,N_20194,N_21774);
nand U25816 (N_25816,N_23375,N_23544);
and U25817 (N_25817,N_22850,N_18966);
or U25818 (N_25818,N_20229,N_18411);
and U25819 (N_25819,N_21362,N_18792);
nand U25820 (N_25820,N_21188,N_19464);
nand U25821 (N_25821,N_21468,N_19263);
xnor U25822 (N_25822,N_22372,N_22053);
or U25823 (N_25823,N_20259,N_21648);
and U25824 (N_25824,N_19178,N_22108);
nor U25825 (N_25825,N_18844,N_22035);
or U25826 (N_25826,N_19684,N_20947);
nor U25827 (N_25827,N_21219,N_18329);
nor U25828 (N_25828,N_23028,N_21241);
nor U25829 (N_25829,N_22493,N_18503);
nor U25830 (N_25830,N_18113,N_22379);
nand U25831 (N_25831,N_20800,N_18987);
nor U25832 (N_25832,N_20720,N_19230);
and U25833 (N_25833,N_22968,N_20236);
and U25834 (N_25834,N_20587,N_18047);
nand U25835 (N_25835,N_23496,N_23633);
xnor U25836 (N_25836,N_22104,N_20853);
or U25837 (N_25837,N_19674,N_22988);
xnor U25838 (N_25838,N_21777,N_22931);
xor U25839 (N_25839,N_23506,N_18132);
nand U25840 (N_25840,N_23079,N_20507);
or U25841 (N_25841,N_22762,N_19162);
and U25842 (N_25842,N_19541,N_19148);
and U25843 (N_25843,N_21138,N_23800);
and U25844 (N_25844,N_20453,N_21758);
xnor U25845 (N_25845,N_18261,N_20018);
and U25846 (N_25846,N_18663,N_21575);
or U25847 (N_25847,N_19497,N_18586);
or U25848 (N_25848,N_20001,N_18936);
and U25849 (N_25849,N_22101,N_21489);
or U25850 (N_25850,N_23309,N_21166);
nand U25851 (N_25851,N_23549,N_21937);
or U25852 (N_25852,N_19515,N_20135);
or U25853 (N_25853,N_18520,N_22963);
nand U25854 (N_25854,N_22708,N_18388);
and U25855 (N_25855,N_22467,N_19990);
or U25856 (N_25856,N_18886,N_23828);
nand U25857 (N_25857,N_18146,N_20009);
nor U25858 (N_25858,N_18908,N_23771);
nand U25859 (N_25859,N_22681,N_19309);
nand U25860 (N_25860,N_18927,N_21007);
and U25861 (N_25861,N_23971,N_18445);
and U25862 (N_25862,N_22538,N_18544);
nand U25863 (N_25863,N_23121,N_22149);
nor U25864 (N_25864,N_18049,N_18126);
or U25865 (N_25865,N_18916,N_20788);
and U25866 (N_25866,N_18917,N_18088);
and U25867 (N_25867,N_23457,N_20694);
nor U25868 (N_25868,N_20599,N_23930);
nand U25869 (N_25869,N_18944,N_20424);
and U25870 (N_25870,N_18757,N_18250);
or U25871 (N_25871,N_20020,N_18794);
and U25872 (N_25872,N_20457,N_21983);
or U25873 (N_25873,N_22024,N_21715);
nand U25874 (N_25874,N_20730,N_23489);
nand U25875 (N_25875,N_19601,N_22907);
nand U25876 (N_25876,N_18945,N_19925);
and U25877 (N_25877,N_21055,N_22657);
xor U25878 (N_25878,N_21966,N_21470);
xor U25879 (N_25879,N_22869,N_23479);
nand U25880 (N_25880,N_21806,N_19604);
xnor U25881 (N_25881,N_18330,N_18949);
and U25882 (N_25882,N_20482,N_22174);
xnor U25883 (N_25883,N_21942,N_21246);
xnor U25884 (N_25884,N_20459,N_20151);
and U25885 (N_25885,N_20292,N_18129);
and U25886 (N_25886,N_21428,N_22384);
nor U25887 (N_25887,N_21589,N_18415);
or U25888 (N_25888,N_22123,N_18995);
nor U25889 (N_25889,N_21202,N_18718);
nand U25890 (N_25890,N_22584,N_20471);
nand U25891 (N_25891,N_20807,N_22245);
and U25892 (N_25892,N_20734,N_21549);
nand U25893 (N_25893,N_23868,N_18554);
nand U25894 (N_25894,N_18324,N_20782);
xor U25895 (N_25895,N_19424,N_22683);
and U25896 (N_25896,N_18998,N_23627);
nor U25897 (N_25897,N_19042,N_21239);
nand U25898 (N_25898,N_22129,N_22103);
nand U25899 (N_25899,N_20203,N_23016);
or U25900 (N_25900,N_19610,N_18027);
nor U25901 (N_25901,N_19264,N_21473);
and U25902 (N_25902,N_23604,N_19105);
and U25903 (N_25903,N_18811,N_23997);
xor U25904 (N_25904,N_19072,N_19736);
or U25905 (N_25905,N_20529,N_20307);
or U25906 (N_25906,N_21340,N_19520);
nand U25907 (N_25907,N_22488,N_22355);
nor U25908 (N_25908,N_22499,N_21322);
nor U25909 (N_25909,N_18361,N_22751);
nand U25910 (N_25910,N_21083,N_20998);
nand U25911 (N_25911,N_20597,N_19396);
nand U25912 (N_25912,N_19493,N_23649);
nor U25913 (N_25913,N_18333,N_22616);
nor U25914 (N_25914,N_23552,N_21496);
nor U25915 (N_25915,N_18259,N_18506);
and U25916 (N_25916,N_21338,N_21443);
nand U25917 (N_25917,N_22347,N_18833);
or U25918 (N_25918,N_19081,N_21948);
nor U25919 (N_25919,N_18184,N_20404);
and U25920 (N_25920,N_22302,N_20375);
nor U25921 (N_25921,N_22857,N_18123);
and U25922 (N_25922,N_19652,N_18537);
nand U25923 (N_25923,N_18115,N_20297);
nor U25924 (N_25924,N_23495,N_21230);
or U25925 (N_25925,N_21417,N_20814);
xor U25926 (N_25926,N_21483,N_21901);
nor U25927 (N_25927,N_18034,N_23934);
xor U25928 (N_25928,N_18280,N_18940);
and U25929 (N_25929,N_22041,N_18926);
nor U25930 (N_25930,N_18650,N_23538);
nor U25931 (N_25931,N_22537,N_19620);
xor U25932 (N_25932,N_18426,N_18699);
xnor U25933 (N_25933,N_18517,N_21685);
or U25934 (N_25934,N_19706,N_19913);
nand U25935 (N_25935,N_18127,N_18283);
xnor U25936 (N_25936,N_22991,N_19781);
xor U25937 (N_25937,N_22257,N_20939);
or U25938 (N_25938,N_18272,N_23577);
or U25939 (N_25939,N_20915,N_23369);
or U25940 (N_25940,N_20688,N_22168);
or U25941 (N_25941,N_22468,N_22528);
nor U25942 (N_25942,N_18466,N_19452);
and U25943 (N_25943,N_19298,N_20964);
xnor U25944 (N_25944,N_23237,N_21792);
nor U25945 (N_25945,N_19056,N_21254);
and U25946 (N_25946,N_18513,N_19582);
nand U25947 (N_25947,N_20864,N_18630);
nand U25948 (N_25948,N_18878,N_19829);
and U25949 (N_25949,N_19277,N_19739);
or U25950 (N_25950,N_19911,N_21539);
and U25951 (N_25951,N_19171,N_21412);
and U25952 (N_25952,N_19708,N_23297);
xnor U25953 (N_25953,N_19415,N_23550);
xor U25954 (N_25954,N_21099,N_20655);
or U25955 (N_25955,N_21027,N_20616);
or U25956 (N_25956,N_21707,N_21934);
xnor U25957 (N_25957,N_23945,N_19083);
nand U25958 (N_25958,N_18160,N_20107);
nor U25959 (N_25959,N_19033,N_21905);
nor U25960 (N_25960,N_19212,N_21682);
nand U25961 (N_25961,N_18932,N_19179);
nand U25962 (N_25962,N_22166,N_23612);
xor U25963 (N_25963,N_22050,N_18187);
and U25964 (N_25964,N_18254,N_21477);
nor U25965 (N_25965,N_23027,N_23480);
and U25966 (N_25966,N_23846,N_19376);
nand U25967 (N_25967,N_19159,N_18527);
nor U25968 (N_25968,N_23439,N_22682);
nor U25969 (N_25969,N_23512,N_19022);
or U25970 (N_25970,N_22760,N_18602);
xnor U25971 (N_25971,N_20940,N_19763);
nor U25972 (N_25972,N_20681,N_18983);
xor U25973 (N_25973,N_19732,N_18472);
nand U25974 (N_25974,N_21012,N_21793);
or U25975 (N_25975,N_23791,N_19220);
and U25976 (N_25976,N_22065,N_21879);
and U25977 (N_25977,N_23957,N_22150);
nand U25978 (N_25978,N_21045,N_23680);
and U25979 (N_25979,N_23974,N_21256);
and U25980 (N_25980,N_20765,N_21799);
nor U25981 (N_25981,N_20927,N_20871);
nand U25982 (N_25982,N_22505,N_22974);
xnor U25983 (N_25983,N_21555,N_19735);
or U25984 (N_25984,N_22614,N_18285);
or U25985 (N_25985,N_22746,N_19891);
xor U25986 (N_25986,N_18063,N_19390);
or U25987 (N_25987,N_19215,N_18242);
or U25988 (N_25988,N_21699,N_22972);
or U25989 (N_25989,N_18321,N_18213);
xnor U25990 (N_25990,N_18740,N_18301);
nor U25991 (N_25991,N_23741,N_18595);
or U25992 (N_25992,N_18186,N_20481);
xor U25993 (N_25993,N_20937,N_20573);
nand U25994 (N_25994,N_21553,N_21101);
and U25995 (N_25995,N_23965,N_19884);
and U25996 (N_25996,N_19676,N_19118);
nand U25997 (N_25997,N_22498,N_19431);
and U25998 (N_25998,N_19342,N_21996);
and U25999 (N_25999,N_18946,N_22648);
xnor U26000 (N_26000,N_20476,N_22339);
or U26001 (N_26001,N_22529,N_20709);
nand U26002 (N_26002,N_19691,N_19285);
nand U26003 (N_26003,N_18620,N_19000);
or U26004 (N_26004,N_23174,N_19223);
nor U26005 (N_26005,N_23087,N_23435);
and U26006 (N_26006,N_21847,N_18078);
nor U26007 (N_26007,N_23977,N_23124);
nor U26008 (N_26008,N_20809,N_21710);
xor U26009 (N_26009,N_21021,N_22829);
xor U26010 (N_26010,N_23288,N_23712);
xnor U26011 (N_26011,N_22503,N_22479);
nand U26012 (N_26012,N_20916,N_22374);
and U26013 (N_26013,N_21379,N_20874);
xnor U26014 (N_26014,N_19317,N_22154);
or U26015 (N_26015,N_23272,N_21403);
and U26016 (N_26016,N_22377,N_19878);
nor U26017 (N_26017,N_19614,N_21828);
nand U26018 (N_26018,N_21335,N_23218);
and U26019 (N_26019,N_19370,N_18875);
xor U26020 (N_26020,N_20806,N_18136);
nor U26021 (N_26021,N_20588,N_20218);
nor U26022 (N_26022,N_20946,N_22195);
nor U26023 (N_26023,N_20131,N_21713);
nand U26024 (N_26024,N_23696,N_23746);
and U26025 (N_26025,N_21617,N_20133);
or U26026 (N_26026,N_21472,N_18658);
or U26027 (N_26027,N_20396,N_20111);
or U26028 (N_26028,N_21759,N_21304);
or U26029 (N_26029,N_19408,N_22440);
nor U26030 (N_26030,N_23529,N_20949);
nand U26031 (N_26031,N_23652,N_18702);
or U26032 (N_26032,N_22578,N_19681);
or U26033 (N_26033,N_22403,N_18847);
or U26034 (N_26034,N_21494,N_18164);
nor U26035 (N_26035,N_18020,N_18075);
nand U26036 (N_26036,N_20821,N_18114);
nand U26037 (N_26037,N_18222,N_23047);
or U26038 (N_26038,N_20515,N_18322);
xnor U26039 (N_26039,N_22151,N_19976);
or U26040 (N_26040,N_22521,N_23964);
or U26041 (N_26041,N_21049,N_21524);
nor U26042 (N_26042,N_18158,N_23748);
and U26043 (N_26043,N_22404,N_23862);
xnor U26044 (N_26044,N_23843,N_21457);
nor U26045 (N_26045,N_19270,N_19097);
nor U26046 (N_26046,N_22442,N_21716);
or U26047 (N_26047,N_18823,N_18555);
nand U26048 (N_26048,N_19364,N_21696);
nand U26049 (N_26049,N_23019,N_19354);
xor U26050 (N_26050,N_22775,N_22697);
xor U26051 (N_26051,N_22727,N_22545);
nor U26052 (N_26052,N_22402,N_18396);
xnor U26053 (N_26053,N_18251,N_18491);
xnor U26054 (N_26054,N_23415,N_23607);
nor U26055 (N_26055,N_19319,N_18848);
nor U26056 (N_26056,N_22297,N_22785);
and U26057 (N_26057,N_19740,N_18058);
and U26058 (N_26058,N_23051,N_18832);
or U26059 (N_26059,N_21849,N_23322);
and U26060 (N_26060,N_19640,N_21459);
or U26061 (N_26061,N_23092,N_18350);
and U26062 (N_26062,N_19965,N_20178);
and U26063 (N_26063,N_23010,N_20038);
nor U26064 (N_26064,N_22912,N_22818);
or U26065 (N_26065,N_18807,N_18076);
nor U26066 (N_26066,N_19063,N_20673);
and U26067 (N_26067,N_20555,N_23132);
nand U26068 (N_26068,N_22361,N_23044);
nor U26069 (N_26069,N_22487,N_20291);
nand U26070 (N_26070,N_19093,N_18573);
nor U26071 (N_26071,N_21518,N_21312);
nand U26072 (N_26072,N_22742,N_18813);
nand U26073 (N_26073,N_19141,N_23902);
xor U26074 (N_26074,N_21413,N_21402);
or U26075 (N_26075,N_22788,N_18022);
nand U26076 (N_26076,N_18684,N_18031);
nor U26077 (N_26077,N_19339,N_20127);
nor U26078 (N_26078,N_20445,N_20854);
xnor U26079 (N_26079,N_20816,N_18760);
or U26080 (N_26080,N_22246,N_20087);
nand U26081 (N_26081,N_19707,N_21855);
xor U26082 (N_26082,N_19603,N_21182);
nor U26083 (N_26083,N_22812,N_21065);
and U26084 (N_26084,N_23302,N_21172);
xnor U26085 (N_26085,N_23808,N_20672);
and U26086 (N_26086,N_23143,N_23209);
or U26087 (N_26087,N_22509,N_20913);
xnor U26088 (N_26088,N_19391,N_22497);
and U26089 (N_26089,N_20922,N_18720);
and U26090 (N_26090,N_19843,N_23602);
and U26091 (N_26091,N_19696,N_19858);
nand U26092 (N_26092,N_19460,N_19748);
and U26093 (N_26093,N_21640,N_19360);
nor U26094 (N_26094,N_22776,N_22127);
xor U26095 (N_26095,N_18677,N_21818);
nor U26096 (N_26096,N_20461,N_21080);
nand U26097 (N_26097,N_21852,N_22277);
nand U26098 (N_26098,N_21883,N_19948);
nand U26099 (N_26099,N_23739,N_18179);
nand U26100 (N_26100,N_23485,N_23043);
nand U26101 (N_26101,N_22158,N_20411);
nor U26102 (N_26102,N_22539,N_22017);
nor U26103 (N_26103,N_19560,N_18107);
or U26104 (N_26104,N_22425,N_21863);
and U26105 (N_26105,N_21740,N_22036);
and U26106 (N_26106,N_21789,N_22500);
or U26107 (N_26107,N_23935,N_20954);
nor U26108 (N_26108,N_18005,N_18297);
xor U26109 (N_26109,N_19777,N_23557);
or U26110 (N_26110,N_20463,N_22139);
xnor U26111 (N_26111,N_22378,N_22946);
nand U26112 (N_26112,N_18868,N_18064);
and U26113 (N_26113,N_20129,N_18626);
xnor U26114 (N_26114,N_18840,N_23581);
or U26115 (N_26115,N_20478,N_19348);
and U26116 (N_26116,N_18557,N_18954);
xor U26117 (N_26117,N_21890,N_23565);
and U26118 (N_26118,N_22411,N_18013);
nand U26119 (N_26119,N_20518,N_18582);
nor U26120 (N_26120,N_22352,N_18446);
xnor U26121 (N_26121,N_21397,N_20658);
xnor U26122 (N_26122,N_19101,N_20176);
nor U26123 (N_26123,N_22285,N_23381);
xnor U26124 (N_26124,N_18428,N_23953);
or U26125 (N_26125,N_18087,N_23213);
or U26126 (N_26126,N_23507,N_21851);
xor U26127 (N_26127,N_19195,N_18335);
nand U26128 (N_26128,N_19812,N_19653);
or U26129 (N_26129,N_20691,N_18993);
nand U26130 (N_26130,N_21273,N_21249);
nand U26131 (N_26131,N_18366,N_22551);
and U26132 (N_26132,N_22837,N_18857);
and U26133 (N_26133,N_21209,N_21178);
xnor U26134 (N_26134,N_22417,N_20917);
nand U26135 (N_26135,N_21387,N_20132);
or U26136 (N_26136,N_21493,N_23576);
nand U26137 (N_26137,N_23760,N_20520);
nand U26138 (N_26138,N_21621,N_22391);
and U26139 (N_26139,N_19673,N_20423);
nor U26140 (N_26140,N_19775,N_22100);
nor U26141 (N_26141,N_21836,N_23186);
xor U26142 (N_26142,N_19504,N_22533);
or U26143 (N_26143,N_22273,N_20621);
and U26144 (N_26144,N_23621,N_23993);
nand U26145 (N_26145,N_20333,N_18379);
nand U26146 (N_26146,N_22207,N_21563);
and U26147 (N_26147,N_21078,N_22536);
nor U26148 (N_26148,N_23991,N_23619);
nor U26149 (N_26149,N_19410,N_19487);
nand U26150 (N_26150,N_23350,N_18795);
nor U26151 (N_26151,N_23978,N_23463);
xor U26152 (N_26152,N_18971,N_21729);
nor U26153 (N_26153,N_18831,N_21330);
nand U26154 (N_26154,N_23065,N_19789);
nand U26155 (N_26155,N_19994,N_19227);
nand U26156 (N_26156,N_21971,N_21435);
and U26157 (N_26157,N_21869,N_19524);
nor U26158 (N_26158,N_18545,N_19624);
and U26159 (N_26159,N_21326,N_23078);
nand U26160 (N_26160,N_22096,N_21684);
nand U26161 (N_26161,N_23130,N_21709);
nor U26162 (N_26162,N_19273,N_23814);
nor U26163 (N_26163,N_19764,N_18581);
and U26164 (N_26164,N_22923,N_21751);
or U26165 (N_26165,N_19710,N_22663);
or U26166 (N_26166,N_22598,N_19051);
or U26167 (N_26167,N_18716,N_18614);
xnor U26168 (N_26168,N_19496,N_20228);
nor U26169 (N_26169,N_21887,N_20451);
nand U26170 (N_26170,N_19030,N_18450);
nand U26171 (N_26171,N_19169,N_21126);
nor U26172 (N_26172,N_22567,N_21619);
xor U26173 (N_26173,N_23085,N_22971);
nor U26174 (N_26174,N_22555,N_23656);
xnor U26175 (N_26175,N_20897,N_19459);
or U26176 (N_26176,N_21165,N_18791);
nand U26177 (N_26177,N_20747,N_20784);
xnor U26178 (N_26178,N_19841,N_21024);
and U26179 (N_26179,N_19823,N_19389);
xnor U26180 (N_26180,N_20474,N_19964);
or U26181 (N_26181,N_19399,N_18399);
nor U26182 (N_26182,N_18091,N_18001);
or U26183 (N_26183,N_18970,N_21816);
nor U26184 (N_26184,N_20647,N_23459);
and U26185 (N_26185,N_23694,N_21274);
or U26186 (N_26186,N_21742,N_20172);
nand U26187 (N_26187,N_23563,N_19386);
xnor U26188 (N_26188,N_19936,N_23059);
and U26189 (N_26189,N_19927,N_18575);
nor U26190 (N_26190,N_22114,N_22249);
or U26191 (N_26191,N_21306,N_19865);
nor U26192 (N_26192,N_19758,N_23319);
or U26193 (N_26193,N_20999,N_19622);
or U26194 (N_26194,N_22646,N_20651);
nor U26195 (N_26195,N_20360,N_20106);
nand U26196 (N_26196,N_19111,N_22678);
nor U26197 (N_26197,N_18231,N_23775);
nand U26198 (N_26198,N_23511,N_20258);
nand U26199 (N_26199,N_21432,N_18352);
nor U26200 (N_26200,N_22314,N_23629);
and U26201 (N_26201,N_21813,N_18959);
and U26202 (N_26202,N_19090,N_21558);
or U26203 (N_26203,N_20628,N_18413);
or U26204 (N_26204,N_22634,N_22253);
nor U26205 (N_26205,N_23225,N_18899);
and U26206 (N_26206,N_18546,N_21960);
nor U26207 (N_26207,N_23471,N_21223);
and U26208 (N_26208,N_21456,N_18579);
xnor U26209 (N_26209,N_21746,N_18382);
nand U26210 (N_26210,N_20802,N_21399);
xor U26211 (N_26211,N_21020,N_22072);
and U26212 (N_26212,N_22152,N_22619);
and U26213 (N_26213,N_22356,N_21271);
nand U26214 (N_26214,N_20416,N_18754);
nand U26215 (N_26215,N_20779,N_18765);
xnor U26216 (N_26216,N_21109,N_19890);
and U26217 (N_26217,N_21534,N_18189);
nor U26218 (N_26218,N_23614,N_22623);
nor U26219 (N_26219,N_19394,N_22801);
xnor U26220 (N_26220,N_20993,N_20137);
and U26221 (N_26221,N_18711,N_21154);
or U26222 (N_26222,N_21651,N_23061);
or U26223 (N_26223,N_23967,N_23281);
or U26224 (N_26224,N_20192,N_19182);
nor U26225 (N_26225,N_22839,N_23610);
and U26226 (N_26226,N_20268,N_19245);
or U26227 (N_26227,N_20640,N_23293);
nand U26228 (N_26228,N_19021,N_20830);
and U26229 (N_26229,N_21218,N_23687);
xor U26230 (N_26230,N_21701,N_22832);
nor U26231 (N_26231,N_23665,N_23211);
and U26232 (N_26232,N_23344,N_23969);
nor U26233 (N_26233,N_23236,N_22685);
nor U26234 (N_26234,N_21904,N_18622);
and U26235 (N_26235,N_18623,N_23832);
xor U26236 (N_26236,N_19639,N_20359);
and U26237 (N_26237,N_18842,N_22636);
nor U26238 (N_26238,N_18077,N_18931);
xnor U26239 (N_26239,N_19768,N_23433);
nand U26240 (N_26240,N_23534,N_22318);
and U26241 (N_26241,N_22004,N_19575);
or U26242 (N_26242,N_18458,N_22596);
and U26243 (N_26243,N_19349,N_20352);
nand U26244 (N_26244,N_20909,N_19798);
nor U26245 (N_26245,N_21928,N_23399);
nor U26246 (N_26246,N_21689,N_21003);
nor U26247 (N_26247,N_20450,N_21215);
xnor U26248 (N_26248,N_21268,N_22846);
or U26249 (N_26249,N_18818,N_20801);
nand U26250 (N_26250,N_19720,N_21008);
or U26251 (N_26251,N_23278,N_18938);
nor U26252 (N_26252,N_18133,N_21323);
xor U26253 (N_26253,N_21041,N_21317);
or U26254 (N_26254,N_22120,N_22758);
nand U26255 (N_26255,N_20446,N_21184);
or U26256 (N_26256,N_18093,N_23432);
nand U26257 (N_26257,N_20627,N_19899);
xor U26258 (N_26258,N_23142,N_22478);
xnor U26259 (N_26259,N_23336,N_20383);
or U26260 (N_26260,N_21367,N_22908);
or U26261 (N_26261,N_19375,N_18062);
or U26262 (N_26262,N_19352,N_20065);
nand U26263 (N_26263,N_19498,N_19261);
and U26264 (N_26264,N_18438,N_21454);
or U26265 (N_26265,N_22077,N_20320);
xor U26266 (N_26266,N_21994,N_20037);
xor U26267 (N_26267,N_20314,N_21196);
xor U26268 (N_26268,N_23609,N_20090);
nor U26269 (N_26269,N_19537,N_23931);
nand U26270 (N_26270,N_21912,N_21321);
and U26271 (N_26271,N_20708,N_22054);
nand U26272 (N_26272,N_19163,N_23896);
xor U26273 (N_26273,N_21084,N_18704);
nand U26274 (N_26274,N_23998,N_18495);
nor U26275 (N_26275,N_23097,N_18202);
xnor U26276 (N_26276,N_22269,N_22736);
nor U26277 (N_26277,N_19125,N_18033);
nand U26278 (N_26278,N_20831,N_20006);
and U26279 (N_26279,N_23182,N_21586);
nand U26280 (N_26280,N_20758,N_23936);
nand U26281 (N_26281,N_19246,N_18092);
nand U26282 (N_26282,N_20251,N_20527);
and U26283 (N_26283,N_18292,N_22430);
nor U26284 (N_26284,N_18253,N_19112);
xnor U26285 (N_26285,N_20480,N_19703);
and U26286 (N_26286,N_23848,N_19851);
nand U26287 (N_26287,N_21334,N_21112);
and U26288 (N_26288,N_19596,N_20880);
xor U26289 (N_26289,N_23363,N_23378);
nor U26290 (N_26290,N_19581,N_19519);
or U26291 (N_26291,N_18615,N_22716);
nand U26292 (N_26292,N_21066,N_22143);
and U26293 (N_26293,N_20580,N_23210);
nor U26294 (N_26294,N_22990,N_20027);
nor U26295 (N_26295,N_21022,N_19869);
nand U26296 (N_26296,N_20510,N_21695);
xor U26297 (N_26297,N_22782,N_22357);
and U26298 (N_26298,N_19052,N_18777);
and U26299 (N_26299,N_23035,N_19765);
nor U26300 (N_26300,N_23443,N_21600);
nand U26301 (N_26301,N_20181,N_20490);
xnor U26302 (N_26302,N_23313,N_22091);
xor U26303 (N_26303,N_19128,N_21790);
and U26304 (N_26304,N_23797,N_21827);
nand U26305 (N_26305,N_19287,N_22573);
xnor U26306 (N_26306,N_20405,N_22897);
or U26307 (N_26307,N_19544,N_19249);
nor U26308 (N_26308,N_23438,N_20598);
xor U26309 (N_26309,N_22833,N_18234);
and U26310 (N_26310,N_22658,N_20475);
or U26311 (N_26311,N_23231,N_22992);
nand U26312 (N_26312,N_22061,N_21832);
nand U26313 (N_26313,N_22662,N_23664);
and U26314 (N_26314,N_18860,N_22995);
xnor U26315 (N_26315,N_18820,N_18625);
xor U26316 (N_26316,N_19377,N_22341);
and U26317 (N_26317,N_19977,N_22799);
xor U26318 (N_26318,N_20572,N_22786);
nor U26319 (N_26319,N_23384,N_18021);
nand U26320 (N_26320,N_22524,N_22383);
nor U26321 (N_26321,N_22074,N_23175);
nor U26322 (N_26322,N_19472,N_21810);
or U26323 (N_26323,N_18229,N_22012);
xor U26324 (N_26324,N_21465,N_18102);
xor U26325 (N_26325,N_18529,N_19664);
nor U26326 (N_26326,N_22645,N_23040);
nor U26327 (N_26327,N_19886,N_19895);
nor U26328 (N_26328,N_20270,N_22794);
nor U26329 (N_26329,N_22640,N_20344);
or U26330 (N_26330,N_23138,N_23670);
or U26331 (N_26331,N_21416,N_18894);
or U26332 (N_26332,N_19492,N_23958);
or U26333 (N_26333,N_23203,N_18553);
nor U26334 (N_26334,N_20894,N_18067);
and U26335 (N_26335,N_20530,N_21884);
xnor U26336 (N_26336,N_22160,N_20316);
xor U26337 (N_26337,N_21325,N_18617);
nor U26338 (N_26338,N_19919,N_22090);
xnor U26339 (N_26339,N_21750,N_18542);
or U26340 (N_26340,N_20240,N_21908);
nand U26341 (N_26341,N_23994,N_20965);
xor U26342 (N_26342,N_21853,N_19268);
nand U26343 (N_26343,N_20421,N_21116);
and U26344 (N_26344,N_20836,N_22547);
or U26345 (N_26345,N_21997,N_23648);
or U26346 (N_26346,N_21450,N_19409);
nor U26347 (N_26347,N_23636,N_18309);
nor U26348 (N_26348,N_19183,N_18505);
or U26349 (N_26349,N_20859,N_22476);
nand U26350 (N_26350,N_22439,N_20789);
nor U26351 (N_26351,N_19578,N_20855);
xor U26352 (N_26352,N_23220,N_20230);
and U26353 (N_26353,N_20973,N_23131);
nor U26354 (N_26354,N_20878,N_21155);
or U26355 (N_26355,N_18871,N_23112);
or U26356 (N_26356,N_21208,N_23430);
and U26357 (N_26357,N_20325,N_20179);
xor U26358 (N_26358,N_21180,N_18090);
nor U26359 (N_26359,N_19473,N_19216);
and U26360 (N_26360,N_23926,N_23677);
or U26361 (N_26361,N_19426,N_19335);
xor U26362 (N_26362,N_23311,N_22913);
xor U26363 (N_26363,N_23342,N_21349);
xnor U26364 (N_26364,N_22060,N_20930);
xor U26365 (N_26365,N_19935,N_22496);
nor U26366 (N_26366,N_21848,N_20030);
nor U26367 (N_26367,N_20158,N_20639);
xor U26368 (N_26368,N_19522,N_21656);
and U26369 (N_26369,N_23566,N_22666);
or U26370 (N_26370,N_19340,N_18342);
and U26371 (N_26371,N_18023,N_22750);
or U26372 (N_26372,N_20525,N_21587);
nand U26373 (N_26373,N_23685,N_21319);
xnor U26374 (N_26374,N_19025,N_18784);
xnor U26375 (N_26375,N_19407,N_19479);
nor U26376 (N_26376,N_22262,N_22125);
nor U26377 (N_26377,N_22070,N_23845);
nor U26378 (N_26378,N_22656,N_18235);
xor U26379 (N_26379,N_21930,N_18631);
or U26380 (N_26380,N_21314,N_23655);
nor U26381 (N_26381,N_21915,N_19306);
nand U26382 (N_26382,N_22550,N_18159);
or U26383 (N_26383,N_18994,N_19868);
nand U26384 (N_26384,N_18854,N_19495);
and U26385 (N_26385,N_19373,N_20242);
xnor U26386 (N_26386,N_18752,N_22058);
nand U26387 (N_26387,N_23916,N_23055);
or U26388 (N_26388,N_22335,N_22557);
nor U26389 (N_26389,N_18695,N_20828);
nand U26390 (N_26390,N_21745,N_22161);
xor U26391 (N_26391,N_19471,N_21010);
and U26392 (N_26392,N_18915,N_18441);
or U26393 (N_26393,N_18389,N_21420);
nand U26394 (N_26394,N_20409,N_21108);
and U26395 (N_26395,N_18605,N_20199);
and U26396 (N_26396,N_21650,N_22082);
nand U26397 (N_26397,N_20767,N_19145);
xor U26398 (N_26398,N_20187,N_22841);
nand U26399 (N_26399,N_19548,N_23197);
nand U26400 (N_26400,N_22308,N_18888);
nand U26401 (N_26401,N_18385,N_22363);
nand U26402 (N_26402,N_20358,N_20346);
or U26403 (N_26403,N_20614,N_21179);
and U26404 (N_26404,N_22701,N_21721);
or U26405 (N_26405,N_22512,N_20942);
or U26406 (N_26406,N_22525,N_20742);
nor U26407 (N_26407,N_21168,N_18914);
or U26408 (N_26408,N_19134,N_20449);
nand U26409 (N_26409,N_22627,N_19325);
nand U26410 (N_26410,N_18678,N_18578);
nor U26411 (N_26411,N_19820,N_23635);
xor U26412 (N_26412,N_19160,N_18736);
xnor U26413 (N_26413,N_22747,N_21205);
and U26414 (N_26414,N_19929,N_23767);
xnor U26415 (N_26415,N_19949,N_22250);
or U26416 (N_26416,N_22400,N_23623);
and U26417 (N_26417,N_23073,N_23833);
or U26418 (N_26418,N_22454,N_18165);
and U26419 (N_26419,N_23316,N_19697);
xnor U26420 (N_26420,N_20167,N_19941);
xnor U26421 (N_26421,N_23569,N_19221);
or U26422 (N_26422,N_23167,N_21846);
or U26423 (N_26423,N_21019,N_19226);
nand U26424 (N_26424,N_18853,N_19509);
and U26425 (N_26425,N_18443,N_22960);
and U26426 (N_26426,N_21237,N_22933);
and U26427 (N_26427,N_22586,N_21229);
and U26428 (N_26428,N_19700,N_22987);
xnor U26429 (N_26429,N_23528,N_18239);
nand U26430 (N_26430,N_19276,N_18191);
nor U26431 (N_26431,N_22719,N_20393);
nand U26432 (N_26432,N_21903,N_22157);
xnor U26433 (N_26433,N_19058,N_20057);
or U26434 (N_26434,N_23080,N_22905);
nand U26435 (N_26435,N_18948,N_18769);
xor U26436 (N_26436,N_23009,N_18082);
nor U26437 (N_26437,N_21255,N_20301);
or U26438 (N_26438,N_22643,N_18434);
nor U26439 (N_26439,N_20285,N_19028);
or U26440 (N_26440,N_18040,N_23223);
and U26441 (N_26441,N_20595,N_22281);
and U26442 (N_26442,N_19076,N_18599);
nand U26443 (N_26443,N_22489,N_18347);
nor U26444 (N_26444,N_18999,N_19347);
nor U26445 (N_26445,N_19136,N_22600);
nor U26446 (N_26446,N_19980,N_18449);
nand U26447 (N_26447,N_18273,N_18362);
xnor U26448 (N_26448,N_18884,N_18120);
xor U26449 (N_26449,N_21542,N_21546);
or U26450 (N_26450,N_23519,N_20059);
xor U26451 (N_26451,N_19235,N_23093);
and U26452 (N_26452,N_23162,N_18668);
or U26453 (N_26453,N_22178,N_18523);
or U26454 (N_26454,N_23287,N_21559);
and U26455 (N_26455,N_20364,N_19872);
xnor U26456 (N_26456,N_18666,N_23717);
nor U26457 (N_26457,N_21913,N_20294);
nor U26458 (N_26458,N_22078,N_20469);
xor U26459 (N_26459,N_22186,N_19292);
and U26460 (N_26460,N_23164,N_23711);
nand U26461 (N_26461,N_22821,N_22593);
and U26462 (N_26462,N_22007,N_23744);
and U26463 (N_26463,N_20620,N_19420);
or U26464 (N_26464,N_21186,N_19594);
and U26465 (N_26465,N_18571,N_20503);
nor U26466 (N_26466,N_19468,N_18486);
nor U26467 (N_26467,N_19669,N_23101);
nor U26468 (N_26468,N_23887,N_22119);
and U26469 (N_26469,N_18920,N_21447);
and U26470 (N_26470,N_18108,N_18464);
nand U26471 (N_26471,N_23042,N_21697);
xor U26472 (N_26472,N_20085,N_18514);
xnor U26473 (N_26473,N_22958,N_22994);
nor U26474 (N_26474,N_22085,N_18425);
nand U26475 (N_26475,N_19333,N_23265);
nand U26476 (N_26476,N_19726,N_20350);
nand U26477 (N_26477,N_19787,N_21410);
nor U26478 (N_26478,N_18834,N_18758);
or U26479 (N_26479,N_20962,N_21072);
nor U26480 (N_26480,N_20356,N_22936);
nand U26481 (N_26481,N_22491,N_22381);
and U26482 (N_26482,N_22456,N_23486);
xnor U26483 (N_26483,N_21476,N_21993);
nor U26484 (N_26484,N_21148,N_20650);
nor U26485 (N_26485,N_21320,N_19200);
and U26486 (N_26486,N_19143,N_21974);
nor U26487 (N_26487,N_20753,N_19835);
and U26488 (N_26488,N_18437,N_23400);
nand U26489 (N_26489,N_23440,N_21584);
and U26490 (N_26490,N_20883,N_21807);
xor U26491 (N_26491,N_21487,N_23347);
nor U26492 (N_26492,N_20147,N_19368);
nor U26493 (N_26493,N_22961,N_21503);
and U26494 (N_26494,N_18494,N_19290);
xnor U26495 (N_26495,N_21359,N_19142);
and U26496 (N_26496,N_21344,N_19167);
nor U26497 (N_26497,N_21906,N_18314);
xnor U26498 (N_26498,N_20439,N_22172);
and U26499 (N_26499,N_22660,N_18705);
or U26500 (N_26500,N_18766,N_21139);
xnor U26501 (N_26501,N_20848,N_20824);
nand U26502 (N_26502,N_21596,N_23508);
and U26503 (N_26503,N_19746,N_22805);
and U26504 (N_26504,N_19625,N_19433);
xor U26505 (N_26505,N_18500,N_18675);
and U26506 (N_26506,N_20005,N_18319);
xnor U26507 (N_26507,N_22311,N_20877);
xnor U26508 (N_26508,N_21602,N_22970);
or U26509 (N_26509,N_23861,N_19301);
nor U26510 (N_26510,N_19825,N_20532);
nand U26511 (N_26511,N_23940,N_23464);
or U26512 (N_26512,N_20630,N_19077);
nor U26513 (N_26513,N_18768,N_22469);
nor U26514 (N_26514,N_21409,N_20262);
nor U26515 (N_26515,N_20849,N_18455);
or U26516 (N_26516,N_22523,N_19993);
xnor U26517 (N_26517,N_18534,N_18781);
xor U26518 (N_26518,N_22735,N_23827);
or U26519 (N_26519,N_20341,N_21151);
or U26520 (N_26520,N_22981,N_20437);
or U26521 (N_26521,N_21667,N_18215);
xor U26522 (N_26522,N_21159,N_18294);
and U26523 (N_26523,N_20124,N_20571);
nor U26524 (N_26524,N_19856,N_18964);
nor U26525 (N_26525,N_20487,N_22706);
and U26526 (N_26526,N_20384,N_20422);
nand U26527 (N_26527,N_19840,N_20456);
nor U26528 (N_26528,N_19006,N_22813);
or U26529 (N_26529,N_19958,N_20724);
xnor U26530 (N_26530,N_23497,N_22959);
and U26531 (N_26531,N_20105,N_23134);
nand U26532 (N_26532,N_19501,N_21749);
xor U26533 (N_26533,N_18606,N_21979);
xor U26534 (N_26534,N_23663,N_19766);
xnor U26535 (N_26535,N_19075,N_21687);
xnor U26536 (N_26536,N_19779,N_19329);
nand U26537 (N_26537,N_21850,N_21840);
xnor U26538 (N_26538,N_20140,N_22703);
xnor U26539 (N_26539,N_20044,N_22415);
and U26540 (N_26540,N_18796,N_22251);
and U26541 (N_26541,N_20757,N_21889);
xnor U26542 (N_26542,N_22237,N_22310);
or U26543 (N_26543,N_23525,N_23638);
xor U26544 (N_26544,N_18431,N_19909);
xor U26545 (N_26545,N_22305,N_21512);
nand U26546 (N_26546,N_19630,N_22777);
nand U26547 (N_26547,N_21953,N_22601);
nand U26548 (N_26548,N_22221,N_22741);
and U26549 (N_26549,N_18921,N_21955);
and U26550 (N_26550,N_20579,N_23632);
nand U26551 (N_26551,N_22769,N_18183);
or U26552 (N_26552,N_21623,N_23707);
nand U26553 (N_26553,N_19446,N_23444);
nor U26554 (N_26554,N_18628,N_19557);
nand U26555 (N_26555,N_20713,N_18570);
or U26556 (N_26556,N_23276,N_20731);
xnor U26557 (N_26557,N_23539,N_21466);
nand U26558 (N_26558,N_18851,N_20602);
or U26559 (N_26559,N_20441,N_19054);
nand U26560 (N_26560,N_19607,N_18802);
nor U26561 (N_26561,N_22700,N_19045);
nand U26562 (N_26562,N_20624,N_23651);
and U26563 (N_26563,N_20511,N_21737);
or U26564 (N_26564,N_19535,N_23067);
and U26565 (N_26565,N_21615,N_21449);
and U26566 (N_26566,N_20710,N_22605);
and U26567 (N_26567,N_18783,N_23151);
xnor U26568 (N_26568,N_22891,N_20408);
and U26569 (N_26569,N_23230,N_23616);
and U26570 (N_26570,N_20012,N_21297);
or U26571 (N_26571,N_22450,N_21963);
nor U26572 (N_26572,N_21896,N_19844);
or U26573 (N_26573,N_20493,N_23253);
nor U26574 (N_26574,N_19879,N_21213);
and U26575 (N_26575,N_19140,N_21437);
and U26576 (N_26576,N_21860,N_23815);
xor U26577 (N_26577,N_20982,N_23551);
and U26578 (N_26578,N_23466,N_20183);
and U26579 (N_26579,N_20492,N_22180);
nand U26580 (N_26580,N_18046,N_22628);
xor U26581 (N_26581,N_18315,N_23076);
xnor U26582 (N_26582,N_19334,N_22106);
nand U26583 (N_26583,N_18423,N_20186);
nor U26584 (N_26584,N_18481,N_23340);
xor U26585 (N_26585,N_20649,N_21210);
xnor U26586 (N_26586,N_23262,N_23380);
nor U26587 (N_26587,N_19896,N_18406);
or U26588 (N_26588,N_20975,N_21826);
nand U26589 (N_26589,N_19313,N_20956);
and U26590 (N_26590,N_21817,N_20901);
nor U26591 (N_26591,N_20521,N_20175);
nor U26592 (N_26592,N_21727,N_19715);
xor U26593 (N_26593,N_22615,N_21736);
xnor U26594 (N_26594,N_20335,N_20080);
nor U26595 (N_26595,N_22006,N_18026);
nand U26596 (N_26596,N_23853,N_23491);
xnor U26597 (N_26597,N_23445,N_20562);
nand U26598 (N_26598,N_22838,N_18103);
nand U26599 (N_26599,N_23437,N_21348);
nor U26600 (N_26600,N_19430,N_20275);
or U26601 (N_26601,N_22113,N_19164);
or U26602 (N_26602,N_18372,N_22338);
and U26603 (N_26603,N_23158,N_22808);
xnor U26604 (N_26604,N_21822,N_21053);
xor U26605 (N_26605,N_22603,N_19613);
or U26606 (N_26606,N_19284,N_19330);
xor U26607 (N_26607,N_23522,N_20398);
and U26608 (N_26608,N_23927,N_18968);
or U26609 (N_26609,N_21678,N_22604);
and U26610 (N_26610,N_22588,N_21052);
nor U26611 (N_26611,N_18192,N_23049);
nand U26612 (N_26612,N_21573,N_22188);
or U26613 (N_26613,N_21479,N_21781);
and U26614 (N_26614,N_19135,N_23221);
xor U26615 (N_26615,N_18100,N_20787);
xnor U26616 (N_26616,N_23750,N_21595);
or U26617 (N_26617,N_20021,N_19036);
xnor U26618 (N_26618,N_19483,N_23689);
or U26619 (N_26619,N_20177,N_21341);
nand U26620 (N_26620,N_18593,N_20738);
or U26621 (N_26621,N_21644,N_21117);
and U26622 (N_26622,N_22083,N_21015);
nor U26623 (N_26623,N_18044,N_18059);
xor U26624 (N_26624,N_23222,N_22860);
nor U26625 (N_26625,N_21163,N_21978);
xnor U26626 (N_26626,N_18672,N_19467);
and U26627 (N_26627,N_21984,N_20073);
xnor U26628 (N_26628,N_23362,N_19039);
or U26629 (N_26629,N_19445,N_21834);
and U26630 (N_26630,N_19963,N_18950);
nor U26631 (N_26631,N_23774,N_22073);
and U26632 (N_26632,N_21421,N_21766);
and U26633 (N_26633,N_21625,N_18006);
xnor U26634 (N_26634,N_22765,N_19412);
xnor U26635 (N_26635,N_23358,N_23646);
or U26636 (N_26636,N_19930,N_18071);
or U26637 (N_26637,N_18679,N_18010);
nor U26638 (N_26638,N_23521,N_21277);
nor U26639 (N_26639,N_19793,N_20370);
nand U26640 (N_26640,N_22098,N_18152);
nor U26641 (N_26641,N_18690,N_20361);
and U26642 (N_26642,N_19018,N_20061);
nor U26643 (N_26643,N_23268,N_18902);
nand U26644 (N_26644,N_19811,N_21862);
and U26645 (N_26645,N_18744,N_18200);
or U26646 (N_26646,N_20244,N_20625);
and U26647 (N_26647,N_23377,N_21965);
or U26648 (N_26648,N_23547,N_23427);
nor U26649 (N_26649,N_22694,N_21808);
nand U26650 (N_26650,N_23618,N_20231);
or U26651 (N_26651,N_21547,N_22975);
xnor U26652 (N_26652,N_18084,N_18986);
nor U26653 (N_26653,N_20149,N_21295);
xor U26654 (N_26654,N_19003,N_21722);
xor U26655 (N_26655,N_21545,N_23963);
or U26656 (N_26656,N_19699,N_23764);
nor U26657 (N_26657,N_23989,N_22187);
and U26658 (N_26658,N_20637,N_21370);
xnor U26659 (N_26659,N_19514,N_20032);
nor U26660 (N_26660,N_22664,N_19621);
xor U26661 (N_26661,N_18687,N_20250);
or U26662 (N_26662,N_23168,N_21444);
nor U26663 (N_26663,N_18137,N_23229);
nor U26664 (N_26664,N_18714,N_22204);
or U26665 (N_26665,N_21217,N_22219);
nor U26666 (N_26666,N_19667,N_21267);
and U26667 (N_26667,N_19588,N_19201);
xnor U26668 (N_26668,N_22111,N_21375);
xnor U26669 (N_26669,N_19314,N_19792);
xnor U26670 (N_26670,N_18655,N_23801);
nor U26671 (N_26671,N_20952,N_18142);
nand U26672 (N_26672,N_23011,N_20204);
nor U26673 (N_26673,N_20950,N_23295);
or U26674 (N_26674,N_18808,N_23873);
and U26675 (N_26675,N_18002,N_23706);
nor U26676 (N_26676,N_21471,N_18907);
nor U26677 (N_26677,N_21250,N_23212);
or U26678 (N_26678,N_19632,N_19281);
or U26679 (N_26679,N_23749,N_19893);
nor U26680 (N_26680,N_21131,N_23893);
xor U26681 (N_26681,N_21645,N_18647);
or U26682 (N_26682,N_21355,N_22847);
or U26683 (N_26683,N_22870,N_19871);
or U26684 (N_26684,N_23216,N_21485);
xor U26685 (N_26685,N_22115,N_22176);
nor U26686 (N_26686,N_23490,N_23530);
nand U26687 (N_26687,N_21044,N_19580);
and U26688 (N_26688,N_21728,N_19874);
or U26689 (N_26689,N_23768,N_22810);
or U26690 (N_26690,N_18304,N_21939);
and U26691 (N_26691,N_20146,N_19849);
or U26692 (N_26692,N_19094,N_21961);
or U26693 (N_26693,N_22575,N_23647);
and U26694 (N_26694,N_19322,N_20201);
nor U26695 (N_26695,N_22518,N_19608);
nor U26696 (N_26696,N_19126,N_23125);
xnor U26697 (N_26697,N_23773,N_21442);
and U26698 (N_26698,N_19754,N_22568);
nor U26699 (N_26699,N_23881,N_23626);
nand U26700 (N_26700,N_18698,N_21455);
nand U26701 (N_26701,N_21411,N_21204);
and U26702 (N_26702,N_21106,N_23105);
nand U26703 (N_26703,N_22519,N_23299);
nand U26704 (N_26704,N_19190,N_21245);
or U26705 (N_26705,N_23951,N_18845);
nor U26706 (N_26706,N_20617,N_23867);
xor U26707 (N_26707,N_23979,N_21098);
or U26708 (N_26708,N_19892,N_18407);
nor U26709 (N_26709,N_18973,N_21585);
nor U26710 (N_26710,N_22989,N_22342);
nand U26711 (N_26711,N_19503,N_23734);
or U26712 (N_26712,N_20363,N_18585);
nor U26713 (N_26713,N_21952,N_18827);
nor U26714 (N_26714,N_23909,N_22407);
xnor U26715 (N_26715,N_21762,N_19228);
or U26716 (N_26716,N_22164,N_18722);
xnor U26717 (N_26717,N_18639,N_20267);
and U26718 (N_26718,N_23558,N_18016);
or U26719 (N_26719,N_23031,N_18621);
or U26720 (N_26720,N_21353,N_20283);
and U26721 (N_26721,N_18790,N_21195);
or U26722 (N_26722,N_18318,N_23804);
xor U26723 (N_26723,N_21260,N_18776);
and U26724 (N_26724,N_18028,N_22389);
xnor U26725 (N_26725,N_18473,N_23000);
nand U26726 (N_26726,N_23615,N_22192);
or U26727 (N_26727,N_23123,N_20846);
or U26728 (N_26728,N_18447,N_23755);
nor U26729 (N_26729,N_21257,N_21082);
nand U26730 (N_26730,N_18353,N_21854);
or U26731 (N_26731,N_23137,N_23233);
or U26732 (N_26732,N_18364,N_18334);
nand U26733 (N_26733,N_18045,N_23424);
nor U26734 (N_26734,N_23122,N_23863);
or U26735 (N_26735,N_21877,N_22358);
and U26736 (N_26736,N_23421,N_20928);
and U26737 (N_26737,N_19484,N_18576);
xnor U26738 (N_26738,N_20296,N_19769);
or U26739 (N_26739,N_20661,N_19807);
and U26740 (N_26740,N_23452,N_20099);
nand U26741 (N_26741,N_23352,N_22027);
xor U26742 (N_26742,N_18937,N_19704);
xor U26743 (N_26743,N_23672,N_18054);
nor U26744 (N_26744,N_22964,N_23608);
xor U26745 (N_26745,N_22132,N_20966);
or U26746 (N_26746,N_22432,N_20535);
nand U26747 (N_26747,N_20777,N_22563);
xnor U26748 (N_26748,N_22081,N_22284);
or U26749 (N_26749,N_20419,N_21893);
and U26750 (N_26750,N_19104,N_19716);
or U26751 (N_26751,N_23368,N_21157);
nor U26752 (N_26752,N_22934,N_22131);
nand U26753 (N_26753,N_21513,N_19677);
nand U26754 (N_26754,N_21324,N_21384);
and U26755 (N_26755,N_18761,N_21247);
or U26756 (N_26756,N_21907,N_23722);
nor U26757 (N_26757,N_20264,N_20660);
nor U26758 (N_26758,N_19346,N_23389);
nand U26759 (N_26759,N_23503,N_22756);
nor U26760 (N_26760,N_22441,N_23324);
or U26761 (N_26761,N_22359,N_23057);
and U26762 (N_26762,N_23039,N_21845);
and U26763 (N_26763,N_20737,N_20766);
or U26764 (N_26764,N_19687,N_18507);
nand U26765 (N_26765,N_22712,N_18412);
nor U26766 (N_26766,N_18405,N_22884);
or U26767 (N_26767,N_21973,N_23982);
or U26768 (N_26768,N_20086,N_22332);
or U26769 (N_26769,N_20055,N_18236);
nand U26770 (N_26770,N_23425,N_21804);
xor U26771 (N_26771,N_20775,N_18893);
nand U26772 (N_26772,N_23591,N_22010);
nor U26773 (N_26773,N_22473,N_19280);
nand U26774 (N_26774,N_19536,N_19600);
nor U26775 (N_26775,N_18502,N_20633);
nand U26776 (N_26776,N_19721,N_21096);
nand U26777 (N_26777,N_18732,N_19427);
nor U26778 (N_26778,N_19117,N_23487);
or U26779 (N_26779,N_20019,N_19070);
or U26780 (N_26780,N_23729,N_21510);
and U26781 (N_26781,N_21757,N_22554);
nor U26782 (N_26782,N_22611,N_19015);
xnor U26783 (N_26783,N_23745,N_23317);
or U26784 (N_26784,N_19405,N_20911);
nand U26785 (N_26785,N_20512,N_20349);
and U26786 (N_26786,N_22620,N_22943);
nand U26787 (N_26787,N_18313,N_23637);
and U26788 (N_26788,N_19791,N_19175);
xnor U26789 (N_26789,N_22759,N_22797);
xor U26790 (N_26790,N_22924,N_19401);
or U26791 (N_26791,N_18519,N_22707);
and U26792 (N_26792,N_22037,N_22698);
or U26793 (N_26793,N_20256,N_22875);
nand U26794 (N_26794,N_19722,N_21497);
nor U26795 (N_26795,N_20903,N_22858);
xor U26796 (N_26796,N_23966,N_20096);
and U26797 (N_26797,N_22128,N_20206);
nand U26798 (N_26798,N_18979,N_20860);
or U26799 (N_26799,N_18377,N_22121);
nor U26800 (N_26800,N_22231,N_23721);
or U26801 (N_26801,N_20120,N_22283);
nand U26802 (N_26802,N_22492,N_22956);
and U26803 (N_26803,N_18296,N_21194);
or U26804 (N_26804,N_23999,N_21313);
and U26805 (N_26805,N_19642,N_22714);
xnor U26806 (N_26806,N_22066,N_20263);
nand U26807 (N_26807,N_21207,N_22408);
and U26808 (N_26808,N_23903,N_22999);
xor U26809 (N_26809,N_21261,N_19955);
xor U26810 (N_26810,N_21111,N_20632);
nand U26811 (N_26811,N_19933,N_23329);
and U26812 (N_26812,N_23388,N_19303);
or U26813 (N_26813,N_22239,N_20271);
or U26814 (N_26814,N_19574,N_19208);
or U26815 (N_26815,N_22460,N_20223);
nor U26816 (N_26816,N_18955,N_20116);
xor U26817 (N_26817,N_18862,N_22631);
nor U26818 (N_26818,N_20852,N_21264);
and U26819 (N_26819,N_23402,N_20434);
and U26820 (N_26820,N_20712,N_21606);
nor U26821 (N_26821,N_21404,N_21067);
and U26822 (N_26822,N_21398,N_22695);
nand U26823 (N_26823,N_19120,N_21831);
xnor U26824 (N_26824,N_22033,N_23895);
nor U26825 (N_26825,N_21156,N_22126);
nor U26826 (N_26826,N_21333,N_20885);
or U26827 (N_26827,N_21927,N_18387);
nand U26828 (N_26828,N_19444,N_23312);
xnor U26829 (N_26829,N_19889,N_22345);
or U26830 (N_26830,N_22543,N_18106);
or U26831 (N_26831,N_22418,N_22583);
nor U26832 (N_26832,N_18247,N_23387);
or U26833 (N_26833,N_21738,N_19367);
xor U26834 (N_26834,N_18470,N_19266);
nor U26835 (N_26835,N_23371,N_22717);
or U26836 (N_26836,N_23332,N_18276);
nor U26837 (N_26837,N_20313,N_23780);
or U26838 (N_26838,N_22579,N_19177);
nand U26839 (N_26839,N_18957,N_22349);
nor U26840 (N_26840,N_18065,N_22474);
nor U26841 (N_26841,N_18642,N_18307);
or U26842 (N_26842,N_21371,N_18012);
nor U26843 (N_26843,N_23089,N_19885);
or U26844 (N_26844,N_21414,N_21654);
xnor U26845 (N_26845,N_20211,N_19418);
and U26846 (N_26846,N_18806,N_23643);
or U26847 (N_26847,N_19605,N_23671);
and U26848 (N_26848,N_23620,N_19695);
nand U26849 (N_26849,N_18692,N_20936);
nor U26850 (N_26850,N_19474,N_20876);
or U26851 (N_26851,N_20559,N_22515);
and U26852 (N_26852,N_21292,N_21127);
and U26853 (N_26853,N_18975,N_23595);
and U26854 (N_26854,N_23772,N_18960);
or U26855 (N_26855,N_22484,N_23403);
xnor U26856 (N_26856,N_23310,N_20347);
nor U26857 (N_26857,N_21142,N_23069);
nand U26858 (N_26858,N_19549,N_20539);
and U26859 (N_26859,N_20241,N_23792);
nand U26860 (N_26860,N_19300,N_19979);
nor U26861 (N_26861,N_20026,N_22135);
or U26862 (N_26862,N_23888,N_22130);
or U26863 (N_26863,N_18739,N_21279);
and U26864 (N_26864,N_18648,N_20117);
nand U26865 (N_26865,N_18230,N_21107);
or U26866 (N_26866,N_21636,N_18882);
nor U26867 (N_26867,N_21394,N_18662);
and U26868 (N_26868,N_19727,N_21240);
and U26869 (N_26869,N_22842,N_19771);
nand U26870 (N_26870,N_22141,N_22153);
nor U26871 (N_26871,N_23315,N_20516);
nor U26872 (N_26872,N_18633,N_21191);
and U26873 (N_26873,N_22530,N_22191);
or U26874 (N_26874,N_21462,N_19982);
nand U26875 (N_26875,N_18069,N_23766);
or U26876 (N_26876,N_23147,N_21276);
or U26877 (N_26877,N_22475,N_22556);
or U26878 (N_26878,N_22738,N_23083);
xor U26879 (N_26879,N_18943,N_22513);
nor U26880 (N_26880,N_23408,N_20136);
xnor U26881 (N_26881,N_21692,N_21363);
nand U26882 (N_26882,N_18508,N_22928);
xnor U26883 (N_26883,N_19638,N_22255);
and U26884 (N_26884,N_20088,N_20540);
and U26885 (N_26885,N_19132,N_20015);
nand U26886 (N_26886,N_21657,N_18584);
and U26887 (N_26887,N_23594,N_22009);
xnor U26888 (N_26888,N_20773,N_21980);
nor U26889 (N_26889,N_21870,N_21969);
nor U26890 (N_26890,N_18151,N_18788);
nand U26891 (N_26891,N_19592,N_23968);
and U26892 (N_26892,N_20180,N_23870);
xor U26893 (N_26893,N_18604,N_20906);
and U26894 (N_26894,N_21504,N_22410);
and U26895 (N_26895,N_18801,N_21069);
or U26896 (N_26896,N_21043,N_21985);
nand U26897 (N_26897,N_20050,N_18442);
or U26898 (N_26898,N_19694,N_21647);
xnor U26899 (N_26899,N_22622,N_22001);
xnor U26900 (N_26900,N_23947,N_21236);
or U26901 (N_26901,N_22647,N_20317);
nor U26902 (N_26902,N_22653,N_23855);
or U26903 (N_26903,N_20497,N_20653);
nand U26904 (N_26904,N_21881,N_20626);
nand U26905 (N_26905,N_19343,N_23053);
nand U26906 (N_26906,N_19254,N_23406);
nand U26907 (N_26907,N_18787,N_18670);
and U26908 (N_26908,N_22699,N_21270);
xor U26909 (N_26909,N_18816,N_20070);
nor U26910 (N_26910,N_23821,N_22011);
xor U26911 (N_26911,N_19053,N_22739);
and U26912 (N_26912,N_19595,N_20031);
xor U26913 (N_26913,N_19122,N_22300);
nor U26914 (N_26914,N_21611,N_20153);
and U26915 (N_26915,N_19552,N_21577);
nand U26916 (N_26916,N_23784,N_22200);
nand U26917 (N_26917,N_21023,N_19310);
and U26918 (N_26918,N_22819,N_20558);
nand U26919 (N_26919,N_21474,N_21675);
nand U26920 (N_26920,N_23385,N_18785);
or U26921 (N_26921,N_19756,N_19365);
or U26922 (N_26922,N_23448,N_20698);
nand U26923 (N_26923,N_23877,N_20987);
nor U26924 (N_26924,N_21998,N_22258);
or U26925 (N_26925,N_18536,N_21567);
or U26926 (N_26926,N_21164,N_23356);
xor U26927 (N_26927,N_22585,N_19799);
xnor U26928 (N_26928,N_22560,N_23429);
and U26929 (N_26929,N_22630,N_22016);
and U26930 (N_26930,N_21812,N_20988);
and U26931 (N_26931,N_21018,N_21086);
and U26932 (N_26932,N_22602,N_19383);
or U26933 (N_26933,N_23454,N_20522);
xnor U26934 (N_26934,N_22670,N_22110);
or U26935 (N_26935,N_20613,N_21669);
nand U26936 (N_26936,N_21769,N_21206);
or U26937 (N_26937,N_22392,N_18877);
xnor U26938 (N_26938,N_21089,N_22323);
nor U26939 (N_26939,N_21597,N_18686);
nor U26940 (N_26940,N_21232,N_22757);
nor U26941 (N_26941,N_19384,N_23822);
or U26942 (N_26942,N_19643,N_20233);
and U26943 (N_26943,N_18649,N_20302);
xnor U26944 (N_26944,N_20665,N_21532);
or U26945 (N_26945,N_19152,N_19558);
and U26946 (N_26946,N_22935,N_22502);
and U26947 (N_26947,N_23116,N_18338);
nand U26948 (N_26948,N_18373,N_23805);
nor U26949 (N_26949,N_22893,N_20165);
and U26950 (N_26950,N_18421,N_18682);
nor U26951 (N_26951,N_18919,N_19598);
nand U26952 (N_26952,N_22962,N_23117);
or U26953 (N_26953,N_20679,N_23970);
xor U26954 (N_26954,N_20703,N_20657);
or U26955 (N_26955,N_19485,N_21635);
nor U26956 (N_26956,N_21422,N_18701);
xor U26957 (N_26957,N_20594,N_19797);
nand U26958 (N_26958,N_23537,N_23420);
nor U26959 (N_26959,N_23396,N_18196);
nor U26960 (N_26960,N_22879,N_21823);
xor U26961 (N_26961,N_23884,N_18061);
nor U26962 (N_26962,N_19530,N_22194);
xnor U26963 (N_26963,N_18198,N_18659);
and U26964 (N_26964,N_22482,N_22709);
or U26965 (N_26965,N_23070,N_23984);
xnor U26966 (N_26966,N_22898,N_18863);
or U26967 (N_26967,N_19017,N_23259);
nand U26968 (N_26968,N_19106,N_19834);
nor U26969 (N_26969,N_21303,N_19041);
nand U26970 (N_26970,N_21898,N_21798);
nand U26971 (N_26971,N_23856,N_21068);
and U26972 (N_26972,N_18965,N_18408);
xor U26973 (N_26973,N_22896,N_22177);
or U26974 (N_26974,N_22882,N_23275);
xor U26975 (N_26975,N_21283,N_20664);
nor U26976 (N_26976,N_23546,N_22770);
nand U26977 (N_26977,N_20924,N_18459);
nand U26978 (N_26978,N_18728,N_18079);
or U26979 (N_26979,N_21244,N_23269);
and U26980 (N_26980,N_20663,N_21791);
nor U26981 (N_26981,N_23107,N_19767);
or U26982 (N_26982,N_20972,N_22532);
nor U26983 (N_26983,N_20078,N_20749);
nand U26984 (N_26984,N_18221,N_21076);
nand U26985 (N_26985,N_22724,N_22595);
nand U26986 (N_26986,N_22768,N_23279);
and U26987 (N_26987,N_23826,N_23483);
nand U26988 (N_26988,N_23939,N_21290);
nor U26989 (N_26989,N_19645,N_22767);
or U26990 (N_26990,N_23515,N_19341);
nor U26991 (N_26991,N_23562,N_23778);
and U26992 (N_26992,N_22889,N_23449);
xnor U26993 (N_26993,N_23639,N_18742);
xnor U26994 (N_26994,N_18420,N_18070);
nand U26995 (N_26995,N_22571,N_19049);
and U26996 (N_26996,N_21070,N_20835);
and U26997 (N_26997,N_19566,N_18829);
nand U26998 (N_26998,N_23834,N_21658);
or U26999 (N_26999,N_21124,N_20686);
nand U27000 (N_27000,N_19968,N_22686);
nor U27001 (N_27001,N_20794,N_22657);
and U27002 (N_27002,N_21131,N_18594);
nor U27003 (N_27003,N_19560,N_20493);
xnor U27004 (N_27004,N_19566,N_18552);
nor U27005 (N_27005,N_20089,N_21343);
nor U27006 (N_27006,N_19616,N_23919);
xnor U27007 (N_27007,N_23564,N_19058);
and U27008 (N_27008,N_20285,N_22009);
nor U27009 (N_27009,N_23775,N_22261);
xnor U27010 (N_27010,N_19781,N_22154);
or U27011 (N_27011,N_18302,N_18660);
xnor U27012 (N_27012,N_22855,N_22172);
nor U27013 (N_27013,N_18884,N_20729);
or U27014 (N_27014,N_22557,N_20116);
or U27015 (N_27015,N_23033,N_19380);
or U27016 (N_27016,N_20241,N_21305);
xnor U27017 (N_27017,N_21987,N_19763);
or U27018 (N_27018,N_20445,N_19864);
or U27019 (N_27019,N_22926,N_19122);
nand U27020 (N_27020,N_18075,N_19642);
nor U27021 (N_27021,N_22015,N_22126);
or U27022 (N_27022,N_22743,N_20163);
and U27023 (N_27023,N_23638,N_20019);
nand U27024 (N_27024,N_22477,N_20293);
and U27025 (N_27025,N_21553,N_18334);
and U27026 (N_27026,N_21535,N_20944);
and U27027 (N_27027,N_18105,N_22444);
xnor U27028 (N_27028,N_23913,N_22716);
or U27029 (N_27029,N_18191,N_22863);
nand U27030 (N_27030,N_20404,N_21262);
or U27031 (N_27031,N_23966,N_18418);
xor U27032 (N_27032,N_23689,N_20807);
nand U27033 (N_27033,N_20603,N_21702);
and U27034 (N_27034,N_20612,N_18209);
xnor U27035 (N_27035,N_18590,N_23142);
and U27036 (N_27036,N_22391,N_20782);
nand U27037 (N_27037,N_19789,N_18726);
xnor U27038 (N_27038,N_20325,N_20185);
or U27039 (N_27039,N_23720,N_23463);
or U27040 (N_27040,N_18078,N_23255);
nor U27041 (N_27041,N_20784,N_19876);
nor U27042 (N_27042,N_21895,N_22885);
xnor U27043 (N_27043,N_22467,N_23848);
nor U27044 (N_27044,N_20587,N_19600);
nand U27045 (N_27045,N_18753,N_19032);
or U27046 (N_27046,N_22102,N_21277);
nand U27047 (N_27047,N_23994,N_18139);
and U27048 (N_27048,N_19048,N_18525);
or U27049 (N_27049,N_20128,N_18916);
nand U27050 (N_27050,N_19803,N_22887);
or U27051 (N_27051,N_23308,N_19568);
nand U27052 (N_27052,N_23505,N_19138);
nor U27053 (N_27053,N_22832,N_22468);
xnor U27054 (N_27054,N_23699,N_22002);
or U27055 (N_27055,N_18342,N_23248);
nor U27056 (N_27056,N_23734,N_22009);
nand U27057 (N_27057,N_22030,N_21071);
or U27058 (N_27058,N_19534,N_21118);
xnor U27059 (N_27059,N_20470,N_23502);
nor U27060 (N_27060,N_23662,N_19759);
nand U27061 (N_27061,N_23714,N_19150);
xor U27062 (N_27062,N_21493,N_18483);
nor U27063 (N_27063,N_23971,N_18493);
nor U27064 (N_27064,N_19416,N_23367);
nand U27065 (N_27065,N_22593,N_22228);
and U27066 (N_27066,N_18686,N_18356);
nand U27067 (N_27067,N_18419,N_20608);
nand U27068 (N_27068,N_23037,N_22981);
nand U27069 (N_27069,N_21538,N_23810);
and U27070 (N_27070,N_21074,N_21960);
and U27071 (N_27071,N_22828,N_19093);
nor U27072 (N_27072,N_21363,N_19155);
nor U27073 (N_27073,N_18957,N_20520);
nor U27074 (N_27074,N_18608,N_21732);
or U27075 (N_27075,N_20598,N_22493);
xnor U27076 (N_27076,N_21580,N_21034);
xnor U27077 (N_27077,N_21828,N_20708);
nand U27078 (N_27078,N_21489,N_20219);
xor U27079 (N_27079,N_21518,N_23917);
and U27080 (N_27080,N_18806,N_19694);
xor U27081 (N_27081,N_22648,N_19707);
nand U27082 (N_27082,N_18816,N_19472);
xnor U27083 (N_27083,N_22291,N_20193);
or U27084 (N_27084,N_23789,N_23588);
and U27085 (N_27085,N_20255,N_21823);
nand U27086 (N_27086,N_23768,N_20576);
or U27087 (N_27087,N_22278,N_21868);
nor U27088 (N_27088,N_18173,N_22249);
nand U27089 (N_27089,N_22636,N_19460);
nor U27090 (N_27090,N_19135,N_21823);
xor U27091 (N_27091,N_23679,N_19122);
nand U27092 (N_27092,N_20835,N_21951);
nand U27093 (N_27093,N_21429,N_21386);
nand U27094 (N_27094,N_19735,N_22595);
xor U27095 (N_27095,N_18544,N_23958);
nor U27096 (N_27096,N_23701,N_20852);
and U27097 (N_27097,N_18013,N_22289);
xnor U27098 (N_27098,N_22096,N_22648);
nand U27099 (N_27099,N_19659,N_18868);
nand U27100 (N_27100,N_21324,N_18086);
nand U27101 (N_27101,N_23246,N_18508);
and U27102 (N_27102,N_21055,N_22522);
xnor U27103 (N_27103,N_22239,N_23113);
xnor U27104 (N_27104,N_21161,N_18340);
nand U27105 (N_27105,N_19292,N_19946);
xor U27106 (N_27106,N_21435,N_21969);
nand U27107 (N_27107,N_22618,N_19831);
and U27108 (N_27108,N_21869,N_18667);
xnor U27109 (N_27109,N_19936,N_20351);
nor U27110 (N_27110,N_23370,N_22849);
nor U27111 (N_27111,N_20303,N_23381);
nand U27112 (N_27112,N_18724,N_20352);
and U27113 (N_27113,N_18032,N_23953);
or U27114 (N_27114,N_18073,N_19286);
or U27115 (N_27115,N_20518,N_21429);
xnor U27116 (N_27116,N_20801,N_23663);
nor U27117 (N_27117,N_21080,N_20946);
and U27118 (N_27118,N_20798,N_19495);
xor U27119 (N_27119,N_18187,N_23420);
or U27120 (N_27120,N_18419,N_18652);
and U27121 (N_27121,N_22426,N_18809);
nor U27122 (N_27122,N_18424,N_18362);
nand U27123 (N_27123,N_18639,N_22057);
and U27124 (N_27124,N_23911,N_19370);
and U27125 (N_27125,N_21834,N_18321);
nor U27126 (N_27126,N_23527,N_22241);
and U27127 (N_27127,N_22102,N_18714);
xor U27128 (N_27128,N_22745,N_21057);
and U27129 (N_27129,N_22880,N_23208);
xnor U27130 (N_27130,N_21244,N_23226);
or U27131 (N_27131,N_18508,N_19173);
nor U27132 (N_27132,N_21048,N_22186);
and U27133 (N_27133,N_20232,N_22086);
nand U27134 (N_27134,N_18275,N_21593);
or U27135 (N_27135,N_23593,N_22904);
nor U27136 (N_27136,N_21057,N_22787);
xor U27137 (N_27137,N_22539,N_23144);
and U27138 (N_27138,N_20525,N_20252);
nor U27139 (N_27139,N_22619,N_21794);
nor U27140 (N_27140,N_20282,N_19838);
nor U27141 (N_27141,N_22502,N_19753);
nand U27142 (N_27142,N_19732,N_19828);
xor U27143 (N_27143,N_22795,N_19146);
or U27144 (N_27144,N_23718,N_20045);
nand U27145 (N_27145,N_22729,N_23237);
and U27146 (N_27146,N_21174,N_21265);
xnor U27147 (N_27147,N_22964,N_22227);
nor U27148 (N_27148,N_20634,N_18791);
and U27149 (N_27149,N_23911,N_21740);
or U27150 (N_27150,N_19076,N_23622);
or U27151 (N_27151,N_21750,N_23471);
nand U27152 (N_27152,N_20228,N_21725);
or U27153 (N_27153,N_21364,N_21983);
nor U27154 (N_27154,N_21054,N_21118);
or U27155 (N_27155,N_18674,N_22811);
xor U27156 (N_27156,N_19746,N_21812);
and U27157 (N_27157,N_23498,N_20841);
nand U27158 (N_27158,N_19023,N_21222);
nor U27159 (N_27159,N_18809,N_22867);
nor U27160 (N_27160,N_19074,N_18085);
xnor U27161 (N_27161,N_19180,N_18693);
nor U27162 (N_27162,N_22466,N_22695);
or U27163 (N_27163,N_21908,N_21437);
or U27164 (N_27164,N_22543,N_22362);
nand U27165 (N_27165,N_19907,N_19839);
and U27166 (N_27166,N_19585,N_22568);
and U27167 (N_27167,N_20786,N_20386);
xor U27168 (N_27168,N_18788,N_20234);
nor U27169 (N_27169,N_22299,N_23972);
nand U27170 (N_27170,N_20564,N_18322);
nand U27171 (N_27171,N_23536,N_23328);
and U27172 (N_27172,N_19299,N_22697);
or U27173 (N_27173,N_21459,N_20387);
nand U27174 (N_27174,N_18875,N_23128);
xor U27175 (N_27175,N_18807,N_19162);
and U27176 (N_27176,N_19801,N_19381);
or U27177 (N_27177,N_18628,N_21713);
nand U27178 (N_27178,N_18766,N_22961);
xnor U27179 (N_27179,N_18868,N_20957);
nor U27180 (N_27180,N_22551,N_22249);
nand U27181 (N_27181,N_20312,N_23976);
or U27182 (N_27182,N_22616,N_19002);
nor U27183 (N_27183,N_19340,N_20866);
nor U27184 (N_27184,N_19777,N_19637);
nor U27185 (N_27185,N_19566,N_19392);
nor U27186 (N_27186,N_18396,N_23445);
xnor U27187 (N_27187,N_20079,N_20369);
and U27188 (N_27188,N_18077,N_20702);
nor U27189 (N_27189,N_23333,N_19554);
and U27190 (N_27190,N_23030,N_20919);
xor U27191 (N_27191,N_21121,N_22471);
and U27192 (N_27192,N_22884,N_23433);
nor U27193 (N_27193,N_23191,N_19701);
xor U27194 (N_27194,N_22026,N_21941);
and U27195 (N_27195,N_23893,N_19707);
or U27196 (N_27196,N_22868,N_18117);
or U27197 (N_27197,N_18141,N_23185);
nand U27198 (N_27198,N_18431,N_20211);
nand U27199 (N_27199,N_18479,N_21603);
xor U27200 (N_27200,N_23306,N_20351);
nor U27201 (N_27201,N_18111,N_22266);
nor U27202 (N_27202,N_21775,N_23403);
or U27203 (N_27203,N_18036,N_21907);
nor U27204 (N_27204,N_23588,N_21874);
nor U27205 (N_27205,N_21788,N_21680);
xnor U27206 (N_27206,N_23833,N_20202);
nand U27207 (N_27207,N_23545,N_18015);
nand U27208 (N_27208,N_21226,N_21191);
xor U27209 (N_27209,N_20556,N_19416);
nor U27210 (N_27210,N_21584,N_18142);
nand U27211 (N_27211,N_21685,N_19182);
xnor U27212 (N_27212,N_21198,N_20065);
nor U27213 (N_27213,N_21926,N_22063);
and U27214 (N_27214,N_19413,N_20289);
nor U27215 (N_27215,N_20136,N_21359);
and U27216 (N_27216,N_19798,N_20990);
and U27217 (N_27217,N_21706,N_19848);
or U27218 (N_27218,N_22423,N_22812);
xor U27219 (N_27219,N_18517,N_22443);
or U27220 (N_27220,N_22018,N_21286);
nor U27221 (N_27221,N_21392,N_19382);
nor U27222 (N_27222,N_22247,N_20263);
or U27223 (N_27223,N_22505,N_20121);
nand U27224 (N_27224,N_23266,N_19800);
nor U27225 (N_27225,N_18349,N_21710);
or U27226 (N_27226,N_23850,N_22454);
nor U27227 (N_27227,N_18991,N_20139);
or U27228 (N_27228,N_18363,N_18998);
xor U27229 (N_27229,N_23799,N_21353);
or U27230 (N_27230,N_18546,N_22023);
and U27231 (N_27231,N_22422,N_21584);
nor U27232 (N_27232,N_18087,N_20310);
or U27233 (N_27233,N_21879,N_19981);
xor U27234 (N_27234,N_19377,N_19893);
and U27235 (N_27235,N_21595,N_22997);
nand U27236 (N_27236,N_21864,N_22499);
xnor U27237 (N_27237,N_19498,N_23257);
nor U27238 (N_27238,N_19977,N_21909);
xor U27239 (N_27239,N_22793,N_21005);
nor U27240 (N_27240,N_23541,N_21089);
nand U27241 (N_27241,N_23253,N_22576);
nand U27242 (N_27242,N_19460,N_20995);
xnor U27243 (N_27243,N_19652,N_19649);
nand U27244 (N_27244,N_19666,N_18577);
or U27245 (N_27245,N_19069,N_18563);
xnor U27246 (N_27246,N_20426,N_18743);
or U27247 (N_27247,N_20844,N_23933);
and U27248 (N_27248,N_18851,N_18455);
xor U27249 (N_27249,N_22588,N_21286);
xor U27250 (N_27250,N_22317,N_19226);
nor U27251 (N_27251,N_19396,N_19234);
or U27252 (N_27252,N_22740,N_21374);
nand U27253 (N_27253,N_19978,N_18004);
nor U27254 (N_27254,N_21213,N_21099);
xnor U27255 (N_27255,N_21789,N_20519);
nand U27256 (N_27256,N_20145,N_21767);
and U27257 (N_27257,N_23053,N_21764);
nor U27258 (N_27258,N_22653,N_21645);
xor U27259 (N_27259,N_19851,N_18285);
or U27260 (N_27260,N_23700,N_19526);
nand U27261 (N_27261,N_21789,N_19743);
and U27262 (N_27262,N_22930,N_20121);
nor U27263 (N_27263,N_18364,N_23911);
and U27264 (N_27264,N_19808,N_21754);
nor U27265 (N_27265,N_22716,N_21225);
or U27266 (N_27266,N_21440,N_20198);
or U27267 (N_27267,N_19610,N_19394);
and U27268 (N_27268,N_18506,N_19082);
nand U27269 (N_27269,N_19061,N_19939);
or U27270 (N_27270,N_22405,N_23114);
xor U27271 (N_27271,N_21812,N_23093);
nor U27272 (N_27272,N_21726,N_19339);
xnor U27273 (N_27273,N_20619,N_19472);
or U27274 (N_27274,N_23912,N_21669);
xnor U27275 (N_27275,N_22959,N_19707);
or U27276 (N_27276,N_19198,N_20066);
nand U27277 (N_27277,N_21130,N_18714);
nor U27278 (N_27278,N_21317,N_21437);
xnor U27279 (N_27279,N_20829,N_21315);
nor U27280 (N_27280,N_23405,N_22870);
nand U27281 (N_27281,N_22682,N_21519);
xnor U27282 (N_27282,N_19758,N_19431);
and U27283 (N_27283,N_19224,N_21728);
or U27284 (N_27284,N_22923,N_23209);
nand U27285 (N_27285,N_23678,N_21492);
nand U27286 (N_27286,N_23613,N_19284);
xnor U27287 (N_27287,N_22889,N_18496);
nor U27288 (N_27288,N_22016,N_22753);
nor U27289 (N_27289,N_23739,N_18415);
and U27290 (N_27290,N_21608,N_23982);
nand U27291 (N_27291,N_20461,N_21858);
and U27292 (N_27292,N_18746,N_20754);
and U27293 (N_27293,N_22481,N_23712);
nor U27294 (N_27294,N_19417,N_19948);
nand U27295 (N_27295,N_22830,N_22776);
or U27296 (N_27296,N_22187,N_19891);
nand U27297 (N_27297,N_18776,N_21478);
nor U27298 (N_27298,N_22773,N_19537);
or U27299 (N_27299,N_21917,N_20985);
and U27300 (N_27300,N_23576,N_22251);
nand U27301 (N_27301,N_22018,N_18866);
nand U27302 (N_27302,N_23158,N_19092);
or U27303 (N_27303,N_23927,N_18440);
and U27304 (N_27304,N_23959,N_19728);
or U27305 (N_27305,N_22966,N_21588);
and U27306 (N_27306,N_18720,N_23839);
or U27307 (N_27307,N_19498,N_20813);
and U27308 (N_27308,N_23549,N_21271);
nor U27309 (N_27309,N_19022,N_19512);
or U27310 (N_27310,N_21425,N_20051);
nand U27311 (N_27311,N_22345,N_18983);
nor U27312 (N_27312,N_22821,N_21478);
and U27313 (N_27313,N_19752,N_22951);
nor U27314 (N_27314,N_21474,N_22372);
xnor U27315 (N_27315,N_19147,N_18497);
or U27316 (N_27316,N_20734,N_23473);
xor U27317 (N_27317,N_23083,N_21716);
or U27318 (N_27318,N_18367,N_20971);
and U27319 (N_27319,N_19738,N_23914);
xor U27320 (N_27320,N_19898,N_18799);
nor U27321 (N_27321,N_21896,N_20578);
or U27322 (N_27322,N_20940,N_22695);
or U27323 (N_27323,N_20596,N_19580);
or U27324 (N_27324,N_18076,N_23627);
xor U27325 (N_27325,N_23361,N_23382);
nor U27326 (N_27326,N_22687,N_20208);
nand U27327 (N_27327,N_22664,N_21260);
nor U27328 (N_27328,N_19759,N_20527);
xnor U27329 (N_27329,N_23120,N_20044);
nand U27330 (N_27330,N_20135,N_23062);
and U27331 (N_27331,N_22910,N_18704);
xnor U27332 (N_27332,N_22969,N_21896);
xor U27333 (N_27333,N_19305,N_19512);
or U27334 (N_27334,N_18271,N_18505);
xnor U27335 (N_27335,N_21386,N_21472);
nand U27336 (N_27336,N_22411,N_21181);
or U27337 (N_27337,N_22740,N_21863);
and U27338 (N_27338,N_19654,N_23989);
nor U27339 (N_27339,N_21458,N_19364);
xnor U27340 (N_27340,N_20469,N_23749);
and U27341 (N_27341,N_22017,N_20476);
and U27342 (N_27342,N_23972,N_18732);
nor U27343 (N_27343,N_19024,N_22304);
nor U27344 (N_27344,N_20246,N_22267);
xnor U27345 (N_27345,N_21956,N_23681);
or U27346 (N_27346,N_20109,N_22713);
nor U27347 (N_27347,N_23420,N_23516);
xnor U27348 (N_27348,N_21184,N_21339);
nor U27349 (N_27349,N_19731,N_23317);
xnor U27350 (N_27350,N_23486,N_22175);
and U27351 (N_27351,N_20002,N_18866);
nor U27352 (N_27352,N_21752,N_20079);
or U27353 (N_27353,N_21526,N_21498);
and U27354 (N_27354,N_21581,N_19419);
nand U27355 (N_27355,N_18632,N_21204);
xnor U27356 (N_27356,N_19416,N_23849);
and U27357 (N_27357,N_21405,N_21632);
nand U27358 (N_27358,N_22706,N_18131);
nor U27359 (N_27359,N_22724,N_21092);
or U27360 (N_27360,N_23796,N_20649);
or U27361 (N_27361,N_19603,N_18659);
and U27362 (N_27362,N_18348,N_19837);
nand U27363 (N_27363,N_23522,N_21028);
nand U27364 (N_27364,N_21745,N_20134);
and U27365 (N_27365,N_23357,N_18363);
xor U27366 (N_27366,N_23043,N_20158);
nand U27367 (N_27367,N_18778,N_22464);
or U27368 (N_27368,N_23145,N_21177);
or U27369 (N_27369,N_21268,N_19372);
nor U27370 (N_27370,N_23889,N_19337);
nand U27371 (N_27371,N_18792,N_21640);
nor U27372 (N_27372,N_19497,N_18293);
xnor U27373 (N_27373,N_18891,N_22006);
or U27374 (N_27374,N_18934,N_20038);
xnor U27375 (N_27375,N_21133,N_19812);
xnor U27376 (N_27376,N_20045,N_22921);
nand U27377 (N_27377,N_22383,N_18592);
xnor U27378 (N_27378,N_21360,N_22832);
and U27379 (N_27379,N_21215,N_23745);
xor U27380 (N_27380,N_22366,N_22712);
nor U27381 (N_27381,N_20392,N_22837);
nand U27382 (N_27382,N_23418,N_19800);
and U27383 (N_27383,N_18228,N_18478);
or U27384 (N_27384,N_23957,N_20119);
nor U27385 (N_27385,N_23395,N_22253);
and U27386 (N_27386,N_19397,N_23556);
xor U27387 (N_27387,N_22322,N_18459);
or U27388 (N_27388,N_18912,N_23952);
and U27389 (N_27389,N_21918,N_23429);
xor U27390 (N_27390,N_21184,N_21907);
and U27391 (N_27391,N_22093,N_22290);
and U27392 (N_27392,N_22187,N_21201);
or U27393 (N_27393,N_20749,N_21184);
or U27394 (N_27394,N_23442,N_18938);
or U27395 (N_27395,N_19585,N_21707);
and U27396 (N_27396,N_20953,N_20615);
xnor U27397 (N_27397,N_19203,N_23769);
and U27398 (N_27398,N_19695,N_22096);
nor U27399 (N_27399,N_23201,N_23596);
nor U27400 (N_27400,N_20264,N_18213);
or U27401 (N_27401,N_23340,N_23312);
xor U27402 (N_27402,N_22713,N_22802);
or U27403 (N_27403,N_22196,N_22223);
nand U27404 (N_27404,N_22961,N_19991);
xnor U27405 (N_27405,N_23088,N_22885);
xnor U27406 (N_27406,N_19512,N_23128);
nand U27407 (N_27407,N_23164,N_19985);
nor U27408 (N_27408,N_22339,N_22599);
nand U27409 (N_27409,N_21204,N_18875);
or U27410 (N_27410,N_20605,N_19737);
xnor U27411 (N_27411,N_22418,N_19965);
nor U27412 (N_27412,N_22947,N_19177);
or U27413 (N_27413,N_21724,N_21799);
or U27414 (N_27414,N_22698,N_20566);
and U27415 (N_27415,N_20188,N_20716);
nand U27416 (N_27416,N_20713,N_19885);
nor U27417 (N_27417,N_22095,N_22034);
nand U27418 (N_27418,N_23424,N_23477);
nand U27419 (N_27419,N_18747,N_18997);
or U27420 (N_27420,N_23779,N_22622);
xnor U27421 (N_27421,N_22969,N_22024);
and U27422 (N_27422,N_18795,N_19231);
nand U27423 (N_27423,N_19147,N_18225);
xnor U27424 (N_27424,N_21184,N_22497);
nand U27425 (N_27425,N_19517,N_18474);
xnor U27426 (N_27426,N_21916,N_19749);
nor U27427 (N_27427,N_20317,N_18672);
nor U27428 (N_27428,N_18778,N_19573);
xor U27429 (N_27429,N_21986,N_21543);
xor U27430 (N_27430,N_22612,N_22235);
xnor U27431 (N_27431,N_19353,N_18025);
nor U27432 (N_27432,N_21125,N_22220);
and U27433 (N_27433,N_21764,N_20866);
or U27434 (N_27434,N_22622,N_18883);
or U27435 (N_27435,N_18473,N_19686);
nand U27436 (N_27436,N_23275,N_21382);
xnor U27437 (N_27437,N_18481,N_18901);
or U27438 (N_27438,N_19521,N_20116);
nor U27439 (N_27439,N_23603,N_20317);
nor U27440 (N_27440,N_19216,N_21704);
or U27441 (N_27441,N_18774,N_18252);
and U27442 (N_27442,N_22972,N_23941);
xnor U27443 (N_27443,N_21902,N_18309);
nor U27444 (N_27444,N_23714,N_21635);
xnor U27445 (N_27445,N_18248,N_20536);
xor U27446 (N_27446,N_20870,N_20097);
xor U27447 (N_27447,N_21204,N_22585);
or U27448 (N_27448,N_22840,N_23695);
and U27449 (N_27449,N_19864,N_21081);
nand U27450 (N_27450,N_22222,N_23531);
nor U27451 (N_27451,N_19989,N_23687);
or U27452 (N_27452,N_20813,N_19451);
nand U27453 (N_27453,N_21765,N_21263);
xnor U27454 (N_27454,N_19511,N_21598);
nand U27455 (N_27455,N_20250,N_19444);
and U27456 (N_27456,N_22182,N_20155);
nand U27457 (N_27457,N_19278,N_18426);
nand U27458 (N_27458,N_20540,N_18486);
nor U27459 (N_27459,N_18722,N_22050);
and U27460 (N_27460,N_19697,N_22587);
or U27461 (N_27461,N_21248,N_23100);
and U27462 (N_27462,N_22213,N_18265);
xor U27463 (N_27463,N_18234,N_23385);
xor U27464 (N_27464,N_20687,N_19316);
or U27465 (N_27465,N_22715,N_22348);
nor U27466 (N_27466,N_19417,N_19640);
xor U27467 (N_27467,N_18486,N_22936);
nand U27468 (N_27468,N_22943,N_23749);
xor U27469 (N_27469,N_23062,N_20172);
xor U27470 (N_27470,N_23876,N_19768);
nor U27471 (N_27471,N_23208,N_18437);
or U27472 (N_27472,N_23216,N_23303);
or U27473 (N_27473,N_22166,N_19064);
xor U27474 (N_27474,N_22854,N_18166);
or U27475 (N_27475,N_21075,N_23653);
nand U27476 (N_27476,N_19470,N_19917);
xor U27477 (N_27477,N_22846,N_22570);
or U27478 (N_27478,N_20250,N_18867);
xnor U27479 (N_27479,N_23579,N_20966);
or U27480 (N_27480,N_18844,N_21791);
nand U27481 (N_27481,N_22842,N_20187);
nand U27482 (N_27482,N_21976,N_21409);
and U27483 (N_27483,N_20318,N_21542);
nand U27484 (N_27484,N_22862,N_19185);
or U27485 (N_27485,N_22133,N_21233);
nand U27486 (N_27486,N_18355,N_22465);
and U27487 (N_27487,N_23781,N_19993);
nor U27488 (N_27488,N_20314,N_19528);
or U27489 (N_27489,N_23382,N_20732);
nand U27490 (N_27490,N_23157,N_19109);
xnor U27491 (N_27491,N_18587,N_18935);
or U27492 (N_27492,N_20735,N_19733);
or U27493 (N_27493,N_23360,N_20659);
xor U27494 (N_27494,N_23908,N_18590);
nand U27495 (N_27495,N_18027,N_19516);
nor U27496 (N_27496,N_20555,N_20157);
nand U27497 (N_27497,N_22051,N_21395);
or U27498 (N_27498,N_22029,N_21591);
and U27499 (N_27499,N_21179,N_23214);
xnor U27500 (N_27500,N_19385,N_19178);
nor U27501 (N_27501,N_19566,N_22003);
and U27502 (N_27502,N_23371,N_22954);
xor U27503 (N_27503,N_23331,N_19009);
nand U27504 (N_27504,N_23604,N_23372);
and U27505 (N_27505,N_20626,N_18878);
nand U27506 (N_27506,N_20866,N_21860);
and U27507 (N_27507,N_22659,N_18803);
xnor U27508 (N_27508,N_19336,N_21323);
nand U27509 (N_27509,N_18039,N_18145);
and U27510 (N_27510,N_20728,N_22927);
and U27511 (N_27511,N_20856,N_23977);
or U27512 (N_27512,N_21425,N_19019);
and U27513 (N_27513,N_19643,N_20512);
xnor U27514 (N_27514,N_20992,N_18898);
or U27515 (N_27515,N_21831,N_19772);
and U27516 (N_27516,N_20867,N_19915);
or U27517 (N_27517,N_22114,N_21604);
and U27518 (N_27518,N_23836,N_23180);
nor U27519 (N_27519,N_22317,N_19520);
nor U27520 (N_27520,N_18861,N_21952);
or U27521 (N_27521,N_21504,N_20703);
nand U27522 (N_27522,N_19346,N_20740);
nor U27523 (N_27523,N_18094,N_20062);
and U27524 (N_27524,N_21735,N_20565);
nand U27525 (N_27525,N_23321,N_23645);
nand U27526 (N_27526,N_18014,N_23700);
xor U27527 (N_27527,N_21226,N_22069);
nor U27528 (N_27528,N_19836,N_22840);
or U27529 (N_27529,N_23087,N_20112);
and U27530 (N_27530,N_20550,N_18871);
or U27531 (N_27531,N_23745,N_18653);
nand U27532 (N_27532,N_20913,N_21126);
xor U27533 (N_27533,N_22478,N_19263);
nor U27534 (N_27534,N_20861,N_21811);
nand U27535 (N_27535,N_21342,N_20904);
nor U27536 (N_27536,N_19440,N_21142);
nor U27537 (N_27537,N_21749,N_19455);
or U27538 (N_27538,N_20539,N_19564);
or U27539 (N_27539,N_22984,N_21733);
and U27540 (N_27540,N_22702,N_20611);
and U27541 (N_27541,N_20306,N_18267);
or U27542 (N_27542,N_21906,N_21689);
and U27543 (N_27543,N_22729,N_18703);
nand U27544 (N_27544,N_21071,N_23090);
nor U27545 (N_27545,N_19772,N_23172);
nand U27546 (N_27546,N_21089,N_23078);
or U27547 (N_27547,N_19743,N_20150);
nand U27548 (N_27548,N_20347,N_22691);
or U27549 (N_27549,N_18735,N_22092);
nand U27550 (N_27550,N_21013,N_21770);
nand U27551 (N_27551,N_20148,N_19102);
or U27552 (N_27552,N_21249,N_20682);
or U27553 (N_27553,N_21962,N_19526);
xor U27554 (N_27554,N_21668,N_22965);
or U27555 (N_27555,N_20668,N_22859);
or U27556 (N_27556,N_21080,N_19462);
nor U27557 (N_27557,N_21581,N_22438);
or U27558 (N_27558,N_19977,N_21506);
xor U27559 (N_27559,N_20162,N_23989);
nand U27560 (N_27560,N_19943,N_21126);
nand U27561 (N_27561,N_18315,N_22824);
or U27562 (N_27562,N_19046,N_21783);
and U27563 (N_27563,N_23772,N_23388);
nand U27564 (N_27564,N_20824,N_20837);
and U27565 (N_27565,N_23094,N_20903);
xor U27566 (N_27566,N_22436,N_21252);
nand U27567 (N_27567,N_22311,N_20796);
or U27568 (N_27568,N_23147,N_19609);
and U27569 (N_27569,N_20179,N_21977);
xor U27570 (N_27570,N_21637,N_20539);
nor U27571 (N_27571,N_23666,N_21448);
nor U27572 (N_27572,N_18096,N_21770);
xnor U27573 (N_27573,N_23426,N_23109);
or U27574 (N_27574,N_22203,N_18693);
and U27575 (N_27575,N_23617,N_20365);
and U27576 (N_27576,N_18950,N_20720);
and U27577 (N_27577,N_23359,N_23143);
and U27578 (N_27578,N_18875,N_21534);
nor U27579 (N_27579,N_18974,N_20153);
and U27580 (N_27580,N_22807,N_22101);
or U27581 (N_27581,N_21722,N_22064);
or U27582 (N_27582,N_19518,N_22924);
nor U27583 (N_27583,N_19156,N_19845);
nor U27584 (N_27584,N_21240,N_19894);
and U27585 (N_27585,N_18561,N_23889);
nand U27586 (N_27586,N_20270,N_20913);
or U27587 (N_27587,N_23176,N_18453);
and U27588 (N_27588,N_18267,N_19867);
or U27589 (N_27589,N_22687,N_23329);
or U27590 (N_27590,N_20714,N_18424);
nor U27591 (N_27591,N_18490,N_19424);
xnor U27592 (N_27592,N_22482,N_18985);
xor U27593 (N_27593,N_21954,N_23243);
nand U27594 (N_27594,N_22610,N_19572);
and U27595 (N_27595,N_18838,N_21243);
and U27596 (N_27596,N_22029,N_21637);
nand U27597 (N_27597,N_19536,N_19584);
nand U27598 (N_27598,N_22318,N_23936);
nand U27599 (N_27599,N_20271,N_20135);
or U27600 (N_27600,N_21049,N_22239);
and U27601 (N_27601,N_19668,N_23547);
xor U27602 (N_27602,N_22986,N_20326);
xnor U27603 (N_27603,N_18324,N_18779);
nand U27604 (N_27604,N_21083,N_18299);
nor U27605 (N_27605,N_21610,N_18685);
and U27606 (N_27606,N_23096,N_21113);
nand U27607 (N_27607,N_23531,N_22669);
xnor U27608 (N_27608,N_20225,N_23419);
nand U27609 (N_27609,N_22851,N_20930);
or U27610 (N_27610,N_23552,N_21914);
nand U27611 (N_27611,N_22499,N_22233);
xnor U27612 (N_27612,N_22444,N_23627);
and U27613 (N_27613,N_18449,N_23470);
xnor U27614 (N_27614,N_20750,N_18088);
nand U27615 (N_27615,N_23302,N_23240);
nor U27616 (N_27616,N_22215,N_21166);
xnor U27617 (N_27617,N_22285,N_19943);
nand U27618 (N_27618,N_23294,N_21021);
xnor U27619 (N_27619,N_22774,N_19455);
xor U27620 (N_27620,N_20375,N_19824);
xor U27621 (N_27621,N_18020,N_20608);
nand U27622 (N_27622,N_21759,N_19703);
and U27623 (N_27623,N_21525,N_20742);
xor U27624 (N_27624,N_20255,N_23913);
xor U27625 (N_27625,N_19345,N_18033);
or U27626 (N_27626,N_21095,N_21316);
nand U27627 (N_27627,N_23527,N_23457);
and U27628 (N_27628,N_20199,N_23839);
xor U27629 (N_27629,N_23266,N_20804);
nand U27630 (N_27630,N_18353,N_20293);
nand U27631 (N_27631,N_23195,N_23087);
and U27632 (N_27632,N_19375,N_23535);
or U27633 (N_27633,N_19133,N_21706);
and U27634 (N_27634,N_19029,N_23301);
xnor U27635 (N_27635,N_20424,N_21419);
or U27636 (N_27636,N_22935,N_22825);
and U27637 (N_27637,N_22815,N_19257);
nor U27638 (N_27638,N_20222,N_23826);
and U27639 (N_27639,N_19830,N_22720);
and U27640 (N_27640,N_23964,N_18754);
or U27641 (N_27641,N_21442,N_22175);
nand U27642 (N_27642,N_22662,N_22989);
and U27643 (N_27643,N_23263,N_20550);
xor U27644 (N_27644,N_18604,N_23596);
nor U27645 (N_27645,N_18053,N_23108);
nand U27646 (N_27646,N_19089,N_23167);
nor U27647 (N_27647,N_20504,N_22073);
and U27648 (N_27648,N_23707,N_19210);
and U27649 (N_27649,N_18474,N_20318);
nor U27650 (N_27650,N_21039,N_18143);
nor U27651 (N_27651,N_23166,N_22621);
and U27652 (N_27652,N_19191,N_19772);
xnor U27653 (N_27653,N_19704,N_18262);
or U27654 (N_27654,N_20014,N_20449);
and U27655 (N_27655,N_18259,N_20963);
or U27656 (N_27656,N_22217,N_22788);
or U27657 (N_27657,N_23084,N_21923);
xor U27658 (N_27658,N_21978,N_18407);
and U27659 (N_27659,N_22502,N_18489);
or U27660 (N_27660,N_21352,N_21704);
and U27661 (N_27661,N_20945,N_23029);
nor U27662 (N_27662,N_21298,N_21384);
xor U27663 (N_27663,N_23426,N_18909);
nand U27664 (N_27664,N_20545,N_21961);
nor U27665 (N_27665,N_18145,N_18183);
nor U27666 (N_27666,N_23973,N_21104);
xor U27667 (N_27667,N_22371,N_18378);
and U27668 (N_27668,N_22427,N_18691);
nor U27669 (N_27669,N_21184,N_20182);
and U27670 (N_27670,N_22761,N_21759);
or U27671 (N_27671,N_22050,N_19867);
nand U27672 (N_27672,N_18649,N_23859);
xor U27673 (N_27673,N_21627,N_20335);
xnor U27674 (N_27674,N_21353,N_18276);
xnor U27675 (N_27675,N_21056,N_23140);
and U27676 (N_27676,N_20340,N_18005);
xnor U27677 (N_27677,N_22167,N_18376);
nand U27678 (N_27678,N_22603,N_20776);
nand U27679 (N_27679,N_20820,N_23585);
nor U27680 (N_27680,N_22444,N_19691);
and U27681 (N_27681,N_23345,N_19052);
xor U27682 (N_27682,N_19835,N_20355);
xnor U27683 (N_27683,N_22292,N_21432);
xor U27684 (N_27684,N_18079,N_21586);
and U27685 (N_27685,N_20534,N_19315);
nor U27686 (N_27686,N_19488,N_18874);
xor U27687 (N_27687,N_18370,N_23502);
nor U27688 (N_27688,N_18693,N_18832);
xnor U27689 (N_27689,N_20385,N_22474);
nor U27690 (N_27690,N_18839,N_21903);
nor U27691 (N_27691,N_23796,N_21868);
xnor U27692 (N_27692,N_20245,N_21287);
nor U27693 (N_27693,N_20076,N_19564);
nand U27694 (N_27694,N_23003,N_20155);
xnor U27695 (N_27695,N_19886,N_18125);
and U27696 (N_27696,N_22952,N_19106);
nor U27697 (N_27697,N_21976,N_20033);
xor U27698 (N_27698,N_22307,N_22553);
nor U27699 (N_27699,N_21520,N_18052);
xnor U27700 (N_27700,N_20890,N_23864);
nor U27701 (N_27701,N_23099,N_18386);
nand U27702 (N_27702,N_21027,N_21239);
or U27703 (N_27703,N_23296,N_19714);
xor U27704 (N_27704,N_18414,N_20552);
nor U27705 (N_27705,N_22719,N_23913);
nor U27706 (N_27706,N_20631,N_22768);
xnor U27707 (N_27707,N_18853,N_23730);
or U27708 (N_27708,N_19512,N_21049);
or U27709 (N_27709,N_18728,N_22709);
and U27710 (N_27710,N_19884,N_20303);
xor U27711 (N_27711,N_19363,N_18677);
nor U27712 (N_27712,N_22145,N_22985);
or U27713 (N_27713,N_21855,N_22911);
xor U27714 (N_27714,N_23623,N_22581);
or U27715 (N_27715,N_21706,N_18681);
xor U27716 (N_27716,N_20136,N_23102);
nand U27717 (N_27717,N_22666,N_22366);
and U27718 (N_27718,N_20322,N_19050);
nor U27719 (N_27719,N_18956,N_23734);
xor U27720 (N_27720,N_19491,N_21186);
or U27721 (N_27721,N_19733,N_23266);
nor U27722 (N_27722,N_21243,N_22969);
nand U27723 (N_27723,N_20502,N_18863);
xor U27724 (N_27724,N_20058,N_23056);
nand U27725 (N_27725,N_22271,N_22344);
nand U27726 (N_27726,N_18777,N_20510);
or U27727 (N_27727,N_20362,N_19068);
nand U27728 (N_27728,N_19114,N_19442);
xor U27729 (N_27729,N_23809,N_21968);
nand U27730 (N_27730,N_23193,N_18473);
xor U27731 (N_27731,N_20794,N_21323);
and U27732 (N_27732,N_18580,N_20612);
and U27733 (N_27733,N_20808,N_23787);
xor U27734 (N_27734,N_23871,N_18253);
nand U27735 (N_27735,N_18269,N_21401);
xnor U27736 (N_27736,N_19057,N_20951);
and U27737 (N_27737,N_19812,N_23323);
or U27738 (N_27738,N_21170,N_23685);
xnor U27739 (N_27739,N_20385,N_22276);
xnor U27740 (N_27740,N_23059,N_19683);
or U27741 (N_27741,N_23460,N_21748);
nand U27742 (N_27742,N_18266,N_18719);
xnor U27743 (N_27743,N_23059,N_19101);
and U27744 (N_27744,N_20307,N_18092);
xor U27745 (N_27745,N_23483,N_18301);
or U27746 (N_27746,N_21794,N_21250);
xnor U27747 (N_27747,N_20991,N_23769);
nor U27748 (N_27748,N_18650,N_21595);
or U27749 (N_27749,N_23080,N_19980);
nor U27750 (N_27750,N_23098,N_23078);
and U27751 (N_27751,N_18849,N_18619);
or U27752 (N_27752,N_21623,N_22002);
and U27753 (N_27753,N_22846,N_21012);
xor U27754 (N_27754,N_21783,N_18087);
and U27755 (N_27755,N_21339,N_21007);
nand U27756 (N_27756,N_22317,N_18025);
xnor U27757 (N_27757,N_19720,N_18706);
nor U27758 (N_27758,N_19622,N_20429);
nand U27759 (N_27759,N_21696,N_23882);
or U27760 (N_27760,N_19377,N_21777);
and U27761 (N_27761,N_23464,N_23783);
and U27762 (N_27762,N_20518,N_19039);
and U27763 (N_27763,N_20723,N_18686);
and U27764 (N_27764,N_19976,N_22047);
nor U27765 (N_27765,N_23242,N_19525);
and U27766 (N_27766,N_19767,N_19200);
nand U27767 (N_27767,N_22533,N_21890);
nand U27768 (N_27768,N_23433,N_18276);
nor U27769 (N_27769,N_19131,N_21559);
or U27770 (N_27770,N_20500,N_21641);
nand U27771 (N_27771,N_23783,N_20163);
and U27772 (N_27772,N_22242,N_21331);
nor U27773 (N_27773,N_22180,N_21335);
nor U27774 (N_27774,N_23541,N_23768);
nand U27775 (N_27775,N_18885,N_19171);
nor U27776 (N_27776,N_23172,N_23193);
or U27777 (N_27777,N_20026,N_19864);
xor U27778 (N_27778,N_22365,N_19495);
nor U27779 (N_27779,N_23706,N_23243);
xnor U27780 (N_27780,N_20282,N_23413);
nand U27781 (N_27781,N_18751,N_20312);
and U27782 (N_27782,N_20038,N_22724);
xor U27783 (N_27783,N_20394,N_21114);
nor U27784 (N_27784,N_23044,N_18111);
nor U27785 (N_27785,N_21981,N_21179);
nor U27786 (N_27786,N_23055,N_23517);
xnor U27787 (N_27787,N_18563,N_21349);
xnor U27788 (N_27788,N_19133,N_22621);
nand U27789 (N_27789,N_20447,N_18451);
and U27790 (N_27790,N_19989,N_20012);
nor U27791 (N_27791,N_23969,N_18049);
nand U27792 (N_27792,N_20861,N_21617);
nor U27793 (N_27793,N_23223,N_21039);
nand U27794 (N_27794,N_21955,N_18795);
nor U27795 (N_27795,N_20564,N_20043);
nor U27796 (N_27796,N_19925,N_20395);
or U27797 (N_27797,N_20750,N_23152);
xor U27798 (N_27798,N_21498,N_19323);
xor U27799 (N_27799,N_21945,N_21680);
and U27800 (N_27800,N_22319,N_21053);
nand U27801 (N_27801,N_20265,N_18756);
nand U27802 (N_27802,N_18118,N_21949);
nor U27803 (N_27803,N_18720,N_22170);
nor U27804 (N_27804,N_18524,N_19161);
nor U27805 (N_27805,N_22889,N_22869);
or U27806 (N_27806,N_19962,N_21275);
or U27807 (N_27807,N_20951,N_18215);
nor U27808 (N_27808,N_20760,N_19268);
nand U27809 (N_27809,N_21943,N_18037);
or U27810 (N_27810,N_22485,N_22482);
nor U27811 (N_27811,N_21865,N_19463);
nor U27812 (N_27812,N_22825,N_18883);
and U27813 (N_27813,N_19071,N_20514);
and U27814 (N_27814,N_19131,N_23793);
xor U27815 (N_27815,N_22963,N_20340);
nor U27816 (N_27816,N_19965,N_22948);
or U27817 (N_27817,N_21135,N_22000);
nor U27818 (N_27818,N_20728,N_22936);
xor U27819 (N_27819,N_20217,N_20242);
xor U27820 (N_27820,N_22902,N_19886);
and U27821 (N_27821,N_20036,N_22238);
and U27822 (N_27822,N_22082,N_22147);
nand U27823 (N_27823,N_23840,N_19679);
and U27824 (N_27824,N_21163,N_23093);
or U27825 (N_27825,N_18974,N_22187);
nand U27826 (N_27826,N_19626,N_19476);
nand U27827 (N_27827,N_23165,N_20550);
nand U27828 (N_27828,N_22980,N_23111);
nand U27829 (N_27829,N_20391,N_21351);
or U27830 (N_27830,N_23699,N_18704);
xor U27831 (N_27831,N_20830,N_18010);
and U27832 (N_27832,N_22237,N_19931);
nand U27833 (N_27833,N_23522,N_19009);
xor U27834 (N_27834,N_20858,N_21096);
nor U27835 (N_27835,N_23052,N_20514);
nor U27836 (N_27836,N_22353,N_23631);
nand U27837 (N_27837,N_21675,N_23434);
nor U27838 (N_27838,N_22849,N_18466);
and U27839 (N_27839,N_21193,N_21876);
nand U27840 (N_27840,N_20108,N_18222);
and U27841 (N_27841,N_18437,N_20081);
nor U27842 (N_27842,N_23119,N_21556);
nor U27843 (N_27843,N_18350,N_20281);
or U27844 (N_27844,N_20991,N_19097);
nor U27845 (N_27845,N_23432,N_18389);
or U27846 (N_27846,N_22971,N_23499);
or U27847 (N_27847,N_22153,N_18200);
nor U27848 (N_27848,N_19374,N_18028);
and U27849 (N_27849,N_19548,N_19488);
nor U27850 (N_27850,N_19478,N_22352);
nor U27851 (N_27851,N_18050,N_19269);
and U27852 (N_27852,N_21674,N_21078);
nor U27853 (N_27853,N_19061,N_23356);
nor U27854 (N_27854,N_20581,N_19210);
xnor U27855 (N_27855,N_22118,N_21792);
and U27856 (N_27856,N_22778,N_20777);
or U27857 (N_27857,N_20786,N_19320);
nand U27858 (N_27858,N_19147,N_22304);
xor U27859 (N_27859,N_18240,N_21526);
and U27860 (N_27860,N_19534,N_21627);
and U27861 (N_27861,N_23322,N_21865);
and U27862 (N_27862,N_22085,N_19460);
nand U27863 (N_27863,N_19596,N_20659);
or U27864 (N_27864,N_19532,N_20309);
nor U27865 (N_27865,N_18810,N_19695);
xnor U27866 (N_27866,N_22238,N_20690);
nor U27867 (N_27867,N_23772,N_23527);
nand U27868 (N_27868,N_23766,N_19594);
nor U27869 (N_27869,N_20026,N_20046);
and U27870 (N_27870,N_19852,N_19403);
nand U27871 (N_27871,N_19403,N_21299);
xnor U27872 (N_27872,N_22107,N_22538);
nand U27873 (N_27873,N_19523,N_19878);
and U27874 (N_27874,N_22105,N_20220);
and U27875 (N_27875,N_21864,N_22942);
xnor U27876 (N_27876,N_23735,N_23378);
or U27877 (N_27877,N_23849,N_22553);
and U27878 (N_27878,N_18445,N_22119);
nand U27879 (N_27879,N_22564,N_18757);
and U27880 (N_27880,N_18031,N_20505);
nand U27881 (N_27881,N_21063,N_23436);
xnor U27882 (N_27882,N_18371,N_20970);
xnor U27883 (N_27883,N_22238,N_19243);
and U27884 (N_27884,N_23865,N_20161);
or U27885 (N_27885,N_18355,N_22311);
nand U27886 (N_27886,N_20104,N_23379);
nor U27887 (N_27887,N_19883,N_20819);
nand U27888 (N_27888,N_19146,N_22828);
and U27889 (N_27889,N_20889,N_21382);
nor U27890 (N_27890,N_18820,N_22257);
nand U27891 (N_27891,N_18909,N_23895);
and U27892 (N_27892,N_20138,N_23998);
or U27893 (N_27893,N_22965,N_18368);
xor U27894 (N_27894,N_22381,N_20436);
xor U27895 (N_27895,N_22762,N_19929);
nor U27896 (N_27896,N_19460,N_22487);
nand U27897 (N_27897,N_18926,N_22192);
nor U27898 (N_27898,N_18140,N_23271);
nand U27899 (N_27899,N_22076,N_23974);
nor U27900 (N_27900,N_23367,N_19315);
nand U27901 (N_27901,N_18053,N_19878);
and U27902 (N_27902,N_22798,N_21618);
nand U27903 (N_27903,N_22047,N_22613);
nand U27904 (N_27904,N_22286,N_20703);
and U27905 (N_27905,N_21258,N_19874);
nor U27906 (N_27906,N_23480,N_18635);
nor U27907 (N_27907,N_21900,N_23850);
or U27908 (N_27908,N_23284,N_19008);
nand U27909 (N_27909,N_22904,N_23127);
nand U27910 (N_27910,N_19599,N_23495);
or U27911 (N_27911,N_22725,N_19532);
nor U27912 (N_27912,N_19657,N_19146);
nand U27913 (N_27913,N_19521,N_19353);
and U27914 (N_27914,N_23732,N_21663);
nor U27915 (N_27915,N_23215,N_21653);
xor U27916 (N_27916,N_21762,N_20711);
and U27917 (N_27917,N_21357,N_20034);
nand U27918 (N_27918,N_20831,N_23955);
nand U27919 (N_27919,N_22145,N_21246);
xnor U27920 (N_27920,N_19834,N_19046);
xnor U27921 (N_27921,N_21503,N_20633);
and U27922 (N_27922,N_21949,N_20867);
xnor U27923 (N_27923,N_19949,N_19601);
nor U27924 (N_27924,N_18307,N_23152);
or U27925 (N_27925,N_20466,N_21757);
and U27926 (N_27926,N_18724,N_21644);
xor U27927 (N_27927,N_21322,N_21346);
and U27928 (N_27928,N_19578,N_21145);
nor U27929 (N_27929,N_21471,N_22597);
nand U27930 (N_27930,N_21818,N_19791);
or U27931 (N_27931,N_22337,N_22605);
nor U27932 (N_27932,N_21084,N_18091);
nor U27933 (N_27933,N_23097,N_20118);
or U27934 (N_27934,N_20890,N_22272);
xnor U27935 (N_27935,N_19443,N_18086);
and U27936 (N_27936,N_18717,N_19087);
xor U27937 (N_27937,N_20838,N_18792);
nand U27938 (N_27938,N_18657,N_23242);
xor U27939 (N_27939,N_19240,N_20981);
nand U27940 (N_27940,N_22693,N_21669);
and U27941 (N_27941,N_23157,N_18087);
or U27942 (N_27942,N_20848,N_21570);
xnor U27943 (N_27943,N_18457,N_23349);
xnor U27944 (N_27944,N_19803,N_21147);
or U27945 (N_27945,N_20654,N_21612);
or U27946 (N_27946,N_22389,N_23627);
nand U27947 (N_27947,N_19896,N_18750);
xor U27948 (N_27948,N_22106,N_18830);
nand U27949 (N_27949,N_19878,N_19032);
nor U27950 (N_27950,N_23490,N_20045);
or U27951 (N_27951,N_21435,N_23114);
nor U27952 (N_27952,N_20101,N_18065);
and U27953 (N_27953,N_18493,N_22524);
nand U27954 (N_27954,N_21653,N_21901);
xor U27955 (N_27955,N_19379,N_22619);
or U27956 (N_27956,N_21911,N_23666);
nand U27957 (N_27957,N_19678,N_19635);
xnor U27958 (N_27958,N_18429,N_20945);
and U27959 (N_27959,N_20649,N_19995);
nand U27960 (N_27960,N_21137,N_23261);
or U27961 (N_27961,N_21328,N_23296);
nor U27962 (N_27962,N_23729,N_18043);
nor U27963 (N_27963,N_22099,N_21415);
nand U27964 (N_27964,N_23748,N_21085);
nand U27965 (N_27965,N_19524,N_18748);
nand U27966 (N_27966,N_21123,N_23965);
xnor U27967 (N_27967,N_18775,N_23586);
nor U27968 (N_27968,N_19079,N_22815);
nor U27969 (N_27969,N_20131,N_18480);
xnor U27970 (N_27970,N_23536,N_19934);
nor U27971 (N_27971,N_23687,N_18130);
xnor U27972 (N_27972,N_22585,N_22907);
xor U27973 (N_27973,N_20679,N_19459);
or U27974 (N_27974,N_22046,N_20271);
and U27975 (N_27975,N_22620,N_18229);
nor U27976 (N_27976,N_20377,N_20996);
nor U27977 (N_27977,N_21226,N_23503);
and U27978 (N_27978,N_21134,N_20368);
xnor U27979 (N_27979,N_22641,N_21442);
xnor U27980 (N_27980,N_20654,N_20612);
or U27981 (N_27981,N_18257,N_18422);
and U27982 (N_27982,N_21281,N_20521);
and U27983 (N_27983,N_21001,N_21612);
or U27984 (N_27984,N_18192,N_21029);
nor U27985 (N_27985,N_22284,N_21620);
xnor U27986 (N_27986,N_21545,N_18038);
nor U27987 (N_27987,N_19652,N_23137);
nor U27988 (N_27988,N_20949,N_19013);
nor U27989 (N_27989,N_21792,N_20761);
xnor U27990 (N_27990,N_20447,N_18351);
nand U27991 (N_27991,N_20788,N_21610);
or U27992 (N_27992,N_23478,N_23095);
or U27993 (N_27993,N_19402,N_22749);
nor U27994 (N_27994,N_21250,N_21512);
nand U27995 (N_27995,N_22630,N_22760);
nand U27996 (N_27996,N_23951,N_19981);
nor U27997 (N_27997,N_20035,N_23330);
and U27998 (N_27998,N_22474,N_18996);
and U27999 (N_27999,N_18771,N_21878);
or U28000 (N_28000,N_18169,N_21109);
xnor U28001 (N_28001,N_23413,N_22347);
nand U28002 (N_28002,N_19422,N_21035);
nand U28003 (N_28003,N_19381,N_20471);
nor U28004 (N_28004,N_22564,N_22555);
and U28005 (N_28005,N_18134,N_21974);
nor U28006 (N_28006,N_19299,N_19903);
xnor U28007 (N_28007,N_22231,N_18686);
nor U28008 (N_28008,N_21018,N_18780);
nand U28009 (N_28009,N_20895,N_18846);
and U28010 (N_28010,N_21393,N_19033);
nor U28011 (N_28011,N_18150,N_18228);
nand U28012 (N_28012,N_21805,N_23379);
xor U28013 (N_28013,N_18902,N_21488);
nand U28014 (N_28014,N_23648,N_19221);
nand U28015 (N_28015,N_20333,N_19210);
nor U28016 (N_28016,N_22606,N_19069);
nor U28017 (N_28017,N_20225,N_19214);
nor U28018 (N_28018,N_23252,N_21853);
nor U28019 (N_28019,N_23534,N_20060);
and U28020 (N_28020,N_19499,N_23352);
xor U28021 (N_28021,N_21362,N_19176);
and U28022 (N_28022,N_23896,N_20132);
or U28023 (N_28023,N_20110,N_21822);
and U28024 (N_28024,N_23176,N_18326);
nor U28025 (N_28025,N_22678,N_18737);
or U28026 (N_28026,N_18410,N_18318);
xor U28027 (N_28027,N_18946,N_19438);
nor U28028 (N_28028,N_20855,N_20040);
nor U28029 (N_28029,N_22509,N_18933);
and U28030 (N_28030,N_23676,N_19000);
nand U28031 (N_28031,N_23671,N_21902);
xnor U28032 (N_28032,N_18398,N_20866);
and U28033 (N_28033,N_22803,N_23352);
xnor U28034 (N_28034,N_19377,N_21998);
and U28035 (N_28035,N_18038,N_23608);
nor U28036 (N_28036,N_23803,N_21007);
or U28037 (N_28037,N_18443,N_23113);
nand U28038 (N_28038,N_21203,N_22540);
nor U28039 (N_28039,N_22569,N_18862);
nand U28040 (N_28040,N_22957,N_21920);
nand U28041 (N_28041,N_19667,N_21019);
nor U28042 (N_28042,N_23924,N_19972);
and U28043 (N_28043,N_18120,N_21991);
or U28044 (N_28044,N_21296,N_21171);
nor U28045 (N_28045,N_18141,N_21472);
or U28046 (N_28046,N_23063,N_18280);
or U28047 (N_28047,N_23452,N_22653);
xor U28048 (N_28048,N_22243,N_23085);
xnor U28049 (N_28049,N_20248,N_18943);
xor U28050 (N_28050,N_19862,N_21674);
or U28051 (N_28051,N_21392,N_20356);
xnor U28052 (N_28052,N_20056,N_19358);
nor U28053 (N_28053,N_19385,N_21568);
or U28054 (N_28054,N_21452,N_19834);
xnor U28055 (N_28055,N_22411,N_18838);
xor U28056 (N_28056,N_22172,N_21101);
or U28057 (N_28057,N_23260,N_18605);
nand U28058 (N_28058,N_19797,N_22290);
nand U28059 (N_28059,N_20704,N_22294);
xnor U28060 (N_28060,N_19800,N_23067);
xor U28061 (N_28061,N_22210,N_23648);
nor U28062 (N_28062,N_18793,N_21200);
nor U28063 (N_28063,N_23605,N_23727);
and U28064 (N_28064,N_22432,N_20361);
and U28065 (N_28065,N_22030,N_18344);
and U28066 (N_28066,N_20891,N_20997);
nor U28067 (N_28067,N_20606,N_18028);
nor U28068 (N_28068,N_20997,N_21557);
xnor U28069 (N_28069,N_20453,N_21671);
nand U28070 (N_28070,N_18066,N_19834);
xnor U28071 (N_28071,N_19665,N_19542);
xor U28072 (N_28072,N_23199,N_20238);
nor U28073 (N_28073,N_22697,N_19028);
nand U28074 (N_28074,N_22183,N_20097);
nand U28075 (N_28075,N_20590,N_18958);
nor U28076 (N_28076,N_19178,N_21071);
nand U28077 (N_28077,N_18260,N_18714);
nor U28078 (N_28078,N_20848,N_20840);
nand U28079 (N_28079,N_19608,N_18877);
or U28080 (N_28080,N_23101,N_18207);
or U28081 (N_28081,N_23202,N_23340);
nand U28082 (N_28082,N_18496,N_19077);
or U28083 (N_28083,N_19173,N_23061);
xor U28084 (N_28084,N_19118,N_20790);
xor U28085 (N_28085,N_21518,N_22357);
nand U28086 (N_28086,N_23739,N_21616);
xnor U28087 (N_28087,N_22955,N_21636);
or U28088 (N_28088,N_20598,N_18129);
or U28089 (N_28089,N_23816,N_18270);
nor U28090 (N_28090,N_20461,N_18713);
xor U28091 (N_28091,N_18637,N_22985);
nor U28092 (N_28092,N_18845,N_22796);
and U28093 (N_28093,N_20247,N_22836);
xnor U28094 (N_28094,N_21545,N_21558);
nor U28095 (N_28095,N_21957,N_21322);
nand U28096 (N_28096,N_21146,N_20842);
nor U28097 (N_28097,N_21435,N_18257);
nor U28098 (N_28098,N_19472,N_20603);
or U28099 (N_28099,N_19053,N_21072);
or U28100 (N_28100,N_20286,N_23192);
and U28101 (N_28101,N_18070,N_20908);
xnor U28102 (N_28102,N_22202,N_20345);
or U28103 (N_28103,N_22820,N_19220);
and U28104 (N_28104,N_18840,N_19935);
xor U28105 (N_28105,N_20650,N_21631);
nand U28106 (N_28106,N_20988,N_19299);
and U28107 (N_28107,N_21241,N_20159);
and U28108 (N_28108,N_23782,N_21319);
nand U28109 (N_28109,N_21606,N_20142);
xor U28110 (N_28110,N_20692,N_20970);
nand U28111 (N_28111,N_22165,N_20781);
or U28112 (N_28112,N_23127,N_19613);
xor U28113 (N_28113,N_19309,N_22156);
xnor U28114 (N_28114,N_21934,N_18415);
nand U28115 (N_28115,N_22500,N_21419);
or U28116 (N_28116,N_23587,N_19522);
nor U28117 (N_28117,N_19080,N_21263);
xnor U28118 (N_28118,N_22688,N_23121);
and U28119 (N_28119,N_20383,N_19326);
xnor U28120 (N_28120,N_21278,N_21587);
and U28121 (N_28121,N_22229,N_22371);
or U28122 (N_28122,N_20090,N_21743);
nand U28123 (N_28123,N_21617,N_19954);
and U28124 (N_28124,N_21299,N_18875);
nor U28125 (N_28125,N_21343,N_18995);
xor U28126 (N_28126,N_23665,N_22772);
or U28127 (N_28127,N_18632,N_18624);
xor U28128 (N_28128,N_21645,N_18375);
nand U28129 (N_28129,N_19007,N_19747);
xor U28130 (N_28130,N_22218,N_23612);
xor U28131 (N_28131,N_20433,N_18465);
nand U28132 (N_28132,N_22305,N_22014);
and U28133 (N_28133,N_19511,N_20207);
or U28134 (N_28134,N_19076,N_18959);
and U28135 (N_28135,N_19855,N_21454);
xor U28136 (N_28136,N_19570,N_20964);
or U28137 (N_28137,N_22535,N_23087);
and U28138 (N_28138,N_18388,N_18783);
or U28139 (N_28139,N_22897,N_21591);
nand U28140 (N_28140,N_22499,N_23869);
nand U28141 (N_28141,N_21526,N_21338);
or U28142 (N_28142,N_18188,N_20938);
or U28143 (N_28143,N_20086,N_23736);
and U28144 (N_28144,N_18115,N_20128);
xor U28145 (N_28145,N_22340,N_19514);
or U28146 (N_28146,N_19891,N_19640);
and U28147 (N_28147,N_19287,N_19140);
nor U28148 (N_28148,N_23239,N_19125);
and U28149 (N_28149,N_23258,N_22676);
xor U28150 (N_28150,N_23236,N_20784);
nand U28151 (N_28151,N_23060,N_21180);
and U28152 (N_28152,N_22799,N_18518);
or U28153 (N_28153,N_22893,N_19118);
nand U28154 (N_28154,N_23037,N_21765);
and U28155 (N_28155,N_19567,N_23456);
xnor U28156 (N_28156,N_23683,N_20962);
xnor U28157 (N_28157,N_22552,N_18662);
xnor U28158 (N_28158,N_23330,N_20904);
and U28159 (N_28159,N_18058,N_21187);
and U28160 (N_28160,N_21165,N_21990);
xnor U28161 (N_28161,N_21035,N_23990);
nand U28162 (N_28162,N_18270,N_21311);
or U28163 (N_28163,N_21133,N_18140);
and U28164 (N_28164,N_22531,N_19587);
xor U28165 (N_28165,N_23238,N_21266);
or U28166 (N_28166,N_20052,N_22336);
xor U28167 (N_28167,N_23184,N_22323);
nor U28168 (N_28168,N_18272,N_18964);
nand U28169 (N_28169,N_23401,N_19520);
nand U28170 (N_28170,N_23418,N_23479);
nand U28171 (N_28171,N_20588,N_18292);
nor U28172 (N_28172,N_22942,N_19885);
or U28173 (N_28173,N_21093,N_20151);
nor U28174 (N_28174,N_20918,N_22310);
nor U28175 (N_28175,N_18744,N_18691);
xor U28176 (N_28176,N_21114,N_18200);
nand U28177 (N_28177,N_23534,N_21135);
or U28178 (N_28178,N_18623,N_22421);
nand U28179 (N_28179,N_22744,N_23900);
or U28180 (N_28180,N_18081,N_20935);
xnor U28181 (N_28181,N_22781,N_23694);
nor U28182 (N_28182,N_18775,N_20102);
nor U28183 (N_28183,N_19008,N_19807);
and U28184 (N_28184,N_21514,N_18160);
or U28185 (N_28185,N_21177,N_22176);
xnor U28186 (N_28186,N_23255,N_18874);
or U28187 (N_28187,N_23444,N_23220);
xnor U28188 (N_28188,N_19054,N_20043);
or U28189 (N_28189,N_20779,N_20736);
nor U28190 (N_28190,N_20597,N_20664);
xnor U28191 (N_28191,N_19154,N_20930);
or U28192 (N_28192,N_19058,N_18830);
nand U28193 (N_28193,N_19071,N_22662);
nor U28194 (N_28194,N_20502,N_21122);
and U28195 (N_28195,N_19576,N_22202);
xnor U28196 (N_28196,N_20655,N_21023);
nor U28197 (N_28197,N_19092,N_21932);
nand U28198 (N_28198,N_20684,N_21662);
and U28199 (N_28199,N_23332,N_18748);
or U28200 (N_28200,N_20532,N_20912);
nor U28201 (N_28201,N_20098,N_19504);
nor U28202 (N_28202,N_20579,N_21218);
xnor U28203 (N_28203,N_22647,N_18745);
and U28204 (N_28204,N_21934,N_18119);
nand U28205 (N_28205,N_18748,N_21626);
nand U28206 (N_28206,N_23367,N_20285);
xor U28207 (N_28207,N_20292,N_23717);
or U28208 (N_28208,N_23591,N_22116);
xor U28209 (N_28209,N_22187,N_19668);
and U28210 (N_28210,N_20955,N_23926);
and U28211 (N_28211,N_20570,N_20706);
nand U28212 (N_28212,N_20238,N_21629);
or U28213 (N_28213,N_23633,N_23786);
xnor U28214 (N_28214,N_22334,N_22795);
or U28215 (N_28215,N_19487,N_19779);
and U28216 (N_28216,N_21867,N_22293);
nor U28217 (N_28217,N_18314,N_22271);
or U28218 (N_28218,N_21712,N_23867);
nor U28219 (N_28219,N_21743,N_21555);
nor U28220 (N_28220,N_20373,N_21610);
and U28221 (N_28221,N_20016,N_22412);
and U28222 (N_28222,N_21598,N_22341);
or U28223 (N_28223,N_19189,N_20427);
or U28224 (N_28224,N_20401,N_20977);
nand U28225 (N_28225,N_22752,N_21988);
or U28226 (N_28226,N_20616,N_22387);
nor U28227 (N_28227,N_21828,N_23172);
and U28228 (N_28228,N_20728,N_21272);
and U28229 (N_28229,N_19830,N_21029);
or U28230 (N_28230,N_21972,N_23630);
nor U28231 (N_28231,N_23085,N_23691);
and U28232 (N_28232,N_21432,N_19106);
xor U28233 (N_28233,N_18133,N_23407);
xor U28234 (N_28234,N_21106,N_22418);
xnor U28235 (N_28235,N_23398,N_21087);
or U28236 (N_28236,N_21158,N_21849);
xnor U28237 (N_28237,N_22154,N_23698);
nor U28238 (N_28238,N_22064,N_18752);
nor U28239 (N_28239,N_23634,N_21965);
nor U28240 (N_28240,N_18263,N_23277);
and U28241 (N_28241,N_20726,N_20243);
nand U28242 (N_28242,N_22251,N_20766);
xnor U28243 (N_28243,N_20191,N_23854);
xor U28244 (N_28244,N_22476,N_20765);
nor U28245 (N_28245,N_18692,N_21555);
or U28246 (N_28246,N_21614,N_18345);
nor U28247 (N_28247,N_18953,N_20333);
or U28248 (N_28248,N_23951,N_21965);
or U28249 (N_28249,N_19531,N_23042);
and U28250 (N_28250,N_19753,N_18512);
xor U28251 (N_28251,N_21535,N_22633);
or U28252 (N_28252,N_23634,N_22584);
nor U28253 (N_28253,N_19614,N_22611);
xnor U28254 (N_28254,N_20496,N_20485);
or U28255 (N_28255,N_20208,N_22049);
xnor U28256 (N_28256,N_19854,N_22068);
xnor U28257 (N_28257,N_21623,N_18708);
nand U28258 (N_28258,N_20181,N_19795);
xor U28259 (N_28259,N_19989,N_21847);
and U28260 (N_28260,N_23471,N_19963);
or U28261 (N_28261,N_21270,N_19621);
or U28262 (N_28262,N_21794,N_23490);
nor U28263 (N_28263,N_19469,N_19474);
xor U28264 (N_28264,N_18779,N_19376);
nand U28265 (N_28265,N_20729,N_18442);
and U28266 (N_28266,N_23349,N_22052);
or U28267 (N_28267,N_23073,N_23573);
nand U28268 (N_28268,N_21807,N_20365);
nor U28269 (N_28269,N_22870,N_21202);
or U28270 (N_28270,N_21911,N_18958);
nand U28271 (N_28271,N_21343,N_18478);
xor U28272 (N_28272,N_20431,N_18435);
nand U28273 (N_28273,N_20495,N_22055);
or U28274 (N_28274,N_20837,N_23895);
and U28275 (N_28275,N_23166,N_23664);
nand U28276 (N_28276,N_21583,N_19195);
and U28277 (N_28277,N_23424,N_22968);
nand U28278 (N_28278,N_20134,N_19024);
nor U28279 (N_28279,N_19288,N_18487);
or U28280 (N_28280,N_21908,N_23539);
xnor U28281 (N_28281,N_22266,N_20156);
and U28282 (N_28282,N_23278,N_21298);
nand U28283 (N_28283,N_23220,N_19684);
nand U28284 (N_28284,N_22651,N_22165);
xor U28285 (N_28285,N_22180,N_18576);
and U28286 (N_28286,N_22499,N_21844);
nor U28287 (N_28287,N_18861,N_18443);
nand U28288 (N_28288,N_18938,N_22840);
or U28289 (N_28289,N_20253,N_20373);
nand U28290 (N_28290,N_22498,N_22435);
and U28291 (N_28291,N_20999,N_21205);
nand U28292 (N_28292,N_19617,N_21450);
nor U28293 (N_28293,N_23472,N_21931);
xor U28294 (N_28294,N_20534,N_20796);
xnor U28295 (N_28295,N_23916,N_20040);
and U28296 (N_28296,N_19208,N_23465);
nand U28297 (N_28297,N_20967,N_21240);
or U28298 (N_28298,N_21203,N_22099);
nor U28299 (N_28299,N_19740,N_22429);
xor U28300 (N_28300,N_21529,N_23748);
and U28301 (N_28301,N_20820,N_19653);
nand U28302 (N_28302,N_18466,N_22878);
nor U28303 (N_28303,N_20713,N_19758);
xor U28304 (N_28304,N_23639,N_23743);
and U28305 (N_28305,N_22398,N_22728);
or U28306 (N_28306,N_19265,N_20634);
xnor U28307 (N_28307,N_22253,N_21655);
and U28308 (N_28308,N_19718,N_21179);
or U28309 (N_28309,N_22350,N_19996);
nand U28310 (N_28310,N_21274,N_18592);
and U28311 (N_28311,N_21496,N_19621);
and U28312 (N_28312,N_21790,N_22843);
or U28313 (N_28313,N_22617,N_20724);
nor U28314 (N_28314,N_22552,N_19856);
xnor U28315 (N_28315,N_19673,N_18488);
xor U28316 (N_28316,N_23001,N_19874);
and U28317 (N_28317,N_21599,N_20259);
nand U28318 (N_28318,N_20860,N_22925);
xnor U28319 (N_28319,N_22815,N_22760);
or U28320 (N_28320,N_18978,N_18941);
xor U28321 (N_28321,N_18998,N_18067);
and U28322 (N_28322,N_19469,N_21808);
nand U28323 (N_28323,N_19667,N_21319);
xnor U28324 (N_28324,N_20721,N_21513);
or U28325 (N_28325,N_20909,N_20594);
nand U28326 (N_28326,N_18601,N_21000);
and U28327 (N_28327,N_23557,N_19941);
nand U28328 (N_28328,N_19822,N_18472);
and U28329 (N_28329,N_22604,N_21202);
nor U28330 (N_28330,N_19373,N_21468);
or U28331 (N_28331,N_22233,N_21173);
and U28332 (N_28332,N_18066,N_22789);
nor U28333 (N_28333,N_22816,N_19488);
nand U28334 (N_28334,N_18950,N_21832);
xnor U28335 (N_28335,N_20530,N_22247);
nand U28336 (N_28336,N_22158,N_19622);
nand U28337 (N_28337,N_22409,N_22796);
or U28338 (N_28338,N_21241,N_20825);
or U28339 (N_28339,N_21970,N_18038);
nand U28340 (N_28340,N_18306,N_18603);
xor U28341 (N_28341,N_21116,N_20806);
and U28342 (N_28342,N_22700,N_18025);
nor U28343 (N_28343,N_22589,N_23806);
and U28344 (N_28344,N_19295,N_19907);
nor U28345 (N_28345,N_20088,N_18632);
nand U28346 (N_28346,N_19196,N_19953);
or U28347 (N_28347,N_22751,N_20177);
or U28348 (N_28348,N_19294,N_21834);
nor U28349 (N_28349,N_23341,N_23217);
and U28350 (N_28350,N_23131,N_21029);
or U28351 (N_28351,N_20152,N_23555);
nor U28352 (N_28352,N_23223,N_19068);
or U28353 (N_28353,N_21035,N_20532);
nor U28354 (N_28354,N_19668,N_22551);
and U28355 (N_28355,N_19619,N_20760);
or U28356 (N_28356,N_18930,N_23645);
xnor U28357 (N_28357,N_18369,N_18623);
or U28358 (N_28358,N_20903,N_23292);
or U28359 (N_28359,N_20927,N_18084);
or U28360 (N_28360,N_23138,N_21742);
and U28361 (N_28361,N_23152,N_22670);
nand U28362 (N_28362,N_23922,N_23883);
or U28363 (N_28363,N_21758,N_23996);
or U28364 (N_28364,N_21564,N_19453);
nor U28365 (N_28365,N_20637,N_18924);
xnor U28366 (N_28366,N_19398,N_21272);
nand U28367 (N_28367,N_18815,N_21498);
nor U28368 (N_28368,N_22028,N_21566);
nand U28369 (N_28369,N_20854,N_18662);
nand U28370 (N_28370,N_22285,N_23647);
xnor U28371 (N_28371,N_22244,N_22643);
and U28372 (N_28372,N_21815,N_21261);
xnor U28373 (N_28373,N_22315,N_19730);
xnor U28374 (N_28374,N_19804,N_21452);
nand U28375 (N_28375,N_20541,N_22459);
nor U28376 (N_28376,N_18485,N_23218);
xor U28377 (N_28377,N_22371,N_18028);
nand U28378 (N_28378,N_22168,N_21531);
nor U28379 (N_28379,N_21057,N_20299);
nand U28380 (N_28380,N_21842,N_20264);
nand U28381 (N_28381,N_22944,N_19208);
and U28382 (N_28382,N_18382,N_19384);
xor U28383 (N_28383,N_21473,N_19631);
and U28384 (N_28384,N_22917,N_20824);
xnor U28385 (N_28385,N_23311,N_19014);
nand U28386 (N_28386,N_23435,N_22211);
nand U28387 (N_28387,N_22706,N_19419);
and U28388 (N_28388,N_19642,N_18486);
or U28389 (N_28389,N_19878,N_20814);
nand U28390 (N_28390,N_23786,N_21746);
or U28391 (N_28391,N_21581,N_20033);
xnor U28392 (N_28392,N_23211,N_23614);
nor U28393 (N_28393,N_20972,N_23180);
xnor U28394 (N_28394,N_18308,N_23191);
nor U28395 (N_28395,N_20496,N_18245);
nand U28396 (N_28396,N_22909,N_18659);
or U28397 (N_28397,N_23613,N_22966);
and U28398 (N_28398,N_23653,N_22977);
nand U28399 (N_28399,N_21182,N_22032);
nand U28400 (N_28400,N_20680,N_22501);
or U28401 (N_28401,N_19734,N_19544);
xnor U28402 (N_28402,N_21360,N_22986);
nor U28403 (N_28403,N_23864,N_23459);
xor U28404 (N_28404,N_18764,N_19406);
nor U28405 (N_28405,N_19539,N_18283);
and U28406 (N_28406,N_22479,N_18733);
or U28407 (N_28407,N_18811,N_20927);
and U28408 (N_28408,N_18856,N_20484);
nor U28409 (N_28409,N_23671,N_20897);
and U28410 (N_28410,N_20856,N_20336);
xnor U28411 (N_28411,N_23381,N_19320);
or U28412 (N_28412,N_22427,N_23188);
or U28413 (N_28413,N_20213,N_20493);
nor U28414 (N_28414,N_18922,N_21846);
and U28415 (N_28415,N_20564,N_21180);
or U28416 (N_28416,N_18378,N_23369);
nor U28417 (N_28417,N_19536,N_21846);
nor U28418 (N_28418,N_22116,N_21736);
nor U28419 (N_28419,N_22828,N_22127);
and U28420 (N_28420,N_19975,N_20189);
nor U28421 (N_28421,N_19432,N_19890);
xor U28422 (N_28422,N_23842,N_19005);
nor U28423 (N_28423,N_21103,N_19984);
or U28424 (N_28424,N_20933,N_18375);
nor U28425 (N_28425,N_21171,N_19207);
xor U28426 (N_28426,N_22491,N_21390);
or U28427 (N_28427,N_18043,N_21353);
or U28428 (N_28428,N_23429,N_19952);
or U28429 (N_28429,N_21982,N_18133);
and U28430 (N_28430,N_18023,N_18367);
or U28431 (N_28431,N_23299,N_19831);
nor U28432 (N_28432,N_20660,N_23038);
nand U28433 (N_28433,N_20029,N_20885);
nor U28434 (N_28434,N_20056,N_22553);
or U28435 (N_28435,N_18434,N_18100);
xnor U28436 (N_28436,N_23968,N_20099);
and U28437 (N_28437,N_21484,N_19368);
xor U28438 (N_28438,N_23181,N_23889);
nand U28439 (N_28439,N_23916,N_20613);
xnor U28440 (N_28440,N_19443,N_23253);
nor U28441 (N_28441,N_18122,N_23440);
or U28442 (N_28442,N_21910,N_22939);
or U28443 (N_28443,N_19842,N_21636);
nor U28444 (N_28444,N_20078,N_20196);
xnor U28445 (N_28445,N_19146,N_21512);
nor U28446 (N_28446,N_22122,N_19257);
or U28447 (N_28447,N_22938,N_18459);
nor U28448 (N_28448,N_18415,N_23048);
nand U28449 (N_28449,N_21060,N_18442);
and U28450 (N_28450,N_19536,N_21464);
nor U28451 (N_28451,N_23726,N_23441);
nor U28452 (N_28452,N_22267,N_18735);
nor U28453 (N_28453,N_20915,N_20745);
or U28454 (N_28454,N_23843,N_22371);
nor U28455 (N_28455,N_20975,N_18178);
nor U28456 (N_28456,N_22657,N_23844);
nor U28457 (N_28457,N_19996,N_22155);
and U28458 (N_28458,N_21035,N_19697);
xnor U28459 (N_28459,N_22586,N_22244);
nand U28460 (N_28460,N_18805,N_18915);
nor U28461 (N_28461,N_22165,N_18174);
and U28462 (N_28462,N_22204,N_18922);
and U28463 (N_28463,N_18717,N_18461);
and U28464 (N_28464,N_21556,N_20454);
or U28465 (N_28465,N_20195,N_19548);
and U28466 (N_28466,N_20272,N_22040);
or U28467 (N_28467,N_22894,N_21874);
and U28468 (N_28468,N_21717,N_23953);
xnor U28469 (N_28469,N_18736,N_23496);
xor U28470 (N_28470,N_20541,N_18937);
and U28471 (N_28471,N_18495,N_21704);
or U28472 (N_28472,N_20979,N_21421);
xnor U28473 (N_28473,N_18625,N_19797);
nor U28474 (N_28474,N_19834,N_19201);
or U28475 (N_28475,N_20384,N_23970);
nor U28476 (N_28476,N_23959,N_23174);
or U28477 (N_28477,N_22251,N_21149);
xor U28478 (N_28478,N_23611,N_20852);
and U28479 (N_28479,N_20988,N_22697);
or U28480 (N_28480,N_18507,N_23330);
or U28481 (N_28481,N_22632,N_21587);
nand U28482 (N_28482,N_22077,N_21759);
or U28483 (N_28483,N_19930,N_20078);
and U28484 (N_28484,N_21061,N_19854);
or U28485 (N_28485,N_18462,N_21491);
nor U28486 (N_28486,N_21528,N_22583);
or U28487 (N_28487,N_22890,N_20178);
nor U28488 (N_28488,N_22086,N_20169);
and U28489 (N_28489,N_19211,N_19578);
or U28490 (N_28490,N_20344,N_23511);
nor U28491 (N_28491,N_22018,N_20622);
xnor U28492 (N_28492,N_18482,N_23971);
and U28493 (N_28493,N_18493,N_19192);
or U28494 (N_28494,N_22099,N_21622);
and U28495 (N_28495,N_18970,N_22768);
xnor U28496 (N_28496,N_21033,N_18348);
and U28497 (N_28497,N_20000,N_19460);
and U28498 (N_28498,N_21667,N_19431);
xnor U28499 (N_28499,N_19244,N_20444);
or U28500 (N_28500,N_23230,N_21328);
or U28501 (N_28501,N_19217,N_23335);
xnor U28502 (N_28502,N_19810,N_22073);
nor U28503 (N_28503,N_23727,N_19569);
and U28504 (N_28504,N_21962,N_22176);
nand U28505 (N_28505,N_23847,N_22415);
and U28506 (N_28506,N_21985,N_21051);
xnor U28507 (N_28507,N_18030,N_21286);
nand U28508 (N_28508,N_22049,N_20698);
nand U28509 (N_28509,N_22725,N_19591);
or U28510 (N_28510,N_20587,N_20781);
xor U28511 (N_28511,N_22521,N_22626);
nor U28512 (N_28512,N_18934,N_20684);
or U28513 (N_28513,N_19577,N_23281);
nor U28514 (N_28514,N_20685,N_20506);
or U28515 (N_28515,N_21984,N_22940);
xnor U28516 (N_28516,N_23937,N_20420);
and U28517 (N_28517,N_20616,N_22934);
or U28518 (N_28518,N_18550,N_22362);
xor U28519 (N_28519,N_20502,N_19396);
and U28520 (N_28520,N_18542,N_23315);
and U28521 (N_28521,N_19973,N_23416);
xor U28522 (N_28522,N_23070,N_20108);
nor U28523 (N_28523,N_20536,N_23059);
xnor U28524 (N_28524,N_18786,N_23071);
and U28525 (N_28525,N_22989,N_18143);
nor U28526 (N_28526,N_20529,N_19539);
or U28527 (N_28527,N_19623,N_23789);
or U28528 (N_28528,N_23074,N_19991);
xnor U28529 (N_28529,N_20441,N_19104);
and U28530 (N_28530,N_21989,N_22410);
nand U28531 (N_28531,N_23385,N_23265);
nor U28532 (N_28532,N_21004,N_19133);
nor U28533 (N_28533,N_22245,N_23993);
and U28534 (N_28534,N_21036,N_21538);
nor U28535 (N_28535,N_21982,N_20708);
or U28536 (N_28536,N_23417,N_21182);
and U28537 (N_28537,N_23808,N_21661);
and U28538 (N_28538,N_20319,N_23175);
or U28539 (N_28539,N_21043,N_18977);
or U28540 (N_28540,N_21003,N_20434);
nor U28541 (N_28541,N_18306,N_21364);
or U28542 (N_28542,N_23298,N_23517);
or U28543 (N_28543,N_23058,N_21805);
xnor U28544 (N_28544,N_21850,N_20352);
or U28545 (N_28545,N_23582,N_18716);
or U28546 (N_28546,N_18233,N_20929);
xor U28547 (N_28547,N_22199,N_23557);
and U28548 (N_28548,N_21001,N_19362);
and U28549 (N_28549,N_22926,N_18669);
and U28550 (N_28550,N_22808,N_21503);
xor U28551 (N_28551,N_21089,N_19220);
nor U28552 (N_28552,N_22208,N_18404);
xor U28553 (N_28553,N_21990,N_22613);
xnor U28554 (N_28554,N_22752,N_18813);
nor U28555 (N_28555,N_19331,N_19734);
xnor U28556 (N_28556,N_23063,N_20777);
xnor U28557 (N_28557,N_22173,N_18069);
nor U28558 (N_28558,N_18914,N_21391);
nor U28559 (N_28559,N_22589,N_18393);
or U28560 (N_28560,N_23401,N_18703);
nand U28561 (N_28561,N_21663,N_20674);
and U28562 (N_28562,N_22529,N_22590);
or U28563 (N_28563,N_20589,N_19203);
or U28564 (N_28564,N_21785,N_18819);
nor U28565 (N_28565,N_23161,N_18717);
nor U28566 (N_28566,N_21259,N_23672);
xor U28567 (N_28567,N_20029,N_22368);
and U28568 (N_28568,N_19812,N_20580);
nand U28569 (N_28569,N_20505,N_20287);
and U28570 (N_28570,N_19440,N_18971);
and U28571 (N_28571,N_19427,N_21869);
nand U28572 (N_28572,N_23869,N_20635);
nor U28573 (N_28573,N_22755,N_22563);
or U28574 (N_28574,N_22039,N_23655);
and U28575 (N_28575,N_19175,N_18849);
nor U28576 (N_28576,N_20319,N_23779);
nor U28577 (N_28577,N_23747,N_23435);
xor U28578 (N_28578,N_18157,N_23010);
or U28579 (N_28579,N_20886,N_23164);
xor U28580 (N_28580,N_23030,N_18092);
or U28581 (N_28581,N_18910,N_19064);
and U28582 (N_28582,N_21761,N_19373);
and U28583 (N_28583,N_21783,N_22092);
and U28584 (N_28584,N_20002,N_18991);
xor U28585 (N_28585,N_23323,N_20390);
and U28586 (N_28586,N_20394,N_18652);
xor U28587 (N_28587,N_21961,N_18872);
nand U28588 (N_28588,N_19145,N_20494);
or U28589 (N_28589,N_19875,N_20845);
or U28590 (N_28590,N_23664,N_22185);
nor U28591 (N_28591,N_20565,N_18676);
and U28592 (N_28592,N_21727,N_18011);
xnor U28593 (N_28593,N_22448,N_22740);
and U28594 (N_28594,N_18209,N_21750);
nor U28595 (N_28595,N_23495,N_22966);
xnor U28596 (N_28596,N_23084,N_22183);
and U28597 (N_28597,N_18607,N_19957);
xnor U28598 (N_28598,N_19212,N_20784);
xnor U28599 (N_28599,N_20747,N_23895);
nor U28600 (N_28600,N_23400,N_23915);
xor U28601 (N_28601,N_20270,N_18665);
xnor U28602 (N_28602,N_23348,N_22503);
and U28603 (N_28603,N_20221,N_22807);
xor U28604 (N_28604,N_18311,N_21508);
nand U28605 (N_28605,N_23048,N_21649);
nand U28606 (N_28606,N_22038,N_18494);
xor U28607 (N_28607,N_23211,N_18876);
nand U28608 (N_28608,N_18241,N_18253);
and U28609 (N_28609,N_21646,N_22018);
xor U28610 (N_28610,N_19095,N_19976);
xnor U28611 (N_28611,N_23860,N_20786);
nor U28612 (N_28612,N_22846,N_20382);
nor U28613 (N_28613,N_23991,N_19479);
xor U28614 (N_28614,N_21436,N_22833);
nand U28615 (N_28615,N_18536,N_21481);
nor U28616 (N_28616,N_23210,N_22520);
nand U28617 (N_28617,N_18098,N_19736);
nor U28618 (N_28618,N_21251,N_20215);
and U28619 (N_28619,N_19642,N_21232);
or U28620 (N_28620,N_22135,N_19808);
nor U28621 (N_28621,N_22550,N_23561);
nand U28622 (N_28622,N_23303,N_19258);
or U28623 (N_28623,N_22113,N_18729);
xor U28624 (N_28624,N_22334,N_18103);
xnor U28625 (N_28625,N_18284,N_21750);
and U28626 (N_28626,N_23241,N_21780);
xor U28627 (N_28627,N_18598,N_21243);
or U28628 (N_28628,N_20265,N_22901);
nor U28629 (N_28629,N_19261,N_23046);
xor U28630 (N_28630,N_19309,N_22949);
or U28631 (N_28631,N_22830,N_22359);
nor U28632 (N_28632,N_18694,N_19172);
or U28633 (N_28633,N_18292,N_20479);
or U28634 (N_28634,N_21555,N_22796);
nand U28635 (N_28635,N_21924,N_22657);
or U28636 (N_28636,N_18732,N_23782);
and U28637 (N_28637,N_18445,N_19513);
and U28638 (N_28638,N_21286,N_22228);
xnor U28639 (N_28639,N_20409,N_19025);
or U28640 (N_28640,N_18567,N_20096);
nor U28641 (N_28641,N_21071,N_22553);
nor U28642 (N_28642,N_21514,N_20151);
xor U28643 (N_28643,N_22337,N_22667);
xnor U28644 (N_28644,N_20750,N_22780);
nand U28645 (N_28645,N_19897,N_21303);
nor U28646 (N_28646,N_23225,N_21481);
or U28647 (N_28647,N_22127,N_22345);
or U28648 (N_28648,N_19409,N_20807);
or U28649 (N_28649,N_20824,N_19813);
nor U28650 (N_28650,N_19127,N_19042);
nand U28651 (N_28651,N_22184,N_18184);
xor U28652 (N_28652,N_19701,N_20152);
xnor U28653 (N_28653,N_20053,N_20154);
or U28654 (N_28654,N_23883,N_23034);
or U28655 (N_28655,N_19228,N_20369);
nor U28656 (N_28656,N_22915,N_18828);
nand U28657 (N_28657,N_19160,N_23726);
nor U28658 (N_28658,N_19947,N_23530);
xor U28659 (N_28659,N_21663,N_22107);
and U28660 (N_28660,N_21851,N_20880);
and U28661 (N_28661,N_21258,N_19863);
nor U28662 (N_28662,N_19590,N_23030);
nor U28663 (N_28663,N_21183,N_18240);
xnor U28664 (N_28664,N_21367,N_23576);
or U28665 (N_28665,N_19576,N_23270);
and U28666 (N_28666,N_20204,N_18223);
nor U28667 (N_28667,N_20952,N_19875);
nand U28668 (N_28668,N_22532,N_22457);
xnor U28669 (N_28669,N_19868,N_22620);
or U28670 (N_28670,N_18948,N_19673);
nand U28671 (N_28671,N_19985,N_23391);
xnor U28672 (N_28672,N_21898,N_19384);
nand U28673 (N_28673,N_20725,N_18868);
xnor U28674 (N_28674,N_22129,N_22901);
xor U28675 (N_28675,N_21525,N_19974);
nor U28676 (N_28676,N_21224,N_18754);
nand U28677 (N_28677,N_23958,N_19627);
nand U28678 (N_28678,N_19807,N_19994);
or U28679 (N_28679,N_21975,N_22311);
nor U28680 (N_28680,N_22175,N_20161);
xor U28681 (N_28681,N_20459,N_20316);
nor U28682 (N_28682,N_22843,N_20648);
nand U28683 (N_28683,N_20827,N_19697);
nor U28684 (N_28684,N_23455,N_21348);
or U28685 (N_28685,N_19542,N_23839);
or U28686 (N_28686,N_23951,N_19579);
nand U28687 (N_28687,N_19343,N_22278);
xnor U28688 (N_28688,N_21548,N_20590);
nor U28689 (N_28689,N_21414,N_21123);
nand U28690 (N_28690,N_23714,N_23718);
xnor U28691 (N_28691,N_21193,N_22441);
and U28692 (N_28692,N_23514,N_19067);
nor U28693 (N_28693,N_23636,N_19329);
nand U28694 (N_28694,N_23225,N_18299);
or U28695 (N_28695,N_20191,N_19134);
or U28696 (N_28696,N_22690,N_23524);
nand U28697 (N_28697,N_23147,N_23164);
nor U28698 (N_28698,N_20875,N_21888);
and U28699 (N_28699,N_19064,N_18725);
xor U28700 (N_28700,N_21210,N_21325);
or U28701 (N_28701,N_22295,N_18036);
or U28702 (N_28702,N_19894,N_23873);
xor U28703 (N_28703,N_19601,N_22181);
or U28704 (N_28704,N_20559,N_18714);
xnor U28705 (N_28705,N_22609,N_20172);
or U28706 (N_28706,N_23426,N_23483);
xnor U28707 (N_28707,N_19322,N_21848);
xnor U28708 (N_28708,N_21275,N_20844);
and U28709 (N_28709,N_18474,N_20339);
xnor U28710 (N_28710,N_18454,N_21601);
nand U28711 (N_28711,N_19546,N_21984);
xor U28712 (N_28712,N_23733,N_19436);
and U28713 (N_28713,N_18096,N_19319);
and U28714 (N_28714,N_18742,N_21792);
and U28715 (N_28715,N_18421,N_20702);
or U28716 (N_28716,N_21499,N_23444);
nand U28717 (N_28717,N_21873,N_20423);
nor U28718 (N_28718,N_18397,N_18145);
or U28719 (N_28719,N_23160,N_18128);
and U28720 (N_28720,N_23113,N_22211);
nor U28721 (N_28721,N_22346,N_23196);
nand U28722 (N_28722,N_18736,N_23721);
xor U28723 (N_28723,N_19383,N_18027);
nor U28724 (N_28724,N_20965,N_20738);
and U28725 (N_28725,N_19055,N_22934);
nand U28726 (N_28726,N_23649,N_22024);
and U28727 (N_28727,N_23665,N_19479);
nand U28728 (N_28728,N_22249,N_20137);
nor U28729 (N_28729,N_23441,N_23584);
nand U28730 (N_28730,N_22835,N_18866);
or U28731 (N_28731,N_20317,N_20625);
or U28732 (N_28732,N_20942,N_23012);
xnor U28733 (N_28733,N_18034,N_23690);
and U28734 (N_28734,N_20237,N_21932);
nor U28735 (N_28735,N_21584,N_23081);
or U28736 (N_28736,N_22610,N_23643);
and U28737 (N_28737,N_18037,N_21565);
and U28738 (N_28738,N_20958,N_23608);
nor U28739 (N_28739,N_21966,N_21479);
and U28740 (N_28740,N_19807,N_18002);
and U28741 (N_28741,N_19531,N_22565);
or U28742 (N_28742,N_23591,N_22495);
or U28743 (N_28743,N_18175,N_23541);
nand U28744 (N_28744,N_23522,N_18378);
or U28745 (N_28745,N_22127,N_19614);
or U28746 (N_28746,N_19062,N_22800);
and U28747 (N_28747,N_18453,N_23837);
nor U28748 (N_28748,N_18905,N_18366);
nand U28749 (N_28749,N_18353,N_22338);
xor U28750 (N_28750,N_21413,N_19276);
nor U28751 (N_28751,N_20181,N_18973);
or U28752 (N_28752,N_20966,N_19222);
or U28753 (N_28753,N_20565,N_21235);
and U28754 (N_28754,N_22850,N_21773);
and U28755 (N_28755,N_20039,N_18313);
or U28756 (N_28756,N_20511,N_19442);
and U28757 (N_28757,N_23456,N_21513);
nand U28758 (N_28758,N_22826,N_20055);
nor U28759 (N_28759,N_18584,N_23048);
xnor U28760 (N_28760,N_23349,N_22702);
xnor U28761 (N_28761,N_20921,N_20619);
nand U28762 (N_28762,N_23246,N_19769);
and U28763 (N_28763,N_20793,N_20582);
nand U28764 (N_28764,N_18111,N_18363);
xnor U28765 (N_28765,N_21330,N_21415);
or U28766 (N_28766,N_18398,N_20887);
nor U28767 (N_28767,N_18876,N_22935);
nand U28768 (N_28768,N_20916,N_21319);
or U28769 (N_28769,N_20692,N_23714);
xor U28770 (N_28770,N_22477,N_22716);
and U28771 (N_28771,N_20103,N_23093);
and U28772 (N_28772,N_21358,N_20112);
or U28773 (N_28773,N_21752,N_21763);
xor U28774 (N_28774,N_22989,N_21639);
or U28775 (N_28775,N_18116,N_19628);
nand U28776 (N_28776,N_20870,N_23321);
xnor U28777 (N_28777,N_22058,N_19681);
xnor U28778 (N_28778,N_22382,N_20071);
nand U28779 (N_28779,N_18500,N_23602);
xor U28780 (N_28780,N_21298,N_19515);
xnor U28781 (N_28781,N_19531,N_20941);
or U28782 (N_28782,N_23965,N_20692);
or U28783 (N_28783,N_21365,N_20236);
nand U28784 (N_28784,N_19065,N_19288);
nor U28785 (N_28785,N_18736,N_20546);
or U28786 (N_28786,N_20609,N_23476);
nor U28787 (N_28787,N_21845,N_21834);
and U28788 (N_28788,N_23412,N_21642);
nand U28789 (N_28789,N_19739,N_18964);
nor U28790 (N_28790,N_19213,N_22872);
nor U28791 (N_28791,N_23687,N_22775);
and U28792 (N_28792,N_21536,N_19521);
xnor U28793 (N_28793,N_22749,N_23416);
nor U28794 (N_28794,N_19705,N_23559);
and U28795 (N_28795,N_20741,N_20776);
xnor U28796 (N_28796,N_22111,N_23995);
nand U28797 (N_28797,N_18898,N_18297);
nor U28798 (N_28798,N_20742,N_22293);
nor U28799 (N_28799,N_22357,N_19500);
and U28800 (N_28800,N_19854,N_18887);
or U28801 (N_28801,N_23161,N_21729);
nand U28802 (N_28802,N_21413,N_18207);
nor U28803 (N_28803,N_20793,N_22672);
nor U28804 (N_28804,N_21551,N_23062);
or U28805 (N_28805,N_20564,N_18185);
or U28806 (N_28806,N_18843,N_23829);
or U28807 (N_28807,N_22836,N_20382);
or U28808 (N_28808,N_19176,N_18081);
and U28809 (N_28809,N_20075,N_20043);
nand U28810 (N_28810,N_22305,N_18152);
or U28811 (N_28811,N_21863,N_23858);
or U28812 (N_28812,N_19343,N_21690);
nor U28813 (N_28813,N_18311,N_19006);
or U28814 (N_28814,N_21614,N_18697);
or U28815 (N_28815,N_22620,N_22065);
or U28816 (N_28816,N_20931,N_23478);
or U28817 (N_28817,N_23011,N_20236);
nor U28818 (N_28818,N_22784,N_20847);
and U28819 (N_28819,N_21447,N_18497);
and U28820 (N_28820,N_22867,N_18991);
xor U28821 (N_28821,N_22313,N_19212);
xnor U28822 (N_28822,N_21326,N_18684);
or U28823 (N_28823,N_20048,N_21162);
nor U28824 (N_28824,N_22792,N_18099);
or U28825 (N_28825,N_19317,N_23842);
xor U28826 (N_28826,N_21861,N_20376);
xor U28827 (N_28827,N_20238,N_19038);
nor U28828 (N_28828,N_18955,N_23275);
xor U28829 (N_28829,N_22685,N_22912);
nand U28830 (N_28830,N_23306,N_18627);
and U28831 (N_28831,N_19805,N_18828);
nand U28832 (N_28832,N_19963,N_22837);
or U28833 (N_28833,N_21374,N_22307);
nor U28834 (N_28834,N_20310,N_22350);
nand U28835 (N_28835,N_20409,N_21539);
xnor U28836 (N_28836,N_21530,N_18495);
and U28837 (N_28837,N_20799,N_22083);
and U28838 (N_28838,N_21022,N_18235);
xor U28839 (N_28839,N_22571,N_18691);
or U28840 (N_28840,N_23612,N_21221);
or U28841 (N_28841,N_22429,N_22381);
nand U28842 (N_28842,N_19555,N_23878);
nor U28843 (N_28843,N_23774,N_21572);
or U28844 (N_28844,N_19536,N_22733);
xnor U28845 (N_28845,N_21732,N_20639);
xnor U28846 (N_28846,N_19414,N_21335);
and U28847 (N_28847,N_20572,N_22085);
and U28848 (N_28848,N_23553,N_19155);
and U28849 (N_28849,N_23229,N_21748);
nor U28850 (N_28850,N_18121,N_20783);
nand U28851 (N_28851,N_19184,N_23985);
or U28852 (N_28852,N_18297,N_23800);
xor U28853 (N_28853,N_21485,N_19129);
nor U28854 (N_28854,N_18471,N_23848);
xnor U28855 (N_28855,N_21107,N_22147);
nand U28856 (N_28856,N_22686,N_21265);
and U28857 (N_28857,N_20932,N_18785);
nand U28858 (N_28858,N_18331,N_22056);
or U28859 (N_28859,N_22685,N_22059);
nor U28860 (N_28860,N_21302,N_22081);
xnor U28861 (N_28861,N_21443,N_18404);
or U28862 (N_28862,N_23127,N_19500);
xor U28863 (N_28863,N_18188,N_22930);
nand U28864 (N_28864,N_19563,N_22028);
nand U28865 (N_28865,N_23989,N_22703);
nand U28866 (N_28866,N_22351,N_21035);
nor U28867 (N_28867,N_22425,N_18106);
nor U28868 (N_28868,N_19971,N_21040);
nor U28869 (N_28869,N_19156,N_19958);
and U28870 (N_28870,N_23093,N_21492);
and U28871 (N_28871,N_23448,N_18661);
and U28872 (N_28872,N_21872,N_18475);
or U28873 (N_28873,N_18657,N_20633);
or U28874 (N_28874,N_22044,N_21912);
nor U28875 (N_28875,N_23663,N_18562);
xnor U28876 (N_28876,N_20010,N_19508);
nor U28877 (N_28877,N_19434,N_21442);
nor U28878 (N_28878,N_18171,N_18357);
nor U28879 (N_28879,N_21053,N_23431);
nor U28880 (N_28880,N_23670,N_19385);
nand U28881 (N_28881,N_23758,N_22951);
or U28882 (N_28882,N_22522,N_18741);
nor U28883 (N_28883,N_23484,N_20457);
nand U28884 (N_28884,N_21976,N_18182);
nand U28885 (N_28885,N_22940,N_19145);
xnor U28886 (N_28886,N_20926,N_23294);
nand U28887 (N_28887,N_22554,N_18470);
or U28888 (N_28888,N_22952,N_21245);
and U28889 (N_28889,N_22113,N_18768);
nand U28890 (N_28890,N_23100,N_22343);
or U28891 (N_28891,N_21936,N_22298);
or U28892 (N_28892,N_20739,N_22574);
nor U28893 (N_28893,N_21408,N_22029);
nor U28894 (N_28894,N_21695,N_21032);
nor U28895 (N_28895,N_21475,N_20304);
or U28896 (N_28896,N_21947,N_22529);
xor U28897 (N_28897,N_20681,N_19099);
or U28898 (N_28898,N_23357,N_20590);
nand U28899 (N_28899,N_21498,N_23551);
xnor U28900 (N_28900,N_21256,N_19025);
and U28901 (N_28901,N_23545,N_18822);
or U28902 (N_28902,N_18106,N_23342);
nand U28903 (N_28903,N_20166,N_22216);
nand U28904 (N_28904,N_21633,N_20030);
nand U28905 (N_28905,N_21040,N_22506);
nor U28906 (N_28906,N_18479,N_18576);
nor U28907 (N_28907,N_22026,N_21621);
or U28908 (N_28908,N_23325,N_22831);
xnor U28909 (N_28909,N_21532,N_22508);
xnor U28910 (N_28910,N_19491,N_21176);
nand U28911 (N_28911,N_23809,N_22697);
and U28912 (N_28912,N_20763,N_22246);
nor U28913 (N_28913,N_20028,N_23355);
xor U28914 (N_28914,N_23115,N_23967);
and U28915 (N_28915,N_18547,N_23964);
nor U28916 (N_28916,N_21759,N_20567);
xnor U28917 (N_28917,N_21842,N_20290);
nand U28918 (N_28918,N_20862,N_23437);
nand U28919 (N_28919,N_20077,N_20971);
or U28920 (N_28920,N_22146,N_22248);
and U28921 (N_28921,N_18116,N_18362);
or U28922 (N_28922,N_23066,N_22048);
xor U28923 (N_28923,N_18044,N_23316);
xnor U28924 (N_28924,N_23996,N_18559);
nor U28925 (N_28925,N_21793,N_23710);
nor U28926 (N_28926,N_22626,N_20619);
nand U28927 (N_28927,N_23850,N_18210);
xor U28928 (N_28928,N_19095,N_18209);
nor U28929 (N_28929,N_23172,N_18733);
or U28930 (N_28930,N_23472,N_23118);
nor U28931 (N_28931,N_19843,N_21085);
and U28932 (N_28932,N_23609,N_21999);
nor U28933 (N_28933,N_21254,N_20993);
and U28934 (N_28934,N_23831,N_20271);
nor U28935 (N_28935,N_20717,N_22028);
and U28936 (N_28936,N_22301,N_20796);
xnor U28937 (N_28937,N_22823,N_22204);
nor U28938 (N_28938,N_23526,N_19396);
and U28939 (N_28939,N_20206,N_22345);
nand U28940 (N_28940,N_19902,N_22973);
or U28941 (N_28941,N_19567,N_22695);
xor U28942 (N_28942,N_18266,N_18184);
xnor U28943 (N_28943,N_20400,N_22693);
or U28944 (N_28944,N_18059,N_18287);
and U28945 (N_28945,N_20507,N_19709);
or U28946 (N_28946,N_21482,N_19703);
xnor U28947 (N_28947,N_21750,N_19276);
xor U28948 (N_28948,N_19116,N_22217);
xnor U28949 (N_28949,N_18316,N_22855);
nand U28950 (N_28950,N_20663,N_20151);
nand U28951 (N_28951,N_18054,N_22235);
nor U28952 (N_28952,N_21157,N_22996);
xnor U28953 (N_28953,N_23192,N_21083);
nand U28954 (N_28954,N_19739,N_20263);
or U28955 (N_28955,N_21141,N_21006);
or U28956 (N_28956,N_19239,N_21359);
and U28957 (N_28957,N_20350,N_23583);
and U28958 (N_28958,N_18738,N_20574);
and U28959 (N_28959,N_19296,N_19174);
nand U28960 (N_28960,N_23488,N_20745);
nor U28961 (N_28961,N_21462,N_19980);
and U28962 (N_28962,N_21246,N_23707);
nor U28963 (N_28963,N_22340,N_20309);
and U28964 (N_28964,N_22920,N_18788);
nor U28965 (N_28965,N_18950,N_20809);
nor U28966 (N_28966,N_18776,N_22216);
nand U28967 (N_28967,N_21651,N_20616);
and U28968 (N_28968,N_23013,N_19196);
nor U28969 (N_28969,N_22617,N_18462);
and U28970 (N_28970,N_18845,N_19577);
or U28971 (N_28971,N_20980,N_20748);
xnor U28972 (N_28972,N_23593,N_21710);
xnor U28973 (N_28973,N_18000,N_20403);
or U28974 (N_28974,N_23767,N_21295);
nor U28975 (N_28975,N_21500,N_22935);
xnor U28976 (N_28976,N_22473,N_23185);
nand U28977 (N_28977,N_23972,N_21391);
nand U28978 (N_28978,N_23813,N_20715);
nand U28979 (N_28979,N_20183,N_21517);
xor U28980 (N_28980,N_21396,N_21662);
nor U28981 (N_28981,N_18126,N_19593);
xor U28982 (N_28982,N_21633,N_22711);
nor U28983 (N_28983,N_19577,N_19018);
and U28984 (N_28984,N_20283,N_22749);
xor U28985 (N_28985,N_19250,N_21368);
xor U28986 (N_28986,N_22068,N_18535);
or U28987 (N_28987,N_22211,N_23737);
nor U28988 (N_28988,N_20916,N_19409);
xor U28989 (N_28989,N_19249,N_19098);
xnor U28990 (N_28990,N_22099,N_23936);
and U28991 (N_28991,N_23848,N_19572);
nand U28992 (N_28992,N_23120,N_22519);
or U28993 (N_28993,N_22506,N_21089);
and U28994 (N_28994,N_21401,N_19069);
xnor U28995 (N_28995,N_19399,N_21071);
xor U28996 (N_28996,N_21299,N_19143);
xnor U28997 (N_28997,N_23269,N_21484);
nand U28998 (N_28998,N_20214,N_23717);
and U28999 (N_28999,N_23564,N_23434);
or U29000 (N_29000,N_22764,N_19079);
nand U29001 (N_29001,N_20691,N_22468);
and U29002 (N_29002,N_22846,N_20807);
nor U29003 (N_29003,N_22563,N_23838);
nor U29004 (N_29004,N_18172,N_19327);
and U29005 (N_29005,N_20281,N_21626);
xnor U29006 (N_29006,N_20445,N_23772);
nand U29007 (N_29007,N_18103,N_23962);
nand U29008 (N_29008,N_21506,N_18862);
or U29009 (N_29009,N_21026,N_22326);
and U29010 (N_29010,N_22591,N_22433);
and U29011 (N_29011,N_23407,N_20099);
or U29012 (N_29012,N_19090,N_18627);
and U29013 (N_29013,N_23072,N_21685);
xnor U29014 (N_29014,N_21224,N_23678);
xnor U29015 (N_29015,N_23431,N_20473);
nand U29016 (N_29016,N_19982,N_22265);
nand U29017 (N_29017,N_18344,N_21665);
xnor U29018 (N_29018,N_20757,N_19414);
xnor U29019 (N_29019,N_23009,N_21795);
nand U29020 (N_29020,N_19752,N_19205);
nor U29021 (N_29021,N_23190,N_23944);
and U29022 (N_29022,N_20009,N_23374);
nand U29023 (N_29023,N_22192,N_20648);
nand U29024 (N_29024,N_20548,N_18394);
nand U29025 (N_29025,N_22503,N_23054);
nor U29026 (N_29026,N_20043,N_18472);
nand U29027 (N_29027,N_18587,N_19235);
or U29028 (N_29028,N_20011,N_23252);
xnor U29029 (N_29029,N_19444,N_23442);
and U29030 (N_29030,N_18668,N_19093);
nor U29031 (N_29031,N_18751,N_21543);
and U29032 (N_29032,N_19902,N_22516);
nand U29033 (N_29033,N_22581,N_23825);
and U29034 (N_29034,N_18154,N_19163);
nor U29035 (N_29035,N_22698,N_23176);
or U29036 (N_29036,N_18735,N_20511);
or U29037 (N_29037,N_19849,N_18177);
nor U29038 (N_29038,N_22726,N_23749);
and U29039 (N_29039,N_21639,N_22168);
or U29040 (N_29040,N_23865,N_21730);
xor U29041 (N_29041,N_21808,N_18892);
and U29042 (N_29042,N_23561,N_20278);
xor U29043 (N_29043,N_18434,N_20223);
and U29044 (N_29044,N_19155,N_22011);
nand U29045 (N_29045,N_23794,N_20382);
nand U29046 (N_29046,N_22009,N_21572);
nor U29047 (N_29047,N_22003,N_23834);
and U29048 (N_29048,N_22911,N_18697);
xor U29049 (N_29049,N_20301,N_19687);
or U29050 (N_29050,N_20328,N_23599);
nor U29051 (N_29051,N_20695,N_22116);
nor U29052 (N_29052,N_20480,N_22412);
nor U29053 (N_29053,N_20871,N_23633);
nor U29054 (N_29054,N_18086,N_20387);
nand U29055 (N_29055,N_19729,N_18811);
nor U29056 (N_29056,N_18262,N_22540);
and U29057 (N_29057,N_21262,N_22069);
or U29058 (N_29058,N_23247,N_21009);
nor U29059 (N_29059,N_20074,N_19615);
xor U29060 (N_29060,N_21831,N_19582);
nor U29061 (N_29061,N_22597,N_18984);
and U29062 (N_29062,N_20767,N_23408);
and U29063 (N_29063,N_18707,N_19097);
nand U29064 (N_29064,N_22025,N_23117);
xor U29065 (N_29065,N_22788,N_19776);
or U29066 (N_29066,N_20678,N_21964);
nor U29067 (N_29067,N_21077,N_18178);
nand U29068 (N_29068,N_20554,N_21552);
nand U29069 (N_29069,N_21245,N_23117);
nor U29070 (N_29070,N_20541,N_20631);
nand U29071 (N_29071,N_20640,N_23961);
nor U29072 (N_29072,N_21545,N_19087);
nand U29073 (N_29073,N_22283,N_18775);
and U29074 (N_29074,N_21762,N_23814);
nor U29075 (N_29075,N_18144,N_21476);
and U29076 (N_29076,N_22143,N_21619);
and U29077 (N_29077,N_21669,N_20092);
nand U29078 (N_29078,N_23794,N_20991);
or U29079 (N_29079,N_20865,N_18262);
and U29080 (N_29080,N_22181,N_20425);
nor U29081 (N_29081,N_20928,N_20499);
or U29082 (N_29082,N_22059,N_22608);
and U29083 (N_29083,N_22746,N_18218);
nand U29084 (N_29084,N_23983,N_18419);
nor U29085 (N_29085,N_21360,N_20378);
xnor U29086 (N_29086,N_22803,N_18052);
nand U29087 (N_29087,N_19811,N_19195);
xnor U29088 (N_29088,N_18269,N_18546);
xnor U29089 (N_29089,N_19362,N_20160);
and U29090 (N_29090,N_19141,N_21726);
or U29091 (N_29091,N_22650,N_21343);
nand U29092 (N_29092,N_22591,N_20313);
and U29093 (N_29093,N_21602,N_21839);
or U29094 (N_29094,N_23388,N_19472);
or U29095 (N_29095,N_20634,N_20740);
and U29096 (N_29096,N_18039,N_19063);
nand U29097 (N_29097,N_21360,N_22391);
or U29098 (N_29098,N_23457,N_20597);
and U29099 (N_29099,N_22303,N_20784);
xor U29100 (N_29100,N_22951,N_21907);
nand U29101 (N_29101,N_23881,N_22595);
xor U29102 (N_29102,N_20511,N_21147);
xnor U29103 (N_29103,N_18204,N_18707);
xor U29104 (N_29104,N_18278,N_18392);
or U29105 (N_29105,N_21992,N_18552);
nand U29106 (N_29106,N_22461,N_22273);
and U29107 (N_29107,N_18324,N_21013);
xor U29108 (N_29108,N_19632,N_18218);
or U29109 (N_29109,N_18693,N_20624);
nand U29110 (N_29110,N_23848,N_22350);
or U29111 (N_29111,N_20112,N_19205);
nand U29112 (N_29112,N_18230,N_19988);
xnor U29113 (N_29113,N_19015,N_20030);
xnor U29114 (N_29114,N_19351,N_18468);
or U29115 (N_29115,N_20029,N_23729);
or U29116 (N_29116,N_19548,N_22772);
or U29117 (N_29117,N_21551,N_21316);
and U29118 (N_29118,N_22726,N_20627);
and U29119 (N_29119,N_19181,N_21016);
xor U29120 (N_29120,N_19579,N_23814);
and U29121 (N_29121,N_19642,N_21117);
or U29122 (N_29122,N_21030,N_23201);
nand U29123 (N_29123,N_23159,N_22285);
nand U29124 (N_29124,N_20659,N_20209);
nand U29125 (N_29125,N_23187,N_21450);
and U29126 (N_29126,N_18639,N_20218);
xor U29127 (N_29127,N_18543,N_21415);
nor U29128 (N_29128,N_20761,N_23341);
xor U29129 (N_29129,N_20616,N_19932);
xnor U29130 (N_29130,N_20861,N_22916);
and U29131 (N_29131,N_18717,N_21711);
xor U29132 (N_29132,N_21927,N_23094);
and U29133 (N_29133,N_19865,N_23520);
and U29134 (N_29134,N_19159,N_20451);
nor U29135 (N_29135,N_21547,N_18686);
xnor U29136 (N_29136,N_21811,N_21621);
and U29137 (N_29137,N_23250,N_23649);
or U29138 (N_29138,N_18912,N_23009);
nor U29139 (N_29139,N_19551,N_19523);
and U29140 (N_29140,N_20980,N_22066);
xor U29141 (N_29141,N_18022,N_23692);
nor U29142 (N_29142,N_19981,N_22473);
and U29143 (N_29143,N_18520,N_22778);
and U29144 (N_29144,N_19191,N_23381);
nor U29145 (N_29145,N_21658,N_19840);
xor U29146 (N_29146,N_21005,N_23652);
and U29147 (N_29147,N_19325,N_18660);
nor U29148 (N_29148,N_21856,N_23410);
nand U29149 (N_29149,N_21087,N_23095);
nor U29150 (N_29150,N_20520,N_19979);
or U29151 (N_29151,N_18680,N_20633);
xor U29152 (N_29152,N_21823,N_21582);
nor U29153 (N_29153,N_18637,N_19604);
nor U29154 (N_29154,N_18748,N_21338);
nand U29155 (N_29155,N_19479,N_18793);
nand U29156 (N_29156,N_21848,N_22310);
xnor U29157 (N_29157,N_18100,N_21161);
xor U29158 (N_29158,N_18296,N_22405);
or U29159 (N_29159,N_22293,N_23283);
nand U29160 (N_29160,N_23281,N_23135);
xnor U29161 (N_29161,N_22475,N_18911);
nand U29162 (N_29162,N_20807,N_19445);
xor U29163 (N_29163,N_21576,N_23997);
or U29164 (N_29164,N_20494,N_19431);
or U29165 (N_29165,N_23330,N_22275);
and U29166 (N_29166,N_20861,N_19002);
or U29167 (N_29167,N_20394,N_18284);
xor U29168 (N_29168,N_22586,N_19777);
xor U29169 (N_29169,N_21081,N_22310);
nand U29170 (N_29170,N_18234,N_19391);
and U29171 (N_29171,N_21620,N_22144);
and U29172 (N_29172,N_21352,N_21456);
xor U29173 (N_29173,N_20716,N_22114);
xnor U29174 (N_29174,N_22701,N_19658);
xnor U29175 (N_29175,N_23924,N_20735);
or U29176 (N_29176,N_19660,N_22997);
nor U29177 (N_29177,N_22434,N_22975);
nor U29178 (N_29178,N_18871,N_21124);
xnor U29179 (N_29179,N_20148,N_20754);
xor U29180 (N_29180,N_22753,N_23150);
nand U29181 (N_29181,N_20645,N_20922);
nor U29182 (N_29182,N_18843,N_19276);
nand U29183 (N_29183,N_18416,N_20579);
nor U29184 (N_29184,N_18765,N_21064);
nand U29185 (N_29185,N_20393,N_21837);
nand U29186 (N_29186,N_22932,N_19403);
nor U29187 (N_29187,N_22241,N_21858);
nand U29188 (N_29188,N_20246,N_20066);
xnor U29189 (N_29189,N_20856,N_20544);
xor U29190 (N_29190,N_18117,N_19996);
or U29191 (N_29191,N_22425,N_20675);
or U29192 (N_29192,N_20268,N_21659);
nor U29193 (N_29193,N_23596,N_23676);
or U29194 (N_29194,N_22518,N_20288);
nand U29195 (N_29195,N_19010,N_23077);
nor U29196 (N_29196,N_18510,N_23935);
xor U29197 (N_29197,N_18178,N_22384);
nor U29198 (N_29198,N_23275,N_22773);
or U29199 (N_29199,N_21290,N_18224);
nor U29200 (N_29200,N_22804,N_19868);
and U29201 (N_29201,N_19286,N_22728);
nand U29202 (N_29202,N_23316,N_19781);
or U29203 (N_29203,N_22241,N_23625);
nor U29204 (N_29204,N_18238,N_18164);
and U29205 (N_29205,N_23384,N_19821);
and U29206 (N_29206,N_20346,N_21058);
or U29207 (N_29207,N_22978,N_20270);
or U29208 (N_29208,N_18856,N_21305);
and U29209 (N_29209,N_20671,N_19451);
and U29210 (N_29210,N_18785,N_22864);
or U29211 (N_29211,N_20179,N_21251);
xor U29212 (N_29212,N_21967,N_23679);
or U29213 (N_29213,N_18020,N_19154);
and U29214 (N_29214,N_23016,N_21637);
nor U29215 (N_29215,N_19985,N_22081);
and U29216 (N_29216,N_20265,N_19278);
or U29217 (N_29217,N_23346,N_22311);
nor U29218 (N_29218,N_21999,N_22906);
nand U29219 (N_29219,N_18789,N_21688);
xnor U29220 (N_29220,N_23177,N_20500);
and U29221 (N_29221,N_23816,N_18580);
and U29222 (N_29222,N_19442,N_23293);
nand U29223 (N_29223,N_20631,N_22237);
and U29224 (N_29224,N_19491,N_23043);
nor U29225 (N_29225,N_18267,N_20204);
nand U29226 (N_29226,N_22841,N_22314);
xor U29227 (N_29227,N_23637,N_21216);
and U29228 (N_29228,N_22177,N_20580);
or U29229 (N_29229,N_23188,N_18922);
or U29230 (N_29230,N_23188,N_21230);
and U29231 (N_29231,N_18096,N_23295);
and U29232 (N_29232,N_20504,N_23303);
nor U29233 (N_29233,N_20080,N_22073);
xnor U29234 (N_29234,N_20968,N_19838);
or U29235 (N_29235,N_18860,N_21465);
or U29236 (N_29236,N_18062,N_18425);
and U29237 (N_29237,N_20406,N_22026);
and U29238 (N_29238,N_19931,N_22350);
xor U29239 (N_29239,N_18886,N_21424);
or U29240 (N_29240,N_20535,N_21187);
xor U29241 (N_29241,N_19162,N_21051);
xnor U29242 (N_29242,N_23769,N_23434);
and U29243 (N_29243,N_23860,N_23925);
or U29244 (N_29244,N_23031,N_20332);
or U29245 (N_29245,N_23269,N_20648);
or U29246 (N_29246,N_20000,N_18603);
nor U29247 (N_29247,N_23661,N_19004);
nand U29248 (N_29248,N_20673,N_20697);
xnor U29249 (N_29249,N_18984,N_18147);
nor U29250 (N_29250,N_22921,N_19384);
nor U29251 (N_29251,N_20327,N_18924);
and U29252 (N_29252,N_21493,N_21051);
and U29253 (N_29253,N_22724,N_20907);
nand U29254 (N_29254,N_21606,N_19228);
or U29255 (N_29255,N_19166,N_23451);
or U29256 (N_29256,N_23247,N_18920);
and U29257 (N_29257,N_21723,N_18685);
nand U29258 (N_29258,N_19343,N_22926);
or U29259 (N_29259,N_22227,N_22015);
and U29260 (N_29260,N_19322,N_18655);
nand U29261 (N_29261,N_22031,N_20686);
nor U29262 (N_29262,N_22894,N_19008);
nor U29263 (N_29263,N_20199,N_23398);
or U29264 (N_29264,N_20502,N_20334);
nor U29265 (N_29265,N_22277,N_23259);
and U29266 (N_29266,N_22170,N_22322);
nor U29267 (N_29267,N_19418,N_20874);
nor U29268 (N_29268,N_23028,N_18236);
nor U29269 (N_29269,N_23450,N_21441);
or U29270 (N_29270,N_22926,N_18795);
or U29271 (N_29271,N_23395,N_18545);
or U29272 (N_29272,N_23808,N_18521);
nand U29273 (N_29273,N_21028,N_20502);
and U29274 (N_29274,N_23177,N_23537);
and U29275 (N_29275,N_18481,N_20050);
nor U29276 (N_29276,N_21622,N_22316);
nand U29277 (N_29277,N_22236,N_22764);
or U29278 (N_29278,N_20145,N_22973);
and U29279 (N_29279,N_21372,N_18451);
nor U29280 (N_29280,N_19713,N_23643);
nor U29281 (N_29281,N_21958,N_22581);
xnor U29282 (N_29282,N_23528,N_23533);
or U29283 (N_29283,N_23650,N_23154);
or U29284 (N_29284,N_19741,N_22823);
xor U29285 (N_29285,N_22253,N_20719);
nand U29286 (N_29286,N_20942,N_22895);
nor U29287 (N_29287,N_20479,N_23290);
nor U29288 (N_29288,N_18746,N_18977);
nor U29289 (N_29289,N_19147,N_18106);
nor U29290 (N_29290,N_20975,N_18712);
nand U29291 (N_29291,N_22602,N_18263);
and U29292 (N_29292,N_21731,N_23674);
xor U29293 (N_29293,N_19323,N_18866);
xor U29294 (N_29294,N_23313,N_20421);
and U29295 (N_29295,N_19333,N_20507);
xor U29296 (N_29296,N_19369,N_19646);
or U29297 (N_29297,N_23166,N_20003);
or U29298 (N_29298,N_19202,N_23500);
or U29299 (N_29299,N_21493,N_20892);
or U29300 (N_29300,N_23486,N_21693);
xnor U29301 (N_29301,N_23181,N_21302);
nor U29302 (N_29302,N_23187,N_21345);
or U29303 (N_29303,N_23087,N_21568);
or U29304 (N_29304,N_21664,N_18550);
and U29305 (N_29305,N_18868,N_18607);
or U29306 (N_29306,N_23063,N_23632);
nor U29307 (N_29307,N_22295,N_23714);
and U29308 (N_29308,N_19582,N_23191);
or U29309 (N_29309,N_21653,N_19186);
or U29310 (N_29310,N_20861,N_19917);
nor U29311 (N_29311,N_18506,N_19956);
or U29312 (N_29312,N_18911,N_19580);
nand U29313 (N_29313,N_22799,N_19290);
and U29314 (N_29314,N_23384,N_18571);
nor U29315 (N_29315,N_19175,N_18125);
xnor U29316 (N_29316,N_21694,N_18707);
xnor U29317 (N_29317,N_22455,N_19564);
nand U29318 (N_29318,N_18512,N_18702);
xnor U29319 (N_29319,N_19947,N_22214);
or U29320 (N_29320,N_18729,N_22152);
and U29321 (N_29321,N_19555,N_22031);
nand U29322 (N_29322,N_21980,N_20415);
or U29323 (N_29323,N_21970,N_19330);
nor U29324 (N_29324,N_19620,N_22606);
or U29325 (N_29325,N_18126,N_21326);
nand U29326 (N_29326,N_20907,N_19127);
and U29327 (N_29327,N_22358,N_20949);
nand U29328 (N_29328,N_20036,N_19277);
nand U29329 (N_29329,N_20284,N_22081);
nand U29330 (N_29330,N_20667,N_20100);
nor U29331 (N_29331,N_22615,N_20281);
xnor U29332 (N_29332,N_21782,N_19679);
or U29333 (N_29333,N_18164,N_23868);
xnor U29334 (N_29334,N_20363,N_23831);
nand U29335 (N_29335,N_18448,N_19438);
nor U29336 (N_29336,N_23904,N_23634);
nor U29337 (N_29337,N_23495,N_18529);
nor U29338 (N_29338,N_20148,N_18497);
and U29339 (N_29339,N_22235,N_18236);
and U29340 (N_29340,N_21420,N_19099);
nand U29341 (N_29341,N_22138,N_23083);
nand U29342 (N_29342,N_21246,N_23596);
or U29343 (N_29343,N_21002,N_18386);
nand U29344 (N_29344,N_21035,N_19045);
xnor U29345 (N_29345,N_23765,N_20832);
nand U29346 (N_29346,N_23721,N_21703);
nand U29347 (N_29347,N_22280,N_19056);
nand U29348 (N_29348,N_18608,N_20732);
nand U29349 (N_29349,N_21471,N_22954);
nor U29350 (N_29350,N_18143,N_22364);
nor U29351 (N_29351,N_18966,N_23779);
nor U29352 (N_29352,N_21976,N_19121);
nand U29353 (N_29353,N_20599,N_23042);
xnor U29354 (N_29354,N_19152,N_21492);
nand U29355 (N_29355,N_20030,N_20270);
xor U29356 (N_29356,N_19018,N_22765);
and U29357 (N_29357,N_19187,N_18655);
nand U29358 (N_29358,N_20817,N_19088);
nor U29359 (N_29359,N_18607,N_23473);
or U29360 (N_29360,N_20139,N_23020);
xor U29361 (N_29361,N_18525,N_23216);
nand U29362 (N_29362,N_22769,N_21487);
nor U29363 (N_29363,N_18556,N_21203);
nor U29364 (N_29364,N_21412,N_19065);
or U29365 (N_29365,N_23779,N_19822);
or U29366 (N_29366,N_19037,N_21416);
nor U29367 (N_29367,N_18277,N_21381);
and U29368 (N_29368,N_18605,N_18579);
or U29369 (N_29369,N_20582,N_20537);
or U29370 (N_29370,N_20347,N_22238);
nor U29371 (N_29371,N_19531,N_23603);
or U29372 (N_29372,N_21369,N_21768);
and U29373 (N_29373,N_19524,N_19287);
xor U29374 (N_29374,N_20546,N_23281);
nand U29375 (N_29375,N_21524,N_18085);
or U29376 (N_29376,N_18941,N_22816);
xor U29377 (N_29377,N_21098,N_20004);
or U29378 (N_29378,N_23799,N_20565);
nand U29379 (N_29379,N_19070,N_22580);
and U29380 (N_29380,N_21185,N_21985);
nor U29381 (N_29381,N_21358,N_21819);
or U29382 (N_29382,N_20296,N_23197);
and U29383 (N_29383,N_19361,N_21260);
nor U29384 (N_29384,N_18690,N_19655);
or U29385 (N_29385,N_21148,N_23326);
nand U29386 (N_29386,N_23190,N_22967);
or U29387 (N_29387,N_18799,N_22240);
nor U29388 (N_29388,N_19238,N_19801);
nor U29389 (N_29389,N_23902,N_22322);
xnor U29390 (N_29390,N_19160,N_21169);
xor U29391 (N_29391,N_22863,N_23225);
nor U29392 (N_29392,N_18764,N_20411);
or U29393 (N_29393,N_22610,N_18213);
nor U29394 (N_29394,N_20503,N_20676);
xor U29395 (N_29395,N_18439,N_19315);
xor U29396 (N_29396,N_23394,N_22595);
nand U29397 (N_29397,N_23769,N_18483);
or U29398 (N_29398,N_18059,N_18430);
xnor U29399 (N_29399,N_22203,N_23372);
xnor U29400 (N_29400,N_20245,N_23525);
nor U29401 (N_29401,N_19126,N_23863);
nor U29402 (N_29402,N_18673,N_18054);
xnor U29403 (N_29403,N_20264,N_21009);
nand U29404 (N_29404,N_19491,N_23870);
or U29405 (N_29405,N_23308,N_21697);
nand U29406 (N_29406,N_19774,N_20715);
or U29407 (N_29407,N_22763,N_18406);
xnor U29408 (N_29408,N_23932,N_20017);
and U29409 (N_29409,N_18874,N_21003);
and U29410 (N_29410,N_19679,N_23574);
nor U29411 (N_29411,N_23016,N_19106);
and U29412 (N_29412,N_19423,N_18400);
nand U29413 (N_29413,N_18243,N_23758);
xor U29414 (N_29414,N_18348,N_23717);
xor U29415 (N_29415,N_23436,N_23358);
and U29416 (N_29416,N_21585,N_18688);
nand U29417 (N_29417,N_21788,N_19119);
nand U29418 (N_29418,N_21057,N_23125);
nor U29419 (N_29419,N_19774,N_22345);
xnor U29420 (N_29420,N_19833,N_19756);
xnor U29421 (N_29421,N_23197,N_19416);
nor U29422 (N_29422,N_23185,N_21411);
nor U29423 (N_29423,N_23682,N_19937);
xor U29424 (N_29424,N_22888,N_21469);
and U29425 (N_29425,N_20701,N_23121);
or U29426 (N_29426,N_19323,N_19805);
or U29427 (N_29427,N_23404,N_23479);
and U29428 (N_29428,N_18787,N_23289);
and U29429 (N_29429,N_20221,N_20720);
xnor U29430 (N_29430,N_22194,N_19915);
nor U29431 (N_29431,N_22791,N_22575);
nor U29432 (N_29432,N_22305,N_21763);
and U29433 (N_29433,N_19195,N_22107);
and U29434 (N_29434,N_22548,N_19227);
and U29435 (N_29435,N_19069,N_23387);
nor U29436 (N_29436,N_20905,N_23069);
xnor U29437 (N_29437,N_23422,N_19607);
or U29438 (N_29438,N_18444,N_21924);
nor U29439 (N_29439,N_22702,N_18117);
or U29440 (N_29440,N_23495,N_22753);
nand U29441 (N_29441,N_19541,N_21879);
nand U29442 (N_29442,N_18146,N_21122);
nand U29443 (N_29443,N_21520,N_20666);
and U29444 (N_29444,N_23255,N_20091);
and U29445 (N_29445,N_23391,N_19507);
or U29446 (N_29446,N_20916,N_22986);
xnor U29447 (N_29447,N_20734,N_18522);
or U29448 (N_29448,N_21472,N_23398);
nor U29449 (N_29449,N_21134,N_21094);
or U29450 (N_29450,N_18088,N_22554);
xnor U29451 (N_29451,N_22554,N_21884);
xnor U29452 (N_29452,N_22931,N_19974);
nand U29453 (N_29453,N_22163,N_19770);
and U29454 (N_29454,N_20481,N_22421);
or U29455 (N_29455,N_22451,N_20373);
xor U29456 (N_29456,N_19853,N_22653);
xor U29457 (N_29457,N_23921,N_21263);
nand U29458 (N_29458,N_19104,N_23301);
nor U29459 (N_29459,N_19727,N_20622);
nand U29460 (N_29460,N_18966,N_21844);
xnor U29461 (N_29461,N_20496,N_21380);
and U29462 (N_29462,N_20933,N_20771);
nor U29463 (N_29463,N_22994,N_20705);
nor U29464 (N_29464,N_22183,N_20225);
nor U29465 (N_29465,N_21051,N_23918);
xor U29466 (N_29466,N_19329,N_23105);
nand U29467 (N_29467,N_23808,N_20053);
nand U29468 (N_29468,N_22948,N_20672);
or U29469 (N_29469,N_22581,N_18044);
and U29470 (N_29470,N_20006,N_21125);
xor U29471 (N_29471,N_18515,N_22634);
or U29472 (N_29472,N_22983,N_20858);
and U29473 (N_29473,N_23188,N_20025);
or U29474 (N_29474,N_23796,N_21315);
and U29475 (N_29475,N_18113,N_22569);
nor U29476 (N_29476,N_18650,N_18868);
nand U29477 (N_29477,N_21136,N_20911);
xor U29478 (N_29478,N_20387,N_22009);
nor U29479 (N_29479,N_23804,N_18971);
nand U29480 (N_29480,N_20300,N_21195);
nand U29481 (N_29481,N_18985,N_20143);
nor U29482 (N_29482,N_23921,N_18450);
nand U29483 (N_29483,N_19053,N_21788);
or U29484 (N_29484,N_23006,N_19791);
nand U29485 (N_29485,N_23619,N_23523);
nand U29486 (N_29486,N_19487,N_22036);
or U29487 (N_29487,N_19297,N_19104);
and U29488 (N_29488,N_22802,N_22729);
nor U29489 (N_29489,N_23225,N_23321);
nand U29490 (N_29490,N_21969,N_21953);
nand U29491 (N_29491,N_21492,N_23434);
nand U29492 (N_29492,N_23693,N_23863);
nand U29493 (N_29493,N_18540,N_21197);
or U29494 (N_29494,N_21218,N_20735);
or U29495 (N_29495,N_22315,N_20216);
or U29496 (N_29496,N_19413,N_21287);
nand U29497 (N_29497,N_20199,N_19163);
nand U29498 (N_29498,N_23587,N_23393);
or U29499 (N_29499,N_22319,N_18141);
xnor U29500 (N_29500,N_18640,N_22310);
and U29501 (N_29501,N_19915,N_23386);
nor U29502 (N_29502,N_20460,N_21907);
nor U29503 (N_29503,N_20670,N_18107);
nor U29504 (N_29504,N_19374,N_20710);
or U29505 (N_29505,N_21137,N_18599);
nand U29506 (N_29506,N_19694,N_19519);
nand U29507 (N_29507,N_23613,N_18954);
or U29508 (N_29508,N_23841,N_19194);
and U29509 (N_29509,N_19544,N_21795);
xnor U29510 (N_29510,N_18319,N_22169);
xnor U29511 (N_29511,N_20237,N_21091);
nor U29512 (N_29512,N_18359,N_18565);
xor U29513 (N_29513,N_20116,N_22642);
nand U29514 (N_29514,N_22703,N_20527);
and U29515 (N_29515,N_23623,N_19821);
nand U29516 (N_29516,N_18836,N_20588);
and U29517 (N_29517,N_20996,N_20901);
nor U29518 (N_29518,N_19527,N_19249);
or U29519 (N_29519,N_18876,N_23579);
nor U29520 (N_29520,N_19569,N_20381);
nor U29521 (N_29521,N_19249,N_22197);
or U29522 (N_29522,N_22882,N_21322);
and U29523 (N_29523,N_18935,N_23845);
or U29524 (N_29524,N_21093,N_20153);
nand U29525 (N_29525,N_21943,N_20554);
or U29526 (N_29526,N_18694,N_20737);
nand U29527 (N_29527,N_21687,N_19935);
and U29528 (N_29528,N_19434,N_22260);
or U29529 (N_29529,N_23430,N_20162);
nand U29530 (N_29530,N_21925,N_19897);
nand U29531 (N_29531,N_21627,N_19401);
nor U29532 (N_29532,N_20084,N_21467);
nand U29533 (N_29533,N_18779,N_19139);
nor U29534 (N_29534,N_22823,N_19721);
xor U29535 (N_29535,N_21672,N_20806);
xor U29536 (N_29536,N_23002,N_20224);
nor U29537 (N_29537,N_21318,N_22914);
and U29538 (N_29538,N_22917,N_18564);
nor U29539 (N_29539,N_20576,N_22156);
and U29540 (N_29540,N_23899,N_20630);
and U29541 (N_29541,N_20920,N_22706);
or U29542 (N_29542,N_19072,N_21010);
or U29543 (N_29543,N_18975,N_20146);
xor U29544 (N_29544,N_20429,N_22570);
and U29545 (N_29545,N_20434,N_22699);
or U29546 (N_29546,N_22581,N_21864);
nor U29547 (N_29547,N_18424,N_20267);
xor U29548 (N_29548,N_19021,N_18396);
nor U29549 (N_29549,N_18050,N_20919);
or U29550 (N_29550,N_20601,N_18067);
or U29551 (N_29551,N_23323,N_19172);
and U29552 (N_29552,N_18042,N_20450);
nor U29553 (N_29553,N_23051,N_22674);
nand U29554 (N_29554,N_22865,N_22369);
nand U29555 (N_29555,N_18191,N_18148);
xor U29556 (N_29556,N_20008,N_21543);
and U29557 (N_29557,N_20863,N_23331);
or U29558 (N_29558,N_19445,N_18030);
or U29559 (N_29559,N_20445,N_18655);
or U29560 (N_29560,N_22734,N_23970);
nor U29561 (N_29561,N_22367,N_20740);
or U29562 (N_29562,N_22698,N_20710);
xor U29563 (N_29563,N_23773,N_21722);
nand U29564 (N_29564,N_19167,N_20009);
and U29565 (N_29565,N_20163,N_19698);
and U29566 (N_29566,N_20055,N_23042);
nand U29567 (N_29567,N_22382,N_19964);
and U29568 (N_29568,N_19555,N_21840);
or U29569 (N_29569,N_21239,N_18822);
nand U29570 (N_29570,N_22242,N_19815);
or U29571 (N_29571,N_19316,N_22253);
and U29572 (N_29572,N_23658,N_23484);
nand U29573 (N_29573,N_20272,N_22564);
nor U29574 (N_29574,N_21871,N_18660);
and U29575 (N_29575,N_18998,N_21660);
xnor U29576 (N_29576,N_20054,N_20683);
nor U29577 (N_29577,N_22690,N_20295);
nand U29578 (N_29578,N_19505,N_23872);
or U29579 (N_29579,N_22435,N_23219);
xor U29580 (N_29580,N_20728,N_18829);
and U29581 (N_29581,N_20759,N_22716);
and U29582 (N_29582,N_23925,N_22977);
and U29583 (N_29583,N_23005,N_20754);
xor U29584 (N_29584,N_19016,N_20717);
nand U29585 (N_29585,N_21322,N_21141);
nand U29586 (N_29586,N_22802,N_21582);
and U29587 (N_29587,N_21948,N_20406);
nand U29588 (N_29588,N_18323,N_20522);
or U29589 (N_29589,N_21205,N_18294);
or U29590 (N_29590,N_23208,N_23491);
or U29591 (N_29591,N_22416,N_23935);
or U29592 (N_29592,N_21996,N_21398);
nor U29593 (N_29593,N_18926,N_21131);
and U29594 (N_29594,N_19991,N_18773);
or U29595 (N_29595,N_21135,N_22339);
xnor U29596 (N_29596,N_21967,N_20040);
nor U29597 (N_29597,N_21415,N_20512);
nor U29598 (N_29598,N_22785,N_19576);
or U29599 (N_29599,N_19385,N_18689);
nand U29600 (N_29600,N_22510,N_20640);
nand U29601 (N_29601,N_18029,N_22363);
xnor U29602 (N_29602,N_18745,N_18920);
nand U29603 (N_29603,N_21791,N_18626);
or U29604 (N_29604,N_21676,N_19124);
nor U29605 (N_29605,N_18002,N_23584);
and U29606 (N_29606,N_23002,N_18845);
xnor U29607 (N_29607,N_21841,N_22401);
and U29608 (N_29608,N_23195,N_20213);
nor U29609 (N_29609,N_21155,N_18396);
xnor U29610 (N_29610,N_21625,N_18763);
nor U29611 (N_29611,N_21580,N_18150);
nor U29612 (N_29612,N_18527,N_18496);
nor U29613 (N_29613,N_18516,N_22761);
and U29614 (N_29614,N_23421,N_23803);
nor U29615 (N_29615,N_18045,N_19937);
and U29616 (N_29616,N_23154,N_21513);
nor U29617 (N_29617,N_18784,N_19867);
xor U29618 (N_29618,N_20552,N_23385);
xnor U29619 (N_29619,N_19378,N_23197);
or U29620 (N_29620,N_21322,N_21462);
xor U29621 (N_29621,N_19805,N_18293);
nand U29622 (N_29622,N_18400,N_18213);
or U29623 (N_29623,N_18639,N_18557);
or U29624 (N_29624,N_19499,N_22320);
nand U29625 (N_29625,N_21013,N_19235);
nand U29626 (N_29626,N_18006,N_22782);
nor U29627 (N_29627,N_22726,N_21139);
xnor U29628 (N_29628,N_20844,N_23796);
nor U29629 (N_29629,N_20253,N_20835);
and U29630 (N_29630,N_18549,N_18968);
xor U29631 (N_29631,N_23078,N_22890);
nor U29632 (N_29632,N_22405,N_21266);
or U29633 (N_29633,N_23998,N_20010);
nand U29634 (N_29634,N_18611,N_23929);
or U29635 (N_29635,N_22320,N_19770);
xor U29636 (N_29636,N_21944,N_22602);
nand U29637 (N_29637,N_18121,N_22925);
and U29638 (N_29638,N_22898,N_21024);
and U29639 (N_29639,N_23106,N_22209);
xnor U29640 (N_29640,N_23787,N_22285);
and U29641 (N_29641,N_19376,N_18616);
nor U29642 (N_29642,N_22710,N_22206);
nand U29643 (N_29643,N_21654,N_19942);
nand U29644 (N_29644,N_19608,N_23595);
or U29645 (N_29645,N_18074,N_20274);
nor U29646 (N_29646,N_20556,N_19564);
xor U29647 (N_29647,N_23707,N_18891);
xor U29648 (N_29648,N_21471,N_22523);
nor U29649 (N_29649,N_22291,N_21174);
and U29650 (N_29650,N_21805,N_20673);
or U29651 (N_29651,N_21392,N_23732);
xnor U29652 (N_29652,N_18808,N_22503);
xor U29653 (N_29653,N_22400,N_20873);
or U29654 (N_29654,N_22748,N_22954);
xor U29655 (N_29655,N_18884,N_20641);
or U29656 (N_29656,N_23483,N_18409);
nand U29657 (N_29657,N_21912,N_23712);
nor U29658 (N_29658,N_20393,N_19716);
nor U29659 (N_29659,N_21822,N_18955);
or U29660 (N_29660,N_23361,N_22185);
xor U29661 (N_29661,N_22013,N_22004);
xnor U29662 (N_29662,N_19312,N_22702);
xor U29663 (N_29663,N_21066,N_23884);
and U29664 (N_29664,N_22898,N_22632);
nor U29665 (N_29665,N_18484,N_18004);
or U29666 (N_29666,N_20228,N_22035);
xnor U29667 (N_29667,N_20843,N_18739);
or U29668 (N_29668,N_18663,N_22736);
nand U29669 (N_29669,N_22918,N_18196);
xnor U29670 (N_29670,N_23720,N_18893);
nor U29671 (N_29671,N_21557,N_21469);
nand U29672 (N_29672,N_23824,N_23335);
nand U29673 (N_29673,N_21495,N_19820);
nor U29674 (N_29674,N_18079,N_18906);
or U29675 (N_29675,N_18815,N_21079);
and U29676 (N_29676,N_20776,N_23560);
xor U29677 (N_29677,N_21114,N_22264);
nor U29678 (N_29678,N_23610,N_19821);
and U29679 (N_29679,N_18940,N_23701);
nand U29680 (N_29680,N_19364,N_19165);
and U29681 (N_29681,N_23723,N_21521);
xnor U29682 (N_29682,N_21008,N_22131);
xnor U29683 (N_29683,N_21804,N_20346);
and U29684 (N_29684,N_20995,N_19309);
or U29685 (N_29685,N_22205,N_23061);
xor U29686 (N_29686,N_22856,N_20753);
xor U29687 (N_29687,N_19384,N_22670);
xor U29688 (N_29688,N_21488,N_21283);
or U29689 (N_29689,N_19458,N_19075);
xor U29690 (N_29690,N_19076,N_18114);
and U29691 (N_29691,N_22870,N_23252);
xnor U29692 (N_29692,N_20860,N_21065);
xor U29693 (N_29693,N_18118,N_23897);
nand U29694 (N_29694,N_22006,N_21987);
and U29695 (N_29695,N_23237,N_23440);
and U29696 (N_29696,N_22227,N_22507);
or U29697 (N_29697,N_19114,N_23833);
nor U29698 (N_29698,N_23953,N_21496);
nor U29699 (N_29699,N_22448,N_22972);
or U29700 (N_29700,N_18777,N_19282);
and U29701 (N_29701,N_19395,N_20076);
or U29702 (N_29702,N_18728,N_18952);
or U29703 (N_29703,N_22859,N_21834);
xnor U29704 (N_29704,N_23290,N_19466);
nand U29705 (N_29705,N_19988,N_23696);
xor U29706 (N_29706,N_18926,N_18908);
nor U29707 (N_29707,N_22172,N_21283);
or U29708 (N_29708,N_18235,N_18154);
and U29709 (N_29709,N_18459,N_23476);
and U29710 (N_29710,N_20275,N_20775);
or U29711 (N_29711,N_19476,N_21386);
and U29712 (N_29712,N_22725,N_18813);
nand U29713 (N_29713,N_18005,N_20854);
xor U29714 (N_29714,N_20882,N_22376);
or U29715 (N_29715,N_18067,N_19547);
nand U29716 (N_29716,N_18269,N_18010);
nor U29717 (N_29717,N_23913,N_23666);
nor U29718 (N_29718,N_18639,N_20932);
xor U29719 (N_29719,N_18098,N_21137);
xnor U29720 (N_29720,N_19035,N_20502);
nand U29721 (N_29721,N_23685,N_20165);
and U29722 (N_29722,N_22345,N_22518);
or U29723 (N_29723,N_20771,N_18896);
nand U29724 (N_29724,N_21551,N_20746);
nor U29725 (N_29725,N_20779,N_19301);
and U29726 (N_29726,N_23260,N_22649);
and U29727 (N_29727,N_20532,N_19922);
nor U29728 (N_29728,N_23080,N_21100);
or U29729 (N_29729,N_20499,N_19424);
or U29730 (N_29730,N_20452,N_18001);
and U29731 (N_29731,N_23820,N_19058);
or U29732 (N_29732,N_20039,N_19552);
nand U29733 (N_29733,N_21969,N_21731);
or U29734 (N_29734,N_21697,N_19845);
and U29735 (N_29735,N_21506,N_18219);
and U29736 (N_29736,N_23010,N_20225);
nor U29737 (N_29737,N_20129,N_22570);
and U29738 (N_29738,N_19470,N_23057);
xnor U29739 (N_29739,N_18767,N_22985);
nor U29740 (N_29740,N_19832,N_22309);
nor U29741 (N_29741,N_23018,N_21520);
and U29742 (N_29742,N_18615,N_20846);
nand U29743 (N_29743,N_21802,N_21207);
or U29744 (N_29744,N_20839,N_20951);
or U29745 (N_29745,N_22412,N_21864);
and U29746 (N_29746,N_20749,N_23922);
nor U29747 (N_29747,N_21397,N_23582);
nand U29748 (N_29748,N_18418,N_18046);
and U29749 (N_29749,N_21934,N_22404);
nor U29750 (N_29750,N_19398,N_22533);
and U29751 (N_29751,N_20597,N_22556);
nand U29752 (N_29752,N_23899,N_22799);
or U29753 (N_29753,N_21803,N_22754);
or U29754 (N_29754,N_22601,N_19463);
and U29755 (N_29755,N_21386,N_22255);
nand U29756 (N_29756,N_18276,N_21739);
or U29757 (N_29757,N_20834,N_20414);
and U29758 (N_29758,N_23459,N_21772);
nand U29759 (N_29759,N_21748,N_20885);
xnor U29760 (N_29760,N_23173,N_23675);
xor U29761 (N_29761,N_19803,N_23825);
and U29762 (N_29762,N_19997,N_21808);
and U29763 (N_29763,N_23439,N_23778);
nand U29764 (N_29764,N_18412,N_20826);
xor U29765 (N_29765,N_22297,N_22487);
xor U29766 (N_29766,N_21898,N_18080);
and U29767 (N_29767,N_21319,N_22541);
nand U29768 (N_29768,N_23875,N_19928);
nand U29769 (N_29769,N_19184,N_19822);
xor U29770 (N_29770,N_18573,N_19746);
or U29771 (N_29771,N_18307,N_18591);
or U29772 (N_29772,N_18540,N_20117);
xnor U29773 (N_29773,N_21781,N_23533);
or U29774 (N_29774,N_20208,N_23435);
nand U29775 (N_29775,N_19014,N_18776);
nand U29776 (N_29776,N_22930,N_21802);
nor U29777 (N_29777,N_19655,N_18922);
nand U29778 (N_29778,N_22441,N_19294);
and U29779 (N_29779,N_21523,N_21257);
and U29780 (N_29780,N_22691,N_23483);
or U29781 (N_29781,N_21159,N_20173);
xnor U29782 (N_29782,N_20391,N_23593);
nand U29783 (N_29783,N_21264,N_21666);
and U29784 (N_29784,N_20161,N_19000);
nand U29785 (N_29785,N_22387,N_21867);
nand U29786 (N_29786,N_21856,N_19969);
or U29787 (N_29787,N_22477,N_18896);
and U29788 (N_29788,N_21415,N_20710);
nand U29789 (N_29789,N_23263,N_23078);
xnor U29790 (N_29790,N_22221,N_19447);
or U29791 (N_29791,N_18596,N_22559);
nor U29792 (N_29792,N_23562,N_21936);
nor U29793 (N_29793,N_21573,N_18154);
and U29794 (N_29794,N_19322,N_22940);
or U29795 (N_29795,N_18847,N_18106);
nand U29796 (N_29796,N_22887,N_20207);
xor U29797 (N_29797,N_21652,N_21536);
and U29798 (N_29798,N_18014,N_22410);
or U29799 (N_29799,N_23728,N_21582);
and U29800 (N_29800,N_23144,N_19006);
xor U29801 (N_29801,N_20163,N_21676);
and U29802 (N_29802,N_19843,N_18989);
nand U29803 (N_29803,N_20303,N_23486);
and U29804 (N_29804,N_18285,N_23195);
or U29805 (N_29805,N_20590,N_20443);
nand U29806 (N_29806,N_19936,N_22378);
nand U29807 (N_29807,N_19162,N_20452);
and U29808 (N_29808,N_19692,N_18501);
and U29809 (N_29809,N_22795,N_18459);
and U29810 (N_29810,N_23349,N_22712);
nor U29811 (N_29811,N_18896,N_21217);
nand U29812 (N_29812,N_21327,N_21810);
nand U29813 (N_29813,N_19410,N_22205);
nand U29814 (N_29814,N_19155,N_22160);
xor U29815 (N_29815,N_22054,N_23322);
xor U29816 (N_29816,N_22641,N_21443);
nand U29817 (N_29817,N_19666,N_20543);
or U29818 (N_29818,N_19222,N_23079);
nor U29819 (N_29819,N_23340,N_22596);
nor U29820 (N_29820,N_20404,N_22355);
and U29821 (N_29821,N_20779,N_23114);
nand U29822 (N_29822,N_20155,N_22416);
nand U29823 (N_29823,N_19003,N_23597);
and U29824 (N_29824,N_19821,N_20665);
nand U29825 (N_29825,N_19700,N_18689);
or U29826 (N_29826,N_19378,N_19916);
nor U29827 (N_29827,N_22787,N_22948);
xor U29828 (N_29828,N_23620,N_18843);
or U29829 (N_29829,N_23455,N_18022);
nand U29830 (N_29830,N_23283,N_21113);
nand U29831 (N_29831,N_20212,N_19491);
and U29832 (N_29832,N_23636,N_21591);
nand U29833 (N_29833,N_20091,N_19080);
and U29834 (N_29834,N_23272,N_20759);
nand U29835 (N_29835,N_20283,N_18294);
and U29836 (N_29836,N_21327,N_18626);
and U29837 (N_29837,N_23972,N_20734);
nand U29838 (N_29838,N_23999,N_20247);
nand U29839 (N_29839,N_22556,N_20664);
and U29840 (N_29840,N_22908,N_19230);
nor U29841 (N_29841,N_23531,N_23213);
xor U29842 (N_29842,N_18975,N_23200);
nand U29843 (N_29843,N_22550,N_21050);
xor U29844 (N_29844,N_22549,N_20380);
and U29845 (N_29845,N_22626,N_23057);
nor U29846 (N_29846,N_21568,N_20722);
and U29847 (N_29847,N_22908,N_23570);
nand U29848 (N_29848,N_23917,N_18273);
and U29849 (N_29849,N_22933,N_22367);
or U29850 (N_29850,N_18380,N_18083);
and U29851 (N_29851,N_18783,N_18383);
or U29852 (N_29852,N_19090,N_22325);
nor U29853 (N_29853,N_21979,N_18132);
nor U29854 (N_29854,N_23383,N_23999);
and U29855 (N_29855,N_18452,N_21977);
and U29856 (N_29856,N_19803,N_18587);
xnor U29857 (N_29857,N_23884,N_22953);
nor U29858 (N_29858,N_21960,N_18464);
nor U29859 (N_29859,N_18736,N_21339);
and U29860 (N_29860,N_22244,N_23176);
nor U29861 (N_29861,N_18259,N_23119);
xor U29862 (N_29862,N_20520,N_18682);
nor U29863 (N_29863,N_21014,N_23204);
and U29864 (N_29864,N_23445,N_23309);
nand U29865 (N_29865,N_18811,N_23210);
nand U29866 (N_29866,N_19762,N_18124);
nand U29867 (N_29867,N_22024,N_21709);
nor U29868 (N_29868,N_23211,N_18140);
and U29869 (N_29869,N_21797,N_18379);
nand U29870 (N_29870,N_19448,N_19392);
or U29871 (N_29871,N_22888,N_21990);
nand U29872 (N_29872,N_21968,N_20430);
xor U29873 (N_29873,N_23374,N_21209);
nand U29874 (N_29874,N_22543,N_18394);
nor U29875 (N_29875,N_19403,N_18696);
xor U29876 (N_29876,N_20474,N_20231);
xnor U29877 (N_29877,N_22407,N_23837);
xnor U29878 (N_29878,N_21218,N_19490);
and U29879 (N_29879,N_18800,N_20284);
or U29880 (N_29880,N_18409,N_19168);
nor U29881 (N_29881,N_18382,N_23960);
or U29882 (N_29882,N_21498,N_22619);
and U29883 (N_29883,N_22440,N_23697);
nor U29884 (N_29884,N_23285,N_19003);
and U29885 (N_29885,N_22277,N_20035);
nor U29886 (N_29886,N_22131,N_21557);
xnor U29887 (N_29887,N_23928,N_21351);
and U29888 (N_29888,N_18842,N_22328);
nand U29889 (N_29889,N_23602,N_22507);
xnor U29890 (N_29890,N_23559,N_19581);
xor U29891 (N_29891,N_23014,N_20393);
or U29892 (N_29892,N_22307,N_20681);
or U29893 (N_29893,N_20085,N_20539);
or U29894 (N_29894,N_21567,N_23850);
nor U29895 (N_29895,N_19995,N_22430);
nor U29896 (N_29896,N_23291,N_20103);
or U29897 (N_29897,N_20343,N_19577);
and U29898 (N_29898,N_19809,N_20749);
nor U29899 (N_29899,N_21358,N_21634);
or U29900 (N_29900,N_18668,N_19088);
nand U29901 (N_29901,N_19039,N_21769);
or U29902 (N_29902,N_19468,N_23810);
or U29903 (N_29903,N_23509,N_22884);
nand U29904 (N_29904,N_20136,N_19572);
and U29905 (N_29905,N_18608,N_19842);
nand U29906 (N_29906,N_20588,N_21262);
xor U29907 (N_29907,N_21725,N_19340);
nand U29908 (N_29908,N_22120,N_21147);
xnor U29909 (N_29909,N_23962,N_23594);
and U29910 (N_29910,N_19372,N_21828);
and U29911 (N_29911,N_22021,N_21911);
and U29912 (N_29912,N_20027,N_22679);
nand U29913 (N_29913,N_18444,N_18398);
or U29914 (N_29914,N_19072,N_20046);
nor U29915 (N_29915,N_19195,N_19354);
nor U29916 (N_29916,N_22557,N_22344);
or U29917 (N_29917,N_21586,N_20543);
xnor U29918 (N_29918,N_18375,N_22463);
xor U29919 (N_29919,N_23137,N_20491);
nor U29920 (N_29920,N_21966,N_22802);
nand U29921 (N_29921,N_20895,N_18743);
xor U29922 (N_29922,N_18395,N_20216);
xnor U29923 (N_29923,N_18828,N_18214);
xor U29924 (N_29924,N_19876,N_18092);
or U29925 (N_29925,N_20198,N_22991);
xor U29926 (N_29926,N_23856,N_22634);
nor U29927 (N_29927,N_18872,N_22371);
and U29928 (N_29928,N_22109,N_22814);
nor U29929 (N_29929,N_22947,N_22424);
or U29930 (N_29930,N_23560,N_21353);
xor U29931 (N_29931,N_20404,N_19157);
and U29932 (N_29932,N_18725,N_23372);
nand U29933 (N_29933,N_21406,N_18898);
nand U29934 (N_29934,N_21788,N_20068);
or U29935 (N_29935,N_19133,N_20557);
nor U29936 (N_29936,N_18059,N_18561);
nor U29937 (N_29937,N_20382,N_22478);
nand U29938 (N_29938,N_21907,N_18894);
nand U29939 (N_29939,N_18569,N_20069);
or U29940 (N_29940,N_18293,N_22149);
or U29941 (N_29941,N_18876,N_18220);
nor U29942 (N_29942,N_18957,N_18013);
and U29943 (N_29943,N_22244,N_22525);
xnor U29944 (N_29944,N_23062,N_20914);
xor U29945 (N_29945,N_23374,N_21711);
or U29946 (N_29946,N_18459,N_23026);
nand U29947 (N_29947,N_20763,N_21858);
xor U29948 (N_29948,N_21162,N_21026);
and U29949 (N_29949,N_20026,N_22170);
nor U29950 (N_29950,N_23128,N_22088);
nor U29951 (N_29951,N_20192,N_22247);
nor U29952 (N_29952,N_19706,N_20997);
xnor U29953 (N_29953,N_21464,N_18806);
and U29954 (N_29954,N_20070,N_20379);
or U29955 (N_29955,N_21809,N_18103);
nand U29956 (N_29956,N_23042,N_19989);
nand U29957 (N_29957,N_23232,N_22431);
nand U29958 (N_29958,N_21485,N_19889);
nor U29959 (N_29959,N_23151,N_18834);
xor U29960 (N_29960,N_20542,N_21567);
or U29961 (N_29961,N_18031,N_19560);
and U29962 (N_29962,N_23919,N_22923);
xnor U29963 (N_29963,N_20572,N_21726);
nor U29964 (N_29964,N_20333,N_19846);
nor U29965 (N_29965,N_23870,N_18040);
xnor U29966 (N_29966,N_23808,N_19243);
xnor U29967 (N_29967,N_19866,N_20498);
and U29968 (N_29968,N_21445,N_21628);
and U29969 (N_29969,N_22735,N_20767);
nand U29970 (N_29970,N_22180,N_18491);
nand U29971 (N_29971,N_23864,N_22025);
nand U29972 (N_29972,N_23120,N_23663);
nand U29973 (N_29973,N_22415,N_19907);
nand U29974 (N_29974,N_23517,N_20429);
xnor U29975 (N_29975,N_19566,N_21180);
and U29976 (N_29976,N_22684,N_22331);
nand U29977 (N_29977,N_18502,N_18436);
xnor U29978 (N_29978,N_20697,N_22427);
or U29979 (N_29979,N_18861,N_19626);
nand U29980 (N_29980,N_23435,N_18944);
or U29981 (N_29981,N_20178,N_23107);
nand U29982 (N_29982,N_22317,N_20989);
nor U29983 (N_29983,N_19943,N_20987);
or U29984 (N_29984,N_23823,N_18567);
nand U29985 (N_29985,N_20380,N_22027);
nor U29986 (N_29986,N_23184,N_21693);
nand U29987 (N_29987,N_20563,N_18940);
nand U29988 (N_29988,N_21411,N_19060);
nand U29989 (N_29989,N_21506,N_22117);
xnor U29990 (N_29990,N_22057,N_21271);
nor U29991 (N_29991,N_19222,N_19799);
nand U29992 (N_29992,N_20872,N_21404);
nand U29993 (N_29993,N_23712,N_18807);
xor U29994 (N_29994,N_23333,N_20288);
or U29995 (N_29995,N_21047,N_22311);
or U29996 (N_29996,N_19332,N_21889);
nor U29997 (N_29997,N_21367,N_22057);
nand U29998 (N_29998,N_23580,N_21357);
and U29999 (N_29999,N_18787,N_21079);
and UO_0 (O_0,N_29899,N_28500);
and UO_1 (O_1,N_29975,N_24501);
and UO_2 (O_2,N_24796,N_26526);
nor UO_3 (O_3,N_26380,N_27398);
and UO_4 (O_4,N_28664,N_29143);
nor UO_5 (O_5,N_28349,N_27041);
and UO_6 (O_6,N_24704,N_27380);
nor UO_7 (O_7,N_24282,N_24544);
nand UO_8 (O_8,N_26221,N_28192);
nand UO_9 (O_9,N_26143,N_27943);
nor UO_10 (O_10,N_24791,N_26436);
xor UO_11 (O_11,N_27909,N_25401);
nand UO_12 (O_12,N_25268,N_26356);
xnor UO_13 (O_13,N_25005,N_29208);
and UO_14 (O_14,N_28739,N_26432);
nand UO_15 (O_15,N_29538,N_29668);
nand UO_16 (O_16,N_24143,N_27706);
xnor UO_17 (O_17,N_28060,N_24406);
or UO_18 (O_18,N_27040,N_27712);
nor UO_19 (O_19,N_25118,N_26282);
and UO_20 (O_20,N_28508,N_27583);
and UO_21 (O_21,N_28259,N_29068);
or UO_22 (O_22,N_27905,N_25151);
and UO_23 (O_23,N_29060,N_24500);
or UO_24 (O_24,N_25932,N_27359);
and UO_25 (O_25,N_24570,N_27485);
or UO_26 (O_26,N_26346,N_27999);
or UO_27 (O_27,N_28662,N_29412);
nor UO_28 (O_28,N_27028,N_28417);
nor UO_29 (O_29,N_26111,N_28533);
and UO_30 (O_30,N_27879,N_24977);
and UO_31 (O_31,N_28269,N_25235);
xnor UO_32 (O_32,N_29358,N_28496);
nor UO_33 (O_33,N_27839,N_24163);
xnor UO_34 (O_34,N_28590,N_27813);
or UO_35 (O_35,N_27316,N_24793);
and UO_36 (O_36,N_27295,N_24777);
nand UO_37 (O_37,N_25606,N_27548);
nand UO_38 (O_38,N_27489,N_27928);
nand UO_39 (O_39,N_27244,N_29070);
xor UO_40 (O_40,N_28938,N_27387);
nor UO_41 (O_41,N_25247,N_26600);
nand UO_42 (O_42,N_24205,N_24764);
xor UO_43 (O_43,N_27253,N_28431);
nand UO_44 (O_44,N_24494,N_28412);
nand UO_45 (O_45,N_25298,N_27033);
nor UO_46 (O_46,N_29253,N_25971);
xor UO_47 (O_47,N_28965,N_25747);
and UO_48 (O_48,N_25210,N_25446);
nor UO_49 (O_49,N_29173,N_27546);
or UO_50 (O_50,N_26530,N_28109);
and UO_51 (O_51,N_29431,N_29234);
or UO_52 (O_52,N_29245,N_25748);
and UO_53 (O_53,N_25437,N_24925);
and UO_54 (O_54,N_25583,N_26595);
xnor UO_55 (O_55,N_29804,N_28993);
or UO_56 (O_56,N_29266,N_27200);
nor UO_57 (O_57,N_28405,N_29995);
nand UO_58 (O_58,N_26792,N_24723);
nand UO_59 (O_59,N_26786,N_29388);
nand UO_60 (O_60,N_25432,N_25662);
nor UO_61 (O_61,N_24424,N_28261);
or UO_62 (O_62,N_24467,N_25564);
or UO_63 (O_63,N_26696,N_26212);
nand UO_64 (O_64,N_25811,N_24292);
and UO_65 (O_65,N_24952,N_29507);
nand UO_66 (O_66,N_26387,N_24693);
or UO_67 (O_67,N_25907,N_25391);
nand UO_68 (O_68,N_24134,N_27037);
nand UO_69 (O_69,N_27711,N_24595);
xor UO_70 (O_70,N_24060,N_25261);
and UO_71 (O_71,N_26107,N_26078);
or UO_72 (O_72,N_28146,N_25392);
or UO_73 (O_73,N_25678,N_28848);
xnor UO_74 (O_74,N_25043,N_29398);
and UO_75 (O_75,N_27845,N_27978);
nor UO_76 (O_76,N_25368,N_26177);
and UO_77 (O_77,N_29905,N_26395);
or UO_78 (O_78,N_28206,N_26896);
nand UO_79 (O_79,N_25930,N_25554);
and UO_80 (O_80,N_26878,N_29894);
nand UO_81 (O_81,N_29593,N_29048);
and UO_82 (O_82,N_26016,N_29961);
or UO_83 (O_83,N_26331,N_26853);
and UO_84 (O_84,N_26376,N_26516);
or UO_85 (O_85,N_28277,N_24170);
nand UO_86 (O_86,N_28438,N_25617);
and UO_87 (O_87,N_26303,N_27927);
or UO_88 (O_88,N_26049,N_25040);
nand UO_89 (O_89,N_29135,N_27347);
and UO_90 (O_90,N_24183,N_27341);
nor UO_91 (O_91,N_29564,N_29373);
xor UO_92 (O_92,N_24632,N_28542);
nand UO_93 (O_93,N_24728,N_26843);
xor UO_94 (O_94,N_27973,N_28086);
xnor UO_95 (O_95,N_27588,N_26525);
xnor UO_96 (O_96,N_25100,N_29998);
nor UO_97 (O_97,N_29230,N_26003);
xnor UO_98 (O_98,N_25683,N_29973);
nand UO_99 (O_99,N_26233,N_26392);
nand UO_100 (O_100,N_24833,N_28850);
xnor UO_101 (O_101,N_26827,N_28199);
nand UO_102 (O_102,N_26673,N_26535);
or UO_103 (O_103,N_29891,N_29274);
or UO_104 (O_104,N_26446,N_26637);
nand UO_105 (O_105,N_25305,N_25624);
or UO_106 (O_106,N_27024,N_26183);
xor UO_107 (O_107,N_27611,N_27190);
or UO_108 (O_108,N_25963,N_24617);
and UO_109 (O_109,N_24225,N_24253);
xnor UO_110 (O_110,N_28760,N_24257);
and UO_111 (O_111,N_25122,N_25902);
nand UO_112 (O_112,N_27268,N_24047);
xor UO_113 (O_113,N_24882,N_24584);
and UO_114 (O_114,N_29183,N_25433);
or UO_115 (O_115,N_29424,N_27188);
nand UO_116 (O_116,N_28375,N_26803);
nand UO_117 (O_117,N_25503,N_26857);
nand UO_118 (O_118,N_29236,N_27364);
and UO_119 (O_119,N_24107,N_28224);
nor UO_120 (O_120,N_25762,N_29484);
xor UO_121 (O_121,N_28725,N_28562);
nand UO_122 (O_122,N_29697,N_27699);
xnor UO_123 (O_123,N_28550,N_27592);
nand UO_124 (O_124,N_27587,N_26531);
nor UO_125 (O_125,N_26597,N_28386);
xnor UO_126 (O_126,N_24930,N_26201);
nand UO_127 (O_127,N_29608,N_25360);
xor UO_128 (O_128,N_25652,N_25817);
nand UO_129 (O_129,N_25450,N_29103);
nand UO_130 (O_130,N_28291,N_29807);
and UO_131 (O_131,N_26155,N_25011);
nor UO_132 (O_132,N_28377,N_26189);
or UO_133 (O_133,N_24733,N_26678);
nor UO_134 (O_134,N_24069,N_25862);
and UO_135 (O_135,N_26650,N_29683);
and UO_136 (O_136,N_29286,N_27785);
nor UO_137 (O_137,N_28221,N_24711);
and UO_138 (O_138,N_27768,N_25426);
nand UO_139 (O_139,N_26795,N_25160);
or UO_140 (O_140,N_26855,N_29893);
nor UO_141 (O_141,N_28359,N_25171);
nand UO_142 (O_142,N_27258,N_27513);
or UO_143 (O_143,N_26998,N_25327);
and UO_144 (O_144,N_26912,N_26515);
nand UO_145 (O_145,N_24752,N_25867);
or UO_146 (O_146,N_24110,N_24524);
nor UO_147 (O_147,N_24030,N_27018);
or UO_148 (O_148,N_29156,N_24781);
nor UO_149 (O_149,N_26042,N_25253);
or UO_150 (O_150,N_29205,N_26945);
or UO_151 (O_151,N_27922,N_27545);
or UO_152 (O_152,N_28731,N_28632);
nor UO_153 (O_153,N_25701,N_25256);
or UO_154 (O_154,N_26937,N_29297);
nand UO_155 (O_155,N_28378,N_28583);
or UO_156 (O_156,N_29671,N_26137);
nand UO_157 (O_157,N_26716,N_27171);
xor UO_158 (O_158,N_24363,N_26226);
nand UO_159 (O_159,N_24399,N_25243);
or UO_160 (O_160,N_27824,N_27348);
nor UO_161 (O_161,N_25017,N_24440);
and UO_162 (O_162,N_24997,N_28812);
or UO_163 (O_163,N_29127,N_27735);
xnor UO_164 (O_164,N_28801,N_25124);
nand UO_165 (O_165,N_24883,N_28132);
or UO_166 (O_166,N_29523,N_27882);
xor UO_167 (O_167,N_27697,N_29916);
nand UO_168 (O_168,N_25129,N_25948);
nand UO_169 (O_169,N_24434,N_27919);
or UO_170 (O_170,N_28872,N_26369);
nor UO_171 (O_171,N_27958,N_29741);
xor UO_172 (O_172,N_27720,N_28331);
nor UO_173 (O_173,N_28644,N_24928);
nor UO_174 (O_174,N_27772,N_27032);
xor UO_175 (O_175,N_27254,N_29067);
or UO_176 (O_176,N_24398,N_29501);
nor UO_177 (O_177,N_28433,N_28276);
xor UO_178 (O_178,N_28079,N_26690);
xnor UO_179 (O_179,N_27769,N_26804);
or UO_180 (O_180,N_25047,N_26501);
xor UO_181 (O_181,N_25180,N_28507);
and UO_182 (O_182,N_28975,N_29685);
and UO_183 (O_183,N_26254,N_29781);
xor UO_184 (O_184,N_27576,N_28671);
xnor UO_185 (O_185,N_25396,N_28946);
nor UO_186 (O_186,N_25533,N_24940);
nor UO_187 (O_187,N_29919,N_29256);
nor UO_188 (O_188,N_29394,N_28751);
and UO_189 (O_189,N_28484,N_29906);
and UO_190 (O_190,N_29980,N_24583);
nor UO_191 (O_191,N_24235,N_24348);
nand UO_192 (O_192,N_28587,N_25280);
nand UO_193 (O_193,N_24094,N_24630);
and UO_194 (O_194,N_26301,N_26944);
xnor UO_195 (O_195,N_28350,N_29838);
xor UO_196 (O_196,N_27644,N_28044);
and UO_197 (O_197,N_24820,N_28286);
nand UO_198 (O_198,N_29992,N_29371);
or UO_199 (O_199,N_27161,N_26499);
or UO_200 (O_200,N_26680,N_28636);
nor UO_201 (O_201,N_25894,N_24835);
xor UO_202 (O_202,N_24233,N_26020);
or UO_203 (O_203,N_28399,N_27416);
or UO_204 (O_204,N_24392,N_24957);
or UO_205 (O_205,N_29452,N_24732);
nand UO_206 (O_206,N_25535,N_26075);
and UO_207 (O_207,N_26490,N_26845);
and UO_208 (O_208,N_28290,N_24393);
nor UO_209 (O_209,N_26713,N_26908);
nand UO_210 (O_210,N_24580,N_24284);
nand UO_211 (O_211,N_28035,N_29822);
or UO_212 (O_212,N_24346,N_29531);
nand UO_213 (O_213,N_26262,N_25381);
nor UO_214 (O_214,N_28177,N_29719);
xor UO_215 (O_215,N_27551,N_29739);
or UO_216 (O_216,N_24412,N_26149);
or UO_217 (O_217,N_24070,N_27271);
nor UO_218 (O_218,N_28619,N_29235);
nor UO_219 (O_219,N_28793,N_24989);
and UO_220 (O_220,N_28081,N_29199);
nand UO_221 (O_221,N_29753,N_24378);
nor UO_222 (O_222,N_24578,N_27304);
and UO_223 (O_223,N_27723,N_27305);
and UO_224 (O_224,N_27232,N_28136);
nand UO_225 (O_225,N_24079,N_25479);
or UO_226 (O_226,N_28050,N_27433);
nor UO_227 (O_227,N_26176,N_24809);
and UO_228 (O_228,N_24980,N_28789);
nor UO_229 (O_229,N_26846,N_26310);
or UO_230 (O_230,N_25187,N_27595);
nand UO_231 (O_231,N_24371,N_29698);
xor UO_232 (O_232,N_27532,N_26796);
or UO_233 (O_233,N_24784,N_26314);
nand UO_234 (O_234,N_26780,N_29986);
xor UO_235 (O_235,N_28232,N_28572);
nor UO_236 (O_236,N_27678,N_24615);
and UO_237 (O_237,N_27367,N_28532);
and UO_238 (O_238,N_25164,N_29788);
and UO_239 (O_239,N_25715,N_25289);
or UO_240 (O_240,N_27047,N_28077);
or UO_241 (O_241,N_25008,N_26565);
nand UO_242 (O_242,N_26882,N_27636);
or UO_243 (O_243,N_26194,N_25226);
nor UO_244 (O_244,N_28011,N_24324);
nor UO_245 (O_245,N_26179,N_29492);
nand UO_246 (O_246,N_29572,N_28309);
and UO_247 (O_247,N_29359,N_29567);
xor UO_248 (O_248,N_26390,N_24267);
xor UO_249 (O_249,N_28641,N_29415);
and UO_250 (O_250,N_24579,N_27336);
xor UO_251 (O_251,N_28231,N_25219);
nand UO_252 (O_252,N_26089,N_27464);
nor UO_253 (O_253,N_26811,N_28296);
and UO_254 (O_254,N_24926,N_25599);
nand UO_255 (O_255,N_26311,N_28905);
nor UO_256 (O_256,N_26283,N_24754);
xnor UO_257 (O_257,N_27076,N_26835);
nand UO_258 (O_258,N_27102,N_29469);
nor UO_259 (O_259,N_28229,N_25240);
or UO_260 (O_260,N_25369,N_29882);
and UO_261 (O_261,N_28479,N_28769);
nand UO_262 (O_262,N_25451,N_29666);
nor UO_263 (O_263,N_27748,N_25355);
nor UO_264 (O_264,N_26997,N_29691);
or UO_265 (O_265,N_24289,N_27997);
and UO_266 (O_266,N_27508,N_25032);
nand UO_267 (O_267,N_24484,N_27278);
nand UO_268 (O_268,N_27781,N_27281);
and UO_269 (O_269,N_29699,N_28063);
xor UO_270 (O_270,N_25552,N_24843);
nand UO_271 (O_271,N_24439,N_25816);
or UO_272 (O_272,N_26570,N_28429);
or UO_273 (O_273,N_26767,N_25014);
and UO_274 (O_274,N_24016,N_24731);
and UO_275 (O_275,N_27405,N_27060);
xnor UO_276 (O_276,N_27079,N_29852);
and UO_277 (O_277,N_26222,N_27426);
nor UO_278 (O_278,N_27753,N_25972);
and UO_279 (O_279,N_29485,N_28200);
nor UO_280 (O_280,N_25419,N_26590);
or UO_281 (O_281,N_27414,N_24441);
nor UO_282 (O_282,N_25818,N_25515);
nor UO_283 (O_283,N_26156,N_26861);
xnor UO_284 (O_284,N_27695,N_26290);
xor UO_285 (O_285,N_29249,N_27120);
or UO_286 (O_286,N_26748,N_25382);
and UO_287 (O_287,N_28033,N_25096);
and UO_288 (O_288,N_24574,N_26017);
nand UO_289 (O_289,N_29096,N_29262);
nand UO_290 (O_290,N_26900,N_26759);
nand UO_291 (O_291,N_27467,N_27389);
or UO_292 (O_292,N_29648,N_25260);
and UO_293 (O_293,N_24126,N_28266);
or UO_294 (O_294,N_26326,N_27631);
nor UO_295 (O_295,N_28202,N_27771);
nor UO_296 (O_296,N_29464,N_26308);
nor UO_297 (O_297,N_29247,N_25721);
xor UO_298 (O_298,N_24050,N_26231);
and UO_299 (O_299,N_28088,N_25635);
xor UO_300 (O_300,N_27170,N_29499);
xor UO_301 (O_301,N_27984,N_25820);
nand UO_302 (O_302,N_28312,N_26350);
nand UO_303 (O_303,N_24291,N_24566);
and UO_304 (O_304,N_29563,N_27247);
nand UO_305 (O_305,N_25949,N_25499);
xor UO_306 (O_306,N_26498,N_25542);
nand UO_307 (O_307,N_26132,N_28008);
or UO_308 (O_308,N_29312,N_29372);
and UO_309 (O_309,N_27174,N_26408);
nand UO_310 (O_310,N_28788,N_29057);
or UO_311 (O_311,N_24388,N_28874);
nand UO_312 (O_312,N_25984,N_24465);
or UO_313 (O_313,N_25150,N_26812);
nor UO_314 (O_314,N_26227,N_28581);
nor UO_315 (O_315,N_27091,N_25457);
xor UO_316 (O_316,N_26193,N_25083);
or UO_317 (O_317,N_24770,N_24769);
or UO_318 (O_318,N_25329,N_24314);
nand UO_319 (O_319,N_24181,N_27815);
and UO_320 (O_320,N_28890,N_27825);
or UO_321 (O_321,N_24258,N_29665);
nor UO_322 (O_322,N_26445,N_26976);
and UO_323 (O_323,N_28169,N_28345);
xor UO_324 (O_324,N_25955,N_28714);
or UO_325 (O_325,N_25836,N_25854);
nor UO_326 (O_326,N_27698,N_28054);
or UO_327 (O_327,N_24674,N_24224);
and UO_328 (O_328,N_29308,N_27123);
and UO_329 (O_329,N_27945,N_27320);
xnor UO_330 (O_330,N_28148,N_27312);
nand UO_331 (O_331,N_29032,N_29042);
nor UO_332 (O_332,N_26466,N_28381);
or UO_333 (O_333,N_27435,N_28299);
nor UO_334 (O_334,N_29958,N_24360);
or UO_335 (O_335,N_29138,N_24705);
and UO_336 (O_336,N_29092,N_28629);
nand UO_337 (O_337,N_27383,N_24647);
and UO_338 (O_338,N_29251,N_27614);
or UO_339 (O_339,N_24073,N_27786);
nand UO_340 (O_340,N_29511,N_29692);
or UO_341 (O_341,N_26933,N_27732);
nor UO_342 (O_342,N_24415,N_27780);
nor UO_343 (O_343,N_28219,N_24101);
and UO_344 (O_344,N_24072,N_28028);
xor UO_345 (O_345,N_28185,N_29586);
or UO_346 (O_346,N_27809,N_26405);
nor UO_347 (O_347,N_26011,N_28810);
xnor UO_348 (O_348,N_26139,N_28434);
nand UO_349 (O_349,N_28711,N_29159);
nand UO_350 (O_350,N_24933,N_29900);
or UO_351 (O_351,N_28451,N_24480);
and UO_352 (O_352,N_25675,N_24600);
and UO_353 (O_353,N_26109,N_24007);
nand UO_354 (O_354,N_28693,N_25117);
nor UO_355 (O_355,N_28866,N_28647);
nand UO_356 (O_356,N_24191,N_28411);
or UO_357 (O_357,N_29447,N_27301);
or UO_358 (O_358,N_28330,N_28995);
or UO_359 (O_359,N_24368,N_25506);
nor UO_360 (O_360,N_24066,N_24210);
nor UO_361 (O_361,N_26142,N_29053);
and UO_362 (O_362,N_28716,N_29599);
xnor UO_363 (O_363,N_27070,N_27382);
nor UO_364 (O_364,N_29420,N_29016);
and UO_365 (O_365,N_25656,N_28509);
nor UO_366 (O_366,N_28677,N_29207);
or UO_367 (O_367,N_24032,N_29170);
nand UO_368 (O_368,N_26551,N_28924);
nor UO_369 (O_369,N_29456,N_26777);
or UO_370 (O_370,N_29473,N_29907);
nand UO_371 (O_371,N_25839,N_28141);
nand UO_372 (O_372,N_27556,N_28165);
nand UO_373 (O_373,N_27319,N_25075);
or UO_374 (O_374,N_25567,N_25245);
nor UO_375 (O_375,N_24238,N_28197);
nand UO_376 (O_376,N_26019,N_25562);
or UO_377 (O_377,N_28317,N_26297);
xor UO_378 (O_378,N_25945,N_28821);
nand UO_379 (O_379,N_29267,N_28503);
nor UO_380 (O_380,N_25141,N_24771);
nor UO_381 (O_381,N_26862,N_27891);
or UO_382 (O_382,N_25814,N_24495);
and UO_383 (O_383,N_27523,N_27075);
and UO_384 (O_384,N_26919,N_25629);
and UO_385 (O_385,N_25900,N_26292);
nand UO_386 (O_386,N_25258,N_27671);
xnor UO_387 (O_387,N_26035,N_29397);
xor UO_388 (O_388,N_28875,N_28845);
nor UO_389 (O_389,N_26118,N_29097);
or UO_390 (O_390,N_28740,N_25486);
xor UO_391 (O_391,N_25544,N_25592);
and UO_392 (O_392,N_26245,N_25349);
nand UO_393 (O_393,N_26722,N_29843);
nor UO_394 (O_394,N_26877,N_26553);
nor UO_395 (O_395,N_29816,N_25222);
and UO_396 (O_396,N_25317,N_28006);
or UO_397 (O_397,N_25680,N_28745);
nand UO_398 (O_398,N_29912,N_25527);
or UO_399 (O_399,N_25670,N_26665);
or UO_400 (O_400,N_26963,N_26410);
xor UO_401 (O_401,N_26477,N_27555);
nor UO_402 (O_402,N_26363,N_29494);
and UO_403 (O_403,N_27519,N_27952);
and UO_404 (O_404,N_24335,N_24535);
or UO_405 (O_405,N_24538,N_24092);
and UO_406 (O_406,N_29524,N_25959);
or UO_407 (O_407,N_25078,N_27888);
nand UO_408 (O_408,N_28355,N_28954);
and UO_409 (O_409,N_24902,N_27242);
nor UO_410 (O_410,N_26925,N_26216);
nand UO_411 (O_411,N_24816,N_25135);
or UO_412 (O_412,N_29659,N_24559);
and UO_413 (O_413,N_24744,N_25571);
nand UO_414 (O_414,N_25602,N_27954);
xnor UO_415 (O_415,N_27757,N_27220);
xor UO_416 (O_416,N_26732,N_24985);
and UO_417 (O_417,N_26148,N_25837);
and UO_418 (O_418,N_27949,N_27245);
xor UO_419 (O_419,N_28736,N_28002);
or UO_420 (O_420,N_27897,N_29968);
and UO_421 (O_421,N_28908,N_27071);
and UO_422 (O_422,N_28152,N_25330);
or UO_423 (O_423,N_27443,N_29033);
nand UO_424 (O_424,N_28482,N_27297);
and UO_425 (O_425,N_28163,N_25434);
or UO_426 (O_426,N_24259,N_28419);
and UO_427 (O_427,N_25545,N_27452);
nor UO_428 (O_428,N_26204,N_24068);
xnor UO_429 (O_429,N_29214,N_25332);
nand UO_430 (O_430,N_25466,N_27550);
or UO_431 (O_431,N_27558,N_26728);
and UO_432 (O_432,N_26624,N_25018);
xor UO_433 (O_433,N_29121,N_29962);
and UO_434 (O_434,N_27828,N_24180);
or UO_435 (O_435,N_28452,N_24539);
nor UO_436 (O_436,N_27101,N_26999);
nor UO_437 (O_437,N_26213,N_26655);
or UO_438 (O_438,N_26284,N_27350);
xnor UO_439 (O_439,N_24536,N_28753);
nand UO_440 (O_440,N_26230,N_24353);
and UO_441 (O_441,N_29688,N_26141);
or UO_442 (O_442,N_29377,N_26966);
nand UO_443 (O_443,N_24215,N_24694);
and UO_444 (O_444,N_26105,N_25229);
or UO_445 (O_445,N_27777,N_27783);
and UO_446 (O_446,N_27417,N_28670);
nor UO_447 (O_447,N_29503,N_28588);
and UO_448 (O_448,N_26724,N_27539);
xor UO_449 (O_449,N_29851,N_28042);
or UO_450 (O_450,N_25732,N_24420);
or UO_451 (O_451,N_25312,N_27422);
nand UO_452 (O_452,N_29509,N_26385);
nor UO_453 (O_453,N_26625,N_27237);
nor UO_454 (O_454,N_25607,N_27862);
or UO_455 (O_455,N_25573,N_24760);
or UO_456 (O_456,N_24942,N_26569);
and UO_457 (O_457,N_29418,N_28067);
nor UO_458 (O_458,N_24206,N_26652);
or UO_459 (O_459,N_25104,N_28837);
nand UO_460 (O_460,N_25851,N_24199);
or UO_461 (O_461,N_26903,N_24626);
and UO_462 (O_462,N_25576,N_27151);
and UO_463 (O_463,N_25859,N_27477);
xor UO_464 (O_464,N_27648,N_28339);
nand UO_465 (O_465,N_24741,N_25668);
nand UO_466 (O_466,N_28649,N_28594);
nand UO_467 (O_467,N_28806,N_28110);
xor UO_468 (O_468,N_25128,N_27603);
xor UO_469 (O_469,N_24890,N_26805);
nand UO_470 (O_470,N_27722,N_24884);
or UO_471 (O_471,N_25755,N_29984);
and UO_472 (O_472,N_29265,N_26327);
nand UO_473 (O_473,N_28696,N_27444);
and UO_474 (O_474,N_25553,N_28688);
xor UO_475 (O_475,N_24148,N_28226);
nand UO_476 (O_476,N_29113,N_28818);
nand UO_477 (O_477,N_25543,N_24065);
nand UO_478 (O_478,N_24246,N_25526);
nor UO_479 (O_479,N_24774,N_29284);
nand UO_480 (O_480,N_26129,N_28880);
and UO_481 (O_481,N_26083,N_27798);
or UO_482 (O_482,N_29395,N_26634);
nor UO_483 (O_483,N_28668,N_29756);
nand UO_484 (O_484,N_25136,N_26415);
nor UO_485 (O_485,N_25379,N_29433);
or UO_486 (O_486,N_28175,N_27049);
nor UO_487 (O_487,N_29180,N_24596);
and UO_488 (O_488,N_29201,N_24988);
and UO_489 (O_489,N_27600,N_27817);
xor UO_490 (O_490,N_28406,N_28173);
nor UO_491 (O_491,N_26099,N_28285);
or UO_492 (O_492,N_26951,N_24487);
nand UO_493 (O_493,N_29336,N_29796);
nor UO_494 (O_494,N_27038,N_25735);
and UO_495 (O_495,N_24976,N_26091);
or UO_496 (O_496,N_28023,N_25711);
nor UO_497 (O_497,N_27008,N_28105);
and UO_498 (O_498,N_24603,N_26286);
nand UO_499 (O_499,N_27335,N_28613);
xnor UO_500 (O_500,N_25665,N_25266);
nor UO_501 (O_501,N_28524,N_25212);
and UO_502 (O_502,N_26867,N_27841);
nor UO_503 (O_503,N_27223,N_29941);
and UO_504 (O_504,N_27796,N_24842);
nor UO_505 (O_505,N_28974,N_24577);
nor UO_506 (O_506,N_26989,N_26199);
nor UO_507 (O_507,N_25962,N_25190);
nand UO_508 (O_508,N_29667,N_26729);
xor UO_509 (O_509,N_24682,N_29014);
nand UO_510 (O_510,N_25509,N_24317);
nand UO_511 (O_511,N_24250,N_29078);
nor UO_512 (O_512,N_28732,N_28362);
and UO_513 (O_513,N_27266,N_29226);
xnor UO_514 (O_514,N_24543,N_25203);
nor UO_515 (O_515,N_28699,N_26398);
nor UO_516 (O_516,N_29109,N_26317);
or UO_517 (O_517,N_28346,N_29309);
xnor UO_518 (O_518,N_27360,N_28672);
nand UO_519 (O_519,N_27229,N_27202);
or UO_520 (O_520,N_24433,N_29740);
nand UO_521 (O_521,N_28321,N_24167);
nor UO_522 (O_522,N_27080,N_26952);
xnor UO_523 (O_523,N_29824,N_26585);
or UO_524 (O_524,N_26287,N_25643);
nand UO_525 (O_525,N_24061,N_26828);
or UO_526 (O_526,N_25548,N_24507);
nor UO_527 (O_527,N_29031,N_24868);
nand UO_528 (O_528,N_25992,N_25581);
or UO_529 (O_529,N_24290,N_28007);
or UO_530 (O_530,N_25045,N_29512);
nand UO_531 (O_531,N_29211,N_25055);
xnor UO_532 (O_532,N_29561,N_24160);
nor UO_533 (O_533,N_27868,N_28213);
nand UO_534 (O_534,N_27212,N_29736);
nor UO_535 (O_535,N_27338,N_28529);
nand UO_536 (O_536,N_29064,N_28166);
nor UO_537 (O_537,N_29058,N_26394);
and UO_538 (O_538,N_25677,N_27052);
nor UO_539 (O_539,N_26497,N_26586);
xnor UO_540 (O_540,N_24027,N_29310);
nor UO_541 (O_541,N_26787,N_25989);
nor UO_542 (O_542,N_25452,N_27626);
and UO_543 (O_543,N_26617,N_28000);
or UO_544 (O_544,N_25609,N_24018);
and UO_545 (O_545,N_25560,N_29546);
and UO_546 (O_546,N_28655,N_26626);
nand UO_547 (O_547,N_26603,N_24384);
xnor UO_548 (O_548,N_24528,N_26145);
xnor UO_549 (O_549,N_29562,N_28743);
or UO_550 (O_550,N_28846,N_27669);
xor UO_551 (O_551,N_24223,N_24075);
nor UO_552 (O_552,N_25259,N_24742);
nand UO_553 (O_553,N_28642,N_25402);
and UO_554 (O_554,N_24877,N_28034);
xor UO_555 (O_555,N_29602,N_28335);
or UO_556 (O_556,N_27890,N_25608);
nand UO_557 (O_557,N_29396,N_24643);
and UO_558 (O_558,N_25956,N_25507);
xor UO_559 (O_559,N_26540,N_25633);
or UO_560 (O_560,N_28620,N_26476);
or UO_561 (O_561,N_25698,N_24776);
nor UO_562 (O_562,N_24227,N_24678);
and UO_563 (O_563,N_26444,N_25975);
or UO_564 (O_564,N_27843,N_29856);
and UO_565 (O_565,N_25281,N_29017);
or UO_566 (O_566,N_28133,N_27988);
nand UO_567 (O_567,N_24436,N_25423);
nand UO_568 (O_568,N_29744,N_28506);
and UO_569 (O_569,N_27264,N_26768);
or UO_570 (O_570,N_29294,N_26929);
or UO_571 (O_571,N_28172,N_26758);
nand UO_572 (O_572,N_27313,N_27496);
nor UO_573 (O_573,N_28260,N_26029);
nand UO_574 (O_574,N_25766,N_28304);
nor UO_575 (O_575,N_25438,N_28680);
xor UO_576 (O_576,N_24099,N_25132);
or UO_577 (O_577,N_25910,N_29551);
or UO_578 (O_578,N_25714,N_26077);
nand UO_579 (O_579,N_28920,N_27222);
nand UO_580 (O_580,N_28064,N_29268);
xnor UO_581 (O_581,N_24795,N_27185);
or UO_582 (O_582,N_29332,N_26884);
or UO_583 (O_583,N_26991,N_27492);
nor UO_584 (O_584,N_25057,N_25659);
or UO_585 (O_585,N_25493,N_29462);
and UO_586 (O_586,N_25895,N_29743);
nor UO_587 (O_587,N_24935,N_27153);
or UO_588 (O_588,N_29533,N_25950);
and UO_589 (O_589,N_27022,N_29453);
nor UO_590 (O_590,N_29603,N_28264);
or UO_591 (O_591,N_29970,N_25425);
or UO_592 (O_592,N_29411,N_29313);
nor UO_593 (O_593,N_24758,N_24182);
and UO_594 (O_594,N_25925,N_24709);
xnor UO_595 (O_595,N_26070,N_24716);
or UO_596 (O_596,N_27447,N_26518);
nand UO_597 (O_597,N_28819,N_29333);
nor UO_598 (O_598,N_24703,N_28698);
and UO_599 (O_599,N_26428,N_28786);
or UO_600 (O_600,N_26833,N_28678);
nand UO_601 (O_601,N_29197,N_25084);
nor UO_602 (O_602,N_24866,N_27344);
or UO_603 (O_603,N_28939,N_24525);
xor UO_604 (O_604,N_28841,N_24876);
and UO_605 (O_605,N_24858,N_24811);
nand UO_606 (O_606,N_27323,N_24599);
or UO_607 (O_607,N_24380,N_29393);
or UO_608 (O_608,N_28075,N_24475);
and UO_609 (O_609,N_29246,N_27125);
xor UO_610 (O_610,N_26810,N_27953);
or UO_611 (O_611,N_29560,N_25905);
nand UO_612 (O_612,N_25142,N_26253);
or UO_613 (O_613,N_24240,N_28847);
xor UO_614 (O_614,N_29325,N_25134);
nand UO_615 (O_615,N_28528,N_24056);
nor UO_616 (O_616,N_24715,N_24144);
and UO_617 (O_617,N_26773,N_25563);
and UO_618 (O_618,N_28831,N_25422);
nor UO_619 (O_619,N_27442,N_25759);
xor UO_620 (O_620,N_26184,N_24028);
and UO_621 (O_621,N_28448,N_27448);
and UO_622 (O_622,N_25990,N_25464);
nand UO_623 (O_623,N_24836,N_24906);
nand UO_624 (O_624,N_25865,N_26157);
or UO_625 (O_625,N_24969,N_26645);
xnor UO_626 (O_626,N_26411,N_25522);
nand UO_627 (O_627,N_29553,N_28998);
nand UO_628 (O_628,N_24520,N_24533);
nor UO_629 (O_629,N_24262,N_24278);
xor UO_630 (O_630,N_25985,N_24560);
or UO_631 (O_631,N_26291,N_27203);
nand UO_632 (O_632,N_28795,N_29077);
nor UO_633 (O_633,N_29496,N_25082);
or UO_634 (O_634,N_29348,N_26948);
xor UO_635 (O_635,N_25681,N_29072);
xnor UO_636 (O_636,N_28738,N_29079);
and UO_637 (O_637,N_27472,N_26880);
or UO_638 (O_638,N_24145,N_25341);
nor UO_639 (O_639,N_26472,N_28083);
nand UO_640 (O_640,N_29747,N_24395);
or UO_641 (O_641,N_27754,N_27007);
xnor UO_642 (O_642,N_27230,N_27415);
nor UO_643 (O_643,N_25734,N_24102);
or UO_644 (O_644,N_28403,N_29171);
nor UO_645 (O_645,N_28036,N_27895);
nor UO_646 (O_646,N_27429,N_24921);
xnor UO_647 (O_647,N_26574,N_27094);
or UO_648 (O_648,N_27226,N_25058);
and UO_649 (O_649,N_29999,N_28945);
nand UO_650 (O_650,N_24043,N_24285);
xor UO_651 (O_651,N_27792,N_26894);
and UO_652 (O_652,N_25822,N_27759);
nand UO_653 (O_653,N_28244,N_24443);
or UO_654 (O_654,N_28679,N_26924);
or UO_655 (O_655,N_29877,N_27738);
nand UO_656 (O_656,N_29287,N_26694);
and UO_657 (O_657,N_25170,N_25685);
and UO_658 (O_658,N_28640,N_29335);
xnor UO_659 (O_659,N_28784,N_29223);
and UO_660 (O_660,N_28947,N_29327);
or UO_661 (O_661,N_28194,N_25269);
or UO_662 (O_662,N_25185,N_27450);
nand UO_663 (O_663,N_27111,N_24222);
nor UO_664 (O_664,N_25676,N_26100);
nor UO_665 (O_665,N_25080,N_26985);
nor UO_666 (O_666,N_27001,N_27178);
nand UO_667 (O_667,N_27369,N_26299);
and UO_668 (O_668,N_26856,N_29965);
xnor UO_669 (O_669,N_27917,N_24807);
nand UO_670 (O_670,N_29351,N_26192);
xnor UO_671 (O_671,N_24518,N_24124);
xor UO_672 (O_672,N_26909,N_27659);
nand UO_673 (O_673,N_27186,N_27993);
nor UO_674 (O_674,N_29026,N_28342);
or UO_675 (O_675,N_26235,N_26270);
nor UO_676 (O_676,N_29772,N_29887);
or UO_677 (O_677,N_26584,N_25821);
and UO_678 (O_678,N_28545,N_29592);
nor UO_679 (O_679,N_27138,N_29352);
nor UO_680 (O_680,N_28987,N_29518);
nand UO_681 (O_681,N_25306,N_29059);
or UO_682 (O_682,N_29018,N_26050);
and UO_683 (O_683,N_25167,N_27651);
and UO_684 (O_684,N_28959,N_28469);
and UO_685 (O_685,N_26923,N_27749);
or UO_686 (O_686,N_24710,N_26580);
nand UO_687 (O_687,N_27842,N_25686);
nand UO_688 (O_688,N_25999,N_26920);
and UO_689 (O_689,N_28896,N_27916);
and UO_690 (O_690,N_27941,N_28635);
and UO_691 (O_691,N_29291,N_24863);
or UO_692 (O_692,N_29200,N_26269);
and UO_693 (O_693,N_29357,N_26334);
and UO_694 (O_694,N_25241,N_28849);
nor UO_695 (O_695,N_24759,N_24171);
or UO_696 (O_696,N_24916,N_25429);
nor UO_697 (O_697,N_25644,N_25311);
and UO_698 (O_698,N_24648,N_26409);
nand UO_699 (O_699,N_25850,N_26116);
nand UO_700 (O_700,N_25359,N_24681);
nand UO_701 (O_701,N_24555,N_28774);
or UO_702 (O_702,N_26972,N_28567);
or UO_703 (O_703,N_24367,N_24377);
and UO_704 (O_704,N_26134,N_26800);
or UO_705 (O_705,N_25209,N_25877);
xor UO_706 (O_706,N_27156,N_29093);
xnor UO_707 (O_707,N_28316,N_26737);
xor UO_708 (O_708,N_25880,N_24328);
and UO_709 (O_709,N_27036,N_26940);
nor UO_710 (O_710,N_28765,N_28937);
nor UO_711 (O_711,N_28314,N_24153);
and UO_712 (O_712,N_24294,N_25540);
or UO_713 (O_713,N_24327,N_26140);
nor UO_714 (O_714,N_24476,N_27358);
and UO_715 (O_715,N_28176,N_26246);
or UO_716 (O_716,N_24519,N_25469);
xnor UO_717 (O_717,N_24558,N_27756);
nand UO_718 (O_718,N_29979,N_29924);
xnor UO_719 (O_719,N_25297,N_27218);
xor UO_720 (O_720,N_25896,N_24904);
and UO_721 (O_721,N_27566,N_26417);
xor UO_722 (O_722,N_25794,N_26439);
or UO_723 (O_723,N_27986,N_25671);
nand UO_724 (O_724,N_25931,N_24311);
or UO_725 (O_725,N_28923,N_28340);
nand UO_726 (O_726,N_26293,N_28395);
nand UO_727 (O_727,N_29846,N_27765);
or UO_728 (O_728,N_29936,N_29322);
nand UO_729 (O_729,N_29382,N_28393);
or UO_730 (O_730,N_24019,N_29726);
or UO_731 (O_731,N_24091,N_26053);
xnor UO_732 (O_732,N_24684,N_27675);
nor UO_733 (O_733,N_25374,N_27340);
or UO_734 (O_734,N_28313,N_28142);
or UO_735 (O_735,N_25657,N_27441);
nor UO_736 (O_736,N_29557,N_28673);
xor UO_737 (O_737,N_29552,N_26829);
and UO_738 (O_738,N_27616,N_24428);
and UO_739 (O_739,N_29375,N_29777);
and UO_740 (O_740,N_24639,N_27349);
or UO_741 (O_741,N_27043,N_24251);
nor UO_742 (O_742,N_27553,N_28440);
and UO_743 (O_743,N_24383,N_25569);
nor UO_744 (O_744,N_28311,N_29381);
nand UO_745 (O_745,N_28247,N_29337);
nor UO_746 (O_746,N_26263,N_28230);
or UO_747 (O_747,N_27995,N_26256);
nand UO_748 (O_748,N_26481,N_26375);
and UO_749 (O_749,N_28783,N_24840);
nor UO_750 (O_750,N_26990,N_24837);
nor UO_751 (O_751,N_24880,N_25362);
or UO_752 (O_752,N_24114,N_29362);
or UO_753 (O_753,N_24817,N_29706);
and UO_754 (O_754,N_25216,N_29880);
or UO_755 (O_755,N_24719,N_25250);
and UO_756 (O_756,N_26068,N_29702);
nand UO_757 (O_757,N_28935,N_25666);
and UO_758 (O_758,N_25758,N_28191);
xnor UO_759 (O_759,N_27290,N_26763);
or UO_760 (O_760,N_27408,N_27767);
nor UO_761 (O_761,N_29755,N_24242);
nand UO_762 (O_762,N_27180,N_26699);
nor UO_763 (O_763,N_27666,N_28323);
nor UO_764 (O_764,N_29547,N_29071);
and UO_765 (O_765,N_25244,N_28371);
nand UO_766 (O_766,N_25757,N_26683);
and UO_767 (O_767,N_29010,N_25386);
and UO_768 (O_768,N_29353,N_27597);
and UO_769 (O_769,N_28627,N_28842);
or UO_770 (O_770,N_28450,N_25781);
nand UO_771 (O_771,N_28408,N_29775);
or UO_772 (O_772,N_26527,N_28305);
nor UO_773 (O_773,N_28214,N_25251);
xnor UO_774 (O_774,N_25472,N_26224);
and UO_775 (O_775,N_25183,N_28637);
or UO_776 (O_776,N_26797,N_27148);
nand UO_777 (O_777,N_24334,N_25965);
nand UO_778 (O_778,N_24416,N_27179);
and UO_779 (O_779,N_25769,N_29716);
xnor UO_780 (O_780,N_24209,N_24459);
xor UO_781 (O_781,N_29949,N_29589);
and UO_782 (O_782,N_27646,N_26755);
or UO_783 (O_783,N_26686,N_26902);
or UO_784 (O_784,N_29556,N_29278);
nand UO_785 (O_785,N_25852,N_26636);
or UO_786 (O_786,N_26834,N_27751);
or UO_787 (O_787,N_24983,N_29387);
and UO_788 (O_788,N_28615,N_26571);
or UO_789 (O_789,N_29890,N_24999);
or UO_790 (O_790,N_26465,N_28467);
nor UO_791 (O_791,N_25291,N_25443);
and UO_792 (O_792,N_29935,N_27337);
nand UO_793 (O_793,N_27624,N_29790);
nor UO_794 (O_794,N_24722,N_27996);
xnor UO_795 (O_795,N_26992,N_24714);
nand UO_796 (O_796,N_26449,N_28979);
nor UO_797 (O_797,N_26542,N_27964);
or UO_798 (O_798,N_26816,N_26702);
nor UO_799 (O_799,N_28128,N_27676);
xor UO_800 (O_800,N_28624,N_24309);
or UO_801 (O_801,N_29757,N_24505);
nand UO_802 (O_802,N_29952,N_26067);
xor UO_803 (O_803,N_25691,N_29090);
xor UO_804 (O_804,N_25052,N_29141);
and UO_805 (O_805,N_29717,N_25835);
nand UO_806 (O_806,N_25514,N_24821);
xnor UO_807 (O_807,N_27643,N_29202);
or UO_808 (O_808,N_25130,N_27109);
xnor UO_809 (O_809,N_28584,N_28445);
nand UO_810 (O_810,N_27847,N_27096);
nor UO_811 (O_811,N_28130,N_24772);
xor UO_812 (O_812,N_29252,N_26519);
nor UO_813 (O_813,N_29920,N_25785);
nand UO_814 (O_814,N_29855,N_28056);
nor UO_815 (O_815,N_26858,N_28762);
and UO_816 (O_816,N_29673,N_28726);
xor UO_817 (O_817,N_24618,N_27507);
xnor UO_818 (O_818,N_24271,N_25384);
xnor UO_819 (O_819,N_24913,N_27262);
or UO_820 (O_820,N_27691,N_26885);
nand UO_821 (O_821,N_24201,N_24532);
nor UO_822 (O_822,N_25081,N_27957);
nand UO_823 (O_823,N_27088,N_27029);
nor UO_824 (O_824,N_29175,N_24673);
and UO_825 (O_825,N_25086,N_27770);
nor UO_826 (O_826,N_26178,N_28265);
nor UO_827 (O_827,N_28423,N_28724);
or UO_828 (O_828,N_24548,N_26400);
and UO_829 (O_829,N_25322,N_29844);
or UO_830 (O_830,N_28361,N_27221);
xor UO_831 (O_831,N_29007,N_25847);
nand UO_832 (O_832,N_26784,N_27243);
nand UO_833 (O_833,N_25538,N_28106);
nor UO_834 (O_834,N_24510,N_24049);
xor UO_835 (O_835,N_26079,N_29797);
xor UO_836 (O_836,N_25658,N_24657);
or UO_837 (O_837,N_29149,N_29318);
or UO_838 (O_838,N_25424,N_27835);
xnor UO_839 (O_839,N_28435,N_25459);
nand UO_840 (O_840,N_26543,N_29776);
nand UO_841 (O_841,N_27650,N_25873);
and UO_842 (O_842,N_25504,N_27371);
xor UO_843 (O_843,N_27705,N_28980);
nor UO_844 (O_844,N_28207,N_28598);
nand UO_845 (O_845,N_27725,N_27124);
nor UO_846 (O_846,N_26196,N_27902);
or UO_847 (O_847,N_25952,N_24351);
and UO_848 (O_848,N_28483,N_24838);
xor UO_849 (O_849,N_26333,N_25169);
and UO_850 (O_850,N_24423,N_24979);
nor UO_851 (O_851,N_27025,N_25611);
xor UO_852 (O_852,N_25600,N_28135);
nand UO_853 (O_853,N_28883,N_25770);
xnor UO_854 (O_854,N_25650,N_29862);
nor UO_855 (O_855,N_27284,N_29783);
and UO_856 (O_856,N_24404,N_25155);
nor UO_857 (O_857,N_28701,N_28459);
and UO_858 (O_858,N_25938,N_28015);
nand UO_859 (O_859,N_28878,N_28888);
nand UO_860 (O_860,N_27939,N_29259);
or UO_861 (O_861,N_29884,N_29649);
nand UO_862 (O_862,N_26243,N_27165);
nand UO_863 (O_863,N_26653,N_26962);
xnor UO_864 (O_864,N_25351,N_26646);
xnor UO_865 (O_865,N_27209,N_26761);
nand UO_866 (O_866,N_25557,N_26006);
xor UO_867 (O_867,N_29206,N_28097);
nor UO_868 (O_868,N_26957,N_29570);
xor UO_869 (O_869,N_24812,N_29516);
xnor UO_870 (O_870,N_24839,N_25739);
or UO_871 (O_871,N_24850,N_24829);
or UO_872 (O_872,N_24059,N_29445);
and UO_873 (O_873,N_27574,N_26707);
nor UO_874 (O_874,N_25006,N_24039);
nor UO_875 (O_875,N_26239,N_27623);
xnor UO_876 (O_876,N_29111,N_28621);
nor UO_877 (O_877,N_28616,N_25301);
nand UO_878 (O_878,N_25340,N_28196);
and UO_879 (O_879,N_27822,N_29813);
nor UO_880 (O_880,N_28853,N_27859);
and UO_881 (O_881,N_29784,N_24389);
or UO_882 (O_882,N_28009,N_29495);
or UO_883 (O_883,N_27282,N_25470);
xor UO_884 (O_884,N_27317,N_29020);
or UO_885 (O_885,N_27885,N_29653);
xor UO_886 (O_886,N_27034,N_25885);
nor UO_887 (O_887,N_29299,N_27019);
nor UO_888 (O_888,N_29427,N_29129);
or UO_889 (O_889,N_25919,N_29857);
xor UO_890 (O_890,N_24844,N_26364);
and UO_891 (O_891,N_29728,N_29497);
xnor UO_892 (O_892,N_25689,N_26131);
and UO_893 (O_893,N_25709,N_26996);
or UO_894 (O_894,N_24084,N_25586);
xor UO_895 (O_895,N_26007,N_28273);
nand UO_896 (O_896,N_25870,N_25841);
nor UO_897 (O_897,N_27858,N_26071);
xor UO_898 (O_898,N_24470,N_26977);
or UO_899 (O_899,N_24308,N_25660);
xor UO_900 (O_900,N_28222,N_27510);
or UO_901 (O_901,N_28058,N_28369);
or UO_902 (O_902,N_27629,N_28218);
and UO_903 (O_903,N_26341,N_24905);
or UO_904 (O_904,N_28162,N_27602);
or UO_905 (O_905,N_27004,N_28771);
nand UO_906 (O_906,N_29940,N_27568);
xnor UO_907 (O_907,N_29454,N_29836);
nor UO_908 (O_908,N_24594,N_24720);
nand UO_909 (O_909,N_24672,N_27950);
nor UO_910 (O_910,N_26442,N_28887);
or UO_911 (O_911,N_26606,N_26307);
xor UO_912 (O_912,N_25860,N_27175);
or UO_913 (O_913,N_24725,N_29805);
nand UO_914 (O_914,N_29137,N_24692);
nand UO_915 (O_915,N_28882,N_25195);
or UO_916 (O_916,N_27421,N_26315);
nand UO_917 (O_917,N_26691,N_25914);
xnor UO_918 (O_918,N_25906,N_26506);
nor UO_919 (O_919,N_26122,N_29645);
or UO_920 (O_920,N_29929,N_26238);
or UO_921 (O_921,N_28685,N_25532);
xor UO_922 (O_922,N_27141,N_26313);
nor UO_923 (O_923,N_26384,N_24726);
xor UO_924 (O_924,N_24097,N_26370);
xnor UO_925 (O_925,N_26095,N_24450);
and UO_926 (O_926,N_27224,N_29798);
xor UO_927 (O_927,N_25202,N_27627);
nor UO_928 (O_928,N_27883,N_25062);
xor UO_929 (O_929,N_26576,N_25510);
nand UO_930 (O_930,N_29634,N_27594);
or UO_931 (O_931,N_27493,N_26581);
nand UO_932 (O_932,N_27228,N_25805);
nand UO_933 (O_933,N_29241,N_26549);
nor UO_934 (O_934,N_25319,N_26660);
or UO_935 (O_935,N_27605,N_28487);
or UO_936 (O_936,N_27856,N_29361);
and UO_937 (O_937,N_25304,N_25090);
nor UO_938 (O_938,N_27488,N_26599);
xor UO_939 (O_939,N_28858,N_27805);
xnor UO_940 (O_940,N_29027,N_24790);
xor UO_941 (O_941,N_27351,N_25825);
nor UO_942 (O_942,N_26163,N_27030);
nor UO_943 (O_943,N_24899,N_25491);
nor UO_944 (O_944,N_25565,N_27635);
nand UO_945 (O_945,N_27830,N_25716);
or UO_946 (O_946,N_29931,N_24955);
nand UO_947 (O_947,N_27656,N_26228);
xor UO_948 (O_948,N_29232,N_28144);
xnor UO_949 (O_949,N_29969,N_29276);
nand UO_950 (O_950,N_28723,N_24254);
nor UO_951 (O_951,N_28122,N_24125);
nor UO_952 (O_952,N_25347,N_26842);
nand UO_953 (O_953,N_24037,N_27571);
and UO_954 (O_954,N_24451,N_27194);
nor UO_955 (O_955,N_28092,N_29881);
nand UO_956 (O_956,N_29749,N_28076);
nor UO_957 (O_957,N_26778,N_28473);
nor UO_958 (O_958,N_24625,N_27930);
or UO_959 (O_959,N_25603,N_29957);
and UO_960 (O_960,N_24664,N_28952);
nand UO_961 (O_961,N_28658,N_26032);
and UO_962 (O_962,N_28481,N_25441);
or UO_963 (O_963,N_24403,N_28690);
and UO_964 (O_964,N_25856,N_29789);
or UO_965 (O_965,N_28953,N_24826);
nor UO_966 (O_966,N_26488,N_29177);
nand UO_967 (O_967,N_27863,N_29117);
and UO_968 (O_968,N_29288,N_28103);
xor UO_969 (O_969,N_26347,N_25807);
and UO_970 (O_970,N_25844,N_27976);
xnor UO_971 (O_971,N_27412,N_28392);
xnor UO_972 (O_972,N_27788,N_25767);
and UO_973 (O_973,N_28712,N_24136);
nor UO_974 (O_974,N_26073,N_27009);
nor UO_975 (O_975,N_29700,N_29875);
nand UO_976 (O_976,N_29023,N_29534);
xnor UO_977 (O_977,N_25038,N_29663);
nand UO_978 (O_978,N_24104,N_24264);
xnor UO_979 (O_979,N_28527,N_28019);
and UO_980 (O_980,N_28827,N_24336);
nand UO_981 (O_981,N_26150,N_25756);
and UO_982 (O_982,N_24919,N_26779);
nor UO_983 (O_983,N_28488,N_24001);
nor UO_984 (O_984,N_25257,N_29510);
nor UO_985 (O_985,N_25126,N_25285);
and UO_986 (O_986,N_26191,N_27640);
nor UO_987 (O_987,N_28095,N_25294);
and UO_988 (O_988,N_27356,N_25630);
and UO_989 (O_989,N_28282,N_24331);
nor UO_990 (O_990,N_28217,N_27283);
nor UO_991 (O_991,N_28969,N_24867);
nand UO_992 (O_992,N_28308,N_25815);
xor UO_993 (O_993,N_25605,N_25242);
and UO_994 (O_994,N_26854,N_28870);
and UO_995 (O_995,N_27776,N_29181);
and UO_996 (O_996,N_24608,N_26354);
and UO_997 (O_997,N_29347,N_28228);
nand UO_998 (O_998,N_27998,N_24806);
xor UO_999 (O_999,N_29392,N_28032);
or UO_1000 (O_1000,N_24005,N_27573);
xor UO_1001 (O_1001,N_27610,N_26708);
and UO_1002 (O_1002,N_24671,N_24083);
or UO_1003 (O_1003,N_24286,N_27601);
and UO_1004 (O_1004,N_25783,N_24200);
or UO_1005 (O_1005,N_29596,N_26815);
nand UO_1006 (O_1006,N_25373,N_27399);
or UO_1007 (O_1007,N_25288,N_26890);
xnor UO_1008 (O_1008,N_24409,N_26125);
xor UO_1009 (O_1009,N_24149,N_25284);
nor UO_1010 (O_1010,N_29635,N_27086);
xnor UO_1011 (O_1011,N_28049,N_28918);
xnor UO_1012 (O_1012,N_27081,N_27144);
xor UO_1013 (O_1013,N_28836,N_28639);
xor UO_1014 (O_1014,N_29629,N_25556);
or UO_1015 (O_1015,N_29303,N_25993);
nand UO_1016 (O_1016,N_29419,N_27820);
xor UO_1017 (O_1017,N_24797,N_29426);
and UO_1018 (O_1018,N_26839,N_27498);
nand UO_1019 (O_1019,N_25352,N_24295);
nand UO_1020 (O_1020,N_25370,N_25414);
xor UO_1021 (O_1021,N_29904,N_24020);
or UO_1022 (O_1022,N_28605,N_29425);
and UO_1023 (O_1023,N_29896,N_26040);
nor UO_1024 (O_1024,N_25483,N_26895);
nor UO_1025 (O_1025,N_27272,N_27663);
xnor UO_1026 (O_1026,N_24571,N_27578);
and UO_1027 (O_1027,N_26502,N_26982);
xor UO_1028 (O_1028,N_25921,N_28186);
nor UO_1029 (O_1029,N_27721,N_28430);
and UO_1030 (O_1030,N_26455,N_24865);
nand UO_1031 (O_1031,N_27802,N_27291);
xnor UO_1032 (O_1032,N_26172,N_24815);
and UO_1033 (O_1033,N_26830,N_29465);
xnor UO_1034 (O_1034,N_26859,N_29389);
nor UO_1035 (O_1035,N_25833,N_25577);
and UO_1036 (O_1036,N_27490,N_25761);
xor UO_1037 (O_1037,N_29472,N_29100);
or UO_1038 (O_1038,N_25121,N_29421);
nand UO_1039 (O_1039,N_26133,N_25070);
and UO_1040 (O_1040,N_27502,N_25302);
or UO_1041 (O_1041,N_27818,N_26352);
and UO_1042 (O_1042,N_26338,N_26752);
or UO_1043 (O_1043,N_24332,N_27596);
or UO_1044 (O_1044,N_29221,N_29967);
nor UO_1045 (O_1045,N_29806,N_24984);
nand UO_1046 (O_1046,N_25728,N_29174);
nand UO_1047 (O_1047,N_28134,N_28234);
xnor UO_1048 (O_1048,N_24687,N_24918);
and UO_1049 (O_1049,N_28521,N_24627);
nor UO_1050 (O_1050,N_29674,N_24003);
and UO_1051 (O_1051,N_24967,N_29210);
and UO_1052 (O_1052,N_28324,N_25638);
xor UO_1053 (O_1053,N_25061,N_27324);
xnor UO_1054 (O_1054,N_24683,N_24298);
or UO_1055 (O_1055,N_28418,N_24386);
and UO_1056 (O_1056,N_26101,N_24679);
nand UO_1057 (O_1057,N_27332,N_25596);
nor UO_1058 (O_1058,N_29614,N_24446);
nand UO_1059 (O_1059,N_28427,N_27840);
nand UO_1060 (O_1060,N_29976,N_26555);
and UO_1061 (O_1061,N_27000,N_26168);
nand UO_1062 (O_1062,N_25521,N_27106);
nor UO_1063 (O_1063,N_26561,N_27016);
nand UO_1064 (O_1064,N_26418,N_28402);
or UO_1065 (O_1065,N_24036,N_29408);
nand UO_1066 (O_1066,N_27773,N_29440);
nor UO_1067 (O_1067,N_28337,N_29476);
nand UO_1068 (O_1068,N_29298,N_28021);
or UO_1069 (O_1069,N_25922,N_29098);
nor UO_1070 (O_1070,N_26881,N_28258);
xnor UO_1071 (O_1071,N_26165,N_26743);
nor UO_1072 (O_1072,N_26873,N_26781);
and UO_1073 (O_1073,N_28065,N_28687);
xor UO_1074 (O_1074,N_26044,N_29933);
nand UO_1075 (O_1075,N_28820,N_24602);
nand UO_1076 (O_1076,N_29316,N_27850);
and UO_1077 (O_1077,N_26544,N_29342);
nand UO_1078 (O_1078,N_27966,N_25406);
xnor UO_1079 (O_1079,N_24792,N_27169);
nand UO_1080 (O_1080,N_29917,N_25487);
or UO_1081 (O_1081,N_27216,N_24146);
or UO_1082 (O_1082,N_27826,N_28117);
and UO_1083 (O_1083,N_26577,N_24413);
xor UO_1084 (O_1084,N_26941,N_24176);
nor UO_1085 (O_1085,N_26692,N_27938);
or UO_1086 (O_1086,N_27694,N_29987);
nand UO_1087 (O_1087,N_25248,N_29315);
nand UO_1088 (O_1088,N_29194,N_29356);
nand UO_1089 (O_1089,N_28899,N_29466);
nand UO_1090 (O_1090,N_28425,N_25792);
and UO_1091 (O_1091,N_26479,N_24202);
xor UO_1092 (O_1092,N_25928,N_24661);
and UO_1093 (O_1093,N_28432,N_24860);
nand UO_1094 (O_1094,N_28501,N_24425);
nand UO_1095 (O_1095,N_25188,N_29248);
nand UO_1096 (O_1096,N_25941,N_26500);
xor UO_1097 (O_1097,N_29504,N_27585);
nor UO_1098 (O_1098,N_25763,N_29611);
nor UO_1099 (O_1099,N_29283,N_29763);
nand UO_1100 (O_1100,N_29101,N_26914);
xor UO_1101 (O_1101,N_29542,N_24652);
nor UO_1102 (O_1102,N_29434,N_26278);
and UO_1103 (O_1103,N_27763,N_24814);
or UO_1104 (O_1104,N_24799,N_27615);
nor UO_1105 (O_1105,N_29468,N_25827);
nand UO_1106 (O_1106,N_27095,N_25232);
xor UO_1107 (O_1107,N_28708,N_29158);
and UO_1108 (O_1108,N_25462,N_28515);
nand UO_1109 (O_1109,N_26901,N_27549);
nand UO_1110 (O_1110,N_25356,N_28449);
or UO_1111 (O_1111,N_24137,N_25738);
xnor UO_1112 (O_1112,N_25520,N_28310);
nor UO_1113 (O_1113,N_25206,N_25316);
or UO_1114 (O_1114,N_25186,N_27234);
and UO_1115 (O_1115,N_24330,N_29554);
and UO_1116 (O_1116,N_29436,N_25404);
and UO_1117 (O_1117,N_24151,N_24557);
and UO_1118 (O_1118,N_29624,N_27302);
or UO_1119 (O_1119,N_28766,N_24221);
xor UO_1120 (O_1120,N_29147,N_29686);
nor UO_1121 (O_1121,N_26648,N_28675);
and UO_1122 (O_1122,N_24531,N_24508);
and UO_1123 (O_1123,N_24680,N_26537);
nand UO_1124 (O_1124,N_27823,N_27256);
nand UO_1125 (O_1125,N_29888,N_28700);
xnor UO_1126 (O_1126,N_24034,N_26206);
or UO_1127 (O_1127,N_24012,N_29065);
xor UO_1128 (O_1128,N_25233,N_27126);
and UO_1129 (O_1129,N_26654,N_28099);
xor UO_1130 (O_1130,N_28843,N_26434);
and UO_1131 (O_1131,N_27346,N_26559);
xor UO_1132 (O_1132,N_24750,N_27413);
nor UO_1133 (O_1133,N_28591,N_25189);
xor UO_1134 (O_1134,N_24396,N_29062);
and UO_1135 (O_1135,N_28930,N_24458);
or UO_1136 (O_1136,N_27747,N_26069);
or UO_1137 (O_1137,N_25218,N_28476);
xor UO_1138 (O_1138,N_27766,N_28704);
xnor UO_1139 (O_1139,N_27068,N_25768);
nand UO_1140 (O_1140,N_29847,N_26248);
or UO_1141 (O_1141,N_25537,N_27391);
xnor UO_1142 (O_1142,N_27806,N_25604);
xnor UO_1143 (O_1143,N_24478,N_26661);
and UO_1144 (O_1144,N_27470,N_25804);
nor UO_1145 (O_1145,N_25830,N_27015);
xnor UO_1146 (O_1146,N_28241,N_26023);
and UO_1147 (O_1147,N_24197,N_28683);
or UO_1148 (O_1148,N_29019,N_26509);
nand UO_1149 (O_1149,N_24646,N_27547);
and UO_1150 (O_1150,N_24949,N_25313);
and UO_1151 (O_1151,N_27778,N_27664);
and UO_1152 (O_1152,N_26823,N_25407);
nand UO_1153 (O_1153,N_26045,N_28902);
nor UO_1154 (O_1154,N_24275,N_29066);
nor UO_1155 (O_1155,N_27881,N_27913);
and UO_1156 (O_1156,N_26693,N_26922);
and UO_1157 (O_1157,N_24612,N_26173);
and UO_1158 (O_1158,N_26836,N_28112);
xor UO_1159 (O_1159,N_27238,N_27710);
nand UO_1160 (O_1160,N_29793,N_29021);
nor UO_1161 (O_1161,N_26429,N_27811);
nand UO_1162 (O_1162,N_29597,N_29655);
xnor UO_1163 (O_1163,N_24302,N_28917);
or UO_1164 (O_1164,N_28485,N_28999);
or UO_1165 (O_1165,N_29761,N_29854);
nand UO_1166 (O_1166,N_29152,N_26412);
nor UO_1167 (O_1167,N_29988,N_29733);
nor UO_1168 (O_1168,N_29821,N_27837);
nor UO_1169 (O_1169,N_24063,N_25148);
nor UO_1170 (O_1170,N_25042,N_25622);
nand UO_1171 (O_1171,N_24472,N_25598);
and UO_1172 (O_1172,N_24768,N_28977);
or UO_1173 (O_1173,N_28120,N_28287);
and UO_1174 (O_1174,N_27821,N_24338);
nand UO_1175 (O_1175,N_25549,N_29120);
xor UO_1176 (O_1176,N_24530,N_25651);
and UO_1177 (O_1177,N_29849,N_28895);
xnor UO_1178 (O_1178,N_28444,N_25772);
xor UO_1179 (O_1179,N_25505,N_29837);
xnor UO_1180 (O_1180,N_27157,N_24268);
xor UO_1181 (O_1181,N_28301,N_26260);
nand UO_1182 (O_1182,N_24444,N_26762);
xor UO_1183 (O_1183,N_27569,N_28160);
xor UO_1184 (O_1184,N_25023,N_27542);
nor UO_1185 (O_1185,N_26414,N_26799);
and UO_1186 (O_1186,N_28728,N_24717);
nand UO_1187 (O_1187,N_26959,N_25593);
or UO_1188 (O_1188,N_25149,N_25009);
nor UO_1189 (O_1189,N_29140,N_28022);
nand UO_1190 (O_1190,N_28455,N_27058);
nand UO_1191 (O_1191,N_25120,N_27861);
nor UO_1192 (O_1192,N_29815,N_29945);
and UO_1193 (O_1193,N_28426,N_28096);
xnor UO_1194 (O_1194,N_27384,N_26887);
nand UO_1195 (O_1195,N_27211,N_24488);
nand UO_1196 (O_1196,N_29483,N_24263);
and UO_1197 (O_1197,N_27474,N_24008);
or UO_1198 (O_1198,N_26939,N_29922);
nor UO_1199 (O_1199,N_27453,N_25594);
xnor UO_1200 (O_1200,N_25274,N_29690);
nand UO_1201 (O_1201,N_29344,N_27503);
xor UO_1202 (O_1202,N_29850,N_28599);
or UO_1203 (O_1203,N_27808,N_26514);
or UO_1204 (O_1204,N_26619,N_25421);
nand UO_1205 (O_1205,N_26607,N_25300);
xnor UO_1206 (O_1206,N_29930,N_29369);
nand UO_1207 (O_1207,N_28571,N_29346);
and UO_1208 (O_1208,N_25336,N_28886);
and UO_1209 (O_1209,N_25191,N_25354);
xor UO_1210 (O_1210,N_24212,N_26651);
nand UO_1211 (O_1211,N_29578,N_26064);
and UO_1212 (O_1212,N_29270,N_28962);
xnor UO_1213 (O_1213,N_29481,N_29513);
xor UO_1214 (O_1214,N_25595,N_27819);
and UO_1215 (O_1215,N_28041,N_24755);
and UO_1216 (O_1216,N_29041,N_29139);
nand UO_1217 (O_1217,N_27362,N_28538);
xor UO_1218 (O_1218,N_27504,N_29791);
and UO_1219 (O_1219,N_24255,N_24994);
and UO_1220 (O_1220,N_28879,N_27739);
or UO_1221 (O_1221,N_28554,N_28066);
and UO_1222 (O_1222,N_25939,N_25988);
xor UO_1223 (O_1223,N_29154,N_26473);
or UO_1224 (O_1224,N_24565,N_26685);
and UO_1225 (O_1225,N_24706,N_27654);
or UO_1226 (O_1226,N_24447,N_27066);
nor UO_1227 (O_1227,N_25723,N_27520);
xnor UO_1228 (O_1228,N_29128,N_26591);
or UO_1229 (O_1229,N_29703,N_26589);
xor UO_1230 (O_1230,N_26545,N_29003);
and UO_1231 (O_1231,N_25627,N_25555);
nand UO_1232 (O_1232,N_25154,N_27201);
and UO_1233 (O_1233,N_29530,N_27003);
nand UO_1234 (O_1234,N_29802,N_24590);
and UO_1235 (O_1235,N_25980,N_29678);
and UO_1236 (O_1236,N_24131,N_27707);
xor UO_1237 (O_1237,N_26620,N_26734);
nor UO_1238 (O_1238,N_27561,N_24875);
and UO_1239 (O_1239,N_27321,N_27962);
nand UO_1240 (O_1240,N_29172,N_28757);
or UO_1241 (O_1241,N_24591,N_24629);
xnor UO_1242 (O_1242,N_24564,N_24497);
or UO_1243 (O_1243,N_29081,N_26154);
nor UO_1244 (O_1244,N_28409,N_29801);
and UO_1245 (O_1245,N_24468,N_28250);
xor UO_1246 (O_1246,N_26554,N_28462);
or UO_1247 (O_1247,N_29319,N_26973);
xor UO_1248 (O_1248,N_28297,N_25740);
xor UO_1249 (O_1249,N_27050,N_26642);
xnor UO_1250 (O_1250,N_28436,N_27681);
or UO_1251 (O_1251,N_26727,N_29520);
and UO_1252 (O_1252,N_25703,N_29727);
xnor UO_1253 (O_1253,N_26751,N_26746);
nand UO_1254 (O_1254,N_26082,N_26014);
xor UO_1255 (O_1255,N_28558,N_28171);
xor UO_1256 (O_1256,N_24374,N_27866);
or UO_1257 (O_1257,N_26520,N_29573);
and UO_1258 (O_1258,N_27331,N_26893);
xnor UO_1259 (O_1259,N_24031,N_25645);
or UO_1260 (O_1260,N_27196,N_24142);
nor UO_1261 (O_1261,N_29575,N_24132);
nor UO_1262 (O_1262,N_27342,N_26849);
or UO_1263 (O_1263,N_27900,N_25828);
nand UO_1264 (O_1264,N_24178,N_24272);
xor UO_1265 (O_1265,N_25398,N_29639);
nor UO_1266 (O_1266,N_24515,N_24934);
xnor UO_1267 (O_1267,N_28579,N_26090);
and UO_1268 (O_1268,N_27500,N_28573);
xnor UO_1269 (O_1269,N_25139,N_27875);
and UO_1270 (O_1270,N_26241,N_27674);
xnor UO_1271 (O_1271,N_27530,N_28889);
or UO_1272 (O_1272,N_24243,N_29293);
nor UO_1273 (O_1273,N_29124,N_28178);
nand UO_1274 (O_1274,N_26930,N_29566);
xor UO_1275 (O_1275,N_24213,N_29613);
xor UO_1276 (O_1276,N_25774,N_29689);
xnor UO_1277 (O_1277,N_26512,N_27322);
or UO_1278 (O_1278,N_28763,N_27260);
nor UO_1279 (O_1279,N_26393,N_25321);
or UO_1280 (O_1280,N_26041,N_28944);
and UO_1281 (O_1281,N_29676,N_25159);
or UO_1282 (O_1282,N_26627,N_26170);
or UO_1283 (O_1283,N_28799,N_29413);
or UO_1284 (O_1284,N_27872,N_28600);
or UO_1285 (O_1285,N_27864,N_26240);
and UO_1286 (O_1286,N_29618,N_27948);
xnor UO_1287 (O_1287,N_27959,N_26288);
nor UO_1288 (O_1288,N_27394,N_27991);
and UO_1289 (O_1289,N_26821,N_29946);
and UO_1290 (O_1290,N_28385,N_28082);
xnor UO_1291 (O_1291,N_27612,N_25940);
or UO_1292 (O_1292,N_26203,N_29273);
nor UO_1293 (O_1293,N_29825,N_25974);
nor UO_1294 (O_1294,N_26120,N_28614);
xor UO_1295 (O_1295,N_27273,N_29993);
nor UO_1296 (O_1296,N_29028,N_25394);
and UO_1297 (O_1297,N_27259,N_24387);
nand UO_1298 (O_1298,N_26865,N_26719);
nor UO_1299 (O_1299,N_29189,N_25575);
xor UO_1300 (O_1300,N_27078,N_28121);
xnor UO_1301 (O_1301,N_24130,N_27658);
or UO_1302 (O_1302,N_29422,N_27208);
or UO_1303 (O_1303,N_29043,N_28502);
nand UO_1304 (O_1304,N_24273,N_27446);
and UO_1305 (O_1305,N_24845,N_29220);
nor UO_1306 (O_1306,N_28458,N_29134);
nand UO_1307 (O_1307,N_24234,N_27269);
or UO_1308 (O_1308,N_28894,N_25276);
nand UO_1309 (O_1309,N_26538,N_28747);
and UO_1310 (O_1310,N_24641,N_25348);
nor UO_1311 (O_1311,N_27103,N_27918);
nand UO_1312 (O_1312,N_25162,N_26932);
xnor UO_1313 (O_1313,N_29379,N_25777);
or UO_1314 (O_1314,N_24822,N_27263);
nand UO_1315 (O_1315,N_24105,N_27577);
nand UO_1316 (O_1316,N_29529,N_24297);
nand UO_1317 (O_1317,N_28919,N_27409);
xor UO_1318 (O_1318,N_29942,N_25205);
nand UO_1319 (O_1319,N_29024,N_26483);
and UO_1320 (O_1320,N_24893,N_26435);
or UO_1321 (O_1321,N_27154,N_28179);
nor UO_1322 (O_1322,N_27014,N_29656);
nand UO_1323 (O_1323,N_25440,N_28111);
xnor UO_1324 (O_1324,N_24011,N_27761);
and UO_1325 (O_1325,N_26458,N_24697);
xnor UO_1326 (O_1326,N_26850,N_29363);
and UO_1327 (O_1327,N_26316,N_25140);
nor UO_1328 (O_1328,N_28574,N_27713);
nor UO_1329 (O_1329,N_26123,N_28472);
and UO_1330 (O_1330,N_26528,N_28824);
xor UO_1331 (O_1331,N_24499,N_25307);
xnor UO_1332 (O_1332,N_28494,N_29146);
nand UO_1333 (O_1333,N_24828,N_25580);
nand UO_1334 (O_1334,N_24947,N_25977);
and UO_1335 (O_1335,N_25737,N_29045);
nor UO_1336 (O_1336,N_26573,N_29926);
or UO_1337 (O_1337,N_25861,N_28569);
and UO_1338 (O_1338,N_26638,N_28480);
nand UO_1339 (O_1339,N_25872,N_24659);
or UO_1340 (O_1340,N_28932,N_24090);
xor UO_1341 (O_1341,N_26462,N_24963);
nor UO_1342 (O_1342,N_28963,N_27288);
and UO_1343 (O_1343,N_27758,N_25693);
and UO_1344 (O_1344,N_24241,N_25529);
or UO_1345 (O_1345,N_26236,N_29095);
or UO_1346 (O_1346,N_24509,N_28352);
nor UO_1347 (O_1347,N_26892,N_25717);
nand UO_1348 (O_1348,N_25579,N_24972);
xor UO_1349 (O_1349,N_24569,N_29069);
or UO_1350 (O_1350,N_27733,N_28150);
or UO_1351 (O_1351,N_24198,N_28174);
nand UO_1352 (O_1352,N_25111,N_28489);
xor UO_1353 (O_1353,N_27062,N_28823);
or UO_1354 (O_1354,N_26162,N_29165);
xnor UO_1355 (O_1355,N_24207,N_28443);
or UO_1356 (O_1356,N_28153,N_24847);
nand UO_1357 (O_1357,N_29203,N_24400);
nand UO_1358 (O_1358,N_28421,N_26675);
or UO_1359 (O_1359,N_29898,N_27065);
nand UO_1360 (O_1360,N_26039,N_25114);
nor UO_1361 (O_1361,N_25476,N_29762);
xnor UO_1362 (O_1362,N_26421,N_29008);
xnor UO_1363 (O_1363,N_29428,N_29320);
and UO_1364 (O_1364,N_25299,N_25951);
and UO_1365 (O_1365,N_24397,N_27912);
nor UO_1366 (O_1366,N_26249,N_27657);
and UO_1367 (O_1367,N_27159,N_25550);
and UO_1368 (O_1368,N_29222,N_29193);
nor UO_1369 (O_1369,N_29108,N_24794);
xor UO_1370 (O_1370,N_24944,N_26725);
nor UO_1371 (O_1371,N_26774,N_25236);
or UO_1372 (O_1372,N_28604,N_25385);
nor UO_1373 (O_1373,N_29918,N_29355);
or UO_1374 (O_1374,N_26431,N_24909);
xor UO_1375 (O_1375,N_28656,N_27162);
or UO_1376 (O_1376,N_25710,N_26043);
or UO_1377 (O_1377,N_24605,N_27055);
or UO_1378 (O_1378,N_24922,N_26185);
or UO_1379 (O_1379,N_27110,N_24248);
and UO_1380 (O_1380,N_25161,N_26063);
nand UO_1381 (O_1381,N_25339,N_27880);
nand UO_1382 (O_1382,N_24024,N_27907);
and UO_1383 (O_1383,N_27884,N_29429);
and UO_1384 (O_1384,N_26319,N_25376);
nor UO_1385 (O_1385,N_26489,N_29819);
and UO_1386 (O_1386,N_24296,N_29687);
nand UO_1387 (O_1387,N_26657,N_28659);
xnor UO_1388 (O_1388,N_29305,N_28475);
nor UO_1389 (O_1389,N_25393,N_28190);
nand UO_1390 (O_1390,N_26459,N_25970);
nand UO_1391 (O_1391,N_24688,N_27637);
or UO_1392 (O_1392,N_25375,N_27128);
and UO_1393 (O_1393,N_25641,N_25655);
and UO_1394 (O_1394,N_26061,N_28320);
nand UO_1395 (O_1395,N_24753,N_26868);
xor UO_1396 (O_1396,N_27210,N_24506);
nor UO_1397 (O_1397,N_29669,N_25455);
or UO_1398 (O_1398,N_29657,N_28553);
or UO_1399 (O_1399,N_24831,N_28692);
or UO_1400 (O_1400,N_27164,N_24196);
nand UO_1401 (O_1401,N_26355,N_24846);
and UO_1402 (O_1402,N_25176,N_26272);
nand UO_1403 (O_1403,N_29442,N_27372);
nor UO_1404 (O_1404,N_27069,N_26931);
nor UO_1405 (O_1405,N_26566,N_25620);
or UO_1406 (O_1406,N_25720,N_26546);
xnor UO_1407 (O_1407,N_28832,N_28989);
and UO_1408 (O_1408,N_29748,N_24862);
and UO_1409 (O_1409,N_28913,N_26791);
nor UO_1410 (O_1410,N_26557,N_29002);
and UO_1411 (O_1411,N_25915,N_28270);
or UO_1412 (O_1412,N_27113,N_26190);
nand UO_1413 (O_1413,N_25342,N_28561);
and UO_1414 (O_1414,N_28539,N_27737);
or UO_1415 (O_1415,N_27684,N_29519);
and UO_1416 (O_1416,N_26343,N_25387);
and UO_1417 (O_1417,N_29913,N_29715);
and UO_1418 (O_1418,N_29004,N_27606);
or UO_1419 (O_1419,N_25654,N_27145);
xor UO_1420 (O_1420,N_24089,N_28546);
and UO_1421 (O_1421,N_25791,N_27468);
nor UO_1422 (O_1422,N_28029,N_24100);
or UO_1423 (O_1423,N_26891,N_24813);
and UO_1424 (O_1424,N_28343,N_28802);
xnor UO_1425 (O_1425,N_24076,N_26820);
or UO_1426 (O_1426,N_24098,N_25787);
and UO_1427 (O_1427,N_25864,N_24663);
nand UO_1428 (O_1428,N_25101,N_28522);
or UO_1429 (O_1429,N_24239,N_28326);
and UO_1430 (O_1430,N_27683,N_27715);
xor UO_1431 (O_1431,N_27860,N_28568);
nor UO_1432 (O_1432,N_26872,N_24004);
xnor UO_1433 (O_1433,N_29354,N_25831);
or UO_1434 (O_1434,N_28446,N_24927);
and UO_1435 (O_1435,N_24937,N_25143);
xor UO_1436 (O_1436,N_26285,N_27021);
nor UO_1437 (O_1437,N_28118,N_29414);
xor UO_1438 (O_1438,N_24853,N_25074);
nand UO_1439 (O_1439,N_24249,N_26866);
and UO_1440 (O_1440,N_24322,N_28860);
or UO_1441 (O_1441,N_27056,N_27961);
xnor UO_1442 (O_1442,N_27286,N_24418);
xor UO_1443 (O_1443,N_27097,N_29280);
xnor UO_1444 (O_1444,N_24522,N_29548);
nand UO_1445 (O_1445,N_24789,N_28239);
xnor UO_1446 (O_1446,N_27115,N_24053);
or UO_1447 (O_1447,N_28498,N_29006);
and UO_1448 (O_1448,N_24666,N_28622);
xor UO_1449 (O_1449,N_26644,N_26717);
xor UO_1450 (O_1450,N_26641,N_25502);
and UO_1451 (O_1451,N_25619,N_25909);
or UO_1452 (O_1452,N_24917,N_28547);
and UO_1453 (O_1453,N_24385,N_29889);
xnor UO_1454 (O_1454,N_26152,N_28684);
nor UO_1455 (O_1455,N_25795,N_24991);
nand UO_1456 (O_1456,N_28742,N_29652);
xnor UO_1457 (O_1457,N_24587,N_29615);
xnor UO_1458 (O_1458,N_25325,N_28353);
nand UO_1459 (O_1459,N_25454,N_28750);
or UO_1460 (O_1460,N_25109,N_26764);
nor UO_1461 (O_1461,N_27908,N_26374);
or UO_1462 (O_1462,N_29227,N_27044);
nand UO_1463 (O_1463,N_24058,N_28943);
nor UO_1464 (O_1464,N_24175,N_26371);
and UO_1465 (O_1465,N_28100,N_24359);
or UO_1466 (O_1466,N_24000,N_29953);
and UO_1467 (O_1467,N_25326,N_27598);
and UO_1468 (O_1468,N_28439,N_28300);
nand UO_1469 (O_1469,N_28576,N_24892);
xnor UO_1470 (O_1470,N_24929,N_24637);
and UO_1471 (O_1471,N_28119,N_28903);
nand UO_1472 (O_1472,N_25524,N_29044);
and UO_1473 (O_1473,N_24394,N_29125);
nor UO_1474 (O_1474,N_26793,N_27693);
nor UO_1475 (O_1475,N_25916,N_29300);
and UO_1476 (O_1476,N_24834,N_25089);
nor UO_1477 (O_1477,N_29587,N_27466);
nand UO_1478 (O_1478,N_28634,N_27630);
nor UO_1479 (O_1479,N_28643,N_29627);
and UO_1480 (O_1480,N_28564,N_25679);
nor UO_1481 (O_1481,N_24974,N_28158);
and UO_1482 (O_1482,N_28718,N_28951);
xor UO_1483 (O_1483,N_25287,N_28984);
and UO_1484 (O_1484,N_29384,N_25310);
nor UO_1485 (O_1485,N_26851,N_26171);
xor UO_1486 (O_1486,N_28373,N_29959);
or UO_1487 (O_1487,N_25699,N_27536);
nor UO_1488 (O_1488,N_28252,N_27160);
nor UO_1489 (O_1489,N_26916,N_26046);
nand UO_1490 (O_1490,N_26379,N_28607);
or UO_1491 (O_1491,N_27213,N_25923);
and UO_1492 (O_1492,N_28927,N_25221);
nor UO_1493 (O_1493,N_26096,N_27206);
xor UO_1494 (O_1494,N_24430,N_25478);
or UO_1495 (O_1495,N_25790,N_27687);
xnor UO_1496 (O_1496,N_27647,N_28360);
or UO_1497 (O_1497,N_27105,N_26726);
or UO_1498 (O_1498,N_24064,N_27832);
xor UO_1499 (O_1499,N_29911,N_26749);
or UO_1500 (O_1500,N_24471,N_28394);
xor UO_1501 (O_1501,N_29479,N_26917);
or UO_1502 (O_1502,N_29972,N_28761);
xor UO_1503 (O_1503,N_27345,N_24581);
nand UO_1504 (O_1504,N_28746,N_25551);
xnor UO_1505 (O_1505,N_25056,N_28651);
and UO_1506 (O_1506,N_24319,N_28988);
xor UO_1507 (O_1507,N_28601,N_28420);
or UO_1508 (O_1508,N_29540,N_24607);
nor UO_1509 (O_1509,N_27714,N_26533);
or UO_1510 (O_1510,N_28867,N_28512);
or UO_1511 (O_1511,N_29460,N_29606);
xor UO_1512 (O_1512,N_24116,N_26721);
nor UO_1513 (O_1513,N_26523,N_25408);
and UO_1514 (O_1514,N_26813,N_26169);
xnor UO_1515 (O_1515,N_25156,N_26632);
and UO_1516 (O_1516,N_28633,N_27855);
xnor UO_1517 (O_1517,N_29430,N_28183);
nor UO_1518 (O_1518,N_28544,N_26621);
nor UO_1519 (O_1519,N_29921,N_25007);
nand UO_1520 (O_1520,N_25223,N_26438);
xor UO_1521 (O_1521,N_28139,N_26318);
or UO_1522 (O_1522,N_29470,N_27436);
or UO_1523 (O_1523,N_26847,N_28344);
nor UO_1524 (O_1524,N_25481,N_28667);
nand UO_1525 (O_1525,N_28238,N_25797);
nand UO_1526 (O_1526,N_25137,N_27315);
nor UO_1527 (O_1527,N_24133,N_28749);
and UO_1528 (O_1528,N_27072,N_24038);
nor UO_1529 (O_1529,N_26128,N_25127);
xnor UO_1530 (O_1530,N_26667,N_28341);
and UO_1531 (O_1531,N_27921,N_27276);
xnor UO_1532 (O_1532,N_29334,N_25345);
nand UO_1533 (O_1533,N_26059,N_24074);
nand UO_1534 (O_1534,N_27017,N_25102);
nand UO_1535 (O_1535,N_26631,N_28876);
xnor UO_1536 (O_1536,N_24158,N_27368);
and UO_1537 (O_1537,N_25275,N_26389);
and UO_1538 (O_1538,N_29435,N_29239);
nand UO_1539 (O_1539,N_25066,N_29000);
or UO_1540 (O_1540,N_24265,N_24152);
or UO_1541 (O_1541,N_25871,N_27876);
and UO_1542 (O_1542,N_25444,N_24078);
and UO_1543 (O_1543,N_25934,N_24411);
xnor UO_1544 (O_1544,N_26548,N_28790);
xor UO_1545 (O_1545,N_28030,N_28777);
or UO_1546 (O_1546,N_26383,N_24567);
nor UO_1547 (O_1547,N_28754,N_29955);
or UO_1548 (O_1548,N_24168,N_27970);
nor UO_1549 (O_1549,N_25019,N_28674);
and UO_1550 (O_1550,N_26359,N_29527);
xor UO_1551 (O_1551,N_27628,N_28422);
or UO_1552 (O_1552,N_25157,N_26084);
or UO_1553 (O_1553,N_25416,N_26103);
nor UO_1554 (O_1554,N_29576,N_26247);
nor UO_1555 (O_1555,N_28817,N_28358);
or UO_1556 (O_1556,N_27853,N_27562);
nor UO_1557 (O_1557,N_29681,N_27166);
and UO_1558 (O_1558,N_24819,N_25277);
and UO_1559 (O_1559,N_27411,N_28552);
and UO_1560 (O_1560,N_27807,N_26217);
nor UO_1561 (O_1561,N_29670,N_28347);
and UO_1562 (O_1562,N_25810,N_28526);
or UO_1563 (O_1563,N_28826,N_24410);
nor UO_1564 (O_1564,N_29914,N_25343);
and UO_1565 (O_1565,N_26257,N_26018);
and UO_1566 (O_1566,N_29923,N_25123);
or UO_1567 (O_1567,N_28437,N_24481);
or UO_1568 (O_1568,N_29555,N_26452);
or UO_1569 (O_1569,N_24665,N_24305);
xor UO_1570 (O_1570,N_27688,N_29402);
xnor UO_1571 (O_1571,N_25911,N_28891);
and UO_1572 (O_1572,N_25572,N_29133);
or UO_1573 (O_1573,N_24230,N_29759);
xnor UO_1574 (O_1574,N_24218,N_29486);
xor UO_1575 (O_1575,N_25901,N_24734);
xor UO_1576 (O_1576,N_25024,N_26358);
xnor UO_1577 (O_1577,N_25413,N_25254);
nand UO_1578 (O_1578,N_27023,N_27696);
and UO_1579 (O_1579,N_25601,N_27439);
nand UO_1580 (O_1580,N_25001,N_24006);
nand UO_1581 (O_1581,N_29532,N_27108);
or UO_1582 (O_1582,N_26237,N_28854);
nand UO_1583 (O_1583,N_25237,N_28597);
nand UO_1584 (O_1584,N_29990,N_28492);
xor UO_1585 (O_1585,N_28005,N_25113);
nand UO_1586 (O_1586,N_24585,N_27960);
or UO_1587 (O_1587,N_28580,N_25182);
xnor UO_1588 (O_1588,N_27274,N_24879);
or UO_1589 (O_1589,N_28256,N_26054);
nor UO_1590 (O_1590,N_27217,N_29982);
or UO_1591 (O_1591,N_25442,N_26229);
nand UO_1592 (O_1592,N_27904,N_27844);
nand UO_1593 (O_1593,N_25361,N_27277);
and UO_1594 (O_1594,N_26587,N_26608);
and UO_1595 (O_1595,N_29675,N_24621);
or UO_1596 (O_1596,N_28537,N_28225);
xor UO_1597 (O_1597,N_25399,N_27515);
xnor UO_1598 (O_1598,N_26508,N_29012);
xor UO_1599 (O_1599,N_26669,N_24427);
or UO_1600 (O_1600,N_27967,N_29474);
and UO_1601 (O_1601,N_28274,N_27894);
xor UO_1602 (O_1602,N_28565,N_27494);
xor UO_1603 (O_1603,N_25445,N_26879);
nor UO_1604 (O_1604,N_24379,N_24086);
nor UO_1605 (O_1605,N_27423,N_24217);
or UO_1606 (O_1606,N_25115,N_25415);
xnor UO_1607 (O_1607,N_27491,N_28069);
nand UO_1608 (O_1608,N_27718,N_28155);
or UO_1609 (O_1609,N_24849,N_26065);
nand UO_1610 (O_1610,N_26244,N_28859);
nand UO_1611 (O_1611,N_28949,N_26776);
xor UO_1612 (O_1612,N_29528,N_24293);
and UO_1613 (O_1613,N_29448,N_26463);
or UO_1614 (O_1614,N_27621,N_25878);
xnor UO_1615 (O_1615,N_25039,N_25764);
xnor UO_1616 (O_1616,N_25388,N_26302);
nand UO_1617 (O_1617,N_27483,N_27755);
xor UO_1618 (O_1618,N_26493,N_25461);
xor UO_1619 (O_1619,N_27462,N_29820);
or UO_1620 (O_1620,N_24576,N_27374);
nand UO_1621 (O_1621,N_26663,N_29050);
or UO_1622 (O_1622,N_24655,N_27158);
xnor UO_1623 (O_1623,N_26496,N_29089);
or UO_1624 (O_1624,N_29764,N_29450);
and UO_1625 (O_1625,N_26733,N_26094);
or UO_1626 (O_1626,N_24650,N_25771);
nor UO_1627 (O_1627,N_25891,N_28830);
and UO_1628 (O_1628,N_29321,N_24326);
and UO_1629 (O_1629,N_25418,N_25344);
nand UO_1630 (O_1630,N_28383,N_26753);
nand UO_1631 (O_1631,N_25875,N_25866);
xnor UO_1632 (O_1632,N_26967,N_27240);
and UO_1633 (O_1633,N_27328,N_25308);
xor UO_1634 (O_1634,N_24483,N_27427);
nand UO_1635 (O_1635,N_28164,N_26360);
nor UO_1636 (O_1636,N_26423,N_26336);
and UO_1637 (O_1637,N_29609,N_25812);
nor UO_1638 (O_1638,N_24118,N_29257);
nand UO_1639 (O_1639,N_28043,N_29539);
nor UO_1640 (O_1640,N_24161,N_26822);
nor UO_1641 (O_1641,N_29620,N_24951);
and UO_1642 (O_1642,N_26187,N_29323);
nor UO_1643 (O_1643,N_27898,N_25796);
and UO_1644 (O_1644,N_25320,N_28892);
xor UO_1645 (O_1645,N_28401,N_27163);
nor UO_1646 (O_1646,N_27476,N_28460);
xnor UO_1647 (O_1647,N_28967,N_24214);
or UO_1648 (O_1648,N_27632,N_25334);
nand UO_1649 (O_1649,N_25105,N_29034);
xnor UO_1650 (O_1650,N_24457,N_28098);
nor UO_1651 (O_1651,N_27035,N_28292);
and UO_1652 (O_1652,N_25204,N_26232);
or UO_1653 (O_1653,N_26938,N_28464);
nand UO_1654 (O_1654,N_29705,N_26532);
nand UO_1655 (O_1655,N_29277,N_26568);
xor UO_1656 (O_1656,N_24635,N_25168);
xnor UO_1657 (O_1657,N_29830,N_25095);
xnor UO_1658 (O_1658,N_28713,N_24081);
xor UO_1659 (O_1659,N_28803,N_27385);
nor UO_1660 (O_1660,N_26072,N_29565);
or UO_1661 (O_1661,N_28540,N_27172);
and UO_1662 (O_1662,N_26697,N_27887);
nand UO_1663 (O_1663,N_28901,N_28267);
nor UO_1664 (O_1664,N_25918,N_27287);
or UO_1665 (O_1665,N_25020,N_27619);
xnor UO_1666 (O_1666,N_24620,N_28839);
or UO_1667 (O_1667,N_29339,N_24859);
and UO_1668 (O_1668,N_28104,N_25589);
nand UO_1669 (O_1669,N_29863,N_28596);
nor UO_1670 (O_1670,N_27390,N_27122);
and UO_1671 (O_1671,N_29463,N_25669);
and UO_1672 (O_1672,N_27478,N_28281);
or UO_1673 (O_1673,N_24490,N_25309);
or UO_1674 (O_1674,N_29403,N_24573);
xor UO_1675 (O_1675,N_27946,N_24964);
or UO_1676 (O_1676,N_27309,N_24120);
and UO_1677 (O_1677,N_25868,N_27430);
and UO_1678 (O_1678,N_24651,N_26113);
nand UO_1679 (O_1679,N_26705,N_28251);
nor UO_1680 (O_1680,N_27525,N_26250);
nand UO_1681 (O_1681,N_27343,N_24194);
and UO_1682 (O_1682,N_25753,N_29897);
nand UO_1683 (O_1683,N_29915,N_26598);
and UO_1684 (O_1684,N_28016,N_24442);
and UO_1685 (O_1685,N_27225,N_25648);
or UO_1686 (O_1686,N_26401,N_25966);
and UO_1687 (O_1687,N_24422,N_28233);
xor UO_1688 (O_1688,N_29865,N_26806);
or UO_1689 (O_1689,N_27048,N_24491);
nand UO_1690 (O_1690,N_25786,N_29750);
nor UO_1691 (O_1691,N_26772,N_27487);
or UO_1692 (O_1692,N_25467,N_27053);
xor UO_1693 (O_1693,N_26658,N_25682);
or UO_1694 (O_1694,N_28127,N_25358);
nor UO_1695 (O_1695,N_26076,N_24582);
nand UO_1696 (O_1696,N_26684,N_27971);
xnor UO_1697 (O_1697,N_28534,N_25093);
xor UO_1698 (O_1698,N_25742,N_27560);
nand UO_1699 (O_1699,N_29640,N_27085);
or UO_1700 (O_1700,N_25044,N_24087);
or UO_1701 (O_1701,N_26074,N_26397);
xnor UO_1702 (O_1702,N_25724,N_28248);
or UO_1703 (O_1703,N_24953,N_26905);
or UO_1704 (O_1704,N_28325,N_27006);
or UO_1705 (O_1705,N_29444,N_29475);
or UO_1706 (O_1706,N_24864,N_24640);
and UO_1707 (O_1707,N_24093,N_26649);
or UO_1708 (O_1708,N_24127,N_27136);
xnor UO_1709 (O_1709,N_26188,N_29991);
and UO_1710 (O_1710,N_29795,N_28804);
or UO_1711 (O_1711,N_26027,N_26086);
or UO_1712 (O_1712,N_29997,N_27073);
nand UO_1713 (O_1713,N_29730,N_27012);
or UO_1714 (O_1714,N_25133,N_24623);
nor UO_1715 (O_1715,N_28997,N_25036);
nor UO_1716 (O_1716,N_29800,N_29178);
nor UO_1717 (O_1717,N_29374,N_27395);
and UO_1718 (O_1718,N_28856,N_25364);
xnor UO_1719 (O_1719,N_24610,N_26731);
xor UO_1720 (O_1720,N_26021,N_26558);
nand UO_1721 (O_1721,N_26332,N_24938);
and UO_1722 (O_1722,N_26144,N_25201);
and UO_1723 (O_1723,N_25460,N_25752);
nor UO_1724 (O_1724,N_29760,N_24724);
and UO_1725 (O_1725,N_28181,N_26478);
or UO_1726 (O_1726,N_26594,N_24463);
and UO_1727 (O_1727,N_25411,N_29467);
xor UO_1728 (O_1728,N_27935,N_25696);
and UO_1729 (O_1729,N_24270,N_29001);
or UO_1730 (O_1730,N_28904,N_24749);
or UO_1731 (O_1731,N_27425,N_28928);
nor UO_1732 (O_1732,N_28755,N_26197);
nand UO_1733 (O_1733,N_26056,N_24636);
nor UO_1734 (O_1734,N_25367,N_25069);
nand UO_1735 (O_1735,N_24701,N_25642);
or UO_1736 (O_1736,N_28400,N_28089);
xor UO_1737 (O_1737,N_29224,N_24252);
or UO_1738 (O_1738,N_28776,N_25050);
nor UO_1739 (O_1739,N_27511,N_24310);
and UO_1740 (O_1740,N_24968,N_29841);
or UO_1741 (O_1741,N_29161,N_24345);
and UO_1742 (O_1742,N_27782,N_25722);
or UO_1743 (O_1743,N_26802,N_25775);
xnor UO_1744 (O_1744,N_25231,N_29619);
or UO_1745 (O_1745,N_24173,N_25073);
nor UO_1746 (O_1746,N_26622,N_27499);
nor UO_1747 (O_1747,N_26300,N_29932);
nor UO_1748 (O_1748,N_27974,N_27177);
or UO_1749 (O_1749,N_28958,N_28424);
xor UO_1750 (O_1750,N_26969,N_25144);
or UO_1751 (O_1751,N_26404,N_26467);
or UO_1752 (O_1752,N_27410,N_24529);
xnor UO_1753 (O_1753,N_26926,N_25458);
nor UO_1754 (O_1754,N_24634,N_24713);
nand UO_1755 (O_1755,N_28897,N_26348);
nand UO_1756 (O_1756,N_28933,N_27275);
and UO_1757 (O_1757,N_24993,N_27593);
nand UO_1758 (O_1758,N_27618,N_25690);
nand UO_1759 (O_1759,N_27176,N_27851);
and UO_1760 (O_1760,N_26087,N_25991);
or UO_1761 (O_1761,N_27137,N_25719);
xor UO_1762 (O_1762,N_28161,N_28814);
nand UO_1763 (O_1763,N_27233,N_29711);
or UO_1764 (O_1764,N_26954,N_27810);
nor UO_1765 (O_1765,N_24489,N_27729);
or UO_1766 (O_1766,N_26425,N_24067);
and UO_1767 (O_1767,N_24546,N_28834);
xor UO_1768 (O_1768,N_26440,N_29013);
or UO_1769 (O_1769,N_29417,N_29508);
and UO_1770 (O_1770,N_26980,N_26106);
nand UO_1771 (O_1771,N_24188,N_29765);
nor UO_1772 (O_1772,N_29679,N_25328);
xor UO_1773 (O_1773,N_26563,N_29502);
nand UO_1774 (O_1774,N_24174,N_27800);
and UO_1775 (O_1775,N_25855,N_25262);
or UO_1776 (O_1776,N_25103,N_25453);
or UO_1777 (O_1777,N_28781,N_27937);
xnor UO_1778 (O_1778,N_29823,N_27325);
nand UO_1779 (O_1779,N_26593,N_24169);
and UO_1780 (O_1780,N_28772,N_26357);
nor UO_1781 (O_1781,N_24287,N_28478);
or UO_1782 (O_1782,N_24872,N_26055);
and UO_1783 (O_1783,N_29082,N_25230);
and UO_1784 (O_1784,N_28210,N_26809);
nor UO_1785 (O_1785,N_27797,N_26840);
xnor UO_1786 (O_1786,N_26426,N_25947);
xor UO_1787 (O_1787,N_27608,N_24782);
and UO_1788 (O_1788,N_29480,N_28389);
nand UO_1789 (O_1789,N_25112,N_28840);
xnor UO_1790 (O_1790,N_27147,N_29864);
or UO_1791 (O_1791,N_28123,N_24907);
xor UO_1792 (O_1792,N_27554,N_24945);
xnor UO_1793 (O_1793,N_26918,N_28168);
nand UO_1794 (O_1794,N_27093,N_24156);
xor UO_1795 (O_1795,N_24894,N_25587);
nor UO_1796 (O_1796,N_25271,N_24870);
nor UO_1797 (O_1797,N_29083,N_29376);
nor UO_1798 (O_1798,N_27403,N_26736);
nor UO_1799 (O_1799,N_24111,N_26744);
nand UO_1800 (O_1800,N_28140,N_25849);
xor UO_1801 (O_1801,N_28156,N_25498);
nor UO_1802 (O_1802,N_24455,N_24575);
nor UO_1803 (O_1803,N_28807,N_29292);
or UO_1804 (O_1804,N_28334,N_24633);
or UO_1805 (O_1805,N_28628,N_25881);
nand UO_1806 (O_1806,N_26640,N_27251);
nor UO_1807 (O_1807,N_25869,N_26013);
or UO_1808 (O_1808,N_28295,N_24044);
xnor UO_1809 (O_1809,N_28208,N_26330);
or UO_1810 (O_1810,N_26399,N_27903);
nor UO_1811 (O_1811,N_29723,N_28093);
xor UO_1812 (O_1812,N_27746,N_28453);
nand UO_1813 (O_1813,N_29768,N_28566);
nand UO_1814 (O_1814,N_25727,N_26889);
xnor UO_1815 (O_1815,N_24162,N_28212);
and UO_1816 (O_1816,N_25252,N_27104);
nor UO_1817 (O_1817,N_28835,N_26539);
nor UO_1818 (O_1818,N_27708,N_26037);
xor UO_1819 (O_1819,N_28862,N_27541);
xnor UO_1820 (O_1820,N_28441,N_26921);
and UO_1821 (O_1821,N_29622,N_25597);
or UO_1822 (O_1822,N_29632,N_26666);
or UO_1823 (O_1823,N_27140,N_28039);
or UO_1824 (O_1824,N_24888,N_28061);
nor UO_1825 (O_1825,N_29341,N_27235);
nand UO_1826 (O_1826,N_25346,N_26604);
nand UO_1827 (O_1827,N_28477,N_27353);
xor UO_1828 (O_1828,N_25184,N_29701);
nor UO_1829 (O_1829,N_29874,N_24119);
nand UO_1830 (O_1830,N_26615,N_27924);
xor UO_1831 (O_1831,N_24304,N_25528);
and UO_1832 (O_1832,N_25092,N_29729);
and UO_1833 (O_1833,N_29908,N_25863);
xor UO_1834 (O_1834,N_25076,N_26280);
xnor UO_1835 (O_1835,N_24915,N_26618);
xnor UO_1836 (O_1836,N_29709,N_25021);
nand UO_1837 (O_1837,N_29939,N_28981);
nor UO_1838 (O_1838,N_27790,N_27968);
nor UO_1839 (O_1839,N_26386,N_29049);
nand UO_1840 (O_1840,N_24667,N_27020);
or UO_1841 (O_1841,N_26022,N_29051);
xnor UO_1842 (O_1842,N_28497,N_24417);
and UO_1843 (O_1843,N_24825,N_29944);
xnor UO_1844 (O_1844,N_26309,N_26062);
nor UO_1845 (O_1845,N_28608,N_26485);
xnor UO_1846 (O_1846,N_24848,N_24800);
or UO_1847 (O_1847,N_27042,N_29878);
and UO_1848 (O_1848,N_25094,N_29583);
or UO_1849 (O_1849,N_28575,N_27090);
nor UO_1850 (O_1850,N_25067,N_29338);
nand UO_1851 (O_1851,N_27730,N_24159);
or UO_1852 (O_1852,N_28676,N_26521);
xnor UO_1853 (O_1853,N_28606,N_26335);
and UO_1854 (O_1854,N_25568,N_28551);
and UO_1855 (O_1855,N_24025,N_25033);
nand UO_1856 (O_1856,N_29242,N_24260);
and UO_1857 (O_1857,N_25531,N_27565);
xor UO_1858 (O_1858,N_28697,N_29902);
and UO_1859 (O_1859,N_25725,N_24660);
nor UO_1860 (O_1860,N_28051,N_24365);
or UO_1861 (O_1861,N_27977,N_28364);
or UO_1862 (O_1862,N_26494,N_28861);
xor UO_1863 (O_1863,N_28108,N_29176);
or UO_1864 (O_1864,N_29244,N_27865);
nor UO_1865 (O_1865,N_28530,N_25405);
nor UO_1866 (O_1866,N_25779,N_28557);
or UO_1867 (O_1867,N_24462,N_28914);
and UO_1868 (O_1868,N_26863,N_27559);
nand UO_1869 (O_1869,N_25649,N_24541);
nor UO_1870 (O_1870,N_25516,N_27719);
nand UO_1871 (O_1871,N_28592,N_26572);
nand UO_1872 (O_1872,N_27388,N_27187);
and UO_1873 (O_1873,N_28037,N_26274);
nor UO_1874 (O_1874,N_28618,N_28851);
xor UO_1875 (O_1875,N_24948,N_29187);
nor UO_1876 (O_1876,N_25193,N_28068);
and UO_1877 (O_1877,N_24128,N_25380);
and UO_1878 (O_1878,N_26704,N_28387);
and UO_1879 (O_1879,N_28570,N_29073);
nor UO_1880 (O_1880,N_26031,N_28511);
and UO_1881 (O_1881,N_29738,N_25879);
or UO_1882 (O_1882,N_29365,N_24358);
nor UO_1883 (O_1883,N_25751,N_26093);
xor UO_1884 (O_1884,N_27219,N_24712);
and UO_1885 (O_1885,N_27026,N_24962);
and UO_1886 (O_1886,N_24041,N_26710);
xor UO_1887 (O_1887,N_26480,N_28603);
xnor UO_1888 (O_1888,N_25846,N_26986);
xnor UO_1889 (O_1889,N_24534,N_24593);
or UO_1890 (O_1890,N_25484,N_25004);
nand UO_1891 (O_1891,N_26225,N_28505);
nand UO_1892 (O_1892,N_29954,N_25694);
and UO_1893 (O_1893,N_29275,N_25981);
xnor UO_1894 (O_1894,N_27397,N_29228);
xnor UO_1895 (O_1895,N_27064,N_29517);
or UO_1896 (O_1896,N_29110,N_27246);
nand UO_1897 (O_1897,N_24337,N_29260);
and UO_1898 (O_1898,N_27184,N_24954);
xnor UO_1899 (O_1899,N_27198,N_25801);
xnor UO_1900 (O_1900,N_28873,N_26153);
or UO_1901 (O_1901,N_25823,N_24164);
or UO_1902 (O_1902,N_28107,N_27972);
nand UO_1903 (O_1903,N_29792,N_27214);
xor UO_1904 (O_1904,N_29808,N_24810);
nor UO_1905 (O_1905,N_27734,N_26935);
and UO_1906 (O_1906,N_27431,N_26899);
or UO_1907 (O_1907,N_26886,N_29047);
nand UO_1908 (O_1908,N_25314,N_25295);
xor UO_1909 (O_1909,N_27146,N_28911);
nor UO_1910 (O_1910,N_29157,N_24023);
or UO_1911 (O_1911,N_24504,N_29438);
and UO_1912 (O_1912,N_25546,N_28468);
xnor UO_1913 (O_1913,N_25315,N_27480);
or UO_1914 (O_1914,N_27933,N_27906);
nand UO_1915 (O_1915,N_24307,N_28990);
and UO_1916 (O_1916,N_26060,N_24941);
xor UO_1917 (O_1917,N_25702,N_26771);
xor UO_1918 (O_1918,N_29150,N_28510);
and UO_1919 (O_1919,N_25333,N_25687);
or UO_1920 (O_1920,N_27607,N_28816);
nand UO_1921 (O_1921,N_29910,N_26223);
nand UO_1922 (O_1922,N_26534,N_27599);
nor UO_1923 (O_1923,N_27310,N_27529);
xor UO_1924 (O_1924,N_29780,N_24861);
and UO_1925 (O_1925,N_24088,N_24707);
nor UO_1926 (O_1926,N_28442,N_24117);
and UO_1927 (O_1927,N_29102,N_27434);
xor UO_1928 (O_1928,N_25888,N_25718);
nand UO_1929 (O_1929,N_28773,N_25889);
nand UO_1930 (O_1930,N_25765,N_28415);
nand UO_1931 (O_1931,N_24656,N_28013);
nand UO_1932 (O_1932,N_27402,N_29638);
nand UO_1933 (O_1933,N_29989,N_29773);
and UO_1934 (O_1934,N_27609,N_25898);
xnor UO_1935 (O_1935,N_28535,N_28785);
or UO_1936 (O_1936,N_28242,N_29903);
xor UO_1937 (O_1937,N_28556,N_27057);
nand UO_1938 (O_1938,N_26613,N_28593);
nand UO_1939 (O_1939,N_24970,N_24344);
nor UO_1940 (O_1940,N_29610,N_25447);
and UO_1941 (O_1941,N_25667,N_27173);
and UO_1942 (O_1942,N_25022,N_27846);
nand UO_1943 (O_1943,N_26745,N_24592);
and UO_1944 (O_1944,N_25799,N_28638);
xor UO_1945 (O_1945,N_24873,N_24165);
or UO_1946 (O_1946,N_24306,N_28279);
or UO_1947 (O_1947,N_26934,N_29712);
nand UO_1948 (O_1948,N_24960,N_24340);
xor UO_1949 (O_1949,N_24554,N_29385);
nor UO_1950 (O_1950,N_24226,N_28332);
nor UO_1951 (O_1951,N_26208,N_26289);
xor UO_1952 (O_1952,N_25539,N_25793);
xor UO_1953 (O_1953,N_24740,N_24015);
or UO_1954 (O_1954,N_25051,N_29409);
xor UO_1955 (O_1955,N_28964,N_24830);
or UO_1956 (O_1956,N_25838,N_24738);
nor UO_1957 (O_1957,N_28796,N_27133);
xor UO_1958 (O_1958,N_27544,N_25220);
nand UO_1959 (O_1959,N_26114,N_25634);
and UO_1960 (O_1960,N_27590,N_28800);
or UO_1961 (O_1961,N_27497,N_24473);
nand UO_1962 (O_1962,N_26382,N_25420);
xor UO_1963 (O_1963,N_26825,N_29054);
and UO_1964 (O_1964,N_25034,N_25255);
and UO_1965 (O_1965,N_26268,N_26321);
or UO_1966 (O_1966,N_28689,N_25924);
nand UO_1967 (O_1967,N_27191,N_29994);
or UO_1968 (O_1968,N_25754,N_27789);
xor UO_1969 (O_1969,N_24896,N_24761);
and UO_1970 (O_1970,N_29144,N_27365);
and UO_1971 (O_1971,N_28407,N_24349);
xor UO_1972 (O_1972,N_27378,N_24300);
or UO_1973 (O_1973,N_28157,N_24057);
xnor UO_1974 (O_1974,N_24685,N_25175);
or UO_1975 (O_1975,N_26639,N_24354);
xor UO_1976 (O_1976,N_29522,N_29340);
or UO_1977 (O_1977,N_28868,N_24147);
xor UO_1978 (O_1978,N_29895,N_26709);
nor UO_1979 (O_1979,N_26182,N_26092);
nand UO_1980 (O_1980,N_27552,N_29302);
nand UO_1981 (O_1981,N_27744,N_24675);
nand UO_1982 (O_1982,N_29832,N_27990);
nor UO_1983 (O_1983,N_24177,N_25708);
xnor UO_1984 (O_1984,N_26742,N_24645);
and UO_1985 (O_1985,N_25621,N_28253);
or UO_1986 (O_1986,N_28126,N_27132);
xnor UO_1987 (O_1987,N_25942,N_26454);
or UO_1988 (O_1988,N_25283,N_25953);
nor UO_1989 (O_1989,N_28915,N_29301);
or UO_1990 (O_1990,N_28719,N_25653);
nor UO_1991 (O_1991,N_27652,N_28881);
nand UO_1992 (O_1992,N_24891,N_24982);
nor UO_1993 (O_1993,N_27774,N_25640);
or UO_1994 (O_1994,N_24628,N_26656);
or UO_1995 (O_1995,N_26329,N_25214);
or UO_1996 (O_1996,N_26413,N_26112);
or UO_1997 (O_1997,N_24138,N_25435);
and UO_1998 (O_1998,N_24245,N_25745);
and UO_1999 (O_1999,N_24851,N_24971);
and UO_2000 (O_2000,N_28758,N_24748);
and UO_2001 (O_2001,N_29179,N_27572);
xnor UO_2002 (O_2002,N_29086,N_26469);
nor UO_2003 (O_2003,N_28246,N_28254);
nand UO_2004 (O_2004,N_26339,N_26575);
xor UO_2005 (O_2005,N_27731,N_26161);
xor UO_2006 (O_2006,N_26464,N_26960);
and UO_2007 (O_2007,N_29661,N_25983);
and UO_2008 (O_2008,N_28372,N_24486);
and UO_2009 (O_2009,N_28085,N_28906);
nand UO_2010 (O_2010,N_28391,N_24690);
and UO_2011 (O_2011,N_26381,N_26081);
nand UO_2012 (O_2012,N_29722,N_26788);
nand UO_2013 (O_2013,N_27604,N_29848);
xor UO_2014 (O_2014,N_29399,N_25110);
or UO_2015 (O_2015,N_28236,N_29449);
or UO_2016 (O_2016,N_26789,N_25664);
or UO_2017 (O_2017,N_28909,N_28184);
nand UO_2018 (O_2018,N_25840,N_26668);
or UO_2019 (O_2019,N_27992,N_29814);
nand UO_2020 (O_2020,N_29543,N_25618);
or UO_2021 (O_2021,N_29901,N_29625);
and UO_2022 (O_2022,N_28756,N_24517);
nor UO_2023 (O_2023,N_29477,N_24370);
nand UO_2024 (O_2024,N_24787,N_24140);
xnor UO_2025 (O_2025,N_25249,N_27633);
nand UO_2026 (O_2026,N_26002,N_29794);
xnor UO_2027 (O_2027,N_29845,N_24986);
nor UO_2028 (O_2028,N_28322,N_26503);
nor UO_2029 (O_2029,N_24553,N_28808);
nand UO_2030 (O_2030,N_28062,N_26739);
xnor UO_2031 (O_2031,N_28306,N_26927);
xnor UO_2032 (O_2032,N_29112,N_27518);
or UO_2033 (O_2033,N_24654,N_29184);
xnor UO_2034 (O_2034,N_26513,N_27454);
xnor UO_2035 (O_2035,N_29771,N_25031);
or UO_2036 (O_2036,N_29459,N_26672);
or UO_2037 (O_2037,N_25087,N_27289);
xnor UO_2038 (O_2038,N_28585,N_28249);
and UO_2039 (O_2039,N_24421,N_26564);
and UO_2040 (O_2040,N_28159,N_29950);
or UO_2041 (O_2041,N_28871,N_27661);
and UO_2042 (O_2042,N_28170,N_24739);
or UO_2043 (O_2043,N_25147,N_29063);
nand UO_2044 (O_2044,N_26988,N_27570);
and UO_2045 (O_2045,N_27660,N_24276);
nand UO_2046 (O_2046,N_28017,N_27914);
or UO_2047 (O_2047,N_28775,N_29662);
and UO_2048 (O_2048,N_25063,N_29774);
nor UO_2049 (O_2049,N_27639,N_25199);
nand UO_2050 (O_2050,N_28960,N_24547);
nand UO_2051 (O_2051,N_25318,N_24932);
or UO_2052 (O_2052,N_29818,N_28354);
nand UO_2053 (O_2053,N_25936,N_28187);
xnor UO_2054 (O_2054,N_26782,N_25829);
and UO_2055 (O_2055,N_27980,N_27878);
or UO_2056 (O_2056,N_28991,N_26738);
nor UO_2057 (O_2057,N_27182,N_24568);
nand UO_2058 (O_2058,N_24341,N_26324);
nand UO_2059 (O_2059,N_24010,N_26579);
or UO_2060 (O_2060,N_28268,N_24051);
and UO_2061 (O_2061,N_28471,N_27083);
or UO_2062 (O_2062,N_29104,N_28983);
nor UO_2063 (O_2063,N_24155,N_26756);
nor UO_2064 (O_2064,N_26769,N_28516);
nor UO_2065 (O_2065,N_26852,N_27031);
nor UO_2066 (O_2066,N_28586,N_26198);
nor UO_2067 (O_2067,N_26294,N_26628);
and UO_2068 (O_2068,N_29595,N_28653);
nand UO_2069 (O_2069,N_26507,N_24261);
or UO_2070 (O_2070,N_24350,N_29213);
nor UO_2071 (O_2071,N_28577,N_29169);
and UO_2072 (O_2072,N_28893,N_24702);
and UO_2073 (O_2073,N_27318,N_28302);
or UO_2074 (O_2074,N_24545,N_28936);
nor UO_2075 (O_2075,N_28102,N_27183);
xor UO_2076 (O_2076,N_27589,N_26151);
and UO_2077 (O_2077,N_24185,N_26754);
nor UO_2078 (O_2078,N_28992,N_24033);
and UO_2079 (O_2079,N_24312,N_24452);
and UO_2080 (O_2080,N_24046,N_24924);
and UO_2081 (O_2081,N_28059,N_28630);
or UO_2082 (O_2082,N_29107,N_27874);
nor UO_2083 (O_2083,N_28900,N_28048);
or UO_2084 (O_2084,N_24613,N_25064);
xor UO_2085 (O_2085,N_26030,N_27975);
xor UO_2086 (O_2086,N_25107,N_26121);
and UO_2087 (O_2087,N_24887,N_24561);
nand UO_2088 (O_2088,N_24454,N_26325);
nand UO_2089 (O_2089,N_28966,N_27672);
xor UO_2090 (O_2090,N_25197,N_28828);
nand UO_2091 (O_2091,N_25475,N_27512);
or UO_2092 (O_2092,N_27195,N_25417);
and UO_2093 (O_2093,N_24779,N_29646);
nand UO_2094 (O_2094,N_25350,N_28665);
or UO_2095 (O_2095,N_28336,N_25227);
or UO_2096 (O_2096,N_27257,N_26601);
nor UO_2097 (O_2097,N_25547,N_28536);
or UO_2098 (O_2098,N_26034,N_28289);
xnor UO_2099 (O_2099,N_24013,N_25208);
nor UO_2100 (O_2100,N_29636,N_24978);
nand UO_2101 (O_2101,N_27535,N_28014);
or UO_2102 (O_2102,N_25780,N_25448);
nand UO_2103 (O_2103,N_24961,N_24466);
or UO_2104 (O_2104,N_26517,N_24229);
xor UO_2105 (O_2105,N_24818,N_24788);
and UO_2106 (O_2106,N_28805,N_29885);
and UO_2107 (O_2107,N_26259,N_26495);
nor UO_2108 (O_2108,N_29290,N_29654);
and UO_2109 (O_2109,N_27087,N_28792);
and UO_2110 (O_2110,N_29876,N_25035);
or UO_2111 (O_2111,N_28205,N_27432);
nor UO_2112 (O_2112,N_26205,N_25969);
nor UO_2113 (O_2113,N_25937,N_25264);
or UO_2114 (O_2114,N_26979,N_28646);
or UO_2115 (O_2115,N_26372,N_27506);
nand UO_2116 (O_2116,N_27686,N_29471);
nor UO_2117 (O_2117,N_26051,N_28727);
or UO_2118 (O_2118,N_26609,N_26629);
nand UO_2119 (O_2119,N_25912,N_29612);
nor UO_2120 (O_2120,N_29219,N_28333);
nand UO_2121 (O_2121,N_24718,N_24786);
and UO_2122 (O_2122,N_26790,N_25179);
nand UO_2123 (O_2123,N_29094,N_26328);
nand UO_2124 (O_2124,N_27563,N_25746);
and UO_2125 (O_2125,N_29737,N_28031);
and UO_2126 (O_2126,N_26277,N_29693);
and UO_2127 (O_2127,N_27027,N_29826);
xnor UO_2128 (O_2128,N_28994,N_28523);
and UO_2129 (O_2129,N_25646,N_27955);
or UO_2130 (O_2130,N_24601,N_24112);
or UO_2131 (O_2131,N_29088,N_27270);
and UO_2132 (O_2132,N_24321,N_25065);
nand UO_2133 (O_2133,N_25588,N_28549);
or UO_2134 (O_2134,N_27373,N_27524);
xor UO_2135 (O_2135,N_27889,N_26770);
nand UO_2136 (O_2136,N_27690,N_27311);
xnor UO_2137 (O_2137,N_29787,N_27709);
nand UO_2138 (O_2138,N_29360,N_25010);
xor UO_2139 (O_2139,N_24474,N_27827);
or UO_2140 (O_2140,N_28884,N_27726);
nand UO_2141 (O_2141,N_24477,N_28885);
xor UO_2142 (O_2142,N_25436,N_26124);
nand UO_2143 (O_2143,N_24186,N_28262);
and UO_2144 (O_2144,N_25000,N_24743);
xnor UO_2145 (O_2145,N_29080,N_29559);
and UO_2146 (O_2146,N_26757,N_24381);
xor UO_2147 (O_2147,N_27329,N_25449);
or UO_2148 (O_2148,N_28072,N_24987);
or UO_2149 (O_2149,N_24315,N_27591);
and UO_2150 (O_2150,N_25997,N_29643);
nor UO_2151 (O_2151,N_28223,N_28829);
and UO_2152 (O_2152,N_27131,N_27682);
xor UO_2153 (O_2153,N_27685,N_25088);
or UO_2154 (O_2154,N_26110,N_25211);
and UO_2155 (O_2155,N_27084,N_28970);
nor UO_2156 (O_2156,N_29574,N_24274);
nand UO_2157 (O_2157,N_25585,N_24453);
xor UO_2158 (O_2158,N_29451,N_26681);
xnor UO_2159 (O_2159,N_27625,N_28428);
or UO_2160 (O_2160,N_27495,N_29036);
xor UO_2161 (O_2161,N_25265,N_29745);
nand UO_2162 (O_2162,N_27197,N_24881);
xnor UO_2163 (O_2163,N_27670,N_25485);
nand UO_2164 (O_2164,N_26345,N_25628);
nor UO_2165 (O_2165,N_29650,N_29037);
or UO_2166 (O_2166,N_26202,N_28298);
or UO_2167 (O_2167,N_24737,N_28328);
nand UO_2168 (O_2168,N_25377,N_27794);
xor UO_2169 (O_2169,N_29590,N_25456);
nor UO_2170 (O_2170,N_25744,N_26038);
or UO_2171 (O_2171,N_29879,N_28195);
and UO_2172 (O_2172,N_26871,N_25857);
xnor UO_2173 (O_2173,N_25789,N_24910);
or UO_2174 (O_2174,N_26146,N_29754);
nor UO_2175 (O_2175,N_26005,N_24959);
nand UO_2176 (O_2176,N_25125,N_29166);
nand UO_2177 (O_2177,N_29074,N_24823);
nand UO_2178 (O_2178,N_24035,N_27745);
and UO_2179 (O_2179,N_24062,N_26138);
and UO_2180 (O_2180,N_28263,N_25286);
xor UO_2181 (O_2181,N_26664,N_26349);
nor UO_2182 (O_2182,N_29974,N_26936);
xor UO_2183 (O_2183,N_27540,N_24614);
and UO_2184 (O_2184,N_28466,N_25705);
or UO_2185 (O_2185,N_28366,N_29927);
xor UO_2186 (O_2186,N_29487,N_29582);
nand UO_2187 (O_2187,N_26814,N_25403);
xnor UO_2188 (O_2188,N_24832,N_26471);
or UO_2189 (O_2189,N_24493,N_28010);
xnor UO_2190 (O_2190,N_28180,N_26883);
nand UO_2191 (O_2191,N_27303,N_27114);
or UO_2192 (O_2192,N_29380,N_28721);
nand UO_2193 (O_2193,N_29192,N_24751);
xnor UO_2194 (O_2194,N_29866,N_25904);
and UO_2195 (O_2195,N_28151,N_28985);
nand UO_2196 (O_2196,N_26712,N_26838);
nand UO_2197 (O_2197,N_24801,N_25615);
xnor UO_2198 (O_2198,N_28929,N_28852);
nand UO_2199 (O_2199,N_27645,N_25196);
nand UO_2200 (O_2200,N_24802,N_25518);
or UO_2201 (O_2201,N_25731,N_25882);
nand UO_2202 (O_2202,N_28555,N_28811);
or UO_2203 (O_2203,N_24981,N_27082);
or UO_2204 (O_2204,N_27461,N_28940);
or UO_2205 (O_2205,N_29871,N_25886);
xor UO_2206 (O_2206,N_29126,N_24995);
nor UO_2207 (O_2207,N_25060,N_26211);
nor UO_2208 (O_2208,N_26605,N_26671);
xnor UO_2209 (O_2209,N_28329,N_26888);
nand UO_2210 (O_2210,N_28020,N_28057);
xor UO_2211 (O_2211,N_25773,N_25412);
xor UO_2212 (O_2212,N_27129,N_24372);
and UO_2213 (O_2213,N_24082,N_29423);
nor UO_2214 (O_2214,N_29525,N_29934);
nor UO_2215 (O_2215,N_29087,N_24115);
and UO_2216 (O_2216,N_29782,N_26841);
xor UO_2217 (O_2217,N_27481,N_24045);
or UO_2218 (O_2218,N_29708,N_26560);
xor UO_2219 (O_2219,N_29343,N_25508);
nand UO_2220 (O_2220,N_29858,N_25002);
nor UO_2221 (O_2221,N_24445,N_29598);
and UO_2222 (O_2222,N_27702,N_27215);
or UO_2223 (O_2223,N_27816,N_24479);
xnor UO_2224 (O_2224,N_24730,N_27760);
xor UO_2225 (O_2225,N_29713,N_28396);
and UO_2226 (O_2226,N_26643,N_25029);
and UO_2227 (O_2227,N_25806,N_25636);
nand UO_2228 (O_2228,N_25409,N_27667);
xor UO_2229 (O_2229,N_26735,N_26964);
nor UO_2230 (O_2230,N_28972,N_29076);
nor UO_2231 (O_2231,N_25929,N_28374);
and UO_2232 (O_2232,N_26004,N_28722);
and UO_2233 (O_2233,N_27039,N_24598);
and UO_2234 (O_2234,N_27150,N_29664);
or UO_2235 (O_2235,N_25079,N_27689);
or UO_2236 (O_2236,N_27892,N_25958);
xor UO_2237 (O_2237,N_27728,N_29811);
xnor UO_2238 (O_2238,N_29182,N_29407);
and UO_2239 (O_2239,N_26864,N_25920);
or UO_2240 (O_2240,N_24901,N_24002);
nand UO_2241 (O_2241,N_26677,N_24208);
xnor UO_2242 (O_2242,N_25673,N_29766);
nor UO_2243 (O_2243,N_28957,N_27061);
nor UO_2244 (O_2244,N_25152,N_26968);
or UO_2245 (O_2245,N_26943,N_28493);
or UO_2246 (O_2246,N_28457,N_24923);
and UO_2247 (O_2247,N_25632,N_27910);
or UO_2248 (O_2248,N_26295,N_29264);
nor UO_2249 (O_2249,N_29155,N_28404);
or UO_2250 (O_2250,N_26052,N_28243);
xor UO_2251 (O_2251,N_27261,N_29364);
nand UO_2252 (O_2252,N_27249,N_25238);
and UO_2253 (O_2253,N_28748,N_25808);
xor UO_2254 (O_2254,N_25303,N_29964);
nand UO_2255 (O_2255,N_26024,N_24339);
or UO_2256 (O_2256,N_25003,N_26460);
and UO_2257 (O_2257,N_27456,N_24220);
xnor UO_2258 (O_2258,N_25273,N_27662);
nand UO_2259 (O_2259,N_29607,N_26057);
nor UO_2260 (O_2260,N_24095,N_28220);
nor UO_2261 (O_2261,N_29148,N_26995);
and UO_2262 (O_2262,N_27327,N_24677);
nor UO_2263 (O_2263,N_28087,N_29162);
xor UO_2264 (O_2264,N_28413,N_26482);
nand UO_2265 (O_2265,N_29118,N_27812);
nor UO_2266 (O_2266,N_29404,N_25097);
nor UO_2267 (O_2267,N_25733,N_27655);
nor UO_2268 (O_2268,N_26219,N_27942);
nand UO_2269 (O_2269,N_26468,N_24333);
or UO_2270 (O_2270,N_28024,N_24658);
and UO_2271 (O_2271,N_29779,N_29714);
nand UO_2272 (O_2272,N_24542,N_27963);
or UO_2273 (O_2273,N_28278,N_27306);
nor UO_2274 (O_2274,N_28609,N_24280);
nor UO_2275 (O_2275,N_29046,N_27775);
and UO_2276 (O_2276,N_25400,N_26180);
nand UO_2277 (O_2277,N_24767,N_28003);
or UO_2278 (O_2278,N_24619,N_25612);
or UO_2279 (O_2279,N_24644,N_29799);
xor UO_2280 (O_2280,N_26630,N_25954);
nor UO_2281 (O_2281,N_25015,N_27424);
nor UO_2282 (O_2282,N_28046,N_24342);
nor UO_2283 (O_2283,N_24316,N_25530);
or UO_2284 (O_2284,N_29604,N_25292);
and UO_2285 (O_2285,N_28710,N_29585);
nand UO_2286 (O_2286,N_26119,N_29812);
nor UO_2287 (O_2287,N_25946,N_27459);
and UO_2288 (O_2288,N_24992,N_27779);
nand UO_2289 (O_2289,N_26010,N_26167);
and UO_2290 (O_2290,N_27298,N_29446);
xor UO_2291 (O_2291,N_25234,N_29623);
nor UO_2292 (O_2292,N_27673,N_24662);
or UO_2293 (O_2293,N_29151,N_26209);
xnor UO_2294 (O_2294,N_25037,N_26337);
nand UO_2295 (O_2295,N_27736,N_27152);
or UO_2296 (O_2296,N_27533,N_28080);
and UO_2297 (O_2297,N_26220,N_28090);
nor UO_2298 (O_2298,N_29296,N_24203);
nand UO_2299 (O_2299,N_28729,N_25843);
xnor UO_2300 (O_2300,N_24854,N_26913);
xnor UO_2301 (O_2301,N_27956,N_29130);
nor UO_2302 (O_2302,N_27167,N_27473);
and UO_2303 (O_2303,N_29506,N_29785);
nor UO_2304 (O_2304,N_29204,N_26200);
nor UO_2305 (O_2305,N_29580,N_27296);
nand UO_2306 (O_2306,N_28365,N_28833);
nor UO_2307 (O_2307,N_26524,N_28348);
nand UO_2308 (O_2308,N_26008,N_24122);
nand UO_2309 (O_2309,N_29571,N_25365);
and UO_2310 (O_2310,N_29368,N_26978);
or UO_2311 (O_2311,N_26279,N_29123);
xor UO_2312 (O_2312,N_25887,N_25465);
or UO_2313 (O_2313,N_26312,N_29391);
xor UO_2314 (O_2314,N_28857,N_29218);
nor UO_2315 (O_2315,N_25496,N_28864);
xor UO_2316 (O_2316,N_28844,N_25876);
and UO_2317 (O_2317,N_29295,N_28318);
xnor UO_2318 (O_2318,N_27366,N_29682);
and UO_2319 (O_2319,N_27537,N_28490);
or UO_2320 (O_2320,N_29886,N_24113);
or UO_2321 (O_2321,N_28070,N_27354);
nand UO_2322 (O_2322,N_27801,N_28912);
and UO_2323 (O_2323,N_25976,N_29869);
nor UO_2324 (O_2324,N_29647,N_25800);
xor UO_2325 (O_2325,N_29948,N_27580);
and UO_2326 (O_2326,N_27893,N_29324);
or UO_2327 (O_2327,N_25085,N_24408);
and UO_2328 (O_2328,N_25899,N_26306);
xor UO_2329 (O_2329,N_28091,N_26058);
or UO_2330 (O_2330,N_25059,N_26602);
xor UO_2331 (O_2331,N_28084,N_27326);
xor UO_2332 (O_2332,N_26801,N_28791);
nand UO_2333 (O_2333,N_29626,N_29498);
and UO_2334 (O_2334,N_29039,N_27896);
nand UO_2335 (O_2335,N_29217,N_28294);
or UO_2336 (O_2336,N_26088,N_29326);
xor UO_2337 (O_2337,N_29225,N_27743);
nand UO_2338 (O_2338,N_27965,N_29569);
xnor UO_2339 (O_2339,N_25511,N_28504);
nand UO_2340 (O_2340,N_26824,N_29579);
nand UO_2341 (O_2341,N_26837,N_25071);
or UO_2342 (O_2342,N_29584,N_24426);
xnor UO_2343 (O_2343,N_27940,N_28996);
nand UO_2344 (O_2344,N_28942,N_26510);
or UO_2345 (O_2345,N_27791,N_29307);
nand UO_2346 (O_2346,N_29488,N_27300);
nand UO_2347 (O_2347,N_29416,N_24376);
nor UO_2348 (O_2348,N_27982,N_25145);
and UO_2349 (O_2349,N_28978,N_24616);
xor UO_2350 (O_2350,N_28759,N_25684);
nand UO_2351 (O_2351,N_26264,N_28602);
or UO_2352 (O_2352,N_27418,N_29684);
and UO_2353 (O_2353,N_25713,N_27469);
and UO_2354 (O_2354,N_27923,N_29641);
nor UO_2355 (O_2355,N_28971,N_26012);
nor UO_2356 (O_2356,N_29250,N_26447);
or UO_2357 (O_2357,N_28822,N_27074);
and UO_2358 (O_2358,N_25091,N_26102);
and UO_2359 (O_2359,N_26015,N_28797);
and UO_2360 (O_2360,N_26818,N_24900);
and UO_2361 (O_2361,N_24256,N_24150);
xor UO_2362 (O_2362,N_26159,N_25335);
nand UO_2363 (O_2363,N_24219,N_27784);
nand UO_2364 (O_2364,N_24357,N_27987);
or UO_2365 (O_2365,N_24766,N_29651);
nor UO_2366 (O_2366,N_28779,N_29052);
nor UO_2367 (O_2367,N_27741,N_26353);
and UO_2368 (O_2368,N_25192,N_27098);
xnor UO_2369 (O_2369,N_26695,N_27013);
or UO_2370 (O_2370,N_27981,N_27205);
nand UO_2371 (O_2371,N_26215,N_28380);
or UO_2372 (O_2372,N_29167,N_29116);
or UO_2373 (O_2373,N_29981,N_25559);
nand UO_2374 (O_2374,N_26275,N_28012);
or UO_2375 (O_2375,N_29829,N_29304);
or UO_2376 (O_2376,N_26388,N_25293);
xor UO_2377 (O_2377,N_27045,N_25026);
or UO_2378 (O_2378,N_26210,N_24366);
and UO_2379 (O_2379,N_25427,N_27357);
or UO_2380 (O_2380,N_27925,N_24708);
nor UO_2381 (O_2381,N_24871,N_29269);
nor UO_2382 (O_2382,N_29725,N_28209);
nand UO_2383 (O_2383,N_26740,N_27926);
or UO_2384 (O_2384,N_26674,N_26511);
xor UO_2385 (O_2385,N_24017,N_25482);
nand UO_2386 (O_2386,N_28129,N_26265);
nor UO_2387 (O_2387,N_24736,N_25046);
xor UO_2388 (O_2388,N_24460,N_27231);
and UO_2389 (O_2389,N_25337,N_24563);
and UO_2390 (O_2390,N_26703,N_26164);
or UO_2391 (O_2391,N_29168,N_26907);
nor UO_2392 (O_2392,N_27255,N_25217);
xor UO_2393 (O_2393,N_29216,N_24552);
and UO_2394 (O_2394,N_26687,N_29526);
or UO_2395 (O_2395,N_27653,N_24055);
nand UO_2396 (O_2396,N_26422,N_25494);
and UO_2397 (O_2397,N_27475,N_27579);
or UO_2398 (O_2398,N_24756,N_28582);
xnor UO_2399 (O_2399,N_26098,N_28741);
or UO_2400 (O_2400,N_27107,N_24973);
and UO_2401 (O_2401,N_29600,N_25480);
xnor UO_2402 (O_2402,N_24597,N_25146);
or UO_2403 (O_2403,N_26305,N_27517);
and UO_2404 (O_2404,N_28288,N_24216);
or UO_2405 (O_2405,N_29038,N_25824);
and UO_2406 (O_2406,N_26367,N_27877);
or UO_2407 (O_2407,N_25108,N_28235);
or UO_2408 (O_2408,N_29892,N_26946);
and UO_2409 (O_2409,N_28543,N_27294);
and UO_2410 (O_2410,N_24686,N_25492);
xor UO_2411 (O_2411,N_24244,N_26298);
nor UO_2412 (O_2412,N_25163,N_27400);
and UO_2413 (O_2413,N_25246,N_25488);
nor UO_2414 (O_2414,N_27692,N_29707);
and UO_2415 (O_2415,N_24405,N_24232);
and UO_2416 (O_2416,N_26242,N_24375);
or UO_2417 (O_2417,N_28968,N_28734);
nor UO_2418 (O_2418,N_29680,N_29514);
or UO_2419 (O_2419,N_25225,N_24195);
and UO_2420 (O_2420,N_27011,N_26567);
nor UO_2421 (O_2421,N_25497,N_28813);
or UO_2422 (O_2422,N_25961,N_25582);
nor UO_2423 (O_2423,N_24550,N_25389);
xor UO_2424 (O_2424,N_24798,N_28925);
and UO_2425 (O_2425,N_29642,N_28211);
nand UO_2426 (O_2426,N_24179,N_26807);
nor UO_2427 (O_2427,N_28661,N_29860);
or UO_2428 (O_2428,N_29925,N_24669);
nor UO_2429 (O_2429,N_28703,N_25590);
nand UO_2430 (O_2430,N_27063,N_26984);
and UO_2431 (O_2431,N_26720,N_27677);
nor UO_2432 (O_2432,N_28357,N_29867);
nor UO_2433 (O_2433,N_28863,N_28666);
nor UO_2434 (O_2434,N_26616,N_24464);
xor UO_2435 (O_2435,N_25525,N_26296);
nand UO_2436 (O_2436,N_28855,N_29282);
nor UO_2437 (O_2437,N_28055,N_25776);
or UO_2438 (O_2438,N_29400,N_27280);
nor UO_2439 (O_2439,N_29489,N_28926);
or UO_2440 (O_2440,N_29694,N_25967);
nor UO_2441 (O_2441,N_24456,N_29817);
nor UO_2442 (O_2442,N_24885,N_25943);
nor UO_2443 (O_2443,N_28215,N_26971);
and UO_2444 (O_2444,N_29099,N_28237);
or UO_2445 (O_2445,N_27869,N_27379);
or UO_2446 (O_2446,N_26915,N_26958);
or UO_2447 (O_2447,N_27241,N_29644);
xor UO_2448 (O_2448,N_25692,N_27668);
xor UO_2449 (O_2449,N_24727,N_28203);
xor UO_2450 (O_2450,N_24052,N_29311);
nor UO_2451 (O_2451,N_26402,N_26366);
xor UO_2452 (O_2452,N_27936,N_26994);
xor UO_2453 (O_2453,N_25267,N_27279);
and UO_2454 (O_2454,N_27838,N_26433);
or UO_2455 (O_2455,N_24549,N_28610);
or UO_2456 (O_2456,N_29491,N_27642);
or UO_2457 (O_2457,N_25357,N_24325);
nand UO_2458 (O_2458,N_27931,N_27386);
or UO_2459 (O_2459,N_25884,N_27445);
or UO_2460 (O_2460,N_24184,N_24735);
or UO_2461 (O_2461,N_24313,N_26267);
nor UO_2462 (O_2462,N_25290,N_26760);
xor UO_2463 (O_2463,N_26351,N_24042);
nor UO_2464 (O_2464,N_24691,N_28764);
and UO_2465 (O_2465,N_27005,N_28397);
xor UO_2466 (O_2466,N_29198,N_29828);
nor UO_2467 (O_2467,N_28327,N_29009);
nor UO_2468 (O_2468,N_26775,N_28921);
nor UO_2469 (O_2469,N_26974,N_25741);
nor UO_2470 (O_2470,N_27449,N_25704);
or UO_2471 (O_2471,N_24390,N_26906);
or UO_2472 (O_2472,N_26635,N_24943);
nand UO_2473 (O_2473,N_26218,N_24502);
nand UO_2474 (O_2474,N_28809,N_29285);
and UO_2475 (O_2475,N_25626,N_29786);
xnor UO_2476 (O_2476,N_28303,N_29558);
nor UO_2477 (O_2477,N_27482,N_25802);
and UO_2478 (O_2478,N_27581,N_25378);
nor UO_2479 (O_2479,N_25517,N_27134);
nand UO_2480 (O_2480,N_26975,N_28447);
or UO_2481 (O_2481,N_28931,N_27455);
nand UO_2482 (O_2482,N_28654,N_27803);
xnor UO_2483 (O_2483,N_26679,N_24936);
nor UO_2484 (O_2484,N_29971,N_25614);
or UO_2485 (O_2485,N_26174,N_29238);
xnor UO_2486 (O_2486,N_25473,N_24785);
xor UO_2487 (O_2487,N_28182,N_27089);
nor UO_2488 (O_2488,N_25331,N_25489);
nor UO_2489 (O_2489,N_28941,N_25706);
nor UO_2490 (O_2490,N_29977,N_28004);
nand UO_2491 (O_2491,N_28319,N_25395);
nor UO_2492 (O_2492,N_29535,N_26255);
nand UO_2493 (O_2493,N_28491,N_24204);
xnor UO_2494 (O_2494,N_24765,N_29386);
xnor UO_2495 (O_2495,N_27979,N_28463);
xor UO_2496 (O_2496,N_24438,N_24911);
xor UO_2497 (O_2497,N_26583,N_29022);
nand UO_2498 (O_2498,N_27983,N_25153);
and UO_2499 (O_2499,N_27501,N_28018);
nor UO_2500 (O_2500,N_28116,N_28456);
and UO_2501 (O_2501,N_29040,N_28461);
nand UO_2502 (O_2502,N_28101,N_26552);
nand UO_2503 (O_2503,N_26487,N_28705);
nor UO_2504 (O_2504,N_26950,N_24511);
nand UO_2505 (O_2505,N_27308,N_25172);
or UO_2506 (O_2506,N_24123,N_29317);
nor UO_2507 (O_2507,N_25897,N_29672);
and UO_2508 (O_2508,N_27848,N_24431);
nand UO_2509 (O_2509,N_24096,N_27665);
nand UO_2510 (O_2510,N_27740,N_25558);
and UO_2511 (O_2511,N_25661,N_24562);
nand UO_2512 (O_2512,N_26158,N_24805);
nor UO_2513 (O_2513,N_24496,N_27886);
or UO_2514 (O_2514,N_26025,N_27361);
nand UO_2515 (O_2515,N_26304,N_28950);
xor UO_2516 (O_2516,N_29545,N_25028);
or UO_2517 (O_2517,N_28934,N_28686);
nor UO_2518 (O_2518,N_24622,N_26965);
nand UO_2519 (O_2519,N_27871,N_29209);
nor UO_2520 (O_2520,N_27457,N_28737);
xnor UO_2521 (O_2521,N_29281,N_27100);
xor UO_2522 (O_2522,N_27355,N_24482);
nand UO_2523 (O_2523,N_25397,N_25501);
xnor UO_2524 (O_2524,N_28363,N_26765);
nand UO_2525 (O_2525,N_24355,N_26147);
nand UO_2526 (O_2526,N_25712,N_27564);
xor UO_2527 (O_2527,N_29505,N_28660);
nand UO_2528 (O_2528,N_28956,N_24676);
or UO_2529 (O_2529,N_24903,N_27911);
nand UO_2530 (O_2530,N_24288,N_29025);
and UO_2531 (O_2531,N_26066,N_27121);
nand UO_2532 (O_2532,N_29055,N_28204);
nand UO_2533 (O_2533,N_29105,N_27392);
nand UO_2534 (O_2534,N_29331,N_25371);
nor UO_2535 (O_2535,N_26276,N_25272);
xor UO_2536 (O_2536,N_27189,N_26450);
and UO_2537 (O_2537,N_24551,N_24432);
xnor UO_2538 (O_2538,N_26715,N_24014);
or UO_2539 (O_2539,N_28147,N_29544);
xor UO_2540 (O_2540,N_25239,N_24950);
nor UO_2541 (O_2541,N_29254,N_25390);
nand UO_2542 (O_2542,N_26430,N_25053);
nor UO_2543 (O_2543,N_25048,N_28916);
and UO_2544 (O_2544,N_27458,N_26036);
or UO_2545 (O_2545,N_26647,N_26611);
xor UO_2546 (O_2546,N_29966,N_27267);
or UO_2547 (O_2547,N_24649,N_26448);
nand UO_2548 (O_2548,N_29084,N_27557);
nor UO_2549 (O_2549,N_27920,N_24803);
and UO_2550 (O_2550,N_25173,N_28384);
and UO_2551 (O_2551,N_24347,N_28695);
nand UO_2552 (O_2552,N_26505,N_28612);
xnor UO_2553 (O_2553,N_24303,N_29258);
or UO_2554 (O_2554,N_25372,N_24448);
or UO_2555 (O_2555,N_25883,N_24391);
nor UO_2556 (O_2556,N_25027,N_27870);
or UO_2557 (O_2557,N_27951,N_27059);
or UO_2558 (O_2558,N_26474,N_29271);
and UO_2559 (O_2559,N_25996,N_26942);
xor UO_2560 (O_2560,N_29366,N_27463);
nand UO_2561 (O_2561,N_25729,N_27750);
nor UO_2562 (O_2562,N_24746,N_25174);
or UO_2563 (O_2563,N_24773,N_28465);
and UO_2564 (O_2564,N_29145,N_25944);
and UO_2565 (O_2565,N_27762,N_25736);
or UO_2566 (O_2566,N_24318,N_28815);
or UO_2567 (O_2567,N_28798,N_27067);
xnor UO_2568 (O_2568,N_29541,N_26320);
nor UO_2569 (O_2569,N_25178,N_29229);
nor UO_2570 (O_2570,N_26794,N_24588);
and UO_2571 (O_2571,N_25463,N_27516);
nor UO_2572 (O_2572,N_26783,N_24975);
xor UO_2573 (O_2573,N_27586,N_26416);
nand UO_2574 (O_2574,N_26362,N_25282);
or UO_2575 (O_2575,N_24762,N_24364);
or UO_2576 (O_2576,N_24435,N_28625);
xnor UO_2577 (O_2577,N_27002,N_28518);
nand UO_2578 (O_2578,N_29742,N_25892);
nor UO_2579 (O_2579,N_28382,N_25933);
nand UO_2580 (O_2580,N_29106,N_29500);
nor UO_2581 (O_2581,N_27460,N_24187);
or UO_2582 (O_2582,N_24965,N_28865);
nor UO_2583 (O_2583,N_27314,N_26441);
nand UO_2584 (O_2584,N_25138,N_25584);
nand UO_2585 (O_2585,N_24745,N_29261);
nand UO_2586 (O_2586,N_26427,N_29630);
and UO_2587 (O_2587,N_24931,N_24419);
nor UO_2588 (O_2588,N_26457,N_24172);
and UO_2589 (O_2589,N_28707,N_27401);
and UO_2590 (O_2590,N_28652,N_28131);
nor UO_2591 (O_2591,N_27119,N_25760);
nor UO_2592 (O_2592,N_28778,N_24606);
or UO_2593 (O_2593,N_24077,N_26541);
xnor UO_2594 (O_2594,N_26981,N_26396);
and UO_2595 (O_2595,N_27428,N_27932);
nand UO_2596 (O_2596,N_24586,N_26860);
xnor UO_2597 (O_2597,N_26491,N_26529);
and UO_2598 (O_2598,N_27680,N_27505);
xnor UO_2599 (O_2599,N_27420,N_29345);
nand UO_2600 (O_2600,N_26676,N_24237);
nand UO_2601 (O_2601,N_28520,N_26419);
nand UO_2602 (O_2602,N_25979,N_26688);
xor UO_2603 (O_2603,N_27613,N_24009);
nand UO_2604 (O_2604,N_28733,N_25534);
nand UO_2605 (O_2605,N_28517,N_25926);
and UO_2606 (O_2606,N_26108,N_25913);
xnor UO_2607 (O_2607,N_28414,N_28216);
nand UO_2608 (O_2608,N_27199,N_24361);
and UO_2609 (O_2609,N_24190,N_28410);
nand UO_2610 (O_2610,N_29367,N_26080);
or UO_2611 (O_2611,N_27526,N_26365);
or UO_2612 (O_2612,N_25623,N_28681);
xnor UO_2613 (O_2613,N_28825,N_29521);
nor UO_2614 (O_2614,N_26271,N_29617);
xnor UO_2615 (O_2615,N_26486,N_25278);
or UO_2616 (O_2616,N_27934,N_28188);
nand UO_2617 (O_2617,N_29710,N_28631);
and UO_2618 (O_2618,N_27527,N_25566);
nor UO_2619 (O_2619,N_28025,N_25353);
and UO_2620 (O_2620,N_24040,N_25964);
nor UO_2621 (O_2621,N_29616,N_25263);
or UO_2622 (O_2622,N_24878,N_29075);
and UO_2623 (O_2623,N_26437,N_27534);
nor UO_2624 (O_2624,N_26701,N_29401);
or UO_2625 (O_2625,N_24236,N_29406);
xnor UO_2626 (O_2626,N_24852,N_25013);
or UO_2627 (O_2627,N_27252,N_24526);
nor UO_2628 (O_2628,N_29114,N_26718);
or UO_2629 (O_2629,N_25012,N_29943);
xor UO_2630 (O_2630,N_29240,N_24624);
xor UO_2631 (O_2631,N_25165,N_26166);
xnor UO_2632 (O_2632,N_29410,N_25688);
or UO_2633 (O_2633,N_26961,N_28767);
nor UO_2634 (O_2634,N_26484,N_28124);
nor UO_2635 (O_2635,N_29458,N_27471);
xnor UO_2636 (O_2636,N_25106,N_29803);
and UO_2637 (O_2637,N_24869,N_24054);
or UO_2638 (O_2638,N_25726,N_29537);
nand UO_2639 (O_2639,N_27404,N_25430);
nand UO_2640 (O_2640,N_24747,N_26130);
nand UO_2641 (O_2641,N_28623,N_28245);
or UO_2642 (O_2642,N_25468,N_24141);
or UO_2643 (O_2643,N_25968,N_25995);
or UO_2644 (O_2644,N_27307,N_29631);
nor UO_2645 (O_2645,N_25363,N_28663);
and UO_2646 (O_2646,N_29724,N_24402);
or UO_2647 (O_2647,N_28388,N_25957);
xnor UO_2648 (O_2648,N_27787,N_25834);
xor UO_2649 (O_2649,N_28284,N_27099);
xnor UO_2650 (O_2650,N_27330,N_26706);
nand UO_2651 (O_2651,N_28356,N_25098);
nor UO_2652 (O_2652,N_26420,N_28548);
nand UO_2653 (O_2653,N_28744,N_29835);
nor UO_2654 (O_2654,N_29493,N_27575);
xnor UO_2655 (O_2655,N_24247,N_24699);
xor UO_2656 (O_2656,N_24537,N_25674);
or UO_2657 (O_2657,N_27010,N_24269);
xor UO_2658 (O_2658,N_27901,N_29735);
and UO_2659 (O_2659,N_28768,N_28531);
nor UO_2660 (O_2660,N_29482,N_28114);
nand UO_2661 (O_2661,N_28907,N_26949);
nor UO_2662 (O_2662,N_24757,N_24958);
nand UO_2663 (O_2663,N_27567,N_27873);
nand UO_2664 (O_2664,N_26808,N_25428);
xor UO_2665 (O_2665,N_27333,N_24841);
nand UO_2666 (O_2666,N_29441,N_26562);
xnor UO_2667 (O_2667,N_25782,N_29231);
or UO_2668 (O_2668,N_25474,N_26470);
or UO_2669 (O_2669,N_29131,N_25637);
or UO_2670 (O_2670,N_27944,N_24824);
xnor UO_2671 (O_2671,N_26322,N_29581);
nor UO_2672 (O_2672,N_29279,N_26456);
xnor UO_2673 (O_2673,N_24469,N_29695);
or UO_2674 (O_2674,N_28315,N_26798);
or UO_2675 (O_2675,N_29951,N_27638);
and UO_2676 (O_2676,N_24362,N_24281);
nand UO_2677 (O_2677,N_24513,N_27227);
xnor UO_2678 (O_2678,N_26175,N_25908);
nor UO_2679 (O_2679,N_27814,N_29330);
nor UO_2680 (O_2680,N_26127,N_26126);
xor UO_2681 (O_2681,N_26831,N_29056);
and UO_2682 (O_2682,N_25784,N_27112);
and UO_2683 (O_2683,N_28271,N_27742);
and UO_2684 (O_2684,N_29164,N_29030);
and UO_2685 (O_2685,N_29868,N_25574);
nand UO_2686 (O_2686,N_24700,N_25490);
nor UO_2687 (O_2687,N_25207,N_27419);
or UO_2688 (O_2688,N_24856,N_29637);
and UO_2689 (O_2689,N_24109,N_28094);
nor UO_2690 (O_2690,N_27381,N_27704);
or UO_2691 (O_2691,N_28560,N_29035);
and UO_2692 (O_2692,N_28193,N_29591);
nor UO_2693 (O_2693,N_25832,N_25743);
nand UO_2694 (O_2694,N_27451,N_29872);
nand UO_2695 (O_2695,N_24231,N_27899);
or UO_2696 (O_2696,N_29237,N_29349);
nor UO_2697 (O_2697,N_29840,N_24914);
xor UO_2698 (O_2698,N_26911,N_29677);
nand UO_2699 (O_2699,N_29978,N_27207);
and UO_2700 (O_2700,N_29660,N_28293);
or UO_2701 (O_2701,N_27514,N_28368);
xor UO_2702 (O_2702,N_27854,N_27717);
and UO_2703 (O_2703,N_27634,N_24512);
or UO_2704 (O_2704,N_24157,N_26009);
xor UO_2705 (O_2705,N_24775,N_27969);
or UO_2706 (O_2706,N_28922,N_28589);
nor UO_2707 (O_2707,N_26947,N_28910);
xor UO_2708 (O_2708,N_25616,N_29810);
nand UO_2709 (O_2709,N_28073,N_26614);
nand UO_2710 (O_2710,N_25695,N_24356);
nand UO_2711 (O_2711,N_24193,N_25523);
nor UO_2712 (O_2712,N_28986,N_27521);
nand UO_2713 (O_2713,N_26711,N_25982);
nand UO_2714 (O_2714,N_28275,N_24277);
nor UO_2715 (O_2715,N_24503,N_24912);
nor UO_2716 (O_2716,N_25119,N_24323);
xor UO_2717 (O_2717,N_29272,N_29153);
xnor UO_2718 (O_2718,N_24898,N_29601);
xnor UO_2719 (O_2719,N_24729,N_27716);
and UO_2720 (O_2720,N_29658,N_27831);
or UO_2721 (O_2721,N_27046,N_26953);
xor UO_2722 (O_2722,N_26407,N_27406);
and UO_2723 (O_2723,N_24778,N_29432);
nand UO_2724 (O_2724,N_27393,N_26623);
xor UO_2725 (O_2725,N_29314,N_26195);
and UO_2726 (O_2726,N_27465,N_27149);
and UO_2727 (O_2727,N_25803,N_24343);
and UO_2728 (O_2728,N_29751,N_24266);
and UO_2729 (O_2729,N_24121,N_26550);
and UO_2730 (O_2730,N_24166,N_25158);
nand UO_2731 (O_2731,N_28709,N_26875);
nand UO_2732 (O_2732,N_29732,N_27915);
and UO_2733 (O_2733,N_29960,N_25798);
nor UO_2734 (O_2734,N_25826,N_26406);
nor UO_2735 (O_2735,N_26596,N_28145);
or UO_2736 (O_2736,N_27620,N_27989);
nor UO_2737 (O_2737,N_24897,N_26266);
nor UO_2738 (O_2738,N_24572,N_27799);
and UO_2739 (O_2739,N_25663,N_25819);
xor UO_2740 (O_2740,N_26403,N_29577);
or UO_2741 (O_2741,N_29122,N_28143);
nand UO_2742 (O_2742,N_24998,N_26844);
xor UO_2743 (O_2743,N_28650,N_24698);
and UO_2744 (O_2744,N_28045,N_27396);
nor UO_2745 (O_2745,N_25987,N_24874);
nand UO_2746 (O_2746,N_27127,N_26461);
nor UO_2747 (O_2747,N_28948,N_29378);
or UO_2748 (O_2748,N_29185,N_28720);
and UO_2749 (O_2749,N_29190,N_27117);
nand UO_2750 (O_2750,N_25068,N_28201);
or UO_2751 (O_2751,N_25512,N_25960);
nand UO_2752 (O_2752,N_29839,N_28617);
or UO_2753 (O_2753,N_26536,N_25973);
nand UO_2754 (O_2754,N_24695,N_27135);
xnor UO_2755 (O_2755,N_24021,N_24401);
nand UO_2756 (O_2756,N_26258,N_28379);
nand UO_2757 (O_2757,N_27370,N_29191);
and UO_2758 (O_2758,N_28198,N_29770);
nor UO_2759 (O_2759,N_28398,N_24485);
xnor UO_2760 (O_2760,N_25030,N_24106);
nor UO_2761 (O_2761,N_28307,N_29861);
and UO_2762 (O_2762,N_28376,N_27622);
and UO_2763 (O_2763,N_24990,N_29827);
nand UO_2764 (O_2764,N_27116,N_27092);
nand UO_2765 (O_2765,N_27376,N_24804);
nor UO_2766 (O_2766,N_28715,N_29621);
or UO_2767 (O_2767,N_25788,N_24154);
or UO_2768 (O_2768,N_25054,N_24301);
xnor UO_2769 (O_2769,N_26633,N_29212);
nor UO_2770 (O_2770,N_26588,N_28682);
nand UO_2771 (O_2771,N_28154,N_27727);
nand UO_2772 (O_2772,N_26207,N_25439);
xnor UO_2773 (O_2773,N_29439,N_26714);
and UO_2774 (O_2774,N_29243,N_27239);
and UO_2775 (O_2775,N_25049,N_27764);
and UO_2776 (O_2776,N_27440,N_29549);
and UO_2777 (O_2777,N_27236,N_24299);
xor UO_2778 (O_2778,N_25730,N_25631);
nor UO_2779 (O_2779,N_25215,N_24071);
nand UO_2780 (O_2780,N_26897,N_25431);
nand UO_2781 (O_2781,N_29956,N_26281);
nor UO_2782 (O_2782,N_24889,N_29996);
and UO_2783 (O_2783,N_26047,N_24139);
xnor UO_2784 (O_2784,N_25809,N_28525);
nor UO_2785 (O_2785,N_26700,N_27833);
nor UO_2786 (O_2786,N_29704,N_27834);
nand UO_2787 (O_2787,N_24920,N_29461);
and UO_2788 (O_2788,N_26214,N_29594);
nand UO_2789 (O_2789,N_25697,N_27538);
or UO_2790 (O_2790,N_29928,N_26342);
or UO_2791 (O_2791,N_27617,N_29136);
or UO_2792 (O_2792,N_24080,N_26323);
nand UO_2793 (O_2793,N_29870,N_26492);
nand UO_2794 (O_2794,N_25672,N_24540);
nor UO_2795 (O_2795,N_27377,N_24129);
xnor UO_2796 (O_2796,N_29350,N_29721);
or UO_2797 (O_2797,N_29328,N_29834);
or UO_2798 (O_2798,N_29390,N_26698);
xor UO_2799 (O_2799,N_29718,N_26136);
or UO_2800 (O_2800,N_26373,N_25041);
nand UO_2801 (O_2801,N_25471,N_24382);
nor UO_2802 (O_2802,N_27836,N_26785);
and UO_2803 (O_2803,N_24279,N_25927);
and UO_2804 (O_2804,N_24895,N_26368);
nand UO_2805 (O_2805,N_26033,N_29195);
nor UO_2806 (O_2806,N_26874,N_29778);
and UO_2807 (O_2807,N_24414,N_26443);
or UO_2808 (O_2808,N_29809,N_24611);
or UO_2809 (O_2809,N_24492,N_26848);
nor UO_2810 (O_2810,N_29947,N_27051);
and UO_2811 (O_2811,N_28717,N_28338);
nor UO_2812 (O_2812,N_25213,N_29119);
nand UO_2813 (O_2813,N_25477,N_29215);
nor UO_2814 (O_2814,N_27204,N_29160);
nand UO_2815 (O_2815,N_29306,N_26556);
nand UO_2816 (O_2816,N_29536,N_24026);
and UO_2817 (O_2817,N_29490,N_28283);
nor UO_2818 (O_2818,N_29746,N_24521);
and UO_2819 (O_2819,N_26181,N_24996);
nor UO_2820 (O_2820,N_25639,N_28513);
and UO_2821 (O_2821,N_28694,N_24956);
nor UO_2822 (O_2822,N_24516,N_24189);
xnor UO_2823 (O_2823,N_25198,N_26117);
xor UO_2824 (O_2824,N_29163,N_28495);
xor UO_2825 (O_2825,N_24449,N_26612);
and UO_2826 (O_2826,N_25986,N_29758);
nand UO_2827 (O_2827,N_25610,N_25200);
xor UO_2828 (O_2828,N_24631,N_27479);
and UO_2829 (O_2829,N_25513,N_26504);
nand UO_2830 (O_2830,N_26955,N_29767);
and UO_2831 (O_2831,N_29752,N_27486);
xnor UO_2832 (O_2832,N_29188,N_24808);
nor UO_2833 (O_2833,N_28559,N_25561);
nor UO_2834 (O_2834,N_28078,N_27752);
nand UO_2835 (O_2835,N_27375,N_29263);
xor UO_2836 (O_2836,N_29061,N_29909);
nor UO_2837 (O_2837,N_29550,N_27339);
nor UO_2838 (O_2838,N_26582,N_27265);
nand UO_2839 (O_2839,N_28780,N_24228);
and UO_2840 (O_2840,N_27334,N_29029);
or UO_2841 (O_2841,N_28645,N_28706);
nand UO_2842 (O_2842,N_25541,N_27701);
and UO_2843 (O_2843,N_24721,N_27929);
nor UO_2844 (O_2844,N_27193,N_29478);
and UO_2845 (O_2845,N_26340,N_29457);
and UO_2846 (O_2846,N_28691,N_28390);
nor UO_2847 (O_2847,N_24192,N_29329);
and UO_2848 (O_2848,N_29132,N_26251);
and UO_2849 (O_2849,N_27139,N_25578);
xor UO_2850 (O_2850,N_26723,N_27407);
xor UO_2851 (O_2851,N_25935,N_26361);
nor UO_2852 (O_2852,N_27849,N_28240);
and UO_2853 (O_2853,N_25647,N_25194);
and UO_2854 (O_2854,N_26662,N_24352);
and UO_2855 (O_2855,N_25998,N_29985);
or UO_2856 (O_2856,N_25917,N_26817);
and UO_2857 (O_2857,N_25591,N_28115);
or UO_2858 (O_2858,N_28578,N_27703);
and UO_2859 (O_2859,N_26659,N_28367);
nand UO_2860 (O_2860,N_28669,N_25903);
nand UO_2861 (O_2861,N_28782,N_29628);
or UO_2862 (O_2862,N_27437,N_29515);
or UO_2863 (O_2863,N_24670,N_26234);
or UO_2864 (O_2864,N_24329,N_27804);
or UO_2865 (O_2865,N_26956,N_28648);
or UO_2866 (O_2866,N_27649,N_29142);
xor UO_2867 (O_2867,N_28787,N_24429);
xnor UO_2868 (O_2868,N_26160,N_27582);
nor UO_2869 (O_2869,N_29115,N_28735);
nand UO_2870 (O_2870,N_28973,N_25858);
xnor UO_2871 (O_2871,N_28626,N_29842);
or UO_2872 (O_2872,N_26252,N_29696);
nand UO_2873 (O_2873,N_27528,N_24855);
or UO_2874 (O_2874,N_24946,N_27292);
nand UO_2875 (O_2875,N_28752,N_25224);
nand UO_2876 (O_2876,N_24696,N_27795);
and UO_2877 (O_2877,N_24437,N_27522);
and UO_2878 (O_2878,N_24461,N_29455);
nor UO_2879 (O_2879,N_28280,N_25853);
or UO_2880 (O_2880,N_28595,N_27867);
nand UO_2881 (O_2881,N_24780,N_29568);
and UO_2882 (O_2882,N_29370,N_26898);
xor UO_2883 (O_2883,N_26766,N_29963);
nor UO_2884 (O_2884,N_26819,N_27724);
or UO_2885 (O_2885,N_25778,N_25994);
and UO_2886 (O_2886,N_25700,N_28370);
or UO_2887 (O_2887,N_28898,N_24211);
nor UO_2888 (O_2888,N_28976,N_28040);
and UO_2889 (O_2889,N_29443,N_27985);
nor UO_2890 (O_2890,N_26097,N_25177);
nand UO_2891 (O_2891,N_26826,N_28053);
nor UO_2892 (O_2892,N_24642,N_24283);
xnor UO_2893 (O_2893,N_27118,N_28027);
and UO_2894 (O_2894,N_27248,N_27438);
or UO_2895 (O_2895,N_25228,N_25893);
or UO_2896 (O_2896,N_27077,N_24108);
nor UO_2897 (O_2897,N_27054,N_29633);
or UO_2898 (O_2898,N_25016,N_28470);
or UO_2899 (O_2899,N_25410,N_28519);
and UO_2900 (O_2900,N_27142,N_26000);
and UO_2901 (O_2901,N_27947,N_26424);
or UO_2902 (O_2902,N_25131,N_28071);
nand UO_2903 (O_2903,N_24689,N_24022);
or UO_2904 (O_2904,N_26085,N_27641);
or UO_2905 (O_2905,N_24320,N_24668);
nor UO_2906 (O_2906,N_28052,N_25279);
and UO_2907 (O_2907,N_28272,N_26391);
xnor UO_2908 (O_2908,N_27299,N_29437);
and UO_2909 (O_2909,N_24527,N_26689);
nand UO_2910 (O_2910,N_28125,N_27363);
and UO_2911 (O_2911,N_29769,N_28227);
or UO_2912 (O_2912,N_27793,N_29883);
xor UO_2913 (O_2913,N_25842,N_29091);
nand UO_2914 (O_2914,N_26682,N_29937);
or UO_2915 (O_2915,N_24966,N_25296);
and UO_2916 (O_2916,N_24514,N_29833);
or UO_2917 (O_2917,N_28416,N_24029);
xor UO_2918 (O_2918,N_25383,N_27285);
nand UO_2919 (O_2919,N_28514,N_25749);
and UO_2920 (O_2920,N_27994,N_29605);
and UO_2921 (O_2921,N_26592,N_25495);
xnor UO_2922 (O_2922,N_26670,N_25166);
and UO_2923 (O_2923,N_26135,N_26451);
and UO_2924 (O_2924,N_26104,N_25077);
xor UO_2925 (O_2925,N_27700,N_27852);
xor UO_2926 (O_2926,N_28074,N_25890);
nor UO_2927 (O_2927,N_27531,N_26876);
nor UO_2928 (O_2928,N_29011,N_24609);
nand UO_2929 (O_2929,N_24827,N_24369);
nand UO_2930 (O_2930,N_24373,N_24498);
or UO_2931 (O_2931,N_26547,N_26904);
nand UO_2932 (O_2932,N_25978,N_25366);
and UO_2933 (O_2933,N_26987,N_29005);
and UO_2934 (O_2934,N_25536,N_25570);
nand UO_2935 (O_2935,N_29289,N_28563);
nand UO_2936 (O_2936,N_27293,N_29831);
nand UO_2937 (O_2937,N_25707,N_24939);
nand UO_2938 (O_2938,N_29233,N_29731);
nand UO_2939 (O_2939,N_26910,N_26001);
and UO_2940 (O_2940,N_24407,N_24085);
nor UO_2941 (O_2941,N_25500,N_24638);
nor UO_2942 (O_2942,N_25845,N_26750);
nor UO_2943 (O_2943,N_27168,N_26832);
or UO_2944 (O_2944,N_28499,N_29196);
nor UO_2945 (O_2945,N_28167,N_28454);
or UO_2946 (O_2946,N_28955,N_28113);
nand UO_2947 (O_2947,N_25323,N_28149);
nor UO_2948 (O_2948,N_27509,N_26026);
xnor UO_2949 (O_2949,N_26453,N_26730);
or UO_2950 (O_2950,N_26747,N_29405);
xor UO_2951 (O_2951,N_25338,N_24763);
nor UO_2952 (O_2952,N_28486,N_27130);
nor UO_2953 (O_2953,N_27484,N_26610);
or UO_2954 (O_2954,N_27584,N_28838);
xnor UO_2955 (O_2955,N_26983,N_27143);
nand UO_2956 (O_2956,N_25270,N_24523);
nor UO_2957 (O_2957,N_29186,N_26993);
or UO_2958 (O_2958,N_26344,N_28255);
and UO_2959 (O_2959,N_27829,N_28869);
or UO_2960 (O_2960,N_26261,N_28137);
nor UO_2961 (O_2961,N_29853,N_25072);
nor UO_2962 (O_2962,N_28001,N_27181);
nor UO_2963 (O_2963,N_28657,N_28702);
nand UO_2964 (O_2964,N_28877,N_25519);
nand UO_2965 (O_2965,N_25613,N_28611);
xnor UO_2966 (O_2966,N_24857,N_24604);
nand UO_2967 (O_2967,N_27192,N_25874);
nand UO_2968 (O_2968,N_28730,N_26522);
and UO_2969 (O_2969,N_28982,N_28047);
xnor UO_2970 (O_2970,N_27250,N_25025);
xor UO_2971 (O_2971,N_26578,N_26928);
xnor UO_2972 (O_2972,N_24908,N_27543);
or UO_2973 (O_2973,N_27857,N_25625);
or UO_2974 (O_2974,N_25116,N_24103);
nand UO_2975 (O_2975,N_26115,N_26970);
and UO_2976 (O_2976,N_25324,N_26273);
nand UO_2977 (O_2977,N_26870,N_28474);
xor UO_2978 (O_2978,N_29015,N_28026);
xnor UO_2979 (O_2979,N_28351,N_29734);
nor UO_2980 (O_2980,N_29383,N_25099);
xor UO_2981 (O_2981,N_28770,N_26741);
or UO_2982 (O_2982,N_26186,N_25750);
and UO_2983 (O_2983,N_29255,N_27155);
nand UO_2984 (O_2984,N_28794,N_26028);
and UO_2985 (O_2985,N_29085,N_28038);
xnor UO_2986 (O_2986,N_24783,N_26869);
or UO_2987 (O_2987,N_26377,N_29983);
nor UO_2988 (O_2988,N_24589,N_28257);
nand UO_2989 (O_2989,N_29859,N_28189);
nand UO_2990 (O_2990,N_26378,N_25181);
or UO_2991 (O_2991,N_25813,N_28961);
or UO_2992 (O_2992,N_29873,N_26475);
nor UO_2993 (O_2993,N_28138,N_25848);
nor UO_2994 (O_2994,N_24556,N_26048);
xor UO_2995 (O_2995,N_24135,N_27352);
nand UO_2996 (O_2996,N_28541,N_29588);
or UO_2997 (O_2997,N_29938,N_24886);
xor UO_2998 (O_2998,N_27679,N_24048);
and UO_2999 (O_2999,N_24653,N_29720);
or UO_3000 (O_3000,N_25712,N_26290);
nor UO_3001 (O_3001,N_29234,N_29253);
or UO_3002 (O_3002,N_26677,N_25399);
nand UO_3003 (O_3003,N_24553,N_27157);
nor UO_3004 (O_3004,N_26436,N_26411);
xor UO_3005 (O_3005,N_26415,N_28487);
or UO_3006 (O_3006,N_27113,N_28896);
or UO_3007 (O_3007,N_27808,N_29084);
nor UO_3008 (O_3008,N_25965,N_28295);
or UO_3009 (O_3009,N_24412,N_24146);
xnor UO_3010 (O_3010,N_24530,N_24448);
nand UO_3011 (O_3011,N_25575,N_27460);
and UO_3012 (O_3012,N_27152,N_26509);
or UO_3013 (O_3013,N_28384,N_25031);
nor UO_3014 (O_3014,N_24581,N_25645);
xnor UO_3015 (O_3015,N_27687,N_24420);
or UO_3016 (O_3016,N_24961,N_28289);
xor UO_3017 (O_3017,N_28006,N_25191);
and UO_3018 (O_3018,N_25624,N_26568);
xor UO_3019 (O_3019,N_26824,N_25991);
and UO_3020 (O_3020,N_27546,N_26894);
xnor UO_3021 (O_3021,N_29590,N_24227);
nand UO_3022 (O_3022,N_25674,N_27889);
or UO_3023 (O_3023,N_26922,N_29574);
nor UO_3024 (O_3024,N_25995,N_26548);
nor UO_3025 (O_3025,N_25655,N_26292);
nor UO_3026 (O_3026,N_26356,N_25773);
nor UO_3027 (O_3027,N_25574,N_29167);
and UO_3028 (O_3028,N_28277,N_29932);
and UO_3029 (O_3029,N_27009,N_29502);
xor UO_3030 (O_3030,N_28080,N_28801);
or UO_3031 (O_3031,N_25225,N_27436);
nand UO_3032 (O_3032,N_26918,N_24210);
xnor UO_3033 (O_3033,N_27623,N_24000);
or UO_3034 (O_3034,N_26107,N_28446);
nand UO_3035 (O_3035,N_25450,N_28162);
nand UO_3036 (O_3036,N_24779,N_27841);
xnor UO_3037 (O_3037,N_26430,N_27407);
nand UO_3038 (O_3038,N_28229,N_26079);
nor UO_3039 (O_3039,N_24252,N_26782);
nor UO_3040 (O_3040,N_25273,N_24110);
or UO_3041 (O_3041,N_26008,N_26024);
and UO_3042 (O_3042,N_29366,N_24017);
and UO_3043 (O_3043,N_27682,N_24110);
nor UO_3044 (O_3044,N_28362,N_26932);
or UO_3045 (O_3045,N_29040,N_24385);
or UO_3046 (O_3046,N_27673,N_25122);
and UO_3047 (O_3047,N_24615,N_28203);
and UO_3048 (O_3048,N_29329,N_29082);
nor UO_3049 (O_3049,N_24529,N_28617);
xnor UO_3050 (O_3050,N_24792,N_27294);
xnor UO_3051 (O_3051,N_24900,N_28969);
nand UO_3052 (O_3052,N_26675,N_28166);
nand UO_3053 (O_3053,N_27326,N_27162);
and UO_3054 (O_3054,N_24598,N_29316);
nor UO_3055 (O_3055,N_27929,N_24305);
xor UO_3056 (O_3056,N_26819,N_28825);
and UO_3057 (O_3057,N_27378,N_25146);
nand UO_3058 (O_3058,N_24173,N_26051);
xor UO_3059 (O_3059,N_29025,N_24829);
nor UO_3060 (O_3060,N_25382,N_27631);
and UO_3061 (O_3061,N_28688,N_24204);
nand UO_3062 (O_3062,N_27267,N_28791);
or UO_3063 (O_3063,N_25011,N_24860);
nand UO_3064 (O_3064,N_24175,N_29086);
xor UO_3065 (O_3065,N_24775,N_27678);
nor UO_3066 (O_3066,N_26753,N_24885);
or UO_3067 (O_3067,N_28301,N_27789);
or UO_3068 (O_3068,N_28893,N_27310);
xnor UO_3069 (O_3069,N_29396,N_24648);
nor UO_3070 (O_3070,N_26388,N_25831);
or UO_3071 (O_3071,N_24946,N_27273);
nor UO_3072 (O_3072,N_28071,N_26292);
nor UO_3073 (O_3073,N_26362,N_29419);
nand UO_3074 (O_3074,N_28957,N_24368);
and UO_3075 (O_3075,N_27683,N_24720);
and UO_3076 (O_3076,N_26359,N_27656);
or UO_3077 (O_3077,N_28807,N_29064);
or UO_3078 (O_3078,N_24555,N_28707);
nor UO_3079 (O_3079,N_28031,N_26510);
nand UO_3080 (O_3080,N_25229,N_25744);
nand UO_3081 (O_3081,N_28133,N_26963);
xnor UO_3082 (O_3082,N_24201,N_28379);
and UO_3083 (O_3083,N_26334,N_24062);
and UO_3084 (O_3084,N_26305,N_29172);
and UO_3085 (O_3085,N_28835,N_29967);
or UO_3086 (O_3086,N_25929,N_24167);
nand UO_3087 (O_3087,N_28741,N_27799);
xnor UO_3088 (O_3088,N_29375,N_24365);
nor UO_3089 (O_3089,N_26125,N_25940);
nand UO_3090 (O_3090,N_24092,N_28766);
or UO_3091 (O_3091,N_29541,N_24894);
nor UO_3092 (O_3092,N_25446,N_28708);
nand UO_3093 (O_3093,N_28927,N_26582);
or UO_3094 (O_3094,N_24889,N_25345);
and UO_3095 (O_3095,N_26877,N_25607);
xnor UO_3096 (O_3096,N_29566,N_28436);
or UO_3097 (O_3097,N_26782,N_29576);
nor UO_3098 (O_3098,N_25081,N_25438);
and UO_3099 (O_3099,N_26864,N_24919);
or UO_3100 (O_3100,N_24812,N_29206);
or UO_3101 (O_3101,N_29893,N_29201);
and UO_3102 (O_3102,N_27284,N_27078);
xnor UO_3103 (O_3103,N_29704,N_26266);
or UO_3104 (O_3104,N_28357,N_28947);
xor UO_3105 (O_3105,N_29395,N_25438);
or UO_3106 (O_3106,N_25305,N_29732);
or UO_3107 (O_3107,N_29982,N_24322);
nor UO_3108 (O_3108,N_28000,N_24384);
xnor UO_3109 (O_3109,N_27472,N_26732);
nor UO_3110 (O_3110,N_28161,N_27286);
xor UO_3111 (O_3111,N_24948,N_25918);
nor UO_3112 (O_3112,N_27315,N_24260);
nor UO_3113 (O_3113,N_25257,N_28734);
xnor UO_3114 (O_3114,N_25909,N_24431);
or UO_3115 (O_3115,N_27405,N_29989);
or UO_3116 (O_3116,N_26594,N_29766);
xnor UO_3117 (O_3117,N_29383,N_25199);
and UO_3118 (O_3118,N_27882,N_26094);
and UO_3119 (O_3119,N_28327,N_27520);
xor UO_3120 (O_3120,N_27909,N_27472);
or UO_3121 (O_3121,N_27979,N_25695);
or UO_3122 (O_3122,N_25210,N_29071);
or UO_3123 (O_3123,N_25971,N_28360);
and UO_3124 (O_3124,N_29107,N_24300);
nand UO_3125 (O_3125,N_25359,N_26680);
nand UO_3126 (O_3126,N_25092,N_29258);
or UO_3127 (O_3127,N_29617,N_29486);
nand UO_3128 (O_3128,N_28774,N_28348);
nand UO_3129 (O_3129,N_29951,N_26941);
nand UO_3130 (O_3130,N_26250,N_28569);
nor UO_3131 (O_3131,N_26749,N_29337);
or UO_3132 (O_3132,N_28865,N_26991);
and UO_3133 (O_3133,N_29318,N_28779);
or UO_3134 (O_3134,N_24567,N_27807);
nand UO_3135 (O_3135,N_24832,N_29740);
and UO_3136 (O_3136,N_28361,N_27077);
xnor UO_3137 (O_3137,N_28030,N_29094);
nor UO_3138 (O_3138,N_26228,N_27393);
nor UO_3139 (O_3139,N_27106,N_26497);
nand UO_3140 (O_3140,N_26143,N_26361);
xor UO_3141 (O_3141,N_27359,N_27082);
and UO_3142 (O_3142,N_29026,N_27410);
or UO_3143 (O_3143,N_26353,N_26409);
xnor UO_3144 (O_3144,N_26626,N_28553);
and UO_3145 (O_3145,N_25976,N_28082);
or UO_3146 (O_3146,N_27575,N_27874);
xor UO_3147 (O_3147,N_25313,N_24847);
nand UO_3148 (O_3148,N_24192,N_27722);
nand UO_3149 (O_3149,N_26467,N_28184);
xor UO_3150 (O_3150,N_26045,N_25004);
and UO_3151 (O_3151,N_26558,N_28252);
nor UO_3152 (O_3152,N_25339,N_29363);
nor UO_3153 (O_3153,N_27652,N_28837);
or UO_3154 (O_3154,N_28152,N_28165);
or UO_3155 (O_3155,N_25849,N_27167);
nand UO_3156 (O_3156,N_25025,N_24137);
xnor UO_3157 (O_3157,N_29192,N_28664);
or UO_3158 (O_3158,N_26635,N_28848);
or UO_3159 (O_3159,N_29192,N_29339);
and UO_3160 (O_3160,N_26352,N_24745);
or UO_3161 (O_3161,N_29841,N_25803);
xnor UO_3162 (O_3162,N_25659,N_27406);
or UO_3163 (O_3163,N_25865,N_29071);
nor UO_3164 (O_3164,N_27408,N_27209);
xnor UO_3165 (O_3165,N_28129,N_29530);
and UO_3166 (O_3166,N_29498,N_28484);
nand UO_3167 (O_3167,N_25342,N_24515);
and UO_3168 (O_3168,N_25670,N_28564);
xor UO_3169 (O_3169,N_25380,N_25215);
nor UO_3170 (O_3170,N_26460,N_24359);
nor UO_3171 (O_3171,N_27555,N_29084);
nor UO_3172 (O_3172,N_27817,N_25638);
xor UO_3173 (O_3173,N_26912,N_24746);
or UO_3174 (O_3174,N_26935,N_25043);
or UO_3175 (O_3175,N_28487,N_28113);
and UO_3176 (O_3176,N_26515,N_28416);
or UO_3177 (O_3177,N_29659,N_29777);
or UO_3178 (O_3178,N_29680,N_25195);
or UO_3179 (O_3179,N_27478,N_29760);
and UO_3180 (O_3180,N_25301,N_28780);
or UO_3181 (O_3181,N_26231,N_26746);
nor UO_3182 (O_3182,N_29169,N_29428);
xnor UO_3183 (O_3183,N_27050,N_27794);
nor UO_3184 (O_3184,N_24442,N_29095);
nor UO_3185 (O_3185,N_27853,N_25808);
or UO_3186 (O_3186,N_27028,N_28535);
xor UO_3187 (O_3187,N_25146,N_25867);
nand UO_3188 (O_3188,N_24315,N_25232);
nand UO_3189 (O_3189,N_26069,N_26914);
or UO_3190 (O_3190,N_25150,N_26513);
or UO_3191 (O_3191,N_28444,N_29048);
nor UO_3192 (O_3192,N_27112,N_25500);
nor UO_3193 (O_3193,N_28456,N_24366);
nor UO_3194 (O_3194,N_29958,N_28219);
xnor UO_3195 (O_3195,N_24492,N_28558);
nor UO_3196 (O_3196,N_24007,N_25930);
xor UO_3197 (O_3197,N_24694,N_29118);
or UO_3198 (O_3198,N_27242,N_25995);
nand UO_3199 (O_3199,N_25164,N_27693);
xor UO_3200 (O_3200,N_25664,N_27479);
nand UO_3201 (O_3201,N_24765,N_28064);
and UO_3202 (O_3202,N_27776,N_28672);
nand UO_3203 (O_3203,N_27314,N_24898);
xor UO_3204 (O_3204,N_28208,N_25861);
nand UO_3205 (O_3205,N_28330,N_28899);
and UO_3206 (O_3206,N_29945,N_25101);
or UO_3207 (O_3207,N_26020,N_24522);
and UO_3208 (O_3208,N_26376,N_29219);
nor UO_3209 (O_3209,N_25594,N_27610);
xor UO_3210 (O_3210,N_26885,N_29773);
xor UO_3211 (O_3211,N_24876,N_24154);
or UO_3212 (O_3212,N_26320,N_26373);
or UO_3213 (O_3213,N_26288,N_25786);
nor UO_3214 (O_3214,N_27703,N_29637);
xnor UO_3215 (O_3215,N_28860,N_27242);
xnor UO_3216 (O_3216,N_27265,N_27771);
nand UO_3217 (O_3217,N_29225,N_29048);
or UO_3218 (O_3218,N_29801,N_24726);
or UO_3219 (O_3219,N_28691,N_25876);
or UO_3220 (O_3220,N_27138,N_29521);
and UO_3221 (O_3221,N_28898,N_26570);
nand UO_3222 (O_3222,N_26739,N_26726);
nand UO_3223 (O_3223,N_25430,N_24339);
and UO_3224 (O_3224,N_24591,N_28933);
or UO_3225 (O_3225,N_25073,N_27923);
nand UO_3226 (O_3226,N_28620,N_29501);
and UO_3227 (O_3227,N_24226,N_25836);
or UO_3228 (O_3228,N_29602,N_29735);
or UO_3229 (O_3229,N_26225,N_25355);
nor UO_3230 (O_3230,N_25276,N_25421);
nand UO_3231 (O_3231,N_24326,N_25525);
or UO_3232 (O_3232,N_24228,N_27505);
nor UO_3233 (O_3233,N_26576,N_27425);
nor UO_3234 (O_3234,N_29112,N_25719);
nor UO_3235 (O_3235,N_29379,N_26649);
and UO_3236 (O_3236,N_27803,N_29856);
and UO_3237 (O_3237,N_29876,N_26561);
xnor UO_3238 (O_3238,N_29861,N_29821);
and UO_3239 (O_3239,N_27841,N_24432);
and UO_3240 (O_3240,N_24116,N_25711);
or UO_3241 (O_3241,N_26365,N_24802);
nand UO_3242 (O_3242,N_25018,N_28638);
nand UO_3243 (O_3243,N_28684,N_25190);
or UO_3244 (O_3244,N_24418,N_29099);
xor UO_3245 (O_3245,N_24300,N_27210);
xnor UO_3246 (O_3246,N_25968,N_29824);
xor UO_3247 (O_3247,N_25620,N_25270);
xor UO_3248 (O_3248,N_29949,N_24571);
nand UO_3249 (O_3249,N_29566,N_27949);
nor UO_3250 (O_3250,N_24140,N_27816);
nand UO_3251 (O_3251,N_27162,N_29447);
nand UO_3252 (O_3252,N_24930,N_29937);
or UO_3253 (O_3253,N_26819,N_24944);
nor UO_3254 (O_3254,N_26147,N_25150);
nand UO_3255 (O_3255,N_27478,N_27668);
and UO_3256 (O_3256,N_25990,N_24473);
or UO_3257 (O_3257,N_26399,N_28664);
xor UO_3258 (O_3258,N_27786,N_25991);
or UO_3259 (O_3259,N_28015,N_29634);
nand UO_3260 (O_3260,N_28490,N_24289);
nor UO_3261 (O_3261,N_29373,N_28150);
xnor UO_3262 (O_3262,N_29770,N_26918);
and UO_3263 (O_3263,N_28314,N_25004);
xnor UO_3264 (O_3264,N_26169,N_28128);
and UO_3265 (O_3265,N_26906,N_25278);
nand UO_3266 (O_3266,N_28423,N_27939);
xor UO_3267 (O_3267,N_28878,N_27210);
and UO_3268 (O_3268,N_29285,N_27039);
xor UO_3269 (O_3269,N_24050,N_26344);
and UO_3270 (O_3270,N_27428,N_28538);
nand UO_3271 (O_3271,N_24525,N_26615);
and UO_3272 (O_3272,N_24948,N_28294);
xor UO_3273 (O_3273,N_27092,N_24015);
or UO_3274 (O_3274,N_29401,N_27054);
nand UO_3275 (O_3275,N_25873,N_29575);
nor UO_3276 (O_3276,N_27730,N_27403);
nor UO_3277 (O_3277,N_26026,N_24746);
and UO_3278 (O_3278,N_29761,N_24421);
nand UO_3279 (O_3279,N_24071,N_24539);
xnor UO_3280 (O_3280,N_25056,N_24788);
and UO_3281 (O_3281,N_28880,N_29536);
and UO_3282 (O_3282,N_29355,N_24760);
or UO_3283 (O_3283,N_27078,N_28975);
nor UO_3284 (O_3284,N_28710,N_29690);
nor UO_3285 (O_3285,N_25419,N_27150);
nand UO_3286 (O_3286,N_27615,N_25114);
or UO_3287 (O_3287,N_26947,N_29094);
nand UO_3288 (O_3288,N_25495,N_26470);
nor UO_3289 (O_3289,N_28647,N_28218);
nand UO_3290 (O_3290,N_28187,N_29050);
nor UO_3291 (O_3291,N_27657,N_26653);
nand UO_3292 (O_3292,N_26017,N_26634);
nand UO_3293 (O_3293,N_26222,N_26898);
xor UO_3294 (O_3294,N_25016,N_28771);
nand UO_3295 (O_3295,N_24565,N_24494);
and UO_3296 (O_3296,N_27794,N_26597);
and UO_3297 (O_3297,N_27517,N_28675);
and UO_3298 (O_3298,N_27603,N_28028);
nor UO_3299 (O_3299,N_28181,N_25768);
xor UO_3300 (O_3300,N_25464,N_26885);
or UO_3301 (O_3301,N_25885,N_25844);
and UO_3302 (O_3302,N_28944,N_29763);
or UO_3303 (O_3303,N_28614,N_29065);
and UO_3304 (O_3304,N_26204,N_25770);
or UO_3305 (O_3305,N_26196,N_29805);
and UO_3306 (O_3306,N_28938,N_25380);
and UO_3307 (O_3307,N_26323,N_24471);
or UO_3308 (O_3308,N_29463,N_24736);
or UO_3309 (O_3309,N_29659,N_25245);
or UO_3310 (O_3310,N_26764,N_26137);
nand UO_3311 (O_3311,N_25505,N_28475);
and UO_3312 (O_3312,N_27110,N_29209);
and UO_3313 (O_3313,N_26218,N_29241);
xor UO_3314 (O_3314,N_28332,N_24949);
and UO_3315 (O_3315,N_28413,N_28625);
or UO_3316 (O_3316,N_29775,N_26257);
and UO_3317 (O_3317,N_26090,N_26660);
nand UO_3318 (O_3318,N_28282,N_27722);
or UO_3319 (O_3319,N_27492,N_28915);
xor UO_3320 (O_3320,N_28235,N_25233);
and UO_3321 (O_3321,N_28550,N_27168);
or UO_3322 (O_3322,N_27962,N_27024);
or UO_3323 (O_3323,N_29715,N_25175);
xnor UO_3324 (O_3324,N_25248,N_25897);
and UO_3325 (O_3325,N_25326,N_24992);
and UO_3326 (O_3326,N_28993,N_24992);
nand UO_3327 (O_3327,N_27167,N_25080);
or UO_3328 (O_3328,N_29806,N_24974);
nand UO_3329 (O_3329,N_24532,N_24318);
xnor UO_3330 (O_3330,N_29491,N_26333);
or UO_3331 (O_3331,N_27963,N_24353);
and UO_3332 (O_3332,N_25666,N_26346);
nand UO_3333 (O_3333,N_27631,N_28092);
or UO_3334 (O_3334,N_25347,N_29925);
xor UO_3335 (O_3335,N_29483,N_26296);
xor UO_3336 (O_3336,N_29469,N_29945);
nand UO_3337 (O_3337,N_29290,N_27901);
nor UO_3338 (O_3338,N_26408,N_29667);
xnor UO_3339 (O_3339,N_27940,N_26932);
and UO_3340 (O_3340,N_24660,N_26278);
or UO_3341 (O_3341,N_27433,N_28157);
and UO_3342 (O_3342,N_24438,N_26336);
and UO_3343 (O_3343,N_24748,N_29739);
and UO_3344 (O_3344,N_25220,N_26670);
xnor UO_3345 (O_3345,N_26674,N_28761);
and UO_3346 (O_3346,N_26959,N_25561);
nand UO_3347 (O_3347,N_29183,N_26469);
and UO_3348 (O_3348,N_27415,N_25876);
xor UO_3349 (O_3349,N_27765,N_27872);
nor UO_3350 (O_3350,N_28104,N_27117);
nor UO_3351 (O_3351,N_26578,N_27518);
nand UO_3352 (O_3352,N_29945,N_24492);
xor UO_3353 (O_3353,N_27514,N_29670);
or UO_3354 (O_3354,N_28979,N_27969);
nand UO_3355 (O_3355,N_26616,N_28773);
nor UO_3356 (O_3356,N_27250,N_26197);
nand UO_3357 (O_3357,N_27327,N_27101);
nor UO_3358 (O_3358,N_25259,N_26916);
xnor UO_3359 (O_3359,N_26009,N_29870);
and UO_3360 (O_3360,N_29605,N_27876);
and UO_3361 (O_3361,N_28324,N_27922);
xor UO_3362 (O_3362,N_26183,N_26524);
and UO_3363 (O_3363,N_28327,N_25845);
xor UO_3364 (O_3364,N_29484,N_24527);
xnor UO_3365 (O_3365,N_28011,N_26456);
and UO_3366 (O_3366,N_27276,N_27246);
and UO_3367 (O_3367,N_25616,N_25492);
xor UO_3368 (O_3368,N_28312,N_25210);
or UO_3369 (O_3369,N_26219,N_26067);
or UO_3370 (O_3370,N_27444,N_24648);
or UO_3371 (O_3371,N_27883,N_25716);
xor UO_3372 (O_3372,N_26121,N_25220);
nand UO_3373 (O_3373,N_28207,N_24879);
nand UO_3374 (O_3374,N_28638,N_24524);
xnor UO_3375 (O_3375,N_27179,N_29005);
nor UO_3376 (O_3376,N_26569,N_29737);
nand UO_3377 (O_3377,N_28521,N_27761);
nand UO_3378 (O_3378,N_25734,N_28572);
nor UO_3379 (O_3379,N_28065,N_27667);
or UO_3380 (O_3380,N_24283,N_28766);
nor UO_3381 (O_3381,N_24099,N_27654);
nor UO_3382 (O_3382,N_27561,N_25492);
or UO_3383 (O_3383,N_25795,N_28982);
nand UO_3384 (O_3384,N_24686,N_26657);
xor UO_3385 (O_3385,N_24241,N_28042);
or UO_3386 (O_3386,N_29221,N_25136);
nor UO_3387 (O_3387,N_29403,N_27933);
or UO_3388 (O_3388,N_29755,N_25732);
and UO_3389 (O_3389,N_26102,N_26049);
or UO_3390 (O_3390,N_25950,N_27044);
nor UO_3391 (O_3391,N_28338,N_28795);
and UO_3392 (O_3392,N_26656,N_24120);
nand UO_3393 (O_3393,N_25877,N_29270);
nand UO_3394 (O_3394,N_29092,N_27433);
and UO_3395 (O_3395,N_26109,N_26405);
and UO_3396 (O_3396,N_28566,N_26880);
xor UO_3397 (O_3397,N_29378,N_24725);
nand UO_3398 (O_3398,N_27212,N_26917);
nand UO_3399 (O_3399,N_29418,N_25172);
xnor UO_3400 (O_3400,N_24408,N_25699);
and UO_3401 (O_3401,N_27319,N_25859);
nor UO_3402 (O_3402,N_26233,N_29034);
xor UO_3403 (O_3403,N_24256,N_29002);
and UO_3404 (O_3404,N_28988,N_29307);
nor UO_3405 (O_3405,N_28422,N_24065);
or UO_3406 (O_3406,N_27494,N_27235);
or UO_3407 (O_3407,N_25288,N_25804);
or UO_3408 (O_3408,N_24938,N_24702);
or UO_3409 (O_3409,N_29082,N_27036);
nor UO_3410 (O_3410,N_25502,N_28612);
nor UO_3411 (O_3411,N_24513,N_29681);
and UO_3412 (O_3412,N_25840,N_26903);
and UO_3413 (O_3413,N_24117,N_29295);
nor UO_3414 (O_3414,N_25802,N_27147);
and UO_3415 (O_3415,N_25715,N_29976);
xor UO_3416 (O_3416,N_25839,N_29628);
and UO_3417 (O_3417,N_29120,N_28875);
xor UO_3418 (O_3418,N_28765,N_27409);
or UO_3419 (O_3419,N_27431,N_25958);
or UO_3420 (O_3420,N_25400,N_28553);
nand UO_3421 (O_3421,N_27642,N_28766);
xor UO_3422 (O_3422,N_26604,N_26704);
or UO_3423 (O_3423,N_29925,N_24518);
or UO_3424 (O_3424,N_27782,N_24115);
nor UO_3425 (O_3425,N_29414,N_29118);
or UO_3426 (O_3426,N_24607,N_29136);
or UO_3427 (O_3427,N_27953,N_24128);
xnor UO_3428 (O_3428,N_26151,N_28225);
and UO_3429 (O_3429,N_28570,N_29916);
and UO_3430 (O_3430,N_25344,N_28549);
or UO_3431 (O_3431,N_25039,N_25501);
xor UO_3432 (O_3432,N_26082,N_24373);
and UO_3433 (O_3433,N_24485,N_29414);
and UO_3434 (O_3434,N_25120,N_28853);
or UO_3435 (O_3435,N_25551,N_25292);
or UO_3436 (O_3436,N_29992,N_24269);
and UO_3437 (O_3437,N_29647,N_28165);
or UO_3438 (O_3438,N_25182,N_27361);
nor UO_3439 (O_3439,N_24566,N_28443);
and UO_3440 (O_3440,N_24840,N_26922);
xnor UO_3441 (O_3441,N_26889,N_27655);
nand UO_3442 (O_3442,N_24986,N_26093);
xnor UO_3443 (O_3443,N_26528,N_26808);
nand UO_3444 (O_3444,N_25496,N_28572);
nand UO_3445 (O_3445,N_28562,N_28171);
nand UO_3446 (O_3446,N_29035,N_24196);
nand UO_3447 (O_3447,N_24107,N_28470);
nor UO_3448 (O_3448,N_29752,N_26230);
nand UO_3449 (O_3449,N_25375,N_28544);
nor UO_3450 (O_3450,N_24011,N_25194);
nand UO_3451 (O_3451,N_26793,N_26360);
nor UO_3452 (O_3452,N_28810,N_24198);
nor UO_3453 (O_3453,N_29220,N_29006);
nand UO_3454 (O_3454,N_26204,N_28996);
or UO_3455 (O_3455,N_25504,N_27216);
nand UO_3456 (O_3456,N_27114,N_29655);
nand UO_3457 (O_3457,N_24430,N_29602);
or UO_3458 (O_3458,N_29702,N_28178);
or UO_3459 (O_3459,N_28617,N_26131);
xnor UO_3460 (O_3460,N_26263,N_24702);
and UO_3461 (O_3461,N_27555,N_29381);
xor UO_3462 (O_3462,N_28220,N_24941);
nor UO_3463 (O_3463,N_26138,N_24908);
or UO_3464 (O_3464,N_25170,N_24449);
nand UO_3465 (O_3465,N_26756,N_26586);
nor UO_3466 (O_3466,N_27340,N_25826);
or UO_3467 (O_3467,N_24791,N_27382);
nor UO_3468 (O_3468,N_29686,N_26665);
xnor UO_3469 (O_3469,N_24771,N_29574);
nor UO_3470 (O_3470,N_24332,N_26385);
nand UO_3471 (O_3471,N_26728,N_29565);
xor UO_3472 (O_3472,N_28880,N_26565);
nor UO_3473 (O_3473,N_26040,N_28657);
nor UO_3474 (O_3474,N_24053,N_25702);
nand UO_3475 (O_3475,N_29860,N_25557);
nor UO_3476 (O_3476,N_26149,N_24658);
and UO_3477 (O_3477,N_25003,N_26860);
and UO_3478 (O_3478,N_27856,N_25526);
nand UO_3479 (O_3479,N_27630,N_25935);
or UO_3480 (O_3480,N_27728,N_27215);
and UO_3481 (O_3481,N_25711,N_25538);
xnor UO_3482 (O_3482,N_26286,N_29519);
nor UO_3483 (O_3483,N_26143,N_26077);
and UO_3484 (O_3484,N_28401,N_26155);
or UO_3485 (O_3485,N_26576,N_28664);
xor UO_3486 (O_3486,N_28802,N_27397);
or UO_3487 (O_3487,N_25942,N_28182);
and UO_3488 (O_3488,N_26526,N_25386);
and UO_3489 (O_3489,N_24218,N_27555);
nor UO_3490 (O_3490,N_24670,N_24369);
xor UO_3491 (O_3491,N_28134,N_25172);
and UO_3492 (O_3492,N_28702,N_28050);
nor UO_3493 (O_3493,N_29954,N_25385);
xnor UO_3494 (O_3494,N_29828,N_29175);
or UO_3495 (O_3495,N_28644,N_29845);
nor UO_3496 (O_3496,N_25543,N_29168);
and UO_3497 (O_3497,N_29563,N_29277);
nand UO_3498 (O_3498,N_24097,N_26850);
and UO_3499 (O_3499,N_24283,N_29805);
endmodule