module basic_3000_30000_3500_6_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_964,In_467);
nor U1 (N_1,In_487,In_446);
xnor U2 (N_2,In_2412,In_320);
nand U3 (N_3,In_1362,In_201);
nand U4 (N_4,In_1354,In_594);
nor U5 (N_5,In_1745,In_191);
nand U6 (N_6,In_2939,In_628);
or U7 (N_7,In_2820,In_2961);
and U8 (N_8,In_2036,In_491);
nand U9 (N_9,In_225,In_2078);
or U10 (N_10,In_1669,In_1792);
nand U11 (N_11,In_1475,In_2760);
nor U12 (N_12,In_1161,In_389);
or U13 (N_13,In_1197,In_1743);
xor U14 (N_14,In_2902,In_1205);
xor U15 (N_15,In_58,In_40);
and U16 (N_16,In_2013,In_1509);
xor U17 (N_17,In_97,In_2573);
nor U18 (N_18,In_439,In_277);
nor U19 (N_19,In_131,In_848);
nor U20 (N_20,In_256,In_2827);
nor U21 (N_21,In_755,In_2201);
nor U22 (N_22,In_2814,In_1382);
or U23 (N_23,In_1346,In_2192);
xnor U24 (N_24,In_2246,In_2987);
nor U25 (N_25,In_2588,In_987);
nand U26 (N_26,In_994,In_285);
or U27 (N_27,In_1704,In_2023);
and U28 (N_28,In_1414,In_856);
xor U29 (N_29,In_2066,In_773);
or U30 (N_30,In_1785,In_2236);
and U31 (N_31,In_1646,In_45);
xnor U32 (N_32,In_2449,In_2697);
nand U33 (N_33,In_378,In_1962);
or U34 (N_34,In_2642,In_1891);
nand U35 (N_35,In_2934,In_2223);
and U36 (N_36,In_1630,In_612);
xor U37 (N_37,In_681,In_1210);
or U38 (N_38,In_319,In_2615);
nor U39 (N_39,In_128,In_1367);
xor U40 (N_40,In_1181,In_957);
and U41 (N_41,In_2206,In_2275);
nor U42 (N_42,In_2751,In_2346);
and U43 (N_43,In_1040,In_2297);
xnor U44 (N_44,In_728,In_995);
or U45 (N_45,In_1126,In_824);
and U46 (N_46,In_1165,In_1659);
nor U47 (N_47,In_2869,In_413);
xnor U48 (N_48,In_151,In_1162);
or U49 (N_49,In_2128,In_948);
nor U50 (N_50,In_1811,In_2841);
or U51 (N_51,In_461,In_1959);
or U52 (N_52,In_377,In_1653);
or U53 (N_53,In_1264,In_1964);
nor U54 (N_54,In_1731,In_2423);
and U55 (N_55,In_163,In_65);
or U56 (N_56,In_1960,In_2606);
or U57 (N_57,In_1238,In_571);
xor U58 (N_58,In_214,In_2837);
xnor U59 (N_59,In_1520,In_203);
xor U60 (N_60,In_2115,In_1784);
nand U61 (N_61,In_2187,In_1584);
xnor U62 (N_62,In_2565,In_2469);
nor U63 (N_63,In_423,In_313);
xor U64 (N_64,In_933,In_1045);
nand U65 (N_65,In_1466,In_2408);
and U66 (N_66,In_1936,In_2217);
or U67 (N_67,In_295,In_1693);
xnor U68 (N_68,In_1638,In_325);
nor U69 (N_69,In_1775,In_2307);
nand U70 (N_70,In_1338,In_2477);
nor U71 (N_71,In_1231,In_1364);
nand U72 (N_72,In_2547,In_2755);
nor U73 (N_73,In_1433,In_798);
nor U74 (N_74,In_144,In_1881);
nand U75 (N_75,In_963,In_1718);
and U76 (N_76,In_2543,In_2222);
nor U77 (N_77,In_2124,In_509);
and U78 (N_78,In_85,In_1921);
or U79 (N_79,In_260,In_958);
xnor U80 (N_80,In_1139,In_35);
nand U81 (N_81,In_1858,In_1472);
xor U82 (N_82,In_54,In_1948);
nor U83 (N_83,In_2836,In_1174);
and U84 (N_84,In_2185,In_323);
nand U85 (N_85,In_1122,In_2501);
or U86 (N_86,In_1402,In_1533);
nand U87 (N_87,In_2823,In_2004);
or U88 (N_88,In_2510,In_2541);
nand U89 (N_89,In_1110,In_481);
or U90 (N_90,In_1285,In_1783);
nor U91 (N_91,In_2105,In_2978);
nand U92 (N_92,In_101,In_1493);
xor U93 (N_93,In_826,In_741);
xor U94 (N_94,In_2070,In_1813);
or U95 (N_95,In_1305,In_2988);
or U96 (N_96,In_768,In_109);
xor U97 (N_97,In_2917,In_1702);
xnor U98 (N_98,In_1739,In_2787);
nand U99 (N_99,In_1989,In_2673);
nor U100 (N_100,In_2754,In_838);
nor U101 (N_101,In_813,In_2694);
or U102 (N_102,In_2738,In_789);
and U103 (N_103,In_1986,In_684);
and U104 (N_104,In_2003,In_662);
nor U105 (N_105,In_412,In_1882);
or U106 (N_106,In_2047,In_1768);
xnor U107 (N_107,In_2896,In_837);
or U108 (N_108,In_2269,In_1932);
and U109 (N_109,In_244,In_447);
nor U110 (N_110,In_125,In_2957);
nor U111 (N_111,In_1085,In_1298);
nor U112 (N_112,In_2445,In_2624);
xnor U113 (N_113,In_2798,In_1257);
nand U114 (N_114,In_2998,In_978);
nor U115 (N_115,In_479,In_2895);
or U116 (N_116,In_2635,In_660);
xor U117 (N_117,In_1939,In_2580);
or U118 (N_118,In_2639,In_1381);
and U119 (N_119,In_2537,In_1824);
nand U120 (N_120,In_2599,In_2968);
and U121 (N_121,In_137,In_2671);
and U122 (N_122,In_2420,In_832);
and U123 (N_123,In_827,In_259);
nor U124 (N_124,In_1322,In_67);
nor U125 (N_125,In_213,In_272);
nand U126 (N_126,In_1913,In_1129);
nand U127 (N_127,In_1571,In_921);
nor U128 (N_128,In_2052,In_1582);
nand U129 (N_129,In_230,In_1919);
nand U130 (N_130,In_1312,In_11);
or U131 (N_131,In_115,In_1725);
xor U132 (N_132,In_2970,In_513);
or U133 (N_133,In_956,In_2308);
nand U134 (N_134,In_2190,In_120);
and U135 (N_135,In_2109,In_440);
or U136 (N_136,In_2072,In_1395);
xor U137 (N_137,In_76,In_1209);
and U138 (N_138,In_1855,In_1862);
nor U139 (N_139,In_2750,In_1606);
and U140 (N_140,In_945,In_2782);
or U141 (N_141,In_1325,In_1689);
nand U142 (N_142,In_2597,In_2436);
or U143 (N_143,In_1971,In_1415);
nor U144 (N_144,In_1546,In_2323);
xor U145 (N_145,In_673,In_1608);
and U146 (N_146,In_1189,In_274);
nand U147 (N_147,In_2773,In_2886);
nand U148 (N_148,In_2908,In_1452);
and U149 (N_149,In_2168,In_2688);
nor U150 (N_150,In_2370,In_1044);
nand U151 (N_151,In_2108,In_2058);
or U152 (N_152,In_1931,In_533);
and U153 (N_153,In_2144,In_1972);
and U154 (N_154,In_1933,In_414);
or U155 (N_155,In_1042,In_1898);
and U156 (N_156,In_383,In_2653);
xnor U157 (N_157,In_1192,In_627);
nor U158 (N_158,In_502,In_693);
nor U159 (N_159,In_2858,In_2355);
and U160 (N_160,In_2389,In_672);
nor U161 (N_161,In_2561,In_1570);
xnor U162 (N_162,In_2162,In_1559);
nor U163 (N_163,In_2527,In_843);
or U164 (N_164,In_1769,In_1518);
nand U165 (N_165,In_658,In_477);
and U166 (N_166,In_2329,In_405);
nand U167 (N_167,In_2595,In_2045);
nand U168 (N_168,In_1761,In_62);
nor U169 (N_169,In_550,In_1900);
nor U170 (N_170,In_2708,In_2009);
xor U171 (N_171,In_241,In_1899);
and U172 (N_172,In_2517,In_1666);
nor U173 (N_173,In_124,In_936);
or U174 (N_174,In_872,In_1937);
nand U175 (N_175,In_1539,In_1097);
nand U176 (N_176,In_2163,In_1757);
nor U177 (N_177,In_2320,In_90);
nor U178 (N_178,In_38,In_2313);
or U179 (N_179,In_1534,In_2359);
nor U180 (N_180,In_1039,In_44);
xor U181 (N_181,In_2812,In_2690);
nor U182 (N_182,In_2431,In_2172);
nor U183 (N_183,In_2603,In_2404);
nand U184 (N_184,In_2055,In_2270);
and U185 (N_185,In_2110,In_1998);
and U186 (N_186,In_2267,In_2796);
or U187 (N_187,In_404,In_165);
nor U188 (N_188,In_685,In_2202);
and U189 (N_189,In_1526,In_2845);
and U190 (N_190,In_1572,In_1328);
xnor U191 (N_191,In_1084,In_1537);
nor U192 (N_192,In_2979,In_489);
or U193 (N_193,In_71,In_2347);
xor U194 (N_194,In_703,In_1755);
nand U195 (N_195,In_2513,In_1934);
and U196 (N_196,In_1625,In_2214);
or U197 (N_197,In_2067,In_1491);
and U198 (N_198,In_1014,In_1116);
and U199 (N_199,In_305,In_1842);
xor U200 (N_200,In_1615,In_2038);
nor U201 (N_201,In_2646,In_1236);
nor U202 (N_202,In_2973,In_2175);
xor U203 (N_203,In_522,In_2799);
and U204 (N_204,In_951,In_356);
nor U205 (N_205,In_39,In_1549);
nor U206 (N_206,In_663,In_2479);
and U207 (N_207,In_2789,In_2197);
nor U208 (N_208,In_2061,In_2676);
xor U209 (N_209,In_2865,In_456);
nand U210 (N_210,In_136,In_417);
and U211 (N_211,In_1123,In_1379);
xnor U212 (N_212,In_1887,In_188);
and U213 (N_213,In_1418,In_910);
xnor U214 (N_214,In_877,In_1383);
nand U215 (N_215,In_2963,In_1973);
nand U216 (N_216,In_1166,In_424);
nor U217 (N_217,In_2576,In_2638);
nand U218 (N_218,In_2314,In_1480);
or U219 (N_219,In_2169,In_1476);
and U220 (N_220,In_196,In_1249);
nand U221 (N_221,In_2393,In_1851);
and U222 (N_222,In_2416,In_2553);
and U223 (N_223,In_1431,In_1007);
nand U224 (N_224,In_1635,In_2919);
and U225 (N_225,In_1751,In_1233);
xor U226 (N_226,In_2873,In_2195);
and U227 (N_227,In_633,In_1499);
or U228 (N_228,In_155,In_1911);
or U229 (N_229,In_527,In_2016);
xnor U230 (N_230,In_238,In_716);
nand U231 (N_231,In_1034,In_326);
and U232 (N_232,In_2288,In_1797);
and U233 (N_233,In_2994,In_1309);
or U234 (N_234,In_1096,In_1175);
and U235 (N_235,In_46,In_1154);
nand U236 (N_236,In_2732,In_1623);
and U237 (N_237,In_640,In_1894);
nor U238 (N_238,In_1023,In_270);
nor U239 (N_239,In_499,In_2361);
or U240 (N_240,In_1113,In_205);
xnor U241 (N_241,In_2680,In_1202);
nand U242 (N_242,In_2198,In_867);
nand U243 (N_243,In_2867,In_2103);
nor U244 (N_244,In_1070,In_2051);
nand U245 (N_245,In_2304,In_772);
nor U246 (N_246,In_2578,In_1760);
nor U247 (N_247,In_381,In_687);
and U248 (N_248,In_403,In_1287);
nand U249 (N_249,In_2667,In_606);
nor U250 (N_250,In_1482,In_2659);
nor U251 (N_251,In_1676,In_2443);
nor U252 (N_252,In_587,In_2399);
and U253 (N_253,In_806,In_2749);
or U254 (N_254,In_2180,In_985);
nand U255 (N_255,In_1341,In_2560);
or U256 (N_256,In_1829,In_1050);
or U257 (N_257,In_2158,In_1943);
and U258 (N_258,In_1944,In_742);
nor U259 (N_259,In_1140,In_1917);
nor U260 (N_260,In_1796,In_754);
and U261 (N_261,In_2480,In_445);
xnor U262 (N_262,In_862,In_2181);
nand U263 (N_263,In_1598,In_431);
nor U264 (N_264,In_661,In_746);
or U265 (N_265,In_2330,In_1317);
xor U266 (N_266,In_1263,In_949);
nand U267 (N_267,In_586,In_118);
and U268 (N_268,In_2113,In_81);
nor U269 (N_269,In_2118,In_2126);
nand U270 (N_270,In_829,In_1353);
nand U271 (N_271,In_2063,In_1759);
and U272 (N_272,In_2995,In_1552);
nor U273 (N_273,In_63,In_740);
xnor U274 (N_274,In_1201,In_2208);
nor U275 (N_275,In_1164,In_2127);
nor U276 (N_276,In_1244,In_1949);
or U277 (N_277,In_1701,In_1600);
nor U278 (N_278,In_2752,In_1333);
or U279 (N_279,In_2005,In_2074);
or U280 (N_280,In_950,In_1650);
xnor U281 (N_281,In_2859,In_2306);
or U282 (N_282,In_600,In_722);
and U283 (N_283,In_1009,In_2333);
xnor U284 (N_284,In_184,In_1270);
nand U285 (N_285,In_222,In_273);
nor U286 (N_286,In_1788,In_52);
or U287 (N_287,In_2327,In_940);
nand U288 (N_288,In_1372,In_625);
or U289 (N_289,In_2631,In_654);
nand U290 (N_290,In_1710,In_2952);
nand U291 (N_291,In_327,In_2101);
xnor U292 (N_292,In_1074,In_2784);
nor U293 (N_293,In_296,In_1684);
nor U294 (N_294,In_2097,In_1246);
nand U295 (N_295,In_1284,In_1321);
nand U296 (N_296,In_1531,In_2766);
and U297 (N_297,In_2834,In_2381);
nand U298 (N_298,In_2929,In_1920);
and U299 (N_299,In_2022,In_2001);
xor U300 (N_300,In_1016,In_6);
and U301 (N_301,In_917,In_2286);
nor U302 (N_302,In_1611,In_2473);
xnor U303 (N_303,In_2511,In_1473);
and U304 (N_304,In_466,In_2460);
nand U305 (N_305,In_2419,In_1734);
and U306 (N_306,In_26,In_737);
nor U307 (N_307,In_408,In_31);
and U308 (N_308,In_1738,In_2388);
or U309 (N_309,In_1506,In_175);
nand U310 (N_310,In_1727,In_2540);
nor U311 (N_311,In_421,In_1432);
xor U312 (N_312,In_1425,In_2364);
nand U313 (N_313,In_1063,In_392);
and U314 (N_314,In_2215,In_1683);
nor U315 (N_315,In_1370,In_2133);
xor U316 (N_316,In_2077,In_849);
xor U317 (N_317,In_1218,In_1868);
nand U318 (N_318,In_2941,In_2098);
nor U319 (N_319,In_1416,In_1407);
xor U320 (N_320,In_459,In_1156);
and U321 (N_321,In_2685,In_2619);
nor U322 (N_322,In_449,In_2387);
and U323 (N_323,In_161,In_2535);
or U324 (N_324,In_1400,In_472);
or U325 (N_325,In_1885,In_1524);
xnor U326 (N_326,In_651,In_1670);
and U327 (N_327,In_2592,In_2139);
xnor U328 (N_328,In_1765,In_1294);
nand U329 (N_329,In_2674,In_2644);
or U330 (N_330,In_2049,In_1131);
xor U331 (N_331,In_1545,In_2122);
nand U332 (N_332,In_898,In_825);
xnor U333 (N_333,In_64,In_552);
and U334 (N_334,In_1267,In_409);
and U335 (N_335,In_1588,In_1691);
and U336 (N_336,In_2526,In_536);
nand U337 (N_337,In_2675,In_2735);
nor U338 (N_338,In_2153,In_396);
xor U339 (N_339,In_1836,In_2769);
nor U340 (N_340,In_2946,In_2062);
nand U341 (N_341,In_180,In_2825);
xor U342 (N_342,In_2844,In_79);
nand U343 (N_343,In_1922,In_2522);
nand U344 (N_344,In_1951,In_2587);
xnor U345 (N_345,In_1368,In_2012);
and U346 (N_346,In_2807,In_1032);
and U347 (N_347,In_1248,In_756);
and U348 (N_348,In_2090,In_518);
and U349 (N_349,In_762,In_217);
xnor U350 (N_350,In_300,In_2373);
xor U351 (N_351,In_710,In_873);
nand U352 (N_352,In_2462,In_1150);
nand U353 (N_353,In_194,In_100);
or U354 (N_354,In_1791,In_2475);
xnor U355 (N_355,In_23,In_232);
or U356 (N_356,In_1490,In_2997);
or U357 (N_357,In_1709,In_1143);
xor U358 (N_358,In_1215,In_1144);
nor U359 (N_359,In_2885,In_726);
nand U360 (N_360,In_360,In_1777);
and U361 (N_361,In_521,In_2779);
nand U362 (N_362,In_2811,In_3);
or U363 (N_363,In_1436,In_468);
and U364 (N_364,In_271,In_2745);
nand U365 (N_365,In_1581,In_1983);
nand U366 (N_366,In_2343,In_2372);
nand U367 (N_367,In_2380,In_1928);
nor U368 (N_368,In_601,In_1121);
xnor U369 (N_369,In_869,In_2200);
and U370 (N_370,In_1186,In_442);
xor U371 (N_371,In_1619,In_349);
nand U372 (N_372,In_1345,In_1396);
xor U373 (N_373,In_1057,In_2991);
nand U374 (N_374,In_1974,In_564);
and U375 (N_375,In_1655,In_493);
nor U376 (N_376,In_1182,In_1035);
xor U377 (N_377,In_1066,In_2935);
nand U378 (N_378,In_344,In_1946);
and U379 (N_379,In_152,In_769);
or U380 (N_380,In_2657,In_2669);
and U381 (N_381,In_2803,In_558);
nand U382 (N_382,In_1266,In_858);
nor U383 (N_383,In_2360,In_2203);
or U384 (N_384,In_237,In_2089);
xnor U385 (N_385,In_610,In_671);
nand U386 (N_386,In_724,In_1318);
nor U387 (N_387,In_1498,In_1277);
or U388 (N_388,In_1487,In_250);
nor U389 (N_389,In_840,In_1782);
nor U390 (N_390,In_1258,In_1105);
or U391 (N_391,In_2140,In_2944);
nand U392 (N_392,In_365,In_2582);
nor U393 (N_393,In_1966,In_1153);
nor U394 (N_394,In_293,In_2876);
and U395 (N_395,In_939,In_140);
nor U396 (N_396,In_547,In_2188);
and U397 (N_397,In_452,In_433);
nor U398 (N_398,In_387,In_2171);
xnor U399 (N_399,In_1477,In_1580);
xor U400 (N_400,In_2672,In_264);
nand U401 (N_401,In_2032,In_1622);
nor U402 (N_402,In_1820,In_704);
or U403 (N_403,In_1896,In_2562);
or U404 (N_404,In_534,In_1527);
nor U405 (N_405,In_1386,In_1827);
or U406 (N_406,In_2174,In_2441);
nand U407 (N_407,In_331,In_1320);
nor U408 (N_408,In_690,In_1401);
or U409 (N_409,In_595,In_2602);
xor U410 (N_410,In_2641,In_2383);
xnor U411 (N_411,In_894,In_596);
xnor U412 (N_412,In_2239,In_799);
or U413 (N_413,In_2046,In_164);
nor U414 (N_414,In_1628,In_2989);
nor U415 (N_415,In_650,In_246);
and U416 (N_416,In_2268,In_1224);
nand U417 (N_417,In_620,In_2992);
or U418 (N_418,In_2287,In_1594);
or U419 (N_419,In_678,In_2808);
nand U420 (N_420,In_2965,In_1102);
nor U421 (N_421,In_761,In_2753);
nand U422 (N_422,In_1686,In_80);
nand U423 (N_423,In_707,In_2913);
and U424 (N_424,In_2699,In_2147);
or U425 (N_425,In_2775,In_993);
nor U426 (N_426,In_566,In_2583);
or U427 (N_427,In_511,In_388);
or U428 (N_428,In_1682,In_2628);
nor U429 (N_429,In_2593,In_683);
or U430 (N_430,In_2618,In_2901);
and U431 (N_431,In_460,In_2468);
nand U432 (N_432,In_2345,In_2506);
nor U433 (N_433,In_1523,In_1601);
nand U434 (N_434,In_1004,In_1672);
or U435 (N_435,In_169,In_1111);
nand U436 (N_436,In_2733,In_2783);
xor U437 (N_437,In_2568,In_1819);
and U438 (N_438,In_1076,In_542);
nor U439 (N_439,In_299,In_1350);
or U440 (N_440,In_1344,In_354);
or U441 (N_441,In_592,In_2455);
nor U442 (N_442,In_2508,In_1200);
and U443 (N_443,In_765,In_361);
nand U444 (N_444,In_1587,In_297);
or U445 (N_445,In_1474,In_1468);
and U446 (N_446,In_2059,In_1947);
nand U447 (N_447,In_2428,In_795);
xor U448 (N_448,In_330,In_967);
or U449 (N_449,In_1230,In_1025);
xnor U450 (N_450,In_2940,In_1618);
xor U451 (N_451,In_2154,In_2034);
xor U452 (N_452,In_2846,In_2539);
nand U453 (N_453,In_1749,In_2427);
and U454 (N_454,In_2465,In_870);
xor U455 (N_455,In_1918,In_2930);
xor U456 (N_456,In_339,In_589);
or U457 (N_457,In_2977,In_2528);
xor U458 (N_458,In_1495,In_418);
nand U459 (N_459,In_1310,In_842);
or U460 (N_460,In_2972,In_2880);
and U461 (N_461,In_2092,In_914);
nand U462 (N_462,In_506,In_27);
nand U463 (N_463,In_1507,In_2847);
nor U464 (N_464,In_1026,In_1326);
and U465 (N_465,In_1137,In_2525);
xnor U466 (N_466,In_2073,In_2456);
nor U467 (N_467,In_757,In_551);
nor U468 (N_468,In_322,In_2810);
nand U469 (N_469,In_351,In_1825);
and U470 (N_470,In_178,In_252);
xor U471 (N_471,In_1845,In_2881);
nand U472 (N_472,In_657,In_1914);
nand U473 (N_473,In_1187,In_2926);
nand U474 (N_474,In_1926,In_2569);
nor U475 (N_475,In_2550,In_739);
nor U476 (N_476,In_2969,In_1109);
nand U477 (N_477,In_1390,In_119);
or U478 (N_478,In_1560,In_1794);
or U479 (N_479,In_2234,In_2353);
and U480 (N_480,In_2656,In_1366);
nand U481 (N_481,In_1235,In_2204);
or U482 (N_482,In_2910,In_1038);
nand U483 (N_483,In_1217,In_1985);
nor U484 (N_484,In_2832,In_2960);
xnor U485 (N_485,In_187,In_2878);
nor U486 (N_486,In_2405,In_1463);
xor U487 (N_487,In_1758,In_133);
nor U488 (N_488,In_1872,In_1251);
xnor U489 (N_489,In_2700,In_1117);
nand U490 (N_490,In_2871,In_495);
nand U491 (N_491,In_2040,In_2363);
and U492 (N_492,In_1048,In_1078);
and U493 (N_493,In_556,In_2484);
or U494 (N_494,In_931,In_1799);
xnor U495 (N_495,In_1954,In_1673);
and U496 (N_496,In_268,In_2491);
or U497 (N_497,In_590,In_1100);
nand U498 (N_498,In_242,In_48);
and U499 (N_499,In_7,In_454);
and U500 (N_500,In_1744,In_709);
nor U501 (N_501,In_1801,In_2397);
nand U502 (N_502,In_1766,In_820);
or U503 (N_503,In_2261,In_1252);
xor U504 (N_504,In_2184,In_2617);
nor U505 (N_505,In_2626,In_1343);
nor U506 (N_506,In_766,In_2678);
and U507 (N_507,In_996,In_1963);
nand U508 (N_508,In_503,In_2520);
xnor U509 (N_509,In_111,In_510);
nand U510 (N_510,In_1391,In_2911);
nor U511 (N_511,In_2454,In_777);
and U512 (N_512,In_694,In_355);
nand U513 (N_513,In_1207,In_1736);
xor U514 (N_514,In_2207,In_1281);
and U515 (N_515,In_2481,In_1211);
nand U516 (N_516,In_2645,In_2627);
and U517 (N_517,In_2156,In_1365);
nand U518 (N_518,In_1445,In_385);
nand U519 (N_519,In_20,In_2736);
nand U520 (N_520,In_2664,In_2927);
and U521 (N_521,In_1632,In_2464);
xnor U522 (N_522,In_338,In_2037);
xor U523 (N_523,In_1185,In_1804);
or U524 (N_524,In_1363,In_366);
xor U525 (N_525,In_1591,In_937);
and U526 (N_526,In_2851,In_2131);
nor U527 (N_527,In_578,In_2262);
nand U528 (N_528,In_0,In_653);
nand U529 (N_529,In_2494,In_374);
nand U530 (N_530,In_2600,In_1003);
nor U531 (N_531,In_2292,In_1654);
and U532 (N_532,In_1429,In_168);
and U533 (N_533,In_2855,In_583);
nand U534 (N_534,In_1553,In_480);
nand U535 (N_535,In_1748,In_2875);
xnor U536 (N_536,In_1860,In_1107);
nand U537 (N_537,In_853,In_1663);
nand U538 (N_538,In_1773,In_2483);
or U539 (N_539,In_212,In_2717);
or U540 (N_540,In_2610,In_2316);
xnor U541 (N_541,In_686,In_1082);
nand U542 (N_542,In_478,In_1120);
or U543 (N_543,In_2570,In_1815);
and U544 (N_544,In_721,In_2702);
or U545 (N_545,In_1389,In_60);
nor U546 (N_546,In_2874,In_1599);
nor U547 (N_547,In_1172,In_962);
xnor U548 (N_548,In_2196,In_2452);
and U549 (N_549,In_1133,In_84);
and U550 (N_550,In_516,In_1525);
nor U551 (N_551,In_2945,In_2060);
xor U552 (N_552,In_2064,In_1104);
nor U553 (N_553,In_1030,In_200);
or U554 (N_554,In_1075,In_2791);
or U555 (N_555,In_1451,In_2538);
or U556 (N_556,In_59,In_735);
nor U557 (N_557,In_920,In_1846);
nand U558 (N_558,In_1607,In_1462);
nor U559 (N_559,In_171,In_16);
nor U560 (N_560,In_2637,In_810);
xor U561 (N_561,In_2245,In_736);
nor U562 (N_562,In_2492,In_1750);
or U563 (N_563,In_2354,In_1576);
or U564 (N_564,In_2647,In_2956);
xnor U565 (N_565,In_1817,In_783);
and U566 (N_566,In_802,In_2311);
xor U567 (N_567,In_682,In_2209);
xnor U568 (N_568,In_695,In_1837);
nor U569 (N_569,In_1575,In_559);
nor U570 (N_570,In_1214,In_1022);
nand U571 (N_571,In_2725,In_307);
or U572 (N_572,In_733,In_975);
nor U573 (N_573,In_778,In_1589);
or U574 (N_574,In_292,In_342);
and U575 (N_575,In_138,In_1696);
and U576 (N_576,In_1295,In_1644);
nand U577 (N_577,In_822,In_2719);
nand U578 (N_578,In_2589,In_543);
and U579 (N_579,In_395,In_1510);
nor U580 (N_580,In_1260,In_635);
nand U581 (N_581,In_2607,In_705);
xnor U582 (N_582,In_2658,In_1812);
nor U583 (N_583,In_2007,In_420);
xor U584 (N_584,In_880,In_130);
nand U585 (N_585,In_352,In_1636);
nor U586 (N_586,In_2757,In_482);
or U587 (N_587,In_1411,In_343);
nor U588 (N_588,In_372,In_306);
nand U589 (N_589,In_889,In_1062);
or U590 (N_590,In_1604,In_1456);
and U591 (N_591,In_913,In_93);
or U592 (N_592,In_2574,In_605);
or U593 (N_593,In_139,In_2247);
and U594 (N_594,In_2813,In_2795);
or U595 (N_595,In_611,In_2332);
nand U596 (N_596,In_553,In_4);
or U597 (N_597,In_1980,In_2923);
or U598 (N_598,In_1543,In_2936);
and U599 (N_599,In_473,In_2438);
and U600 (N_600,In_1544,In_647);
and U601 (N_601,In_1823,In_1033);
or U602 (N_602,In_95,In_1015);
and U603 (N_603,In_841,In_1558);
or U604 (N_604,In_1661,In_1020);
xor U605 (N_605,In_1671,In_546);
nand U606 (N_606,In_1511,In_1232);
or U607 (N_607,In_2777,In_1657);
or U608 (N_608,In_743,In_2737);
nand U609 (N_609,In_2564,In_2212);
xor U610 (N_610,In_1315,In_2763);
xnor U611 (N_611,In_2143,In_1127);
xnor U612 (N_612,In_1303,In_2720);
xnor U613 (N_613,In_1726,In_2982);
or U614 (N_614,In_1844,In_1225);
nand U615 (N_615,In_2019,In_2242);
and U616 (N_616,In_970,In_1668);
xnor U617 (N_617,In_2723,In_725);
xnor U618 (N_618,In_2244,In_1957);
xnor U619 (N_619,In_126,In_1828);
or U620 (N_620,In_1010,In_729);
and U621 (N_621,In_1037,In_1583);
or U622 (N_622,In_2852,In_2544);
nor U623 (N_623,In_753,In_2430);
and U624 (N_624,In_334,In_127);
and U625 (N_625,In_895,In_2451);
and U626 (N_626,In_1551,In_2938);
and U627 (N_627,In_839,In_1904);
and U628 (N_628,In_1574,In_441);
xnor U629 (N_629,In_1877,In_186);
nor U630 (N_630,In_540,In_2374);
nor U631 (N_631,In_665,In_2029);
nor U632 (N_632,In_2686,In_2897);
nand U633 (N_633,In_526,In_2955);
nor U634 (N_634,In_2705,In_1046);
and U635 (N_635,In_823,In_2031);
and U636 (N_636,In_1072,In_1586);
xor U637 (N_637,In_269,In_142);
or U638 (N_638,In_55,In_267);
or U639 (N_639,In_2011,In_1134);
xor U640 (N_640,In_2914,In_1515);
nand U641 (N_641,In_2334,In_770);
or U642 (N_642,In_145,In_2684);
xor U643 (N_643,In_1849,In_1464);
nor U644 (N_644,In_793,In_2150);
xnor U645 (N_645,In_1203,In_386);
nand U646 (N_646,In_56,In_676);
or U647 (N_647,In_779,In_132);
and U648 (N_648,In_2395,In_2033);
nand U649 (N_649,In_861,In_1221);
nor U650 (N_650,In_1198,In_2707);
and U651 (N_651,In_2410,In_670);
xnor U652 (N_652,In_2764,In_999);
or U653 (N_653,In_29,In_1094);
or U654 (N_654,In_2229,In_2839);
nor U655 (N_655,In_2050,In_2931);
xor U656 (N_656,In_1912,In_2259);
nand U657 (N_657,In_2170,In_2160);
and U658 (N_658,In_561,In_1324);
nand U659 (N_659,In_254,In_2790);
or U660 (N_660,In_2794,In_1340);
xor U661 (N_661,In_1724,In_2277);
xnor U662 (N_662,In_2925,In_2444);
nor U663 (N_663,In_2742,In_816);
nand U664 (N_664,In_1713,In_639);
nor U665 (N_665,In_2407,In_2780);
nor U666 (N_666,In_1633,In_677);
and U667 (N_667,In_1119,In_317);
and U668 (N_668,In_1276,In_1250);
nor U669 (N_669,In_143,In_1457);
xor U670 (N_670,In_1716,In_1746);
nand U671 (N_671,In_2849,In_744);
nor U672 (N_672,In_2053,In_2227);
and U673 (N_673,In_2924,In_1279);
xnor U674 (N_674,In_1561,In_2826);
xnor U675 (N_675,In_1711,In_831);
xnor U676 (N_676,In_284,In_1529);
or U677 (N_677,In_15,In_675);
nand U678 (N_678,In_2102,In_900);
nor U679 (N_679,In_645,In_2903);
or U680 (N_680,In_2282,In_1878);
or U681 (N_681,In_453,In_2258);
nand U682 (N_682,In_465,In_934);
or U683 (N_683,In_1687,In_2146);
and U684 (N_684,In_549,In_1443);
xor U685 (N_685,In_505,In_1419);
nor U686 (N_686,In_1332,In_249);
nor U687 (N_687,In_1360,In_1754);
and U688 (N_688,In_2530,In_1779);
nor U689 (N_689,In_2000,In_854);
or U690 (N_690,In_57,In_2433);
nor U691 (N_691,In_1115,In_2035);
xor U692 (N_692,In_1055,In_2191);
and U693 (N_693,In_1781,In_923);
nor U694 (N_694,In_2414,In_1516);
nand U695 (N_695,In_2727,In_1643);
nand U696 (N_696,In_2422,In_2152);
nor U697 (N_697,In_150,In_2224);
nand U698 (N_698,In_2401,In_227);
or U699 (N_699,In_847,In_2630);
and U700 (N_700,In_2248,In_1421);
nor U701 (N_701,In_2819,In_1347);
or U702 (N_702,In_2243,In_2488);
nand U703 (N_703,In_603,In_1147);
xor U704 (N_704,In_1261,In_2087);
and U705 (N_705,In_642,In_1908);
nand U706 (N_706,In_173,In_2302);
xnor U707 (N_707,In_255,In_312);
xnor U708 (N_708,In_979,In_2909);
nor U709 (N_709,In_104,In_1005);
or U710 (N_710,In_2778,In_2280);
and U711 (N_711,In_580,In_135);
nand U712 (N_712,In_1564,In_2816);
xor U713 (N_713,In_1194,In_1956);
and U714 (N_714,In_160,In_720);
or U715 (N_715,In_604,In_416);
nor U716 (N_716,In_852,In_1697);
xor U717 (N_717,In_253,In_830);
or U718 (N_718,In_2716,In_2842);
xnor U719 (N_719,In_2643,In_2125);
nor U720 (N_720,In_315,In_2500);
xor U721 (N_721,In_953,In_464);
and U722 (N_722,In_930,In_1158);
or U723 (N_723,In_1798,In_117);
and U724 (N_724,In_1169,In_1641);
or U725 (N_725,In_2083,In_34);
nand U726 (N_726,In_182,In_422);
nand U727 (N_727,In_2164,In_2116);
nor U728 (N_728,In_2756,In_2376);
nand U729 (N_729,In_2335,In_2378);
xor U730 (N_730,In_2274,In_2106);
nand U731 (N_731,In_1380,In_1705);
nor U732 (N_732,In_463,In_713);
nand U733 (N_733,In_485,In_1245);
and U734 (N_734,In_1563,In_2590);
and U735 (N_735,In_2613,In_2683);
nand U736 (N_736,In_2567,In_1873);
nand U737 (N_737,In_291,In_2860);
nor U738 (N_738,In_174,In_1925);
and U739 (N_739,In_807,In_1991);
nand U740 (N_740,In_1297,In_2495);
or U741 (N_741,In_907,In_1616);
nand U742 (N_742,In_2840,In_1387);
nor U743 (N_743,In_2272,In_1027);
xor U744 (N_744,In_597,In_265);
nor U745 (N_745,In_1047,In_1275);
xor U746 (N_746,In_2326,In_2273);
and U747 (N_747,In_879,In_1609);
xor U748 (N_748,In_1852,In_2421);
or U749 (N_749,In_42,In_1149);
nor U750 (N_750,In_613,In_2663);
nand U751 (N_751,In_122,In_2640);
xor U752 (N_752,In_882,In_1067);
nor U753 (N_753,In_1530,In_202);
xor U754 (N_754,In_314,In_1167);
nand U755 (N_755,In_2890,In_1196);
nand U756 (N_756,In_2802,In_992);
nand U757 (N_757,In_2028,In_763);
xor U758 (N_758,In_2216,In_562);
and U759 (N_759,In_2496,In_2682);
and U760 (N_760,In_1388,In_1603);
nand U761 (N_761,In_1871,In_2281);
and U762 (N_762,In_804,In_2253);
xnor U763 (N_763,In_2015,In_809);
and U764 (N_764,In_49,In_1335);
or U765 (N_765,In_2797,In_508);
and U766 (N_766,In_22,In_1296);
xor U767 (N_767,In_251,In_2369);
or U768 (N_768,In_2030,In_749);
and U769 (N_769,In_1674,In_290);
xor U770 (N_770,In_116,In_1688);
nor U771 (N_771,In_1907,In_1348);
xor U772 (N_772,In_2591,In_2554);
xor U773 (N_773,In_759,In_2149);
xnor U774 (N_774,In_2830,In_1195);
nor U775 (N_775,In_598,In_2559);
nor U776 (N_776,In_828,In_2251);
nor U777 (N_777,In_239,In_375);
or U778 (N_778,In_1000,In_1639);
nand U779 (N_779,In_2231,In_2069);
xor U780 (N_780,In_2505,In_1053);
or U781 (N_781,In_764,In_2446);
xor U782 (N_782,In_2691,In_398);
nand U783 (N_783,In_2655,In_2386);
or U784 (N_784,In_614,In_2829);
xor U785 (N_785,In_2984,In_2838);
and U786 (N_786,In_1486,In_1492);
or U787 (N_787,In_2226,In_618);
xnor U788 (N_788,In_2396,In_303);
and U789 (N_789,In_1213,In_1789);
nand U790 (N_790,In_2114,In_332);
nor U791 (N_791,In_1428,In_1722);
nor U792 (N_792,In_897,In_1578);
and U793 (N_793,In_581,In_474);
xor U794 (N_794,In_2950,In_1384);
or U795 (N_795,In_1961,In_2767);
nor U796 (N_796,In_1547,In_1620);
or U797 (N_797,In_458,In_1417);
nor U798 (N_798,In_2512,In_2817);
nor U799 (N_799,In_815,In_426);
nor U800 (N_800,In_946,In_2864);
and U801 (N_801,In_711,In_1703);
or U802 (N_802,In_311,In_1660);
xor U803 (N_803,In_229,In_698);
nand U804 (N_804,In_2809,In_565);
nand U805 (N_805,In_2879,In_2835);
nor U806 (N_806,In_771,In_425);
xnor U807 (N_807,In_1454,In_1093);
or U808 (N_808,In_490,In_1863);
xnor U809 (N_809,In_1448,In_2218);
nor U810 (N_810,In_641,In_2556);
and U811 (N_811,In_2241,In_2629);
nor U812 (N_812,In_2870,In_1359);
xnor U813 (N_813,In_2279,In_1838);
or U814 (N_814,In_308,In_1489);
xnor U815 (N_815,In_2176,In_983);
nand U816 (N_816,In_2662,In_2557);
xnor U817 (N_817,In_2476,In_1496);
xnor U818 (N_818,In_1369,In_2358);
nor U819 (N_819,In_1699,In_1967);
nor U820 (N_820,In_345,In_1857);
or U821 (N_821,In_2621,In_2493);
and U822 (N_822,In_2325,In_792);
nand U823 (N_823,In_2948,In_1145);
or U824 (N_824,In_2765,In_984);
nor U825 (N_825,In_750,In_9);
or U826 (N_826,In_1987,In_1651);
nand U827 (N_827,In_1191,In_1774);
or U828 (N_828,In_469,In_519);
and U829 (N_829,In_2585,In_1929);
nor U830 (N_830,In_107,In_156);
and U831 (N_831,In_248,In_1708);
and U832 (N_832,In_1188,In_643);
nor U833 (N_833,In_2843,In_2167);
or U834 (N_834,In_243,In_2804);
nor U835 (N_835,In_745,In_656);
or U836 (N_836,In_833,In_68);
and U837 (N_837,In_2713,In_335);
or U838 (N_838,In_1706,In_228);
nor U839 (N_839,In_954,In_1897);
and U840 (N_840,In_2474,In_524);
nor U841 (N_841,In_1114,In_569);
nor U842 (N_842,In_1698,In_2324);
xnor U843 (N_843,In_1135,In_2301);
nor U844 (N_844,In_730,In_224);
nor U845 (N_845,In_2666,In_538);
nor U846 (N_846,In_2548,In_902);
nor U847 (N_847,In_1762,In_579);
nor U848 (N_848,In_37,In_2689);
nand U849 (N_849,In_1839,In_1627);
xnor U850 (N_850,In_1854,In_929);
or U851 (N_851,In_1642,In_1596);
and U852 (N_852,In_1790,In_1274);
xnor U853 (N_853,In_197,In_1645);
nor U854 (N_854,In_2435,In_2687);
or U855 (N_855,In_1223,In_436);
and U856 (N_856,In_348,In_588);
xor U857 (N_857,In_2237,In_531);
or U858 (N_858,In_1621,In_18);
or U859 (N_859,In_2437,In_1568);
nand U860 (N_860,In_2677,In_1927);
nand U861 (N_861,In_402,In_1807);
nand U862 (N_862,In_626,In_876);
or U863 (N_863,In_2785,In_2356);
or U864 (N_864,In_1890,In_1314);
and U865 (N_865,In_2021,In_696);
or U866 (N_866,In_443,In_1938);
nor U867 (N_867,In_2993,In_788);
xor U868 (N_868,In_190,In_362);
or U869 (N_869,In_92,In_110);
nor U870 (N_870,In_916,In_2623);
nand U871 (N_871,In_932,In_36);
nand U872 (N_872,In_1753,In_177);
nand U873 (N_873,In_393,In_1301);
nand U874 (N_874,In_483,In_886);
nand U875 (N_875,In_591,In_411);
or U876 (N_876,In_1735,In_2962);
xor U877 (N_877,In_1485,In_2704);
nand U878 (N_878,In_2365,In_1629);
or U879 (N_879,In_61,In_1859);
or U880 (N_880,In_86,In_714);
or U881 (N_881,In_1061,In_2774);
or U882 (N_882,In_952,In_2088);
and U883 (N_883,In_935,In_2971);
xor U884 (N_884,In_1880,In_1870);
and U885 (N_885,In_1124,In_496);
nand U886 (N_886,In_146,In_1741);
or U887 (N_887,In_2601,In_2555);
nor U888 (N_888,In_2220,In_2470);
nor U889 (N_889,In_977,In_450);
nor U890 (N_890,In_2418,In_112);
nor U891 (N_891,In_2714,In_1377);
or U892 (N_892,In_1184,In_1997);
xnor U893 (N_893,In_2425,In_288);
nand U894 (N_894,In_922,In_2848);
or U895 (N_895,In_2254,In_1780);
or U896 (N_896,In_2290,In_968);
xor U897 (N_897,In_2822,In_2786);
and U898 (N_898,In_134,In_1313);
and U899 (N_899,In_874,In_2893);
nand U900 (N_900,In_1283,In_1299);
and U901 (N_901,In_316,In_2921);
nor U902 (N_902,In_1086,In_938);
nand U903 (N_903,In_497,In_2747);
nand U904 (N_904,In_2792,In_283);
xnor U905 (N_905,In_1803,In_462);
and U906 (N_906,In_888,In_1021);
nand U907 (N_907,In_1555,In_1406);
xnor U908 (N_908,In_892,In_1867);
nand U909 (N_909,In_2503,In_340);
nor U910 (N_910,In_2331,In_944);
xor U911 (N_911,In_1426,In_2291);
nand U912 (N_912,In_498,In_2429);
nor U913 (N_913,In_5,In_1982);
nand U914 (N_914,In_2768,In_738);
nand U915 (N_915,In_1652,In_2315);
nor U916 (N_916,In_2660,In_2718);
nor U917 (N_917,In_2928,In_2039);
nor U918 (N_918,In_2831,In_905);
and U919 (N_919,In_2384,In_1869);
xor U920 (N_920,In_2772,In_1770);
and U921 (N_921,In_2104,In_1157);
and U922 (N_922,In_2478,In_2730);
nand U923 (N_923,In_364,In_2442);
xor U924 (N_924,In_717,In_2303);
or U925 (N_925,In_2111,In_2349);
and U926 (N_926,In_2762,In_2265);
xor U927 (N_927,In_1193,In_1602);
nand U928 (N_928,In_1995,In_2828);
or U929 (N_929,In_2112,In_1573);
and U930 (N_930,In_2085,In_1293);
nor U931 (N_931,In_2949,In_646);
nor U932 (N_932,In_1423,In_2065);
nand U933 (N_933,In_791,In_2696);
nor U934 (N_934,In_24,In_1695);
or U935 (N_935,In_2352,In_2536);
and U936 (N_936,In_2625,In_226);
xnor U937 (N_937,In_906,In_103);
and U938 (N_938,In_2096,In_1521);
and U939 (N_939,In_1018,In_575);
or U940 (N_940,In_557,In_1532);
or U941 (N_941,In_2605,In_2382);
xor U942 (N_942,In_262,In_836);
xor U943 (N_943,In_1895,In_1984);
nand U944 (N_944,In_2081,In_1334);
nand U945 (N_945,In_166,In_1019);
and U946 (N_946,In_2027,In_1752);
or U947 (N_947,In_1742,In_634);
xnor U948 (N_948,In_2854,In_278);
and U949 (N_949,In_21,In_47);
nor U950 (N_950,In_2056,In_666);
nor U951 (N_951,In_1730,In_172);
nand U952 (N_952,In_1950,In_1028);
nand U953 (N_953,In_2857,In_2734);
and U954 (N_954,In_1467,In_2518);
or U955 (N_955,In_2514,In_2394);
nand U956 (N_956,In_1099,In_1269);
nand U957 (N_957,In_2604,In_371);
nor U958 (N_958,In_544,In_1065);
or U959 (N_959,In_2729,In_2542);
nand U960 (N_960,In_2199,In_220);
xor U961 (N_961,In_2999,In_688);
or U962 (N_962,In_2741,In_1447);
nand U963 (N_963,In_457,In_548);
nand U964 (N_964,In_1397,In_2145);
xor U965 (N_965,In_2284,In_1355);
and U966 (N_966,In_1556,In_2482);
and U967 (N_967,In_621,In_500);
and U968 (N_968,In_83,In_624);
nand U969 (N_969,In_2233,In_567);
or U970 (N_970,In_619,In_2119);
and U971 (N_971,In_1612,In_2781);
and U972 (N_972,In_233,In_1884);
and U973 (N_973,In_1677,In_437);
and U974 (N_974,In_1330,In_1958);
nand U975 (N_975,In_1247,In_1273);
xnor U976 (N_976,In_702,In_2411);
and U977 (N_977,In_369,In_1631);
nor U978 (N_978,In_1795,In_1945);
nor U979 (N_979,In_1159,In_75);
xnor U980 (N_980,In_2091,In_141);
nand U981 (N_981,In_2042,In_333);
nand U982 (N_982,In_2552,In_2135);
and U983 (N_983,In_2983,In_167);
xor U984 (N_984,In_2980,In_2256);
and U985 (N_985,In_1268,In_2193);
nor U986 (N_986,In_2453,In_488);
and U987 (N_987,In_1241,In_1909);
or U988 (N_988,In_2210,In_2579);
nand U989 (N_989,In_2120,In_2079);
nand U990 (N_990,In_2439,In_2889);
nand U991 (N_991,In_2951,In_1528);
nor U992 (N_992,In_2912,In_959);
or U993 (N_993,In_1413,In_286);
nor U994 (N_994,In_30,In_78);
or U995 (N_995,In_1595,In_1069);
xnor U996 (N_996,In_982,In_1148);
xnor U997 (N_997,In_884,In_2532);
nand U998 (N_998,In_2366,In_1438);
nor U999 (N_999,In_1715,In_2891);
and U1000 (N_1000,In_801,In_2434);
and U1001 (N_1001,In_1747,In_2636);
or U1002 (N_1002,In_1590,In_231);
nor U1003 (N_1003,In_28,In_419);
and U1004 (N_1004,In_2413,In_2633);
or U1005 (N_1005,In_1288,In_2899);
nand U1006 (N_1006,In_2134,In_1071);
or U1007 (N_1007,In_1132,In_2771);
nor U1008 (N_1008,In_2486,In_1557);
xor U1009 (N_1009,In_2551,In_216);
nand U1010 (N_1010,In_2080,In_585);
xnor U1011 (N_1011,In_1444,In_2888);
and U1012 (N_1012,In_623,In_878);
xor U1013 (N_1013,In_593,In_969);
nor U1014 (N_1014,In_887,In_1519);
xor U1015 (N_1015,In_207,In_2776);
and U1016 (N_1016,In_2318,In_179);
nor U1017 (N_1017,In_2966,In_2932);
nor U1018 (N_1018,In_310,In_1992);
xnor U1019 (N_1019,In_1393,In_397);
nor U1020 (N_1020,In_2260,In_91);
xnor U1021 (N_1021,In_96,In_1969);
or U1022 (N_1022,In_767,In_1548);
or U1023 (N_1023,In_1017,In_2726);
or U1024 (N_1024,In_14,In_981);
nor U1025 (N_1025,In_723,In_1146);
xor U1026 (N_1026,In_1222,In_1876);
nand U1027 (N_1027,In_2598,In_1204);
nor U1028 (N_1028,In_2581,In_2406);
nand U1029 (N_1029,In_1242,In_850);
nand U1030 (N_1030,In_1538,In_12);
or U1031 (N_1031,In_2856,In_2342);
and U1032 (N_1032,In_570,In_1719);
nand U1033 (N_1033,In_1289,In_1080);
xor U1034 (N_1034,In_1403,In_401);
xor U1035 (N_1035,In_2612,In_353);
nor U1036 (N_1036,In_2868,In_664);
nand U1037 (N_1037,In_2609,In_599);
nand U1038 (N_1038,In_1787,In_183);
nor U1039 (N_1039,In_2390,In_1378);
nor U1040 (N_1040,In_918,In_708);
or U1041 (N_1041,In_2173,In_2905);
nand U1042 (N_1042,In_1843,In_2575);
nor U1043 (N_1043,In_2947,In_2515);
xnor U1044 (N_1044,In_2759,In_1554);
nor U1045 (N_1045,In_2906,In_2377);
nand U1046 (N_1046,In_2793,In_2976);
and U1047 (N_1047,In_1190,In_911);
nand U1048 (N_1048,In_1729,In_1179);
nand U1049 (N_1049,In_1605,In_615);
or U1050 (N_1050,In_2457,In_1455);
nand U1051 (N_1051,In_576,In_2264);
xnor U1052 (N_1052,In_1865,In_2041);
and U1053 (N_1053,In_896,In_1720);
nand U1054 (N_1054,In_1723,In_2312);
and U1055 (N_1055,In_2898,In_198);
nor U1056 (N_1056,In_2328,In_2534);
and U1057 (N_1057,In_1952,In_2339);
or U1058 (N_1058,In_2161,In_1256);
xnor U1059 (N_1059,In_1434,In_890);
and U1060 (N_1060,In_1505,In_1239);
xnor U1061 (N_1061,In_19,In_2461);
xnor U1062 (N_1062,In_492,In_697);
nand U1063 (N_1063,In_435,In_1008);
or U1064 (N_1064,In_1562,In_1199);
and U1065 (N_1065,In_321,In_211);
and U1066 (N_1066,In_1458,In_1680);
and U1067 (N_1067,In_2743,In_2679);
and U1068 (N_1068,In_1308,In_1358);
and U1069 (N_1069,In_428,In_2758);
or U1070 (N_1070,In_616,In_1404);
or U1071 (N_1071,In_1579,In_2739);
or U1072 (N_1072,In_245,In_1170);
nand U1073 (N_1073,In_1291,In_1437);
or U1074 (N_1074,In_1081,In_470);
nand U1075 (N_1075,In_2294,In_2205);
nand U1076 (N_1076,In_1656,In_814);
nand U1077 (N_1077,In_391,In_2137);
xor U1078 (N_1078,In_1990,In_1041);
nor U1079 (N_1079,In_2235,In_2132);
nor U1080 (N_1080,In_399,In_1778);
xnor U1081 (N_1081,In_2296,In_747);
nor U1082 (N_1082,In_2620,In_1307);
nor U1083 (N_1083,In_1376,In_1565);
nand U1084 (N_1084,In_1142,In_512);
xnor U1085 (N_1085,In_2448,In_2148);
or U1086 (N_1086,In_1001,In_147);
xor U1087 (N_1087,In_235,In_1278);
xor U1088 (N_1088,In_1965,In_1771);
nand U1089 (N_1089,In_1151,In_1690);
xnor U1090 (N_1090,In_2509,In_844);
and U1091 (N_1091,In_2350,In_1058);
xor U1092 (N_1092,In_2006,In_276);
nor U1093 (N_1093,In_2348,In_574);
or U1094 (N_1094,In_1883,In_347);
nor U1095 (N_1095,In_1024,In_785);
and U1096 (N_1096,In_2487,In_195);
or U1097 (N_1097,In_2100,In_2155);
nor U1098 (N_1098,In_88,In_857);
xnor U1099 (N_1099,In_1536,In_659);
nor U1100 (N_1100,In_148,In_2907);
xor U1101 (N_1101,In_680,In_357);
xnor U1102 (N_1102,In_2044,In_2129);
nand U1103 (N_1103,In_2278,In_486);
nand U1104 (N_1104,In_2489,In_535);
xor U1105 (N_1105,In_2498,In_2614);
xor U1106 (N_1106,In_2002,In_471);
xnor U1107 (N_1107,In_2467,In_2240);
nor U1108 (N_1108,In_924,In_1029);
nand U1109 (N_1109,In_328,In_1955);
and U1110 (N_1110,In_2054,In_774);
nand U1111 (N_1111,In_885,In_2996);
or U1112 (N_1112,In_170,In_2943);
xor U1113 (N_1113,In_407,In_541);
and U1114 (N_1114,In_2648,In_2584);
nand U1115 (N_1115,In_32,In_2850);
and U1116 (N_1116,In_1793,In_1282);
and U1117 (N_1117,In_1776,In_758);
and U1118 (N_1118,In_69,In_863);
nor U1119 (N_1119,In_1271,In_2472);
nor U1120 (N_1120,In_2853,In_928);
xnor U1121 (N_1121,In_370,In_545);
xnor U1122 (N_1122,In_2285,In_608);
or U1123 (N_1123,In_1717,In_1435);
and U1124 (N_1124,In_2424,In_2157);
xnor U1125 (N_1125,In_501,In_2440);
and U1126 (N_1126,In_655,In_1229);
xor U1127 (N_1127,In_1054,In_1471);
nor U1128 (N_1128,In_1597,In_2426);
xor U1129 (N_1129,In_974,In_972);
nor U1130 (N_1130,In_282,In_1930);
and U1131 (N_1131,In_1163,In_2463);
and U1132 (N_1132,In_70,In_2);
nand U1133 (N_1133,In_812,In_689);
and U1134 (N_1134,In_1056,In_236);
or U1135 (N_1135,In_868,In_1624);
nand U1136 (N_1136,In_582,In_573);
xnor U1137 (N_1137,In_430,In_2249);
nand U1138 (N_1138,In_2524,In_2385);
nand U1139 (N_1139,In_379,In_1394);
xor U1140 (N_1140,In_1012,In_1864);
xor U1141 (N_1141,In_410,In_455);
and U1142 (N_1142,In_8,In_834);
or U1143 (N_1143,In_1092,In_438);
and U1144 (N_1144,In_1821,In_2502);
nor U1145 (N_1145,In_989,In_668);
or U1146 (N_1146,In_2884,In_1585);
xnor U1147 (N_1147,In_1300,In_2344);
or U1148 (N_1148,In_77,In_2833);
xnor U1149 (N_1149,In_1465,In_324);
or U1150 (N_1150,In_105,In_2018);
nand U1151 (N_1151,In_1409,In_692);
nor U1152 (N_1152,In_2571,In_2130);
or U1153 (N_1153,In_1083,In_240);
or U1154 (N_1154,In_206,In_1901);
and U1155 (N_1155,In_835,In_336);
nor U1156 (N_1156,In_2159,In_2744);
and U1157 (N_1157,In_797,In_1488);
nand U1158 (N_1158,In_1685,In_1503);
or U1159 (N_1159,In_359,In_803);
nand U1160 (N_1160,In_1649,In_2409);
nor U1161 (N_1161,In_1648,In_712);
or U1162 (N_1162,In_1976,In_1740);
xor U1163 (N_1163,In_1517,In_1567);
nor U1164 (N_1164,In_368,In_2183);
or U1165 (N_1165,In_1732,In_1772);
xor U1166 (N_1166,In_1470,In_2182);
or U1167 (N_1167,In_2117,In_998);
xor U1168 (N_1168,In_1847,In_2398);
nand U1169 (N_1169,In_555,In_2746);
or U1170 (N_1170,In_507,In_1903);
nand U1171 (N_1171,In_2800,In_1808);
and U1172 (N_1172,In_1098,In_1118);
and U1173 (N_1173,In_1280,In_2017);
and U1174 (N_1174,In_2504,In_2712);
xor U1175 (N_1175,In_1504,In_309);
and U1176 (N_1176,In_2228,In_1514);
or U1177 (N_1177,In_158,In_1441);
nand U1178 (N_1178,In_971,In_908);
and U1179 (N_1179,In_2531,In_2321);
and U1180 (N_1180,In_376,In_1006);
or U1181 (N_1181,In_2293,In_2632);
nand U1182 (N_1182,In_1031,In_1848);
and U1183 (N_1183,In_973,In_1091);
nor U1184 (N_1184,In_1853,In_1243);
and U1185 (N_1185,In_1272,In_123);
xnor U1186 (N_1186,In_10,In_382);
nand U1187 (N_1187,In_1306,In_2770);
nor U1188 (N_1188,In_1088,In_2340);
and U1189 (N_1189,In_1634,In_204);
or U1190 (N_1190,In_2920,In_2076);
and U1191 (N_1191,In_2887,In_1329);
xor U1192 (N_1192,In_943,In_2250);
nor U1193 (N_1193,In_304,In_1227);
nand U1194 (N_1194,In_966,In_1721);
nor U1195 (N_1195,In_432,In_2933);
nor U1196 (N_1196,In_346,In_1262);
nand U1197 (N_1197,In_2490,In_1292);
xor U1198 (N_1198,In_2904,In_537);
or U1199 (N_1199,In_2665,In_2151);
nor U1200 (N_1200,In_1180,In_1714);
xor U1201 (N_1201,In_875,In_2761);
or U1202 (N_1202,In_1304,In_1637);
or U1203 (N_1203,In_1226,In_2283);
xor U1204 (N_1204,In_1089,In_1905);
and U1205 (N_1205,In_1036,In_1112);
and U1206 (N_1206,In_2391,In_1459);
nor U1207 (N_1207,In_1349,In_1694);
nor U1208 (N_1208,In_2417,In_2219);
nor U1209 (N_1209,In_2877,In_390);
xnor U1210 (N_1210,In_50,In_2305);
xor U1211 (N_1211,In_99,In_530);
xnor U1212 (N_1212,In_560,In_2010);
xor U1213 (N_1213,In_1183,In_1052);
nor U1214 (N_1214,In_845,In_1640);
nand U1215 (N_1215,In_1856,In_1763);
nand U1216 (N_1216,In_2351,In_715);
or U1217 (N_1217,In_1850,In_1800);
xor U1218 (N_1218,In_775,In_2900);
nand U1219 (N_1219,In_699,In_2068);
nor U1220 (N_1220,In_2392,In_350);
nor U1221 (N_1221,In_400,In_1923);
xor U1222 (N_1222,In_617,In_2008);
xor U1223 (N_1223,In_2701,In_961);
nand U1224 (N_1224,In_669,In_1831);
nand U1225 (N_1225,In_991,In_719);
or U1226 (N_1226,In_261,In_2165);
nor U1227 (N_1227,In_1830,In_1405);
nor U1228 (N_1228,In_2238,In_1136);
nand U1229 (N_1229,In_2654,In_960);
nor U1230 (N_1230,In_221,In_234);
xnor U1231 (N_1231,In_644,In_2616);
nand U1232 (N_1232,In_2075,In_2257);
xor U1233 (N_1233,In_162,In_2310);
nor U1234 (N_1234,In_1399,In_1833);
nand U1235 (N_1235,In_1254,In_1906);
nor U1236 (N_1236,In_629,In_415);
nor U1237 (N_1237,In_193,In_2861);
nor U1238 (N_1238,In_1352,In_1915);
xor U1239 (N_1239,In_1569,In_1902);
xnor U1240 (N_1240,In_2821,In_484);
and U1241 (N_1241,In_1155,In_2709);
xor U1242 (N_1242,In_1893,In_2519);
nor U1243 (N_1243,In_679,In_1327);
or U1244 (N_1244,In_280,In_1614);
nand U1245 (N_1245,In_2450,In_2025);
nand U1246 (N_1246,In_2516,In_727);
nor U1247 (N_1247,In_2724,In_1351);
or U1248 (N_1248,In_294,In_1681);
nand U1249 (N_1249,In_1712,In_1988);
and U1250 (N_1250,In_2138,In_1339);
nand U1251 (N_1251,In_2975,In_909);
xnor U1252 (N_1252,In_691,In_1212);
or U1253 (N_1253,In_927,In_1941);
nand U1254 (N_1254,In_17,In_1125);
nand U1255 (N_1255,In_176,In_1675);
nand U1256 (N_1256,In_732,In_1316);
nand U1257 (N_1257,In_301,In_2954);
nand U1258 (N_1258,In_1707,In_275);
or U1259 (N_1259,In_73,In_2276);
nor U1260 (N_1260,In_1692,In_2459);
nor U1261 (N_1261,In_1512,In_1331);
nand U1262 (N_1262,In_1550,In_2915);
and U1263 (N_1263,In_525,In_2521);
xnor U1264 (N_1264,In_2317,In_865);
nand U1265 (N_1265,In_980,In_2523);
xnor U1266 (N_1266,In_2986,In_494);
or U1267 (N_1267,In_2650,In_1592);
xor U1268 (N_1268,In_1446,In_1240);
and U1269 (N_1269,In_1626,In_380);
and U1270 (N_1270,In_53,In_2611);
or U1271 (N_1271,In_941,In_41);
nand U1272 (N_1272,In_784,In_89);
nor U1273 (N_1273,In_2748,In_1219);
xor U1274 (N_1274,In_2221,In_851);
or U1275 (N_1275,In_1886,In_520);
nand U1276 (N_1276,In_219,In_919);
xnor U1277 (N_1277,In_1566,In_1541);
nor U1278 (N_1278,In_572,In_2596);
nand U1279 (N_1279,In_1970,In_648);
nor U1280 (N_1280,In_302,In_25);
and U1281 (N_1281,In_2497,In_1208);
nor U1282 (N_1282,In_776,In_1999);
nor U1283 (N_1283,In_2942,In_2271);
and U1284 (N_1284,In_218,In_2189);
nor U1285 (N_1285,In_149,In_1522);
nand U1286 (N_1286,In_1361,In_632);
and U1287 (N_1287,In_2594,In_2299);
xor U1288 (N_1288,In_1259,In_1237);
and U1289 (N_1289,In_638,In_2711);
xor U1290 (N_1290,In_2958,In_539);
or U1291 (N_1291,In_1756,In_1484);
nor U1292 (N_1292,In_2866,In_1478);
or U1293 (N_1293,In_434,In_2695);
or U1294 (N_1294,In_2953,In_1430);
and U1295 (N_1295,In_208,In_2485);
nand U1296 (N_1296,In_1981,In_1953);
nand U1297 (N_1297,In_2322,In_114);
nand U1298 (N_1298,In_358,In_1255);
nor U1299 (N_1299,In_1265,In_1916);
and U1300 (N_1300,In_1453,In_819);
and U1301 (N_1301,In_800,In_866);
nand U1302 (N_1302,In_2166,In_1253);
or U1303 (N_1303,In_2563,In_2670);
and U1304 (N_1304,In_2801,In_1577);
and U1305 (N_1305,In_1814,In_988);
nor U1306 (N_1306,In_263,In_860);
nor U1307 (N_1307,In_514,In_2558);
nand U1308 (N_1308,In_154,In_2179);
nor U1309 (N_1309,In_108,In_2634);
xnor U1310 (N_1310,In_1497,In_1535);
and U1311 (N_1311,In_1469,In_2824);
xor U1312 (N_1312,In_2362,In_805);
or U1313 (N_1313,In_2967,In_2892);
xnor U1314 (N_1314,In_947,In_2178);
or U1315 (N_1315,In_786,In_298);
and U1316 (N_1316,In_2319,In_2255);
xnor U1317 (N_1317,In_864,In_2872);
and U1318 (N_1318,In_855,In_2471);
xor U1319 (N_1319,In_2681,In_451);
nor U1320 (N_1320,In_990,In_1806);
xnor U1321 (N_1321,In_796,In_2367);
or U1322 (N_1322,In_2649,In_1662);
nand U1323 (N_1323,In_912,In_1002);
nor U1324 (N_1324,In_2882,In_2295);
nand U1325 (N_1325,In_523,In_636);
and U1326 (N_1326,In_2142,In_2086);
nand U1327 (N_1327,In_2668,In_1178);
nor U1328 (N_1328,In_782,In_1051);
and U1329 (N_1329,In_94,In_1323);
nor U1330 (N_1330,In_2336,In_2622);
or U1331 (N_1331,In_2136,In_1508);
and U1332 (N_1332,In_2545,In_1375);
or U1333 (N_1333,In_2263,In_2710);
and U1334 (N_1334,In_1337,In_1138);
or U1335 (N_1335,In_808,In_66);
nand U1336 (N_1336,In_1374,In_2692);
nand U1337 (N_1337,In_113,In_2740);
xnor U1338 (N_1338,In_2232,In_1079);
xor U1339 (N_1339,In_121,In_2916);
nor U1340 (N_1340,In_787,In_1501);
nor U1341 (N_1341,In_1875,In_2698);
xor U1342 (N_1342,In_2194,In_2883);
or U1343 (N_1343,In_2731,In_637);
nand U1344 (N_1344,In_667,In_1439);
nor U1345 (N_1345,In_1095,In_1979);
or U1346 (N_1346,In_630,In_1542);
nor U1347 (N_1347,In_2499,In_1059);
nor U1348 (N_1348,In_1412,In_223);
or U1349 (N_1349,In_102,In_1502);
or U1350 (N_1350,In_2289,In_2298);
nor U1351 (N_1351,In_1665,In_2141);
xnor U1352 (N_1352,In_1101,In_1410);
and U1353 (N_1353,In_87,In_1398);
and U1354 (N_1354,In_448,In_563);
nor U1355 (N_1355,In_2722,In_373);
xnor U1356 (N_1356,In_2225,In_883);
nor U1357 (N_1357,In_2937,In_2651);
or U1358 (N_1358,In_2024,In_337);
and U1359 (N_1359,In_257,In_444);
or U1360 (N_1360,In_281,In_965);
xor U1361 (N_1361,In_818,In_1924);
nor U1362 (N_1362,In_2082,In_2533);
and U1363 (N_1363,In_1879,In_2266);
and U1364 (N_1364,In_2341,In_1392);
nor U1365 (N_1365,In_2586,In_760);
or U1366 (N_1366,In_2123,In_1679);
xnor U1367 (N_1367,In_266,In_584);
nand U1368 (N_1368,In_2918,In_1593);
or U1369 (N_1369,In_955,In_2507);
xor U1370 (N_1370,In_2703,In_384);
xor U1371 (N_1371,In_2121,In_2338);
nor U1372 (N_1372,In_159,In_394);
or U1373 (N_1373,In_871,In_1610);
nor U1374 (N_1374,In_2922,In_2379);
or U1375 (N_1375,In_1910,In_1786);
or U1376 (N_1376,In_1816,In_153);
nor U1377 (N_1377,In_2300,In_821);
and U1378 (N_1378,In_1177,In_367);
nor U1379 (N_1379,In_2652,In_1385);
xor U1380 (N_1380,In_1171,In_790);
nor U1381 (N_1381,In_1077,In_1128);
nand U1382 (N_1382,In_1087,In_2566);
nand U1383 (N_1383,In_532,In_1073);
nor U1384 (N_1384,In_1,In_1424);
nor U1385 (N_1385,In_406,In_1733);
or U1386 (N_1386,In_2985,In_1667);
nand U1387 (N_1387,In_1866,In_192);
and U1388 (N_1388,In_2375,In_209);
and U1389 (N_1389,In_609,In_1141);
and U1390 (N_1390,In_2805,In_1060);
or U1391 (N_1391,In_1805,In_2959);
or U1392 (N_1392,In_189,In_1540);
nand U1393 (N_1393,In_1420,In_1678);
xor U1394 (N_1394,In_817,In_2862);
and U1395 (N_1395,In_2974,In_82);
nor U1396 (N_1396,In_475,In_1861);
nand U1397 (N_1397,In_554,In_2608);
or U1398 (N_1398,In_2186,In_215);
and U1399 (N_1399,In_2213,In_1173);
nor U1400 (N_1400,In_1935,In_2549);
or U1401 (N_1401,In_1481,In_98);
nand U1402 (N_1402,In_1479,In_199);
xor U1403 (N_1403,In_529,In_1700);
or U1404 (N_1404,In_1889,In_2458);
xor U1405 (N_1405,In_903,In_2806);
or U1406 (N_1406,In_1371,In_2309);
nand U1407 (N_1407,In_1822,In_1220);
nor U1408 (N_1408,In_1513,In_1978);
xnor U1409 (N_1409,In_2337,In_1940);
nand U1410 (N_1410,In_2706,In_2894);
nand U1411 (N_1411,In_157,In_363);
and U1412 (N_1412,In_2715,In_247);
xnor U1413 (N_1413,In_2466,In_1617);
and U1414 (N_1414,In_568,In_1461);
or U1415 (N_1415,In_1064,In_2371);
nand U1416 (N_1416,In_1494,In_752);
nor U1417 (N_1417,In_811,In_891);
xnor U1418 (N_1418,In_2402,In_652);
nand U1419 (N_1419,In_2728,In_504);
nor U1420 (N_1420,In_476,In_1993);
and U1421 (N_1421,In_751,In_2415);
nor U1422 (N_1422,In_577,In_2529);
nand U1423 (N_1423,In_2071,In_718);
xor U1424 (N_1424,In_631,In_2815);
nor U1425 (N_1425,In_1216,In_1290);
or U1426 (N_1426,In_2107,In_899);
xor U1427 (N_1427,In_881,In_2048);
nand U1428 (N_1428,In_329,In_1977);
nor U1429 (N_1429,In_1168,In_427);
xnor U1430 (N_1430,In_1356,In_859);
nand U1431 (N_1431,In_1302,In_2057);
and U1432 (N_1432,In_2693,In_51);
nand U1433 (N_1433,In_1613,In_185);
nor U1434 (N_1434,In_1841,In_2043);
and U1435 (N_1435,In_2577,In_734);
or U1436 (N_1436,In_2211,In_1658);
nor U1437 (N_1437,In_1152,In_1835);
nand U1438 (N_1438,In_2990,In_1013);
nand U1439 (N_1439,In_986,In_1176);
and U1440 (N_1440,In_925,In_1832);
or U1441 (N_1441,In_287,In_1810);
and U1442 (N_1442,In_1106,In_1130);
and U1443 (N_1443,In_2447,In_106);
and U1444 (N_1444,In_649,In_13);
xnor U1445 (N_1445,In_1460,In_1996);
nor U1446 (N_1446,In_2357,In_674);
nor U1447 (N_1447,In_915,In_2403);
nand U1448 (N_1448,In_1336,In_1311);
nand U1449 (N_1449,In_2094,In_1373);
nand U1450 (N_1450,In_289,In_904);
nor U1451 (N_1451,In_1090,In_602);
xor U1452 (N_1452,In_1049,In_901);
xnor U1453 (N_1453,In_1357,In_2661);
and U1454 (N_1454,In_748,In_701);
xnor U1455 (N_1455,In_1228,In_2099);
and U1456 (N_1456,In_2230,In_1500);
and U1457 (N_1457,In_1764,In_846);
xnor U1458 (N_1458,In_1319,In_781);
or U1459 (N_1459,In_279,In_1737);
nand U1460 (N_1460,In_1826,In_2020);
and U1461 (N_1461,In_1011,In_1442);
and U1462 (N_1462,In_1888,In_2981);
nand U1463 (N_1463,In_1968,In_1043);
and U1464 (N_1464,In_33,In_794);
nand U1465 (N_1465,In_258,In_2863);
or U1466 (N_1466,In_1994,In_2432);
nor U1467 (N_1467,In_926,In_515);
or U1468 (N_1468,In_72,In_181);
or U1469 (N_1469,In_210,In_1809);
xnor U1470 (N_1470,In_2026,In_2252);
nand U1471 (N_1471,In_1647,In_2093);
nand U1472 (N_1472,In_2788,In_893);
xnor U1473 (N_1473,In_1767,In_1108);
or U1474 (N_1474,In_74,In_1286);
nor U1475 (N_1475,In_43,In_2400);
nand U1476 (N_1476,In_517,In_2095);
nand U1477 (N_1477,In_1427,In_706);
xor U1478 (N_1478,In_997,In_318);
nand U1479 (N_1479,In_700,In_1103);
nor U1480 (N_1480,In_1408,In_2084);
or U1481 (N_1481,In_1422,In_2721);
xnor U1482 (N_1482,In_976,In_1450);
or U1483 (N_1483,In_2014,In_1728);
and U1484 (N_1484,In_1440,In_1206);
nand U1485 (N_1485,In_1975,In_1449);
or U1486 (N_1486,In_1874,In_1483);
and U1487 (N_1487,In_780,In_622);
and U1488 (N_1488,In_1068,In_129);
xnor U1489 (N_1489,In_2546,In_429);
xnor U1490 (N_1490,In_1342,In_2964);
nor U1491 (N_1491,In_341,In_1942);
and U1492 (N_1492,In_1818,In_1802);
xor U1493 (N_1493,In_2177,In_942);
and U1494 (N_1494,In_2368,In_528);
xnor U1495 (N_1495,In_731,In_1834);
xor U1496 (N_1496,In_1840,In_1160);
nand U1497 (N_1497,In_1234,In_2572);
nand U1498 (N_1498,In_1892,In_607);
xnor U1499 (N_1499,In_2818,In_1664);
nand U1500 (N_1500,In_2748,In_2838);
xnor U1501 (N_1501,In_350,In_1419);
or U1502 (N_1502,In_2560,In_292);
and U1503 (N_1503,In_2900,In_514);
nor U1504 (N_1504,In_876,In_1327);
and U1505 (N_1505,In_1866,In_2371);
or U1506 (N_1506,In_2464,In_1660);
xor U1507 (N_1507,In_698,In_928);
nand U1508 (N_1508,In_2792,In_359);
nand U1509 (N_1509,In_744,In_2246);
and U1510 (N_1510,In_377,In_701);
or U1511 (N_1511,In_724,In_369);
nand U1512 (N_1512,In_976,In_1253);
or U1513 (N_1513,In_1601,In_1039);
nor U1514 (N_1514,In_816,In_1521);
and U1515 (N_1515,In_959,In_2025);
or U1516 (N_1516,In_781,In_339);
xnor U1517 (N_1517,In_2548,In_2257);
nand U1518 (N_1518,In_602,In_2771);
or U1519 (N_1519,In_1003,In_2309);
and U1520 (N_1520,In_954,In_1274);
nand U1521 (N_1521,In_1216,In_1969);
and U1522 (N_1522,In_2002,In_941);
and U1523 (N_1523,In_194,In_2755);
and U1524 (N_1524,In_1541,In_2919);
xnor U1525 (N_1525,In_586,In_413);
nand U1526 (N_1526,In_1533,In_2758);
nand U1527 (N_1527,In_1237,In_946);
xor U1528 (N_1528,In_961,In_2954);
xor U1529 (N_1529,In_2740,In_647);
nand U1530 (N_1530,In_906,In_2202);
nand U1531 (N_1531,In_940,In_565);
xnor U1532 (N_1532,In_530,In_1467);
nand U1533 (N_1533,In_669,In_1038);
nor U1534 (N_1534,In_2053,In_201);
or U1535 (N_1535,In_2482,In_2126);
and U1536 (N_1536,In_255,In_902);
or U1537 (N_1537,In_529,In_134);
nor U1538 (N_1538,In_2191,In_520);
nand U1539 (N_1539,In_1764,In_206);
nand U1540 (N_1540,In_2493,In_597);
nor U1541 (N_1541,In_617,In_163);
xor U1542 (N_1542,In_1918,In_499);
or U1543 (N_1543,In_1515,In_1555);
or U1544 (N_1544,In_932,In_1352);
or U1545 (N_1545,In_2007,In_1352);
and U1546 (N_1546,In_1888,In_235);
xor U1547 (N_1547,In_2358,In_1729);
or U1548 (N_1548,In_2701,In_2680);
or U1549 (N_1549,In_2877,In_1146);
and U1550 (N_1550,In_1613,In_1906);
or U1551 (N_1551,In_722,In_1941);
nand U1552 (N_1552,In_1059,In_88);
or U1553 (N_1553,In_2073,In_146);
and U1554 (N_1554,In_2084,In_1385);
xnor U1555 (N_1555,In_433,In_1100);
or U1556 (N_1556,In_1314,In_2624);
or U1557 (N_1557,In_2778,In_198);
nor U1558 (N_1558,In_963,In_589);
and U1559 (N_1559,In_1991,In_2376);
xnor U1560 (N_1560,In_2961,In_161);
nand U1561 (N_1561,In_2617,In_1604);
xor U1562 (N_1562,In_1907,In_2522);
xor U1563 (N_1563,In_1170,In_819);
or U1564 (N_1564,In_1305,In_1429);
nand U1565 (N_1565,In_2526,In_873);
xor U1566 (N_1566,In_1804,In_208);
xor U1567 (N_1567,In_705,In_1615);
or U1568 (N_1568,In_2141,In_1266);
nor U1569 (N_1569,In_1396,In_1100);
nor U1570 (N_1570,In_1675,In_2929);
and U1571 (N_1571,In_1830,In_2954);
or U1572 (N_1572,In_1167,In_2173);
and U1573 (N_1573,In_810,In_2518);
nand U1574 (N_1574,In_1445,In_2779);
and U1575 (N_1575,In_849,In_1341);
and U1576 (N_1576,In_146,In_288);
and U1577 (N_1577,In_968,In_2224);
or U1578 (N_1578,In_392,In_2425);
xor U1579 (N_1579,In_1519,In_552);
xnor U1580 (N_1580,In_1487,In_1467);
or U1581 (N_1581,In_1595,In_2380);
nand U1582 (N_1582,In_2127,In_383);
or U1583 (N_1583,In_723,In_2938);
nand U1584 (N_1584,In_1664,In_786);
and U1585 (N_1585,In_1678,In_2888);
and U1586 (N_1586,In_1041,In_973);
and U1587 (N_1587,In_2871,In_1256);
or U1588 (N_1588,In_1779,In_1151);
and U1589 (N_1589,In_126,In_2644);
or U1590 (N_1590,In_1250,In_1940);
xor U1591 (N_1591,In_124,In_727);
or U1592 (N_1592,In_2254,In_45);
xnor U1593 (N_1593,In_424,In_2256);
xor U1594 (N_1594,In_1149,In_1717);
nand U1595 (N_1595,In_90,In_1339);
or U1596 (N_1596,In_837,In_1396);
and U1597 (N_1597,In_1672,In_605);
and U1598 (N_1598,In_1245,In_971);
and U1599 (N_1599,In_403,In_2476);
or U1600 (N_1600,In_708,In_523);
nor U1601 (N_1601,In_1356,In_2702);
or U1602 (N_1602,In_996,In_929);
nand U1603 (N_1603,In_2719,In_748);
xor U1604 (N_1604,In_277,In_2818);
and U1605 (N_1605,In_1503,In_2504);
and U1606 (N_1606,In_1948,In_404);
nand U1607 (N_1607,In_2758,In_2429);
xnor U1608 (N_1608,In_2024,In_1199);
and U1609 (N_1609,In_208,In_1089);
nand U1610 (N_1610,In_1354,In_1130);
or U1611 (N_1611,In_1014,In_2580);
nor U1612 (N_1612,In_268,In_1199);
xor U1613 (N_1613,In_680,In_475);
nor U1614 (N_1614,In_641,In_165);
and U1615 (N_1615,In_2008,In_976);
nand U1616 (N_1616,In_15,In_1838);
nor U1617 (N_1617,In_657,In_727);
xnor U1618 (N_1618,In_1915,In_568);
and U1619 (N_1619,In_1210,In_1362);
and U1620 (N_1620,In_2505,In_54);
or U1621 (N_1621,In_1938,In_1381);
xor U1622 (N_1622,In_2957,In_679);
xnor U1623 (N_1623,In_364,In_2872);
or U1624 (N_1624,In_2778,In_1819);
and U1625 (N_1625,In_1623,In_483);
and U1626 (N_1626,In_970,In_681);
xnor U1627 (N_1627,In_1903,In_1714);
or U1628 (N_1628,In_407,In_57);
nand U1629 (N_1629,In_1627,In_1234);
nand U1630 (N_1630,In_2334,In_321);
or U1631 (N_1631,In_1850,In_2741);
nor U1632 (N_1632,In_2273,In_287);
or U1633 (N_1633,In_1381,In_420);
nand U1634 (N_1634,In_814,In_2878);
or U1635 (N_1635,In_2189,In_320);
and U1636 (N_1636,In_1502,In_504);
nor U1637 (N_1637,In_1380,In_414);
or U1638 (N_1638,In_2029,In_2556);
and U1639 (N_1639,In_1106,In_2205);
nand U1640 (N_1640,In_914,In_239);
and U1641 (N_1641,In_110,In_2575);
xor U1642 (N_1642,In_282,In_2526);
and U1643 (N_1643,In_1146,In_249);
xor U1644 (N_1644,In_2960,In_1560);
or U1645 (N_1645,In_150,In_2670);
nor U1646 (N_1646,In_1951,In_920);
nand U1647 (N_1647,In_1494,In_1744);
nand U1648 (N_1648,In_372,In_1471);
nor U1649 (N_1649,In_1057,In_1152);
or U1650 (N_1650,In_439,In_2757);
nand U1651 (N_1651,In_785,In_771);
nand U1652 (N_1652,In_1476,In_956);
or U1653 (N_1653,In_1129,In_1601);
or U1654 (N_1654,In_2501,In_2440);
or U1655 (N_1655,In_1067,In_1086);
xor U1656 (N_1656,In_2579,In_645);
and U1657 (N_1657,In_703,In_1131);
nor U1658 (N_1658,In_2032,In_703);
nor U1659 (N_1659,In_847,In_198);
nor U1660 (N_1660,In_2104,In_1525);
and U1661 (N_1661,In_901,In_211);
and U1662 (N_1662,In_2060,In_2507);
or U1663 (N_1663,In_1695,In_2522);
nand U1664 (N_1664,In_2963,In_2012);
and U1665 (N_1665,In_328,In_471);
and U1666 (N_1666,In_1931,In_2607);
nor U1667 (N_1667,In_2714,In_2207);
nand U1668 (N_1668,In_596,In_1937);
nand U1669 (N_1669,In_186,In_1531);
and U1670 (N_1670,In_335,In_2150);
or U1671 (N_1671,In_1538,In_121);
xnor U1672 (N_1672,In_373,In_2987);
xnor U1673 (N_1673,In_576,In_137);
xnor U1674 (N_1674,In_1569,In_834);
nand U1675 (N_1675,In_1155,In_1946);
and U1676 (N_1676,In_869,In_1716);
nor U1677 (N_1677,In_1028,In_1630);
and U1678 (N_1678,In_980,In_1400);
and U1679 (N_1679,In_1212,In_1232);
and U1680 (N_1680,In_1384,In_994);
or U1681 (N_1681,In_2328,In_978);
xnor U1682 (N_1682,In_1101,In_363);
or U1683 (N_1683,In_603,In_1243);
and U1684 (N_1684,In_381,In_1200);
xnor U1685 (N_1685,In_793,In_1185);
or U1686 (N_1686,In_1484,In_1335);
or U1687 (N_1687,In_753,In_2607);
nand U1688 (N_1688,In_1321,In_2622);
or U1689 (N_1689,In_1648,In_2764);
nand U1690 (N_1690,In_1876,In_2853);
nand U1691 (N_1691,In_1280,In_661);
or U1692 (N_1692,In_2737,In_710);
nand U1693 (N_1693,In_1301,In_745);
nor U1694 (N_1694,In_40,In_2299);
and U1695 (N_1695,In_2085,In_2948);
nor U1696 (N_1696,In_2263,In_1894);
and U1697 (N_1697,In_1222,In_2964);
xnor U1698 (N_1698,In_2862,In_1316);
and U1699 (N_1699,In_1133,In_501);
or U1700 (N_1700,In_2410,In_2646);
nand U1701 (N_1701,In_2318,In_2835);
and U1702 (N_1702,In_1794,In_1445);
nor U1703 (N_1703,In_1284,In_2329);
and U1704 (N_1704,In_219,In_328);
nand U1705 (N_1705,In_2792,In_65);
and U1706 (N_1706,In_2952,In_1215);
xnor U1707 (N_1707,In_633,In_2573);
nand U1708 (N_1708,In_2397,In_225);
and U1709 (N_1709,In_2962,In_1742);
nand U1710 (N_1710,In_832,In_1940);
nand U1711 (N_1711,In_1049,In_1428);
nand U1712 (N_1712,In_258,In_855);
nor U1713 (N_1713,In_2514,In_2134);
xnor U1714 (N_1714,In_17,In_324);
nor U1715 (N_1715,In_2066,In_2627);
nor U1716 (N_1716,In_2451,In_2357);
nor U1717 (N_1717,In_1036,In_968);
nor U1718 (N_1718,In_739,In_93);
nand U1719 (N_1719,In_835,In_1616);
xnor U1720 (N_1720,In_390,In_1156);
or U1721 (N_1721,In_323,In_1527);
and U1722 (N_1722,In_1131,In_688);
or U1723 (N_1723,In_58,In_1695);
or U1724 (N_1724,In_2280,In_917);
nor U1725 (N_1725,In_1618,In_1890);
and U1726 (N_1726,In_980,In_514);
nor U1727 (N_1727,In_1811,In_2112);
and U1728 (N_1728,In_1571,In_2237);
or U1729 (N_1729,In_689,In_2098);
nand U1730 (N_1730,In_367,In_2730);
xnor U1731 (N_1731,In_989,In_1846);
nand U1732 (N_1732,In_2417,In_2845);
xor U1733 (N_1733,In_1298,In_1340);
nor U1734 (N_1734,In_2745,In_1244);
or U1735 (N_1735,In_2582,In_734);
nor U1736 (N_1736,In_2970,In_2931);
nor U1737 (N_1737,In_1120,In_1806);
and U1738 (N_1738,In_2768,In_316);
nand U1739 (N_1739,In_2465,In_2497);
nor U1740 (N_1740,In_2372,In_2877);
and U1741 (N_1741,In_1809,In_50);
or U1742 (N_1742,In_2778,In_2623);
xnor U1743 (N_1743,In_1863,In_2313);
or U1744 (N_1744,In_1918,In_2284);
nand U1745 (N_1745,In_357,In_2564);
and U1746 (N_1746,In_749,In_2407);
nand U1747 (N_1747,In_1428,In_966);
xnor U1748 (N_1748,In_2527,In_2108);
nand U1749 (N_1749,In_2421,In_1061);
or U1750 (N_1750,In_94,In_2362);
and U1751 (N_1751,In_2145,In_559);
xnor U1752 (N_1752,In_1065,In_1057);
or U1753 (N_1753,In_2797,In_2896);
xnor U1754 (N_1754,In_220,In_1616);
and U1755 (N_1755,In_1700,In_2069);
and U1756 (N_1756,In_717,In_2202);
and U1757 (N_1757,In_2402,In_2178);
xor U1758 (N_1758,In_1790,In_2562);
nor U1759 (N_1759,In_964,In_2177);
nor U1760 (N_1760,In_1697,In_2073);
nand U1761 (N_1761,In_2201,In_1473);
nor U1762 (N_1762,In_1227,In_1637);
nand U1763 (N_1763,In_519,In_1914);
xor U1764 (N_1764,In_1378,In_864);
and U1765 (N_1765,In_755,In_1545);
and U1766 (N_1766,In_873,In_1326);
nor U1767 (N_1767,In_1128,In_1505);
or U1768 (N_1768,In_2840,In_118);
nor U1769 (N_1769,In_2117,In_915);
nand U1770 (N_1770,In_894,In_683);
or U1771 (N_1771,In_2875,In_2347);
nor U1772 (N_1772,In_2265,In_1534);
or U1773 (N_1773,In_998,In_888);
or U1774 (N_1774,In_2773,In_1443);
xor U1775 (N_1775,In_2153,In_1625);
or U1776 (N_1776,In_516,In_2428);
nand U1777 (N_1777,In_2365,In_2345);
or U1778 (N_1778,In_2587,In_527);
or U1779 (N_1779,In_192,In_1650);
xnor U1780 (N_1780,In_1676,In_2047);
xnor U1781 (N_1781,In_1296,In_1729);
nand U1782 (N_1782,In_1777,In_2624);
nand U1783 (N_1783,In_2484,In_564);
nand U1784 (N_1784,In_2489,In_203);
nor U1785 (N_1785,In_248,In_411);
or U1786 (N_1786,In_1279,In_2178);
or U1787 (N_1787,In_1818,In_1548);
nor U1788 (N_1788,In_2493,In_942);
or U1789 (N_1789,In_1504,In_2898);
nor U1790 (N_1790,In_2746,In_2219);
nor U1791 (N_1791,In_109,In_500);
nand U1792 (N_1792,In_828,In_2598);
xor U1793 (N_1793,In_1415,In_2409);
nor U1794 (N_1794,In_2554,In_2672);
xor U1795 (N_1795,In_2463,In_2286);
or U1796 (N_1796,In_40,In_1918);
and U1797 (N_1797,In_2215,In_1681);
or U1798 (N_1798,In_149,In_1477);
and U1799 (N_1799,In_2083,In_589);
or U1800 (N_1800,In_321,In_1266);
or U1801 (N_1801,In_1666,In_2397);
or U1802 (N_1802,In_2573,In_2377);
nor U1803 (N_1803,In_2198,In_1288);
xor U1804 (N_1804,In_855,In_1457);
and U1805 (N_1805,In_106,In_1020);
nor U1806 (N_1806,In_231,In_2322);
or U1807 (N_1807,In_1662,In_355);
xor U1808 (N_1808,In_1356,In_2869);
xnor U1809 (N_1809,In_940,In_1336);
and U1810 (N_1810,In_1423,In_1942);
and U1811 (N_1811,In_2215,In_1636);
or U1812 (N_1812,In_2306,In_220);
nand U1813 (N_1813,In_2937,In_1553);
and U1814 (N_1814,In_1295,In_544);
xor U1815 (N_1815,In_2759,In_957);
nor U1816 (N_1816,In_2559,In_2033);
xor U1817 (N_1817,In_2433,In_2556);
and U1818 (N_1818,In_2309,In_1368);
and U1819 (N_1819,In_2043,In_1407);
nand U1820 (N_1820,In_2422,In_1246);
nor U1821 (N_1821,In_2648,In_1957);
xnor U1822 (N_1822,In_1197,In_264);
or U1823 (N_1823,In_27,In_883);
and U1824 (N_1824,In_1318,In_2515);
xnor U1825 (N_1825,In_1016,In_353);
and U1826 (N_1826,In_422,In_531);
or U1827 (N_1827,In_1815,In_77);
xnor U1828 (N_1828,In_2,In_1016);
nor U1829 (N_1829,In_781,In_1346);
nand U1830 (N_1830,In_1482,In_2740);
or U1831 (N_1831,In_1064,In_1188);
or U1832 (N_1832,In_2288,In_2738);
and U1833 (N_1833,In_1676,In_2987);
and U1834 (N_1834,In_239,In_1418);
nand U1835 (N_1835,In_756,In_2169);
nor U1836 (N_1836,In_725,In_1472);
nor U1837 (N_1837,In_965,In_321);
and U1838 (N_1838,In_807,In_1439);
nor U1839 (N_1839,In_1739,In_1686);
or U1840 (N_1840,In_348,In_2734);
and U1841 (N_1841,In_2038,In_2820);
xnor U1842 (N_1842,In_1536,In_42);
nor U1843 (N_1843,In_956,In_24);
or U1844 (N_1844,In_2197,In_1234);
xor U1845 (N_1845,In_1901,In_1907);
or U1846 (N_1846,In_24,In_1149);
or U1847 (N_1847,In_2976,In_1287);
and U1848 (N_1848,In_582,In_1918);
nor U1849 (N_1849,In_44,In_1711);
nor U1850 (N_1850,In_2292,In_1840);
xor U1851 (N_1851,In_2435,In_2410);
or U1852 (N_1852,In_2225,In_256);
nor U1853 (N_1853,In_1678,In_1978);
or U1854 (N_1854,In_2738,In_1397);
nand U1855 (N_1855,In_2374,In_2656);
xnor U1856 (N_1856,In_2412,In_1119);
or U1857 (N_1857,In_1360,In_783);
xor U1858 (N_1858,In_2102,In_1614);
nand U1859 (N_1859,In_1256,In_314);
xnor U1860 (N_1860,In_2415,In_2602);
xor U1861 (N_1861,In_2252,In_14);
nor U1862 (N_1862,In_150,In_144);
nor U1863 (N_1863,In_25,In_1637);
nand U1864 (N_1864,In_1544,In_102);
xor U1865 (N_1865,In_2633,In_1805);
or U1866 (N_1866,In_2056,In_384);
xnor U1867 (N_1867,In_216,In_2576);
and U1868 (N_1868,In_1686,In_593);
nor U1869 (N_1869,In_1841,In_1140);
nor U1870 (N_1870,In_435,In_1588);
or U1871 (N_1871,In_2336,In_1283);
nor U1872 (N_1872,In_1108,In_2496);
nand U1873 (N_1873,In_1871,In_613);
xor U1874 (N_1874,In_216,In_828);
xor U1875 (N_1875,In_548,In_953);
or U1876 (N_1876,In_490,In_1298);
nand U1877 (N_1877,In_178,In_1386);
nor U1878 (N_1878,In_2765,In_2833);
nand U1879 (N_1879,In_731,In_2084);
nor U1880 (N_1880,In_908,In_2903);
nand U1881 (N_1881,In_1850,In_577);
and U1882 (N_1882,In_1692,In_132);
xnor U1883 (N_1883,In_54,In_1622);
and U1884 (N_1884,In_1489,In_610);
nand U1885 (N_1885,In_875,In_2544);
xor U1886 (N_1886,In_1429,In_2659);
or U1887 (N_1887,In_308,In_219);
and U1888 (N_1888,In_1750,In_323);
or U1889 (N_1889,In_1412,In_2307);
and U1890 (N_1890,In_2606,In_978);
or U1891 (N_1891,In_2492,In_153);
xnor U1892 (N_1892,In_2806,In_1577);
nand U1893 (N_1893,In_978,In_234);
or U1894 (N_1894,In_1556,In_213);
xnor U1895 (N_1895,In_2966,In_2124);
nor U1896 (N_1896,In_2332,In_2291);
nand U1897 (N_1897,In_1023,In_1667);
nor U1898 (N_1898,In_2724,In_480);
nor U1899 (N_1899,In_2413,In_319);
or U1900 (N_1900,In_503,In_1908);
xnor U1901 (N_1901,In_2992,In_434);
or U1902 (N_1902,In_2146,In_2363);
and U1903 (N_1903,In_2982,In_2553);
and U1904 (N_1904,In_1859,In_2004);
nand U1905 (N_1905,In_1064,In_259);
or U1906 (N_1906,In_2137,In_940);
nor U1907 (N_1907,In_576,In_1718);
xor U1908 (N_1908,In_862,In_1568);
nor U1909 (N_1909,In_2980,In_947);
xnor U1910 (N_1910,In_1872,In_2077);
nor U1911 (N_1911,In_1444,In_2478);
nor U1912 (N_1912,In_969,In_2974);
xor U1913 (N_1913,In_1982,In_516);
nor U1914 (N_1914,In_2853,In_255);
or U1915 (N_1915,In_706,In_250);
nor U1916 (N_1916,In_1457,In_1049);
nand U1917 (N_1917,In_590,In_2996);
nand U1918 (N_1918,In_2510,In_1202);
nand U1919 (N_1919,In_2980,In_2605);
and U1920 (N_1920,In_116,In_232);
nand U1921 (N_1921,In_2649,In_1583);
nor U1922 (N_1922,In_2536,In_1655);
xor U1923 (N_1923,In_2678,In_2572);
nand U1924 (N_1924,In_1003,In_889);
or U1925 (N_1925,In_2552,In_591);
nand U1926 (N_1926,In_2773,In_22);
nand U1927 (N_1927,In_1031,In_616);
and U1928 (N_1928,In_1314,In_2964);
or U1929 (N_1929,In_849,In_2268);
and U1930 (N_1930,In_1201,In_716);
or U1931 (N_1931,In_1761,In_1516);
and U1932 (N_1932,In_1730,In_1590);
and U1933 (N_1933,In_507,In_2747);
xnor U1934 (N_1934,In_2428,In_848);
xor U1935 (N_1935,In_1246,In_838);
nand U1936 (N_1936,In_136,In_2050);
or U1937 (N_1937,In_579,In_1836);
nand U1938 (N_1938,In_1403,In_1889);
and U1939 (N_1939,In_1108,In_2380);
and U1940 (N_1940,In_2594,In_721);
and U1941 (N_1941,In_228,In_1865);
nand U1942 (N_1942,In_182,In_1835);
or U1943 (N_1943,In_1235,In_1716);
and U1944 (N_1944,In_2321,In_1553);
or U1945 (N_1945,In_2457,In_2206);
and U1946 (N_1946,In_2401,In_548);
nor U1947 (N_1947,In_907,In_303);
xnor U1948 (N_1948,In_470,In_2634);
and U1949 (N_1949,In_1300,In_2399);
nor U1950 (N_1950,In_252,In_190);
nand U1951 (N_1951,In_2420,In_916);
or U1952 (N_1952,In_2118,In_970);
and U1953 (N_1953,In_335,In_47);
xor U1954 (N_1954,In_2997,In_2698);
nor U1955 (N_1955,In_2312,In_2350);
nor U1956 (N_1956,In_1405,In_764);
nor U1957 (N_1957,In_478,In_184);
nor U1958 (N_1958,In_2046,In_252);
or U1959 (N_1959,In_486,In_1093);
nand U1960 (N_1960,In_1443,In_2157);
nor U1961 (N_1961,In_2426,In_2824);
nand U1962 (N_1962,In_2399,In_2205);
nand U1963 (N_1963,In_911,In_1772);
nor U1964 (N_1964,In_1991,In_2728);
nand U1965 (N_1965,In_1094,In_533);
nand U1966 (N_1966,In_2048,In_965);
nand U1967 (N_1967,In_193,In_2184);
and U1968 (N_1968,In_2773,In_2105);
and U1969 (N_1969,In_1849,In_2836);
nor U1970 (N_1970,In_387,In_2218);
and U1971 (N_1971,In_649,In_1338);
or U1972 (N_1972,In_2398,In_2664);
and U1973 (N_1973,In_2355,In_1370);
or U1974 (N_1974,In_2835,In_2289);
xor U1975 (N_1975,In_68,In_1711);
nand U1976 (N_1976,In_1375,In_667);
xor U1977 (N_1977,In_1173,In_2286);
xnor U1978 (N_1978,In_1303,In_144);
xnor U1979 (N_1979,In_1743,In_1855);
xor U1980 (N_1980,In_1901,In_982);
or U1981 (N_1981,In_2172,In_2379);
and U1982 (N_1982,In_1217,In_2772);
nor U1983 (N_1983,In_470,In_488);
or U1984 (N_1984,In_2114,In_276);
xnor U1985 (N_1985,In_390,In_2452);
nand U1986 (N_1986,In_697,In_2603);
nor U1987 (N_1987,In_492,In_1004);
nor U1988 (N_1988,In_523,In_2949);
xnor U1989 (N_1989,In_2464,In_2684);
nor U1990 (N_1990,In_2236,In_1275);
nor U1991 (N_1991,In_2553,In_1026);
and U1992 (N_1992,In_2735,In_1001);
xor U1993 (N_1993,In_1991,In_1683);
and U1994 (N_1994,In_1042,In_108);
or U1995 (N_1995,In_2517,In_1267);
or U1996 (N_1996,In_156,In_323);
xnor U1997 (N_1997,In_2874,In_2456);
nor U1998 (N_1998,In_701,In_2168);
xnor U1999 (N_1999,In_631,In_2705);
nand U2000 (N_2000,In_2834,In_2498);
and U2001 (N_2001,In_773,In_269);
or U2002 (N_2002,In_1912,In_1642);
xnor U2003 (N_2003,In_78,In_1926);
nand U2004 (N_2004,In_2501,In_2738);
nand U2005 (N_2005,In_970,In_1490);
nand U2006 (N_2006,In_2654,In_2568);
nor U2007 (N_2007,In_860,In_1668);
xnor U2008 (N_2008,In_96,In_600);
nor U2009 (N_2009,In_1779,In_2110);
or U2010 (N_2010,In_2804,In_2453);
nor U2011 (N_2011,In_356,In_887);
and U2012 (N_2012,In_72,In_2487);
nor U2013 (N_2013,In_2477,In_220);
xnor U2014 (N_2014,In_100,In_883);
or U2015 (N_2015,In_909,In_2128);
or U2016 (N_2016,In_2221,In_829);
or U2017 (N_2017,In_2794,In_2273);
nand U2018 (N_2018,In_2888,In_2121);
nor U2019 (N_2019,In_1249,In_947);
and U2020 (N_2020,In_1467,In_207);
nor U2021 (N_2021,In_1391,In_64);
or U2022 (N_2022,In_204,In_266);
xor U2023 (N_2023,In_2153,In_1323);
nor U2024 (N_2024,In_1378,In_1192);
and U2025 (N_2025,In_983,In_1398);
nand U2026 (N_2026,In_1125,In_422);
or U2027 (N_2027,In_1106,In_1098);
nor U2028 (N_2028,In_1596,In_163);
or U2029 (N_2029,In_2431,In_943);
nor U2030 (N_2030,In_2019,In_940);
xnor U2031 (N_2031,In_94,In_1677);
or U2032 (N_2032,In_2343,In_2961);
or U2033 (N_2033,In_2372,In_2087);
nor U2034 (N_2034,In_651,In_953);
or U2035 (N_2035,In_993,In_1737);
xor U2036 (N_2036,In_293,In_2239);
and U2037 (N_2037,In_2868,In_1108);
or U2038 (N_2038,In_390,In_973);
nand U2039 (N_2039,In_165,In_219);
and U2040 (N_2040,In_281,In_402);
or U2041 (N_2041,In_1063,In_1285);
xnor U2042 (N_2042,In_2536,In_2108);
nand U2043 (N_2043,In_1907,In_2237);
nand U2044 (N_2044,In_456,In_1769);
nor U2045 (N_2045,In_2314,In_1779);
and U2046 (N_2046,In_815,In_1973);
and U2047 (N_2047,In_2909,In_2076);
or U2048 (N_2048,In_546,In_776);
and U2049 (N_2049,In_2476,In_2389);
nor U2050 (N_2050,In_501,In_285);
nand U2051 (N_2051,In_2408,In_1762);
xor U2052 (N_2052,In_1083,In_2555);
and U2053 (N_2053,In_1440,In_1005);
or U2054 (N_2054,In_2052,In_829);
nor U2055 (N_2055,In_2251,In_2474);
and U2056 (N_2056,In_1971,In_581);
and U2057 (N_2057,In_1877,In_1333);
nand U2058 (N_2058,In_484,In_1369);
nor U2059 (N_2059,In_1507,In_495);
or U2060 (N_2060,In_1776,In_1368);
xor U2061 (N_2061,In_70,In_903);
xnor U2062 (N_2062,In_1646,In_389);
xor U2063 (N_2063,In_1605,In_1928);
xor U2064 (N_2064,In_124,In_1360);
and U2065 (N_2065,In_1184,In_1408);
and U2066 (N_2066,In_1296,In_1555);
nand U2067 (N_2067,In_72,In_314);
nor U2068 (N_2068,In_1367,In_1400);
nand U2069 (N_2069,In_1435,In_2737);
nor U2070 (N_2070,In_1215,In_446);
or U2071 (N_2071,In_32,In_1353);
or U2072 (N_2072,In_1970,In_1975);
xor U2073 (N_2073,In_890,In_2459);
xnor U2074 (N_2074,In_2158,In_2535);
or U2075 (N_2075,In_1515,In_1685);
and U2076 (N_2076,In_309,In_1624);
xnor U2077 (N_2077,In_2628,In_2737);
nand U2078 (N_2078,In_382,In_2560);
xor U2079 (N_2079,In_377,In_834);
and U2080 (N_2080,In_364,In_2722);
nand U2081 (N_2081,In_548,In_1089);
and U2082 (N_2082,In_2039,In_1566);
nand U2083 (N_2083,In_672,In_1135);
or U2084 (N_2084,In_341,In_1402);
or U2085 (N_2085,In_2865,In_1603);
nand U2086 (N_2086,In_2015,In_1902);
nand U2087 (N_2087,In_525,In_2049);
and U2088 (N_2088,In_100,In_2821);
or U2089 (N_2089,In_2840,In_476);
nand U2090 (N_2090,In_189,In_1600);
xor U2091 (N_2091,In_2615,In_2823);
or U2092 (N_2092,In_2307,In_1192);
xor U2093 (N_2093,In_42,In_1951);
and U2094 (N_2094,In_1885,In_1341);
nor U2095 (N_2095,In_1146,In_1554);
or U2096 (N_2096,In_1572,In_2474);
or U2097 (N_2097,In_916,In_1107);
nand U2098 (N_2098,In_1070,In_616);
nand U2099 (N_2099,In_103,In_2308);
and U2100 (N_2100,In_993,In_2933);
nand U2101 (N_2101,In_111,In_2162);
or U2102 (N_2102,In_908,In_2825);
nor U2103 (N_2103,In_2316,In_626);
or U2104 (N_2104,In_398,In_2122);
nor U2105 (N_2105,In_2937,In_2980);
xor U2106 (N_2106,In_1120,In_2359);
xnor U2107 (N_2107,In_97,In_1740);
xor U2108 (N_2108,In_16,In_476);
nor U2109 (N_2109,In_776,In_2682);
and U2110 (N_2110,In_1682,In_788);
nand U2111 (N_2111,In_1181,In_1688);
or U2112 (N_2112,In_460,In_2433);
or U2113 (N_2113,In_783,In_420);
nand U2114 (N_2114,In_101,In_987);
xnor U2115 (N_2115,In_2275,In_1292);
nor U2116 (N_2116,In_994,In_954);
and U2117 (N_2117,In_1817,In_1233);
nor U2118 (N_2118,In_785,In_1106);
or U2119 (N_2119,In_2717,In_1025);
and U2120 (N_2120,In_2012,In_43);
or U2121 (N_2121,In_951,In_1372);
and U2122 (N_2122,In_1549,In_2609);
or U2123 (N_2123,In_2150,In_38);
nand U2124 (N_2124,In_1655,In_2754);
or U2125 (N_2125,In_1107,In_83);
xnor U2126 (N_2126,In_2421,In_1861);
xor U2127 (N_2127,In_1600,In_634);
and U2128 (N_2128,In_2319,In_784);
xnor U2129 (N_2129,In_2530,In_1313);
nand U2130 (N_2130,In_2357,In_805);
xor U2131 (N_2131,In_2308,In_2811);
and U2132 (N_2132,In_2992,In_1134);
and U2133 (N_2133,In_2384,In_285);
or U2134 (N_2134,In_463,In_2283);
nand U2135 (N_2135,In_1580,In_537);
or U2136 (N_2136,In_1803,In_1935);
xnor U2137 (N_2137,In_524,In_1224);
or U2138 (N_2138,In_155,In_777);
xnor U2139 (N_2139,In_590,In_1346);
and U2140 (N_2140,In_1036,In_127);
xor U2141 (N_2141,In_2944,In_674);
or U2142 (N_2142,In_39,In_504);
nand U2143 (N_2143,In_650,In_802);
nand U2144 (N_2144,In_2529,In_2652);
and U2145 (N_2145,In_328,In_1804);
xnor U2146 (N_2146,In_2644,In_1506);
and U2147 (N_2147,In_1209,In_1501);
xnor U2148 (N_2148,In_2378,In_2828);
nand U2149 (N_2149,In_108,In_923);
nand U2150 (N_2150,In_1549,In_543);
nor U2151 (N_2151,In_2700,In_1517);
and U2152 (N_2152,In_159,In_144);
nor U2153 (N_2153,In_2085,In_1732);
nand U2154 (N_2154,In_417,In_39);
and U2155 (N_2155,In_726,In_1759);
or U2156 (N_2156,In_1341,In_252);
and U2157 (N_2157,In_1731,In_612);
nand U2158 (N_2158,In_663,In_69);
nand U2159 (N_2159,In_657,In_395);
nand U2160 (N_2160,In_337,In_1601);
or U2161 (N_2161,In_2803,In_1615);
or U2162 (N_2162,In_2811,In_1637);
and U2163 (N_2163,In_2212,In_837);
nand U2164 (N_2164,In_491,In_1880);
nor U2165 (N_2165,In_2960,In_1146);
or U2166 (N_2166,In_2223,In_1215);
nand U2167 (N_2167,In_1359,In_1381);
nand U2168 (N_2168,In_670,In_1106);
nor U2169 (N_2169,In_574,In_1118);
nor U2170 (N_2170,In_2065,In_185);
or U2171 (N_2171,In_2871,In_301);
and U2172 (N_2172,In_1453,In_890);
and U2173 (N_2173,In_2498,In_191);
xor U2174 (N_2174,In_141,In_678);
nand U2175 (N_2175,In_330,In_1835);
and U2176 (N_2176,In_491,In_22);
xor U2177 (N_2177,In_2447,In_1758);
xnor U2178 (N_2178,In_572,In_187);
or U2179 (N_2179,In_1880,In_2298);
nor U2180 (N_2180,In_1021,In_2618);
nor U2181 (N_2181,In_857,In_1682);
nand U2182 (N_2182,In_1348,In_16);
xnor U2183 (N_2183,In_158,In_1754);
xor U2184 (N_2184,In_200,In_2123);
nand U2185 (N_2185,In_392,In_194);
nor U2186 (N_2186,In_70,In_1307);
nor U2187 (N_2187,In_2447,In_381);
and U2188 (N_2188,In_1140,In_764);
and U2189 (N_2189,In_1951,In_2123);
or U2190 (N_2190,In_790,In_470);
or U2191 (N_2191,In_289,In_2291);
nor U2192 (N_2192,In_1927,In_1155);
nor U2193 (N_2193,In_2431,In_2864);
or U2194 (N_2194,In_2972,In_585);
nand U2195 (N_2195,In_395,In_2323);
and U2196 (N_2196,In_570,In_965);
or U2197 (N_2197,In_480,In_586);
nor U2198 (N_2198,In_2501,In_411);
xor U2199 (N_2199,In_2727,In_2951);
or U2200 (N_2200,In_2210,In_1748);
xor U2201 (N_2201,In_178,In_813);
and U2202 (N_2202,In_263,In_1592);
nor U2203 (N_2203,In_2425,In_386);
nor U2204 (N_2204,In_2928,In_1118);
xor U2205 (N_2205,In_116,In_1416);
nand U2206 (N_2206,In_816,In_1722);
nand U2207 (N_2207,In_160,In_2690);
nor U2208 (N_2208,In_2780,In_2350);
xnor U2209 (N_2209,In_859,In_223);
nor U2210 (N_2210,In_1369,In_1298);
and U2211 (N_2211,In_80,In_1480);
nand U2212 (N_2212,In_2270,In_2079);
nor U2213 (N_2213,In_553,In_2661);
or U2214 (N_2214,In_191,In_589);
or U2215 (N_2215,In_1365,In_52);
nor U2216 (N_2216,In_1592,In_494);
and U2217 (N_2217,In_1325,In_2402);
nand U2218 (N_2218,In_837,In_523);
and U2219 (N_2219,In_2707,In_1812);
xor U2220 (N_2220,In_2326,In_1617);
nand U2221 (N_2221,In_2783,In_473);
or U2222 (N_2222,In_1049,In_2217);
or U2223 (N_2223,In_2973,In_2758);
and U2224 (N_2224,In_1760,In_2316);
nand U2225 (N_2225,In_1670,In_560);
or U2226 (N_2226,In_1452,In_2693);
and U2227 (N_2227,In_1210,In_249);
nor U2228 (N_2228,In_2287,In_1362);
nor U2229 (N_2229,In_69,In_1033);
xnor U2230 (N_2230,In_429,In_2228);
nand U2231 (N_2231,In_2544,In_2858);
and U2232 (N_2232,In_2282,In_1924);
or U2233 (N_2233,In_1542,In_1637);
nand U2234 (N_2234,In_734,In_1496);
nand U2235 (N_2235,In_1645,In_2070);
xor U2236 (N_2236,In_1997,In_345);
nor U2237 (N_2237,In_732,In_343);
nand U2238 (N_2238,In_152,In_2986);
or U2239 (N_2239,In_243,In_472);
or U2240 (N_2240,In_2082,In_609);
nand U2241 (N_2241,In_1143,In_344);
nand U2242 (N_2242,In_755,In_2013);
nand U2243 (N_2243,In_1399,In_2002);
and U2244 (N_2244,In_2153,In_888);
xor U2245 (N_2245,In_485,In_1726);
nand U2246 (N_2246,In_1258,In_721);
and U2247 (N_2247,In_1770,In_468);
xnor U2248 (N_2248,In_1758,In_180);
xnor U2249 (N_2249,In_1180,In_296);
xnor U2250 (N_2250,In_1152,In_1519);
nor U2251 (N_2251,In_41,In_2048);
xnor U2252 (N_2252,In_519,In_1636);
xor U2253 (N_2253,In_1666,In_929);
or U2254 (N_2254,In_1014,In_2579);
or U2255 (N_2255,In_2396,In_1988);
nand U2256 (N_2256,In_1681,In_324);
and U2257 (N_2257,In_1316,In_1224);
nor U2258 (N_2258,In_2477,In_643);
and U2259 (N_2259,In_2935,In_2062);
nor U2260 (N_2260,In_161,In_598);
xor U2261 (N_2261,In_1292,In_1969);
nand U2262 (N_2262,In_378,In_2309);
xor U2263 (N_2263,In_1518,In_556);
and U2264 (N_2264,In_1323,In_1539);
nor U2265 (N_2265,In_50,In_2000);
xor U2266 (N_2266,In_1975,In_2307);
nor U2267 (N_2267,In_1527,In_2000);
nand U2268 (N_2268,In_2369,In_1349);
nor U2269 (N_2269,In_165,In_1084);
xnor U2270 (N_2270,In_2662,In_2604);
nor U2271 (N_2271,In_1086,In_1324);
nand U2272 (N_2272,In_2994,In_962);
and U2273 (N_2273,In_160,In_1762);
xnor U2274 (N_2274,In_2763,In_1610);
xnor U2275 (N_2275,In_129,In_185);
nand U2276 (N_2276,In_1289,In_756);
xor U2277 (N_2277,In_2267,In_1875);
or U2278 (N_2278,In_2079,In_2690);
nand U2279 (N_2279,In_259,In_2002);
and U2280 (N_2280,In_2753,In_657);
and U2281 (N_2281,In_2365,In_1342);
nor U2282 (N_2282,In_2671,In_1950);
nor U2283 (N_2283,In_2534,In_1137);
nor U2284 (N_2284,In_417,In_122);
or U2285 (N_2285,In_427,In_1336);
nor U2286 (N_2286,In_1805,In_1875);
nor U2287 (N_2287,In_248,In_2076);
nand U2288 (N_2288,In_67,In_1218);
and U2289 (N_2289,In_2866,In_230);
nor U2290 (N_2290,In_826,In_2815);
and U2291 (N_2291,In_1638,In_2277);
nor U2292 (N_2292,In_1799,In_799);
xor U2293 (N_2293,In_2070,In_2865);
or U2294 (N_2294,In_1806,In_133);
nor U2295 (N_2295,In_117,In_2348);
and U2296 (N_2296,In_2949,In_420);
nor U2297 (N_2297,In_19,In_541);
and U2298 (N_2298,In_1628,In_490);
xnor U2299 (N_2299,In_1491,In_1839);
and U2300 (N_2300,In_2282,In_2243);
or U2301 (N_2301,In_2816,In_2194);
nand U2302 (N_2302,In_1428,In_1478);
or U2303 (N_2303,In_601,In_2688);
nor U2304 (N_2304,In_1082,In_1566);
nor U2305 (N_2305,In_1519,In_622);
or U2306 (N_2306,In_716,In_1655);
nand U2307 (N_2307,In_495,In_193);
and U2308 (N_2308,In_166,In_2550);
and U2309 (N_2309,In_1755,In_2302);
nand U2310 (N_2310,In_1031,In_2707);
nor U2311 (N_2311,In_492,In_1480);
nor U2312 (N_2312,In_580,In_2717);
and U2313 (N_2313,In_2815,In_2293);
nand U2314 (N_2314,In_428,In_2142);
xnor U2315 (N_2315,In_1787,In_2355);
nor U2316 (N_2316,In_2648,In_885);
nor U2317 (N_2317,In_826,In_911);
and U2318 (N_2318,In_281,In_231);
xnor U2319 (N_2319,In_398,In_1933);
and U2320 (N_2320,In_1621,In_2146);
xnor U2321 (N_2321,In_1591,In_102);
nand U2322 (N_2322,In_187,In_279);
or U2323 (N_2323,In_873,In_722);
nand U2324 (N_2324,In_1465,In_2972);
nor U2325 (N_2325,In_1149,In_1894);
nand U2326 (N_2326,In_2950,In_1850);
xnor U2327 (N_2327,In_367,In_2515);
or U2328 (N_2328,In_1732,In_343);
nor U2329 (N_2329,In_2763,In_2416);
xnor U2330 (N_2330,In_1758,In_470);
xnor U2331 (N_2331,In_96,In_1687);
nand U2332 (N_2332,In_475,In_881);
xnor U2333 (N_2333,In_2418,In_467);
nand U2334 (N_2334,In_1,In_1095);
and U2335 (N_2335,In_1766,In_1832);
nand U2336 (N_2336,In_2884,In_2568);
nand U2337 (N_2337,In_899,In_2080);
or U2338 (N_2338,In_2273,In_1049);
nor U2339 (N_2339,In_2212,In_2741);
and U2340 (N_2340,In_2539,In_114);
and U2341 (N_2341,In_2337,In_567);
or U2342 (N_2342,In_144,In_745);
or U2343 (N_2343,In_2781,In_629);
nor U2344 (N_2344,In_408,In_1100);
xnor U2345 (N_2345,In_149,In_1016);
xnor U2346 (N_2346,In_75,In_90);
nor U2347 (N_2347,In_289,In_2069);
nand U2348 (N_2348,In_75,In_2289);
nor U2349 (N_2349,In_1185,In_1888);
or U2350 (N_2350,In_1647,In_1414);
or U2351 (N_2351,In_2187,In_217);
xnor U2352 (N_2352,In_1010,In_2576);
nor U2353 (N_2353,In_1070,In_580);
or U2354 (N_2354,In_610,In_2882);
nand U2355 (N_2355,In_452,In_729);
xnor U2356 (N_2356,In_2471,In_1322);
and U2357 (N_2357,In_243,In_866);
xor U2358 (N_2358,In_36,In_2385);
and U2359 (N_2359,In_2306,In_2851);
nor U2360 (N_2360,In_1825,In_889);
or U2361 (N_2361,In_1710,In_962);
xor U2362 (N_2362,In_928,In_1060);
and U2363 (N_2363,In_1439,In_2012);
xnor U2364 (N_2364,In_1213,In_1441);
nor U2365 (N_2365,In_1252,In_336);
xor U2366 (N_2366,In_2082,In_2541);
xor U2367 (N_2367,In_1459,In_2710);
nand U2368 (N_2368,In_2028,In_908);
and U2369 (N_2369,In_2924,In_561);
nand U2370 (N_2370,In_195,In_2080);
xor U2371 (N_2371,In_1178,In_2617);
nand U2372 (N_2372,In_691,In_867);
xnor U2373 (N_2373,In_370,In_2465);
or U2374 (N_2374,In_1558,In_1188);
and U2375 (N_2375,In_1147,In_2181);
nor U2376 (N_2376,In_2640,In_1932);
nor U2377 (N_2377,In_515,In_646);
nand U2378 (N_2378,In_1025,In_2369);
or U2379 (N_2379,In_989,In_2737);
nor U2380 (N_2380,In_1206,In_2943);
xor U2381 (N_2381,In_2535,In_429);
and U2382 (N_2382,In_1143,In_1271);
and U2383 (N_2383,In_2074,In_1510);
nor U2384 (N_2384,In_2667,In_1940);
nor U2385 (N_2385,In_1036,In_1620);
nor U2386 (N_2386,In_438,In_631);
and U2387 (N_2387,In_2038,In_2957);
or U2388 (N_2388,In_2418,In_2913);
nor U2389 (N_2389,In_2343,In_1692);
nand U2390 (N_2390,In_2952,In_2456);
xor U2391 (N_2391,In_1892,In_781);
or U2392 (N_2392,In_1057,In_1520);
and U2393 (N_2393,In_1637,In_802);
nand U2394 (N_2394,In_2993,In_625);
or U2395 (N_2395,In_2503,In_961);
or U2396 (N_2396,In_640,In_1244);
xnor U2397 (N_2397,In_2575,In_2648);
nor U2398 (N_2398,In_1641,In_1058);
and U2399 (N_2399,In_1846,In_2627);
nor U2400 (N_2400,In_773,In_302);
xor U2401 (N_2401,In_335,In_73);
and U2402 (N_2402,In_48,In_317);
nand U2403 (N_2403,In_645,In_2502);
nor U2404 (N_2404,In_2670,In_2653);
nand U2405 (N_2405,In_45,In_2803);
nand U2406 (N_2406,In_25,In_1173);
nor U2407 (N_2407,In_1271,In_562);
xor U2408 (N_2408,In_208,In_330);
or U2409 (N_2409,In_83,In_1108);
xor U2410 (N_2410,In_1250,In_2312);
and U2411 (N_2411,In_1252,In_2122);
or U2412 (N_2412,In_1650,In_2102);
or U2413 (N_2413,In_2961,In_891);
nand U2414 (N_2414,In_770,In_1835);
and U2415 (N_2415,In_1505,In_1936);
xnor U2416 (N_2416,In_2048,In_36);
nor U2417 (N_2417,In_601,In_1632);
nor U2418 (N_2418,In_1223,In_1708);
and U2419 (N_2419,In_2098,In_1089);
and U2420 (N_2420,In_1805,In_2015);
nand U2421 (N_2421,In_865,In_570);
xor U2422 (N_2422,In_147,In_893);
or U2423 (N_2423,In_2998,In_2273);
xor U2424 (N_2424,In_648,In_97);
nor U2425 (N_2425,In_2031,In_2174);
and U2426 (N_2426,In_1196,In_2651);
nor U2427 (N_2427,In_39,In_2485);
and U2428 (N_2428,In_1189,In_484);
nand U2429 (N_2429,In_1555,In_2687);
nand U2430 (N_2430,In_441,In_2450);
xor U2431 (N_2431,In_2926,In_1645);
nor U2432 (N_2432,In_1620,In_2856);
nor U2433 (N_2433,In_915,In_2764);
nor U2434 (N_2434,In_2797,In_638);
and U2435 (N_2435,In_933,In_1621);
nand U2436 (N_2436,In_1281,In_1079);
nand U2437 (N_2437,In_1296,In_1683);
nor U2438 (N_2438,In_2628,In_138);
or U2439 (N_2439,In_1288,In_1129);
or U2440 (N_2440,In_1814,In_1359);
xor U2441 (N_2441,In_1375,In_512);
or U2442 (N_2442,In_2410,In_1582);
nand U2443 (N_2443,In_2697,In_285);
or U2444 (N_2444,In_781,In_1161);
nand U2445 (N_2445,In_2072,In_833);
xnor U2446 (N_2446,In_189,In_1013);
nor U2447 (N_2447,In_1007,In_2157);
or U2448 (N_2448,In_402,In_1182);
and U2449 (N_2449,In_1327,In_737);
or U2450 (N_2450,In_310,In_51);
nor U2451 (N_2451,In_1817,In_2552);
xor U2452 (N_2452,In_2144,In_972);
and U2453 (N_2453,In_1712,In_2479);
xor U2454 (N_2454,In_2303,In_1803);
nor U2455 (N_2455,In_2998,In_350);
xor U2456 (N_2456,In_984,In_1017);
nand U2457 (N_2457,In_2862,In_531);
nand U2458 (N_2458,In_1966,In_1818);
xor U2459 (N_2459,In_2855,In_1737);
or U2460 (N_2460,In_2412,In_890);
nand U2461 (N_2461,In_654,In_174);
nor U2462 (N_2462,In_2885,In_1489);
nor U2463 (N_2463,In_1639,In_2058);
nand U2464 (N_2464,In_41,In_1780);
xnor U2465 (N_2465,In_2524,In_1840);
nand U2466 (N_2466,In_520,In_2603);
and U2467 (N_2467,In_1329,In_1500);
xor U2468 (N_2468,In_2929,In_543);
xnor U2469 (N_2469,In_850,In_1580);
xnor U2470 (N_2470,In_1610,In_1372);
xor U2471 (N_2471,In_1434,In_622);
nand U2472 (N_2472,In_54,In_2243);
nor U2473 (N_2473,In_2706,In_467);
or U2474 (N_2474,In_2391,In_1723);
and U2475 (N_2475,In_1703,In_468);
xor U2476 (N_2476,In_720,In_2804);
xnor U2477 (N_2477,In_484,In_146);
and U2478 (N_2478,In_1260,In_699);
and U2479 (N_2479,In_2865,In_2129);
nand U2480 (N_2480,In_648,In_2419);
nand U2481 (N_2481,In_752,In_2137);
or U2482 (N_2482,In_2590,In_1639);
nand U2483 (N_2483,In_1149,In_622);
nor U2484 (N_2484,In_344,In_1394);
and U2485 (N_2485,In_2850,In_1508);
and U2486 (N_2486,In_174,In_71);
or U2487 (N_2487,In_617,In_1446);
nand U2488 (N_2488,In_2889,In_173);
xnor U2489 (N_2489,In_903,In_2494);
nor U2490 (N_2490,In_1930,In_1568);
nor U2491 (N_2491,In_231,In_2147);
xnor U2492 (N_2492,In_526,In_1279);
nand U2493 (N_2493,In_745,In_2997);
nand U2494 (N_2494,In_2891,In_2832);
nand U2495 (N_2495,In_1946,In_2785);
xor U2496 (N_2496,In_1302,In_2275);
xnor U2497 (N_2497,In_1725,In_2718);
nand U2498 (N_2498,In_2360,In_687);
or U2499 (N_2499,In_2904,In_1481);
or U2500 (N_2500,In_1760,In_493);
nor U2501 (N_2501,In_580,In_2312);
or U2502 (N_2502,In_1877,In_1920);
or U2503 (N_2503,In_1282,In_1851);
nor U2504 (N_2504,In_44,In_2144);
and U2505 (N_2505,In_1043,In_2484);
nor U2506 (N_2506,In_1276,In_913);
or U2507 (N_2507,In_2438,In_1134);
nor U2508 (N_2508,In_287,In_2376);
nand U2509 (N_2509,In_2924,In_882);
or U2510 (N_2510,In_2974,In_77);
nand U2511 (N_2511,In_2328,In_2398);
or U2512 (N_2512,In_566,In_2720);
nor U2513 (N_2513,In_472,In_1499);
and U2514 (N_2514,In_1443,In_851);
xnor U2515 (N_2515,In_1924,In_81);
nand U2516 (N_2516,In_203,In_1582);
nor U2517 (N_2517,In_1550,In_955);
and U2518 (N_2518,In_874,In_2767);
xor U2519 (N_2519,In_553,In_1511);
nand U2520 (N_2520,In_2198,In_2);
nor U2521 (N_2521,In_2786,In_1376);
nand U2522 (N_2522,In_1521,In_2689);
nor U2523 (N_2523,In_2798,In_1575);
nor U2524 (N_2524,In_1305,In_335);
nor U2525 (N_2525,In_773,In_126);
or U2526 (N_2526,In_1213,In_2406);
xnor U2527 (N_2527,In_766,In_826);
nand U2528 (N_2528,In_1708,In_2153);
nor U2529 (N_2529,In_321,In_1871);
and U2530 (N_2530,In_651,In_1446);
xor U2531 (N_2531,In_2973,In_1749);
and U2532 (N_2532,In_502,In_256);
and U2533 (N_2533,In_2353,In_1059);
xor U2534 (N_2534,In_934,In_1061);
and U2535 (N_2535,In_1508,In_809);
or U2536 (N_2536,In_2373,In_1993);
or U2537 (N_2537,In_768,In_541);
nor U2538 (N_2538,In_2163,In_2139);
and U2539 (N_2539,In_809,In_2643);
nor U2540 (N_2540,In_1128,In_2691);
and U2541 (N_2541,In_872,In_2512);
nand U2542 (N_2542,In_1723,In_2318);
and U2543 (N_2543,In_593,In_2143);
and U2544 (N_2544,In_2182,In_1130);
xor U2545 (N_2545,In_586,In_1131);
xnor U2546 (N_2546,In_191,In_462);
nand U2547 (N_2547,In_763,In_1555);
and U2548 (N_2548,In_2349,In_1809);
or U2549 (N_2549,In_310,In_707);
or U2550 (N_2550,In_1105,In_2507);
xor U2551 (N_2551,In_284,In_1768);
xor U2552 (N_2552,In_1949,In_2277);
nand U2553 (N_2553,In_421,In_602);
or U2554 (N_2554,In_325,In_1428);
nor U2555 (N_2555,In_564,In_1917);
nor U2556 (N_2556,In_2556,In_831);
and U2557 (N_2557,In_913,In_1227);
nor U2558 (N_2558,In_640,In_1970);
or U2559 (N_2559,In_2379,In_111);
and U2560 (N_2560,In_471,In_448);
nor U2561 (N_2561,In_640,In_700);
xor U2562 (N_2562,In_614,In_2637);
and U2563 (N_2563,In_1146,In_593);
xor U2564 (N_2564,In_2194,In_2006);
nor U2565 (N_2565,In_703,In_1558);
and U2566 (N_2566,In_2204,In_465);
nand U2567 (N_2567,In_216,In_678);
or U2568 (N_2568,In_2568,In_2520);
xnor U2569 (N_2569,In_2982,In_2856);
or U2570 (N_2570,In_829,In_1412);
or U2571 (N_2571,In_1351,In_2326);
nor U2572 (N_2572,In_715,In_1469);
nor U2573 (N_2573,In_1285,In_2235);
nand U2574 (N_2574,In_2403,In_1533);
or U2575 (N_2575,In_1484,In_1773);
or U2576 (N_2576,In_1555,In_2268);
xor U2577 (N_2577,In_2271,In_683);
or U2578 (N_2578,In_854,In_2452);
xnor U2579 (N_2579,In_332,In_1919);
and U2580 (N_2580,In_2383,In_676);
nor U2581 (N_2581,In_1204,In_115);
nor U2582 (N_2582,In_212,In_1550);
and U2583 (N_2583,In_2951,In_1303);
xnor U2584 (N_2584,In_1438,In_74);
xnor U2585 (N_2585,In_2206,In_1086);
and U2586 (N_2586,In_2332,In_1544);
and U2587 (N_2587,In_2836,In_1830);
xnor U2588 (N_2588,In_59,In_999);
nand U2589 (N_2589,In_2027,In_1003);
and U2590 (N_2590,In_1179,In_435);
nor U2591 (N_2591,In_2623,In_519);
nand U2592 (N_2592,In_2817,In_962);
or U2593 (N_2593,In_1504,In_2700);
or U2594 (N_2594,In_2876,In_843);
or U2595 (N_2595,In_500,In_2130);
nand U2596 (N_2596,In_2666,In_660);
or U2597 (N_2597,In_1511,In_1282);
and U2598 (N_2598,In_1904,In_2232);
nor U2599 (N_2599,In_156,In_946);
and U2600 (N_2600,In_2280,In_596);
nand U2601 (N_2601,In_2051,In_2140);
and U2602 (N_2602,In_2350,In_1557);
nand U2603 (N_2603,In_1674,In_1367);
and U2604 (N_2604,In_1309,In_2779);
and U2605 (N_2605,In_267,In_2280);
or U2606 (N_2606,In_2002,In_1981);
nor U2607 (N_2607,In_989,In_905);
and U2608 (N_2608,In_1487,In_1205);
and U2609 (N_2609,In_2034,In_2012);
nor U2610 (N_2610,In_2592,In_693);
or U2611 (N_2611,In_1450,In_216);
or U2612 (N_2612,In_1076,In_1708);
nor U2613 (N_2613,In_2624,In_1885);
nand U2614 (N_2614,In_1459,In_1360);
nand U2615 (N_2615,In_389,In_1005);
and U2616 (N_2616,In_1966,In_2838);
and U2617 (N_2617,In_1364,In_2811);
xnor U2618 (N_2618,In_1675,In_2232);
nor U2619 (N_2619,In_2020,In_1575);
or U2620 (N_2620,In_1716,In_1158);
and U2621 (N_2621,In_2515,In_985);
and U2622 (N_2622,In_2081,In_178);
xor U2623 (N_2623,In_337,In_2173);
nor U2624 (N_2624,In_964,In_2038);
and U2625 (N_2625,In_2826,In_801);
nor U2626 (N_2626,In_2960,In_275);
nand U2627 (N_2627,In_630,In_1595);
or U2628 (N_2628,In_2474,In_2897);
and U2629 (N_2629,In_2984,In_783);
and U2630 (N_2630,In_1040,In_5);
and U2631 (N_2631,In_988,In_35);
nand U2632 (N_2632,In_1391,In_1691);
nand U2633 (N_2633,In_271,In_2706);
nand U2634 (N_2634,In_2848,In_1037);
and U2635 (N_2635,In_1931,In_2493);
xor U2636 (N_2636,In_1861,In_129);
nor U2637 (N_2637,In_2807,In_1813);
and U2638 (N_2638,In_1899,In_1393);
nand U2639 (N_2639,In_992,In_1632);
nand U2640 (N_2640,In_700,In_626);
xnor U2641 (N_2641,In_352,In_2910);
nand U2642 (N_2642,In_537,In_309);
xnor U2643 (N_2643,In_670,In_1363);
and U2644 (N_2644,In_1370,In_357);
or U2645 (N_2645,In_2082,In_2822);
and U2646 (N_2646,In_2607,In_2391);
or U2647 (N_2647,In_2334,In_85);
nor U2648 (N_2648,In_1738,In_1965);
nand U2649 (N_2649,In_2025,In_1319);
nor U2650 (N_2650,In_2611,In_495);
nand U2651 (N_2651,In_2941,In_1658);
and U2652 (N_2652,In_1362,In_2360);
nand U2653 (N_2653,In_1033,In_1912);
nand U2654 (N_2654,In_659,In_23);
nor U2655 (N_2655,In_2009,In_513);
and U2656 (N_2656,In_2892,In_2335);
nor U2657 (N_2657,In_210,In_2394);
xor U2658 (N_2658,In_2436,In_676);
or U2659 (N_2659,In_545,In_540);
and U2660 (N_2660,In_1346,In_1027);
nand U2661 (N_2661,In_1137,In_71);
xor U2662 (N_2662,In_1824,In_870);
or U2663 (N_2663,In_2293,In_1581);
nor U2664 (N_2664,In_1542,In_2445);
or U2665 (N_2665,In_2922,In_345);
and U2666 (N_2666,In_2482,In_1505);
or U2667 (N_2667,In_276,In_561);
nor U2668 (N_2668,In_1411,In_2784);
nand U2669 (N_2669,In_1803,In_1819);
nand U2670 (N_2670,In_912,In_2245);
or U2671 (N_2671,In_255,In_1361);
xnor U2672 (N_2672,In_671,In_157);
or U2673 (N_2673,In_1484,In_2245);
xnor U2674 (N_2674,In_633,In_1620);
nand U2675 (N_2675,In_2803,In_932);
nor U2676 (N_2676,In_218,In_395);
and U2677 (N_2677,In_2050,In_2738);
and U2678 (N_2678,In_2478,In_2674);
xor U2679 (N_2679,In_1036,In_2743);
nand U2680 (N_2680,In_1094,In_1615);
nand U2681 (N_2681,In_1000,In_448);
or U2682 (N_2682,In_1159,In_134);
xnor U2683 (N_2683,In_1724,In_2892);
nor U2684 (N_2684,In_2034,In_1201);
xnor U2685 (N_2685,In_2499,In_314);
and U2686 (N_2686,In_15,In_200);
xnor U2687 (N_2687,In_12,In_542);
or U2688 (N_2688,In_2874,In_1282);
xnor U2689 (N_2689,In_1824,In_2334);
xor U2690 (N_2690,In_624,In_993);
xor U2691 (N_2691,In_719,In_1849);
and U2692 (N_2692,In_1873,In_1688);
and U2693 (N_2693,In_243,In_1773);
nor U2694 (N_2694,In_1062,In_2787);
nor U2695 (N_2695,In_2256,In_1636);
nand U2696 (N_2696,In_1444,In_1490);
or U2697 (N_2697,In_1059,In_1813);
xor U2698 (N_2698,In_1050,In_1114);
nor U2699 (N_2699,In_418,In_1089);
and U2700 (N_2700,In_38,In_1709);
and U2701 (N_2701,In_1883,In_2741);
nor U2702 (N_2702,In_1101,In_1722);
nor U2703 (N_2703,In_2677,In_2622);
and U2704 (N_2704,In_1953,In_2158);
xnor U2705 (N_2705,In_819,In_1382);
or U2706 (N_2706,In_1198,In_1093);
and U2707 (N_2707,In_363,In_2782);
or U2708 (N_2708,In_2409,In_2255);
or U2709 (N_2709,In_1283,In_1325);
nor U2710 (N_2710,In_2986,In_1777);
and U2711 (N_2711,In_2148,In_1775);
nand U2712 (N_2712,In_2548,In_1285);
xor U2713 (N_2713,In_1619,In_1234);
nand U2714 (N_2714,In_291,In_53);
and U2715 (N_2715,In_607,In_1270);
nand U2716 (N_2716,In_2500,In_96);
and U2717 (N_2717,In_176,In_744);
nor U2718 (N_2718,In_47,In_436);
or U2719 (N_2719,In_1763,In_2089);
nor U2720 (N_2720,In_1236,In_555);
xnor U2721 (N_2721,In_209,In_1907);
nor U2722 (N_2722,In_2197,In_1652);
nand U2723 (N_2723,In_2588,In_2029);
xnor U2724 (N_2724,In_2683,In_1579);
or U2725 (N_2725,In_2552,In_1836);
nor U2726 (N_2726,In_2744,In_103);
xor U2727 (N_2727,In_1227,In_2936);
xnor U2728 (N_2728,In_485,In_314);
xor U2729 (N_2729,In_1159,In_1337);
xor U2730 (N_2730,In_1134,In_82);
and U2731 (N_2731,In_2091,In_2584);
and U2732 (N_2732,In_1694,In_350);
nand U2733 (N_2733,In_1205,In_1166);
nor U2734 (N_2734,In_2771,In_2051);
or U2735 (N_2735,In_2493,In_1774);
or U2736 (N_2736,In_117,In_2297);
xnor U2737 (N_2737,In_1782,In_2234);
nand U2738 (N_2738,In_2428,In_1626);
and U2739 (N_2739,In_557,In_2171);
nand U2740 (N_2740,In_795,In_821);
nor U2741 (N_2741,In_376,In_1283);
and U2742 (N_2742,In_1819,In_375);
nor U2743 (N_2743,In_1869,In_1175);
xor U2744 (N_2744,In_261,In_2863);
or U2745 (N_2745,In_1535,In_2616);
xor U2746 (N_2746,In_2475,In_2664);
nand U2747 (N_2747,In_2262,In_42);
and U2748 (N_2748,In_631,In_1710);
nor U2749 (N_2749,In_183,In_1062);
or U2750 (N_2750,In_2668,In_1355);
nor U2751 (N_2751,In_1554,In_701);
and U2752 (N_2752,In_2489,In_2705);
xor U2753 (N_2753,In_1216,In_1162);
or U2754 (N_2754,In_2049,In_1234);
and U2755 (N_2755,In_2048,In_2929);
xor U2756 (N_2756,In_2976,In_1277);
or U2757 (N_2757,In_2729,In_431);
nor U2758 (N_2758,In_2577,In_2299);
nand U2759 (N_2759,In_428,In_1875);
nor U2760 (N_2760,In_255,In_2914);
and U2761 (N_2761,In_2984,In_1787);
nor U2762 (N_2762,In_569,In_1916);
nand U2763 (N_2763,In_733,In_2553);
and U2764 (N_2764,In_2907,In_2786);
or U2765 (N_2765,In_2499,In_1641);
and U2766 (N_2766,In_2029,In_2753);
nand U2767 (N_2767,In_451,In_1451);
nor U2768 (N_2768,In_2977,In_129);
nor U2769 (N_2769,In_2016,In_2874);
and U2770 (N_2770,In_1148,In_1971);
nor U2771 (N_2771,In_1032,In_1889);
nand U2772 (N_2772,In_692,In_1631);
nand U2773 (N_2773,In_2050,In_2170);
xor U2774 (N_2774,In_732,In_401);
nor U2775 (N_2775,In_2343,In_529);
and U2776 (N_2776,In_2136,In_1160);
nor U2777 (N_2777,In_1759,In_1140);
xor U2778 (N_2778,In_2539,In_614);
nor U2779 (N_2779,In_2805,In_2680);
nand U2780 (N_2780,In_1255,In_2070);
and U2781 (N_2781,In_920,In_287);
or U2782 (N_2782,In_1491,In_2932);
and U2783 (N_2783,In_2046,In_930);
or U2784 (N_2784,In_2480,In_2306);
xnor U2785 (N_2785,In_172,In_732);
nand U2786 (N_2786,In_1320,In_1619);
or U2787 (N_2787,In_2164,In_1914);
and U2788 (N_2788,In_82,In_1289);
nor U2789 (N_2789,In_2626,In_1398);
xor U2790 (N_2790,In_957,In_2312);
nor U2791 (N_2791,In_2237,In_2786);
xnor U2792 (N_2792,In_1251,In_2373);
xor U2793 (N_2793,In_1404,In_2789);
xor U2794 (N_2794,In_2749,In_437);
xnor U2795 (N_2795,In_71,In_297);
or U2796 (N_2796,In_247,In_2038);
and U2797 (N_2797,In_1125,In_2746);
xor U2798 (N_2798,In_1924,In_1279);
xor U2799 (N_2799,In_2192,In_242);
or U2800 (N_2800,In_1202,In_488);
nand U2801 (N_2801,In_1379,In_1875);
and U2802 (N_2802,In_1156,In_13);
nor U2803 (N_2803,In_20,In_2415);
nand U2804 (N_2804,In_407,In_658);
nand U2805 (N_2805,In_1745,In_1811);
nor U2806 (N_2806,In_2881,In_2232);
nor U2807 (N_2807,In_2177,In_2725);
xnor U2808 (N_2808,In_816,In_192);
nor U2809 (N_2809,In_1501,In_2126);
and U2810 (N_2810,In_528,In_1474);
and U2811 (N_2811,In_576,In_288);
or U2812 (N_2812,In_1142,In_1562);
or U2813 (N_2813,In_2886,In_1315);
xor U2814 (N_2814,In_1493,In_551);
and U2815 (N_2815,In_2176,In_2597);
or U2816 (N_2816,In_1656,In_1293);
nand U2817 (N_2817,In_727,In_490);
or U2818 (N_2818,In_1469,In_1335);
or U2819 (N_2819,In_1,In_2236);
or U2820 (N_2820,In_990,In_1111);
xor U2821 (N_2821,In_278,In_1751);
and U2822 (N_2822,In_2962,In_132);
and U2823 (N_2823,In_2896,In_501);
and U2824 (N_2824,In_2944,In_160);
and U2825 (N_2825,In_2111,In_1245);
and U2826 (N_2826,In_674,In_1937);
and U2827 (N_2827,In_1059,In_2496);
and U2828 (N_2828,In_2841,In_705);
nor U2829 (N_2829,In_1116,In_1264);
or U2830 (N_2830,In_1105,In_422);
and U2831 (N_2831,In_1555,In_1757);
and U2832 (N_2832,In_278,In_2107);
or U2833 (N_2833,In_1227,In_2393);
nor U2834 (N_2834,In_2097,In_2030);
and U2835 (N_2835,In_2903,In_925);
nand U2836 (N_2836,In_103,In_1484);
nor U2837 (N_2837,In_1346,In_2152);
nor U2838 (N_2838,In_1326,In_1839);
xor U2839 (N_2839,In_2224,In_1159);
xnor U2840 (N_2840,In_1014,In_1890);
or U2841 (N_2841,In_2002,In_2346);
nand U2842 (N_2842,In_1208,In_1640);
and U2843 (N_2843,In_2878,In_258);
nor U2844 (N_2844,In_607,In_2679);
xor U2845 (N_2845,In_383,In_229);
nor U2846 (N_2846,In_2959,In_544);
xnor U2847 (N_2847,In_1200,In_1825);
or U2848 (N_2848,In_1179,In_1111);
xnor U2849 (N_2849,In_2063,In_717);
or U2850 (N_2850,In_2649,In_1803);
or U2851 (N_2851,In_2359,In_1989);
or U2852 (N_2852,In_1580,In_2275);
nor U2853 (N_2853,In_2920,In_699);
xnor U2854 (N_2854,In_153,In_1560);
nand U2855 (N_2855,In_2186,In_2990);
xnor U2856 (N_2856,In_1426,In_2604);
nand U2857 (N_2857,In_727,In_2031);
and U2858 (N_2858,In_595,In_1864);
or U2859 (N_2859,In_2827,In_799);
nor U2860 (N_2860,In_2593,In_1606);
nor U2861 (N_2861,In_1050,In_944);
or U2862 (N_2862,In_148,In_796);
and U2863 (N_2863,In_1265,In_2534);
nor U2864 (N_2864,In_1798,In_1219);
or U2865 (N_2865,In_360,In_878);
nand U2866 (N_2866,In_984,In_485);
xnor U2867 (N_2867,In_1955,In_1997);
nor U2868 (N_2868,In_2637,In_520);
or U2869 (N_2869,In_2294,In_1728);
and U2870 (N_2870,In_2096,In_102);
and U2871 (N_2871,In_2511,In_1206);
and U2872 (N_2872,In_760,In_2565);
or U2873 (N_2873,In_2861,In_1590);
nand U2874 (N_2874,In_1731,In_1050);
nand U2875 (N_2875,In_1182,In_1714);
nand U2876 (N_2876,In_711,In_1030);
or U2877 (N_2877,In_2956,In_306);
nand U2878 (N_2878,In_2458,In_2643);
nand U2879 (N_2879,In_1071,In_1020);
or U2880 (N_2880,In_1255,In_1513);
nor U2881 (N_2881,In_2806,In_2314);
or U2882 (N_2882,In_2546,In_1881);
nand U2883 (N_2883,In_2671,In_2898);
and U2884 (N_2884,In_2532,In_1979);
nor U2885 (N_2885,In_1387,In_1606);
nor U2886 (N_2886,In_694,In_1551);
and U2887 (N_2887,In_1690,In_2496);
and U2888 (N_2888,In_1032,In_1755);
nand U2889 (N_2889,In_1712,In_1851);
or U2890 (N_2890,In_1391,In_1633);
or U2891 (N_2891,In_1008,In_556);
or U2892 (N_2892,In_1751,In_789);
nor U2893 (N_2893,In_2292,In_683);
nor U2894 (N_2894,In_2792,In_1945);
xnor U2895 (N_2895,In_758,In_1045);
or U2896 (N_2896,In_2868,In_472);
nand U2897 (N_2897,In_2370,In_341);
xnor U2898 (N_2898,In_1333,In_217);
nand U2899 (N_2899,In_2647,In_2839);
or U2900 (N_2900,In_1604,In_508);
or U2901 (N_2901,In_1190,In_1466);
xnor U2902 (N_2902,In_83,In_2418);
xnor U2903 (N_2903,In_2186,In_365);
or U2904 (N_2904,In_949,In_39);
or U2905 (N_2905,In_1386,In_2468);
and U2906 (N_2906,In_248,In_1379);
nand U2907 (N_2907,In_136,In_2763);
and U2908 (N_2908,In_1907,In_2279);
nand U2909 (N_2909,In_1280,In_106);
nand U2910 (N_2910,In_1437,In_1479);
nor U2911 (N_2911,In_1696,In_1458);
xor U2912 (N_2912,In_1398,In_2297);
nor U2913 (N_2913,In_1410,In_1876);
nor U2914 (N_2914,In_2401,In_245);
or U2915 (N_2915,In_2787,In_1178);
nor U2916 (N_2916,In_1531,In_1628);
nor U2917 (N_2917,In_2413,In_2697);
and U2918 (N_2918,In_2876,In_579);
nor U2919 (N_2919,In_952,In_1819);
or U2920 (N_2920,In_2294,In_1990);
nand U2921 (N_2921,In_2100,In_1639);
xor U2922 (N_2922,In_648,In_1644);
xnor U2923 (N_2923,In_564,In_2563);
nand U2924 (N_2924,In_1004,In_2045);
nand U2925 (N_2925,In_464,In_575);
and U2926 (N_2926,In_516,In_1388);
or U2927 (N_2927,In_99,In_1336);
xnor U2928 (N_2928,In_2178,In_2661);
nor U2929 (N_2929,In_86,In_1935);
xnor U2930 (N_2930,In_1487,In_2066);
or U2931 (N_2931,In_1427,In_1929);
or U2932 (N_2932,In_322,In_2316);
or U2933 (N_2933,In_2451,In_547);
or U2934 (N_2934,In_975,In_2428);
or U2935 (N_2935,In_2128,In_2046);
or U2936 (N_2936,In_2431,In_703);
nand U2937 (N_2937,In_122,In_1660);
xor U2938 (N_2938,In_2923,In_188);
nand U2939 (N_2939,In_158,In_2931);
nand U2940 (N_2940,In_1185,In_1942);
nor U2941 (N_2941,In_69,In_1183);
xor U2942 (N_2942,In_2221,In_1617);
or U2943 (N_2943,In_588,In_406);
and U2944 (N_2944,In_789,In_2937);
and U2945 (N_2945,In_2201,In_2981);
xor U2946 (N_2946,In_2814,In_1755);
or U2947 (N_2947,In_2547,In_1447);
or U2948 (N_2948,In_1263,In_678);
and U2949 (N_2949,In_927,In_557);
and U2950 (N_2950,In_81,In_1343);
xor U2951 (N_2951,In_1657,In_817);
nor U2952 (N_2952,In_2766,In_1821);
nand U2953 (N_2953,In_185,In_2910);
or U2954 (N_2954,In_2829,In_934);
xor U2955 (N_2955,In_1949,In_877);
and U2956 (N_2956,In_1251,In_2113);
nor U2957 (N_2957,In_439,In_309);
nand U2958 (N_2958,In_2580,In_1160);
and U2959 (N_2959,In_1544,In_2174);
nor U2960 (N_2960,In_1427,In_2105);
nand U2961 (N_2961,In_1195,In_1817);
or U2962 (N_2962,In_818,In_1003);
nor U2963 (N_2963,In_1934,In_2251);
and U2964 (N_2964,In_723,In_2675);
xor U2965 (N_2965,In_57,In_2435);
nand U2966 (N_2966,In_1846,In_1543);
nand U2967 (N_2967,In_686,In_660);
and U2968 (N_2968,In_675,In_2889);
and U2969 (N_2969,In_2445,In_2421);
xor U2970 (N_2970,In_833,In_2560);
nand U2971 (N_2971,In_1847,In_1168);
or U2972 (N_2972,In_2704,In_1196);
nor U2973 (N_2973,In_826,In_2612);
nor U2974 (N_2974,In_1825,In_2124);
xnor U2975 (N_2975,In_1147,In_149);
or U2976 (N_2976,In_2595,In_581);
or U2977 (N_2977,In_1080,In_404);
xnor U2978 (N_2978,In_2578,In_516);
and U2979 (N_2979,In_702,In_1773);
and U2980 (N_2980,In_684,In_975);
xor U2981 (N_2981,In_1378,In_1482);
or U2982 (N_2982,In_216,In_2801);
and U2983 (N_2983,In_606,In_1348);
nor U2984 (N_2984,In_1081,In_763);
nor U2985 (N_2985,In_1938,In_1576);
xor U2986 (N_2986,In_1793,In_1972);
and U2987 (N_2987,In_375,In_1026);
nor U2988 (N_2988,In_1705,In_2022);
and U2989 (N_2989,In_1080,In_1035);
nand U2990 (N_2990,In_116,In_1500);
nand U2991 (N_2991,In_1724,In_2136);
nor U2992 (N_2992,In_1645,In_944);
xnor U2993 (N_2993,In_97,In_1136);
nor U2994 (N_2994,In_2718,In_1052);
or U2995 (N_2995,In_2066,In_2143);
xor U2996 (N_2996,In_1221,In_989);
and U2997 (N_2997,In_754,In_1231);
xnor U2998 (N_2998,In_1849,In_2421);
or U2999 (N_2999,In_1014,In_1153);
nand U3000 (N_3000,In_1976,In_2334);
or U3001 (N_3001,In_972,In_2345);
and U3002 (N_3002,In_303,In_2827);
and U3003 (N_3003,In_2045,In_2234);
xnor U3004 (N_3004,In_1245,In_2958);
or U3005 (N_3005,In_2654,In_1691);
or U3006 (N_3006,In_1309,In_2457);
xor U3007 (N_3007,In_2755,In_187);
and U3008 (N_3008,In_929,In_1525);
nand U3009 (N_3009,In_321,In_1130);
xor U3010 (N_3010,In_362,In_445);
or U3011 (N_3011,In_2461,In_2749);
or U3012 (N_3012,In_1185,In_113);
and U3013 (N_3013,In_1234,In_1872);
nor U3014 (N_3014,In_2267,In_2624);
or U3015 (N_3015,In_2726,In_601);
nor U3016 (N_3016,In_1060,In_2371);
and U3017 (N_3017,In_2049,In_1209);
xnor U3018 (N_3018,In_2572,In_1850);
and U3019 (N_3019,In_2244,In_366);
or U3020 (N_3020,In_2889,In_2143);
nor U3021 (N_3021,In_1205,In_1101);
xnor U3022 (N_3022,In_1283,In_2879);
or U3023 (N_3023,In_1058,In_2854);
xor U3024 (N_3024,In_185,In_971);
and U3025 (N_3025,In_459,In_2223);
nand U3026 (N_3026,In_2790,In_767);
nor U3027 (N_3027,In_2966,In_1312);
nand U3028 (N_3028,In_2476,In_2053);
xnor U3029 (N_3029,In_2207,In_2904);
nand U3030 (N_3030,In_39,In_226);
and U3031 (N_3031,In_17,In_1833);
nor U3032 (N_3032,In_549,In_1234);
or U3033 (N_3033,In_578,In_796);
and U3034 (N_3034,In_192,In_1459);
and U3035 (N_3035,In_1853,In_605);
xor U3036 (N_3036,In_14,In_871);
xor U3037 (N_3037,In_1654,In_1092);
nor U3038 (N_3038,In_1762,In_1860);
nor U3039 (N_3039,In_1591,In_2172);
or U3040 (N_3040,In_1991,In_1969);
and U3041 (N_3041,In_1112,In_2561);
and U3042 (N_3042,In_777,In_2241);
or U3043 (N_3043,In_2946,In_1202);
nor U3044 (N_3044,In_2385,In_2829);
and U3045 (N_3045,In_1800,In_57);
nand U3046 (N_3046,In_2667,In_2548);
xnor U3047 (N_3047,In_2036,In_2163);
xor U3048 (N_3048,In_779,In_336);
nand U3049 (N_3049,In_2629,In_2064);
nor U3050 (N_3050,In_2619,In_2571);
xnor U3051 (N_3051,In_59,In_717);
and U3052 (N_3052,In_2510,In_2399);
nand U3053 (N_3053,In_1504,In_2109);
and U3054 (N_3054,In_2924,In_14);
nand U3055 (N_3055,In_1984,In_2984);
and U3056 (N_3056,In_1343,In_758);
or U3057 (N_3057,In_955,In_1454);
nor U3058 (N_3058,In_2561,In_2875);
nand U3059 (N_3059,In_1710,In_2461);
nand U3060 (N_3060,In_1738,In_2258);
and U3061 (N_3061,In_2856,In_1152);
nor U3062 (N_3062,In_2827,In_1189);
and U3063 (N_3063,In_653,In_2044);
nor U3064 (N_3064,In_929,In_1532);
and U3065 (N_3065,In_2239,In_2150);
nand U3066 (N_3066,In_2468,In_450);
and U3067 (N_3067,In_2016,In_2866);
or U3068 (N_3068,In_2575,In_1616);
or U3069 (N_3069,In_1002,In_2676);
nand U3070 (N_3070,In_2661,In_2800);
or U3071 (N_3071,In_401,In_642);
and U3072 (N_3072,In_2666,In_2815);
nor U3073 (N_3073,In_354,In_2410);
and U3074 (N_3074,In_885,In_2020);
and U3075 (N_3075,In_794,In_2766);
and U3076 (N_3076,In_804,In_2981);
xor U3077 (N_3077,In_1333,In_459);
or U3078 (N_3078,In_2333,In_2340);
nor U3079 (N_3079,In_2531,In_905);
or U3080 (N_3080,In_2493,In_2083);
nor U3081 (N_3081,In_2502,In_2332);
and U3082 (N_3082,In_2590,In_431);
and U3083 (N_3083,In_491,In_2055);
nand U3084 (N_3084,In_1800,In_2118);
nor U3085 (N_3085,In_1788,In_465);
xor U3086 (N_3086,In_1312,In_2463);
xnor U3087 (N_3087,In_2850,In_1976);
and U3088 (N_3088,In_1119,In_2688);
nor U3089 (N_3089,In_2375,In_1145);
and U3090 (N_3090,In_2200,In_2518);
nand U3091 (N_3091,In_2081,In_359);
xor U3092 (N_3092,In_109,In_342);
or U3093 (N_3093,In_1736,In_1509);
nor U3094 (N_3094,In_654,In_1905);
and U3095 (N_3095,In_526,In_122);
xor U3096 (N_3096,In_616,In_291);
nand U3097 (N_3097,In_384,In_2574);
or U3098 (N_3098,In_1743,In_1362);
or U3099 (N_3099,In_611,In_1082);
nand U3100 (N_3100,In_2764,In_1165);
nand U3101 (N_3101,In_2322,In_1637);
nand U3102 (N_3102,In_1303,In_1087);
xor U3103 (N_3103,In_1666,In_625);
and U3104 (N_3104,In_2457,In_527);
nand U3105 (N_3105,In_522,In_1888);
xnor U3106 (N_3106,In_2146,In_2465);
and U3107 (N_3107,In_900,In_1741);
xnor U3108 (N_3108,In_1020,In_1614);
nand U3109 (N_3109,In_343,In_74);
nand U3110 (N_3110,In_600,In_29);
nand U3111 (N_3111,In_1246,In_2952);
or U3112 (N_3112,In_1614,In_429);
nor U3113 (N_3113,In_2433,In_2399);
or U3114 (N_3114,In_1883,In_1393);
xor U3115 (N_3115,In_2420,In_1865);
or U3116 (N_3116,In_1638,In_2917);
nor U3117 (N_3117,In_2459,In_1183);
or U3118 (N_3118,In_2154,In_747);
nor U3119 (N_3119,In_2437,In_2864);
nand U3120 (N_3120,In_2340,In_2745);
xor U3121 (N_3121,In_2398,In_2034);
or U3122 (N_3122,In_2344,In_305);
nor U3123 (N_3123,In_2685,In_767);
nand U3124 (N_3124,In_1662,In_2528);
and U3125 (N_3125,In_1710,In_440);
xor U3126 (N_3126,In_2620,In_889);
or U3127 (N_3127,In_1060,In_987);
nand U3128 (N_3128,In_2057,In_538);
or U3129 (N_3129,In_540,In_316);
xor U3130 (N_3130,In_120,In_1360);
nand U3131 (N_3131,In_1755,In_2656);
nand U3132 (N_3132,In_1228,In_666);
nor U3133 (N_3133,In_94,In_91);
and U3134 (N_3134,In_2905,In_1965);
or U3135 (N_3135,In_2309,In_1182);
nor U3136 (N_3136,In_581,In_2761);
nor U3137 (N_3137,In_2476,In_1078);
nor U3138 (N_3138,In_2630,In_1628);
or U3139 (N_3139,In_1222,In_2104);
nor U3140 (N_3140,In_1194,In_826);
or U3141 (N_3141,In_427,In_1726);
or U3142 (N_3142,In_2633,In_2372);
nand U3143 (N_3143,In_2378,In_1861);
xor U3144 (N_3144,In_1902,In_1824);
and U3145 (N_3145,In_73,In_2847);
xor U3146 (N_3146,In_2469,In_514);
xnor U3147 (N_3147,In_2853,In_2814);
nor U3148 (N_3148,In_916,In_78);
or U3149 (N_3149,In_2879,In_2350);
nor U3150 (N_3150,In_2595,In_1811);
xnor U3151 (N_3151,In_2290,In_356);
nor U3152 (N_3152,In_2647,In_2623);
nand U3153 (N_3153,In_806,In_2383);
xor U3154 (N_3154,In_2597,In_55);
and U3155 (N_3155,In_1064,In_2459);
nor U3156 (N_3156,In_350,In_74);
nand U3157 (N_3157,In_2025,In_672);
nor U3158 (N_3158,In_95,In_322);
nand U3159 (N_3159,In_1048,In_2145);
nor U3160 (N_3160,In_743,In_1822);
xnor U3161 (N_3161,In_94,In_203);
or U3162 (N_3162,In_2731,In_1967);
or U3163 (N_3163,In_1536,In_2051);
nor U3164 (N_3164,In_1622,In_1439);
nor U3165 (N_3165,In_1602,In_2184);
or U3166 (N_3166,In_596,In_1037);
nand U3167 (N_3167,In_845,In_1803);
nor U3168 (N_3168,In_1641,In_1476);
nand U3169 (N_3169,In_1328,In_2138);
and U3170 (N_3170,In_1865,In_1129);
nor U3171 (N_3171,In_2067,In_2901);
or U3172 (N_3172,In_2577,In_2642);
nor U3173 (N_3173,In_925,In_466);
or U3174 (N_3174,In_1018,In_1591);
or U3175 (N_3175,In_1589,In_2923);
nand U3176 (N_3176,In_2360,In_338);
or U3177 (N_3177,In_775,In_1068);
xnor U3178 (N_3178,In_607,In_1192);
and U3179 (N_3179,In_1880,In_346);
nand U3180 (N_3180,In_1098,In_1717);
and U3181 (N_3181,In_1511,In_1766);
or U3182 (N_3182,In_2024,In_727);
and U3183 (N_3183,In_1324,In_2033);
nand U3184 (N_3184,In_2888,In_583);
xnor U3185 (N_3185,In_2287,In_304);
and U3186 (N_3186,In_1241,In_428);
and U3187 (N_3187,In_1779,In_1991);
xor U3188 (N_3188,In_2732,In_2132);
xnor U3189 (N_3189,In_1544,In_1584);
nor U3190 (N_3190,In_76,In_2826);
nand U3191 (N_3191,In_1588,In_2424);
nor U3192 (N_3192,In_1717,In_1460);
or U3193 (N_3193,In_1698,In_435);
and U3194 (N_3194,In_2447,In_1287);
nor U3195 (N_3195,In_2912,In_49);
nor U3196 (N_3196,In_1452,In_1660);
or U3197 (N_3197,In_1251,In_1801);
or U3198 (N_3198,In_1353,In_1889);
xor U3199 (N_3199,In_376,In_1509);
or U3200 (N_3200,In_2709,In_1694);
nor U3201 (N_3201,In_2692,In_2701);
nand U3202 (N_3202,In_1581,In_917);
and U3203 (N_3203,In_2619,In_2051);
or U3204 (N_3204,In_208,In_2971);
or U3205 (N_3205,In_2466,In_2319);
and U3206 (N_3206,In_1158,In_1596);
xor U3207 (N_3207,In_1583,In_1748);
and U3208 (N_3208,In_2804,In_2660);
and U3209 (N_3209,In_2293,In_2952);
nor U3210 (N_3210,In_2455,In_1217);
or U3211 (N_3211,In_1847,In_2436);
or U3212 (N_3212,In_1791,In_213);
and U3213 (N_3213,In_446,In_984);
nor U3214 (N_3214,In_2699,In_629);
xnor U3215 (N_3215,In_2836,In_530);
nor U3216 (N_3216,In_2797,In_466);
or U3217 (N_3217,In_2808,In_1126);
and U3218 (N_3218,In_1689,In_2901);
nor U3219 (N_3219,In_717,In_169);
xnor U3220 (N_3220,In_499,In_2154);
and U3221 (N_3221,In_559,In_937);
and U3222 (N_3222,In_2307,In_1549);
and U3223 (N_3223,In_2818,In_690);
or U3224 (N_3224,In_814,In_2070);
or U3225 (N_3225,In_1867,In_2285);
nor U3226 (N_3226,In_2973,In_2037);
nor U3227 (N_3227,In_2520,In_2348);
nand U3228 (N_3228,In_1300,In_2799);
and U3229 (N_3229,In_1159,In_2743);
nor U3230 (N_3230,In_1992,In_1293);
nor U3231 (N_3231,In_970,In_290);
nand U3232 (N_3232,In_2339,In_1628);
nand U3233 (N_3233,In_699,In_1579);
nor U3234 (N_3234,In_2415,In_307);
nor U3235 (N_3235,In_79,In_1547);
nor U3236 (N_3236,In_965,In_2977);
nand U3237 (N_3237,In_1526,In_2912);
or U3238 (N_3238,In_209,In_2718);
and U3239 (N_3239,In_742,In_1686);
and U3240 (N_3240,In_2318,In_266);
nor U3241 (N_3241,In_2100,In_1844);
and U3242 (N_3242,In_1512,In_2330);
and U3243 (N_3243,In_2877,In_824);
and U3244 (N_3244,In_1471,In_449);
xor U3245 (N_3245,In_1941,In_206);
nor U3246 (N_3246,In_769,In_2355);
and U3247 (N_3247,In_1070,In_2972);
nor U3248 (N_3248,In_1315,In_1808);
xnor U3249 (N_3249,In_947,In_1709);
and U3250 (N_3250,In_2693,In_2471);
and U3251 (N_3251,In_653,In_2031);
xnor U3252 (N_3252,In_434,In_1137);
and U3253 (N_3253,In_1802,In_182);
nand U3254 (N_3254,In_2509,In_970);
nor U3255 (N_3255,In_2772,In_1723);
nor U3256 (N_3256,In_752,In_596);
nand U3257 (N_3257,In_1343,In_628);
xnor U3258 (N_3258,In_1965,In_2848);
nor U3259 (N_3259,In_448,In_254);
or U3260 (N_3260,In_870,In_177);
nand U3261 (N_3261,In_236,In_2311);
nor U3262 (N_3262,In_1823,In_1009);
and U3263 (N_3263,In_131,In_2889);
and U3264 (N_3264,In_1331,In_908);
nand U3265 (N_3265,In_1558,In_2405);
xnor U3266 (N_3266,In_1793,In_688);
xor U3267 (N_3267,In_2810,In_720);
and U3268 (N_3268,In_1302,In_1577);
and U3269 (N_3269,In_1253,In_1122);
xnor U3270 (N_3270,In_1620,In_1279);
and U3271 (N_3271,In_2503,In_799);
nand U3272 (N_3272,In_2293,In_2135);
nand U3273 (N_3273,In_2896,In_466);
nor U3274 (N_3274,In_1246,In_2039);
nor U3275 (N_3275,In_1273,In_1921);
nor U3276 (N_3276,In_2020,In_520);
xnor U3277 (N_3277,In_40,In_1031);
and U3278 (N_3278,In_172,In_1195);
nor U3279 (N_3279,In_711,In_2470);
nand U3280 (N_3280,In_2737,In_2849);
xor U3281 (N_3281,In_282,In_2980);
xnor U3282 (N_3282,In_2581,In_492);
or U3283 (N_3283,In_763,In_567);
nand U3284 (N_3284,In_2672,In_1000);
nor U3285 (N_3285,In_2293,In_2510);
nor U3286 (N_3286,In_1852,In_512);
and U3287 (N_3287,In_2772,In_2331);
or U3288 (N_3288,In_1308,In_230);
or U3289 (N_3289,In_930,In_2317);
nand U3290 (N_3290,In_943,In_1670);
nand U3291 (N_3291,In_543,In_2490);
or U3292 (N_3292,In_2060,In_2710);
and U3293 (N_3293,In_1728,In_2345);
xnor U3294 (N_3294,In_221,In_1425);
nand U3295 (N_3295,In_2275,In_943);
nand U3296 (N_3296,In_2978,In_555);
or U3297 (N_3297,In_338,In_2092);
xor U3298 (N_3298,In_2870,In_1987);
and U3299 (N_3299,In_561,In_927);
xnor U3300 (N_3300,In_2579,In_2167);
nand U3301 (N_3301,In_980,In_366);
or U3302 (N_3302,In_2953,In_2487);
and U3303 (N_3303,In_480,In_1343);
xor U3304 (N_3304,In_1117,In_2173);
nand U3305 (N_3305,In_1848,In_1506);
and U3306 (N_3306,In_1213,In_1503);
and U3307 (N_3307,In_52,In_2907);
and U3308 (N_3308,In_1902,In_1085);
nand U3309 (N_3309,In_2907,In_2942);
nor U3310 (N_3310,In_688,In_179);
or U3311 (N_3311,In_1179,In_946);
nor U3312 (N_3312,In_1965,In_1036);
xor U3313 (N_3313,In_2548,In_2474);
xor U3314 (N_3314,In_806,In_2180);
or U3315 (N_3315,In_1730,In_2435);
xnor U3316 (N_3316,In_1733,In_1601);
nand U3317 (N_3317,In_790,In_1926);
nand U3318 (N_3318,In_351,In_697);
or U3319 (N_3319,In_2059,In_2853);
and U3320 (N_3320,In_1832,In_1066);
xnor U3321 (N_3321,In_2774,In_1885);
or U3322 (N_3322,In_2808,In_2665);
and U3323 (N_3323,In_191,In_2290);
nor U3324 (N_3324,In_1856,In_1950);
nand U3325 (N_3325,In_2180,In_1588);
nor U3326 (N_3326,In_1011,In_2899);
xor U3327 (N_3327,In_2054,In_2888);
nand U3328 (N_3328,In_2156,In_772);
xnor U3329 (N_3329,In_2030,In_2605);
nor U3330 (N_3330,In_583,In_468);
and U3331 (N_3331,In_444,In_1096);
nand U3332 (N_3332,In_1628,In_2535);
and U3333 (N_3333,In_2132,In_1969);
xnor U3334 (N_3334,In_2882,In_1961);
nor U3335 (N_3335,In_1466,In_268);
nand U3336 (N_3336,In_2390,In_1164);
or U3337 (N_3337,In_1886,In_1192);
nand U3338 (N_3338,In_1490,In_543);
xnor U3339 (N_3339,In_607,In_880);
xnor U3340 (N_3340,In_627,In_1789);
nand U3341 (N_3341,In_1928,In_2236);
xnor U3342 (N_3342,In_2928,In_770);
xor U3343 (N_3343,In_1036,In_1305);
nor U3344 (N_3344,In_1347,In_1739);
and U3345 (N_3345,In_905,In_2698);
nand U3346 (N_3346,In_2766,In_2820);
or U3347 (N_3347,In_439,In_566);
nor U3348 (N_3348,In_1092,In_1086);
xnor U3349 (N_3349,In_978,In_347);
nor U3350 (N_3350,In_789,In_2606);
nor U3351 (N_3351,In_63,In_492);
xor U3352 (N_3352,In_1222,In_2130);
or U3353 (N_3353,In_1352,In_1269);
and U3354 (N_3354,In_2511,In_1299);
nor U3355 (N_3355,In_1431,In_1391);
xnor U3356 (N_3356,In_2331,In_2579);
xnor U3357 (N_3357,In_421,In_1757);
xnor U3358 (N_3358,In_2114,In_2998);
nor U3359 (N_3359,In_2123,In_1061);
and U3360 (N_3360,In_2919,In_2461);
xnor U3361 (N_3361,In_369,In_1813);
or U3362 (N_3362,In_1991,In_2977);
or U3363 (N_3363,In_1319,In_1400);
nor U3364 (N_3364,In_2073,In_1018);
and U3365 (N_3365,In_411,In_35);
or U3366 (N_3366,In_1078,In_2605);
nor U3367 (N_3367,In_580,In_1816);
nor U3368 (N_3368,In_471,In_1789);
xor U3369 (N_3369,In_2924,In_182);
nand U3370 (N_3370,In_262,In_416);
and U3371 (N_3371,In_234,In_88);
nand U3372 (N_3372,In_786,In_1565);
xor U3373 (N_3373,In_2720,In_1059);
xnor U3374 (N_3374,In_2472,In_2963);
nand U3375 (N_3375,In_48,In_1319);
nand U3376 (N_3376,In_2517,In_436);
or U3377 (N_3377,In_1969,In_962);
or U3378 (N_3378,In_2703,In_856);
nor U3379 (N_3379,In_1944,In_2927);
and U3380 (N_3380,In_930,In_1974);
and U3381 (N_3381,In_2864,In_1201);
and U3382 (N_3382,In_2496,In_111);
and U3383 (N_3383,In_1802,In_1180);
nand U3384 (N_3384,In_1995,In_1758);
xor U3385 (N_3385,In_2600,In_2496);
xor U3386 (N_3386,In_2650,In_2229);
or U3387 (N_3387,In_1844,In_907);
xnor U3388 (N_3388,In_1151,In_2434);
xor U3389 (N_3389,In_2607,In_2406);
nand U3390 (N_3390,In_1907,In_2172);
nor U3391 (N_3391,In_2470,In_2034);
nand U3392 (N_3392,In_1254,In_1496);
xor U3393 (N_3393,In_673,In_576);
nor U3394 (N_3394,In_355,In_2964);
nand U3395 (N_3395,In_2064,In_1822);
and U3396 (N_3396,In_1218,In_314);
and U3397 (N_3397,In_305,In_186);
and U3398 (N_3398,In_1611,In_411);
and U3399 (N_3399,In_2744,In_2152);
nand U3400 (N_3400,In_419,In_1554);
nor U3401 (N_3401,In_2852,In_224);
or U3402 (N_3402,In_2058,In_252);
xnor U3403 (N_3403,In_2938,In_1372);
nand U3404 (N_3404,In_1316,In_1988);
and U3405 (N_3405,In_1363,In_1891);
and U3406 (N_3406,In_2688,In_1638);
nor U3407 (N_3407,In_1822,In_1116);
and U3408 (N_3408,In_1609,In_1607);
xor U3409 (N_3409,In_1194,In_1547);
or U3410 (N_3410,In_2628,In_1835);
nand U3411 (N_3411,In_1776,In_339);
xor U3412 (N_3412,In_686,In_2012);
xnor U3413 (N_3413,In_1012,In_1114);
and U3414 (N_3414,In_484,In_1089);
and U3415 (N_3415,In_991,In_1956);
nand U3416 (N_3416,In_2051,In_3);
and U3417 (N_3417,In_429,In_2953);
nand U3418 (N_3418,In_880,In_515);
xor U3419 (N_3419,In_1901,In_334);
nor U3420 (N_3420,In_1925,In_512);
nand U3421 (N_3421,In_1222,In_725);
nor U3422 (N_3422,In_2814,In_2060);
and U3423 (N_3423,In_1645,In_819);
or U3424 (N_3424,In_430,In_1304);
or U3425 (N_3425,In_585,In_2314);
nand U3426 (N_3426,In_1516,In_1625);
nor U3427 (N_3427,In_1032,In_2524);
and U3428 (N_3428,In_2289,In_1198);
nor U3429 (N_3429,In_208,In_1925);
xor U3430 (N_3430,In_1457,In_1611);
and U3431 (N_3431,In_381,In_2212);
xor U3432 (N_3432,In_1096,In_1711);
and U3433 (N_3433,In_2639,In_1656);
nor U3434 (N_3434,In_1554,In_1371);
xor U3435 (N_3435,In_1080,In_573);
and U3436 (N_3436,In_926,In_1654);
nand U3437 (N_3437,In_1165,In_1823);
and U3438 (N_3438,In_581,In_2731);
nand U3439 (N_3439,In_89,In_2976);
xnor U3440 (N_3440,In_1791,In_132);
or U3441 (N_3441,In_438,In_1822);
xor U3442 (N_3442,In_1146,In_898);
xnor U3443 (N_3443,In_618,In_1242);
xnor U3444 (N_3444,In_2879,In_516);
nor U3445 (N_3445,In_860,In_921);
nand U3446 (N_3446,In_1503,In_1182);
xnor U3447 (N_3447,In_1792,In_2343);
xor U3448 (N_3448,In_561,In_96);
nor U3449 (N_3449,In_482,In_673);
xor U3450 (N_3450,In_2550,In_1830);
xnor U3451 (N_3451,In_1721,In_2665);
xor U3452 (N_3452,In_1499,In_571);
xor U3453 (N_3453,In_481,In_2532);
xnor U3454 (N_3454,In_2093,In_2071);
and U3455 (N_3455,In_1218,In_138);
and U3456 (N_3456,In_410,In_1713);
and U3457 (N_3457,In_2554,In_1622);
and U3458 (N_3458,In_1418,In_1585);
nor U3459 (N_3459,In_1382,In_2785);
nor U3460 (N_3460,In_613,In_80);
and U3461 (N_3461,In_928,In_2887);
nand U3462 (N_3462,In_1336,In_962);
xnor U3463 (N_3463,In_1013,In_2542);
nand U3464 (N_3464,In_2320,In_1126);
nand U3465 (N_3465,In_2701,In_949);
and U3466 (N_3466,In_2883,In_1315);
or U3467 (N_3467,In_167,In_2047);
nand U3468 (N_3468,In_1838,In_942);
or U3469 (N_3469,In_322,In_2130);
or U3470 (N_3470,In_1978,In_1666);
and U3471 (N_3471,In_1325,In_2382);
or U3472 (N_3472,In_2875,In_1487);
nor U3473 (N_3473,In_675,In_736);
nor U3474 (N_3474,In_1805,In_245);
xor U3475 (N_3475,In_2757,In_765);
or U3476 (N_3476,In_1178,In_2997);
nor U3477 (N_3477,In_896,In_756);
xnor U3478 (N_3478,In_1228,In_599);
nand U3479 (N_3479,In_1643,In_794);
or U3480 (N_3480,In_855,In_433);
or U3481 (N_3481,In_2309,In_170);
and U3482 (N_3482,In_397,In_1928);
xor U3483 (N_3483,In_1155,In_2727);
nand U3484 (N_3484,In_2397,In_1417);
or U3485 (N_3485,In_2222,In_1383);
nor U3486 (N_3486,In_2382,In_2397);
nand U3487 (N_3487,In_1911,In_2299);
or U3488 (N_3488,In_823,In_874);
and U3489 (N_3489,In_1273,In_2329);
nor U3490 (N_3490,In_1900,In_458);
and U3491 (N_3491,In_2060,In_596);
or U3492 (N_3492,In_2378,In_2526);
and U3493 (N_3493,In_2370,In_562);
and U3494 (N_3494,In_226,In_2533);
nand U3495 (N_3495,In_2335,In_1593);
nand U3496 (N_3496,In_664,In_1613);
nand U3497 (N_3497,In_1946,In_2110);
xor U3498 (N_3498,In_1841,In_1915);
xor U3499 (N_3499,In_1288,In_1399);
nand U3500 (N_3500,In_925,In_237);
or U3501 (N_3501,In_2994,In_2722);
or U3502 (N_3502,In_1319,In_2895);
or U3503 (N_3503,In_1923,In_812);
or U3504 (N_3504,In_847,In_418);
nor U3505 (N_3505,In_2587,In_466);
and U3506 (N_3506,In_2539,In_2882);
nand U3507 (N_3507,In_1724,In_1590);
nand U3508 (N_3508,In_1797,In_348);
or U3509 (N_3509,In_244,In_1487);
nand U3510 (N_3510,In_636,In_569);
nor U3511 (N_3511,In_805,In_2248);
and U3512 (N_3512,In_1230,In_1179);
or U3513 (N_3513,In_413,In_259);
nor U3514 (N_3514,In_1287,In_2130);
and U3515 (N_3515,In_610,In_1025);
nor U3516 (N_3516,In_721,In_76);
nand U3517 (N_3517,In_1677,In_1572);
nand U3518 (N_3518,In_2216,In_2285);
and U3519 (N_3519,In_1628,In_2202);
or U3520 (N_3520,In_2634,In_248);
and U3521 (N_3521,In_2041,In_2978);
or U3522 (N_3522,In_1760,In_238);
nor U3523 (N_3523,In_598,In_2107);
nor U3524 (N_3524,In_2555,In_2539);
and U3525 (N_3525,In_576,In_2305);
nand U3526 (N_3526,In_876,In_1948);
nor U3527 (N_3527,In_1108,In_1676);
xor U3528 (N_3528,In_888,In_2630);
xor U3529 (N_3529,In_2169,In_2201);
and U3530 (N_3530,In_1735,In_142);
nor U3531 (N_3531,In_2324,In_1428);
and U3532 (N_3532,In_2985,In_2048);
xnor U3533 (N_3533,In_1712,In_558);
nor U3534 (N_3534,In_393,In_2982);
nor U3535 (N_3535,In_2818,In_2751);
nand U3536 (N_3536,In_1975,In_2700);
xor U3537 (N_3537,In_917,In_2909);
xor U3538 (N_3538,In_1130,In_33);
and U3539 (N_3539,In_243,In_711);
nor U3540 (N_3540,In_1372,In_899);
nor U3541 (N_3541,In_2294,In_1586);
or U3542 (N_3542,In_1984,In_941);
nor U3543 (N_3543,In_2972,In_2747);
nor U3544 (N_3544,In_2076,In_1090);
nor U3545 (N_3545,In_725,In_1228);
and U3546 (N_3546,In_25,In_2326);
or U3547 (N_3547,In_165,In_2447);
nand U3548 (N_3548,In_1013,In_1117);
and U3549 (N_3549,In_2022,In_694);
nand U3550 (N_3550,In_2532,In_841);
nand U3551 (N_3551,In_2665,In_504);
nand U3552 (N_3552,In_186,In_1155);
or U3553 (N_3553,In_855,In_1158);
or U3554 (N_3554,In_1890,In_963);
or U3555 (N_3555,In_152,In_1009);
xor U3556 (N_3556,In_1234,In_1670);
and U3557 (N_3557,In_1988,In_1620);
nand U3558 (N_3558,In_1397,In_541);
xor U3559 (N_3559,In_1603,In_2913);
xnor U3560 (N_3560,In_2568,In_1017);
nor U3561 (N_3561,In_2857,In_155);
xnor U3562 (N_3562,In_2626,In_2590);
xor U3563 (N_3563,In_1760,In_472);
nand U3564 (N_3564,In_1283,In_2793);
nand U3565 (N_3565,In_1147,In_2482);
nand U3566 (N_3566,In_2897,In_746);
and U3567 (N_3567,In_0,In_1083);
xnor U3568 (N_3568,In_2596,In_349);
xor U3569 (N_3569,In_2617,In_2129);
nand U3570 (N_3570,In_2167,In_727);
nor U3571 (N_3571,In_1445,In_2168);
or U3572 (N_3572,In_2440,In_2553);
nand U3573 (N_3573,In_2003,In_315);
and U3574 (N_3574,In_825,In_1145);
xor U3575 (N_3575,In_2987,In_374);
xnor U3576 (N_3576,In_852,In_1316);
or U3577 (N_3577,In_1770,In_39);
nand U3578 (N_3578,In_1367,In_2742);
nand U3579 (N_3579,In_339,In_1842);
and U3580 (N_3580,In_2432,In_1004);
xor U3581 (N_3581,In_2715,In_2711);
or U3582 (N_3582,In_1866,In_1368);
nand U3583 (N_3583,In_2687,In_239);
nand U3584 (N_3584,In_2908,In_1453);
xor U3585 (N_3585,In_1803,In_2652);
nor U3586 (N_3586,In_2270,In_1049);
nand U3587 (N_3587,In_1099,In_822);
and U3588 (N_3588,In_2024,In_2394);
or U3589 (N_3589,In_2715,In_1611);
or U3590 (N_3590,In_2751,In_2056);
nand U3591 (N_3591,In_285,In_304);
and U3592 (N_3592,In_762,In_538);
nand U3593 (N_3593,In_1745,In_196);
nor U3594 (N_3594,In_2432,In_2981);
xor U3595 (N_3595,In_191,In_2028);
nor U3596 (N_3596,In_1886,In_2868);
and U3597 (N_3597,In_1190,In_1187);
xor U3598 (N_3598,In_993,In_2323);
nor U3599 (N_3599,In_797,In_2054);
nand U3600 (N_3600,In_796,In_160);
nor U3601 (N_3601,In_2848,In_2874);
nand U3602 (N_3602,In_2233,In_1624);
xor U3603 (N_3603,In_225,In_1522);
and U3604 (N_3604,In_1808,In_2699);
xnor U3605 (N_3605,In_254,In_2881);
or U3606 (N_3606,In_2406,In_1926);
and U3607 (N_3607,In_121,In_2148);
or U3608 (N_3608,In_1080,In_1688);
xor U3609 (N_3609,In_2325,In_159);
xor U3610 (N_3610,In_1537,In_2806);
and U3611 (N_3611,In_1885,In_292);
nor U3612 (N_3612,In_837,In_2953);
and U3613 (N_3613,In_46,In_2153);
or U3614 (N_3614,In_2173,In_287);
xor U3615 (N_3615,In_2252,In_1502);
nor U3616 (N_3616,In_1999,In_1754);
or U3617 (N_3617,In_1279,In_2826);
xnor U3618 (N_3618,In_1498,In_619);
nor U3619 (N_3619,In_2059,In_338);
xnor U3620 (N_3620,In_112,In_1658);
or U3621 (N_3621,In_345,In_2747);
nor U3622 (N_3622,In_1440,In_2101);
xor U3623 (N_3623,In_1032,In_1386);
nand U3624 (N_3624,In_1231,In_90);
nand U3625 (N_3625,In_1941,In_2003);
and U3626 (N_3626,In_1572,In_2069);
nand U3627 (N_3627,In_250,In_2296);
or U3628 (N_3628,In_2621,In_2690);
nor U3629 (N_3629,In_1772,In_830);
or U3630 (N_3630,In_2466,In_1755);
nand U3631 (N_3631,In_899,In_388);
nor U3632 (N_3632,In_1958,In_2480);
nor U3633 (N_3633,In_2870,In_2730);
nand U3634 (N_3634,In_2193,In_798);
nor U3635 (N_3635,In_444,In_2893);
nor U3636 (N_3636,In_925,In_1353);
xnor U3637 (N_3637,In_557,In_1741);
nor U3638 (N_3638,In_920,In_2818);
or U3639 (N_3639,In_1627,In_159);
nand U3640 (N_3640,In_623,In_2896);
xor U3641 (N_3641,In_1815,In_1622);
or U3642 (N_3642,In_1345,In_49);
xor U3643 (N_3643,In_2463,In_1234);
or U3644 (N_3644,In_1959,In_855);
nand U3645 (N_3645,In_2792,In_24);
nor U3646 (N_3646,In_550,In_2696);
nor U3647 (N_3647,In_1340,In_1972);
and U3648 (N_3648,In_1752,In_2830);
or U3649 (N_3649,In_2237,In_364);
and U3650 (N_3650,In_2491,In_1106);
nor U3651 (N_3651,In_24,In_1248);
nor U3652 (N_3652,In_2015,In_1939);
or U3653 (N_3653,In_2204,In_2222);
nand U3654 (N_3654,In_600,In_242);
and U3655 (N_3655,In_1535,In_398);
and U3656 (N_3656,In_82,In_2682);
nand U3657 (N_3657,In_981,In_2516);
xor U3658 (N_3658,In_1056,In_2413);
xnor U3659 (N_3659,In_2911,In_789);
or U3660 (N_3660,In_970,In_369);
or U3661 (N_3661,In_318,In_540);
or U3662 (N_3662,In_2081,In_1101);
or U3663 (N_3663,In_1504,In_863);
xnor U3664 (N_3664,In_81,In_791);
nand U3665 (N_3665,In_1907,In_184);
and U3666 (N_3666,In_2305,In_33);
nor U3667 (N_3667,In_1504,In_2707);
and U3668 (N_3668,In_675,In_1109);
nor U3669 (N_3669,In_1123,In_203);
xor U3670 (N_3670,In_1083,In_952);
xor U3671 (N_3671,In_504,In_382);
xnor U3672 (N_3672,In_581,In_2900);
nand U3673 (N_3673,In_1614,In_169);
or U3674 (N_3674,In_675,In_1228);
nand U3675 (N_3675,In_213,In_978);
nand U3676 (N_3676,In_2058,In_2760);
and U3677 (N_3677,In_2074,In_2970);
xor U3678 (N_3678,In_2046,In_1334);
or U3679 (N_3679,In_2229,In_1533);
and U3680 (N_3680,In_302,In_430);
or U3681 (N_3681,In_2740,In_1462);
nor U3682 (N_3682,In_1161,In_2726);
xnor U3683 (N_3683,In_935,In_1424);
and U3684 (N_3684,In_243,In_570);
and U3685 (N_3685,In_1410,In_961);
nand U3686 (N_3686,In_424,In_922);
xnor U3687 (N_3687,In_593,In_324);
nor U3688 (N_3688,In_1261,In_2258);
or U3689 (N_3689,In_2823,In_1057);
or U3690 (N_3690,In_810,In_954);
nor U3691 (N_3691,In_2721,In_278);
nor U3692 (N_3692,In_2391,In_2822);
and U3693 (N_3693,In_1543,In_1437);
and U3694 (N_3694,In_398,In_1951);
nor U3695 (N_3695,In_2416,In_1711);
nor U3696 (N_3696,In_308,In_1985);
or U3697 (N_3697,In_1494,In_1879);
nor U3698 (N_3698,In_221,In_2520);
nand U3699 (N_3699,In_1259,In_2817);
xor U3700 (N_3700,In_664,In_2261);
and U3701 (N_3701,In_2637,In_948);
nand U3702 (N_3702,In_2932,In_954);
nand U3703 (N_3703,In_2471,In_2657);
xnor U3704 (N_3704,In_2402,In_2977);
or U3705 (N_3705,In_1009,In_2902);
nor U3706 (N_3706,In_1786,In_2292);
nand U3707 (N_3707,In_397,In_326);
or U3708 (N_3708,In_2875,In_519);
or U3709 (N_3709,In_2535,In_2269);
xnor U3710 (N_3710,In_1799,In_2895);
and U3711 (N_3711,In_1018,In_1837);
nor U3712 (N_3712,In_2521,In_1363);
xnor U3713 (N_3713,In_1461,In_2168);
xnor U3714 (N_3714,In_1056,In_92);
or U3715 (N_3715,In_1825,In_71);
nand U3716 (N_3716,In_1426,In_2116);
xnor U3717 (N_3717,In_1673,In_819);
nor U3718 (N_3718,In_128,In_2227);
nand U3719 (N_3719,In_478,In_2899);
xor U3720 (N_3720,In_2128,In_2535);
and U3721 (N_3721,In_1508,In_965);
nor U3722 (N_3722,In_943,In_2947);
or U3723 (N_3723,In_1190,In_810);
xnor U3724 (N_3724,In_1713,In_981);
xor U3725 (N_3725,In_1156,In_1445);
nor U3726 (N_3726,In_866,In_381);
nor U3727 (N_3727,In_2009,In_1770);
nor U3728 (N_3728,In_2081,In_2337);
or U3729 (N_3729,In_2886,In_194);
nand U3730 (N_3730,In_2971,In_246);
xnor U3731 (N_3731,In_2530,In_1824);
or U3732 (N_3732,In_1181,In_1300);
or U3733 (N_3733,In_1662,In_805);
nand U3734 (N_3734,In_2775,In_129);
nor U3735 (N_3735,In_2933,In_163);
nor U3736 (N_3736,In_441,In_145);
and U3737 (N_3737,In_528,In_47);
nand U3738 (N_3738,In_2393,In_2664);
and U3739 (N_3739,In_793,In_305);
nor U3740 (N_3740,In_2961,In_121);
nand U3741 (N_3741,In_2415,In_2438);
or U3742 (N_3742,In_2968,In_1071);
nor U3743 (N_3743,In_411,In_2768);
or U3744 (N_3744,In_1177,In_659);
xnor U3745 (N_3745,In_848,In_2165);
nand U3746 (N_3746,In_2147,In_2476);
and U3747 (N_3747,In_174,In_2847);
nand U3748 (N_3748,In_161,In_2640);
nand U3749 (N_3749,In_1637,In_2501);
nand U3750 (N_3750,In_2123,In_2833);
nand U3751 (N_3751,In_648,In_2799);
xor U3752 (N_3752,In_2169,In_2352);
xor U3753 (N_3753,In_2125,In_1382);
nor U3754 (N_3754,In_247,In_803);
nand U3755 (N_3755,In_940,In_901);
or U3756 (N_3756,In_2965,In_1161);
and U3757 (N_3757,In_1648,In_1427);
or U3758 (N_3758,In_2321,In_515);
nor U3759 (N_3759,In_2699,In_1488);
and U3760 (N_3760,In_1489,In_1556);
xnor U3761 (N_3761,In_498,In_2589);
nor U3762 (N_3762,In_964,In_2860);
and U3763 (N_3763,In_1078,In_48);
and U3764 (N_3764,In_2025,In_2929);
xnor U3765 (N_3765,In_399,In_1128);
nor U3766 (N_3766,In_1452,In_2591);
or U3767 (N_3767,In_1781,In_1096);
or U3768 (N_3768,In_2824,In_715);
or U3769 (N_3769,In_2750,In_186);
nand U3770 (N_3770,In_958,In_164);
and U3771 (N_3771,In_1529,In_833);
and U3772 (N_3772,In_23,In_516);
or U3773 (N_3773,In_1958,In_921);
or U3774 (N_3774,In_1814,In_2372);
and U3775 (N_3775,In_1420,In_425);
xor U3776 (N_3776,In_221,In_811);
xor U3777 (N_3777,In_2843,In_2007);
nand U3778 (N_3778,In_1475,In_2768);
nand U3779 (N_3779,In_2505,In_1700);
nand U3780 (N_3780,In_383,In_2132);
nand U3781 (N_3781,In_119,In_2727);
and U3782 (N_3782,In_2587,In_1824);
nand U3783 (N_3783,In_798,In_1215);
and U3784 (N_3784,In_2829,In_1759);
or U3785 (N_3785,In_2453,In_1163);
nor U3786 (N_3786,In_2089,In_611);
nand U3787 (N_3787,In_120,In_2660);
nor U3788 (N_3788,In_520,In_1044);
nor U3789 (N_3789,In_1326,In_2632);
xor U3790 (N_3790,In_1350,In_765);
nand U3791 (N_3791,In_1320,In_1794);
xor U3792 (N_3792,In_2732,In_1821);
xor U3793 (N_3793,In_2787,In_70);
nand U3794 (N_3794,In_2656,In_1256);
xnor U3795 (N_3795,In_1671,In_785);
nand U3796 (N_3796,In_670,In_759);
xnor U3797 (N_3797,In_2778,In_840);
and U3798 (N_3798,In_1487,In_1521);
nand U3799 (N_3799,In_2319,In_1107);
and U3800 (N_3800,In_574,In_1382);
or U3801 (N_3801,In_614,In_1743);
nor U3802 (N_3802,In_2016,In_1814);
nand U3803 (N_3803,In_1592,In_2144);
or U3804 (N_3804,In_1556,In_1111);
or U3805 (N_3805,In_1848,In_2853);
nand U3806 (N_3806,In_2185,In_763);
and U3807 (N_3807,In_1932,In_465);
or U3808 (N_3808,In_31,In_2248);
nor U3809 (N_3809,In_2520,In_2400);
nor U3810 (N_3810,In_2031,In_2696);
and U3811 (N_3811,In_434,In_2572);
xnor U3812 (N_3812,In_1670,In_2187);
nor U3813 (N_3813,In_43,In_408);
and U3814 (N_3814,In_2980,In_291);
nor U3815 (N_3815,In_908,In_53);
or U3816 (N_3816,In_498,In_2591);
nand U3817 (N_3817,In_1872,In_853);
nor U3818 (N_3818,In_2175,In_1764);
nor U3819 (N_3819,In_2959,In_960);
or U3820 (N_3820,In_1753,In_1388);
nor U3821 (N_3821,In_2982,In_1950);
and U3822 (N_3822,In_232,In_1792);
or U3823 (N_3823,In_1790,In_2346);
xnor U3824 (N_3824,In_2353,In_2327);
and U3825 (N_3825,In_2556,In_409);
or U3826 (N_3826,In_1247,In_2866);
nor U3827 (N_3827,In_543,In_1701);
or U3828 (N_3828,In_474,In_1878);
nor U3829 (N_3829,In_1269,In_2201);
nor U3830 (N_3830,In_1893,In_1750);
nor U3831 (N_3831,In_1826,In_2459);
nand U3832 (N_3832,In_206,In_2908);
nand U3833 (N_3833,In_2517,In_1470);
nand U3834 (N_3834,In_1173,In_1269);
xnor U3835 (N_3835,In_1291,In_366);
or U3836 (N_3836,In_355,In_2780);
nand U3837 (N_3837,In_416,In_665);
and U3838 (N_3838,In_2393,In_685);
xor U3839 (N_3839,In_172,In_1432);
or U3840 (N_3840,In_1420,In_957);
nor U3841 (N_3841,In_2500,In_319);
and U3842 (N_3842,In_692,In_1404);
nand U3843 (N_3843,In_2142,In_630);
and U3844 (N_3844,In_1033,In_632);
nand U3845 (N_3845,In_808,In_2949);
xor U3846 (N_3846,In_2316,In_2925);
nor U3847 (N_3847,In_1035,In_2324);
or U3848 (N_3848,In_2426,In_2979);
nand U3849 (N_3849,In_708,In_2165);
nor U3850 (N_3850,In_2926,In_1410);
nand U3851 (N_3851,In_2756,In_2733);
nor U3852 (N_3852,In_1023,In_762);
and U3853 (N_3853,In_2191,In_882);
and U3854 (N_3854,In_153,In_1883);
and U3855 (N_3855,In_1641,In_2081);
nor U3856 (N_3856,In_2529,In_42);
nor U3857 (N_3857,In_1847,In_855);
nor U3858 (N_3858,In_2711,In_1374);
and U3859 (N_3859,In_1949,In_2780);
and U3860 (N_3860,In_1763,In_2945);
xnor U3861 (N_3861,In_2099,In_2773);
xor U3862 (N_3862,In_299,In_1790);
nand U3863 (N_3863,In_1105,In_2463);
nand U3864 (N_3864,In_2389,In_952);
and U3865 (N_3865,In_477,In_2588);
and U3866 (N_3866,In_2562,In_2536);
nor U3867 (N_3867,In_470,In_1186);
xnor U3868 (N_3868,In_2615,In_1392);
nor U3869 (N_3869,In_1988,In_1753);
nor U3870 (N_3870,In_619,In_2192);
and U3871 (N_3871,In_1433,In_2074);
nand U3872 (N_3872,In_1069,In_666);
or U3873 (N_3873,In_370,In_385);
nand U3874 (N_3874,In_1831,In_366);
nor U3875 (N_3875,In_1107,In_300);
nand U3876 (N_3876,In_403,In_323);
and U3877 (N_3877,In_2320,In_1385);
and U3878 (N_3878,In_2534,In_2298);
nand U3879 (N_3879,In_1222,In_1854);
and U3880 (N_3880,In_2830,In_2117);
xor U3881 (N_3881,In_1935,In_521);
or U3882 (N_3882,In_33,In_1116);
xor U3883 (N_3883,In_2495,In_107);
or U3884 (N_3884,In_1815,In_952);
nand U3885 (N_3885,In_103,In_690);
nand U3886 (N_3886,In_1481,In_1145);
and U3887 (N_3887,In_383,In_41);
xnor U3888 (N_3888,In_331,In_728);
nor U3889 (N_3889,In_2764,In_2991);
or U3890 (N_3890,In_346,In_989);
nor U3891 (N_3891,In_937,In_204);
and U3892 (N_3892,In_2803,In_1562);
and U3893 (N_3893,In_2675,In_2972);
nand U3894 (N_3894,In_249,In_2805);
nor U3895 (N_3895,In_2573,In_2574);
xnor U3896 (N_3896,In_414,In_1358);
nor U3897 (N_3897,In_224,In_2987);
xor U3898 (N_3898,In_42,In_757);
xor U3899 (N_3899,In_7,In_2169);
or U3900 (N_3900,In_2657,In_357);
xor U3901 (N_3901,In_1500,In_422);
xor U3902 (N_3902,In_602,In_1458);
and U3903 (N_3903,In_1236,In_1306);
nor U3904 (N_3904,In_18,In_1539);
xor U3905 (N_3905,In_430,In_2244);
xor U3906 (N_3906,In_1349,In_2012);
or U3907 (N_3907,In_2452,In_1206);
and U3908 (N_3908,In_2135,In_2217);
nand U3909 (N_3909,In_603,In_2013);
nor U3910 (N_3910,In_428,In_2092);
nor U3911 (N_3911,In_2720,In_118);
nor U3912 (N_3912,In_2966,In_1776);
nand U3913 (N_3913,In_2170,In_2343);
nand U3914 (N_3914,In_636,In_2887);
nand U3915 (N_3915,In_2772,In_546);
nand U3916 (N_3916,In_695,In_867);
xnor U3917 (N_3917,In_1356,In_1203);
and U3918 (N_3918,In_1075,In_544);
nor U3919 (N_3919,In_30,In_428);
nor U3920 (N_3920,In_2496,In_1274);
nor U3921 (N_3921,In_678,In_2195);
and U3922 (N_3922,In_1288,In_806);
nor U3923 (N_3923,In_1891,In_1045);
nand U3924 (N_3924,In_1408,In_2389);
and U3925 (N_3925,In_796,In_900);
nor U3926 (N_3926,In_359,In_1924);
or U3927 (N_3927,In_622,In_705);
nand U3928 (N_3928,In_1357,In_2647);
nand U3929 (N_3929,In_930,In_1400);
nand U3930 (N_3930,In_803,In_2764);
or U3931 (N_3931,In_166,In_2175);
nand U3932 (N_3932,In_1174,In_2463);
xor U3933 (N_3933,In_185,In_483);
nand U3934 (N_3934,In_2764,In_684);
and U3935 (N_3935,In_1094,In_1613);
or U3936 (N_3936,In_2758,In_1111);
xnor U3937 (N_3937,In_2820,In_1245);
xnor U3938 (N_3938,In_320,In_1931);
nor U3939 (N_3939,In_2930,In_1901);
nand U3940 (N_3940,In_1371,In_2700);
xnor U3941 (N_3941,In_377,In_1108);
or U3942 (N_3942,In_1858,In_1598);
or U3943 (N_3943,In_2682,In_480);
nand U3944 (N_3944,In_1536,In_2366);
and U3945 (N_3945,In_1811,In_1124);
nand U3946 (N_3946,In_1036,In_141);
or U3947 (N_3947,In_2096,In_2679);
nand U3948 (N_3948,In_623,In_1710);
nand U3949 (N_3949,In_2982,In_2439);
xnor U3950 (N_3950,In_532,In_2242);
nor U3951 (N_3951,In_2196,In_411);
and U3952 (N_3952,In_1693,In_949);
nor U3953 (N_3953,In_1727,In_2066);
or U3954 (N_3954,In_2792,In_1215);
xor U3955 (N_3955,In_1410,In_2971);
nand U3956 (N_3956,In_338,In_1762);
nand U3957 (N_3957,In_2783,In_1195);
nor U3958 (N_3958,In_2720,In_1853);
and U3959 (N_3959,In_2140,In_1087);
nor U3960 (N_3960,In_1433,In_2610);
or U3961 (N_3961,In_1087,In_2901);
nor U3962 (N_3962,In_337,In_2040);
xor U3963 (N_3963,In_1074,In_290);
xor U3964 (N_3964,In_836,In_2528);
nand U3965 (N_3965,In_2754,In_498);
nand U3966 (N_3966,In_2719,In_2378);
xnor U3967 (N_3967,In_2642,In_1080);
nand U3968 (N_3968,In_233,In_2320);
xor U3969 (N_3969,In_1809,In_2891);
nor U3970 (N_3970,In_2809,In_717);
or U3971 (N_3971,In_2032,In_2988);
or U3972 (N_3972,In_487,In_2571);
or U3973 (N_3973,In_354,In_1230);
or U3974 (N_3974,In_305,In_2969);
and U3975 (N_3975,In_2610,In_1839);
nor U3976 (N_3976,In_2162,In_1134);
nor U3977 (N_3977,In_982,In_126);
xnor U3978 (N_3978,In_2707,In_2224);
nor U3979 (N_3979,In_1322,In_2501);
and U3980 (N_3980,In_487,In_1931);
nor U3981 (N_3981,In_610,In_713);
nor U3982 (N_3982,In_2337,In_1572);
or U3983 (N_3983,In_2228,In_866);
xor U3984 (N_3984,In_2733,In_144);
xnor U3985 (N_3985,In_1770,In_2521);
and U3986 (N_3986,In_1174,In_1319);
nand U3987 (N_3987,In_252,In_2772);
nand U3988 (N_3988,In_824,In_1867);
or U3989 (N_3989,In_2263,In_2963);
xnor U3990 (N_3990,In_1248,In_456);
nor U3991 (N_3991,In_254,In_817);
nand U3992 (N_3992,In_325,In_2286);
xor U3993 (N_3993,In_2551,In_2461);
xnor U3994 (N_3994,In_2338,In_1973);
nor U3995 (N_3995,In_886,In_761);
xnor U3996 (N_3996,In_1159,In_2594);
nor U3997 (N_3997,In_2484,In_1205);
or U3998 (N_3998,In_1707,In_1549);
xor U3999 (N_3999,In_2876,In_1066);
and U4000 (N_4000,In_1028,In_627);
or U4001 (N_4001,In_618,In_1563);
nand U4002 (N_4002,In_1907,In_2435);
nor U4003 (N_4003,In_696,In_2558);
or U4004 (N_4004,In_222,In_2847);
or U4005 (N_4005,In_410,In_1911);
or U4006 (N_4006,In_2127,In_1632);
or U4007 (N_4007,In_434,In_530);
nor U4008 (N_4008,In_1972,In_2788);
nor U4009 (N_4009,In_2324,In_1039);
nor U4010 (N_4010,In_1670,In_2485);
nor U4011 (N_4011,In_367,In_2982);
xnor U4012 (N_4012,In_1716,In_1965);
xnor U4013 (N_4013,In_715,In_2894);
nand U4014 (N_4014,In_105,In_1819);
and U4015 (N_4015,In_2575,In_2304);
and U4016 (N_4016,In_129,In_1592);
nor U4017 (N_4017,In_2564,In_2966);
nand U4018 (N_4018,In_2911,In_2072);
or U4019 (N_4019,In_1419,In_1358);
nor U4020 (N_4020,In_758,In_1712);
xor U4021 (N_4021,In_2306,In_564);
xor U4022 (N_4022,In_2878,In_596);
nor U4023 (N_4023,In_2907,In_458);
nor U4024 (N_4024,In_1828,In_2920);
or U4025 (N_4025,In_1728,In_621);
nor U4026 (N_4026,In_658,In_1935);
or U4027 (N_4027,In_77,In_782);
xor U4028 (N_4028,In_1746,In_1035);
and U4029 (N_4029,In_982,In_1383);
or U4030 (N_4030,In_2429,In_1338);
and U4031 (N_4031,In_2321,In_1011);
nor U4032 (N_4032,In_1385,In_697);
xnor U4033 (N_4033,In_1673,In_2157);
and U4034 (N_4034,In_2350,In_1753);
or U4035 (N_4035,In_1283,In_2941);
nor U4036 (N_4036,In_2451,In_1491);
xnor U4037 (N_4037,In_1418,In_620);
and U4038 (N_4038,In_2072,In_2835);
nand U4039 (N_4039,In_1477,In_1221);
or U4040 (N_4040,In_364,In_2109);
xnor U4041 (N_4041,In_2831,In_1558);
xnor U4042 (N_4042,In_1265,In_1257);
nor U4043 (N_4043,In_1920,In_94);
or U4044 (N_4044,In_2051,In_692);
nand U4045 (N_4045,In_111,In_1634);
nor U4046 (N_4046,In_972,In_2946);
or U4047 (N_4047,In_2239,In_711);
nor U4048 (N_4048,In_767,In_287);
nand U4049 (N_4049,In_2227,In_2473);
xor U4050 (N_4050,In_1709,In_343);
and U4051 (N_4051,In_1703,In_2000);
nand U4052 (N_4052,In_2556,In_1122);
or U4053 (N_4053,In_2702,In_129);
nand U4054 (N_4054,In_661,In_2665);
or U4055 (N_4055,In_2315,In_186);
or U4056 (N_4056,In_1855,In_798);
nand U4057 (N_4057,In_253,In_2378);
nand U4058 (N_4058,In_1863,In_1269);
and U4059 (N_4059,In_2382,In_17);
and U4060 (N_4060,In_2976,In_106);
nor U4061 (N_4061,In_895,In_2093);
xor U4062 (N_4062,In_1405,In_2304);
and U4063 (N_4063,In_2618,In_246);
xor U4064 (N_4064,In_867,In_2073);
nand U4065 (N_4065,In_1976,In_2073);
xor U4066 (N_4066,In_1896,In_773);
nor U4067 (N_4067,In_608,In_478);
xor U4068 (N_4068,In_1169,In_1384);
nand U4069 (N_4069,In_2025,In_844);
nor U4070 (N_4070,In_2509,In_747);
nor U4071 (N_4071,In_1523,In_2871);
xor U4072 (N_4072,In_1227,In_306);
xor U4073 (N_4073,In_2594,In_439);
xnor U4074 (N_4074,In_1301,In_1727);
or U4075 (N_4075,In_995,In_390);
or U4076 (N_4076,In_1172,In_354);
nor U4077 (N_4077,In_1804,In_407);
and U4078 (N_4078,In_1236,In_313);
nand U4079 (N_4079,In_1833,In_1102);
or U4080 (N_4080,In_469,In_1795);
nor U4081 (N_4081,In_1862,In_1526);
xor U4082 (N_4082,In_243,In_490);
nor U4083 (N_4083,In_755,In_2271);
or U4084 (N_4084,In_730,In_238);
nand U4085 (N_4085,In_2538,In_2689);
nor U4086 (N_4086,In_2044,In_149);
nor U4087 (N_4087,In_1332,In_1402);
and U4088 (N_4088,In_2604,In_663);
nand U4089 (N_4089,In_1869,In_1329);
nand U4090 (N_4090,In_307,In_2708);
nor U4091 (N_4091,In_2162,In_2104);
xor U4092 (N_4092,In_2202,In_637);
xnor U4093 (N_4093,In_2812,In_884);
nand U4094 (N_4094,In_1258,In_773);
or U4095 (N_4095,In_147,In_243);
and U4096 (N_4096,In_849,In_2591);
xnor U4097 (N_4097,In_1178,In_2849);
and U4098 (N_4098,In_178,In_2117);
and U4099 (N_4099,In_907,In_1474);
and U4100 (N_4100,In_1050,In_1197);
nor U4101 (N_4101,In_2576,In_2677);
nor U4102 (N_4102,In_2716,In_2161);
nor U4103 (N_4103,In_301,In_213);
nand U4104 (N_4104,In_2033,In_2544);
and U4105 (N_4105,In_2470,In_192);
or U4106 (N_4106,In_1348,In_562);
nand U4107 (N_4107,In_1483,In_1887);
or U4108 (N_4108,In_1841,In_2576);
nand U4109 (N_4109,In_930,In_2261);
xor U4110 (N_4110,In_1703,In_981);
nand U4111 (N_4111,In_2895,In_151);
xor U4112 (N_4112,In_2509,In_817);
nand U4113 (N_4113,In_2710,In_1498);
and U4114 (N_4114,In_625,In_2952);
nand U4115 (N_4115,In_2181,In_730);
or U4116 (N_4116,In_1897,In_1695);
nor U4117 (N_4117,In_1556,In_1621);
xnor U4118 (N_4118,In_1087,In_960);
xor U4119 (N_4119,In_1606,In_1164);
and U4120 (N_4120,In_142,In_296);
nand U4121 (N_4121,In_78,In_49);
or U4122 (N_4122,In_113,In_2425);
or U4123 (N_4123,In_2213,In_2168);
nand U4124 (N_4124,In_42,In_993);
nand U4125 (N_4125,In_1519,In_2477);
nand U4126 (N_4126,In_551,In_2568);
nand U4127 (N_4127,In_305,In_1637);
xnor U4128 (N_4128,In_2460,In_2409);
and U4129 (N_4129,In_2054,In_76);
nand U4130 (N_4130,In_139,In_765);
or U4131 (N_4131,In_557,In_378);
nor U4132 (N_4132,In_254,In_2637);
xnor U4133 (N_4133,In_2071,In_135);
nand U4134 (N_4134,In_2246,In_758);
xnor U4135 (N_4135,In_1755,In_1941);
nand U4136 (N_4136,In_2900,In_2926);
nand U4137 (N_4137,In_209,In_948);
nand U4138 (N_4138,In_668,In_1201);
nor U4139 (N_4139,In_1029,In_1253);
xor U4140 (N_4140,In_1223,In_1407);
xnor U4141 (N_4141,In_1863,In_480);
and U4142 (N_4142,In_787,In_1393);
nor U4143 (N_4143,In_1724,In_990);
xnor U4144 (N_4144,In_1640,In_2923);
and U4145 (N_4145,In_119,In_2941);
nor U4146 (N_4146,In_1256,In_1288);
nand U4147 (N_4147,In_2146,In_2498);
and U4148 (N_4148,In_2366,In_83);
nand U4149 (N_4149,In_1419,In_2638);
nor U4150 (N_4150,In_1330,In_2702);
nor U4151 (N_4151,In_284,In_2273);
nand U4152 (N_4152,In_1618,In_2202);
nand U4153 (N_4153,In_509,In_2939);
or U4154 (N_4154,In_233,In_116);
nor U4155 (N_4155,In_2695,In_1875);
xor U4156 (N_4156,In_538,In_1027);
and U4157 (N_4157,In_2465,In_669);
xor U4158 (N_4158,In_2302,In_2672);
nor U4159 (N_4159,In_143,In_2944);
or U4160 (N_4160,In_1019,In_2001);
nand U4161 (N_4161,In_1297,In_1176);
xor U4162 (N_4162,In_2869,In_2278);
nor U4163 (N_4163,In_1320,In_1814);
xor U4164 (N_4164,In_909,In_1354);
xnor U4165 (N_4165,In_160,In_1591);
xnor U4166 (N_4166,In_2349,In_2977);
nor U4167 (N_4167,In_1494,In_2811);
nor U4168 (N_4168,In_1816,In_2203);
nand U4169 (N_4169,In_1319,In_2603);
and U4170 (N_4170,In_424,In_2147);
and U4171 (N_4171,In_1567,In_295);
nand U4172 (N_4172,In_1462,In_616);
nand U4173 (N_4173,In_2692,In_2874);
nand U4174 (N_4174,In_1040,In_2477);
and U4175 (N_4175,In_2951,In_2967);
xor U4176 (N_4176,In_1261,In_865);
and U4177 (N_4177,In_2813,In_2766);
or U4178 (N_4178,In_1403,In_1372);
or U4179 (N_4179,In_487,In_977);
xor U4180 (N_4180,In_2711,In_2250);
and U4181 (N_4181,In_931,In_1625);
and U4182 (N_4182,In_2182,In_830);
nand U4183 (N_4183,In_2719,In_423);
xnor U4184 (N_4184,In_127,In_2155);
nor U4185 (N_4185,In_94,In_2605);
nor U4186 (N_4186,In_2337,In_2331);
and U4187 (N_4187,In_2147,In_1873);
nand U4188 (N_4188,In_460,In_2847);
and U4189 (N_4189,In_1506,In_1718);
and U4190 (N_4190,In_2565,In_331);
and U4191 (N_4191,In_2638,In_1780);
and U4192 (N_4192,In_78,In_1213);
or U4193 (N_4193,In_1170,In_149);
nor U4194 (N_4194,In_1035,In_483);
or U4195 (N_4195,In_541,In_2102);
and U4196 (N_4196,In_1701,In_113);
nand U4197 (N_4197,In_2544,In_2945);
or U4198 (N_4198,In_2209,In_671);
xor U4199 (N_4199,In_19,In_1455);
nor U4200 (N_4200,In_2724,In_211);
xnor U4201 (N_4201,In_1501,In_2041);
and U4202 (N_4202,In_2621,In_1314);
nor U4203 (N_4203,In_2523,In_687);
or U4204 (N_4204,In_939,In_1295);
nand U4205 (N_4205,In_385,In_1084);
and U4206 (N_4206,In_2485,In_1954);
or U4207 (N_4207,In_378,In_90);
or U4208 (N_4208,In_605,In_1439);
xnor U4209 (N_4209,In_2795,In_241);
or U4210 (N_4210,In_456,In_2414);
or U4211 (N_4211,In_2069,In_2594);
and U4212 (N_4212,In_2165,In_1635);
or U4213 (N_4213,In_867,In_1061);
xnor U4214 (N_4214,In_2142,In_851);
xnor U4215 (N_4215,In_1204,In_2295);
and U4216 (N_4216,In_2988,In_1712);
and U4217 (N_4217,In_137,In_1288);
and U4218 (N_4218,In_755,In_268);
nor U4219 (N_4219,In_1767,In_873);
or U4220 (N_4220,In_1897,In_2200);
nor U4221 (N_4221,In_309,In_1427);
nor U4222 (N_4222,In_2750,In_1860);
nor U4223 (N_4223,In_1262,In_641);
or U4224 (N_4224,In_1991,In_2628);
xor U4225 (N_4225,In_1249,In_1102);
nor U4226 (N_4226,In_34,In_477);
nor U4227 (N_4227,In_349,In_316);
and U4228 (N_4228,In_2599,In_1329);
xor U4229 (N_4229,In_1085,In_2884);
nor U4230 (N_4230,In_1027,In_1999);
or U4231 (N_4231,In_2277,In_830);
xor U4232 (N_4232,In_2273,In_346);
xnor U4233 (N_4233,In_2210,In_1164);
xor U4234 (N_4234,In_2715,In_1083);
and U4235 (N_4235,In_2295,In_21);
xor U4236 (N_4236,In_2237,In_59);
and U4237 (N_4237,In_1302,In_2282);
nor U4238 (N_4238,In_204,In_1929);
or U4239 (N_4239,In_1775,In_1699);
nand U4240 (N_4240,In_2053,In_907);
or U4241 (N_4241,In_20,In_2525);
xnor U4242 (N_4242,In_2929,In_1459);
nand U4243 (N_4243,In_235,In_1420);
xnor U4244 (N_4244,In_2487,In_1505);
and U4245 (N_4245,In_1352,In_2805);
or U4246 (N_4246,In_1389,In_208);
xnor U4247 (N_4247,In_293,In_1202);
nor U4248 (N_4248,In_1571,In_1751);
nor U4249 (N_4249,In_2396,In_620);
nor U4250 (N_4250,In_1077,In_2528);
nor U4251 (N_4251,In_1262,In_363);
and U4252 (N_4252,In_585,In_980);
nand U4253 (N_4253,In_1133,In_1912);
nand U4254 (N_4254,In_1971,In_127);
or U4255 (N_4255,In_501,In_216);
nor U4256 (N_4256,In_1536,In_2252);
xor U4257 (N_4257,In_2628,In_389);
or U4258 (N_4258,In_2723,In_1978);
nor U4259 (N_4259,In_2216,In_74);
or U4260 (N_4260,In_1260,In_1205);
nand U4261 (N_4261,In_2213,In_774);
or U4262 (N_4262,In_272,In_1622);
nor U4263 (N_4263,In_645,In_2259);
xor U4264 (N_4264,In_2801,In_2895);
nand U4265 (N_4265,In_553,In_360);
nand U4266 (N_4266,In_2331,In_1815);
and U4267 (N_4267,In_34,In_1684);
xnor U4268 (N_4268,In_2830,In_2473);
and U4269 (N_4269,In_2431,In_2933);
xor U4270 (N_4270,In_472,In_2106);
and U4271 (N_4271,In_2702,In_138);
xor U4272 (N_4272,In_242,In_767);
and U4273 (N_4273,In_2250,In_2030);
xor U4274 (N_4274,In_1964,In_2067);
nor U4275 (N_4275,In_2827,In_2425);
xnor U4276 (N_4276,In_2926,In_857);
nand U4277 (N_4277,In_2200,In_2662);
and U4278 (N_4278,In_1988,In_1663);
xnor U4279 (N_4279,In_2619,In_1107);
xor U4280 (N_4280,In_2917,In_2515);
nand U4281 (N_4281,In_766,In_882);
xnor U4282 (N_4282,In_147,In_805);
and U4283 (N_4283,In_1608,In_712);
or U4284 (N_4284,In_2980,In_146);
nor U4285 (N_4285,In_1656,In_1071);
nor U4286 (N_4286,In_894,In_2205);
xor U4287 (N_4287,In_176,In_1779);
nor U4288 (N_4288,In_634,In_1536);
nand U4289 (N_4289,In_2612,In_1202);
nor U4290 (N_4290,In_2445,In_2025);
nand U4291 (N_4291,In_432,In_2174);
or U4292 (N_4292,In_1063,In_1786);
nor U4293 (N_4293,In_2954,In_2588);
xor U4294 (N_4294,In_1561,In_1702);
nor U4295 (N_4295,In_1942,In_764);
and U4296 (N_4296,In_25,In_1072);
nor U4297 (N_4297,In_2354,In_1289);
and U4298 (N_4298,In_556,In_958);
xnor U4299 (N_4299,In_1092,In_1857);
xnor U4300 (N_4300,In_782,In_2838);
or U4301 (N_4301,In_112,In_140);
or U4302 (N_4302,In_2949,In_2506);
xnor U4303 (N_4303,In_224,In_262);
nand U4304 (N_4304,In_471,In_2803);
and U4305 (N_4305,In_1801,In_2332);
or U4306 (N_4306,In_2548,In_2963);
or U4307 (N_4307,In_1105,In_2943);
xor U4308 (N_4308,In_1926,In_413);
xor U4309 (N_4309,In_129,In_2772);
nor U4310 (N_4310,In_362,In_122);
or U4311 (N_4311,In_252,In_1422);
or U4312 (N_4312,In_1440,In_413);
and U4313 (N_4313,In_1527,In_1509);
and U4314 (N_4314,In_158,In_438);
nand U4315 (N_4315,In_1150,In_2319);
xnor U4316 (N_4316,In_1801,In_2802);
or U4317 (N_4317,In_1362,In_1880);
or U4318 (N_4318,In_1778,In_663);
nor U4319 (N_4319,In_387,In_674);
xor U4320 (N_4320,In_216,In_457);
nor U4321 (N_4321,In_924,In_866);
nor U4322 (N_4322,In_1794,In_2725);
xor U4323 (N_4323,In_1006,In_2951);
nor U4324 (N_4324,In_987,In_1522);
nor U4325 (N_4325,In_302,In_1843);
xnor U4326 (N_4326,In_2394,In_1508);
or U4327 (N_4327,In_195,In_2481);
nor U4328 (N_4328,In_195,In_2514);
or U4329 (N_4329,In_2258,In_610);
and U4330 (N_4330,In_1158,In_1336);
xor U4331 (N_4331,In_2463,In_2562);
nor U4332 (N_4332,In_1716,In_1258);
nor U4333 (N_4333,In_2062,In_2429);
and U4334 (N_4334,In_1460,In_210);
and U4335 (N_4335,In_269,In_2423);
or U4336 (N_4336,In_1843,In_1538);
nand U4337 (N_4337,In_263,In_2190);
nand U4338 (N_4338,In_1411,In_533);
xnor U4339 (N_4339,In_2665,In_2921);
xor U4340 (N_4340,In_2049,In_2089);
and U4341 (N_4341,In_1070,In_1612);
and U4342 (N_4342,In_1782,In_2549);
xnor U4343 (N_4343,In_1578,In_2526);
nand U4344 (N_4344,In_1833,In_1533);
nand U4345 (N_4345,In_1755,In_2385);
nor U4346 (N_4346,In_476,In_499);
xnor U4347 (N_4347,In_159,In_886);
xnor U4348 (N_4348,In_1728,In_207);
or U4349 (N_4349,In_1125,In_1908);
or U4350 (N_4350,In_460,In_2504);
nor U4351 (N_4351,In_163,In_2330);
nor U4352 (N_4352,In_1534,In_1394);
xnor U4353 (N_4353,In_2425,In_975);
nand U4354 (N_4354,In_1602,In_2367);
or U4355 (N_4355,In_1901,In_2466);
and U4356 (N_4356,In_2376,In_1453);
and U4357 (N_4357,In_2582,In_1589);
xnor U4358 (N_4358,In_2602,In_132);
nor U4359 (N_4359,In_2372,In_2627);
and U4360 (N_4360,In_1411,In_1272);
nand U4361 (N_4361,In_2106,In_1226);
xnor U4362 (N_4362,In_2356,In_1532);
nand U4363 (N_4363,In_2026,In_597);
and U4364 (N_4364,In_191,In_2439);
and U4365 (N_4365,In_2923,In_1362);
nor U4366 (N_4366,In_1472,In_627);
and U4367 (N_4367,In_456,In_2236);
xor U4368 (N_4368,In_445,In_2129);
and U4369 (N_4369,In_467,In_79);
or U4370 (N_4370,In_1133,In_597);
nor U4371 (N_4371,In_1882,In_1546);
nor U4372 (N_4372,In_1733,In_540);
nor U4373 (N_4373,In_2502,In_2629);
nor U4374 (N_4374,In_104,In_2636);
or U4375 (N_4375,In_363,In_331);
nor U4376 (N_4376,In_39,In_1302);
nor U4377 (N_4377,In_677,In_724);
nor U4378 (N_4378,In_2743,In_1728);
or U4379 (N_4379,In_2283,In_1096);
nor U4380 (N_4380,In_383,In_1585);
nand U4381 (N_4381,In_2208,In_2779);
nand U4382 (N_4382,In_1192,In_2389);
xnor U4383 (N_4383,In_481,In_1283);
nor U4384 (N_4384,In_2743,In_2714);
and U4385 (N_4385,In_1649,In_1304);
nand U4386 (N_4386,In_1092,In_2498);
nor U4387 (N_4387,In_1896,In_2567);
nand U4388 (N_4388,In_1274,In_278);
and U4389 (N_4389,In_2572,In_263);
or U4390 (N_4390,In_1085,In_1264);
and U4391 (N_4391,In_991,In_2942);
xor U4392 (N_4392,In_85,In_268);
nor U4393 (N_4393,In_435,In_1934);
nor U4394 (N_4394,In_2368,In_1349);
or U4395 (N_4395,In_726,In_546);
xor U4396 (N_4396,In_97,In_2588);
xor U4397 (N_4397,In_876,In_1443);
nor U4398 (N_4398,In_2348,In_152);
or U4399 (N_4399,In_1474,In_1180);
and U4400 (N_4400,In_1562,In_2112);
and U4401 (N_4401,In_177,In_1181);
and U4402 (N_4402,In_2035,In_2444);
or U4403 (N_4403,In_166,In_1810);
nor U4404 (N_4404,In_1928,In_106);
and U4405 (N_4405,In_1995,In_74);
or U4406 (N_4406,In_1720,In_2572);
and U4407 (N_4407,In_1587,In_1640);
nor U4408 (N_4408,In_2634,In_395);
nand U4409 (N_4409,In_1294,In_998);
nand U4410 (N_4410,In_672,In_541);
or U4411 (N_4411,In_1832,In_790);
nor U4412 (N_4412,In_2175,In_38);
and U4413 (N_4413,In_2893,In_746);
or U4414 (N_4414,In_525,In_1099);
nor U4415 (N_4415,In_584,In_2091);
nor U4416 (N_4416,In_2313,In_856);
and U4417 (N_4417,In_2594,In_419);
or U4418 (N_4418,In_1640,In_1856);
nor U4419 (N_4419,In_926,In_2382);
nand U4420 (N_4420,In_519,In_2081);
and U4421 (N_4421,In_2428,In_1085);
and U4422 (N_4422,In_2145,In_1186);
nand U4423 (N_4423,In_1573,In_826);
or U4424 (N_4424,In_220,In_2313);
and U4425 (N_4425,In_2478,In_2641);
nor U4426 (N_4426,In_553,In_2358);
or U4427 (N_4427,In_94,In_2905);
or U4428 (N_4428,In_567,In_1012);
nor U4429 (N_4429,In_2596,In_1787);
xnor U4430 (N_4430,In_1521,In_2230);
and U4431 (N_4431,In_2603,In_1802);
nand U4432 (N_4432,In_1460,In_2362);
xor U4433 (N_4433,In_1770,In_2393);
nand U4434 (N_4434,In_1678,In_1429);
nand U4435 (N_4435,In_2345,In_209);
nand U4436 (N_4436,In_2588,In_195);
and U4437 (N_4437,In_2546,In_2275);
and U4438 (N_4438,In_2533,In_1862);
xor U4439 (N_4439,In_688,In_2567);
nand U4440 (N_4440,In_2094,In_2973);
and U4441 (N_4441,In_2448,In_2483);
and U4442 (N_4442,In_51,In_2917);
nand U4443 (N_4443,In_2975,In_356);
xnor U4444 (N_4444,In_1610,In_1702);
nand U4445 (N_4445,In_86,In_2297);
and U4446 (N_4446,In_2432,In_1253);
and U4447 (N_4447,In_1896,In_457);
nand U4448 (N_4448,In_60,In_1655);
or U4449 (N_4449,In_370,In_474);
or U4450 (N_4450,In_364,In_742);
nand U4451 (N_4451,In_1528,In_508);
nor U4452 (N_4452,In_2603,In_2428);
nand U4453 (N_4453,In_1579,In_1714);
nand U4454 (N_4454,In_1257,In_1998);
and U4455 (N_4455,In_799,In_2572);
nand U4456 (N_4456,In_1582,In_2635);
nand U4457 (N_4457,In_2621,In_210);
xnor U4458 (N_4458,In_217,In_2849);
nand U4459 (N_4459,In_1268,In_836);
nor U4460 (N_4460,In_1036,In_2569);
nor U4461 (N_4461,In_913,In_19);
nand U4462 (N_4462,In_827,In_2524);
nand U4463 (N_4463,In_1549,In_1292);
nor U4464 (N_4464,In_2749,In_1741);
and U4465 (N_4465,In_2283,In_1025);
nor U4466 (N_4466,In_2000,In_1378);
nor U4467 (N_4467,In_1729,In_2091);
and U4468 (N_4468,In_667,In_2282);
or U4469 (N_4469,In_1653,In_967);
xor U4470 (N_4470,In_934,In_1342);
nor U4471 (N_4471,In_2120,In_1977);
or U4472 (N_4472,In_1569,In_1385);
nand U4473 (N_4473,In_2680,In_738);
nand U4474 (N_4474,In_2026,In_1705);
nor U4475 (N_4475,In_806,In_766);
nand U4476 (N_4476,In_1546,In_2335);
or U4477 (N_4477,In_1015,In_2700);
nor U4478 (N_4478,In_536,In_2367);
or U4479 (N_4479,In_731,In_1608);
nor U4480 (N_4480,In_1409,In_2281);
and U4481 (N_4481,In_725,In_857);
xnor U4482 (N_4482,In_2996,In_2070);
nand U4483 (N_4483,In_859,In_2113);
xor U4484 (N_4484,In_625,In_982);
and U4485 (N_4485,In_1220,In_541);
and U4486 (N_4486,In_1890,In_1370);
or U4487 (N_4487,In_2271,In_174);
or U4488 (N_4488,In_2509,In_600);
and U4489 (N_4489,In_497,In_414);
xnor U4490 (N_4490,In_1730,In_1690);
nor U4491 (N_4491,In_571,In_1567);
and U4492 (N_4492,In_2194,In_2131);
nor U4493 (N_4493,In_1715,In_293);
or U4494 (N_4494,In_2521,In_571);
nand U4495 (N_4495,In_1159,In_1308);
xor U4496 (N_4496,In_2492,In_2643);
xnor U4497 (N_4497,In_2278,In_2765);
and U4498 (N_4498,In_1640,In_1231);
xor U4499 (N_4499,In_2943,In_2369);
nand U4500 (N_4500,In_2473,In_2016);
nor U4501 (N_4501,In_2732,In_2517);
and U4502 (N_4502,In_1653,In_308);
and U4503 (N_4503,In_857,In_341);
nor U4504 (N_4504,In_2106,In_810);
nand U4505 (N_4505,In_1716,In_9);
and U4506 (N_4506,In_1205,In_267);
nand U4507 (N_4507,In_2518,In_623);
nand U4508 (N_4508,In_1742,In_11);
nor U4509 (N_4509,In_1257,In_2533);
nor U4510 (N_4510,In_306,In_2294);
nor U4511 (N_4511,In_62,In_2535);
xnor U4512 (N_4512,In_2419,In_1023);
or U4513 (N_4513,In_2125,In_2947);
and U4514 (N_4514,In_859,In_1265);
or U4515 (N_4515,In_2542,In_1563);
nand U4516 (N_4516,In_1539,In_1624);
or U4517 (N_4517,In_1852,In_2179);
nand U4518 (N_4518,In_2809,In_1743);
xor U4519 (N_4519,In_71,In_2040);
and U4520 (N_4520,In_2365,In_2458);
xnor U4521 (N_4521,In_2862,In_2617);
nor U4522 (N_4522,In_2186,In_584);
and U4523 (N_4523,In_2817,In_752);
xnor U4524 (N_4524,In_2621,In_1259);
nor U4525 (N_4525,In_1227,In_1084);
nor U4526 (N_4526,In_1760,In_2195);
nor U4527 (N_4527,In_2895,In_1307);
and U4528 (N_4528,In_36,In_963);
nor U4529 (N_4529,In_1092,In_299);
and U4530 (N_4530,In_473,In_676);
nor U4531 (N_4531,In_2063,In_2574);
or U4532 (N_4532,In_676,In_1272);
and U4533 (N_4533,In_975,In_28);
nand U4534 (N_4534,In_2598,In_2280);
nor U4535 (N_4535,In_1475,In_1739);
or U4536 (N_4536,In_211,In_1696);
or U4537 (N_4537,In_2220,In_1215);
nor U4538 (N_4538,In_1240,In_2933);
or U4539 (N_4539,In_111,In_1643);
xnor U4540 (N_4540,In_418,In_2111);
and U4541 (N_4541,In_784,In_1532);
xnor U4542 (N_4542,In_1591,In_1932);
xnor U4543 (N_4543,In_141,In_1832);
and U4544 (N_4544,In_566,In_701);
xnor U4545 (N_4545,In_1826,In_769);
xor U4546 (N_4546,In_771,In_2785);
or U4547 (N_4547,In_1139,In_1820);
and U4548 (N_4548,In_980,In_1685);
xor U4549 (N_4549,In_2042,In_2242);
xor U4550 (N_4550,In_1172,In_1453);
nand U4551 (N_4551,In_2212,In_782);
nand U4552 (N_4552,In_2482,In_2961);
nand U4553 (N_4553,In_2679,In_850);
nor U4554 (N_4554,In_28,In_316);
xor U4555 (N_4555,In_2484,In_521);
nand U4556 (N_4556,In_2947,In_304);
and U4557 (N_4557,In_2778,In_603);
and U4558 (N_4558,In_2386,In_26);
xor U4559 (N_4559,In_1424,In_1671);
nor U4560 (N_4560,In_451,In_1326);
and U4561 (N_4561,In_2607,In_534);
or U4562 (N_4562,In_937,In_110);
and U4563 (N_4563,In_1508,In_1270);
or U4564 (N_4564,In_1393,In_2416);
or U4565 (N_4565,In_502,In_1886);
xor U4566 (N_4566,In_1011,In_2815);
and U4567 (N_4567,In_2540,In_2001);
or U4568 (N_4568,In_2668,In_2959);
or U4569 (N_4569,In_585,In_2270);
xor U4570 (N_4570,In_2201,In_1094);
and U4571 (N_4571,In_2475,In_1164);
xnor U4572 (N_4572,In_135,In_927);
or U4573 (N_4573,In_927,In_267);
nor U4574 (N_4574,In_538,In_2485);
or U4575 (N_4575,In_2665,In_1171);
nand U4576 (N_4576,In_1808,In_2052);
nor U4577 (N_4577,In_853,In_1669);
nor U4578 (N_4578,In_153,In_1278);
nand U4579 (N_4579,In_244,In_1095);
nand U4580 (N_4580,In_2294,In_2604);
nand U4581 (N_4581,In_2782,In_1471);
or U4582 (N_4582,In_920,In_1766);
and U4583 (N_4583,In_2273,In_1047);
and U4584 (N_4584,In_1199,In_2716);
and U4585 (N_4585,In_1431,In_104);
nor U4586 (N_4586,In_2189,In_2555);
nand U4587 (N_4587,In_2827,In_2679);
xnor U4588 (N_4588,In_136,In_1527);
or U4589 (N_4589,In_2782,In_682);
xor U4590 (N_4590,In_1612,In_196);
nand U4591 (N_4591,In_2423,In_1949);
or U4592 (N_4592,In_2087,In_20);
nor U4593 (N_4593,In_195,In_1459);
and U4594 (N_4594,In_804,In_828);
xor U4595 (N_4595,In_184,In_789);
nor U4596 (N_4596,In_1259,In_2518);
and U4597 (N_4597,In_1375,In_1619);
nor U4598 (N_4598,In_778,In_464);
nor U4599 (N_4599,In_555,In_1933);
nor U4600 (N_4600,In_868,In_644);
or U4601 (N_4601,In_2522,In_2109);
nor U4602 (N_4602,In_2031,In_2633);
and U4603 (N_4603,In_224,In_1122);
nand U4604 (N_4604,In_1711,In_1648);
nand U4605 (N_4605,In_2913,In_1486);
and U4606 (N_4606,In_1938,In_1761);
nand U4607 (N_4607,In_889,In_2960);
and U4608 (N_4608,In_2917,In_2961);
and U4609 (N_4609,In_1364,In_2455);
xnor U4610 (N_4610,In_954,In_1996);
or U4611 (N_4611,In_1177,In_2509);
xnor U4612 (N_4612,In_2685,In_1287);
and U4613 (N_4613,In_276,In_682);
xnor U4614 (N_4614,In_444,In_136);
nand U4615 (N_4615,In_1211,In_1135);
and U4616 (N_4616,In_2952,In_2125);
nor U4617 (N_4617,In_55,In_2875);
nor U4618 (N_4618,In_463,In_300);
nor U4619 (N_4619,In_450,In_2008);
and U4620 (N_4620,In_1161,In_2995);
or U4621 (N_4621,In_1412,In_2266);
nor U4622 (N_4622,In_2236,In_614);
or U4623 (N_4623,In_1566,In_796);
nor U4624 (N_4624,In_1201,In_1057);
xor U4625 (N_4625,In_2222,In_969);
nand U4626 (N_4626,In_1720,In_2833);
and U4627 (N_4627,In_1338,In_2932);
nor U4628 (N_4628,In_974,In_1496);
xnor U4629 (N_4629,In_2397,In_1611);
xor U4630 (N_4630,In_2122,In_528);
and U4631 (N_4631,In_1268,In_1532);
and U4632 (N_4632,In_236,In_187);
and U4633 (N_4633,In_2280,In_2881);
xor U4634 (N_4634,In_1040,In_2141);
or U4635 (N_4635,In_1894,In_2638);
nor U4636 (N_4636,In_2124,In_2071);
nand U4637 (N_4637,In_2681,In_2036);
or U4638 (N_4638,In_1745,In_1008);
nand U4639 (N_4639,In_1078,In_439);
and U4640 (N_4640,In_352,In_1003);
or U4641 (N_4641,In_537,In_481);
nor U4642 (N_4642,In_532,In_565);
nand U4643 (N_4643,In_726,In_887);
or U4644 (N_4644,In_338,In_619);
xor U4645 (N_4645,In_1553,In_1164);
nor U4646 (N_4646,In_2773,In_975);
nand U4647 (N_4647,In_571,In_1719);
xnor U4648 (N_4648,In_2075,In_0);
xnor U4649 (N_4649,In_2090,In_1805);
or U4650 (N_4650,In_2891,In_96);
and U4651 (N_4651,In_310,In_1796);
xnor U4652 (N_4652,In_858,In_2881);
or U4653 (N_4653,In_838,In_697);
xnor U4654 (N_4654,In_1241,In_586);
nor U4655 (N_4655,In_2715,In_42);
nor U4656 (N_4656,In_2215,In_341);
and U4657 (N_4657,In_543,In_1336);
or U4658 (N_4658,In_2774,In_583);
and U4659 (N_4659,In_424,In_2781);
nor U4660 (N_4660,In_2778,In_2882);
nand U4661 (N_4661,In_560,In_1852);
and U4662 (N_4662,In_446,In_93);
nand U4663 (N_4663,In_209,In_972);
nor U4664 (N_4664,In_100,In_1693);
and U4665 (N_4665,In_1810,In_1031);
and U4666 (N_4666,In_2406,In_1426);
xnor U4667 (N_4667,In_2244,In_465);
and U4668 (N_4668,In_1804,In_1935);
nor U4669 (N_4669,In_2510,In_93);
or U4670 (N_4670,In_2564,In_743);
or U4671 (N_4671,In_89,In_2322);
and U4672 (N_4672,In_2996,In_2648);
xnor U4673 (N_4673,In_2933,In_2508);
nor U4674 (N_4674,In_2295,In_594);
xor U4675 (N_4675,In_730,In_702);
nand U4676 (N_4676,In_1929,In_2634);
nand U4677 (N_4677,In_1740,In_2774);
and U4678 (N_4678,In_1547,In_389);
xnor U4679 (N_4679,In_1176,In_2660);
or U4680 (N_4680,In_298,In_1143);
or U4681 (N_4681,In_0,In_1425);
xnor U4682 (N_4682,In_845,In_1350);
or U4683 (N_4683,In_2286,In_594);
or U4684 (N_4684,In_646,In_2673);
nor U4685 (N_4685,In_2141,In_1203);
and U4686 (N_4686,In_441,In_68);
nand U4687 (N_4687,In_1449,In_538);
and U4688 (N_4688,In_1518,In_1993);
or U4689 (N_4689,In_1120,In_887);
or U4690 (N_4690,In_1604,In_996);
nand U4691 (N_4691,In_204,In_525);
nor U4692 (N_4692,In_511,In_1316);
or U4693 (N_4693,In_1615,In_164);
or U4694 (N_4694,In_1021,In_1551);
nor U4695 (N_4695,In_1807,In_2338);
nor U4696 (N_4696,In_1065,In_774);
xor U4697 (N_4697,In_994,In_1035);
and U4698 (N_4698,In_2124,In_1587);
xor U4699 (N_4699,In_1245,In_465);
or U4700 (N_4700,In_1398,In_301);
and U4701 (N_4701,In_2340,In_446);
and U4702 (N_4702,In_16,In_1039);
or U4703 (N_4703,In_563,In_87);
nand U4704 (N_4704,In_2596,In_2546);
and U4705 (N_4705,In_208,In_2557);
nor U4706 (N_4706,In_2297,In_1207);
or U4707 (N_4707,In_2117,In_1843);
nor U4708 (N_4708,In_2319,In_435);
and U4709 (N_4709,In_997,In_2665);
or U4710 (N_4710,In_794,In_2884);
nor U4711 (N_4711,In_362,In_2381);
and U4712 (N_4712,In_1013,In_914);
nor U4713 (N_4713,In_2149,In_180);
nand U4714 (N_4714,In_266,In_1358);
nor U4715 (N_4715,In_349,In_2843);
nor U4716 (N_4716,In_1116,In_1222);
nor U4717 (N_4717,In_1670,In_1523);
and U4718 (N_4718,In_1118,In_2832);
nand U4719 (N_4719,In_2613,In_491);
or U4720 (N_4720,In_776,In_2823);
xnor U4721 (N_4721,In_709,In_1864);
nor U4722 (N_4722,In_434,In_2253);
and U4723 (N_4723,In_902,In_2617);
or U4724 (N_4724,In_64,In_2051);
and U4725 (N_4725,In_338,In_583);
or U4726 (N_4726,In_349,In_453);
nand U4727 (N_4727,In_2566,In_1800);
nor U4728 (N_4728,In_2764,In_2672);
nor U4729 (N_4729,In_1386,In_2414);
nand U4730 (N_4730,In_2458,In_1904);
and U4731 (N_4731,In_2,In_1376);
or U4732 (N_4732,In_1112,In_2868);
nand U4733 (N_4733,In_1844,In_1202);
and U4734 (N_4734,In_981,In_741);
xnor U4735 (N_4735,In_2144,In_2819);
or U4736 (N_4736,In_2030,In_27);
nand U4737 (N_4737,In_1681,In_727);
nand U4738 (N_4738,In_2040,In_774);
or U4739 (N_4739,In_153,In_1877);
and U4740 (N_4740,In_2844,In_2295);
nand U4741 (N_4741,In_2019,In_1713);
or U4742 (N_4742,In_870,In_264);
and U4743 (N_4743,In_2727,In_1946);
and U4744 (N_4744,In_316,In_1719);
nor U4745 (N_4745,In_41,In_576);
xnor U4746 (N_4746,In_1803,In_986);
or U4747 (N_4747,In_1303,In_841);
and U4748 (N_4748,In_487,In_2726);
and U4749 (N_4749,In_1493,In_2440);
xnor U4750 (N_4750,In_2042,In_153);
or U4751 (N_4751,In_1787,In_1722);
or U4752 (N_4752,In_330,In_1901);
and U4753 (N_4753,In_2907,In_2275);
or U4754 (N_4754,In_236,In_1466);
and U4755 (N_4755,In_970,In_566);
xnor U4756 (N_4756,In_2754,In_1159);
xnor U4757 (N_4757,In_2006,In_2826);
nor U4758 (N_4758,In_1591,In_363);
or U4759 (N_4759,In_218,In_1892);
or U4760 (N_4760,In_1839,In_618);
or U4761 (N_4761,In_1602,In_2716);
or U4762 (N_4762,In_2990,In_2247);
nor U4763 (N_4763,In_323,In_1794);
nor U4764 (N_4764,In_739,In_2535);
nand U4765 (N_4765,In_2359,In_90);
xor U4766 (N_4766,In_2144,In_283);
nor U4767 (N_4767,In_2965,In_2241);
or U4768 (N_4768,In_2712,In_2114);
nor U4769 (N_4769,In_2519,In_714);
nor U4770 (N_4770,In_1744,In_1286);
and U4771 (N_4771,In_421,In_698);
and U4772 (N_4772,In_1790,In_695);
nor U4773 (N_4773,In_2315,In_1731);
and U4774 (N_4774,In_910,In_1457);
xor U4775 (N_4775,In_367,In_941);
nor U4776 (N_4776,In_66,In_1402);
xor U4777 (N_4777,In_1417,In_1770);
nand U4778 (N_4778,In_44,In_1162);
and U4779 (N_4779,In_2039,In_1529);
and U4780 (N_4780,In_1129,In_1757);
nor U4781 (N_4781,In_1410,In_1075);
and U4782 (N_4782,In_173,In_944);
and U4783 (N_4783,In_1725,In_1463);
and U4784 (N_4784,In_355,In_2934);
nand U4785 (N_4785,In_1175,In_1396);
nor U4786 (N_4786,In_1662,In_2739);
nor U4787 (N_4787,In_1816,In_1523);
xor U4788 (N_4788,In_1981,In_1173);
nand U4789 (N_4789,In_2199,In_2710);
nand U4790 (N_4790,In_1728,In_447);
xor U4791 (N_4791,In_1232,In_1751);
nor U4792 (N_4792,In_2754,In_678);
and U4793 (N_4793,In_1984,In_1656);
or U4794 (N_4794,In_734,In_2924);
nor U4795 (N_4795,In_683,In_1430);
nand U4796 (N_4796,In_323,In_2497);
and U4797 (N_4797,In_2905,In_2520);
or U4798 (N_4798,In_2125,In_1829);
xor U4799 (N_4799,In_792,In_2339);
and U4800 (N_4800,In_1008,In_1223);
nand U4801 (N_4801,In_2074,In_2281);
nand U4802 (N_4802,In_50,In_2434);
xor U4803 (N_4803,In_2866,In_1663);
or U4804 (N_4804,In_1669,In_2052);
and U4805 (N_4805,In_2923,In_1335);
or U4806 (N_4806,In_1089,In_1814);
nand U4807 (N_4807,In_1489,In_1824);
nor U4808 (N_4808,In_1487,In_2528);
or U4809 (N_4809,In_554,In_378);
or U4810 (N_4810,In_459,In_2327);
nand U4811 (N_4811,In_1731,In_2456);
or U4812 (N_4812,In_2544,In_2345);
or U4813 (N_4813,In_2367,In_623);
or U4814 (N_4814,In_2981,In_2695);
or U4815 (N_4815,In_1069,In_1731);
nor U4816 (N_4816,In_1293,In_73);
or U4817 (N_4817,In_389,In_2688);
xnor U4818 (N_4818,In_2371,In_129);
xor U4819 (N_4819,In_1555,In_2585);
xor U4820 (N_4820,In_1063,In_2048);
nor U4821 (N_4821,In_1121,In_289);
nor U4822 (N_4822,In_121,In_1231);
xor U4823 (N_4823,In_2540,In_2458);
or U4824 (N_4824,In_2077,In_1588);
xnor U4825 (N_4825,In_2324,In_1806);
xor U4826 (N_4826,In_328,In_2745);
and U4827 (N_4827,In_2326,In_2452);
xnor U4828 (N_4828,In_2206,In_388);
nor U4829 (N_4829,In_1097,In_1566);
nand U4830 (N_4830,In_616,In_398);
xnor U4831 (N_4831,In_2608,In_2376);
and U4832 (N_4832,In_1942,In_2915);
nand U4833 (N_4833,In_2201,In_837);
or U4834 (N_4834,In_2301,In_1036);
nand U4835 (N_4835,In_1914,In_2415);
nor U4836 (N_4836,In_2871,In_2210);
and U4837 (N_4837,In_1515,In_195);
and U4838 (N_4838,In_306,In_2056);
or U4839 (N_4839,In_470,In_2533);
nor U4840 (N_4840,In_2751,In_511);
nand U4841 (N_4841,In_1471,In_1259);
or U4842 (N_4842,In_175,In_2390);
or U4843 (N_4843,In_2108,In_2460);
and U4844 (N_4844,In_906,In_2460);
nand U4845 (N_4845,In_42,In_183);
xor U4846 (N_4846,In_2025,In_1767);
nand U4847 (N_4847,In_592,In_1184);
and U4848 (N_4848,In_1558,In_758);
or U4849 (N_4849,In_2138,In_2917);
nor U4850 (N_4850,In_1798,In_2131);
or U4851 (N_4851,In_2839,In_72);
or U4852 (N_4852,In_2527,In_107);
nor U4853 (N_4853,In_1736,In_2487);
xor U4854 (N_4854,In_1863,In_704);
and U4855 (N_4855,In_609,In_585);
and U4856 (N_4856,In_2397,In_1074);
xnor U4857 (N_4857,In_1950,In_2589);
xnor U4858 (N_4858,In_1158,In_1747);
nor U4859 (N_4859,In_627,In_1153);
or U4860 (N_4860,In_2381,In_1658);
xor U4861 (N_4861,In_1436,In_2762);
nor U4862 (N_4862,In_420,In_2886);
and U4863 (N_4863,In_1578,In_861);
xnor U4864 (N_4864,In_2547,In_2390);
nand U4865 (N_4865,In_1037,In_1882);
xor U4866 (N_4866,In_2515,In_442);
nand U4867 (N_4867,In_2790,In_17);
xnor U4868 (N_4868,In_2623,In_139);
xnor U4869 (N_4869,In_2584,In_2185);
nor U4870 (N_4870,In_342,In_1891);
nor U4871 (N_4871,In_2878,In_2744);
nand U4872 (N_4872,In_2663,In_2120);
nand U4873 (N_4873,In_2488,In_771);
nand U4874 (N_4874,In_2051,In_2236);
nor U4875 (N_4875,In_2175,In_1660);
xor U4876 (N_4876,In_2053,In_2197);
nand U4877 (N_4877,In_1618,In_2504);
or U4878 (N_4878,In_281,In_2581);
and U4879 (N_4879,In_1334,In_2781);
nor U4880 (N_4880,In_2260,In_235);
or U4881 (N_4881,In_364,In_2002);
nor U4882 (N_4882,In_1440,In_2682);
xnor U4883 (N_4883,In_1750,In_1581);
nor U4884 (N_4884,In_920,In_40);
and U4885 (N_4885,In_236,In_2390);
nand U4886 (N_4886,In_1895,In_1454);
nand U4887 (N_4887,In_2780,In_1198);
nor U4888 (N_4888,In_2149,In_1016);
nand U4889 (N_4889,In_558,In_668);
and U4890 (N_4890,In_2703,In_2660);
and U4891 (N_4891,In_188,In_2407);
and U4892 (N_4892,In_1236,In_1185);
nor U4893 (N_4893,In_88,In_2037);
xor U4894 (N_4894,In_573,In_1899);
or U4895 (N_4895,In_2380,In_850);
or U4896 (N_4896,In_932,In_606);
or U4897 (N_4897,In_1323,In_634);
xnor U4898 (N_4898,In_2617,In_2751);
or U4899 (N_4899,In_259,In_970);
nor U4900 (N_4900,In_1967,In_2528);
xor U4901 (N_4901,In_2057,In_1737);
or U4902 (N_4902,In_1414,In_302);
xnor U4903 (N_4903,In_2492,In_213);
xor U4904 (N_4904,In_1931,In_764);
xor U4905 (N_4905,In_2320,In_1283);
or U4906 (N_4906,In_1094,In_2418);
nand U4907 (N_4907,In_61,In_2651);
nor U4908 (N_4908,In_465,In_1215);
nand U4909 (N_4909,In_196,In_827);
or U4910 (N_4910,In_1696,In_2478);
nand U4911 (N_4911,In_2588,In_1564);
or U4912 (N_4912,In_410,In_227);
nand U4913 (N_4913,In_2651,In_2710);
nand U4914 (N_4914,In_2088,In_1221);
and U4915 (N_4915,In_1361,In_1115);
and U4916 (N_4916,In_132,In_1176);
nor U4917 (N_4917,In_73,In_2596);
nor U4918 (N_4918,In_1429,In_1996);
nand U4919 (N_4919,In_2406,In_1260);
xnor U4920 (N_4920,In_1266,In_1776);
or U4921 (N_4921,In_810,In_373);
and U4922 (N_4922,In_2007,In_1430);
nor U4923 (N_4923,In_517,In_1734);
nand U4924 (N_4924,In_1612,In_415);
and U4925 (N_4925,In_2285,In_1282);
or U4926 (N_4926,In_1725,In_2965);
nand U4927 (N_4927,In_2509,In_2073);
and U4928 (N_4928,In_1983,In_1441);
or U4929 (N_4929,In_1602,In_479);
or U4930 (N_4930,In_2731,In_714);
nor U4931 (N_4931,In_2478,In_1889);
and U4932 (N_4932,In_1844,In_2823);
xor U4933 (N_4933,In_1380,In_1767);
nor U4934 (N_4934,In_481,In_606);
xnor U4935 (N_4935,In_2068,In_738);
nand U4936 (N_4936,In_1897,In_22);
and U4937 (N_4937,In_560,In_535);
or U4938 (N_4938,In_308,In_2707);
xor U4939 (N_4939,In_76,In_1520);
nor U4940 (N_4940,In_1291,In_2415);
xnor U4941 (N_4941,In_898,In_1954);
or U4942 (N_4942,In_2549,In_1235);
nand U4943 (N_4943,In_1802,In_282);
nor U4944 (N_4944,In_522,In_2410);
or U4945 (N_4945,In_1796,In_2517);
nor U4946 (N_4946,In_2031,In_1459);
xor U4947 (N_4947,In_2880,In_2719);
nor U4948 (N_4948,In_2804,In_2597);
nor U4949 (N_4949,In_776,In_442);
nor U4950 (N_4950,In_748,In_1757);
nor U4951 (N_4951,In_2694,In_2529);
nand U4952 (N_4952,In_208,In_2914);
nor U4953 (N_4953,In_712,In_1083);
nor U4954 (N_4954,In_244,In_1061);
or U4955 (N_4955,In_972,In_1737);
or U4956 (N_4956,In_207,In_1219);
or U4957 (N_4957,In_1657,In_2784);
and U4958 (N_4958,In_904,In_2476);
and U4959 (N_4959,In_1762,In_2229);
nor U4960 (N_4960,In_286,In_443);
xnor U4961 (N_4961,In_466,In_2606);
nand U4962 (N_4962,In_1395,In_1171);
nand U4963 (N_4963,In_756,In_2209);
and U4964 (N_4964,In_1068,In_189);
nor U4965 (N_4965,In_1730,In_354);
nand U4966 (N_4966,In_388,In_1271);
or U4967 (N_4967,In_1128,In_1484);
xnor U4968 (N_4968,In_66,In_1995);
xnor U4969 (N_4969,In_1777,In_1244);
xnor U4970 (N_4970,In_945,In_80);
nor U4971 (N_4971,In_280,In_1394);
nor U4972 (N_4972,In_321,In_1373);
xnor U4973 (N_4973,In_2369,In_1243);
xnor U4974 (N_4974,In_1295,In_1745);
or U4975 (N_4975,In_349,In_1907);
nor U4976 (N_4976,In_1025,In_122);
xor U4977 (N_4977,In_433,In_1922);
nand U4978 (N_4978,In_759,In_2595);
nand U4979 (N_4979,In_411,In_2929);
and U4980 (N_4980,In_786,In_2702);
nand U4981 (N_4981,In_486,In_2916);
and U4982 (N_4982,In_1212,In_2953);
xnor U4983 (N_4983,In_1208,In_870);
nor U4984 (N_4984,In_2175,In_1740);
nor U4985 (N_4985,In_2527,In_514);
and U4986 (N_4986,In_1796,In_1226);
xnor U4987 (N_4987,In_748,In_1175);
and U4988 (N_4988,In_1767,In_2103);
nor U4989 (N_4989,In_2325,In_2346);
or U4990 (N_4990,In_303,In_2504);
and U4991 (N_4991,In_1236,In_2510);
nand U4992 (N_4992,In_856,In_48);
or U4993 (N_4993,In_369,In_2281);
xor U4994 (N_4994,In_2265,In_693);
and U4995 (N_4995,In_550,In_1135);
nor U4996 (N_4996,In_2864,In_1133);
and U4997 (N_4997,In_1195,In_713);
and U4998 (N_4998,In_2834,In_152);
nor U4999 (N_4999,In_1526,In_2286);
nor U5000 (N_5000,N_4759,N_2315);
and U5001 (N_5001,N_1745,N_3283);
xnor U5002 (N_5002,N_4163,N_3468);
and U5003 (N_5003,N_3389,N_202);
nand U5004 (N_5004,N_3904,N_2793);
and U5005 (N_5005,N_4584,N_820);
nand U5006 (N_5006,N_280,N_1198);
nand U5007 (N_5007,N_52,N_2305);
or U5008 (N_5008,N_2894,N_767);
or U5009 (N_5009,N_214,N_3368);
or U5010 (N_5010,N_3295,N_3620);
nor U5011 (N_5011,N_3116,N_1061);
and U5012 (N_5012,N_3692,N_35);
xor U5013 (N_5013,N_4213,N_3293);
nand U5014 (N_5014,N_4736,N_3621);
and U5015 (N_5015,N_2631,N_2366);
nor U5016 (N_5016,N_4954,N_194);
xor U5017 (N_5017,N_3910,N_1640);
and U5018 (N_5018,N_271,N_1242);
or U5019 (N_5019,N_1513,N_2750);
nand U5020 (N_5020,N_4800,N_903);
nand U5021 (N_5021,N_3960,N_1387);
xnor U5022 (N_5022,N_2938,N_3770);
and U5023 (N_5023,N_3322,N_349);
nor U5024 (N_5024,N_4534,N_1441);
and U5025 (N_5025,N_4009,N_1757);
nand U5026 (N_5026,N_1589,N_4106);
and U5027 (N_5027,N_3426,N_4822);
or U5028 (N_5028,N_1069,N_838);
nor U5029 (N_5029,N_1841,N_4606);
nand U5030 (N_5030,N_1778,N_23);
nor U5031 (N_5031,N_4735,N_2286);
nand U5032 (N_5032,N_219,N_4644);
or U5033 (N_5033,N_4483,N_2173);
nor U5034 (N_5034,N_4064,N_2650);
or U5035 (N_5035,N_2091,N_4783);
xnor U5036 (N_5036,N_646,N_3164);
or U5037 (N_5037,N_147,N_3518);
nand U5038 (N_5038,N_2838,N_3577);
and U5039 (N_5039,N_2893,N_1001);
nor U5040 (N_5040,N_2960,N_2684);
and U5041 (N_5041,N_1569,N_4400);
and U5042 (N_5042,N_910,N_3098);
nor U5043 (N_5043,N_243,N_282);
xor U5044 (N_5044,N_63,N_1895);
or U5045 (N_5045,N_3027,N_1758);
nor U5046 (N_5046,N_2826,N_1169);
and U5047 (N_5047,N_4149,N_990);
nand U5048 (N_5048,N_3392,N_3729);
nand U5049 (N_5049,N_2240,N_2600);
and U5050 (N_5050,N_2117,N_1385);
nand U5051 (N_5051,N_2168,N_4890);
nand U5052 (N_5052,N_2379,N_4674);
and U5053 (N_5053,N_3439,N_539);
nor U5054 (N_5054,N_2055,N_4608);
and U5055 (N_5055,N_432,N_3929);
or U5056 (N_5056,N_4443,N_1455);
and U5057 (N_5057,N_489,N_2234);
nor U5058 (N_5058,N_1431,N_2428);
nor U5059 (N_5059,N_288,N_1178);
nand U5060 (N_5060,N_3131,N_2903);
nor U5061 (N_5061,N_3859,N_4567);
nor U5062 (N_5062,N_2220,N_4270);
or U5063 (N_5063,N_2763,N_3466);
and U5064 (N_5064,N_2436,N_2962);
nor U5065 (N_5065,N_811,N_1678);
and U5066 (N_5066,N_2023,N_3473);
and U5067 (N_5067,N_40,N_2567);
or U5068 (N_5068,N_1496,N_4044);
and U5069 (N_5069,N_203,N_926);
xor U5070 (N_5070,N_3998,N_2710);
or U5071 (N_5071,N_77,N_4175);
nor U5072 (N_5072,N_3252,N_18);
or U5073 (N_5073,N_1764,N_1383);
xnor U5074 (N_5074,N_4335,N_4792);
nand U5075 (N_5075,N_4376,N_200);
or U5076 (N_5076,N_1624,N_4277);
xnor U5077 (N_5077,N_4027,N_1942);
and U5078 (N_5078,N_2515,N_3064);
nand U5079 (N_5079,N_3532,N_4087);
nand U5080 (N_5080,N_4258,N_4439);
nor U5081 (N_5081,N_1480,N_852);
xor U5082 (N_5082,N_3105,N_2804);
nand U5083 (N_5083,N_2657,N_2491);
and U5084 (N_5084,N_30,N_380);
and U5085 (N_5085,N_325,N_4767);
nor U5086 (N_5086,N_2176,N_1988);
nor U5087 (N_5087,N_1986,N_4746);
and U5088 (N_5088,N_163,N_2261);
or U5089 (N_5089,N_2919,N_1313);
xor U5090 (N_5090,N_2051,N_1978);
xor U5091 (N_5091,N_2061,N_4070);
nor U5092 (N_5092,N_2655,N_3488);
xnor U5093 (N_5093,N_130,N_2866);
and U5094 (N_5094,N_3442,N_3284);
and U5095 (N_5095,N_1092,N_4701);
xor U5096 (N_5096,N_4726,N_4816);
nor U5097 (N_5097,N_3206,N_2264);
and U5098 (N_5098,N_4117,N_67);
xor U5099 (N_5099,N_3122,N_840);
nor U5100 (N_5100,N_3655,N_36);
or U5101 (N_5101,N_3,N_659);
xor U5102 (N_5102,N_440,N_892);
nand U5103 (N_5103,N_1052,N_2232);
and U5104 (N_5104,N_2071,N_4743);
nand U5105 (N_5105,N_2449,N_513);
nand U5106 (N_5106,N_3703,N_4224);
nor U5107 (N_5107,N_4773,N_2338);
xor U5108 (N_5108,N_2683,N_3083);
or U5109 (N_5109,N_2251,N_4626);
or U5110 (N_5110,N_3059,N_546);
nand U5111 (N_5111,N_1799,N_698);
nor U5112 (N_5112,N_2699,N_3309);
or U5113 (N_5113,N_4675,N_4705);
or U5114 (N_5114,N_3425,N_4000);
nor U5115 (N_5115,N_3233,N_4324);
and U5116 (N_5116,N_992,N_2689);
or U5117 (N_5117,N_4978,N_102);
and U5118 (N_5118,N_4630,N_1904);
xor U5119 (N_5119,N_4778,N_2309);
nand U5120 (N_5120,N_1167,N_4297);
nor U5121 (N_5121,N_4824,N_536);
xor U5122 (N_5122,N_4672,N_726);
or U5123 (N_5123,N_3208,N_1906);
or U5124 (N_5124,N_3025,N_292);
xor U5125 (N_5125,N_1738,N_810);
and U5126 (N_5126,N_204,N_3776);
xnor U5127 (N_5127,N_207,N_4682);
nor U5128 (N_5128,N_1262,N_1423);
or U5129 (N_5129,N_3816,N_2057);
and U5130 (N_5130,N_385,N_3652);
nor U5131 (N_5131,N_547,N_3218);
nor U5132 (N_5132,N_749,N_1102);
and U5133 (N_5133,N_3300,N_1816);
xor U5134 (N_5134,N_3079,N_2370);
or U5135 (N_5135,N_1989,N_1280);
nor U5136 (N_5136,N_1695,N_2592);
and U5137 (N_5137,N_4751,N_252);
xnor U5138 (N_5138,N_578,N_1950);
or U5139 (N_5139,N_4657,N_1237);
or U5140 (N_5140,N_473,N_4046);
nor U5141 (N_5141,N_4515,N_224);
and U5142 (N_5142,N_1807,N_446);
xor U5143 (N_5143,N_3220,N_4595);
xor U5144 (N_5144,N_1686,N_3661);
nand U5145 (N_5145,N_3282,N_2564);
and U5146 (N_5146,N_277,N_2609);
or U5147 (N_5147,N_2954,N_4467);
nor U5148 (N_5148,N_3727,N_491);
nor U5149 (N_5149,N_4532,N_4947);
nor U5150 (N_5150,N_3850,N_4059);
nor U5151 (N_5151,N_4969,N_3667);
nand U5152 (N_5152,N_3246,N_2636);
and U5153 (N_5153,N_2860,N_293);
nand U5154 (N_5154,N_622,N_3629);
or U5155 (N_5155,N_3747,N_1353);
xnor U5156 (N_5156,N_2832,N_1350);
nor U5157 (N_5157,N_1170,N_4165);
or U5158 (N_5158,N_123,N_2085);
or U5159 (N_5159,N_894,N_2380);
and U5160 (N_5160,N_1495,N_48);
or U5161 (N_5161,N_2394,N_410);
nand U5162 (N_5162,N_2072,N_3782);
and U5163 (N_5163,N_1735,N_3221);
xnor U5164 (N_5164,N_960,N_4642);
nor U5165 (N_5165,N_1563,N_2688);
and U5166 (N_5166,N_4803,N_4358);
and U5167 (N_5167,N_4654,N_2635);
and U5168 (N_5168,N_172,N_4555);
and U5169 (N_5169,N_2303,N_2730);
or U5170 (N_5170,N_765,N_3299);
or U5171 (N_5171,N_4196,N_3409);
nand U5172 (N_5172,N_3176,N_4656);
xor U5173 (N_5173,N_3496,N_1463);
and U5174 (N_5174,N_4507,N_1971);
and U5175 (N_5175,N_3874,N_4756);
and U5176 (N_5176,N_798,N_2170);
or U5177 (N_5177,N_2256,N_4223);
and U5178 (N_5178,N_166,N_471);
or U5179 (N_5179,N_1937,N_4896);
nand U5180 (N_5180,N_1630,N_4770);
nand U5181 (N_5181,N_3965,N_2575);
or U5182 (N_5182,N_3696,N_2197);
xor U5183 (N_5183,N_4075,N_2193);
nand U5184 (N_5184,N_4105,N_3909);
or U5185 (N_5185,N_495,N_4364);
nor U5186 (N_5186,N_1720,N_898);
nand U5187 (N_5187,N_372,N_1367);
xor U5188 (N_5188,N_4340,N_3456);
or U5189 (N_5189,N_653,N_4971);
nor U5190 (N_5190,N_854,N_1450);
xnor U5191 (N_5191,N_3336,N_1004);
and U5192 (N_5192,N_1774,N_4146);
nand U5193 (N_5193,N_3830,N_1299);
xor U5194 (N_5194,N_919,N_3649);
xnor U5195 (N_5195,N_1227,N_1099);
and U5196 (N_5196,N_4333,N_3642);
and U5197 (N_5197,N_1360,N_3080);
or U5198 (N_5198,N_4564,N_3914);
nand U5199 (N_5199,N_3511,N_1055);
or U5200 (N_5200,N_4239,N_1177);
and U5201 (N_5201,N_190,N_296);
or U5202 (N_5202,N_65,N_4872);
and U5203 (N_5203,N_1127,N_752);
and U5204 (N_5204,N_2590,N_3366);
or U5205 (N_5205,N_2225,N_830);
nor U5206 (N_5206,N_1512,N_2668);
xnor U5207 (N_5207,N_4141,N_2922);
and U5208 (N_5208,N_217,N_2870);
nor U5209 (N_5209,N_1230,N_2101);
and U5210 (N_5210,N_4137,N_3582);
nor U5211 (N_5211,N_3418,N_3810);
or U5212 (N_5212,N_356,N_3007);
nand U5213 (N_5213,N_230,N_492);
nor U5214 (N_5214,N_2678,N_654);
or U5215 (N_5215,N_1141,N_4806);
or U5216 (N_5216,N_206,N_3869);
and U5217 (N_5217,N_3695,N_181);
xnor U5218 (N_5218,N_4558,N_3996);
nor U5219 (N_5219,N_2572,N_3811);
xnor U5220 (N_5220,N_861,N_2630);
and U5221 (N_5221,N_3866,N_1708);
and U5222 (N_5222,N_4548,N_3824);
nand U5223 (N_5223,N_989,N_99);
xor U5224 (N_5224,N_3786,N_4817);
and U5225 (N_5225,N_1685,N_629);
and U5226 (N_5226,N_1762,N_2541);
and U5227 (N_5227,N_866,N_3460);
nor U5228 (N_5228,N_1931,N_603);
or U5229 (N_5229,N_4600,N_917);
nor U5230 (N_5230,N_2589,N_3150);
or U5231 (N_5231,N_3651,N_4286);
or U5232 (N_5232,N_4664,N_2840);
or U5233 (N_5233,N_2153,N_996);
xor U5234 (N_5234,N_1244,N_2301);
xor U5235 (N_5235,N_592,N_3444);
or U5236 (N_5236,N_1222,N_2188);
xor U5237 (N_5237,N_2927,N_2440);
and U5238 (N_5238,N_1857,N_2219);
nand U5239 (N_5239,N_1594,N_3019);
and U5240 (N_5240,N_3733,N_1077);
nand U5241 (N_5241,N_4694,N_1608);
or U5242 (N_5242,N_2732,N_981);
and U5243 (N_5243,N_1546,N_4269);
nor U5244 (N_5244,N_4639,N_54);
nor U5245 (N_5245,N_1770,N_1254);
and U5246 (N_5246,N_3804,N_485);
nand U5247 (N_5247,N_883,N_210);
nand U5248 (N_5248,N_4924,N_4869);
or U5249 (N_5249,N_4771,N_2106);
or U5250 (N_5250,N_2496,N_2062);
nor U5251 (N_5251,N_1723,N_428);
or U5252 (N_5252,N_1732,N_3170);
or U5253 (N_5253,N_3448,N_1356);
xnor U5254 (N_5254,N_31,N_2407);
nand U5255 (N_5255,N_3888,N_2983);
nor U5256 (N_5256,N_2302,N_2151);
nor U5257 (N_5257,N_705,N_259);
or U5258 (N_5258,N_1080,N_4949);
or U5259 (N_5259,N_1648,N_4706);
nor U5260 (N_5260,N_167,N_2561);
or U5261 (N_5261,N_3174,N_4347);
and U5262 (N_5262,N_1572,N_3355);
nor U5263 (N_5263,N_1875,N_1521);
nor U5264 (N_5264,N_4876,N_4531);
nand U5265 (N_5265,N_581,N_3891);
and U5266 (N_5266,N_3993,N_3940);
or U5267 (N_5267,N_2160,N_2426);
and U5268 (N_5268,N_523,N_2139);
nand U5269 (N_5269,N_86,N_4111);
nor U5270 (N_5270,N_2836,N_786);
nor U5271 (N_5271,N_1106,N_3343);
and U5272 (N_5272,N_352,N_2772);
nand U5273 (N_5273,N_4368,N_2200);
nand U5274 (N_5274,N_667,N_1924);
xor U5275 (N_5275,N_4912,N_3034);
nor U5276 (N_5276,N_948,N_3084);
nand U5277 (N_5277,N_3104,N_1835);
or U5278 (N_5278,N_848,N_494);
xor U5279 (N_5279,N_2510,N_61);
and U5280 (N_5280,N_1408,N_1456);
nor U5281 (N_5281,N_597,N_3467);
and U5282 (N_5282,N_1053,N_784);
and U5283 (N_5283,N_4257,N_3364);
xor U5284 (N_5284,N_4990,N_2778);
xnor U5285 (N_5285,N_1564,N_1015);
nor U5286 (N_5286,N_3400,N_719);
or U5287 (N_5287,N_4540,N_4903);
xor U5288 (N_5288,N_1851,N_2526);
and U5289 (N_5289,N_4923,N_664);
and U5290 (N_5290,N_1246,N_567);
and U5291 (N_5291,N_3781,N_1331);
nor U5292 (N_5292,N_1128,N_1054);
nor U5293 (N_5293,N_4554,N_4758);
nor U5294 (N_5294,N_312,N_4900);
nand U5295 (N_5295,N_97,N_872);
nor U5296 (N_5296,N_1864,N_4098);
and U5297 (N_5297,N_2326,N_1515);
nand U5298 (N_5298,N_4841,N_3603);
or U5299 (N_5299,N_3507,N_3146);
or U5300 (N_5300,N_1997,N_1211);
or U5301 (N_5301,N_2324,N_1605);
xnor U5302 (N_5302,N_689,N_2137);
nand U5303 (N_5303,N_2692,N_3492);
nand U5304 (N_5304,N_4396,N_2909);
xnor U5305 (N_5305,N_3719,N_2788);
nor U5306 (N_5306,N_758,N_2595);
nor U5307 (N_5307,N_3276,N_4217);
or U5308 (N_5308,N_1878,N_739);
xnor U5309 (N_5309,N_4158,N_970);
or U5310 (N_5310,N_557,N_3580);
or U5311 (N_5311,N_301,N_1591);
xor U5312 (N_5312,N_2296,N_4491);
nand U5313 (N_5313,N_1613,N_4382);
nand U5314 (N_5314,N_965,N_3447);
nor U5315 (N_5315,N_3973,N_3430);
nor U5316 (N_5316,N_968,N_419);
xnor U5317 (N_5317,N_2304,N_1468);
nand U5318 (N_5318,N_2932,N_2079);
nand U5319 (N_5319,N_4320,N_4635);
xor U5320 (N_5320,N_3463,N_3089);
nand U5321 (N_5321,N_1926,N_1288);
xnor U5322 (N_5322,N_3037,N_2457);
and U5323 (N_5323,N_2138,N_4448);
or U5324 (N_5324,N_2529,N_168);
nand U5325 (N_5325,N_1913,N_1990);
xor U5326 (N_5326,N_3662,N_1702);
xor U5327 (N_5327,N_3268,N_3906);
nor U5328 (N_5328,N_2262,N_4240);
xor U5329 (N_5329,N_4742,N_1724);
nand U5330 (N_5330,N_4290,N_4219);
or U5331 (N_5331,N_1345,N_2454);
and U5332 (N_5332,N_3923,N_2291);
nor U5333 (N_5333,N_2930,N_3508);
nor U5334 (N_5334,N_1075,N_855);
xor U5335 (N_5335,N_4025,N_3382);
nand U5336 (N_5336,N_4922,N_158);
nor U5337 (N_5337,N_2968,N_2625);
xor U5338 (N_5338,N_3337,N_2820);
xor U5339 (N_5339,N_1149,N_3552);
nand U5340 (N_5340,N_666,N_768);
nand U5341 (N_5341,N_1575,N_3945);
nor U5342 (N_5342,N_1645,N_3414);
or U5343 (N_5343,N_2142,N_4195);
and U5344 (N_5344,N_778,N_4014);
or U5345 (N_5345,N_2581,N_1527);
xnor U5346 (N_5346,N_4373,N_800);
xnor U5347 (N_5347,N_4113,N_2728);
or U5348 (N_5348,N_3134,N_3204);
xnor U5349 (N_5349,N_3111,N_936);
nor U5350 (N_5350,N_1999,N_2260);
xor U5351 (N_5351,N_151,N_4139);
xor U5352 (N_5352,N_2221,N_1197);
or U5353 (N_5353,N_4090,N_269);
or U5354 (N_5354,N_527,N_381);
or U5355 (N_5355,N_3650,N_3175);
nor U5356 (N_5356,N_3793,N_4218);
nand U5357 (N_5357,N_4619,N_3980);
nand U5358 (N_5358,N_3673,N_4802);
xnor U5359 (N_5359,N_56,N_153);
and U5360 (N_5360,N_3709,N_3068);
nand U5361 (N_5361,N_1005,N_2337);
nand U5362 (N_5362,N_2721,N_1920);
and U5363 (N_5363,N_2654,N_3261);
or U5364 (N_5364,N_803,N_2484);
nand U5365 (N_5365,N_3647,N_451);
nand U5366 (N_5366,N_2317,N_366);
and U5367 (N_5367,N_3628,N_3639);
nand U5368 (N_5368,N_877,N_1947);
nor U5369 (N_5369,N_2560,N_4920);
or U5370 (N_5370,N_3551,N_2474);
or U5371 (N_5371,N_155,N_3234);
and U5372 (N_5372,N_3327,N_740);
nand U5373 (N_5373,N_1095,N_3312);
and U5374 (N_5374,N_1364,N_1315);
xor U5375 (N_5375,N_55,N_3149);
nand U5376 (N_5376,N_3885,N_3437);
and U5377 (N_5377,N_4492,N_3871);
and U5378 (N_5378,N_729,N_1832);
or U5379 (N_5379,N_870,N_3676);
nand U5380 (N_5380,N_3683,N_3592);
nor U5381 (N_5381,N_1418,N_2825);
nor U5382 (N_5382,N_276,N_1899);
xor U5383 (N_5383,N_2281,N_4713);
or U5384 (N_5384,N_2713,N_755);
xnor U5385 (N_5385,N_3503,N_655);
or U5386 (N_5386,N_4037,N_4039);
nand U5387 (N_5387,N_2274,N_891);
and U5388 (N_5388,N_2664,N_1533);
nor U5389 (N_5389,N_3573,N_906);
nand U5390 (N_5390,N_4670,N_1562);
and U5391 (N_5391,N_4084,N_4612);
nor U5392 (N_5392,N_1235,N_4583);
xnor U5393 (N_5393,N_516,N_1873);
or U5394 (N_5394,N_4399,N_1462);
nor U5395 (N_5395,N_1545,N_2864);
xnor U5396 (N_5396,N_1596,N_2390);
or U5397 (N_5397,N_4035,N_1451);
and U5398 (N_5398,N_3354,N_2867);
or U5399 (N_5399,N_4002,N_776);
xnor U5400 (N_5400,N_498,N_1101);
or U5401 (N_5401,N_2438,N_1287);
or U5402 (N_5402,N_2258,N_2435);
xor U5403 (N_5403,N_2391,N_3849);
nor U5404 (N_5404,N_3127,N_2731);
and U5405 (N_5405,N_4268,N_2400);
xor U5406 (N_5406,N_1365,N_2765);
xor U5407 (N_5407,N_3918,N_1829);
xor U5408 (N_5408,N_2330,N_3700);
and U5409 (N_5409,N_50,N_4161);
nand U5410 (N_5410,N_4194,N_3725);
nand U5411 (N_5411,N_3887,N_3254);
xor U5412 (N_5412,N_1973,N_4052);
and U5413 (N_5413,N_687,N_2147);
and U5414 (N_5414,N_2854,N_4814);
xor U5415 (N_5415,N_422,N_949);
nor U5416 (N_5416,N_1517,N_3033);
or U5417 (N_5417,N_1354,N_3273);
and U5418 (N_5418,N_839,N_1039);
or U5419 (N_5419,N_4804,N_4424);
nand U5420 (N_5420,N_3867,N_2796);
or U5421 (N_5421,N_4261,N_264);
nor U5422 (N_5422,N_4580,N_1601);
nand U5423 (N_5423,N_1862,N_1425);
nor U5424 (N_5424,N_2451,N_2026);
and U5425 (N_5425,N_1681,N_4611);
and U5426 (N_5426,N_3385,N_1486);
xor U5427 (N_5427,N_1187,N_4825);
xnor U5428 (N_5428,N_569,N_1290);
and U5429 (N_5429,N_437,N_1771);
xor U5430 (N_5430,N_4663,N_4338);
or U5431 (N_5431,N_1260,N_4589);
nor U5432 (N_5432,N_1998,N_1045);
and U5433 (N_5433,N_4556,N_1506);
nor U5434 (N_5434,N_1697,N_131);
and U5435 (N_5435,N_3749,N_572);
xnor U5436 (N_5436,N_1012,N_4721);
xnor U5437 (N_5437,N_2198,N_663);
nor U5438 (N_5438,N_117,N_2049);
nor U5439 (N_5439,N_430,N_4360);
and U5440 (N_5440,N_3199,N_805);
nand U5441 (N_5441,N_1014,N_3589);
nand U5442 (N_5442,N_3097,N_4099);
xor U5443 (N_5443,N_4594,N_1633);
xnor U5444 (N_5444,N_1954,N_2918);
xnor U5445 (N_5445,N_4536,N_1718);
and U5446 (N_5446,N_3278,N_2881);
or U5447 (N_5447,N_761,N_1877);
nand U5448 (N_5448,N_780,N_3197);
xnor U5449 (N_5449,N_3870,N_4636);
and U5450 (N_5450,N_1112,N_4388);
xnor U5451 (N_5451,N_4957,N_3402);
nand U5452 (N_5452,N_4420,N_637);
and U5453 (N_5453,N_1181,N_2598);
xor U5454 (N_5454,N_1660,N_4357);
nor U5455 (N_5455,N_275,N_790);
and U5456 (N_5456,N_2551,N_3478);
and U5457 (N_5457,N_2633,N_1409);
nand U5458 (N_5458,N_3946,N_624);
xnor U5459 (N_5459,N_2434,N_4355);
xnor U5460 (N_5460,N_1802,N_2404);
xnor U5461 (N_5461,N_3360,N_3132);
nand U5462 (N_5462,N_2339,N_2539);
and U5463 (N_5463,N_4941,N_3223);
xor U5464 (N_5464,N_1719,N_4641);
xor U5465 (N_5465,N_4874,N_1474);
xnor U5466 (N_5466,N_4170,N_1493);
and U5467 (N_5467,N_2773,N_4658);
and U5468 (N_5468,N_1759,N_3229);
and U5469 (N_5469,N_4901,N_3543);
nor U5470 (N_5470,N_4234,N_4319);
nor U5471 (N_5471,N_2476,N_4392);
and U5472 (N_5472,N_195,N_2332);
nor U5473 (N_5473,N_2787,N_844);
and U5474 (N_5474,N_313,N_1598);
and U5475 (N_5475,N_3267,N_345);
and U5476 (N_5476,N_4216,N_3260);
xor U5477 (N_5477,N_3735,N_1714);
or U5478 (N_5478,N_246,N_4461);
nor U5479 (N_5479,N_1094,N_3608);
or U5480 (N_5480,N_3010,N_4982);
and U5481 (N_5481,N_1806,N_1789);
or U5482 (N_5482,N_3003,N_1002);
nand U5483 (N_5483,N_4807,N_3350);
or U5484 (N_5484,N_2523,N_1709);
or U5485 (N_5485,N_4272,N_3305);
nand U5486 (N_5486,N_2127,N_2662);
nor U5487 (N_5487,N_718,N_2898);
nand U5488 (N_5488,N_4991,N_4354);
nor U5489 (N_5489,N_1849,N_2616);
and U5490 (N_5490,N_3520,N_2691);
or U5491 (N_5491,N_1717,N_3399);
nor U5492 (N_5492,N_2421,N_3817);
nand U5493 (N_5493,N_1443,N_4754);
nand U5494 (N_5494,N_2213,N_1979);
and U5495 (N_5495,N_907,N_2629);
nor U5496 (N_5496,N_111,N_2342);
nor U5497 (N_5497,N_474,N_2450);
xnor U5498 (N_5498,N_423,N_4575);
nand U5499 (N_5499,N_2952,N_2674);
xnor U5500 (N_5500,N_3623,N_721);
nand U5501 (N_5501,N_2487,N_1516);
nand U5502 (N_5502,N_4829,N_2527);
or U5503 (N_5503,N_2935,N_1320);
nor U5504 (N_5504,N_3527,N_1908);
nor U5505 (N_5505,N_1531,N_2719);
or U5506 (N_5506,N_1234,N_466);
and U5507 (N_5507,N_2249,N_1957);
or U5508 (N_5508,N_100,N_2549);
nor U5509 (N_5509,N_760,N_771);
xnor U5510 (N_5510,N_3862,N_4516);
nor U5511 (N_5511,N_2288,N_3242);
nand U5512 (N_5512,N_1540,N_2458);
nand U5513 (N_5513,N_1823,N_2174);
nor U5514 (N_5514,N_2970,N_2739);
nor U5515 (N_5515,N_41,N_2039);
xor U5516 (N_5516,N_4383,N_3274);
nand U5517 (N_5517,N_2849,N_993);
xnor U5518 (N_5518,N_3841,N_2333);
nand U5519 (N_5519,N_3051,N_1751);
xnor U5520 (N_5520,N_676,N_4466);
nand U5521 (N_5521,N_3979,N_4119);
nand U5522 (N_5522,N_3748,N_4389);
xnor U5523 (N_5523,N_2708,N_1284);
nor U5524 (N_5524,N_684,N_2532);
and U5525 (N_5525,N_2122,N_414);
xor U5526 (N_5526,N_1482,N_617);
and U5527 (N_5527,N_3765,N_1741);
nor U5528 (N_5528,N_2749,N_27);
or U5529 (N_5529,N_4082,N_2618);
xnor U5530 (N_5530,N_2131,N_3406);
nor U5531 (N_5531,N_7,N_78);
xnor U5532 (N_5532,N_3986,N_1803);
or U5533 (N_5533,N_4775,N_409);
xor U5534 (N_5534,N_2929,N_1532);
nor U5535 (N_5535,N_1834,N_26);
nor U5536 (N_5536,N_1687,N_2516);
or U5537 (N_5537,N_2100,N_3898);
xor U5538 (N_5538,N_808,N_1377);
xnor U5539 (N_5539,N_3332,N_1658);
or U5540 (N_5540,N_1393,N_327);
and U5541 (N_5541,N_2042,N_1064);
or U5542 (N_5542,N_4852,N_4809);
or U5543 (N_5543,N_2382,N_501);
nand U5544 (N_5544,N_1339,N_1529);
and U5545 (N_5545,N_1501,N_2627);
and U5546 (N_5546,N_3412,N_1194);
nor U5547 (N_5547,N_545,N_2953);
nand U5548 (N_5548,N_1189,N_3243);
and U5549 (N_5549,N_4501,N_929);
and U5550 (N_5550,N_685,N_193);
nor U5551 (N_5551,N_1604,N_1573);
and U5552 (N_5552,N_1413,N_4601);
xnor U5553 (N_5553,N_4585,N_4221);
xnor U5554 (N_5554,N_4436,N_2102);
nor U5555 (N_5555,N_208,N_3394);
nand U5556 (N_5556,N_3566,N_2017);
and U5557 (N_5557,N_3882,N_1151);
xor U5558 (N_5558,N_915,N_4255);
nor U5559 (N_5559,N_1577,N_459);
and U5560 (N_5560,N_1297,N_1949);
and U5561 (N_5561,N_606,N_710);
xor U5562 (N_5562,N_1765,N_3110);
and U5563 (N_5563,N_2665,N_3855);
nand U5564 (N_5564,N_2557,N_1172);
and U5565 (N_5565,N_4645,N_3124);
and U5566 (N_5566,N_4761,N_265);
and U5567 (N_5567,N_2253,N_2128);
xnor U5568 (N_5568,N_1553,N_2346);
or U5569 (N_5569,N_1225,N_4652);
nor U5570 (N_5570,N_1378,N_2465);
nand U5571 (N_5571,N_925,N_3494);
nand U5572 (N_5572,N_4162,N_4909);
and U5573 (N_5573,N_4076,N_3147);
nor U5574 (N_5574,N_4692,N_2868);
or U5575 (N_5575,N_4386,N_113);
nor U5576 (N_5576,N_2847,N_3339);
nor U5577 (N_5577,N_3578,N_835);
or U5578 (N_5578,N_4958,N_4779);
nand U5579 (N_5579,N_3549,N_3069);
nor U5580 (N_5580,N_3143,N_3005);
nor U5581 (N_5581,N_1651,N_2495);
and U5582 (N_5582,N_2046,N_1389);
nor U5583 (N_5583,N_240,N_1471);
and U5584 (N_5584,N_4603,N_1164);
nand U5585 (N_5585,N_4381,N_3042);
or U5586 (N_5586,N_1081,N_4884);
and U5587 (N_5587,N_754,N_98);
nor U5588 (N_5588,N_2038,N_4088);
nor U5589 (N_5589,N_3879,N_1996);
nand U5590 (N_5590,N_3801,N_3772);
nand U5591 (N_5591,N_1349,N_2007);
nand U5592 (N_5592,N_2685,N_1333);
and U5593 (N_5593,N_702,N_3029);
or U5594 (N_5594,N_340,N_2372);
and U5595 (N_5595,N_1397,N_3734);
xor U5596 (N_5596,N_1557,N_591);
xor U5597 (N_5597,N_681,N_1637);
and U5598 (N_5598,N_956,N_1798);
or U5599 (N_5599,N_2544,N_47);
nand U5600 (N_5600,N_3371,N_4304);
nor U5601 (N_5601,N_817,N_3311);
nand U5602 (N_5602,N_1440,N_2734);
nor U5603 (N_5603,N_2742,N_4412);
and U5604 (N_5604,N_4812,N_1750);
or U5605 (N_5605,N_650,N_3230);
xor U5606 (N_5606,N_2877,N_462);
or U5607 (N_5607,N_2224,N_3829);
nand U5608 (N_5608,N_1357,N_469);
xor U5609 (N_5609,N_3773,N_1483);
or U5610 (N_5610,N_4932,N_2917);
or U5611 (N_5611,N_429,N_920);
or U5612 (N_5612,N_2669,N_3427);
nand U5613 (N_5613,N_438,N_616);
nand U5614 (N_5614,N_3480,N_2082);
nor U5615 (N_5615,N_3459,N_4660);
nor U5616 (N_5616,N_354,N_3182);
nand U5617 (N_5617,N_1544,N_4292);
and U5618 (N_5618,N_2293,N_2876);
and U5619 (N_5619,N_1071,N_3404);
xnor U5620 (N_5620,N_69,N_2886);
or U5621 (N_5621,N_3762,N_1915);
nor U5622 (N_5622,N_1923,N_1944);
nand U5623 (N_5623,N_4140,N_635);
xnor U5624 (N_5624,N_2941,N_2273);
nand U5625 (N_5625,N_3102,N_3441);
xor U5626 (N_5626,N_4351,N_3484);
or U5627 (N_5627,N_4587,N_371);
nor U5628 (N_5628,N_2902,N_922);
and U5629 (N_5629,N_636,N_1928);
nand U5630 (N_5630,N_2661,N_1917);
nor U5631 (N_5631,N_2851,N_302);
and U5632 (N_5632,N_3476,N_4430);
xor U5633 (N_5633,N_4313,N_2381);
nand U5634 (N_5634,N_3711,N_846);
or U5635 (N_5635,N_2124,N_3001);
nor U5636 (N_5636,N_4478,N_2582);
xor U5637 (N_5637,N_4650,N_1410);
xnor U5638 (N_5638,N_804,N_3333);
nor U5639 (N_5639,N_3959,N_1850);
nand U5640 (N_5640,N_3014,N_4961);
xnor U5641 (N_5641,N_2770,N_4155);
and U5642 (N_5642,N_3777,N_1332);
and U5643 (N_5643,N_79,N_17);
xor U5644 (N_5644,N_2566,N_2933);
xor U5645 (N_5645,N_2183,N_598);
and U5646 (N_5646,N_632,N_3942);
and U5647 (N_5647,N_4838,N_887);
and U5648 (N_5648,N_468,N_1229);
or U5649 (N_5649,N_2360,N_4344);
nand U5650 (N_5650,N_329,N_1416);
xor U5651 (N_5651,N_4243,N_1372);
and U5652 (N_5652,N_4928,N_213);
and U5653 (N_5653,N_4518,N_2624);
nand U5654 (N_5654,N_1549,N_4118);
nand U5655 (N_5655,N_930,N_1017);
xor U5656 (N_5656,N_221,N_2204);
nor U5657 (N_5657,N_3919,N_164);
xor U5658 (N_5658,N_1322,N_4463);
nor U5659 (N_5659,N_2405,N_4863);
nor U5660 (N_5660,N_500,N_2034);
and U5661 (N_5661,N_4683,N_1650);
nand U5662 (N_5662,N_2520,N_1264);
and U5663 (N_5663,N_748,N_699);
and U5664 (N_5664,N_2278,N_3255);
nor U5665 (N_5665,N_3633,N_87);
xor U5666 (N_5666,N_522,N_4985);
or U5667 (N_5667,N_3004,N_3833);
nor U5668 (N_5668,N_3831,N_262);
nor U5669 (N_5669,N_503,N_2716);
nor U5670 (N_5670,N_1051,N_2528);
nand U5671 (N_5671,N_2111,N_571);
and U5672 (N_5672,N_3353,N_1047);
and U5673 (N_5673,N_73,N_245);
or U5674 (N_5674,N_2658,N_2735);
and U5675 (N_5675,N_2759,N_2120);
and U5676 (N_5676,N_3035,N_3522);
and U5677 (N_5677,N_4001,N_412);
or U5678 (N_5678,N_3250,N_3165);
xnor U5679 (N_5679,N_3512,N_4310);
and U5680 (N_5680,N_2356,N_1184);
or U5681 (N_5681,N_3922,N_4850);
and U5682 (N_5682,N_3320,N_972);
nand U5683 (N_5683,N_4615,N_1392);
and U5684 (N_5684,N_1146,N_4588);
xor U5685 (N_5685,N_1180,N_1036);
and U5686 (N_5686,N_255,N_3500);
and U5687 (N_5687,N_1302,N_4254);
or U5688 (N_5688,N_3107,N_985);
nor U5689 (N_5689,N_2764,N_1542);
and U5690 (N_5690,N_2126,N_4418);
xor U5691 (N_5691,N_4541,N_2714);
nand U5692 (N_5692,N_408,N_162);
or U5693 (N_5693,N_4981,N_900);
nand U5694 (N_5694,N_2084,N_4551);
nand U5695 (N_5695,N_4519,N_3171);
nor U5696 (N_5696,N_3114,N_530);
nand U5697 (N_5697,N_2344,N_1479);
or U5698 (N_5698,N_3044,N_4294);
or U5699 (N_5699,N_1025,N_3067);
nor U5700 (N_5700,N_1243,N_3421);
or U5701 (N_5701,N_2977,N_3713);
nor U5702 (N_5702,N_1395,N_4970);
nor U5703 (N_5703,N_982,N_1856);
xnor U5704 (N_5704,N_2989,N_1270);
or U5705 (N_5705,N_96,N_812);
or U5706 (N_5706,N_3446,N_2822);
or U5707 (N_5707,N_3886,N_4505);
xnor U5708 (N_5708,N_2519,N_1006);
or U5709 (N_5709,N_373,N_2105);
nor U5710 (N_5710,N_2226,N_4425);
nor U5711 (N_5711,N_3895,N_4328);
or U5712 (N_5712,N_1508,N_2154);
nand U5713 (N_5713,N_109,N_4891);
nor U5714 (N_5714,N_713,N_3779);
nand U5715 (N_5715,N_361,N_4848);
nor U5716 (N_5716,N_1706,N_3636);
xnor U5717 (N_5717,N_4943,N_1066);
nand U5718 (N_5718,N_4504,N_2823);
or U5719 (N_5719,N_875,N_2110);
or U5720 (N_5720,N_1476,N_2202);
nand U5721 (N_5721,N_3062,N_2858);
xor U5722 (N_5722,N_4729,N_3172);
and U5723 (N_5723,N_1422,N_1940);
nor U5724 (N_5724,N_2944,N_2907);
nand U5725 (N_5725,N_3805,N_2672);
xor U5726 (N_5726,N_3075,N_651);
and U5727 (N_5727,N_4902,N_4006);
nor U5728 (N_5728,N_39,N_1641);
or U5729 (N_5729,N_3984,N_2533);
xnor U5730 (N_5730,N_2092,N_2215);
xor U5731 (N_5731,N_370,N_1525);
nand U5732 (N_5732,N_149,N_1359);
or U5733 (N_5733,N_2508,N_15);
nor U5734 (N_5734,N_1489,N_397);
and U5735 (N_5735,N_2752,N_997);
nor U5736 (N_5736,N_3087,N_3595);
xnor U5737 (N_5737,N_1374,N_4590);
nand U5738 (N_5738,N_3335,N_3534);
xnor U5739 (N_5739,N_3764,N_3205);
xor U5740 (N_5740,N_3189,N_3939);
nand U5741 (N_5741,N_4974,N_3469);
xnor U5742 (N_5742,N_1838,N_4441);
and U5743 (N_5743,N_1276,N_2956);
nand U5744 (N_5744,N_2563,N_3471);
or U5745 (N_5745,N_2211,N_4107);
nand U5746 (N_5746,N_4205,N_1846);
nand U5747 (N_5747,N_415,N_2852);
nand U5748 (N_5748,N_911,N_3860);
nor U5749 (N_5749,N_374,N_3585);
nor U5750 (N_5750,N_3893,N_402);
and U5751 (N_5751,N_1289,N_2891);
or U5752 (N_5752,N_2920,N_2769);
nand U5753 (N_5753,N_794,N_4860);
and U5754 (N_5754,N_2490,N_1379);
nor U5755 (N_5755,N_3851,N_2307);
or U5756 (N_5756,N_2597,N_152);
nor U5757 (N_5757,N_1618,N_1381);
nor U5758 (N_5758,N_4833,N_1593);
nor U5759 (N_5759,N_4939,N_3514);
nand U5760 (N_5760,N_1200,N_3153);
and U5761 (N_5761,N_2118,N_1199);
and U5762 (N_5762,N_1860,N_4450);
or U5763 (N_5763,N_83,N_1205);
xor U5764 (N_5764,N_619,N_4433);
nor U5765 (N_5765,N_3600,N_3266);
and U5766 (N_5766,N_3784,N_2460);
nand U5767 (N_5767,N_1404,N_3292);
xnor U5768 (N_5768,N_3865,N_2345);
and U5769 (N_5769,N_3297,N_4581);
and U5770 (N_5770,N_2890,N_3799);
nor U5771 (N_5771,N_2974,N_3653);
and U5772 (N_5772,N_261,N_933);
nor U5773 (N_5773,N_641,N_1805);
nor U5774 (N_5774,N_3240,N_816);
nor U5775 (N_5775,N_3501,N_4168);
nor U5776 (N_5776,N_1925,N_2943);
and U5777 (N_5777,N_3118,N_4733);
and U5778 (N_5778,N_4053,N_362);
or U5779 (N_5779,N_1932,N_669);
nand U5780 (N_5780,N_4314,N_2963);
nand U5781 (N_5781,N_2856,N_4514);
nand U5782 (N_5782,N_1797,N_336);
and U5783 (N_5783,N_3291,N_1008);
and U5784 (N_5784,N_4295,N_2141);
nor U5785 (N_5785,N_2171,N_1361);
xnor U5786 (N_5786,N_2504,N_3470);
nor U5787 (N_5787,N_2577,N_4525);
or U5788 (N_5788,N_1294,N_1342);
or U5789 (N_5789,N_1370,N_4925);
nand U5790 (N_5790,N_986,N_4130);
and U5791 (N_5791,N_4962,N_2140);
nand U5792 (N_5792,N_4598,N_3050);
and U5793 (N_5793,N_3722,N_3560);
nor U5794 (N_5794,N_376,N_728);
nor U5795 (N_5795,N_1087,N_657);
nand U5796 (N_5796,N_33,N_2348);
and U5797 (N_5797,N_81,N_4413);
nor U5798 (N_5798,N_4398,N_3561);
or U5799 (N_5799,N_4150,N_4708);
xnor U5800 (N_5800,N_978,N_2722);
nor U5801 (N_5801,N_3296,N_4124);
nand U5802 (N_5802,N_1121,N_1338);
and U5803 (N_5803,N_2853,N_1218);
xnor U5804 (N_5804,N_3568,N_4251);
xnor U5805 (N_5805,N_4267,N_53);
and U5806 (N_5806,N_3948,N_1292);
nand U5807 (N_5807,N_2328,N_2588);
xnor U5808 (N_5808,N_2816,N_2888);
nor U5809 (N_5809,N_4322,N_2845);
nor U5810 (N_5810,N_4780,N_3021);
nand U5811 (N_5811,N_4414,N_3617);
nand U5812 (N_5812,N_169,N_2041);
nor U5813 (N_5813,N_2824,N_4741);
and U5814 (N_5814,N_2239,N_2559);
and U5815 (N_5815,N_4610,N_4889);
and U5816 (N_5816,N_4691,N_1343);
nand U5817 (N_5817,N_19,N_3065);
and U5818 (N_5818,N_1824,N_4979);
nand U5819 (N_5819,N_4160,N_3902);
xnor U5820 (N_5820,N_4191,N_3515);
xnor U5821 (N_5821,N_229,N_1722);
nand U5822 (N_5822,N_526,N_2762);
xnor U5823 (N_5823,N_2511,N_733);
and U5824 (N_5824,N_2456,N_1614);
or U5825 (N_5825,N_1556,N_1424);
nor U5826 (N_5826,N_234,N_4417);
nor U5827 (N_5827,N_792,N_1125);
xor U5828 (N_5828,N_4264,N_1804);
nand U5829 (N_5829,N_1202,N_4096);
and U5830 (N_5830,N_3952,N_1683);
and U5831 (N_5831,N_2843,N_3288);
or U5832 (N_5832,N_2591,N_3795);
nand U5833 (N_5833,N_1285,N_4950);
xor U5834 (N_5834,N_2622,N_3052);
xnor U5835 (N_5835,N_399,N_3381);
or U5836 (N_5836,N_4402,N_2936);
nor U5837 (N_5837,N_744,N_1666);
xnor U5838 (N_5838,N_2741,N_706);
nor U5839 (N_5839,N_1324,N_9);
xor U5840 (N_5840,N_1282,N_2012);
xor U5841 (N_5841,N_2376,N_2396);
or U5842 (N_5842,N_1245,N_2536);
and U5843 (N_5843,N_2164,N_3499);
nor U5844 (N_5844,N_1927,N_2703);
xnor U5845 (N_5845,N_3248,N_1238);
and U5846 (N_5846,N_4929,N_1499);
nor U5847 (N_5847,N_741,N_3540);
xor U5848 (N_5848,N_2934,N_2310);
nor U5849 (N_5849,N_1625,N_3279);
nor U5850 (N_5850,N_772,N_3167);
nand U5851 (N_5851,N_4882,N_630);
nand U5852 (N_5852,N_3954,N_456);
and U5853 (N_5853,N_813,N_3349);
and U5854 (N_5854,N_1301,N_2074);
nand U5855 (N_5855,N_3438,N_4993);
xnor U5856 (N_5856,N_2637,N_1621);
nor U5857 (N_5857,N_889,N_1939);
nand U5858 (N_5858,N_2244,N_3550);
nand U5859 (N_5859,N_2420,N_3058);
nor U5860 (N_5860,N_4693,N_3258);
nand U5861 (N_5861,N_3557,N_2308);
and U5862 (N_5862,N_4475,N_1236);
nand U5863 (N_5863,N_2497,N_3968);
nand U5864 (N_5864,N_1673,N_3637);
nand U5865 (N_5865,N_4495,N_1656);
and U5866 (N_5866,N_1179,N_4799);
nor U5867 (N_5867,N_58,N_2694);
xor U5868 (N_5868,N_4868,N_389);
and U5869 (N_5869,N_2647,N_3040);
nand U5870 (N_5870,N_4716,N_4041);
and U5871 (N_5871,N_442,N_661);
nor U5872 (N_5872,N_355,N_1487);
nand U5873 (N_5873,N_4423,N_3796);
or U5874 (N_5874,N_3313,N_3685);
nor U5875 (N_5875,N_4291,N_1458);
nor U5876 (N_5876,N_1140,N_232);
and U5877 (N_5877,N_3181,N_4936);
nor U5878 (N_5878,N_398,N_2412);
xor U5879 (N_5879,N_1689,N_3495);
and U5880 (N_5880,N_2430,N_2485);
or U5881 (N_5881,N_1304,N_2994);
or U5882 (N_5882,N_37,N_3588);
or U5883 (N_5883,N_1152,N_1520);
xor U5884 (N_5884,N_401,N_3990);
xnor U5885 (N_5885,N_3417,N_833);
nor U5886 (N_5886,N_1820,N_3479);
xnor U5887 (N_5887,N_2800,N_132);
xnor U5888 (N_5888,N_4043,N_4886);
or U5889 (N_5889,N_4960,N_1664);
nor U5890 (N_5890,N_32,N_3113);
or U5891 (N_5891,N_1773,N_1380);
nor U5892 (N_5892,N_1163,N_2194);
xor U5893 (N_5893,N_4033,N_1662);
nand U5894 (N_5894,N_3370,N_2104);
xnor U5895 (N_5895,N_4623,N_1642);
xnor U5896 (N_5896,N_127,N_2362);
nand U5897 (N_5897,N_1929,N_946);
nor U5898 (N_5898,N_1067,N_2083);
or U5899 (N_5899,N_2676,N_1185);
nor U5900 (N_5900,N_4772,N_4235);
nor U5901 (N_5901,N_3961,N_4487);
nor U5902 (N_5902,N_233,N_2892);
xnor U5903 (N_5903,N_2088,N_251);
or U5904 (N_5904,N_2385,N_4508);
nor U5905 (N_5905,N_2991,N_4988);
or U5906 (N_5906,N_187,N_1730);
nand U5907 (N_5907,N_351,N_235);
xnor U5908 (N_5908,N_3988,N_3028);
and U5909 (N_5909,N_3324,N_218);
and U5910 (N_5910,N_2790,N_182);
nor U5911 (N_5911,N_2411,N_1881);
and U5912 (N_5912,N_2052,N_1118);
and U5913 (N_5913,N_3880,N_2626);
nor U5914 (N_5914,N_939,N_3048);
xor U5915 (N_5915,N_1273,N_853);
nor U5916 (N_5916,N_272,N_4677);
nand U5917 (N_5917,N_1703,N_3173);
and U5918 (N_5918,N_2166,N_4667);
or U5919 (N_5919,N_3378,N_4282);
and U5920 (N_5920,N_614,N_1272);
or U5921 (N_5921,N_4306,N_763);
nor U5922 (N_5922,N_4085,N_1587);
nand U5923 (N_5923,N_4061,N_3978);
xnor U5924 (N_5924,N_2512,N_4034);
nand U5925 (N_5925,N_3538,N_1784);
xor U5926 (N_5926,N_4776,N_3023);
xor U5927 (N_5927,N_2841,N_834);
xnor U5928 (N_5928,N_3541,N_4369);
and U5929 (N_5929,N_796,N_2747);
nand U5930 (N_5930,N_400,N_20);
and U5931 (N_5931,N_3006,N_4933);
xor U5932 (N_5932,N_2522,N_455);
xnor U5933 (N_5933,N_3590,N_342);
and U5934 (N_5934,N_3346,N_4605);
or U5935 (N_5935,N_1700,N_4572);
xnor U5936 (N_5936,N_3610,N_1042);
xor U5937 (N_5937,N_4676,N_4734);
nand U5938 (N_5938,N_4493,N_80);
xnor U5939 (N_5939,N_328,N_3101);
xor U5940 (N_5940,N_4371,N_4192);
xnor U5941 (N_5941,N_686,N_4078);
or U5942 (N_5942,N_3848,N_1281);
and U5943 (N_5943,N_241,N_3645);
nor U5944 (N_5944,N_3135,N_2611);
nand U5945 (N_5945,N_4821,N_633);
xor U5946 (N_5946,N_3191,N_2784);
or U5947 (N_5947,N_2107,N_4115);
nand U5948 (N_5948,N_3991,N_4167);
nand U5949 (N_5949,N_2265,N_2028);
nand U5950 (N_5950,N_365,N_743);
and U5951 (N_5951,N_4147,N_1033);
and U5952 (N_5952,N_1347,N_2724);
or U5953 (N_5953,N_3330,N_4524);
xor U5954 (N_5954,N_2813,N_4647);
xnor U5955 (N_5955,N_4506,N_3056);
nor U5956 (N_5956,N_4789,N_1415);
or U5957 (N_5957,N_1584,N_1098);
and U5958 (N_5958,N_3835,N_4503);
nand U5959 (N_5959,N_3428,N_4753);
and U5960 (N_5960,N_3213,N_4345);
or U5961 (N_5961,N_1215,N_1813);
nor U5962 (N_5962,N_1744,N_4293);
or U5963 (N_5963,N_3542,N_1900);
or U5964 (N_5964,N_1040,N_524);
nand U5965 (N_5965,N_4377,N_1430);
and U5966 (N_5966,N_1159,N_3970);
and U5967 (N_5967,N_1777,N_1733);
nand U5968 (N_5968,N_3938,N_3675);
nor U5969 (N_5969,N_3046,N_3136);
nand U5970 (N_5970,N_4937,N_3935);
nor U5971 (N_5971,N_3802,N_1113);
xor U5972 (N_5972,N_2831,N_3927);
nor U5973 (N_5973,N_1295,N_3525);
xnor U5974 (N_5974,N_532,N_122);
or U5975 (N_5975,N_1293,N_3187);
or U5976 (N_5976,N_4409,N_827);
or U5977 (N_5977,N_3690,N_2966);
or U5978 (N_5978,N_3775,N_645);
or U5979 (N_5979,N_1311,N_1880);
xor U5980 (N_5980,N_3625,N_3798);
xor U5981 (N_5981,N_4318,N_220);
nor U5982 (N_5982,N_3341,N_599);
nor U5983 (N_5983,N_1020,N_1554);
or U5984 (N_5984,N_1710,N_1126);
xor U5985 (N_5985,N_963,N_2494);
nor U5986 (N_5986,N_3680,N_3256);
nor U5987 (N_5987,N_4229,N_3432);
and U5988 (N_5988,N_3081,N_3086);
and U5989 (N_5989,N_2874,N_1212);
and U5990 (N_5990,N_1548,N_1800);
or U5991 (N_5991,N_943,N_4621);
nand U5992 (N_5992,N_4917,N_3556);
xor U5993 (N_5993,N_2899,N_1962);
nand U5994 (N_5994,N_1884,N_3787);
nor U5995 (N_5995,N_3844,N_4363);
xor U5996 (N_5996,N_2879,N_2601);
and U5997 (N_5997,N_1442,N_2859);
and U5998 (N_5998,N_3930,N_3679);
xor U5999 (N_5999,N_4760,N_1952);
or U6000 (N_6000,N_1830,N_1076);
or U6001 (N_6001,N_3196,N_1110);
xor U6002 (N_6002,N_4245,N_319);
nand U6003 (N_6003,N_1790,N_1902);
nand U6004 (N_6004,N_1490,N_4375);
nor U6005 (N_6005,N_4438,N_2146);
xnor U6006 (N_6006,N_4893,N_2815);
nand U6007 (N_6007,N_1518,N_1019);
or U6008 (N_6008,N_291,N_2108);
and U6009 (N_6009,N_2210,N_1465);
nand U6010 (N_6010,N_4465,N_1810);
xor U6011 (N_6011,N_4440,N_1032);
or U6012 (N_6012,N_639,N_3396);
nor U6013 (N_6013,N_518,N_4056);
nand U6014 (N_6014,N_4091,N_110);
nand U6015 (N_6015,N_3226,N_4737);
or U6016 (N_6016,N_2792,N_4468);
nor U6017 (N_6017,N_703,N_615);
xnor U6018 (N_6018,N_1585,N_3195);
nand U6019 (N_6019,N_8,N_403);
nand U6020 (N_6020,N_2065,N_3721);
nor U6021 (N_6021,N_1444,N_1837);
nor U6022 (N_6022,N_3401,N_3708);
and U6023 (N_6023,N_1844,N_3345);
nor U6024 (N_6024,N_84,N_4108);
and U6025 (N_6025,N_4995,N_314);
nand U6026 (N_6026,N_139,N_2906);
xor U6027 (N_6027,N_1224,N_3236);
xor U6028 (N_6028,N_4831,N_1943);
or U6029 (N_6029,N_538,N_16);
and U6030 (N_6030,N_2144,N_4624);
nor U6031 (N_6031,N_2059,N_3450);
nor U6032 (N_6032,N_2191,N_2250);
and U6033 (N_6033,N_324,N_2727);
or U6034 (N_6034,N_3521,N_4528);
nor U6035 (N_6035,N_2576,N_797);
nand U6036 (N_6036,N_1657,N_1056);
nor U6037 (N_6037,N_2873,N_4560);
nor U6038 (N_6038,N_1481,N_3474);
or U6039 (N_6039,N_3461,N_3145);
nor U6040 (N_6040,N_1994,N_4728);
nand U6041 (N_6041,N_2314,N_2254);
nand U6042 (N_6042,N_334,N_1420);
nor U6043 (N_6043,N_2521,N_2623);
and U6044 (N_6044,N_2921,N_209);
or U6045 (N_6045,N_2500,N_1966);
nor U6046 (N_6046,N_3548,N_1814);
xnor U6047 (N_6047,N_4362,N_4653);
xnor U6048 (N_6048,N_3604,N_4740);
or U6049 (N_6049,N_1606,N_4791);
nor U6050 (N_6050,N_3640,N_4058);
or U6051 (N_6051,N_2185,N_3270);
nor U6052 (N_6052,N_1208,N_528);
nand U6053 (N_6053,N_3315,N_1319);
or U6054 (N_6054,N_2025,N_49);
xor U6055 (N_6055,N_1511,N_3705);
xor U6056 (N_6056,N_3563,N_814);
nand U6057 (N_6057,N_4616,N_966);
nand U6058 (N_6058,N_4845,N_2321);
or U6059 (N_6059,N_4823,N_3200);
nand U6060 (N_6060,N_4303,N_4745);
xnor U6061 (N_6061,N_4004,N_2993);
xor U6062 (N_6062,N_2951,N_1088);
or U6063 (N_6063,N_809,N_3983);
xnor U6064 (N_6064,N_2165,N_2761);
or U6065 (N_6065,N_2964,N_1223);
or U6066 (N_6066,N_2369,N_1155);
xnor U6067 (N_6067,N_4454,N_1671);
or U6068 (N_6068,N_3553,N_2643);
and U6069 (N_6069,N_3012,N_644);
nor U6070 (N_6070,N_534,N_1982);
nor U6071 (N_6071,N_4312,N_3060);
or U6072 (N_6072,N_2818,N_3159);
nor U6073 (N_6073,N_4204,N_878);
and U6074 (N_6074,N_4593,N_4460);
and U6075 (N_6075,N_1576,N_2172);
nor U6076 (N_6076,N_3011,N_3085);
nor U6077 (N_6077,N_3128,N_553);
and U6078 (N_6078,N_1674,N_226);
xor U6079 (N_6079,N_3419,N_4109);
nor U6080 (N_6080,N_709,N_1567);
nand U6081 (N_6081,N_191,N_106);
nand U6082 (N_6082,N_1426,N_4157);
nand U6083 (N_6083,N_2587,N_278);
and U6084 (N_6084,N_1579,N_3808);
xnor U6085 (N_6085,N_3306,N_216);
nor U6086 (N_6086,N_1870,N_4666);
nor U6087 (N_6087,N_1258,N_3013);
nor U6088 (N_6088,N_250,N_1391);
nand U6089 (N_6089,N_1414,N_3000);
xor U6090 (N_6090,N_2480,N_555);
nor U6091 (N_6091,N_3388,N_716);
and U6092 (N_6092,N_4697,N_3944);
xor U6093 (N_6093,N_4916,N_211);
xor U6094 (N_6094,N_1376,N_379);
or U6095 (N_6095,N_1568,N_3605);
and U6096 (N_6096,N_3245,N_3452);
nand U6097 (N_6097,N_3481,N_2781);
nor U6098 (N_6098,N_2387,N_2257);
nor U6099 (N_6099,N_2878,N_330);
or U6100 (N_6100,N_1661,N_4865);
nand U6101 (N_6101,N_1753,N_1639);
nor U6102 (N_6102,N_4565,N_197);
xnor U6103 (N_6103,N_2218,N_3210);
nand U6104 (N_6104,N_519,N_360);
and U6105 (N_6105,N_3975,N_3287);
and U6106 (N_6106,N_1551,N_4537);
xnor U6107 (N_6107,N_696,N_3115);
nor U6108 (N_6108,N_1876,N_4867);
and U6109 (N_6109,N_3539,N_483);
nand U6110 (N_6110,N_4068,N_3347);
nor U6111 (N_6111,N_497,N_4490);
xnor U6112 (N_6112,N_4914,N_2568);
or U6113 (N_6113,N_1314,N_1298);
and U6114 (N_6114,N_283,N_2973);
or U6115 (N_6115,N_2811,N_2189);
xor U6116 (N_6116,N_359,N_1300);
nor U6117 (N_6117,N_3307,N_1911);
nor U6118 (N_6118,N_4332,N_2679);
nand U6119 (N_6119,N_3665,N_4883);
and U6120 (N_6120,N_995,N_1022);
nand U6121 (N_6121,N_43,N_3433);
nor U6122 (N_6122,N_3502,N_4618);
nor U6123 (N_6123,N_4379,N_1173);
xor U6124 (N_6124,N_4185,N_3758);
or U6125 (N_6125,N_3912,N_4348);
nor U6126 (N_6126,N_4462,N_4710);
or U6127 (N_6127,N_3774,N_1206);
and U6128 (N_6128,N_3554,N_1627);
and U6129 (N_6129,N_1505,N_2594);
nand U6130 (N_6130,N_3743,N_2245);
xor U6131 (N_6131,N_2441,N_4953);
nor U6132 (N_6132,N_801,N_634);
and U6133 (N_6133,N_2027,N_3036);
xor U6134 (N_6134,N_2660,N_3926);
and U6135 (N_6135,N_3562,N_2459);
xor U6136 (N_6136,N_802,N_2113);
nand U6137 (N_6137,N_3771,N_1985);
nor U6138 (N_6138,N_2610,N_223);
xor U6139 (N_6139,N_3517,N_3275);
nor U6140 (N_6140,N_2785,N_1131);
xnor U6141 (N_6141,N_2116,N_2325);
nand U6142 (N_6142,N_2680,N_3451);
xor U6143 (N_6143,N_561,N_4456);
nor U6144 (N_6144,N_1123,N_890);
nor U6145 (N_6145,N_4719,N_2940);
xnor U6146 (N_6146,N_3666,N_791);
nor U6147 (N_6147,N_4625,N_1136);
or U6148 (N_6148,N_140,N_4403);
xor U6149 (N_6149,N_3483,N_1084);
and U6150 (N_6150,N_2701,N_2280);
and U6151 (N_6151,N_2488,N_566);
nand U6152 (N_6152,N_1058,N_4669);
xnor U6153 (N_6153,N_1794,N_1592);
nor U6154 (N_6154,N_508,N_3362);
nand U6155 (N_6155,N_3241,N_2004);
nor U6156 (N_6156,N_905,N_3384);
nand U6157 (N_6157,N_3559,N_3767);
nor U6158 (N_6158,N_2704,N_623);
or U6159 (N_6159,N_1897,N_962);
nor U6160 (N_6160,N_998,N_2479);
or U6161 (N_6161,N_4774,N_4275);
nor U6162 (N_6162,N_1721,N_1715);
or U6163 (N_6163,N_868,N_236);
nor U6164 (N_6164,N_1160,N_10);
nor U6165 (N_6165,N_4881,N_2706);
or U6166 (N_6166,N_346,N_1865);
nand U6167 (N_6167,N_2578,N_2808);
and U6168 (N_6168,N_4172,N_3634);
nor U6169 (N_6169,N_951,N_4479);
nor U6170 (N_6170,N_2410,N_1756);
nand U6171 (N_6171,N_4055,N_1693);
and U6172 (N_6172,N_2711,N_1991);
nor U6173 (N_6173,N_480,N_4030);
nand U6174 (N_6174,N_3458,N_1279);
nand U6175 (N_6175,N_2455,N_4184);
xnor U6176 (N_6176,N_783,N_2093);
or U6177 (N_6177,N_4648,N_2829);
nand U6178 (N_6178,N_543,N_4227);
nor U6179 (N_6179,N_3393,N_2311);
xnor U6180 (N_6180,N_4422,N_1672);
nand U6181 (N_6181,N_3140,N_1023);
nand U6182 (N_6182,N_4529,N_1007);
nand U6183 (N_6183,N_1266,N_2834);
or U6184 (N_6184,N_4707,N_1760);
or U6185 (N_6185,N_3574,N_1696);
nand U6186 (N_6186,N_493,N_2717);
nand U6187 (N_6187,N_244,N_2152);
nor U6188 (N_6188,N_1044,N_4356);
and U6189 (N_6189,N_2547,N_4573);
nand U6190 (N_6190,N_1519,N_2895);
or U6191 (N_6191,N_4241,N_1578);
or U6192 (N_6192,N_781,N_228);
nand U6193 (N_6193,N_1460,N_3078);
or U6194 (N_6194,N_2053,N_4126);
and U6195 (N_6195,N_1472,N_4445);
xnor U6196 (N_6196,N_3369,N_4451);
nor U6197 (N_6197,N_2312,N_2295);
nor U6198 (N_6198,N_3321,N_1477);
nor U6199 (N_6199,N_1346,N_1716);
or U6200 (N_6200,N_2565,N_120);
nor U6201 (N_6201,N_1852,N_2802);
nand U6202 (N_6202,N_901,N_4643);
xnor U6203 (N_6203,N_3071,N_4125);
nand U6204 (N_6204,N_4545,N_2425);
nor U6205 (N_6205,N_2355,N_4582);
xor U6206 (N_6206,N_1918,N_4307);
and U6207 (N_6207,N_2276,N_4596);
and U6208 (N_6208,N_1327,N_4499);
xnor U6209 (N_6209,N_2353,N_3900);
xor U6210 (N_6210,N_101,N_1168);
nand U6211 (N_6211,N_3356,N_2323);
and U6212 (N_6212,N_2047,N_4655);
and U6213 (N_6213,N_4154,N_4703);
and U6214 (N_6214,N_3112,N_1701);
nor U6215 (N_6215,N_3043,N_3614);
and U6216 (N_6216,N_2524,N_425);
nand U6217 (N_6217,N_4857,N_4782);
nand U6218 (N_6218,N_2009,N_4523);
nor U6219 (N_6219,N_3932,N_1503);
nor U6220 (N_6220,N_680,N_695);
nor U6221 (N_6221,N_4331,N_1792);
xor U6222 (N_6222,N_2269,N_1597);
and U6223 (N_6223,N_987,N_2755);
xnor U6224 (N_6224,N_2158,N_720);
xnor U6225 (N_6225,N_2509,N_2545);
and U6226 (N_6226,N_1027,N_3868);
and U6227 (N_6227,N_338,N_1034);
nand U6228 (N_6228,N_4566,N_4659);
and U6229 (N_6229,N_1543,N_1175);
and U6230 (N_6230,N_3323,N_2157);
nand U6231 (N_6231,N_4952,N_2359);
nor U6232 (N_6232,N_2709,N_1196);
or U6233 (N_6233,N_3937,N_2693);
or U6234 (N_6234,N_4040,N_1154);
xnor U6235 (N_6235,N_4899,N_1428);
or U6236 (N_6236,N_3455,N_4497);
or U6237 (N_6237,N_0,N_916);
and U6238 (N_6238,N_1629,N_4432);
and U6239 (N_6239,N_725,N_146);
nand U6240 (N_6240,N_3424,N_2871);
nand U6241 (N_6241,N_2392,N_2797);
xor U6242 (N_6242,N_2947,N_3843);
or U6243 (N_6243,N_3472,N_2615);
and U6244 (N_6244,N_192,N_2751);
nor U6245 (N_6245,N_668,N_2904);
or U6246 (N_6246,N_4301,N_580);
and U6247 (N_6247,N_1854,N_1827);
or U6248 (N_6248,N_1892,N_1600);
nand U6249 (N_6249,N_4633,N_3949);
and U6250 (N_6250,N_4407,N_2463);
xor U6251 (N_6251,N_851,N_4135);
or U6252 (N_6252,N_957,N_2848);
and U6253 (N_6253,N_945,N_3088);
nand U6254 (N_6254,N_2159,N_3575);
nand U6255 (N_6255,N_4685,N_1879);
nor U6256 (N_6256,N_4470,N_2409);
nand U6257 (N_6257,N_4604,N_551);
nand U6258 (N_6258,N_4273,N_3031);
or U6259 (N_6259,N_4206,N_2499);
and U6260 (N_6260,N_3682,N_3298);
and U6261 (N_6261,N_387,N_189);
nor U6262 (N_6262,N_4486,N_364);
or U6263 (N_6263,N_1449,N_3358);
or U6264 (N_6264,N_1782,N_2259);
nand U6265 (N_6265,N_2628,N_2002);
and U6266 (N_6266,N_4790,N_4731);
xor U6267 (N_6267,N_1283,N_4712);
xor U6268 (N_6268,N_2897,N_3435);
nand U6269 (N_6269,N_1967,N_188);
and U6270 (N_6270,N_323,N_2531);
xnor U6271 (N_6271,N_1402,N_2402);
and U6272 (N_6272,N_1711,N_3957);
or U6273 (N_6273,N_1626,N_1261);
and U6274 (N_6274,N_2806,N_253);
nor U6275 (N_6275,N_4550,N_2133);
nand U6276 (N_6276,N_873,N_2087);
nor U6277 (N_6277,N_3761,N_514);
xnor U6278 (N_6278,N_4481,N_3915);
and U6279 (N_6279,N_3152,N_2908);
or U6280 (N_6280,N_4934,N_2998);
and U6281 (N_6281,N_640,N_406);
or U6282 (N_6282,N_1470,N_2682);
nor U6283 (N_6283,N_411,N_1636);
nand U6284 (N_6284,N_28,N_2695);
nor U6285 (N_6285,N_4878,N_2415);
and U6286 (N_6286,N_300,N_3141);
and U6287 (N_6287,N_1787,N_2130);
and U6288 (N_6288,N_4426,N_4935);
nor U6289 (N_6289,N_1570,N_711);
nor U6290 (N_6290,N_2599,N_1679);
nand U6291 (N_6291,N_3858,N_1634);
nor U6292 (N_6292,N_620,N_3202);
nor U6293 (N_6293,N_2580,N_885);
nand U6294 (N_6294,N_4764,N_973);
or U6295 (N_6295,N_4847,N_142);
nand U6296 (N_6296,N_4225,N_2030);
or U6297 (N_6297,N_1193,N_266);
and U6298 (N_6298,N_3883,N_1691);
nand U6299 (N_6299,N_3533,N_2378);
xnor U6300 (N_6300,N_1268,N_3407);
or U6301 (N_6301,N_64,N_2032);
xnor U6302 (N_6302,N_4421,N_1698);
xnor U6303 (N_6303,N_29,N_1296);
nor U6304 (N_6304,N_533,N_1534);
nand U6305 (N_6305,N_1665,N_2466);
nand U6306 (N_6306,N_4494,N_2076);
nand U6307 (N_6307,N_1157,N_950);
nor U6308 (N_6308,N_1318,N_2442);
and U6309 (N_6309,N_4634,N_3123);
nor U6310 (N_6310,N_2175,N_2010);
xor U6311 (N_6311,N_3701,N_4271);
and U6312 (N_6312,N_1968,N_3911);
xnor U6313 (N_6313,N_2839,N_449);
xor U6314 (N_6314,N_2447,N_4668);
nand U6315 (N_6315,N_2203,N_3982);
and U6316 (N_6316,N_25,N_1330);
nor U6317 (N_6317,N_4873,N_3657);
xor U6318 (N_6318,N_3664,N_42);
nand U6319 (N_6319,N_4283,N_3828);
nor U6320 (N_6320,N_4057,N_3376);
nand U6321 (N_6321,N_2518,N_4913);
nor U6322 (N_6322,N_3211,N_1142);
and U6323 (N_6323,N_3955,N_2844);
and U6324 (N_6324,N_2275,N_1737);
nor U6325 (N_6325,N_3877,N_2681);
nor U6326 (N_6326,N_3546,N_1308);
xor U6327 (N_6327,N_2180,N_1399);
nand U6328 (N_6328,N_116,N_679);
and U6329 (N_6329,N_3509,N_3168);
or U6330 (N_6330,N_2507,N_3094);
nor U6331 (N_6331,N_2525,N_3694);
and U6332 (N_6332,N_1746,N_4768);
xor U6333 (N_6333,N_1186,N_1466);
and U6334 (N_6334,N_4171,N_173);
or U6335 (N_6335,N_1530,N_4136);
and U6336 (N_6336,N_472,N_3095);
nand U6337 (N_6337,N_322,N_2367);
nor U6338 (N_6338,N_4717,N_4384);
nand U6339 (N_6339,N_1638,N_4285);
or U6340 (N_6340,N_842,N_4844);
or U6341 (N_6341,N_1009,N_3611);
and U6342 (N_6342,N_4103,N_1752);
xnor U6343 (N_6343,N_4049,N_574);
nand U6344 (N_6344,N_1083,N_712);
nand U6345 (N_6345,N_1312,N_4067);
nor U6346 (N_6346,N_2109,N_3120);
and U6347 (N_6347,N_3803,N_4202);
and U6348 (N_6348,N_3789,N_4843);
xnor U6349 (N_6349,N_2981,N_793);
and U6350 (N_6350,N_779,N_2349);
nor U6351 (N_6351,N_959,N_1068);
nor U6352 (N_6352,N_4942,N_2738);
xnor U6353 (N_6353,N_1808,N_931);
or U6354 (N_6354,N_3524,N_1473);
nand U6355 (N_6355,N_2946,N_893);
xor U6356 (N_6356,N_2913,N_4101);
and U6357 (N_6357,N_2056,N_4837);
or U6358 (N_6358,N_3038,N_2640);
nand U6359 (N_6359,N_3490,N_967);
nor U6360 (N_6360,N_4613,N_850);
or U6361 (N_6361,N_2216,N_1565);
or U6362 (N_6362,N_1755,N_2031);
or U6363 (N_6363,N_3756,N_4919);
and U6364 (N_6364,N_3576,N_2686);
xnor U6365 (N_6365,N_2300,N_774);
nor U6366 (N_6366,N_3564,N_2550);
nor U6367 (N_6367,N_2335,N_4997);
xor U6368 (N_6368,N_2842,N_694);
nor U6369 (N_6369,N_2063,N_2556);
xnor U6370 (N_6370,N_62,N_2241);
nor U6371 (N_6371,N_4777,N_1165);
xor U6372 (N_6372,N_2033,N_594);
and U6373 (N_6373,N_3030,N_2068);
xnor U6374 (N_6374,N_2969,N_2605);
xor U6375 (N_6375,N_2923,N_1328);
nand U6376 (N_6376,N_21,N_2807);
and U6377 (N_6377,N_1667,N_4607);
or U6378 (N_6378,N_652,N_4955);
or U6379 (N_6379,N_1953,N_1369);
xor U6380 (N_6380,N_1867,N_45);
nand U6381 (N_6381,N_3760,N_4577);
and U6382 (N_6382,N_4447,N_1948);
and U6383 (N_6383,N_3022,N_270);
nor U6384 (N_6384,N_4173,N_1502);
nor U6385 (N_6385,N_4975,N_2768);
or U6386 (N_6386,N_1031,N_1907);
nand U6387 (N_6387,N_4557,N_2461);
or U6388 (N_6388,N_942,N_4757);
and U6389 (N_6389,N_511,N_1335);
or U6390 (N_6390,N_4248,N_4622);
xor U6391 (N_6391,N_1766,N_1970);
or U6392 (N_6392,N_504,N_2013);
xnor U6393 (N_6393,N_4661,N_2313);
nand U6394 (N_6394,N_1781,N_807);
nand U6395 (N_6395,N_1690,N_4081);
and U6396 (N_6396,N_1965,N_4517);
and U6397 (N_6397,N_731,N_2705);
or U6398 (N_6398,N_4353,N_237);
nand U6399 (N_6399,N_4948,N_4748);
xor U6400 (N_6400,N_1704,N_4977);
and U6401 (N_6401,N_267,N_4446);
nor U6402 (N_6402,N_2584,N_3658);
nand U6403 (N_6403,N_4311,N_769);
and U6404 (N_6404,N_2401,N_88);
or U6405 (N_6405,N_1085,N_2095);
and U6406 (N_6406,N_176,N_3615);
or U6407 (N_6407,N_1074,N_2606);
or U6408 (N_6408,N_4972,N_3338);
xnor U6409 (N_6409,N_2638,N_3766);
or U6410 (N_6410,N_2329,N_2393);
nand U6411 (N_6411,N_141,N_2503);
nand U6412 (N_6412,N_4679,N_467);
xnor U6413 (N_6413,N_4343,N_3875);
and U6414 (N_6414,N_1993,N_4352);
nand U6415 (N_6415,N_3082,N_4186);
and U6416 (N_6416,N_2889,N_3367);
and U6417 (N_6417,N_2089,N_2872);
xor U6418 (N_6418,N_1933,N_1412);
nor U6419 (N_6419,N_2585,N_737);
and U6420 (N_6420,N_4164,N_1538);
or U6421 (N_6421,N_2247,N_2766);
and U6422 (N_6422,N_1217,N_4207);
and U6423 (N_6423,N_3413,N_4066);
nor U6424 (N_6424,N_2386,N_4393);
and U6425 (N_6425,N_2653,N_1405);
or U6426 (N_6426,N_2736,N_3139);
nor U6427 (N_6427,N_4104,N_1726);
and U6428 (N_6428,N_1586,N_896);
or U6429 (N_6429,N_590,N_1037);
xor U6430 (N_6430,N_856,N_4385);
and U6431 (N_6431,N_318,N_1286);
nor U6432 (N_6432,N_1166,N_1018);
nand U6433 (N_6433,N_2470,N_947);
nor U6434 (N_6434,N_4538,N_1417);
or U6435 (N_6435,N_707,N_4281);
nor U6436 (N_6436,N_3814,N_488);
nand U6437 (N_6437,N_2446,N_825);
nor U6438 (N_6438,N_3565,N_4946);
or U6439 (N_6439,N_3627,N_4429);
or U6440 (N_6440,N_4197,N_463);
nor U6441 (N_6441,N_2957,N_4996);
or U6442 (N_6442,N_3947,N_4296);
or U6443 (N_6443,N_22,N_608);
or U6444 (N_6444,N_1063,N_3344);
or U6445 (N_6445,N_154,N_3569);
and U6446 (N_6446,N_2486,N_4765);
and U6447 (N_6447,N_815,N_3924);
and U6448 (N_6448,N_4749,N_2320);
nand U6449 (N_6449,N_175,N_2861);
and U6450 (N_6450,N_4861,N_4013);
nor U6451 (N_6451,N_782,N_2798);
nor U6452 (N_6452,N_3066,N_3908);
xor U6453 (N_6453,N_4276,N_3215);
or U6454 (N_6454,N_85,N_4265);
or U6455 (N_6455,N_3277,N_4391);
nand U6456 (N_6456,N_2707,N_344);
or U6457 (N_6457,N_4586,N_4739);
nand U6458 (N_6458,N_3622,N_4074);
nand U6459 (N_6459,N_4253,N_3913);
nor U6460 (N_6460,N_2535,N_290);
nand U6461 (N_6461,N_1635,N_1433);
or U6462 (N_6462,N_683,N_3289);
nor U6463 (N_6463,N_675,N_1100);
or U6464 (N_6464,N_3429,N_470);
or U6465 (N_6465,N_1607,N_1253);
nand U6466 (N_6466,N_2112,N_2162);
nor U6467 (N_6467,N_404,N_3423);
or U6468 (N_6468,N_3712,N_964);
nor U6469 (N_6469,N_378,N_3702);
xor U6470 (N_6470,N_3504,N_3928);
nand U6471 (N_6471,N_4994,N_3632);
nor U6472 (N_6472,N_4315,N_1599);
or U6473 (N_6473,N_4026,N_1065);
nand U6474 (N_6474,N_2448,N_1922);
and U6475 (N_6475,N_1250,N_1863);
nor U6476 (N_6476,N_1581,N_937);
xor U6477 (N_6477,N_185,N_3166);
xor U6478 (N_6478,N_899,N_2227);
or U6479 (N_6479,N_2021,N_4228);
nand U6480 (N_6480,N_2398,N_4449);
and U6481 (N_6481,N_3061,N_310);
nand U6482 (N_6482,N_3281,N_736);
and U6483 (N_6483,N_1809,N_1097);
nor U6484 (N_6484,N_90,N_2150);
nor U6485 (N_6485,N_3383,N_727);
and U6486 (N_6486,N_1240,N_4183);
nor U6487 (N_6487,N_3818,N_3740);
and U6488 (N_6488,N_3684,N_104);
nor U6489 (N_6489,N_1103,N_4628);
nor U6490 (N_6490,N_818,N_5);
and U6491 (N_6491,N_1675,N_4372);
nand U6492 (N_6492,N_1905,N_4230);
nor U6493 (N_6493,N_826,N_4689);
xor U6494 (N_6494,N_4987,N_670);
xnor U6495 (N_6495,N_3819,N_3857);
or U6496 (N_6496,N_4609,N_4201);
or U6497 (N_6497,N_4024,N_1406);
or U6498 (N_6498,N_2237,N_2201);
xnor U6499 (N_6499,N_3889,N_4350);
xnor U6500 (N_6500,N_1204,N_2791);
or U6501 (N_6501,N_1840,N_3856);
xnor U6502 (N_6502,N_2471,N_4858);
or U6503 (N_6503,N_1783,N_3599);
or U6504 (N_6504,N_3820,N_2602);
and U6505 (N_6505,N_2207,N_4614);
xor U6506 (N_6506,N_4415,N_4849);
nor U6507 (N_6507,N_3310,N_638);
and U6508 (N_6508,N_4266,N_3328);
xnor U6509 (N_6509,N_4840,N_320);
xnor U6510 (N_6510,N_2574,N_3644);
xor U6511 (N_6511,N_2619,N_71);
nor U6512 (N_6512,N_2306,N_3117);
nand U6513 (N_6513,N_2620,N_2986);
and U6514 (N_6514,N_2341,N_413);
and U6515 (N_6515,N_1174,N_4835);
or U6516 (N_6516,N_4457,N_3160);
or U6517 (N_6517,N_724,N_4073);
or U6518 (N_6518,N_3077,N_3809);
and U6519 (N_6519,N_847,N_2475);
and U6520 (N_6520,N_4174,N_2645);
xor U6521 (N_6521,N_3994,N_3791);
and U6522 (N_6522,N_3045,N_4547);
and U6523 (N_6523,N_452,N_3671);
nor U6524 (N_6524,N_1734,N_2035);
nand U6525 (N_6525,N_918,N_4330);
xnor U6526 (N_6526,N_1754,N_4892);
xor U6527 (N_6527,N_4287,N_3351);
xnor U6528 (N_6528,N_1438,N_460);
nand U6529 (N_6529,N_3155,N_4199);
xor U6530 (N_6530,N_3778,N_2812);
or U6531 (N_6531,N_1680,N_1866);
nor U6532 (N_6532,N_4879,N_4110);
nor U6533 (N_6533,N_871,N_4129);
xor U6534 (N_6534,N_4069,N_242);
nand U6535 (N_6535,N_1082,N_750);
and U6536 (N_6536,N_4404,N_3686);
and U6537 (N_6537,N_921,N_1611);
and U6538 (N_6538,N_1344,N_1712);
nand U6539 (N_6539,N_542,N_129);
xnor U6540 (N_6540,N_2925,N_1257);
and U6541 (N_6541,N_2671,N_222);
or U6542 (N_6542,N_1317,N_3884);
nor U6543 (N_6543,N_108,N_4591);
nor U6544 (N_6544,N_3348,N_2094);
and U6545 (N_6545,N_4102,N_977);
xnor U6546 (N_6546,N_4308,N_3074);
or U6547 (N_6547,N_1761,N_1158);
or U6548 (N_6548,N_286,N_179);
nand U6549 (N_6549,N_4151,N_3224);
nand U6550 (N_6550,N_4145,N_4510);
nand U6551 (N_6551,N_1980,N_4416);
and U6552 (N_6552,N_274,N_4687);
and U6553 (N_6553,N_386,N_304);
and U6554 (N_6554,N_2489,N_1914);
and U6555 (N_6555,N_4509,N_554);
nand U6556 (N_6556,N_2331,N_4008);
nand U6557 (N_6557,N_4406,N_2371);
and U6558 (N_6558,N_4542,N_4045);
and U6559 (N_6559,N_4533,N_4665);
and U6560 (N_6560,N_2753,N_2043);
nor U6561 (N_6561,N_2712,N_1394);
or U6562 (N_6562,N_3317,N_3934);
nand U6563 (N_6563,N_1736,N_4474);
nor U6564 (N_6564,N_584,N_1590);
nand U6565 (N_6565,N_4112,N_1309);
and U6566 (N_6566,N_1935,N_2086);
xor U6567 (N_6567,N_2016,N_3096);
and U6568 (N_6568,N_1459,N_3579);
or U6569 (N_6569,N_1382,N_1059);
and U6570 (N_6570,N_3109,N_4051);
or U6571 (N_6571,N_1609,N_4214);
or U6572 (N_6572,N_4498,N_502);
nor U6573 (N_6573,N_4012,N_2805);
and U6574 (N_6574,N_1497,N_863);
nor U6575 (N_6575,N_3183,N_2978);
nand U6576 (N_6576,N_2075,N_205);
xor U6577 (N_6577,N_4725,N_3286);
nand U6578 (N_6578,N_2343,N_3999);
xor U6579 (N_6579,N_908,N_4568);
nand U6580 (N_6580,N_3714,N_2271);
xnor U6581 (N_6581,N_138,N_435);
nand U6582 (N_6582,N_1617,N_2431);
xnor U6583 (N_6583,N_1396,N_3411);
xor U6584 (N_6584,N_2733,N_2417);
xnor U6585 (N_6585,N_2437,N_3216);
and U6586 (N_6586,N_2885,N_4690);
nor U6587 (N_6587,N_4522,N_867);
nand U6588 (N_6588,N_1975,N_2319);
nor U6589 (N_6589,N_148,N_1828);
and U6590 (N_6590,N_4632,N_658);
nand U6591 (N_6591,N_2786,N_3158);
or U6592 (N_6592,N_2996,N_4819);
and U6593 (N_6593,N_913,N_777);
nor U6594 (N_6594,N_393,N_2789);
and U6595 (N_6595,N_3669,N_3374);
nand U6596 (N_6596,N_307,N_507);
and U6597 (N_6597,N_3193,N_1504);
or U6598 (N_6598,N_2222,N_2067);
and U6599 (N_6599,N_974,N_3489);
nor U6600 (N_6600,N_337,N_2373);
or U6601 (N_6601,N_82,N_396);
xor U6602 (N_6602,N_3916,N_2915);
nor U6603 (N_6603,N_3907,N_4317);
nor U6604 (N_6604,N_1432,N_2914);
or U6605 (N_6605,N_2374,N_4700);
nor U6606 (N_6606,N_604,N_1105);
xor U6607 (N_6607,N_3434,N_4279);
and U6608 (N_6608,N_3854,N_602);
and U6609 (N_6609,N_1786,N_1275);
nor U6610 (N_6610,N_2801,N_2429);
nor U6611 (N_6611,N_2297,N_2905);
or U6612 (N_6612,N_4302,N_2363);
and U6613 (N_6613,N_1321,N_3759);
nand U6614 (N_6614,N_303,N_3689);
and U6615 (N_6615,N_2242,N_2236);
nor U6616 (N_6616,N_2011,N_3969);
xnor U6617 (N_6617,N_183,N_2992);
and U6618 (N_6618,N_4794,N_382);
and U6619 (N_6619,N_1742,N_795);
xor U6620 (N_6620,N_2659,N_3391);
or U6621 (N_6621,N_799,N_1403);
xnor U6622 (N_6622,N_2235,N_700);
or U6623 (N_6623,N_1768,N_682);
and U6624 (N_6624,N_4131,N_593);
nand U6625 (N_6625,N_1571,N_1195);
or U6626 (N_6626,N_510,N_4781);
nor U6627 (N_6627,N_3892,N_114);
nand U6628 (N_6628,N_4247,N_4651);
or U6629 (N_6629,N_3041,N_3678);
nor U6630 (N_6630,N_3454,N_991);
nor U6631 (N_6631,N_4464,N_1984);
nor U6632 (N_6632,N_298,N_3558);
nor U6633 (N_6633,N_3231,N_297);
nor U6634 (N_6634,N_1583,N_4233);
nor U6635 (N_6635,N_2408,N_4945);
and U6636 (N_6636,N_1956,N_367);
xor U6637 (N_6637,N_3567,N_3207);
nand U6638 (N_6638,N_1910,N_3738);
nand U6639 (N_6639,N_4699,N_3361);
nand U6640 (N_6640,N_3285,N_3410);
or U6641 (N_6641,N_76,N_822);
nand U6642 (N_6642,N_4190,N_3951);
xnor U6643 (N_6643,N_4089,N_4133);
or U6644 (N_6644,N_2464,N_4959);
nand U6645 (N_6645,N_3941,N_4784);
xnor U6646 (N_6646,N_1232,N_2663);
nand U6647 (N_6647,N_3812,N_4875);
nand U6648 (N_6648,N_2135,N_678);
or U6649 (N_6649,N_2347,N_1526);
or U6650 (N_6650,N_4738,N_3901);
nand U6651 (N_6651,N_59,N_3457);
and U6652 (N_6652,N_3659,N_4885);
nor U6653 (N_6653,N_2939,N_1316);
or U6654 (N_6654,N_2060,N_4484);
xnor U6655 (N_6655,N_2865,N_4570);
and U6656 (N_6656,N_2855,N_1073);
xnor U6657 (N_6657,N_128,N_4640);
or U6658 (N_6658,N_315,N_3656);
or U6659 (N_6659,N_3917,N_1117);
and U6660 (N_6660,N_1188,N_3133);
or U6661 (N_6661,N_2149,N_2255);
nor U6662 (N_6662,N_2209,N_3055);
or U6663 (N_6663,N_759,N_1740);
xor U6664 (N_6664,N_1796,N_225);
xor U6665 (N_6665,N_3594,N_3024);
nor U6666 (N_6666,N_2656,N_1241);
nor U6667 (N_6667,N_4159,N_980);
nand U6668 (N_6668,N_3698,N_2795);
nand U6669 (N_6669,N_3505,N_1041);
or U6670 (N_6670,N_3876,N_4561);
or U6671 (N_6671,N_4305,N_3584);
nand U6672 (N_6672,N_427,N_2243);
or U6673 (N_6673,N_2228,N_558);
nand U6674 (N_6674,N_2292,N_249);
and U6675 (N_6675,N_3431,N_971);
xnor U6676 (N_6676,N_3836,N_4730);
xor U6677 (N_6677,N_2911,N_3956);
and U6678 (N_6678,N_3453,N_4795);
nor U6679 (N_6679,N_4980,N_1616);
or U6680 (N_6680,N_3415,N_1176);
and U6681 (N_6681,N_1026,N_3148);
and U6682 (N_6682,N_570,N_3387);
or U6683 (N_6683,N_4469,N_954);
nor U6684 (N_6684,N_4123,N_426);
nand U6685 (N_6685,N_3178,N_2196);
and U6686 (N_6686,N_1819,N_1162);
or U6687 (N_6687,N_1894,N_2554);
nand U6688 (N_6688,N_2493,N_4546);
nor U6689 (N_6689,N_1352,N_3272);
nand U6690 (N_6690,N_1510,N_757);
and U6691 (N_6691,N_876,N_2726);
and U6692 (N_6692,N_626,N_4144);
xnor U6693 (N_6693,N_3788,N_4062);
nand U6694 (N_6694,N_4489,N_969);
nor U6695 (N_6695,N_2384,N_2700);
and U6696 (N_6696,N_75,N_2350);
nand U6697 (N_6697,N_1868,N_1108);
nor U6698 (N_6698,N_1974,N_1375);
nand U6699 (N_6699,N_2248,N_1869);
or U6700 (N_6700,N_2530,N_2439);
xnor U6701 (N_6701,N_4684,N_857);
nand U6702 (N_6702,N_3247,N_4539);
and U6703 (N_6703,N_520,N_701);
nand U6704 (N_6704,N_2945,N_326);
and U6705 (N_6705,N_4834,N_3616);
xnor U6706 (N_6706,N_4992,N_1946);
xor U6707 (N_6707,N_3899,N_674);
nand U6708 (N_6708,N_2744,N_2022);
xnor U6709 (N_6709,N_2066,N_1452);
nor U6710 (N_6710,N_150,N_4856);
xnor U6711 (N_6711,N_4176,N_4915);
and U6712 (N_6712,N_2199,N_4704);
xor U6713 (N_6713,N_3597,N_143);
or U6714 (N_6714,N_94,N_4114);
xor U6715 (N_6715,N_4077,N_4071);
and U6716 (N_6716,N_238,N_4022);
xnor U6717 (N_6717,N_541,N_1839);
nand U6718 (N_6718,N_2452,N_3736);
xnor U6719 (N_6719,N_2821,N_1329);
nand U6720 (N_6720,N_4793,N_339);
and U6721 (N_6721,N_2961,N_12);
nor U6722 (N_6722,N_1670,N_273);
nand U6723 (N_6723,N_1845,N_2642);
nand U6724 (N_6724,N_4010,N_3648);
nand U6725 (N_6725,N_688,N_333);
nand U6726 (N_6726,N_3635,N_1682);
xnor U6727 (N_6727,N_1855,N_2774);
and U6728 (N_6728,N_3271,N_2453);
nand U6729 (N_6729,N_1659,N_70);
xor U6730 (N_6730,N_3731,N_1478);
and U6731 (N_6731,N_2081,N_2161);
or U6732 (N_6732,N_4521,N_4930);
nor U6733 (N_6733,N_4989,N_1000);
or U6734 (N_6734,N_2982,N_3535);
or U6735 (N_6735,N_3706,N_4888);
nor U6736 (N_6736,N_548,N_2134);
xor U6737 (N_6737,N_568,N_3602);
nand U6738 (N_6738,N_321,N_3198);
nor U6739 (N_6739,N_2987,N_3528);
xnor U6740 (N_6740,N_390,N_4031);
nand U6741 (N_6741,N_4986,N_420);
and U6742 (N_6742,N_3861,N_1210);
xor U6743 (N_6743,N_1826,N_1889);
and U6744 (N_6744,N_3570,N_4327);
and U6745 (N_6745,N_2266,N_2502);
nand U6746 (N_6746,N_2984,N_1124);
xnor U6747 (N_6747,N_309,N_738);
or U6748 (N_6748,N_4543,N_4805);
nand U6749 (N_6749,N_2771,N_4419);
and U6750 (N_6750,N_2696,N_34);
nand U6751 (N_6751,N_3119,N_1559);
and U6752 (N_6752,N_1535,N_2282);
nand U6753 (N_6753,N_517,N_4544);
xor U6754 (N_6754,N_2896,N_4152);
xnor U6755 (N_6755,N_1445,N_1747);
xor U6756 (N_6756,N_4,N_4284);
xnor U6757 (N_6757,N_3227,N_2910);
or U6758 (N_6758,N_2070,N_358);
nor U6759 (N_6759,N_2666,N_662);
xnor U6760 (N_6760,N_665,N_3687);
xnor U6761 (N_6761,N_4178,N_3249);
nor U6762 (N_6762,N_1821,N_2760);
and U6763 (N_6763,N_3583,N_2607);
and U6764 (N_6764,N_3964,N_1050);
and U6765 (N_6765,N_1560,N_1265);
or U6766 (N_6766,N_4122,N_1649);
and U6767 (N_6767,N_3334,N_2187);
or U6768 (N_6768,N_14,N_3717);
nor U6769 (N_6769,N_4189,N_1537);
or U6770 (N_6770,N_2979,N_4359);
xnor U6771 (N_6771,N_1119,N_478);
nand U6772 (N_6772,N_2634,N_1684);
or U6773 (N_6773,N_3498,N_2098);
nor U6774 (N_6774,N_441,N_3763);
and U6775 (N_6775,N_4963,N_2498);
or U6776 (N_6776,N_1093,N_3977);
and U6777 (N_6777,N_565,N_4709);
nor U6778 (N_6778,N_1228,N_2652);
and U6779 (N_6779,N_1728,N_2988);
nand U6780 (N_6780,N_1580,N_3070);
or U6781 (N_6781,N_884,N_607);
nand U6782 (N_6782,N_3881,N_93);
and U6783 (N_6783,N_2675,N_1233);
xor U6784 (N_6784,N_1475,N_3794);
nor U6785 (N_6785,N_764,N_3408);
and U6786 (N_6786,N_369,N_2416);
nor U6787 (N_6787,N_2758,N_1775);
and U6788 (N_6788,N_2477,N_4702);
nor U6789 (N_6789,N_3053,N_3718);
nor U6790 (N_6790,N_3643,N_4220);
nand U6791 (N_6791,N_1362,N_2975);
nor U6792 (N_6792,N_588,N_4444);
or U6793 (N_6793,N_4260,N_2971);
xnor U6794 (N_6794,N_742,N_1748);
xor U6795 (N_6795,N_862,N_2399);
nand U6796 (N_6796,N_1795,N_3130);
nor U6797 (N_6797,N_3190,N_4143);
or U6798 (N_6798,N_2179,N_2125);
nand U6799 (N_6799,N_1812,N_2857);
nand U6800 (N_6800,N_1351,N_3674);
and U6801 (N_6801,N_1945,N_708);
and U6802 (N_6802,N_2283,N_4193);
nand U6803 (N_6803,N_4999,N_556);
nand U6804 (N_6804,N_2217,N_1150);
and U6805 (N_6805,N_2289,N_1727);
xnor U6806 (N_6806,N_3638,N_105);
or U6807 (N_6807,N_934,N_3232);
nand U6808 (N_6808,N_295,N_609);
and U6809 (N_6809,N_4951,N_4880);
nor U6810 (N_6810,N_4169,N_1951);
nand U6811 (N_6811,N_3491,N_3163);
nor U6812 (N_6812,N_1249,N_787);
and U6813 (N_6813,N_3475,N_1550);
nor U6814 (N_6814,N_2882,N_1858);
xor U6815 (N_6815,N_254,N_1898);
nand U6816 (N_6816,N_3326,N_3707);
and U6817 (N_6817,N_1334,N_2155);
nand U6818 (N_6818,N_4862,N_4274);
xnor U6819 (N_6819,N_4859,N_1384);
nor U6820 (N_6820,N_4727,N_4020);
xor U6821 (N_6821,N_2184,N_4148);
xnor U6822 (N_6822,N_1363,N_343);
nor U6823 (N_6823,N_3536,N_3966);
xor U6824 (N_6824,N_159,N_4120);
nor U6825 (N_6825,N_3681,N_4325);
or U6826 (N_6826,N_3598,N_2884);
xnor U6827 (N_6827,N_2354,N_3440);
or U6828 (N_6828,N_3325,N_363);
or U6829 (N_6829,N_3670,N_723);
xnor U6830 (N_6830,N_4374,N_3607);
xor U6831 (N_6831,N_3214,N_2617);
nand U6832 (N_6832,N_4203,N_4842);
or U6833 (N_6833,N_4846,N_1310);
or U6834 (N_6834,N_4629,N_3863);
xnor U6835 (N_6835,N_4671,N_4019);
or U6836 (N_6836,N_2383,N_1887);
nor U6837 (N_6837,N_837,N_610);
and U6838 (N_6838,N_3745,N_4722);
or U6839 (N_6839,N_156,N_4512);
nor U6840 (N_6840,N_1247,N_895);
nor U6841 (N_6841,N_1114,N_484);
or U6842 (N_6842,N_3294,N_3217);
or U6843 (N_6843,N_4681,N_4177);
nor U6844 (N_6844,N_2702,N_3151);
nor U6845 (N_6845,N_4496,N_961);
nand U6846 (N_6846,N_2003,N_923);
nor U6847 (N_6847,N_2299,N_496);
xor U6848 (N_6848,N_454,N_1663);
and U6849 (N_6849,N_4397,N_4968);
and U6850 (N_6850,N_1872,N_3377);
nor U6851 (N_6851,N_704,N_819);
nand U6852 (N_6852,N_4361,N_165);
and U6853 (N_6853,N_3746,N_525);
nor U6854 (N_6854,N_882,N_4263);
nand U6855 (N_6855,N_421,N_2279);
nand U6856 (N_6856,N_747,N_44);
nor U6857 (N_6857,N_1145,N_4128);
xnor U6858 (N_6858,N_2875,N_1251);
nand U6859 (N_6859,N_3755,N_3751);
xor U6860 (N_6860,N_3723,N_3257);
and U6861 (N_6861,N_1464,N_3873);
or U6862 (N_6862,N_4212,N_1552);
nand U6863 (N_6863,N_1972,N_2985);
xor U6864 (N_6864,N_730,N_92);
nand U6865 (N_6865,N_4138,N_2050);
xnor U6866 (N_6866,N_2336,N_2322);
and U6867 (N_6867,N_4222,N_4673);
or U6868 (N_6868,N_118,N_4964);
or U6869 (N_6869,N_434,N_1793);
or U6870 (N_6870,N_2501,N_1713);
nand U6871 (N_6871,N_1030,N_3825);
xnor U6872 (N_6872,N_2163,N_2534);
or U6873 (N_6873,N_3555,N_2573);
and U6874 (N_6874,N_1699,N_4562);
nor U6875 (N_6875,N_3953,N_2513);
nor U6876 (N_6876,N_68,N_3925);
nand U6877 (N_6877,N_2268,N_3510);
nor U6878 (N_6878,N_4744,N_4063);
and U6879 (N_6879,N_1216,N_4553);
nand U6880 (N_6880,N_2208,N_4435);
and U6881 (N_6881,N_2182,N_2794);
and U6882 (N_6882,N_4156,N_3219);
nor U6883 (N_6883,N_648,N_4437);
or U6884 (N_6884,N_215,N_1213);
or U6885 (N_6885,N_4342,N_4323);
xor U6886 (N_6886,N_3265,N_3971);
xor U6887 (N_6887,N_1090,N_1021);
and U6888 (N_6888,N_3728,N_1016);
and U6889 (N_6889,N_458,N_647);
nand U6890 (N_6890,N_2024,N_4907);
xor U6891 (N_6891,N_2967,N_1263);
nand U6892 (N_6892,N_3726,N_2687);
or U6893 (N_6893,N_3302,N_2767);
xnor U6894 (N_6894,N_2427,N_3091);
and U6895 (N_6895,N_531,N_180);
nand U6896 (N_6896,N_1467,N_2537);
or U6897 (N_6897,N_4387,N_1619);
xnor U6898 (N_6898,N_4042,N_789);
xor U6899 (N_6899,N_2780,N_1147);
or U6900 (N_6900,N_773,N_4116);
and U6901 (N_6901,N_4910,N_124);
and U6902 (N_6902,N_612,N_1833);
nor U6903 (N_6903,N_2776,N_3586);
and U6904 (N_6904,N_3697,N_2443);
nand U6905 (N_6905,N_3316,N_3156);
xnor U6906 (N_6906,N_4300,N_512);
or U6907 (N_6907,N_3894,N_859);
and U6908 (N_6908,N_4094,N_1256);
or U6909 (N_6909,N_3259,N_461);
nand U6910 (N_6910,N_691,N_3049);
nor U6911 (N_6911,N_2167,N_521);
xnor U6912 (N_6912,N_3872,N_1107);
nand U6913 (N_6913,N_184,N_4200);
and U6914 (N_6914,N_3571,N_4246);
nor U6915 (N_6915,N_821,N_1631);
xor U6916 (N_6916,N_145,N_4480);
or U6917 (N_6917,N_828,N_2462);
or U6918 (N_6918,N_766,N_3626);
xor U6919 (N_6919,N_285,N_212);
nor U6920 (N_6920,N_2129,N_2673);
xnor U6921 (N_6921,N_1390,N_4897);
nor U6922 (N_6922,N_3314,N_788);
xnor U6923 (N_6923,N_2720,N_4032);
nand U6924 (N_6924,N_1337,N_3443);
nand U6925 (N_6925,N_2757,N_4097);
nand U6926 (N_6926,N_2145,N_3864);
xnor U6927 (N_6927,N_1987,N_2097);
xnor U6928 (N_6928,N_4599,N_4380);
or U6929 (N_6929,N_1623,N_660);
xor U6930 (N_6930,N_4894,N_178);
nor U6931 (N_6931,N_4715,N_2397);
nor U6932 (N_6932,N_4686,N_2745);
xnor U6933 (N_6933,N_1137,N_1977);
xor U6934 (N_6934,N_1776,N_4134);
xor U6935 (N_6935,N_4473,N_4788);
xor U6936 (N_6936,N_133,N_4769);
nor U6937 (N_6937,N_1011,N_4853);
xor U6938 (N_6938,N_2814,N_4459);
nor U6939 (N_6939,N_2926,N_2231);
nor U6940 (N_6940,N_1401,N_2444);
and U6941 (N_6941,N_3194,N_3386);
or U6942 (N_6942,N_1536,N_1484);
or U6943 (N_6943,N_134,N_4571);
xor U6944 (N_6944,N_692,N_4938);
nor U6945 (N_6945,N_2365,N_3375);
xor U6946 (N_6946,N_4278,N_464);
nand U6947 (N_6947,N_3754,N_2639);
nand U6948 (N_6948,N_448,N_3905);
nand U6949 (N_6949,N_4832,N_3380);
or U6950 (N_6950,N_281,N_2483);
xnor U6951 (N_6951,N_4810,N_2229);
or U6952 (N_6952,N_3212,N_4132);
nor U6953 (N_6953,N_3797,N_3704);
and U6954 (N_6954,N_4877,N_3464);
or U6955 (N_6955,N_2361,N_2542);
nor U6956 (N_6956,N_2119,N_126);
nor U6957 (N_6957,N_4410,N_439);
and U6958 (N_6958,N_1901,N_628);
or U6959 (N_6959,N_1739,N_3677);
nand U6960 (N_6960,N_4321,N_3897);
or U6961 (N_6961,N_4678,N_1132);
xor U6962 (N_6962,N_2368,N_1325);
or U6963 (N_6963,N_4602,N_1070);
nor U6964 (N_6964,N_2019,N_3596);
nand U6965 (N_6965,N_2073,N_1561);
and U6966 (N_6966,N_2835,N_1603);
or U6967 (N_6967,N_2514,N_3974);
or U6968 (N_6968,N_2517,N_3936);
nor U6969 (N_6969,N_3826,N_2077);
or U6970 (N_6970,N_2099,N_1602);
nor U6971 (N_6971,N_865,N_1133);
or U6972 (N_6972,N_1043,N_2583);
xor U6973 (N_6973,N_576,N_3253);
xor U6974 (N_6974,N_3373,N_257);
and U6975 (N_6975,N_3154,N_2357);
nor U6976 (N_6976,N_4458,N_2285);
nand U6977 (N_6977,N_1307,N_2799);
nand U6978 (N_6978,N_879,N_1688);
xor U6979 (N_6979,N_444,N_490);
xor U6980 (N_6980,N_4711,N_3162);
nor U6981 (N_6981,N_3715,N_160);
nand U6982 (N_6982,N_3813,N_4559);
or U6983 (N_6983,N_1595,N_3672);
xnor U6984 (N_6984,N_988,N_2327);
nand U6985 (N_6985,N_4378,N_3963);
nor U6986 (N_6986,N_1427,N_2942);
and U6987 (N_6987,N_4574,N_258);
or U6988 (N_6988,N_2223,N_3845);
nand U6989 (N_6989,N_2205,N_1885);
or U6990 (N_6990,N_697,N_107);
or U6991 (N_6991,N_4549,N_453);
xor U6992 (N_6992,N_383,N_4028);
nand U6993 (N_6993,N_1368,N_1366);
nor U6994 (N_6994,N_1893,N_2389);
nor U6995 (N_6995,N_95,N_416);
nand U6996 (N_6996,N_4003,N_3092);
and U6997 (N_6997,N_4983,N_1013);
nand U6998 (N_6998,N_505,N_762);
or U6999 (N_6999,N_3090,N_2136);
xor U7000 (N_7000,N_227,N_3806);
or U7001 (N_7001,N_976,N_2045);
xor U7002 (N_7002,N_3752,N_1120);
nand U7003 (N_7003,N_4256,N_4054);
nor U7004 (N_7004,N_3186,N_4011);
nand U7005 (N_7005,N_677,N_2690);
and U7006 (N_7006,N_2048,N_3303);
xnor U7007 (N_7007,N_2090,N_4262);
xnor U7008 (N_7008,N_1252,N_2177);
or U7009 (N_7009,N_3606,N_2604);
nor U7010 (N_7010,N_3188,N_3251);
and U7011 (N_7011,N_3072,N_284);
or U7012 (N_7012,N_1104,N_2375);
and U7013 (N_7013,N_72,N_4007);
xor U7014 (N_7014,N_51,N_1983);
xnor U7015 (N_7015,N_4142,N_2064);
nand U7016 (N_7016,N_2670,N_289);
xnor U7017 (N_7017,N_2698,N_2980);
xnor U7018 (N_7018,N_2445,N_537);
or U7019 (N_7019,N_2632,N_2069);
nand U7020 (N_7020,N_845,N_4166);
or U7021 (N_7021,N_1303,N_331);
nand U7022 (N_7022,N_4956,N_1882);
xnor U7023 (N_7023,N_1811,N_4226);
and U7024 (N_7024,N_928,N_4349);
and U7025 (N_7025,N_3783,N_2543);
or U7026 (N_7026,N_3340,N_1419);
nor U7027 (N_7027,N_4095,N_2827);
or U7028 (N_7028,N_2612,N_4998);
nor U7029 (N_7029,N_1239,N_2277);
nor U7030 (N_7030,N_1340,N_715);
xor U7031 (N_7031,N_3449,N_375);
and U7032 (N_7032,N_1912,N_1903);
xor U7033 (N_7033,N_1183,N_4931);
nor U7034 (N_7034,N_994,N_3487);
xor U7035 (N_7035,N_4563,N_3646);
or U7036 (N_7036,N_1883,N_1278);
and U7037 (N_7037,N_443,N_2596);
and U7038 (N_7038,N_1407,N_3853);
or U7039 (N_7039,N_4289,N_1498);
xnor U7040 (N_7040,N_4921,N_941);
and U7041 (N_7041,N_1029,N_3613);
and U7042 (N_7042,N_4870,N_3264);
nand U7043 (N_7043,N_2833,N_2667);
nor U7044 (N_7044,N_550,N_1192);
and U7045 (N_7045,N_2190,N_1274);
nand U7046 (N_7046,N_938,N_4244);
or U7047 (N_7047,N_3138,N_1214);
or U7048 (N_7048,N_3739,N_4649);
and U7049 (N_7049,N_2473,N_2037);
or U7050 (N_7050,N_1582,N_348);
and U7051 (N_7051,N_417,N_1485);
or U7052 (N_7052,N_2782,N_121);
nor U7053 (N_7053,N_4579,N_1507);
nor U7054 (N_7054,N_46,N_3976);
nor U7055 (N_7055,N_3581,N_3732);
or U7056 (N_7056,N_3544,N_672);
or U7057 (N_7057,N_1371,N_2803);
or U7058 (N_7058,N_3008,N_186);
xor U7059 (N_7059,N_3920,N_3519);
xor U7060 (N_7060,N_2999,N_2862);
nand U7061 (N_7061,N_3768,N_4826);
or U7062 (N_7062,N_4798,N_2186);
nor U7063 (N_7063,N_4944,N_4181);
xor U7064 (N_7064,N_3026,N_3179);
nor U7065 (N_7065,N_170,N_2569);
nand U7066 (N_7066,N_4714,N_1267);
nand U7067 (N_7067,N_2018,N_656);
and U7068 (N_7068,N_1469,N_3032);
and U7069 (N_7069,N_2284,N_2754);
or U7070 (N_7070,N_2646,N_2931);
or U7071 (N_7071,N_3398,N_1191);
and U7072 (N_7072,N_4127,N_836);
and U7073 (N_7073,N_1791,N_299);
nor U7074 (N_7074,N_3989,N_2252);
xor U7075 (N_7075,N_3660,N_4047);
xnor U7076 (N_7076,N_3365,N_2901);
or U7077 (N_7077,N_1890,N_3506);
and U7078 (N_7078,N_3962,N_3587);
nor U7079 (N_7079,N_4083,N_1130);
xnor U7080 (N_7080,N_479,N_3529);
or U7081 (N_7081,N_3985,N_1861);
or U7082 (N_7082,N_4984,N_2997);
nand U7083 (N_7083,N_3958,N_268);
xnor U7084 (N_7084,N_4048,N_3688);
nand U7085 (N_7085,N_1038,N_4038);
nor U7086 (N_7086,N_1446,N_3002);
or U7087 (N_7087,N_880,N_952);
nor U7088 (N_7088,N_583,N_824);
and U7089 (N_7089,N_3009,N_3209);
nand U7090 (N_7090,N_3269,N_4485);
or U7091 (N_7091,N_1610,N_4093);
and U7092 (N_7092,N_1116,N_559);
nand U7093 (N_7093,N_2729,N_595);
xnor U7094 (N_7094,N_3318,N_3397);
xor U7095 (N_7095,N_888,N_579);
and U7096 (N_7096,N_1448,N_4967);
nand U7097 (N_7097,N_1255,N_979);
or U7098 (N_7098,N_2900,N_1115);
nor U7099 (N_7099,N_897,N_4242);
nor U7100 (N_7100,N_3896,N_2819);
xor U7101 (N_7101,N_335,N_886);
or U7102 (N_7102,N_860,N_3943);
nor U7103 (N_7103,N_2482,N_1494);
nand U7104 (N_7104,N_2603,N_260);
nor U7105 (N_7105,N_2955,N_3663);
xor U7106 (N_7106,N_4927,N_643);
nor U7107 (N_7107,N_2648,N_436);
or U7108 (N_7108,N_3465,N_3839);
xor U7109 (N_7109,N_196,N_2467);
or U7110 (N_7110,N_4752,N_2723);
or U7111 (N_7111,N_2718,N_2272);
nand U7112 (N_7112,N_2641,N_279);
or U7113 (N_7113,N_1221,N_450);
and U7114 (N_7114,N_3619,N_642);
or U7115 (N_7115,N_3612,N_3591);
xor U7116 (N_7116,N_1763,N_4662);
nand U7117 (N_7117,N_1134,N_4576);
nand U7118 (N_7118,N_4018,N_3304);
nor U7119 (N_7119,N_4329,N_2121);
nor U7120 (N_7120,N_4966,N_1046);
nor U7121 (N_7121,N_1896,N_3780);
and U7122 (N_7122,N_560,N_482);
nor U7123 (N_7123,N_3742,N_4976);
nand U7124 (N_7124,N_1817,N_2287);
nor U7125 (N_7125,N_1035,N_940);
and U7126 (N_7126,N_4188,N_4855);
and U7127 (N_7127,N_3593,N_4405);
or U7128 (N_7128,N_2976,N_3225);
nor U7129 (N_7129,N_4811,N_1447);
xnor U7130 (N_7130,N_3228,N_1135);
xor U7131 (N_7131,N_1122,N_3995);
or U7132 (N_7132,N_4427,N_3630);
nor U7133 (N_7133,N_4724,N_136);
nand U7134 (N_7134,N_1528,N_1941);
and U7135 (N_7135,N_1010,N_3807);
and U7136 (N_7136,N_2114,N_2928);
or U7137 (N_7137,N_4965,N_3654);
nand U7138 (N_7138,N_3981,N_433);
or U7139 (N_7139,N_4017,N_4100);
xnor U7140 (N_7140,N_506,N_1936);
nor U7141 (N_7141,N_549,N_1514);
nor U7142 (N_7142,N_3403,N_1219);
and U7143 (N_7143,N_2040,N_975);
nand U7144 (N_7144,N_6,N_2403);
nand U7145 (N_7145,N_829,N_1853);
xor U7146 (N_7146,N_1457,N_4346);
nand U7147 (N_7147,N_1615,N_2887);
and U7148 (N_7148,N_935,N_4252);
xnor U7149 (N_7149,N_1669,N_613);
xnor U7150 (N_7150,N_2364,N_3609);
xor U7151 (N_7151,N_3950,N_770);
xnor U7152 (N_7152,N_3716,N_119);
nand U7153 (N_7153,N_627,N_1306);
xnor U7154 (N_7154,N_1891,N_1779);
xor U7155 (N_7155,N_4482,N_3201);
nor U7156 (N_7156,N_4029,N_2103);
nand U7157 (N_7157,N_4080,N_3357);
nor U7158 (N_7158,N_2054,N_1226);
nor U7159 (N_7159,N_3933,N_596);
nor U7160 (N_7160,N_2395,N_4864);
xor U7161 (N_7161,N_3363,N_1729);
nand U7162 (N_7162,N_4908,N_1111);
nand U7163 (N_7163,N_4637,N_3572);
and U7164 (N_7164,N_4153,N_1842);
nand U7165 (N_7165,N_4395,N_3724);
xnor U7166 (N_7166,N_3800,N_350);
or U7167 (N_7167,N_869,N_1437);
nand U7168 (N_7168,N_3180,N_1731);
or U7169 (N_7169,N_1644,N_4249);
or U7170 (N_7170,N_2351,N_1358);
or U7171 (N_7171,N_3301,N_2080);
xnor U7172 (N_7172,N_1201,N_3815);
and U7173 (N_7173,N_4827,N_2058);
nand U7174 (N_7174,N_1421,N_1995);
or U7175 (N_7175,N_199,N_3516);
and U7176 (N_7176,N_405,N_3157);
nand U7177 (N_7177,N_2143,N_4762);
or U7178 (N_7178,N_600,N_611);
xor U7179 (N_7179,N_3668,N_2267);
xor U7180 (N_7180,N_2850,N_1049);
and U7181 (N_7181,N_4250,N_4259);
nor U7182 (N_7182,N_785,N_2651);
and U7183 (N_7183,N_4732,N_60);
and U7184 (N_7184,N_2014,N_135);
and U7185 (N_7185,N_4973,N_1323);
nor U7186 (N_7186,N_4527,N_953);
or U7187 (N_7187,N_573,N_89);
nor U7188 (N_7188,N_4408,N_144);
and U7189 (N_7189,N_2238,N_621);
and U7190 (N_7190,N_2697,N_958);
nor U7191 (N_7191,N_368,N_4472);
and U7192 (N_7192,N_499,N_4316);
or U7193 (N_7193,N_1767,N_4210);
or U7194 (N_7194,N_3108,N_2558);
xnor U7195 (N_7195,N_1523,N_3129);
or U7196 (N_7196,N_2036,N_1620);
and U7197 (N_7197,N_2132,N_2553);
or U7198 (N_7198,N_2206,N_864);
nand U7199 (N_7199,N_1825,N_858);
xnor U7200 (N_7200,N_3691,N_4488);
and U7201 (N_7201,N_563,N_2290);
xor U7202 (N_7202,N_392,N_4005);
nand U7203 (N_7203,N_3477,N_4366);
xor U7204 (N_7204,N_2614,N_1818);
nand U7205 (N_7205,N_4299,N_746);
and U7206 (N_7206,N_332,N_3618);
nor U7207 (N_7207,N_3792,N_3379);
nor U7208 (N_7208,N_38,N_1871);
or U7209 (N_7209,N_1429,N_904);
nand U7210 (N_7210,N_3753,N_2775);
nand U7211 (N_7211,N_2115,N_11);
and U7212 (N_7212,N_3987,N_1259);
nand U7213 (N_7213,N_3238,N_4179);
nand U7214 (N_7214,N_1434,N_3192);
and U7215 (N_7215,N_3100,N_3631);
nor U7216 (N_7216,N_3530,N_1969);
or U7217 (N_7217,N_1207,N_3840);
or U7218 (N_7218,N_391,N_4336);
xor U7219 (N_7219,N_1522,N_3015);
or U7220 (N_7220,N_3750,N_394);
or U7221 (N_7221,N_2423,N_2178);
xor U7222 (N_7222,N_1934,N_4820);
nor U7223 (N_7223,N_4502,N_3972);
nor U7224 (N_7224,N_4121,N_1500);
nand U7225 (N_7225,N_3416,N_4763);
nand U7226 (N_7226,N_924,N_1743);
or U7227 (N_7227,N_3372,N_198);
nor U7228 (N_7228,N_582,N_2621);
nor U7229 (N_7229,N_4500,N_3903);
or U7230 (N_7230,N_4238,N_4036);
nand U7231 (N_7231,N_457,N_3239);
and U7232 (N_7232,N_1652,N_3486);
and U7233 (N_7233,N_353,N_395);
and U7234 (N_7234,N_2212,N_4180);
and U7235 (N_7235,N_1182,N_4836);
or U7236 (N_7236,N_4337,N_4060);
xor U7237 (N_7237,N_3161,N_2418);
or U7238 (N_7238,N_3047,N_231);
nor U7239 (N_7239,N_4627,N_4926);
nand U7240 (N_7240,N_2006,N_3730);
nand U7241 (N_7241,N_4592,N_751);
and U7242 (N_7242,N_1772,N_388);
and U7243 (N_7243,N_1439,N_1231);
nor U7244 (N_7244,N_171,N_1780);
and U7245 (N_7245,N_529,N_1847);
xnor U7246 (N_7246,N_13,N_3710);
nand U7247 (N_7247,N_2949,N_1622);
xnor U7248 (N_7248,N_4815,N_4452);
nor U7249 (N_7249,N_4830,N_1612);
xnor U7250 (N_7250,N_1815,N_1291);
xnor U7251 (N_7251,N_3531,N_3222);
and U7252 (N_7252,N_3769,N_4569);
xnor U7253 (N_7253,N_2948,N_1348);
nor U7254 (N_7254,N_4021,N_912);
or U7255 (N_7255,N_2468,N_1326);
nor U7256 (N_7256,N_1843,N_4808);
nor U7257 (N_7257,N_1089,N_418);
and U7258 (N_7258,N_1976,N_544);
xnor U7259 (N_7259,N_4453,N_625);
and U7260 (N_7260,N_1547,N_843);
nand U7261 (N_7261,N_3846,N_4288);
xnor U7262 (N_7262,N_3125,N_1964);
xnor U7263 (N_7263,N_3405,N_4578);
nand U7264 (N_7264,N_4898,N_1386);
and U7265 (N_7265,N_1981,N_3790);
nand U7266 (N_7266,N_4434,N_3822);
or U7267 (N_7267,N_2995,N_2506);
xnor U7268 (N_7268,N_1209,N_4208);
or U7269 (N_7269,N_3420,N_4182);
and U7270 (N_7270,N_4904,N_477);
or U7271 (N_7271,N_475,N_3099);
nor U7272 (N_7272,N_2233,N_4801);
xor U7273 (N_7273,N_4680,N_1277);
and U7274 (N_7274,N_535,N_3827);
xnor U7275 (N_7275,N_3744,N_1411);
or U7276 (N_7276,N_2810,N_2916);
nor U7277 (N_7277,N_3237,N_1705);
nor U7278 (N_7278,N_317,N_2571);
or U7279 (N_7279,N_247,N_2958);
nand U7280 (N_7280,N_2743,N_1057);
xor U7281 (N_7281,N_347,N_4187);
and U7282 (N_7282,N_3497,N_1028);
nor U7283 (N_7283,N_3395,N_2740);
nand U7284 (N_7284,N_4309,N_1398);
and U7285 (N_7285,N_2586,N_4079);
nor U7286 (N_7286,N_4718,N_1305);
or U7287 (N_7287,N_4828,N_2817);
nor U7288 (N_7288,N_4617,N_4786);
nand U7289 (N_7289,N_2424,N_690);
and U7290 (N_7290,N_4723,N_552);
xnor U7291 (N_7291,N_4552,N_1588);
nand U7292 (N_7292,N_1836,N_4298);
or U7293 (N_7293,N_874,N_734);
nand U7294 (N_7294,N_125,N_3523);
nand U7295 (N_7295,N_753,N_2478);
nand U7296 (N_7296,N_4895,N_4918);
or U7297 (N_7297,N_3992,N_756);
xor U7298 (N_7298,N_2912,N_311);
and U7299 (N_7299,N_4688,N_4280);
xor U7300 (N_7300,N_1373,N_2562);
or U7301 (N_7301,N_2538,N_4023);
nor U7302 (N_7302,N_649,N_2570);
xnor U7303 (N_7303,N_3184,N_4851);
nand U7304 (N_7304,N_1831,N_4871);
nor U7305 (N_7305,N_4236,N_3054);
nor U7306 (N_7306,N_4750,N_1461);
and U7307 (N_7307,N_3018,N_3641);
or U7308 (N_7308,N_384,N_1785);
and U7309 (N_7309,N_983,N_4050);
xnor U7310 (N_7310,N_2419,N_2316);
xor U7311 (N_7311,N_2377,N_1079);
nor U7312 (N_7312,N_4530,N_673);
nand U7313 (N_7313,N_3493,N_2579);
nand U7314 (N_7314,N_575,N_3785);
xor U7315 (N_7315,N_589,N_2414);
xor U7316 (N_7316,N_487,N_3103);
or U7317 (N_7317,N_717,N_2156);
and U7318 (N_7318,N_3422,N_465);
xnor U7319 (N_7319,N_2783,N_3057);
nor U7320 (N_7320,N_605,N_2552);
or U7321 (N_7321,N_4092,N_3308);
nor U7322 (N_7322,N_2195,N_806);
and U7323 (N_7323,N_1078,N_1341);
nor U7324 (N_7324,N_1848,N_714);
xnor U7325 (N_7325,N_3482,N_1148);
and U7326 (N_7326,N_3693,N_2263);
nand U7327 (N_7327,N_4232,N_1355);
nand U7328 (N_7328,N_3290,N_1509);
and U7329 (N_7329,N_4394,N_1156);
and U7330 (N_7330,N_732,N_1963);
nor U7331 (N_7331,N_4906,N_2298);
and U7332 (N_7332,N_4367,N_4755);
nand U7333 (N_7333,N_2777,N_306);
nand U7334 (N_7334,N_1003,N_3352);
nor U7335 (N_7335,N_2472,N_4940);
nor U7336 (N_7336,N_2,N_3185);
nor U7337 (N_7337,N_294,N_91);
or U7338 (N_7338,N_3342,N_4237);
nand U7339 (N_7339,N_1930,N_4390);
xnor U7340 (N_7340,N_424,N_3017);
nor U7341 (N_7341,N_1492,N_1769);
xnor U7342 (N_7342,N_2837,N_3016);
nand U7343 (N_7343,N_4511,N_2318);
or U7344 (N_7344,N_4646,N_2015);
xor U7345 (N_7345,N_4797,N_2540);
or U7346 (N_7346,N_4620,N_1271);
nand U7347 (N_7347,N_2546,N_832);
nand U7348 (N_7348,N_2959,N_1491);
and U7349 (N_7349,N_1555,N_2388);
or U7350 (N_7350,N_2555,N_2809);
and U7351 (N_7351,N_2756,N_4215);
xnor U7352 (N_7352,N_4597,N_256);
xnor U7353 (N_7353,N_1139,N_3020);
and U7354 (N_7354,N_2924,N_3624);
or U7355 (N_7355,N_2505,N_4520);
or U7356 (N_7356,N_4341,N_2044);
nor U7357 (N_7357,N_2846,N_287);
and U7358 (N_7358,N_476,N_4839);
nor U7359 (N_7359,N_1574,N_2608);
xor U7360 (N_7360,N_3359,N_74);
nor U7361 (N_7361,N_1060,N_4513);
xnor U7362 (N_7362,N_618,N_2649);
or U7363 (N_7363,N_631,N_944);
xor U7364 (N_7364,N_3235,N_66);
xnor U7365 (N_7365,N_4209,N_1109);
xor U7366 (N_7366,N_305,N_1707);
or U7367 (N_7367,N_2746,N_4370);
nor U7368 (N_7368,N_4198,N_1801);
or U7369 (N_7369,N_1788,N_308);
xnor U7370 (N_7370,N_2677,N_1453);
or U7371 (N_7371,N_1558,N_1960);
xnor U7372 (N_7372,N_2965,N_693);
or U7373 (N_7373,N_1203,N_735);
xnor U7374 (N_7374,N_3436,N_3741);
nor U7375 (N_7375,N_377,N_1220);
nor U7376 (N_7376,N_137,N_3852);
nand U7377 (N_7377,N_4476,N_115);
nand U7378 (N_7378,N_4854,N_2123);
and U7379 (N_7379,N_2950,N_3063);
or U7380 (N_7380,N_955,N_2469);
xor U7381 (N_7381,N_1643,N_1129);
nand U7382 (N_7382,N_1190,N_1091);
or U7383 (N_7383,N_248,N_1153);
nor U7384 (N_7384,N_3142,N_3329);
nor U7385 (N_7385,N_3137,N_157);
or U7386 (N_7386,N_849,N_4695);
nor U7387 (N_7387,N_2148,N_2990);
nand U7388 (N_7388,N_1859,N_3390);
nor U7389 (N_7389,N_103,N_4698);
or U7390 (N_7390,N_1725,N_3931);
and U7391 (N_7391,N_1436,N_4747);
and U7392 (N_7392,N_57,N_4818);
nor U7393 (N_7393,N_2748,N_1541);
nand U7394 (N_7394,N_3280,N_2492);
xor U7395 (N_7395,N_2432,N_1959);
or U7396 (N_7396,N_2725,N_3699);
and U7397 (N_7397,N_2000,N_481);
or U7398 (N_7398,N_999,N_4785);
or U7399 (N_7399,N_3106,N_2020);
xnor U7400 (N_7400,N_2828,N_586);
and U7401 (N_7401,N_4072,N_2644);
nand U7402 (N_7402,N_1048,N_2481);
or U7403 (N_7403,N_2230,N_1654);
xnor U7404 (N_7404,N_3601,N_112);
nand U7405 (N_7405,N_4428,N_1628);
or U7406 (N_7406,N_1143,N_445);
xnor U7407 (N_7407,N_3462,N_4339);
nor U7408 (N_7408,N_4911,N_775);
nor U7409 (N_7409,N_4326,N_4411);
xor U7410 (N_7410,N_4787,N_2169);
or U7411 (N_7411,N_1400,N_1647);
nor U7412 (N_7412,N_2029,N_823);
or U7413 (N_7413,N_3967,N_587);
or U7414 (N_7414,N_3545,N_1919);
or U7415 (N_7415,N_4905,N_3547);
nand U7416 (N_7416,N_4442,N_3537);
nor U7417 (N_7417,N_1138,N_177);
nor U7418 (N_7418,N_2715,N_3076);
or U7419 (N_7419,N_1909,N_3821);
nand U7420 (N_7420,N_4696,N_431);
xor U7421 (N_7421,N_2406,N_1692);
or U7422 (N_7422,N_1171,N_1921);
nand U7423 (N_7423,N_540,N_24);
or U7424 (N_7424,N_486,N_316);
and U7425 (N_7425,N_2779,N_201);
nor U7426 (N_7426,N_4086,N_3203);
nand U7427 (N_7427,N_2883,N_1388);
or U7428 (N_7428,N_3737,N_3842);
xnor U7429 (N_7429,N_1653,N_2270);
and U7430 (N_7430,N_3720,N_1024);
nand U7431 (N_7431,N_1668,N_407);
nand U7432 (N_7432,N_4471,N_3263);
xor U7433 (N_7433,N_2830,N_509);
nand U7434 (N_7434,N_3847,N_1248);
nand U7435 (N_7435,N_4477,N_1072);
or U7436 (N_7436,N_2334,N_3445);
nand U7437 (N_7437,N_4015,N_2413);
nor U7438 (N_7438,N_3121,N_1336);
nand U7439 (N_7439,N_3757,N_3890);
xnor U7440 (N_7440,N_2422,N_3319);
nand U7441 (N_7441,N_1096,N_4065);
or U7442 (N_7442,N_4016,N_3093);
nor U7443 (N_7443,N_263,N_1822);
xor U7444 (N_7444,N_3262,N_841);
nand U7445 (N_7445,N_2192,N_2593);
nand U7446 (N_7446,N_3177,N_4638);
and U7447 (N_7447,N_4401,N_1632);
and U7448 (N_7448,N_1269,N_2008);
or U7449 (N_7449,N_2005,N_932);
xnor U7450 (N_7450,N_1677,N_4211);
or U7451 (N_7451,N_3823,N_2433);
nor U7452 (N_7452,N_2613,N_4526);
and U7453 (N_7453,N_2972,N_4796);
or U7454 (N_7454,N_4365,N_357);
or U7455 (N_7455,N_4334,N_4887);
or U7456 (N_7456,N_4535,N_3039);
and U7457 (N_7457,N_1646,N_2863);
or U7458 (N_7458,N_1886,N_1566);
and U7459 (N_7459,N_984,N_3144);
and U7460 (N_7460,N_447,N_161);
and U7461 (N_7461,N_3169,N_1435);
nand U7462 (N_7462,N_239,N_3526);
or U7463 (N_7463,N_1,N_2001);
and U7464 (N_7464,N_4866,N_671);
nand U7465 (N_7465,N_881,N_4720);
nor U7466 (N_7466,N_3921,N_1874);
xor U7467 (N_7467,N_1655,N_174);
and U7468 (N_7468,N_914,N_3832);
xnor U7469 (N_7469,N_831,N_577);
and U7470 (N_7470,N_2737,N_2548);
nand U7471 (N_7471,N_4766,N_3838);
nor U7472 (N_7472,N_1961,N_1539);
and U7473 (N_7473,N_2340,N_1488);
and U7474 (N_7474,N_2294,N_4631);
xnor U7475 (N_7475,N_585,N_1676);
and U7476 (N_7476,N_1992,N_1524);
and U7477 (N_7477,N_722,N_515);
xor U7478 (N_7478,N_1958,N_2352);
nor U7479 (N_7479,N_3997,N_909);
xnor U7480 (N_7480,N_1161,N_1144);
nor U7481 (N_7481,N_4813,N_1062);
nor U7482 (N_7482,N_1916,N_1694);
and U7483 (N_7483,N_2869,N_745);
nor U7484 (N_7484,N_1086,N_1454);
nand U7485 (N_7485,N_2937,N_4231);
or U7486 (N_7486,N_1749,N_4431);
xnor U7487 (N_7487,N_3485,N_3834);
xnor U7488 (N_7488,N_2246,N_2214);
xnor U7489 (N_7489,N_3244,N_3513);
nand U7490 (N_7490,N_3837,N_3126);
nor U7491 (N_7491,N_902,N_2880);
nand U7492 (N_7492,N_1888,N_2078);
nor U7493 (N_7493,N_562,N_2096);
nor U7494 (N_7494,N_927,N_3878);
or U7495 (N_7495,N_341,N_601);
and U7496 (N_7496,N_3073,N_2181);
or U7497 (N_7497,N_564,N_1955);
nor U7498 (N_7498,N_4455,N_3331);
nand U7499 (N_7499,N_2358,N_1938);
nor U7500 (N_7500,N_2980,N_6);
and U7501 (N_7501,N_291,N_1736);
and U7502 (N_7502,N_3759,N_1944);
nor U7503 (N_7503,N_1877,N_1439);
nor U7504 (N_7504,N_3975,N_4984);
xnor U7505 (N_7505,N_4138,N_1513);
nor U7506 (N_7506,N_893,N_552);
nand U7507 (N_7507,N_1836,N_1827);
nand U7508 (N_7508,N_2658,N_1653);
nor U7509 (N_7509,N_491,N_2250);
nor U7510 (N_7510,N_3163,N_1542);
or U7511 (N_7511,N_4573,N_1494);
nor U7512 (N_7512,N_4702,N_3321);
or U7513 (N_7513,N_2620,N_2944);
and U7514 (N_7514,N_4798,N_89);
nor U7515 (N_7515,N_4915,N_4097);
xor U7516 (N_7516,N_269,N_3432);
xnor U7517 (N_7517,N_4662,N_2490);
nor U7518 (N_7518,N_2356,N_3490);
xnor U7519 (N_7519,N_2469,N_3124);
xor U7520 (N_7520,N_3703,N_3523);
or U7521 (N_7521,N_2479,N_3977);
or U7522 (N_7522,N_228,N_1402);
or U7523 (N_7523,N_249,N_725);
nand U7524 (N_7524,N_618,N_1479);
nor U7525 (N_7525,N_1037,N_2704);
or U7526 (N_7526,N_3394,N_918);
or U7527 (N_7527,N_3710,N_2058);
and U7528 (N_7528,N_1369,N_3012);
nor U7529 (N_7529,N_2278,N_4870);
nor U7530 (N_7530,N_2888,N_1843);
nand U7531 (N_7531,N_3999,N_1678);
nand U7532 (N_7532,N_2235,N_4515);
xor U7533 (N_7533,N_2396,N_3182);
nand U7534 (N_7534,N_503,N_495);
nand U7535 (N_7535,N_2884,N_4496);
or U7536 (N_7536,N_1468,N_3974);
nand U7537 (N_7537,N_3261,N_2727);
and U7538 (N_7538,N_4393,N_1356);
and U7539 (N_7539,N_2562,N_2782);
nor U7540 (N_7540,N_1430,N_345);
nor U7541 (N_7541,N_32,N_4145);
or U7542 (N_7542,N_3896,N_719);
xnor U7543 (N_7543,N_4203,N_1941);
or U7544 (N_7544,N_3001,N_168);
nand U7545 (N_7545,N_2225,N_4764);
and U7546 (N_7546,N_2078,N_942);
xnor U7547 (N_7547,N_2153,N_1497);
xnor U7548 (N_7548,N_2301,N_2168);
or U7549 (N_7549,N_4095,N_1966);
nand U7550 (N_7550,N_3238,N_4580);
nand U7551 (N_7551,N_2978,N_3931);
and U7552 (N_7552,N_4494,N_2523);
xnor U7553 (N_7553,N_4387,N_1975);
xor U7554 (N_7554,N_1530,N_3424);
nor U7555 (N_7555,N_1428,N_3774);
nand U7556 (N_7556,N_4339,N_89);
nor U7557 (N_7557,N_1434,N_4962);
nand U7558 (N_7558,N_1871,N_858);
and U7559 (N_7559,N_3942,N_1448);
nor U7560 (N_7560,N_290,N_3029);
xnor U7561 (N_7561,N_4497,N_3605);
nand U7562 (N_7562,N_331,N_110);
nor U7563 (N_7563,N_1150,N_3799);
xnor U7564 (N_7564,N_2297,N_3576);
and U7565 (N_7565,N_782,N_2807);
nand U7566 (N_7566,N_685,N_2549);
nand U7567 (N_7567,N_3495,N_2098);
and U7568 (N_7568,N_3413,N_1110);
or U7569 (N_7569,N_4117,N_3939);
nor U7570 (N_7570,N_3806,N_3533);
nand U7571 (N_7571,N_1359,N_219);
and U7572 (N_7572,N_1572,N_3871);
nand U7573 (N_7573,N_3839,N_4363);
and U7574 (N_7574,N_1582,N_3643);
and U7575 (N_7575,N_4424,N_101);
or U7576 (N_7576,N_501,N_1918);
and U7577 (N_7577,N_1444,N_1366);
xor U7578 (N_7578,N_306,N_4943);
xor U7579 (N_7579,N_2195,N_2044);
nand U7580 (N_7580,N_1924,N_3231);
xnor U7581 (N_7581,N_2269,N_2749);
or U7582 (N_7582,N_3759,N_3960);
nand U7583 (N_7583,N_370,N_1434);
or U7584 (N_7584,N_721,N_946);
nand U7585 (N_7585,N_1342,N_3607);
and U7586 (N_7586,N_3099,N_3344);
or U7587 (N_7587,N_532,N_2530);
nor U7588 (N_7588,N_4782,N_4640);
nand U7589 (N_7589,N_462,N_389);
or U7590 (N_7590,N_3183,N_2876);
and U7591 (N_7591,N_258,N_2401);
nand U7592 (N_7592,N_578,N_3164);
xnor U7593 (N_7593,N_3428,N_3669);
nor U7594 (N_7594,N_2666,N_4905);
and U7595 (N_7595,N_3326,N_4621);
xnor U7596 (N_7596,N_4023,N_383);
nand U7597 (N_7597,N_2079,N_2395);
or U7598 (N_7598,N_283,N_363);
and U7599 (N_7599,N_4473,N_346);
nand U7600 (N_7600,N_1546,N_2651);
nand U7601 (N_7601,N_3556,N_438);
xnor U7602 (N_7602,N_1214,N_2219);
xnor U7603 (N_7603,N_78,N_4266);
and U7604 (N_7604,N_978,N_3035);
nor U7605 (N_7605,N_2734,N_292);
nor U7606 (N_7606,N_2509,N_4359);
nor U7607 (N_7607,N_1881,N_1171);
and U7608 (N_7608,N_3585,N_2463);
or U7609 (N_7609,N_2387,N_23);
or U7610 (N_7610,N_4199,N_3366);
xor U7611 (N_7611,N_264,N_4445);
or U7612 (N_7612,N_4649,N_499);
nor U7613 (N_7613,N_549,N_3116);
nand U7614 (N_7614,N_3864,N_2069);
or U7615 (N_7615,N_1319,N_148);
nor U7616 (N_7616,N_2084,N_1675);
and U7617 (N_7617,N_4423,N_3537);
nor U7618 (N_7618,N_1547,N_2949);
and U7619 (N_7619,N_441,N_2695);
nor U7620 (N_7620,N_1788,N_512);
or U7621 (N_7621,N_2539,N_3027);
nor U7622 (N_7622,N_2169,N_575);
nor U7623 (N_7623,N_491,N_1543);
nor U7624 (N_7624,N_336,N_4481);
nand U7625 (N_7625,N_2535,N_2215);
nand U7626 (N_7626,N_2167,N_2179);
and U7627 (N_7627,N_1995,N_1827);
and U7628 (N_7628,N_593,N_3334);
xnor U7629 (N_7629,N_4954,N_2570);
nand U7630 (N_7630,N_3122,N_4059);
xnor U7631 (N_7631,N_3121,N_1463);
or U7632 (N_7632,N_1999,N_1218);
and U7633 (N_7633,N_774,N_4496);
and U7634 (N_7634,N_335,N_3904);
or U7635 (N_7635,N_1030,N_2507);
and U7636 (N_7636,N_2830,N_377);
or U7637 (N_7637,N_3255,N_3978);
nor U7638 (N_7638,N_3280,N_393);
and U7639 (N_7639,N_3968,N_1325);
nor U7640 (N_7640,N_1473,N_4426);
xor U7641 (N_7641,N_350,N_159);
nand U7642 (N_7642,N_3909,N_1680);
nand U7643 (N_7643,N_216,N_2236);
xnor U7644 (N_7644,N_4477,N_1034);
nand U7645 (N_7645,N_3673,N_1612);
and U7646 (N_7646,N_1452,N_925);
xnor U7647 (N_7647,N_3494,N_950);
nor U7648 (N_7648,N_1461,N_3772);
xnor U7649 (N_7649,N_152,N_4341);
nand U7650 (N_7650,N_1873,N_2305);
nor U7651 (N_7651,N_3996,N_1273);
or U7652 (N_7652,N_4759,N_4058);
nand U7653 (N_7653,N_1674,N_3321);
or U7654 (N_7654,N_3889,N_2156);
nand U7655 (N_7655,N_1082,N_4339);
or U7656 (N_7656,N_998,N_2959);
nor U7657 (N_7657,N_99,N_2120);
nand U7658 (N_7658,N_3369,N_4078);
xor U7659 (N_7659,N_1569,N_3427);
xor U7660 (N_7660,N_334,N_2869);
and U7661 (N_7661,N_1543,N_250);
nand U7662 (N_7662,N_2252,N_1873);
nor U7663 (N_7663,N_3348,N_3856);
and U7664 (N_7664,N_3536,N_2571);
xor U7665 (N_7665,N_4593,N_3256);
nor U7666 (N_7666,N_4487,N_275);
and U7667 (N_7667,N_4219,N_835);
or U7668 (N_7668,N_811,N_427);
xor U7669 (N_7669,N_2572,N_3410);
nand U7670 (N_7670,N_854,N_4754);
nand U7671 (N_7671,N_1648,N_4821);
nor U7672 (N_7672,N_933,N_4879);
or U7673 (N_7673,N_2781,N_4131);
and U7674 (N_7674,N_586,N_3599);
and U7675 (N_7675,N_3127,N_4632);
xnor U7676 (N_7676,N_4783,N_1292);
and U7677 (N_7677,N_3378,N_3618);
or U7678 (N_7678,N_1736,N_636);
nand U7679 (N_7679,N_1435,N_2094);
or U7680 (N_7680,N_4418,N_756);
nor U7681 (N_7681,N_4812,N_3924);
or U7682 (N_7682,N_188,N_3030);
or U7683 (N_7683,N_3035,N_773);
nand U7684 (N_7684,N_1902,N_3309);
or U7685 (N_7685,N_4283,N_1385);
and U7686 (N_7686,N_4424,N_2376);
or U7687 (N_7687,N_4349,N_2001);
nand U7688 (N_7688,N_1103,N_3168);
nor U7689 (N_7689,N_1170,N_1345);
or U7690 (N_7690,N_4538,N_2286);
nor U7691 (N_7691,N_4601,N_2203);
nand U7692 (N_7692,N_4001,N_67);
and U7693 (N_7693,N_555,N_2430);
or U7694 (N_7694,N_812,N_790);
nor U7695 (N_7695,N_2048,N_2475);
or U7696 (N_7696,N_3335,N_2771);
nor U7697 (N_7697,N_1602,N_610);
and U7698 (N_7698,N_1788,N_1005);
nor U7699 (N_7699,N_2886,N_974);
or U7700 (N_7700,N_3909,N_877);
or U7701 (N_7701,N_3081,N_1945);
and U7702 (N_7702,N_3470,N_4425);
and U7703 (N_7703,N_3939,N_2470);
nor U7704 (N_7704,N_3053,N_2342);
or U7705 (N_7705,N_3568,N_2584);
and U7706 (N_7706,N_4800,N_975);
nor U7707 (N_7707,N_2004,N_4783);
xor U7708 (N_7708,N_1509,N_3583);
nor U7709 (N_7709,N_4453,N_1713);
nor U7710 (N_7710,N_4074,N_1059);
nor U7711 (N_7711,N_2700,N_4572);
nor U7712 (N_7712,N_3934,N_1609);
or U7713 (N_7713,N_1353,N_1512);
or U7714 (N_7714,N_3512,N_3501);
and U7715 (N_7715,N_4454,N_2254);
nand U7716 (N_7716,N_4745,N_4997);
xnor U7717 (N_7717,N_3906,N_4418);
xor U7718 (N_7718,N_4082,N_1832);
nand U7719 (N_7719,N_4408,N_1739);
nand U7720 (N_7720,N_1660,N_1250);
nand U7721 (N_7721,N_1866,N_1170);
nand U7722 (N_7722,N_2668,N_739);
and U7723 (N_7723,N_4562,N_1409);
nor U7724 (N_7724,N_1741,N_4638);
and U7725 (N_7725,N_4966,N_1541);
nand U7726 (N_7726,N_674,N_3270);
nor U7727 (N_7727,N_286,N_3708);
or U7728 (N_7728,N_1811,N_2818);
nand U7729 (N_7729,N_1917,N_363);
nand U7730 (N_7730,N_2574,N_1356);
xor U7731 (N_7731,N_2123,N_2464);
nand U7732 (N_7732,N_1959,N_2547);
and U7733 (N_7733,N_1116,N_3840);
nand U7734 (N_7734,N_4755,N_1027);
and U7735 (N_7735,N_4561,N_540);
or U7736 (N_7736,N_2261,N_4078);
or U7737 (N_7737,N_2896,N_3580);
nand U7738 (N_7738,N_4851,N_1484);
and U7739 (N_7739,N_4180,N_38);
nand U7740 (N_7740,N_4700,N_731);
nand U7741 (N_7741,N_4168,N_2447);
and U7742 (N_7742,N_3409,N_4317);
nand U7743 (N_7743,N_4846,N_113);
or U7744 (N_7744,N_4594,N_1135);
and U7745 (N_7745,N_4974,N_1834);
nand U7746 (N_7746,N_2676,N_1462);
and U7747 (N_7747,N_2440,N_4125);
nand U7748 (N_7748,N_2136,N_717);
nor U7749 (N_7749,N_2872,N_896);
xnor U7750 (N_7750,N_1313,N_1617);
or U7751 (N_7751,N_158,N_1981);
and U7752 (N_7752,N_535,N_1551);
or U7753 (N_7753,N_2469,N_2560);
nand U7754 (N_7754,N_4268,N_933);
or U7755 (N_7755,N_2560,N_2865);
nor U7756 (N_7756,N_4891,N_2545);
xnor U7757 (N_7757,N_433,N_735);
xnor U7758 (N_7758,N_4519,N_4339);
nand U7759 (N_7759,N_4680,N_23);
or U7760 (N_7760,N_2157,N_1095);
and U7761 (N_7761,N_3304,N_384);
nand U7762 (N_7762,N_4958,N_3034);
and U7763 (N_7763,N_2698,N_4930);
and U7764 (N_7764,N_3381,N_1971);
nand U7765 (N_7765,N_1698,N_4191);
xor U7766 (N_7766,N_2586,N_3848);
nand U7767 (N_7767,N_377,N_3148);
nand U7768 (N_7768,N_4562,N_3262);
or U7769 (N_7769,N_2253,N_775);
and U7770 (N_7770,N_1428,N_2529);
nand U7771 (N_7771,N_4306,N_2214);
nor U7772 (N_7772,N_2214,N_262);
nor U7773 (N_7773,N_1346,N_777);
nand U7774 (N_7774,N_3160,N_3325);
nor U7775 (N_7775,N_4013,N_2912);
nand U7776 (N_7776,N_1857,N_3041);
nor U7777 (N_7777,N_1456,N_2225);
xnor U7778 (N_7778,N_2345,N_3192);
xnor U7779 (N_7779,N_3719,N_4686);
nor U7780 (N_7780,N_2635,N_3731);
nand U7781 (N_7781,N_1574,N_1409);
nand U7782 (N_7782,N_243,N_1976);
nand U7783 (N_7783,N_2795,N_1252);
xnor U7784 (N_7784,N_2239,N_1549);
nand U7785 (N_7785,N_3292,N_64);
and U7786 (N_7786,N_4572,N_1721);
xor U7787 (N_7787,N_4342,N_373);
and U7788 (N_7788,N_1472,N_3387);
xnor U7789 (N_7789,N_3727,N_4337);
and U7790 (N_7790,N_292,N_2140);
nor U7791 (N_7791,N_4309,N_705);
and U7792 (N_7792,N_4317,N_4444);
xnor U7793 (N_7793,N_2411,N_1725);
and U7794 (N_7794,N_960,N_2670);
or U7795 (N_7795,N_1407,N_2213);
nand U7796 (N_7796,N_2169,N_2979);
nor U7797 (N_7797,N_4930,N_3430);
xor U7798 (N_7798,N_1040,N_4987);
and U7799 (N_7799,N_2247,N_1939);
nand U7800 (N_7800,N_2636,N_2941);
nor U7801 (N_7801,N_4376,N_3459);
nand U7802 (N_7802,N_1085,N_1158);
or U7803 (N_7803,N_317,N_2919);
and U7804 (N_7804,N_332,N_2496);
nor U7805 (N_7805,N_4386,N_4727);
nand U7806 (N_7806,N_4499,N_4583);
or U7807 (N_7807,N_4573,N_3423);
nor U7808 (N_7808,N_1046,N_318);
nor U7809 (N_7809,N_67,N_3474);
or U7810 (N_7810,N_4779,N_4550);
or U7811 (N_7811,N_1528,N_1583);
nand U7812 (N_7812,N_4828,N_1064);
or U7813 (N_7813,N_3729,N_3820);
nand U7814 (N_7814,N_700,N_3908);
nand U7815 (N_7815,N_3809,N_3637);
or U7816 (N_7816,N_408,N_1311);
xnor U7817 (N_7817,N_3039,N_2914);
nor U7818 (N_7818,N_2407,N_4949);
nand U7819 (N_7819,N_2085,N_2040);
nor U7820 (N_7820,N_3309,N_2300);
nand U7821 (N_7821,N_3948,N_4330);
or U7822 (N_7822,N_3258,N_40);
and U7823 (N_7823,N_4450,N_841);
xnor U7824 (N_7824,N_4999,N_1838);
nor U7825 (N_7825,N_2295,N_4900);
xor U7826 (N_7826,N_2176,N_3645);
xnor U7827 (N_7827,N_2388,N_2914);
nand U7828 (N_7828,N_3120,N_3577);
or U7829 (N_7829,N_4363,N_3741);
nand U7830 (N_7830,N_337,N_3481);
or U7831 (N_7831,N_3183,N_3087);
and U7832 (N_7832,N_4326,N_1544);
nand U7833 (N_7833,N_4931,N_3612);
nand U7834 (N_7834,N_4808,N_2778);
nand U7835 (N_7835,N_1210,N_759);
or U7836 (N_7836,N_3249,N_9);
xor U7837 (N_7837,N_3823,N_1434);
nand U7838 (N_7838,N_505,N_4500);
nor U7839 (N_7839,N_972,N_1796);
or U7840 (N_7840,N_3798,N_3984);
and U7841 (N_7841,N_4220,N_3641);
nor U7842 (N_7842,N_4883,N_3035);
nand U7843 (N_7843,N_1305,N_1902);
and U7844 (N_7844,N_3387,N_1755);
and U7845 (N_7845,N_4448,N_796);
and U7846 (N_7846,N_2773,N_4784);
nand U7847 (N_7847,N_4812,N_2788);
and U7848 (N_7848,N_3740,N_3831);
xnor U7849 (N_7849,N_2781,N_2752);
or U7850 (N_7850,N_2955,N_1018);
and U7851 (N_7851,N_2506,N_3012);
xnor U7852 (N_7852,N_4415,N_2307);
nor U7853 (N_7853,N_2969,N_3944);
nor U7854 (N_7854,N_3430,N_3295);
nor U7855 (N_7855,N_695,N_1636);
and U7856 (N_7856,N_1340,N_2477);
and U7857 (N_7857,N_2785,N_1947);
nor U7858 (N_7858,N_1767,N_637);
and U7859 (N_7859,N_3074,N_475);
nor U7860 (N_7860,N_3268,N_4315);
and U7861 (N_7861,N_2830,N_2258);
and U7862 (N_7862,N_341,N_212);
xor U7863 (N_7863,N_1550,N_3940);
or U7864 (N_7864,N_3476,N_1511);
or U7865 (N_7865,N_978,N_173);
and U7866 (N_7866,N_988,N_2000);
or U7867 (N_7867,N_2976,N_4055);
and U7868 (N_7868,N_4779,N_3871);
nor U7869 (N_7869,N_2927,N_2367);
and U7870 (N_7870,N_2893,N_1811);
and U7871 (N_7871,N_1833,N_625);
or U7872 (N_7872,N_4960,N_292);
and U7873 (N_7873,N_1695,N_4080);
xor U7874 (N_7874,N_189,N_1363);
xor U7875 (N_7875,N_3410,N_2422);
nor U7876 (N_7876,N_2925,N_4122);
nor U7877 (N_7877,N_326,N_4085);
nand U7878 (N_7878,N_4413,N_3043);
nor U7879 (N_7879,N_3422,N_537);
nor U7880 (N_7880,N_1681,N_341);
xor U7881 (N_7881,N_2589,N_556);
xor U7882 (N_7882,N_3840,N_4291);
nor U7883 (N_7883,N_3931,N_1032);
or U7884 (N_7884,N_107,N_1875);
or U7885 (N_7885,N_4465,N_51);
nand U7886 (N_7886,N_145,N_195);
nor U7887 (N_7887,N_1895,N_2102);
nand U7888 (N_7888,N_22,N_88);
xor U7889 (N_7889,N_171,N_782);
nand U7890 (N_7890,N_3909,N_1253);
nand U7891 (N_7891,N_3347,N_729);
nand U7892 (N_7892,N_4675,N_4978);
xor U7893 (N_7893,N_1756,N_1640);
xnor U7894 (N_7894,N_690,N_1393);
and U7895 (N_7895,N_4442,N_954);
nor U7896 (N_7896,N_371,N_10);
or U7897 (N_7897,N_3352,N_1130);
nand U7898 (N_7898,N_2102,N_1962);
or U7899 (N_7899,N_960,N_276);
nor U7900 (N_7900,N_4930,N_4437);
and U7901 (N_7901,N_2453,N_516);
and U7902 (N_7902,N_1128,N_3056);
nand U7903 (N_7903,N_23,N_1345);
nand U7904 (N_7904,N_2759,N_2318);
xor U7905 (N_7905,N_3354,N_556);
nor U7906 (N_7906,N_4208,N_4226);
and U7907 (N_7907,N_4181,N_2753);
nand U7908 (N_7908,N_3001,N_2385);
xor U7909 (N_7909,N_3876,N_2746);
xnor U7910 (N_7910,N_922,N_4861);
nand U7911 (N_7911,N_4029,N_4397);
xor U7912 (N_7912,N_1678,N_2353);
nor U7913 (N_7913,N_4244,N_2877);
nor U7914 (N_7914,N_1112,N_4399);
nor U7915 (N_7915,N_979,N_2726);
nand U7916 (N_7916,N_2881,N_3570);
nor U7917 (N_7917,N_3968,N_1195);
nand U7918 (N_7918,N_1197,N_255);
nor U7919 (N_7919,N_4984,N_1911);
nor U7920 (N_7920,N_4820,N_4769);
nand U7921 (N_7921,N_4406,N_2851);
or U7922 (N_7922,N_703,N_211);
or U7923 (N_7923,N_1104,N_602);
and U7924 (N_7924,N_4264,N_4768);
or U7925 (N_7925,N_1337,N_1807);
and U7926 (N_7926,N_2008,N_4746);
or U7927 (N_7927,N_3795,N_4811);
or U7928 (N_7928,N_1827,N_1307);
and U7929 (N_7929,N_3161,N_3019);
xor U7930 (N_7930,N_185,N_3109);
nor U7931 (N_7931,N_1014,N_1355);
nor U7932 (N_7932,N_2766,N_4590);
or U7933 (N_7933,N_1294,N_2288);
nor U7934 (N_7934,N_3731,N_2969);
nand U7935 (N_7935,N_2979,N_35);
or U7936 (N_7936,N_4894,N_1317);
xor U7937 (N_7937,N_4983,N_1492);
or U7938 (N_7938,N_1463,N_2203);
or U7939 (N_7939,N_3542,N_4999);
or U7940 (N_7940,N_2886,N_3222);
xnor U7941 (N_7941,N_2853,N_3180);
or U7942 (N_7942,N_710,N_896);
or U7943 (N_7943,N_3646,N_3129);
xor U7944 (N_7944,N_1706,N_1609);
nor U7945 (N_7945,N_3285,N_982);
nor U7946 (N_7946,N_1769,N_739);
or U7947 (N_7947,N_3299,N_3727);
nor U7948 (N_7948,N_4544,N_1996);
nor U7949 (N_7949,N_1791,N_1166);
or U7950 (N_7950,N_2698,N_791);
nor U7951 (N_7951,N_2483,N_1247);
and U7952 (N_7952,N_394,N_3533);
xor U7953 (N_7953,N_2959,N_1071);
or U7954 (N_7954,N_4562,N_329);
or U7955 (N_7955,N_4515,N_4167);
nand U7956 (N_7956,N_392,N_2692);
or U7957 (N_7957,N_2662,N_2339);
and U7958 (N_7958,N_22,N_2511);
nor U7959 (N_7959,N_4126,N_1134);
xor U7960 (N_7960,N_374,N_2517);
and U7961 (N_7961,N_1703,N_2383);
or U7962 (N_7962,N_3923,N_866);
nor U7963 (N_7963,N_1434,N_1161);
nor U7964 (N_7964,N_1485,N_184);
nor U7965 (N_7965,N_3520,N_1699);
nor U7966 (N_7966,N_3985,N_4726);
nand U7967 (N_7967,N_3838,N_4738);
and U7968 (N_7968,N_1503,N_2138);
nand U7969 (N_7969,N_1155,N_4428);
and U7970 (N_7970,N_2910,N_3703);
xor U7971 (N_7971,N_1905,N_2003);
and U7972 (N_7972,N_4985,N_3690);
nand U7973 (N_7973,N_3804,N_2869);
and U7974 (N_7974,N_1759,N_2132);
and U7975 (N_7975,N_1453,N_4051);
nand U7976 (N_7976,N_1698,N_4950);
nor U7977 (N_7977,N_219,N_2929);
xnor U7978 (N_7978,N_954,N_3064);
or U7979 (N_7979,N_1031,N_996);
nand U7980 (N_7980,N_627,N_1393);
or U7981 (N_7981,N_393,N_2066);
and U7982 (N_7982,N_2165,N_3504);
xnor U7983 (N_7983,N_687,N_1475);
and U7984 (N_7984,N_2472,N_184);
nand U7985 (N_7985,N_3083,N_4710);
nand U7986 (N_7986,N_153,N_4328);
nand U7987 (N_7987,N_3699,N_2878);
nand U7988 (N_7988,N_1708,N_35);
xor U7989 (N_7989,N_4628,N_4504);
nand U7990 (N_7990,N_2521,N_1996);
or U7991 (N_7991,N_1016,N_1963);
or U7992 (N_7992,N_1137,N_2388);
and U7993 (N_7993,N_1790,N_1213);
or U7994 (N_7994,N_2018,N_97);
or U7995 (N_7995,N_2664,N_1524);
or U7996 (N_7996,N_618,N_319);
and U7997 (N_7997,N_3316,N_4399);
and U7998 (N_7998,N_832,N_3963);
nand U7999 (N_7999,N_1772,N_2003);
nor U8000 (N_8000,N_4478,N_4135);
and U8001 (N_8001,N_2509,N_2046);
and U8002 (N_8002,N_724,N_330);
nor U8003 (N_8003,N_668,N_3603);
and U8004 (N_8004,N_1574,N_1726);
nand U8005 (N_8005,N_337,N_2482);
xor U8006 (N_8006,N_2763,N_4767);
nand U8007 (N_8007,N_2792,N_1987);
xor U8008 (N_8008,N_1201,N_4636);
nor U8009 (N_8009,N_2519,N_4141);
xnor U8010 (N_8010,N_460,N_4493);
xnor U8011 (N_8011,N_4767,N_2521);
and U8012 (N_8012,N_2794,N_740);
and U8013 (N_8013,N_1641,N_726);
and U8014 (N_8014,N_2886,N_3304);
and U8015 (N_8015,N_2906,N_2540);
nor U8016 (N_8016,N_1900,N_2751);
and U8017 (N_8017,N_1600,N_4446);
xor U8018 (N_8018,N_4399,N_3033);
nand U8019 (N_8019,N_4053,N_2591);
and U8020 (N_8020,N_3331,N_2108);
nand U8021 (N_8021,N_2786,N_1224);
or U8022 (N_8022,N_2627,N_2706);
xnor U8023 (N_8023,N_3119,N_2445);
nand U8024 (N_8024,N_2105,N_3541);
and U8025 (N_8025,N_4362,N_1659);
xor U8026 (N_8026,N_2621,N_3682);
nor U8027 (N_8027,N_2947,N_1487);
and U8028 (N_8028,N_857,N_577);
xnor U8029 (N_8029,N_869,N_1285);
nor U8030 (N_8030,N_2637,N_4252);
and U8031 (N_8031,N_1003,N_3107);
or U8032 (N_8032,N_4748,N_1617);
nand U8033 (N_8033,N_2381,N_2268);
xor U8034 (N_8034,N_2216,N_4933);
nor U8035 (N_8035,N_2170,N_2263);
or U8036 (N_8036,N_415,N_4970);
nor U8037 (N_8037,N_1214,N_4939);
nor U8038 (N_8038,N_521,N_1043);
or U8039 (N_8039,N_1232,N_3900);
xnor U8040 (N_8040,N_4992,N_2345);
and U8041 (N_8041,N_2260,N_819);
nand U8042 (N_8042,N_986,N_4512);
nor U8043 (N_8043,N_4719,N_1557);
nor U8044 (N_8044,N_1671,N_3925);
xor U8045 (N_8045,N_3077,N_2666);
xor U8046 (N_8046,N_3493,N_2526);
nand U8047 (N_8047,N_2797,N_4888);
or U8048 (N_8048,N_1642,N_2600);
xor U8049 (N_8049,N_4576,N_1268);
nand U8050 (N_8050,N_3485,N_2092);
xor U8051 (N_8051,N_2897,N_2627);
nor U8052 (N_8052,N_2984,N_2414);
xor U8053 (N_8053,N_1534,N_2275);
and U8054 (N_8054,N_3175,N_4909);
nor U8055 (N_8055,N_2349,N_4871);
nor U8056 (N_8056,N_2716,N_3263);
nand U8057 (N_8057,N_2821,N_4806);
and U8058 (N_8058,N_1125,N_2633);
and U8059 (N_8059,N_1761,N_673);
nand U8060 (N_8060,N_4539,N_4626);
or U8061 (N_8061,N_4714,N_4454);
or U8062 (N_8062,N_4408,N_822);
or U8063 (N_8063,N_4125,N_3930);
or U8064 (N_8064,N_2698,N_3899);
and U8065 (N_8065,N_3038,N_161);
xnor U8066 (N_8066,N_1895,N_2067);
or U8067 (N_8067,N_4268,N_3630);
xor U8068 (N_8068,N_4117,N_1836);
and U8069 (N_8069,N_620,N_3215);
or U8070 (N_8070,N_3034,N_556);
xnor U8071 (N_8071,N_3619,N_1078);
xor U8072 (N_8072,N_3515,N_3136);
and U8073 (N_8073,N_1229,N_4268);
nor U8074 (N_8074,N_3009,N_925);
nand U8075 (N_8075,N_3817,N_2494);
nand U8076 (N_8076,N_1328,N_1809);
and U8077 (N_8077,N_3041,N_4335);
nand U8078 (N_8078,N_1075,N_3850);
xor U8079 (N_8079,N_3608,N_4697);
nand U8080 (N_8080,N_2279,N_3859);
nor U8081 (N_8081,N_4126,N_1074);
nand U8082 (N_8082,N_4712,N_3953);
nand U8083 (N_8083,N_838,N_2648);
xor U8084 (N_8084,N_243,N_4664);
xnor U8085 (N_8085,N_4989,N_1180);
nor U8086 (N_8086,N_3262,N_4168);
xor U8087 (N_8087,N_2446,N_4700);
nor U8088 (N_8088,N_4818,N_1095);
nor U8089 (N_8089,N_1732,N_2820);
xor U8090 (N_8090,N_2810,N_2363);
nand U8091 (N_8091,N_150,N_2488);
nor U8092 (N_8092,N_573,N_994);
xnor U8093 (N_8093,N_2769,N_4341);
nor U8094 (N_8094,N_1712,N_3026);
nor U8095 (N_8095,N_277,N_4510);
xor U8096 (N_8096,N_4376,N_2035);
nand U8097 (N_8097,N_4002,N_1932);
xor U8098 (N_8098,N_1092,N_3072);
or U8099 (N_8099,N_4328,N_1159);
or U8100 (N_8100,N_3030,N_656);
nor U8101 (N_8101,N_4978,N_763);
or U8102 (N_8102,N_1744,N_4005);
nor U8103 (N_8103,N_651,N_3234);
nand U8104 (N_8104,N_175,N_2294);
nor U8105 (N_8105,N_4662,N_2741);
nand U8106 (N_8106,N_2092,N_2568);
and U8107 (N_8107,N_1859,N_4068);
nand U8108 (N_8108,N_4539,N_4419);
nor U8109 (N_8109,N_2417,N_2665);
xor U8110 (N_8110,N_1805,N_475);
nand U8111 (N_8111,N_4686,N_887);
nor U8112 (N_8112,N_937,N_580);
nor U8113 (N_8113,N_173,N_499);
nor U8114 (N_8114,N_4449,N_1467);
nand U8115 (N_8115,N_867,N_2774);
nor U8116 (N_8116,N_2734,N_4410);
nand U8117 (N_8117,N_1484,N_4879);
or U8118 (N_8118,N_679,N_2073);
nand U8119 (N_8119,N_763,N_2051);
xor U8120 (N_8120,N_535,N_3225);
and U8121 (N_8121,N_1877,N_1258);
and U8122 (N_8122,N_4976,N_1654);
nand U8123 (N_8123,N_1084,N_2232);
xor U8124 (N_8124,N_604,N_391);
nor U8125 (N_8125,N_2491,N_2609);
and U8126 (N_8126,N_1082,N_3242);
or U8127 (N_8127,N_292,N_573);
nor U8128 (N_8128,N_4533,N_1269);
and U8129 (N_8129,N_685,N_2248);
nor U8130 (N_8130,N_2340,N_675);
xnor U8131 (N_8131,N_791,N_3044);
nor U8132 (N_8132,N_349,N_1256);
xor U8133 (N_8133,N_935,N_3241);
nand U8134 (N_8134,N_4311,N_4019);
nand U8135 (N_8135,N_4701,N_1121);
nor U8136 (N_8136,N_2670,N_3416);
nor U8137 (N_8137,N_4248,N_1821);
and U8138 (N_8138,N_2239,N_4140);
xnor U8139 (N_8139,N_546,N_3768);
nor U8140 (N_8140,N_4938,N_3454);
and U8141 (N_8141,N_3658,N_4598);
and U8142 (N_8142,N_3206,N_3735);
xnor U8143 (N_8143,N_2999,N_3879);
and U8144 (N_8144,N_504,N_1591);
nor U8145 (N_8145,N_2569,N_3183);
nand U8146 (N_8146,N_2427,N_877);
and U8147 (N_8147,N_2296,N_135);
or U8148 (N_8148,N_4124,N_3171);
or U8149 (N_8149,N_1103,N_4527);
nand U8150 (N_8150,N_3503,N_3580);
or U8151 (N_8151,N_2719,N_1005);
or U8152 (N_8152,N_446,N_3737);
xnor U8153 (N_8153,N_2620,N_998);
nand U8154 (N_8154,N_2499,N_2340);
nand U8155 (N_8155,N_2599,N_2439);
and U8156 (N_8156,N_2365,N_2537);
and U8157 (N_8157,N_19,N_3016);
nand U8158 (N_8158,N_2083,N_4339);
and U8159 (N_8159,N_389,N_2645);
xnor U8160 (N_8160,N_284,N_1338);
and U8161 (N_8161,N_451,N_346);
and U8162 (N_8162,N_2999,N_3489);
or U8163 (N_8163,N_808,N_1389);
nor U8164 (N_8164,N_3124,N_2816);
and U8165 (N_8165,N_4478,N_4459);
xor U8166 (N_8166,N_2184,N_4049);
nand U8167 (N_8167,N_2228,N_3057);
nor U8168 (N_8168,N_4555,N_190);
xnor U8169 (N_8169,N_1567,N_344);
nand U8170 (N_8170,N_1679,N_1590);
or U8171 (N_8171,N_1787,N_2612);
or U8172 (N_8172,N_1215,N_3741);
nand U8173 (N_8173,N_677,N_3270);
and U8174 (N_8174,N_3712,N_1212);
and U8175 (N_8175,N_4728,N_2027);
nor U8176 (N_8176,N_3233,N_3036);
nor U8177 (N_8177,N_3406,N_1277);
or U8178 (N_8178,N_3916,N_1140);
nor U8179 (N_8179,N_3310,N_2387);
xor U8180 (N_8180,N_519,N_405);
or U8181 (N_8181,N_4350,N_4975);
and U8182 (N_8182,N_124,N_721);
nand U8183 (N_8183,N_3502,N_3406);
nand U8184 (N_8184,N_3817,N_4724);
xnor U8185 (N_8185,N_1022,N_3430);
xnor U8186 (N_8186,N_3177,N_3074);
and U8187 (N_8187,N_2710,N_3305);
and U8188 (N_8188,N_1566,N_2307);
nand U8189 (N_8189,N_1437,N_1649);
nor U8190 (N_8190,N_4304,N_3079);
nand U8191 (N_8191,N_3269,N_60);
xnor U8192 (N_8192,N_69,N_1648);
xor U8193 (N_8193,N_3562,N_4694);
nor U8194 (N_8194,N_810,N_4440);
nand U8195 (N_8195,N_1061,N_3085);
xor U8196 (N_8196,N_3167,N_4382);
nand U8197 (N_8197,N_1826,N_1980);
or U8198 (N_8198,N_2214,N_935);
nor U8199 (N_8199,N_2533,N_1019);
nor U8200 (N_8200,N_2886,N_3621);
or U8201 (N_8201,N_3224,N_85);
nand U8202 (N_8202,N_3545,N_362);
or U8203 (N_8203,N_2280,N_2745);
xor U8204 (N_8204,N_3994,N_104);
nor U8205 (N_8205,N_4600,N_3512);
nand U8206 (N_8206,N_806,N_4622);
or U8207 (N_8207,N_1052,N_3187);
nor U8208 (N_8208,N_2564,N_4703);
or U8209 (N_8209,N_485,N_2156);
nand U8210 (N_8210,N_3918,N_3894);
and U8211 (N_8211,N_518,N_2958);
or U8212 (N_8212,N_4664,N_806);
nor U8213 (N_8213,N_244,N_2755);
and U8214 (N_8214,N_1953,N_2257);
xor U8215 (N_8215,N_3303,N_3450);
nand U8216 (N_8216,N_3659,N_260);
xnor U8217 (N_8217,N_2374,N_1857);
and U8218 (N_8218,N_4995,N_4010);
nor U8219 (N_8219,N_1294,N_4222);
xnor U8220 (N_8220,N_3021,N_4289);
or U8221 (N_8221,N_4255,N_4148);
nor U8222 (N_8222,N_4370,N_1807);
and U8223 (N_8223,N_2690,N_1192);
nand U8224 (N_8224,N_2646,N_425);
nor U8225 (N_8225,N_2293,N_3332);
xor U8226 (N_8226,N_1584,N_3209);
nor U8227 (N_8227,N_3000,N_1806);
or U8228 (N_8228,N_1006,N_888);
or U8229 (N_8229,N_1297,N_4212);
nor U8230 (N_8230,N_2605,N_4924);
and U8231 (N_8231,N_4896,N_663);
nand U8232 (N_8232,N_4328,N_2583);
or U8233 (N_8233,N_4319,N_4431);
nor U8234 (N_8234,N_4404,N_81);
or U8235 (N_8235,N_2520,N_4972);
xor U8236 (N_8236,N_492,N_3164);
xor U8237 (N_8237,N_470,N_2936);
nand U8238 (N_8238,N_286,N_2648);
xor U8239 (N_8239,N_2040,N_3860);
nor U8240 (N_8240,N_1063,N_2518);
or U8241 (N_8241,N_4756,N_460);
nor U8242 (N_8242,N_3629,N_1108);
or U8243 (N_8243,N_2918,N_4666);
and U8244 (N_8244,N_287,N_928);
nor U8245 (N_8245,N_289,N_1807);
and U8246 (N_8246,N_4222,N_864);
and U8247 (N_8247,N_4538,N_3985);
nand U8248 (N_8248,N_4011,N_3897);
and U8249 (N_8249,N_4243,N_1117);
xnor U8250 (N_8250,N_784,N_531);
nor U8251 (N_8251,N_786,N_352);
and U8252 (N_8252,N_4652,N_2403);
nor U8253 (N_8253,N_2303,N_2289);
nand U8254 (N_8254,N_2554,N_4299);
nor U8255 (N_8255,N_207,N_1908);
and U8256 (N_8256,N_4323,N_547);
and U8257 (N_8257,N_3101,N_1656);
xnor U8258 (N_8258,N_1401,N_851);
nor U8259 (N_8259,N_3779,N_1164);
or U8260 (N_8260,N_90,N_3475);
and U8261 (N_8261,N_450,N_3722);
nor U8262 (N_8262,N_3946,N_933);
nor U8263 (N_8263,N_4762,N_2810);
and U8264 (N_8264,N_2883,N_2757);
xnor U8265 (N_8265,N_2064,N_3875);
or U8266 (N_8266,N_4052,N_1319);
nor U8267 (N_8267,N_1674,N_760);
nor U8268 (N_8268,N_4565,N_2618);
nand U8269 (N_8269,N_565,N_1510);
and U8270 (N_8270,N_2062,N_3734);
or U8271 (N_8271,N_1918,N_2321);
xor U8272 (N_8272,N_4636,N_687);
nor U8273 (N_8273,N_3350,N_4255);
nand U8274 (N_8274,N_555,N_3591);
nand U8275 (N_8275,N_1479,N_1721);
xor U8276 (N_8276,N_2898,N_1156);
nor U8277 (N_8277,N_2836,N_2972);
or U8278 (N_8278,N_374,N_3897);
nor U8279 (N_8279,N_2397,N_3885);
xor U8280 (N_8280,N_2264,N_1874);
or U8281 (N_8281,N_4836,N_1920);
nand U8282 (N_8282,N_1399,N_3413);
or U8283 (N_8283,N_2655,N_4208);
nor U8284 (N_8284,N_4109,N_1000);
and U8285 (N_8285,N_813,N_423);
xnor U8286 (N_8286,N_3271,N_2571);
and U8287 (N_8287,N_2254,N_2104);
xor U8288 (N_8288,N_1862,N_3348);
or U8289 (N_8289,N_3506,N_1278);
nand U8290 (N_8290,N_1917,N_1570);
xnor U8291 (N_8291,N_1216,N_4704);
or U8292 (N_8292,N_964,N_3234);
or U8293 (N_8293,N_280,N_4034);
nand U8294 (N_8294,N_3802,N_423);
and U8295 (N_8295,N_3513,N_2377);
or U8296 (N_8296,N_2456,N_1610);
and U8297 (N_8297,N_1292,N_2228);
and U8298 (N_8298,N_4507,N_4545);
and U8299 (N_8299,N_2302,N_2170);
nand U8300 (N_8300,N_323,N_4502);
or U8301 (N_8301,N_508,N_1738);
and U8302 (N_8302,N_2154,N_185);
nor U8303 (N_8303,N_2055,N_4987);
or U8304 (N_8304,N_897,N_2385);
nor U8305 (N_8305,N_2811,N_4883);
or U8306 (N_8306,N_2360,N_1803);
nor U8307 (N_8307,N_2678,N_782);
or U8308 (N_8308,N_4786,N_2355);
nor U8309 (N_8309,N_1893,N_1734);
nor U8310 (N_8310,N_701,N_3854);
xor U8311 (N_8311,N_1603,N_759);
nor U8312 (N_8312,N_2803,N_2058);
nor U8313 (N_8313,N_2301,N_4750);
nand U8314 (N_8314,N_722,N_3503);
nand U8315 (N_8315,N_4963,N_1263);
and U8316 (N_8316,N_1195,N_4788);
nand U8317 (N_8317,N_2361,N_3829);
nor U8318 (N_8318,N_2912,N_4905);
and U8319 (N_8319,N_1860,N_3803);
and U8320 (N_8320,N_1005,N_1186);
xor U8321 (N_8321,N_4613,N_4839);
nand U8322 (N_8322,N_1195,N_508);
nand U8323 (N_8323,N_399,N_3428);
and U8324 (N_8324,N_3330,N_4905);
xor U8325 (N_8325,N_2145,N_3219);
nor U8326 (N_8326,N_420,N_3052);
nand U8327 (N_8327,N_2,N_4568);
xor U8328 (N_8328,N_1586,N_4053);
nand U8329 (N_8329,N_3852,N_4904);
nand U8330 (N_8330,N_1030,N_2698);
and U8331 (N_8331,N_420,N_4070);
nand U8332 (N_8332,N_4130,N_2254);
xnor U8333 (N_8333,N_4603,N_839);
or U8334 (N_8334,N_4838,N_3285);
or U8335 (N_8335,N_348,N_268);
nor U8336 (N_8336,N_2818,N_2816);
or U8337 (N_8337,N_4529,N_3475);
nor U8338 (N_8338,N_251,N_3581);
nor U8339 (N_8339,N_3558,N_1887);
and U8340 (N_8340,N_4630,N_3769);
xor U8341 (N_8341,N_4635,N_3148);
xor U8342 (N_8342,N_4363,N_1696);
and U8343 (N_8343,N_2067,N_2856);
and U8344 (N_8344,N_3100,N_480);
and U8345 (N_8345,N_3072,N_3113);
xor U8346 (N_8346,N_4559,N_3860);
nor U8347 (N_8347,N_3192,N_478);
xor U8348 (N_8348,N_4093,N_932);
nor U8349 (N_8349,N_3222,N_1430);
nand U8350 (N_8350,N_3798,N_1511);
or U8351 (N_8351,N_973,N_3785);
xor U8352 (N_8352,N_2942,N_3221);
and U8353 (N_8353,N_1887,N_2375);
or U8354 (N_8354,N_4133,N_3299);
xnor U8355 (N_8355,N_4649,N_2212);
or U8356 (N_8356,N_762,N_1931);
nand U8357 (N_8357,N_1613,N_2422);
xor U8358 (N_8358,N_4331,N_579);
nand U8359 (N_8359,N_151,N_3677);
nor U8360 (N_8360,N_1489,N_2677);
or U8361 (N_8361,N_316,N_497);
and U8362 (N_8362,N_4835,N_1056);
or U8363 (N_8363,N_1631,N_3443);
xnor U8364 (N_8364,N_4157,N_4767);
xor U8365 (N_8365,N_1333,N_46);
and U8366 (N_8366,N_3320,N_1891);
xor U8367 (N_8367,N_3347,N_1118);
and U8368 (N_8368,N_1973,N_2512);
nor U8369 (N_8369,N_4650,N_159);
nand U8370 (N_8370,N_2076,N_4927);
xnor U8371 (N_8371,N_2046,N_1293);
nor U8372 (N_8372,N_4745,N_448);
and U8373 (N_8373,N_3616,N_2831);
nor U8374 (N_8374,N_3397,N_3340);
nor U8375 (N_8375,N_991,N_1476);
and U8376 (N_8376,N_3490,N_52);
xor U8377 (N_8377,N_363,N_908);
nor U8378 (N_8378,N_637,N_4133);
or U8379 (N_8379,N_4106,N_534);
nor U8380 (N_8380,N_1017,N_3261);
nor U8381 (N_8381,N_471,N_4057);
or U8382 (N_8382,N_4929,N_1373);
or U8383 (N_8383,N_4246,N_23);
nor U8384 (N_8384,N_3616,N_280);
and U8385 (N_8385,N_4912,N_2732);
nand U8386 (N_8386,N_781,N_3145);
and U8387 (N_8387,N_3713,N_3507);
nand U8388 (N_8388,N_1746,N_1038);
or U8389 (N_8389,N_1856,N_4353);
nor U8390 (N_8390,N_4495,N_724);
or U8391 (N_8391,N_4108,N_954);
or U8392 (N_8392,N_3897,N_1248);
xnor U8393 (N_8393,N_3153,N_1476);
nor U8394 (N_8394,N_391,N_859);
or U8395 (N_8395,N_4949,N_885);
and U8396 (N_8396,N_4116,N_2774);
nor U8397 (N_8397,N_2699,N_1281);
and U8398 (N_8398,N_961,N_4591);
nor U8399 (N_8399,N_1501,N_2200);
and U8400 (N_8400,N_2939,N_4699);
nor U8401 (N_8401,N_2099,N_1066);
nor U8402 (N_8402,N_2753,N_2435);
or U8403 (N_8403,N_76,N_2244);
or U8404 (N_8404,N_3547,N_3926);
and U8405 (N_8405,N_464,N_2968);
nor U8406 (N_8406,N_3132,N_3265);
nor U8407 (N_8407,N_2829,N_3050);
or U8408 (N_8408,N_3920,N_4041);
nand U8409 (N_8409,N_2963,N_2172);
or U8410 (N_8410,N_1340,N_2155);
nand U8411 (N_8411,N_3547,N_2898);
xor U8412 (N_8412,N_2122,N_4878);
nand U8413 (N_8413,N_4254,N_3672);
nor U8414 (N_8414,N_3913,N_1689);
and U8415 (N_8415,N_1442,N_1094);
and U8416 (N_8416,N_558,N_3389);
xnor U8417 (N_8417,N_4687,N_3131);
and U8418 (N_8418,N_4921,N_4087);
xnor U8419 (N_8419,N_4435,N_3447);
nor U8420 (N_8420,N_3197,N_1257);
nand U8421 (N_8421,N_1380,N_2990);
xnor U8422 (N_8422,N_4664,N_253);
or U8423 (N_8423,N_1358,N_183);
and U8424 (N_8424,N_741,N_1708);
xnor U8425 (N_8425,N_4580,N_1596);
or U8426 (N_8426,N_4496,N_2546);
nand U8427 (N_8427,N_2156,N_4245);
nand U8428 (N_8428,N_3515,N_4025);
and U8429 (N_8429,N_4416,N_573);
nor U8430 (N_8430,N_3036,N_4712);
nor U8431 (N_8431,N_664,N_3031);
or U8432 (N_8432,N_1117,N_688);
or U8433 (N_8433,N_2951,N_2606);
nand U8434 (N_8434,N_1840,N_3835);
xnor U8435 (N_8435,N_1794,N_103);
and U8436 (N_8436,N_2638,N_3621);
nor U8437 (N_8437,N_2156,N_57);
xor U8438 (N_8438,N_4289,N_4514);
xnor U8439 (N_8439,N_4864,N_4815);
xnor U8440 (N_8440,N_2359,N_3025);
and U8441 (N_8441,N_1477,N_2553);
or U8442 (N_8442,N_1835,N_2784);
nand U8443 (N_8443,N_689,N_696);
xnor U8444 (N_8444,N_2640,N_1433);
nor U8445 (N_8445,N_4595,N_2747);
nand U8446 (N_8446,N_4698,N_4893);
nor U8447 (N_8447,N_256,N_479);
nor U8448 (N_8448,N_1834,N_450);
and U8449 (N_8449,N_2425,N_438);
xnor U8450 (N_8450,N_1335,N_4952);
and U8451 (N_8451,N_4614,N_3004);
nor U8452 (N_8452,N_1190,N_4099);
or U8453 (N_8453,N_4666,N_1901);
nor U8454 (N_8454,N_2269,N_1488);
xnor U8455 (N_8455,N_4104,N_4587);
or U8456 (N_8456,N_1538,N_4776);
or U8457 (N_8457,N_2950,N_4373);
or U8458 (N_8458,N_4523,N_2535);
nor U8459 (N_8459,N_1177,N_857);
nand U8460 (N_8460,N_3805,N_766);
and U8461 (N_8461,N_2801,N_4303);
nor U8462 (N_8462,N_1147,N_3158);
nand U8463 (N_8463,N_1142,N_4123);
and U8464 (N_8464,N_4760,N_3168);
and U8465 (N_8465,N_4666,N_1443);
nand U8466 (N_8466,N_676,N_3677);
or U8467 (N_8467,N_3586,N_4575);
or U8468 (N_8468,N_3448,N_4143);
xor U8469 (N_8469,N_1306,N_3967);
nand U8470 (N_8470,N_3749,N_352);
nand U8471 (N_8471,N_1853,N_4571);
and U8472 (N_8472,N_1916,N_4197);
nor U8473 (N_8473,N_2427,N_2061);
or U8474 (N_8474,N_1509,N_4628);
or U8475 (N_8475,N_142,N_3500);
nand U8476 (N_8476,N_2301,N_1991);
or U8477 (N_8477,N_495,N_885);
and U8478 (N_8478,N_2051,N_3919);
xor U8479 (N_8479,N_2243,N_2909);
and U8480 (N_8480,N_2882,N_3006);
and U8481 (N_8481,N_1433,N_4138);
xor U8482 (N_8482,N_2823,N_1011);
nand U8483 (N_8483,N_1484,N_4072);
nor U8484 (N_8484,N_1817,N_3908);
nor U8485 (N_8485,N_1759,N_2276);
or U8486 (N_8486,N_4030,N_2276);
xor U8487 (N_8487,N_4640,N_3896);
nor U8488 (N_8488,N_4851,N_4044);
or U8489 (N_8489,N_3610,N_3712);
nor U8490 (N_8490,N_2889,N_2713);
nor U8491 (N_8491,N_2677,N_2927);
or U8492 (N_8492,N_2682,N_53);
xor U8493 (N_8493,N_1302,N_825);
or U8494 (N_8494,N_3404,N_854);
and U8495 (N_8495,N_1125,N_2556);
and U8496 (N_8496,N_4567,N_575);
nor U8497 (N_8497,N_1984,N_2430);
and U8498 (N_8498,N_1723,N_1860);
xnor U8499 (N_8499,N_3370,N_3265);
and U8500 (N_8500,N_3943,N_2889);
nand U8501 (N_8501,N_3863,N_626);
and U8502 (N_8502,N_2830,N_4160);
nor U8503 (N_8503,N_2724,N_194);
nor U8504 (N_8504,N_1251,N_4578);
and U8505 (N_8505,N_777,N_3234);
or U8506 (N_8506,N_4208,N_846);
nand U8507 (N_8507,N_22,N_3866);
and U8508 (N_8508,N_1752,N_1579);
or U8509 (N_8509,N_539,N_755);
and U8510 (N_8510,N_1630,N_2627);
nor U8511 (N_8511,N_4611,N_2030);
xor U8512 (N_8512,N_4565,N_2766);
and U8513 (N_8513,N_4683,N_485);
nor U8514 (N_8514,N_1324,N_1659);
and U8515 (N_8515,N_1981,N_994);
nand U8516 (N_8516,N_3629,N_835);
and U8517 (N_8517,N_370,N_1246);
nor U8518 (N_8518,N_4907,N_1979);
nor U8519 (N_8519,N_541,N_1994);
nor U8520 (N_8520,N_1892,N_3973);
or U8521 (N_8521,N_2665,N_3562);
xor U8522 (N_8522,N_123,N_706);
or U8523 (N_8523,N_2111,N_439);
nand U8524 (N_8524,N_1555,N_3666);
xor U8525 (N_8525,N_394,N_2187);
or U8526 (N_8526,N_4766,N_2235);
nor U8527 (N_8527,N_3831,N_3040);
and U8528 (N_8528,N_67,N_1291);
nor U8529 (N_8529,N_3508,N_4372);
xor U8530 (N_8530,N_1290,N_4775);
nand U8531 (N_8531,N_3921,N_4377);
xnor U8532 (N_8532,N_3385,N_3098);
xnor U8533 (N_8533,N_3556,N_867);
and U8534 (N_8534,N_3084,N_2678);
or U8535 (N_8535,N_2148,N_2043);
nand U8536 (N_8536,N_4616,N_4940);
xnor U8537 (N_8537,N_3599,N_2116);
xnor U8538 (N_8538,N_2244,N_4794);
xor U8539 (N_8539,N_3000,N_4933);
and U8540 (N_8540,N_4898,N_2720);
xnor U8541 (N_8541,N_1529,N_1242);
xor U8542 (N_8542,N_1085,N_1909);
and U8543 (N_8543,N_1356,N_3344);
nand U8544 (N_8544,N_27,N_3070);
or U8545 (N_8545,N_881,N_670);
and U8546 (N_8546,N_3117,N_113);
nand U8547 (N_8547,N_1745,N_1110);
nor U8548 (N_8548,N_2084,N_4319);
xnor U8549 (N_8549,N_3128,N_1276);
nand U8550 (N_8550,N_3695,N_2825);
nor U8551 (N_8551,N_3705,N_951);
nor U8552 (N_8552,N_1377,N_2975);
and U8553 (N_8553,N_1921,N_873);
xnor U8554 (N_8554,N_2353,N_272);
nor U8555 (N_8555,N_3936,N_2463);
and U8556 (N_8556,N_4859,N_3155);
or U8557 (N_8557,N_2925,N_4913);
nor U8558 (N_8558,N_1549,N_895);
or U8559 (N_8559,N_1465,N_2469);
nand U8560 (N_8560,N_3158,N_2831);
nand U8561 (N_8561,N_1655,N_1837);
nor U8562 (N_8562,N_291,N_2752);
nor U8563 (N_8563,N_4086,N_1727);
and U8564 (N_8564,N_1926,N_2319);
nand U8565 (N_8565,N_3089,N_727);
and U8566 (N_8566,N_2634,N_3964);
nand U8567 (N_8567,N_2716,N_4870);
or U8568 (N_8568,N_539,N_3159);
nand U8569 (N_8569,N_2371,N_1664);
or U8570 (N_8570,N_4416,N_1946);
or U8571 (N_8571,N_500,N_2021);
nand U8572 (N_8572,N_3422,N_1334);
and U8573 (N_8573,N_3442,N_551);
and U8574 (N_8574,N_3032,N_3574);
or U8575 (N_8575,N_3199,N_514);
nand U8576 (N_8576,N_2857,N_4540);
nand U8577 (N_8577,N_2446,N_3720);
nor U8578 (N_8578,N_3231,N_1552);
xnor U8579 (N_8579,N_555,N_1829);
and U8580 (N_8580,N_4009,N_3538);
and U8581 (N_8581,N_2691,N_971);
and U8582 (N_8582,N_4364,N_918);
nor U8583 (N_8583,N_112,N_3226);
nor U8584 (N_8584,N_2489,N_1229);
nor U8585 (N_8585,N_4573,N_3740);
or U8586 (N_8586,N_864,N_1814);
xor U8587 (N_8587,N_4588,N_19);
or U8588 (N_8588,N_2628,N_1457);
or U8589 (N_8589,N_241,N_3675);
or U8590 (N_8590,N_2075,N_1631);
and U8591 (N_8591,N_860,N_3447);
and U8592 (N_8592,N_4509,N_4359);
or U8593 (N_8593,N_152,N_1101);
or U8594 (N_8594,N_3384,N_559);
and U8595 (N_8595,N_154,N_3127);
nand U8596 (N_8596,N_2919,N_4160);
and U8597 (N_8597,N_4587,N_1354);
xnor U8598 (N_8598,N_2494,N_3288);
nor U8599 (N_8599,N_1662,N_1117);
nand U8600 (N_8600,N_2739,N_4368);
nor U8601 (N_8601,N_3805,N_1239);
nand U8602 (N_8602,N_1853,N_1663);
nor U8603 (N_8603,N_938,N_3553);
nor U8604 (N_8604,N_117,N_1909);
or U8605 (N_8605,N_4613,N_1917);
nor U8606 (N_8606,N_2904,N_3070);
nand U8607 (N_8607,N_984,N_1718);
or U8608 (N_8608,N_3956,N_2694);
and U8609 (N_8609,N_4788,N_3924);
xor U8610 (N_8610,N_1293,N_1106);
or U8611 (N_8611,N_3219,N_170);
xor U8612 (N_8612,N_98,N_897);
nand U8613 (N_8613,N_916,N_2990);
nand U8614 (N_8614,N_454,N_3100);
or U8615 (N_8615,N_113,N_26);
and U8616 (N_8616,N_705,N_436);
xor U8617 (N_8617,N_215,N_3019);
nor U8618 (N_8618,N_4763,N_2460);
xor U8619 (N_8619,N_3414,N_3646);
or U8620 (N_8620,N_3893,N_4876);
or U8621 (N_8621,N_838,N_2419);
nand U8622 (N_8622,N_4820,N_3384);
or U8623 (N_8623,N_1286,N_1586);
nor U8624 (N_8624,N_687,N_1288);
xnor U8625 (N_8625,N_4079,N_1077);
and U8626 (N_8626,N_440,N_624);
xnor U8627 (N_8627,N_750,N_3749);
and U8628 (N_8628,N_504,N_3170);
and U8629 (N_8629,N_4129,N_1776);
and U8630 (N_8630,N_2962,N_4317);
xnor U8631 (N_8631,N_1059,N_3042);
nand U8632 (N_8632,N_725,N_4194);
nand U8633 (N_8633,N_3533,N_3544);
nand U8634 (N_8634,N_1866,N_1515);
or U8635 (N_8635,N_4236,N_1508);
or U8636 (N_8636,N_2317,N_4974);
nand U8637 (N_8637,N_4147,N_3618);
xnor U8638 (N_8638,N_2324,N_2872);
nand U8639 (N_8639,N_2041,N_2327);
nor U8640 (N_8640,N_3948,N_98);
nor U8641 (N_8641,N_3476,N_2097);
xor U8642 (N_8642,N_1261,N_1140);
nand U8643 (N_8643,N_4824,N_4294);
nand U8644 (N_8644,N_3137,N_2239);
or U8645 (N_8645,N_2771,N_2655);
or U8646 (N_8646,N_845,N_583);
nand U8647 (N_8647,N_4086,N_2879);
and U8648 (N_8648,N_3168,N_2811);
xnor U8649 (N_8649,N_422,N_1638);
nor U8650 (N_8650,N_4377,N_2311);
or U8651 (N_8651,N_754,N_4740);
nand U8652 (N_8652,N_690,N_4127);
or U8653 (N_8653,N_3776,N_3847);
or U8654 (N_8654,N_4716,N_2833);
or U8655 (N_8655,N_4981,N_4992);
or U8656 (N_8656,N_599,N_761);
or U8657 (N_8657,N_622,N_4612);
nand U8658 (N_8658,N_4631,N_666);
or U8659 (N_8659,N_3021,N_1601);
or U8660 (N_8660,N_3107,N_2226);
nand U8661 (N_8661,N_73,N_1675);
or U8662 (N_8662,N_2645,N_683);
xnor U8663 (N_8663,N_2432,N_4102);
and U8664 (N_8664,N_1522,N_1283);
nor U8665 (N_8665,N_3046,N_3990);
xnor U8666 (N_8666,N_2338,N_3863);
or U8667 (N_8667,N_4653,N_990);
xor U8668 (N_8668,N_1861,N_1872);
or U8669 (N_8669,N_2388,N_1484);
or U8670 (N_8670,N_1260,N_3772);
nand U8671 (N_8671,N_4826,N_902);
or U8672 (N_8672,N_3070,N_4324);
xor U8673 (N_8673,N_1415,N_1823);
or U8674 (N_8674,N_2593,N_1637);
nand U8675 (N_8675,N_21,N_1662);
or U8676 (N_8676,N_752,N_794);
and U8677 (N_8677,N_3191,N_2315);
nand U8678 (N_8678,N_3222,N_2527);
nor U8679 (N_8679,N_1138,N_1756);
xnor U8680 (N_8680,N_2465,N_4229);
or U8681 (N_8681,N_4905,N_3883);
nor U8682 (N_8682,N_4789,N_4080);
and U8683 (N_8683,N_1898,N_3511);
nand U8684 (N_8684,N_4028,N_269);
and U8685 (N_8685,N_2666,N_4976);
xnor U8686 (N_8686,N_1321,N_295);
and U8687 (N_8687,N_3905,N_1113);
nor U8688 (N_8688,N_3220,N_2021);
and U8689 (N_8689,N_3832,N_728);
or U8690 (N_8690,N_2026,N_2211);
or U8691 (N_8691,N_192,N_3565);
nand U8692 (N_8692,N_2868,N_4204);
and U8693 (N_8693,N_324,N_506);
nand U8694 (N_8694,N_49,N_4073);
and U8695 (N_8695,N_2844,N_3171);
nor U8696 (N_8696,N_4769,N_1886);
nor U8697 (N_8697,N_4115,N_1231);
xor U8698 (N_8698,N_3134,N_790);
nand U8699 (N_8699,N_1212,N_2528);
and U8700 (N_8700,N_4180,N_2044);
or U8701 (N_8701,N_484,N_1489);
nor U8702 (N_8702,N_1868,N_13);
and U8703 (N_8703,N_3959,N_2774);
xnor U8704 (N_8704,N_3432,N_2078);
nand U8705 (N_8705,N_1389,N_570);
or U8706 (N_8706,N_3685,N_2206);
nor U8707 (N_8707,N_1722,N_3606);
or U8708 (N_8708,N_2025,N_1820);
and U8709 (N_8709,N_4955,N_3750);
nand U8710 (N_8710,N_2844,N_4882);
nand U8711 (N_8711,N_3682,N_1798);
nor U8712 (N_8712,N_3056,N_347);
or U8713 (N_8713,N_806,N_1552);
xnor U8714 (N_8714,N_2423,N_3338);
and U8715 (N_8715,N_966,N_3487);
and U8716 (N_8716,N_4386,N_3527);
and U8717 (N_8717,N_409,N_1997);
nor U8718 (N_8718,N_2848,N_4640);
nor U8719 (N_8719,N_4785,N_421);
or U8720 (N_8720,N_3371,N_216);
nor U8721 (N_8721,N_2307,N_3540);
and U8722 (N_8722,N_4143,N_1743);
and U8723 (N_8723,N_4691,N_4114);
and U8724 (N_8724,N_735,N_4430);
nor U8725 (N_8725,N_3761,N_192);
nor U8726 (N_8726,N_4394,N_4610);
and U8727 (N_8727,N_1131,N_1798);
xnor U8728 (N_8728,N_263,N_4140);
and U8729 (N_8729,N_2740,N_1457);
and U8730 (N_8730,N_1073,N_4576);
xor U8731 (N_8731,N_11,N_1181);
nor U8732 (N_8732,N_2558,N_2546);
and U8733 (N_8733,N_4950,N_3899);
or U8734 (N_8734,N_237,N_606);
and U8735 (N_8735,N_1225,N_920);
xor U8736 (N_8736,N_1726,N_4558);
and U8737 (N_8737,N_2887,N_2297);
xnor U8738 (N_8738,N_658,N_1376);
nand U8739 (N_8739,N_4347,N_798);
and U8740 (N_8740,N_0,N_3603);
and U8741 (N_8741,N_2938,N_4310);
or U8742 (N_8742,N_1730,N_1278);
or U8743 (N_8743,N_1864,N_3268);
nor U8744 (N_8744,N_1328,N_924);
or U8745 (N_8745,N_1708,N_1422);
and U8746 (N_8746,N_1152,N_3557);
xor U8747 (N_8747,N_4161,N_1100);
nor U8748 (N_8748,N_414,N_1722);
and U8749 (N_8749,N_2422,N_1217);
xnor U8750 (N_8750,N_1631,N_2450);
or U8751 (N_8751,N_4571,N_573);
xnor U8752 (N_8752,N_265,N_429);
nor U8753 (N_8753,N_2300,N_869);
nor U8754 (N_8754,N_3747,N_3566);
or U8755 (N_8755,N_2145,N_123);
nor U8756 (N_8756,N_954,N_3307);
or U8757 (N_8757,N_3746,N_1082);
nor U8758 (N_8758,N_537,N_456);
nand U8759 (N_8759,N_1950,N_1614);
and U8760 (N_8760,N_1664,N_1243);
xnor U8761 (N_8761,N_125,N_4290);
or U8762 (N_8762,N_1788,N_2595);
and U8763 (N_8763,N_3668,N_13);
nor U8764 (N_8764,N_1816,N_2821);
or U8765 (N_8765,N_3686,N_1820);
and U8766 (N_8766,N_1148,N_2343);
xor U8767 (N_8767,N_4500,N_2336);
xor U8768 (N_8768,N_1661,N_2444);
nor U8769 (N_8769,N_333,N_4823);
and U8770 (N_8770,N_4683,N_4108);
nor U8771 (N_8771,N_2278,N_2915);
xnor U8772 (N_8772,N_4772,N_2388);
and U8773 (N_8773,N_1986,N_1693);
and U8774 (N_8774,N_3436,N_1167);
or U8775 (N_8775,N_3061,N_4097);
or U8776 (N_8776,N_1515,N_435);
or U8777 (N_8777,N_3438,N_987);
nand U8778 (N_8778,N_3501,N_2742);
nor U8779 (N_8779,N_1942,N_1655);
xor U8780 (N_8780,N_1970,N_2923);
nand U8781 (N_8781,N_3597,N_402);
and U8782 (N_8782,N_3212,N_1630);
nor U8783 (N_8783,N_621,N_4878);
nand U8784 (N_8784,N_640,N_951);
and U8785 (N_8785,N_3389,N_2823);
xor U8786 (N_8786,N_435,N_1811);
nor U8787 (N_8787,N_4130,N_4878);
nor U8788 (N_8788,N_4953,N_4476);
nor U8789 (N_8789,N_789,N_1893);
nor U8790 (N_8790,N_3612,N_4461);
nand U8791 (N_8791,N_2804,N_1993);
nand U8792 (N_8792,N_2138,N_271);
and U8793 (N_8793,N_2390,N_4081);
nor U8794 (N_8794,N_4441,N_1120);
xnor U8795 (N_8795,N_1918,N_1748);
xnor U8796 (N_8796,N_307,N_2213);
or U8797 (N_8797,N_173,N_4375);
nand U8798 (N_8798,N_4346,N_2113);
xnor U8799 (N_8799,N_4258,N_3172);
xor U8800 (N_8800,N_533,N_1503);
or U8801 (N_8801,N_904,N_4906);
nor U8802 (N_8802,N_4935,N_626);
and U8803 (N_8803,N_3373,N_3252);
xnor U8804 (N_8804,N_375,N_3671);
nand U8805 (N_8805,N_1487,N_1378);
and U8806 (N_8806,N_2998,N_4892);
nand U8807 (N_8807,N_3238,N_484);
xor U8808 (N_8808,N_4064,N_4304);
nor U8809 (N_8809,N_2014,N_1509);
nor U8810 (N_8810,N_835,N_4657);
xnor U8811 (N_8811,N_3809,N_4234);
nor U8812 (N_8812,N_3104,N_3095);
or U8813 (N_8813,N_4419,N_4920);
xor U8814 (N_8814,N_4422,N_1800);
xor U8815 (N_8815,N_721,N_401);
or U8816 (N_8816,N_1363,N_4);
or U8817 (N_8817,N_1611,N_1085);
nand U8818 (N_8818,N_3533,N_4571);
and U8819 (N_8819,N_2878,N_830);
xnor U8820 (N_8820,N_1711,N_1832);
or U8821 (N_8821,N_2820,N_908);
nor U8822 (N_8822,N_4601,N_4511);
and U8823 (N_8823,N_3413,N_1267);
and U8824 (N_8824,N_2285,N_392);
nor U8825 (N_8825,N_3896,N_2502);
nand U8826 (N_8826,N_1691,N_705);
nand U8827 (N_8827,N_4090,N_975);
xnor U8828 (N_8828,N_898,N_4821);
and U8829 (N_8829,N_348,N_3186);
nand U8830 (N_8830,N_3913,N_4983);
xnor U8831 (N_8831,N_3822,N_4645);
or U8832 (N_8832,N_4581,N_3114);
and U8833 (N_8833,N_979,N_1549);
or U8834 (N_8834,N_1391,N_3929);
or U8835 (N_8835,N_4109,N_1686);
nand U8836 (N_8836,N_1832,N_1475);
nor U8837 (N_8837,N_2515,N_2365);
nand U8838 (N_8838,N_4549,N_324);
nor U8839 (N_8839,N_543,N_827);
xor U8840 (N_8840,N_3358,N_2403);
xor U8841 (N_8841,N_1050,N_2611);
or U8842 (N_8842,N_4778,N_2428);
and U8843 (N_8843,N_3628,N_3019);
or U8844 (N_8844,N_3075,N_4766);
nor U8845 (N_8845,N_4033,N_706);
or U8846 (N_8846,N_10,N_2296);
and U8847 (N_8847,N_4336,N_3476);
nand U8848 (N_8848,N_3213,N_4141);
xor U8849 (N_8849,N_581,N_1294);
and U8850 (N_8850,N_4173,N_2805);
nand U8851 (N_8851,N_3288,N_2979);
and U8852 (N_8852,N_3141,N_1702);
or U8853 (N_8853,N_70,N_3072);
and U8854 (N_8854,N_1965,N_228);
nor U8855 (N_8855,N_4439,N_1522);
xor U8856 (N_8856,N_1436,N_1109);
xor U8857 (N_8857,N_517,N_4614);
xor U8858 (N_8858,N_949,N_3310);
xnor U8859 (N_8859,N_3841,N_129);
xor U8860 (N_8860,N_3269,N_4470);
xor U8861 (N_8861,N_1476,N_3302);
nor U8862 (N_8862,N_2460,N_1451);
or U8863 (N_8863,N_3578,N_619);
and U8864 (N_8864,N_1115,N_1794);
nor U8865 (N_8865,N_2217,N_3851);
or U8866 (N_8866,N_1409,N_49);
and U8867 (N_8867,N_521,N_968);
or U8868 (N_8868,N_4104,N_2207);
or U8869 (N_8869,N_3135,N_439);
or U8870 (N_8870,N_3773,N_2897);
or U8871 (N_8871,N_1264,N_2491);
and U8872 (N_8872,N_3640,N_2826);
nor U8873 (N_8873,N_1394,N_2981);
or U8874 (N_8874,N_129,N_150);
or U8875 (N_8875,N_1409,N_4209);
nand U8876 (N_8876,N_4118,N_2979);
or U8877 (N_8877,N_71,N_4001);
nand U8878 (N_8878,N_4181,N_4349);
and U8879 (N_8879,N_191,N_3277);
xnor U8880 (N_8880,N_2065,N_1913);
xnor U8881 (N_8881,N_1621,N_1661);
nor U8882 (N_8882,N_2985,N_4436);
nand U8883 (N_8883,N_4441,N_1417);
xnor U8884 (N_8884,N_2371,N_3416);
or U8885 (N_8885,N_3799,N_123);
nor U8886 (N_8886,N_2,N_1822);
and U8887 (N_8887,N_1807,N_3115);
and U8888 (N_8888,N_3452,N_1053);
nor U8889 (N_8889,N_1920,N_1600);
and U8890 (N_8890,N_2660,N_548);
or U8891 (N_8891,N_1990,N_3799);
nand U8892 (N_8892,N_2719,N_1219);
nor U8893 (N_8893,N_2584,N_4991);
nand U8894 (N_8894,N_4584,N_4666);
nor U8895 (N_8895,N_1632,N_1464);
nand U8896 (N_8896,N_4505,N_3464);
xnor U8897 (N_8897,N_411,N_926);
xor U8898 (N_8898,N_1603,N_2711);
xnor U8899 (N_8899,N_4817,N_807);
xnor U8900 (N_8900,N_4924,N_3553);
and U8901 (N_8901,N_4310,N_2626);
and U8902 (N_8902,N_4715,N_988);
xnor U8903 (N_8903,N_2769,N_3612);
nand U8904 (N_8904,N_3046,N_1217);
nand U8905 (N_8905,N_2692,N_1230);
or U8906 (N_8906,N_1649,N_1898);
nor U8907 (N_8907,N_374,N_400);
nor U8908 (N_8908,N_3871,N_2389);
or U8909 (N_8909,N_2077,N_704);
nor U8910 (N_8910,N_56,N_560);
or U8911 (N_8911,N_3992,N_523);
and U8912 (N_8912,N_1491,N_1495);
xor U8913 (N_8913,N_4161,N_2560);
and U8914 (N_8914,N_2734,N_1197);
or U8915 (N_8915,N_609,N_848);
nor U8916 (N_8916,N_4410,N_1258);
xnor U8917 (N_8917,N_627,N_641);
nor U8918 (N_8918,N_4810,N_330);
nor U8919 (N_8919,N_4694,N_2468);
or U8920 (N_8920,N_3797,N_1248);
nand U8921 (N_8921,N_4642,N_3786);
nand U8922 (N_8922,N_4429,N_382);
nor U8923 (N_8923,N_3845,N_4309);
and U8924 (N_8924,N_1620,N_3878);
or U8925 (N_8925,N_1931,N_3892);
xor U8926 (N_8926,N_1069,N_3105);
nor U8927 (N_8927,N_1796,N_1348);
and U8928 (N_8928,N_2279,N_4778);
nand U8929 (N_8929,N_3345,N_3593);
nor U8930 (N_8930,N_2799,N_2574);
nand U8931 (N_8931,N_1105,N_4529);
xor U8932 (N_8932,N_3008,N_2591);
nand U8933 (N_8933,N_1442,N_3050);
nor U8934 (N_8934,N_702,N_4858);
nor U8935 (N_8935,N_2609,N_3353);
nor U8936 (N_8936,N_2693,N_2134);
and U8937 (N_8937,N_1664,N_4225);
xor U8938 (N_8938,N_3099,N_4861);
and U8939 (N_8939,N_53,N_4783);
nand U8940 (N_8940,N_1263,N_3519);
and U8941 (N_8941,N_4267,N_3209);
nor U8942 (N_8942,N_4076,N_4306);
xnor U8943 (N_8943,N_1469,N_415);
xor U8944 (N_8944,N_47,N_1997);
nor U8945 (N_8945,N_4179,N_2054);
and U8946 (N_8946,N_1909,N_3557);
and U8947 (N_8947,N_2110,N_2037);
or U8948 (N_8948,N_4158,N_4141);
nand U8949 (N_8949,N_4654,N_3027);
and U8950 (N_8950,N_3301,N_3477);
nor U8951 (N_8951,N_1668,N_4097);
xor U8952 (N_8952,N_629,N_1059);
nor U8953 (N_8953,N_2203,N_3327);
or U8954 (N_8954,N_1700,N_2579);
nor U8955 (N_8955,N_1451,N_1585);
xnor U8956 (N_8956,N_1922,N_680);
nand U8957 (N_8957,N_2512,N_4035);
nand U8958 (N_8958,N_4567,N_880);
nor U8959 (N_8959,N_3419,N_4103);
nand U8960 (N_8960,N_3318,N_2887);
nor U8961 (N_8961,N_3782,N_2134);
xnor U8962 (N_8962,N_3908,N_2197);
nor U8963 (N_8963,N_1833,N_259);
and U8964 (N_8964,N_2533,N_2095);
and U8965 (N_8965,N_304,N_2157);
nand U8966 (N_8966,N_2014,N_2144);
xor U8967 (N_8967,N_2026,N_4886);
or U8968 (N_8968,N_4922,N_4988);
and U8969 (N_8969,N_4691,N_361);
nand U8970 (N_8970,N_4114,N_4406);
or U8971 (N_8971,N_1914,N_2833);
or U8972 (N_8972,N_4741,N_13);
nand U8973 (N_8973,N_3009,N_4357);
nand U8974 (N_8974,N_3214,N_2304);
nand U8975 (N_8975,N_1052,N_2610);
or U8976 (N_8976,N_2663,N_3669);
and U8977 (N_8977,N_1783,N_2791);
xor U8978 (N_8978,N_104,N_2320);
nand U8979 (N_8979,N_907,N_2099);
nand U8980 (N_8980,N_4862,N_3291);
nor U8981 (N_8981,N_596,N_2895);
nor U8982 (N_8982,N_2878,N_4393);
xor U8983 (N_8983,N_325,N_598);
xnor U8984 (N_8984,N_2774,N_193);
nand U8985 (N_8985,N_4633,N_4086);
and U8986 (N_8986,N_4818,N_1252);
and U8987 (N_8987,N_3888,N_324);
or U8988 (N_8988,N_2974,N_90);
nor U8989 (N_8989,N_3076,N_2494);
and U8990 (N_8990,N_1360,N_1252);
xnor U8991 (N_8991,N_1734,N_3668);
xnor U8992 (N_8992,N_4225,N_1894);
xnor U8993 (N_8993,N_4024,N_4428);
and U8994 (N_8994,N_811,N_4168);
xnor U8995 (N_8995,N_71,N_2787);
nand U8996 (N_8996,N_3343,N_3467);
nand U8997 (N_8997,N_528,N_3103);
nor U8998 (N_8998,N_2829,N_1894);
and U8999 (N_8999,N_2784,N_923);
or U9000 (N_9000,N_523,N_3662);
nor U9001 (N_9001,N_1172,N_3939);
or U9002 (N_9002,N_4555,N_1366);
nor U9003 (N_9003,N_779,N_4554);
or U9004 (N_9004,N_2281,N_4003);
and U9005 (N_9005,N_4384,N_2116);
nand U9006 (N_9006,N_1094,N_1142);
nor U9007 (N_9007,N_3873,N_4373);
and U9008 (N_9008,N_599,N_295);
xor U9009 (N_9009,N_2366,N_305);
and U9010 (N_9010,N_2057,N_80);
nand U9011 (N_9011,N_4696,N_1037);
or U9012 (N_9012,N_469,N_3717);
nand U9013 (N_9013,N_4073,N_1537);
nand U9014 (N_9014,N_607,N_3661);
nor U9015 (N_9015,N_3354,N_2081);
nand U9016 (N_9016,N_2047,N_2044);
xor U9017 (N_9017,N_3162,N_378);
nand U9018 (N_9018,N_4100,N_1240);
or U9019 (N_9019,N_1178,N_3019);
and U9020 (N_9020,N_2049,N_513);
or U9021 (N_9021,N_384,N_1588);
nor U9022 (N_9022,N_2,N_4340);
or U9023 (N_9023,N_469,N_1330);
or U9024 (N_9024,N_4331,N_2482);
and U9025 (N_9025,N_281,N_4971);
and U9026 (N_9026,N_3814,N_3357);
xor U9027 (N_9027,N_1789,N_1509);
nor U9028 (N_9028,N_4215,N_3549);
nor U9029 (N_9029,N_935,N_2382);
xor U9030 (N_9030,N_149,N_2202);
nand U9031 (N_9031,N_2003,N_2122);
nor U9032 (N_9032,N_4716,N_1213);
nor U9033 (N_9033,N_1909,N_306);
or U9034 (N_9034,N_3198,N_3614);
xor U9035 (N_9035,N_4355,N_3450);
xnor U9036 (N_9036,N_1801,N_325);
nor U9037 (N_9037,N_677,N_338);
nand U9038 (N_9038,N_4419,N_2706);
xor U9039 (N_9039,N_2331,N_2128);
nand U9040 (N_9040,N_3545,N_2377);
or U9041 (N_9041,N_4556,N_4269);
xnor U9042 (N_9042,N_3086,N_3379);
and U9043 (N_9043,N_1442,N_1376);
or U9044 (N_9044,N_3682,N_4821);
or U9045 (N_9045,N_678,N_1768);
or U9046 (N_9046,N_2154,N_3096);
nor U9047 (N_9047,N_3404,N_4578);
nand U9048 (N_9048,N_4516,N_859);
nand U9049 (N_9049,N_640,N_882);
xor U9050 (N_9050,N_1721,N_852);
and U9051 (N_9051,N_2075,N_2744);
nand U9052 (N_9052,N_4466,N_773);
or U9053 (N_9053,N_922,N_4543);
or U9054 (N_9054,N_977,N_1908);
nand U9055 (N_9055,N_3280,N_1851);
xor U9056 (N_9056,N_3724,N_96);
and U9057 (N_9057,N_1386,N_2807);
or U9058 (N_9058,N_4423,N_3623);
and U9059 (N_9059,N_3841,N_3530);
xor U9060 (N_9060,N_1936,N_3674);
or U9061 (N_9061,N_368,N_2780);
nand U9062 (N_9062,N_3754,N_450);
nand U9063 (N_9063,N_1807,N_1423);
xor U9064 (N_9064,N_3467,N_4120);
and U9065 (N_9065,N_2111,N_2281);
nor U9066 (N_9066,N_1680,N_3584);
nand U9067 (N_9067,N_4965,N_447);
and U9068 (N_9068,N_1302,N_2510);
nand U9069 (N_9069,N_4705,N_1470);
xnor U9070 (N_9070,N_1814,N_1092);
and U9071 (N_9071,N_269,N_650);
xnor U9072 (N_9072,N_4366,N_2588);
xor U9073 (N_9073,N_1440,N_3153);
and U9074 (N_9074,N_4974,N_3283);
xnor U9075 (N_9075,N_2240,N_267);
nand U9076 (N_9076,N_3669,N_2564);
and U9077 (N_9077,N_3199,N_1696);
nand U9078 (N_9078,N_3928,N_1416);
nor U9079 (N_9079,N_4932,N_2283);
nand U9080 (N_9080,N_4913,N_1230);
and U9081 (N_9081,N_2044,N_3954);
nand U9082 (N_9082,N_2695,N_1429);
and U9083 (N_9083,N_2453,N_3335);
or U9084 (N_9084,N_918,N_2638);
nand U9085 (N_9085,N_899,N_4968);
xnor U9086 (N_9086,N_3437,N_335);
nor U9087 (N_9087,N_2155,N_3202);
or U9088 (N_9088,N_1327,N_4832);
nor U9089 (N_9089,N_1615,N_1619);
nand U9090 (N_9090,N_2366,N_4966);
xor U9091 (N_9091,N_2887,N_1110);
or U9092 (N_9092,N_3296,N_3197);
nor U9093 (N_9093,N_3893,N_4386);
xnor U9094 (N_9094,N_4422,N_2545);
and U9095 (N_9095,N_3241,N_4277);
nand U9096 (N_9096,N_3090,N_455);
and U9097 (N_9097,N_2531,N_698);
or U9098 (N_9098,N_1103,N_4170);
xor U9099 (N_9099,N_2915,N_2944);
or U9100 (N_9100,N_2560,N_4478);
nand U9101 (N_9101,N_2712,N_647);
or U9102 (N_9102,N_2756,N_3105);
or U9103 (N_9103,N_3575,N_2875);
or U9104 (N_9104,N_3406,N_4450);
or U9105 (N_9105,N_1747,N_1866);
or U9106 (N_9106,N_3258,N_4078);
and U9107 (N_9107,N_387,N_3171);
xnor U9108 (N_9108,N_2468,N_2679);
and U9109 (N_9109,N_2119,N_1878);
or U9110 (N_9110,N_2454,N_301);
or U9111 (N_9111,N_2547,N_3268);
and U9112 (N_9112,N_3467,N_3977);
and U9113 (N_9113,N_2957,N_2856);
nand U9114 (N_9114,N_48,N_3752);
nand U9115 (N_9115,N_2314,N_2947);
nor U9116 (N_9116,N_1401,N_3814);
xnor U9117 (N_9117,N_4063,N_1929);
or U9118 (N_9118,N_3841,N_1225);
xor U9119 (N_9119,N_2409,N_4634);
nor U9120 (N_9120,N_4167,N_4075);
nand U9121 (N_9121,N_2764,N_2944);
or U9122 (N_9122,N_4893,N_1543);
nand U9123 (N_9123,N_269,N_3351);
nor U9124 (N_9124,N_1325,N_4123);
nor U9125 (N_9125,N_2261,N_4692);
or U9126 (N_9126,N_4849,N_3711);
nand U9127 (N_9127,N_277,N_3839);
and U9128 (N_9128,N_2770,N_4749);
or U9129 (N_9129,N_3178,N_2759);
nand U9130 (N_9130,N_311,N_3186);
nand U9131 (N_9131,N_1138,N_4725);
and U9132 (N_9132,N_4635,N_4547);
nand U9133 (N_9133,N_559,N_619);
xor U9134 (N_9134,N_1299,N_4263);
or U9135 (N_9135,N_3839,N_2928);
and U9136 (N_9136,N_4492,N_3362);
nor U9137 (N_9137,N_3739,N_3187);
or U9138 (N_9138,N_205,N_2879);
nand U9139 (N_9139,N_1237,N_1571);
nor U9140 (N_9140,N_462,N_2350);
or U9141 (N_9141,N_989,N_13);
nor U9142 (N_9142,N_3929,N_469);
nor U9143 (N_9143,N_1812,N_4683);
xnor U9144 (N_9144,N_3544,N_3019);
nor U9145 (N_9145,N_1034,N_3996);
nor U9146 (N_9146,N_3504,N_142);
nor U9147 (N_9147,N_3663,N_1513);
xnor U9148 (N_9148,N_2049,N_4258);
or U9149 (N_9149,N_2777,N_3372);
nor U9150 (N_9150,N_1402,N_2368);
xor U9151 (N_9151,N_3287,N_697);
nor U9152 (N_9152,N_1325,N_4648);
and U9153 (N_9153,N_3516,N_2291);
and U9154 (N_9154,N_603,N_1022);
nor U9155 (N_9155,N_940,N_1678);
xor U9156 (N_9156,N_1875,N_580);
xnor U9157 (N_9157,N_3835,N_719);
xor U9158 (N_9158,N_2590,N_4872);
and U9159 (N_9159,N_2762,N_814);
or U9160 (N_9160,N_1566,N_1460);
nand U9161 (N_9161,N_3025,N_641);
nor U9162 (N_9162,N_1310,N_2303);
xnor U9163 (N_9163,N_1611,N_2804);
xor U9164 (N_9164,N_646,N_3238);
xor U9165 (N_9165,N_1423,N_4050);
and U9166 (N_9166,N_874,N_231);
xor U9167 (N_9167,N_3127,N_2701);
xnor U9168 (N_9168,N_3092,N_4366);
nand U9169 (N_9169,N_3482,N_3457);
and U9170 (N_9170,N_1858,N_3562);
nor U9171 (N_9171,N_2738,N_977);
nor U9172 (N_9172,N_4182,N_176);
xnor U9173 (N_9173,N_3658,N_1999);
or U9174 (N_9174,N_1400,N_1520);
nor U9175 (N_9175,N_2813,N_3065);
or U9176 (N_9176,N_1977,N_2354);
or U9177 (N_9177,N_3764,N_1304);
or U9178 (N_9178,N_184,N_1551);
and U9179 (N_9179,N_1734,N_54);
and U9180 (N_9180,N_582,N_2098);
xor U9181 (N_9181,N_2758,N_1774);
nand U9182 (N_9182,N_1127,N_1510);
nand U9183 (N_9183,N_4492,N_4465);
and U9184 (N_9184,N_4624,N_1819);
or U9185 (N_9185,N_2399,N_125);
and U9186 (N_9186,N_730,N_3903);
and U9187 (N_9187,N_3313,N_2553);
or U9188 (N_9188,N_1497,N_395);
xnor U9189 (N_9189,N_2034,N_3184);
and U9190 (N_9190,N_4044,N_1584);
and U9191 (N_9191,N_3790,N_2776);
nand U9192 (N_9192,N_1166,N_2855);
nand U9193 (N_9193,N_389,N_3039);
and U9194 (N_9194,N_3016,N_2859);
or U9195 (N_9195,N_2726,N_4146);
xor U9196 (N_9196,N_2666,N_745);
xor U9197 (N_9197,N_4208,N_3812);
nor U9198 (N_9198,N_3005,N_1341);
or U9199 (N_9199,N_2163,N_1927);
or U9200 (N_9200,N_1254,N_3658);
and U9201 (N_9201,N_4966,N_742);
and U9202 (N_9202,N_1945,N_802);
nor U9203 (N_9203,N_3935,N_1014);
nand U9204 (N_9204,N_3610,N_1656);
nor U9205 (N_9205,N_2199,N_4809);
and U9206 (N_9206,N_3730,N_1118);
xnor U9207 (N_9207,N_2621,N_4034);
xnor U9208 (N_9208,N_2562,N_4598);
or U9209 (N_9209,N_3210,N_3192);
nand U9210 (N_9210,N_513,N_3966);
nor U9211 (N_9211,N_1614,N_2755);
nor U9212 (N_9212,N_279,N_1185);
nor U9213 (N_9213,N_83,N_2694);
xnor U9214 (N_9214,N_483,N_2748);
xnor U9215 (N_9215,N_1401,N_3003);
xor U9216 (N_9216,N_2967,N_1174);
or U9217 (N_9217,N_2021,N_3221);
and U9218 (N_9218,N_2267,N_2334);
or U9219 (N_9219,N_1448,N_4004);
nand U9220 (N_9220,N_4125,N_1494);
or U9221 (N_9221,N_260,N_944);
nand U9222 (N_9222,N_3877,N_3549);
or U9223 (N_9223,N_1731,N_2781);
nand U9224 (N_9224,N_4629,N_4581);
and U9225 (N_9225,N_4536,N_2268);
nand U9226 (N_9226,N_3448,N_3937);
nor U9227 (N_9227,N_2587,N_1538);
or U9228 (N_9228,N_858,N_4028);
and U9229 (N_9229,N_2938,N_4587);
and U9230 (N_9230,N_558,N_3696);
and U9231 (N_9231,N_4900,N_2308);
nand U9232 (N_9232,N_1195,N_2336);
or U9233 (N_9233,N_2125,N_4827);
nor U9234 (N_9234,N_425,N_77);
nor U9235 (N_9235,N_1588,N_4950);
nand U9236 (N_9236,N_3890,N_3319);
xor U9237 (N_9237,N_3608,N_3272);
and U9238 (N_9238,N_4156,N_1190);
or U9239 (N_9239,N_4116,N_3333);
and U9240 (N_9240,N_2256,N_2700);
or U9241 (N_9241,N_3116,N_1333);
or U9242 (N_9242,N_555,N_4822);
nand U9243 (N_9243,N_797,N_2483);
xnor U9244 (N_9244,N_887,N_3103);
nor U9245 (N_9245,N_402,N_4060);
xnor U9246 (N_9246,N_3829,N_1543);
nand U9247 (N_9247,N_1937,N_4109);
or U9248 (N_9248,N_1014,N_1918);
xor U9249 (N_9249,N_660,N_4476);
nand U9250 (N_9250,N_560,N_895);
nor U9251 (N_9251,N_4618,N_3018);
nor U9252 (N_9252,N_3358,N_4877);
xnor U9253 (N_9253,N_607,N_3700);
and U9254 (N_9254,N_4107,N_1563);
nor U9255 (N_9255,N_3713,N_3341);
nand U9256 (N_9256,N_4412,N_794);
nor U9257 (N_9257,N_2005,N_2016);
or U9258 (N_9258,N_3640,N_3317);
nor U9259 (N_9259,N_3037,N_1294);
nand U9260 (N_9260,N_3731,N_4821);
or U9261 (N_9261,N_4133,N_3568);
or U9262 (N_9262,N_3856,N_3464);
nor U9263 (N_9263,N_1846,N_757);
nand U9264 (N_9264,N_4414,N_4815);
nand U9265 (N_9265,N_4383,N_2371);
nand U9266 (N_9266,N_828,N_4512);
xnor U9267 (N_9267,N_4893,N_1347);
and U9268 (N_9268,N_2431,N_2642);
or U9269 (N_9269,N_3917,N_894);
nor U9270 (N_9270,N_4159,N_1809);
nand U9271 (N_9271,N_871,N_109);
nor U9272 (N_9272,N_787,N_1108);
xor U9273 (N_9273,N_168,N_1512);
and U9274 (N_9274,N_4444,N_2555);
xnor U9275 (N_9275,N_1071,N_2054);
nand U9276 (N_9276,N_3873,N_2551);
nor U9277 (N_9277,N_1056,N_4262);
and U9278 (N_9278,N_3368,N_831);
and U9279 (N_9279,N_165,N_4458);
xnor U9280 (N_9280,N_2273,N_4049);
and U9281 (N_9281,N_1430,N_2624);
nor U9282 (N_9282,N_2939,N_4551);
or U9283 (N_9283,N_2630,N_1855);
nand U9284 (N_9284,N_4070,N_984);
and U9285 (N_9285,N_1535,N_424);
nor U9286 (N_9286,N_4419,N_638);
nor U9287 (N_9287,N_161,N_2136);
nor U9288 (N_9288,N_3977,N_1796);
and U9289 (N_9289,N_2057,N_1999);
xor U9290 (N_9290,N_4683,N_34);
nor U9291 (N_9291,N_4256,N_2337);
nor U9292 (N_9292,N_3036,N_3866);
nor U9293 (N_9293,N_614,N_2666);
and U9294 (N_9294,N_1593,N_497);
nor U9295 (N_9295,N_4247,N_3223);
nand U9296 (N_9296,N_600,N_3542);
and U9297 (N_9297,N_4145,N_3597);
or U9298 (N_9298,N_2142,N_1232);
nor U9299 (N_9299,N_3463,N_2462);
xnor U9300 (N_9300,N_3241,N_1059);
nor U9301 (N_9301,N_2007,N_82);
and U9302 (N_9302,N_2607,N_1007);
nand U9303 (N_9303,N_2761,N_3420);
or U9304 (N_9304,N_666,N_1686);
xnor U9305 (N_9305,N_4798,N_4464);
and U9306 (N_9306,N_1866,N_3252);
nor U9307 (N_9307,N_2187,N_3531);
nor U9308 (N_9308,N_1778,N_700);
nor U9309 (N_9309,N_996,N_1423);
and U9310 (N_9310,N_72,N_2643);
xor U9311 (N_9311,N_3186,N_3621);
or U9312 (N_9312,N_4699,N_3317);
or U9313 (N_9313,N_314,N_507);
or U9314 (N_9314,N_2114,N_1570);
nor U9315 (N_9315,N_4690,N_3653);
nand U9316 (N_9316,N_4947,N_4105);
xor U9317 (N_9317,N_3525,N_1425);
nand U9318 (N_9318,N_3659,N_4539);
nor U9319 (N_9319,N_2169,N_267);
and U9320 (N_9320,N_3808,N_4458);
or U9321 (N_9321,N_735,N_4647);
nand U9322 (N_9322,N_438,N_2294);
xnor U9323 (N_9323,N_1932,N_808);
or U9324 (N_9324,N_4011,N_3722);
nand U9325 (N_9325,N_2329,N_455);
nor U9326 (N_9326,N_3913,N_3180);
and U9327 (N_9327,N_378,N_2680);
or U9328 (N_9328,N_1031,N_560);
xnor U9329 (N_9329,N_2950,N_1577);
xor U9330 (N_9330,N_3804,N_2293);
xnor U9331 (N_9331,N_4326,N_2797);
nand U9332 (N_9332,N_706,N_2430);
or U9333 (N_9333,N_4174,N_1042);
nand U9334 (N_9334,N_1837,N_1449);
xnor U9335 (N_9335,N_3121,N_4079);
or U9336 (N_9336,N_819,N_3059);
nor U9337 (N_9337,N_2263,N_4350);
nand U9338 (N_9338,N_4816,N_4764);
or U9339 (N_9339,N_1091,N_1968);
xnor U9340 (N_9340,N_4346,N_2086);
and U9341 (N_9341,N_3875,N_4805);
nand U9342 (N_9342,N_4904,N_2804);
and U9343 (N_9343,N_3615,N_2215);
nor U9344 (N_9344,N_2354,N_172);
or U9345 (N_9345,N_2398,N_3827);
and U9346 (N_9346,N_722,N_3352);
and U9347 (N_9347,N_1945,N_1942);
xnor U9348 (N_9348,N_3187,N_2177);
or U9349 (N_9349,N_2790,N_2386);
and U9350 (N_9350,N_2767,N_2041);
xor U9351 (N_9351,N_1431,N_2238);
nand U9352 (N_9352,N_2678,N_244);
nand U9353 (N_9353,N_3526,N_2775);
nand U9354 (N_9354,N_851,N_1178);
or U9355 (N_9355,N_4606,N_1231);
or U9356 (N_9356,N_1142,N_4229);
and U9357 (N_9357,N_3120,N_45);
or U9358 (N_9358,N_3013,N_1210);
xor U9359 (N_9359,N_657,N_4020);
nor U9360 (N_9360,N_1818,N_609);
nand U9361 (N_9361,N_491,N_3985);
and U9362 (N_9362,N_1109,N_3401);
or U9363 (N_9363,N_4062,N_1265);
nand U9364 (N_9364,N_1967,N_4307);
nor U9365 (N_9365,N_2647,N_4329);
nand U9366 (N_9366,N_443,N_845);
or U9367 (N_9367,N_3124,N_1681);
and U9368 (N_9368,N_1131,N_1332);
or U9369 (N_9369,N_228,N_4150);
and U9370 (N_9370,N_435,N_3983);
nor U9371 (N_9371,N_4148,N_2694);
xor U9372 (N_9372,N_639,N_1876);
nor U9373 (N_9373,N_834,N_2760);
and U9374 (N_9374,N_1856,N_1777);
nor U9375 (N_9375,N_3590,N_116);
nor U9376 (N_9376,N_3600,N_1977);
xor U9377 (N_9377,N_4903,N_2029);
nor U9378 (N_9378,N_4265,N_436);
xor U9379 (N_9379,N_1269,N_3190);
and U9380 (N_9380,N_334,N_2207);
xor U9381 (N_9381,N_4672,N_1447);
xor U9382 (N_9382,N_3531,N_579);
xnor U9383 (N_9383,N_2987,N_1426);
or U9384 (N_9384,N_627,N_4121);
nor U9385 (N_9385,N_4340,N_4725);
and U9386 (N_9386,N_460,N_2812);
xnor U9387 (N_9387,N_3367,N_1776);
nand U9388 (N_9388,N_3715,N_4122);
nor U9389 (N_9389,N_4218,N_2479);
nand U9390 (N_9390,N_2701,N_3675);
xor U9391 (N_9391,N_574,N_4885);
nor U9392 (N_9392,N_2698,N_184);
xnor U9393 (N_9393,N_964,N_3836);
and U9394 (N_9394,N_4889,N_26);
and U9395 (N_9395,N_4895,N_1189);
or U9396 (N_9396,N_4133,N_4176);
and U9397 (N_9397,N_760,N_4210);
and U9398 (N_9398,N_4994,N_2620);
xnor U9399 (N_9399,N_2840,N_4690);
or U9400 (N_9400,N_1489,N_4753);
and U9401 (N_9401,N_4825,N_3855);
xor U9402 (N_9402,N_3143,N_3102);
nor U9403 (N_9403,N_3777,N_1267);
nand U9404 (N_9404,N_283,N_241);
xor U9405 (N_9405,N_1344,N_2004);
or U9406 (N_9406,N_2892,N_2083);
or U9407 (N_9407,N_1349,N_4905);
and U9408 (N_9408,N_3954,N_662);
xnor U9409 (N_9409,N_3776,N_1788);
nor U9410 (N_9410,N_3658,N_1410);
and U9411 (N_9411,N_3235,N_698);
and U9412 (N_9412,N_2149,N_4009);
xor U9413 (N_9413,N_3376,N_261);
xnor U9414 (N_9414,N_690,N_4522);
nor U9415 (N_9415,N_569,N_4422);
nor U9416 (N_9416,N_2190,N_1175);
and U9417 (N_9417,N_1267,N_2388);
nor U9418 (N_9418,N_1116,N_1239);
or U9419 (N_9419,N_4380,N_2598);
nor U9420 (N_9420,N_2806,N_1881);
or U9421 (N_9421,N_997,N_1103);
nand U9422 (N_9422,N_2448,N_506);
or U9423 (N_9423,N_2300,N_1117);
or U9424 (N_9424,N_380,N_4928);
and U9425 (N_9425,N_3068,N_2380);
and U9426 (N_9426,N_432,N_2061);
nor U9427 (N_9427,N_4727,N_3994);
and U9428 (N_9428,N_3631,N_2345);
xor U9429 (N_9429,N_4483,N_4892);
xor U9430 (N_9430,N_218,N_4820);
or U9431 (N_9431,N_908,N_2007);
xor U9432 (N_9432,N_1090,N_2540);
xor U9433 (N_9433,N_169,N_2872);
and U9434 (N_9434,N_947,N_3186);
or U9435 (N_9435,N_1161,N_1746);
nor U9436 (N_9436,N_3483,N_1126);
xor U9437 (N_9437,N_1568,N_258);
and U9438 (N_9438,N_3980,N_1204);
nand U9439 (N_9439,N_4376,N_4073);
xor U9440 (N_9440,N_2467,N_349);
or U9441 (N_9441,N_2482,N_4592);
xor U9442 (N_9442,N_4489,N_920);
nand U9443 (N_9443,N_631,N_2342);
xor U9444 (N_9444,N_2175,N_2865);
and U9445 (N_9445,N_2553,N_890);
or U9446 (N_9446,N_1177,N_4673);
or U9447 (N_9447,N_4122,N_4990);
and U9448 (N_9448,N_3733,N_1631);
nor U9449 (N_9449,N_4498,N_262);
xor U9450 (N_9450,N_4786,N_2553);
nand U9451 (N_9451,N_4368,N_2624);
nand U9452 (N_9452,N_2290,N_3209);
or U9453 (N_9453,N_4916,N_3965);
or U9454 (N_9454,N_2290,N_905);
xnor U9455 (N_9455,N_3873,N_353);
and U9456 (N_9456,N_2827,N_1373);
and U9457 (N_9457,N_3379,N_1726);
nor U9458 (N_9458,N_3964,N_199);
or U9459 (N_9459,N_3536,N_3234);
and U9460 (N_9460,N_1804,N_1665);
or U9461 (N_9461,N_1647,N_232);
nand U9462 (N_9462,N_3862,N_1463);
xor U9463 (N_9463,N_3906,N_451);
xnor U9464 (N_9464,N_4158,N_4128);
nor U9465 (N_9465,N_2037,N_84);
nor U9466 (N_9466,N_1684,N_111);
nand U9467 (N_9467,N_3860,N_1092);
nand U9468 (N_9468,N_1547,N_3388);
nor U9469 (N_9469,N_3691,N_143);
and U9470 (N_9470,N_2319,N_26);
or U9471 (N_9471,N_2224,N_4227);
or U9472 (N_9472,N_296,N_1048);
and U9473 (N_9473,N_2683,N_1697);
xnor U9474 (N_9474,N_2458,N_4597);
or U9475 (N_9475,N_4911,N_2933);
or U9476 (N_9476,N_2142,N_4635);
nand U9477 (N_9477,N_4482,N_4306);
xnor U9478 (N_9478,N_4973,N_4533);
and U9479 (N_9479,N_3751,N_4460);
nor U9480 (N_9480,N_3512,N_3389);
nor U9481 (N_9481,N_3319,N_3550);
nor U9482 (N_9482,N_1772,N_3852);
xor U9483 (N_9483,N_764,N_1623);
nand U9484 (N_9484,N_2921,N_3881);
or U9485 (N_9485,N_4391,N_322);
or U9486 (N_9486,N_2235,N_1872);
nor U9487 (N_9487,N_4522,N_2583);
nor U9488 (N_9488,N_299,N_4183);
xnor U9489 (N_9489,N_3517,N_4227);
xor U9490 (N_9490,N_10,N_877);
or U9491 (N_9491,N_1317,N_1628);
nor U9492 (N_9492,N_2217,N_2518);
and U9493 (N_9493,N_4711,N_3787);
or U9494 (N_9494,N_3624,N_96);
and U9495 (N_9495,N_3703,N_1449);
xnor U9496 (N_9496,N_4246,N_1027);
and U9497 (N_9497,N_4051,N_2907);
and U9498 (N_9498,N_4292,N_1831);
or U9499 (N_9499,N_3994,N_1802);
nor U9500 (N_9500,N_3719,N_2020);
or U9501 (N_9501,N_2026,N_2611);
or U9502 (N_9502,N_937,N_3192);
nor U9503 (N_9503,N_146,N_3350);
and U9504 (N_9504,N_2933,N_2902);
xor U9505 (N_9505,N_4735,N_2894);
nand U9506 (N_9506,N_1046,N_4790);
and U9507 (N_9507,N_2491,N_2928);
or U9508 (N_9508,N_2460,N_2579);
nand U9509 (N_9509,N_4787,N_4840);
or U9510 (N_9510,N_2940,N_487);
and U9511 (N_9511,N_1262,N_885);
nand U9512 (N_9512,N_135,N_2739);
nand U9513 (N_9513,N_4619,N_90);
xnor U9514 (N_9514,N_3889,N_2185);
xnor U9515 (N_9515,N_1256,N_1435);
xnor U9516 (N_9516,N_4180,N_1024);
xnor U9517 (N_9517,N_4157,N_2052);
nor U9518 (N_9518,N_1801,N_1804);
nor U9519 (N_9519,N_1843,N_1143);
nand U9520 (N_9520,N_743,N_2551);
or U9521 (N_9521,N_1936,N_4960);
xor U9522 (N_9522,N_3782,N_3594);
nand U9523 (N_9523,N_995,N_2636);
nand U9524 (N_9524,N_4699,N_3144);
nor U9525 (N_9525,N_1577,N_4481);
xor U9526 (N_9526,N_3650,N_3300);
or U9527 (N_9527,N_4864,N_4851);
nand U9528 (N_9528,N_3265,N_1537);
and U9529 (N_9529,N_2139,N_1323);
nor U9530 (N_9530,N_1611,N_1973);
xor U9531 (N_9531,N_555,N_2356);
nor U9532 (N_9532,N_2219,N_4586);
or U9533 (N_9533,N_1920,N_2534);
or U9534 (N_9534,N_57,N_862);
nand U9535 (N_9535,N_3656,N_2592);
nor U9536 (N_9536,N_489,N_2882);
nor U9537 (N_9537,N_1494,N_749);
xor U9538 (N_9538,N_4015,N_4140);
nor U9539 (N_9539,N_2284,N_4575);
and U9540 (N_9540,N_374,N_3506);
nor U9541 (N_9541,N_1909,N_1159);
nor U9542 (N_9542,N_3226,N_1299);
or U9543 (N_9543,N_2851,N_621);
and U9544 (N_9544,N_2257,N_3273);
or U9545 (N_9545,N_697,N_4349);
nor U9546 (N_9546,N_3126,N_3760);
nand U9547 (N_9547,N_2648,N_3387);
xnor U9548 (N_9548,N_3446,N_1935);
or U9549 (N_9549,N_238,N_2640);
or U9550 (N_9550,N_3231,N_3501);
and U9551 (N_9551,N_55,N_1690);
nand U9552 (N_9552,N_3159,N_3938);
nor U9553 (N_9553,N_4520,N_2807);
and U9554 (N_9554,N_954,N_4164);
nor U9555 (N_9555,N_3467,N_3834);
or U9556 (N_9556,N_997,N_1052);
xor U9557 (N_9557,N_336,N_3026);
or U9558 (N_9558,N_788,N_4302);
nand U9559 (N_9559,N_4414,N_3528);
and U9560 (N_9560,N_3846,N_228);
and U9561 (N_9561,N_1549,N_4440);
nand U9562 (N_9562,N_74,N_4191);
nand U9563 (N_9563,N_575,N_1510);
xor U9564 (N_9564,N_1122,N_4518);
nand U9565 (N_9565,N_3877,N_2160);
and U9566 (N_9566,N_279,N_874);
nand U9567 (N_9567,N_4572,N_3747);
nor U9568 (N_9568,N_4382,N_3410);
or U9569 (N_9569,N_2452,N_3624);
and U9570 (N_9570,N_3305,N_2955);
and U9571 (N_9571,N_3469,N_2064);
nand U9572 (N_9572,N_3828,N_4181);
xnor U9573 (N_9573,N_1542,N_2948);
xnor U9574 (N_9574,N_1488,N_4696);
xor U9575 (N_9575,N_216,N_4018);
xnor U9576 (N_9576,N_1519,N_3648);
nand U9577 (N_9577,N_638,N_3340);
and U9578 (N_9578,N_4071,N_176);
and U9579 (N_9579,N_4108,N_4241);
nor U9580 (N_9580,N_1805,N_2057);
and U9581 (N_9581,N_959,N_774);
nor U9582 (N_9582,N_4409,N_1923);
nand U9583 (N_9583,N_2073,N_310);
and U9584 (N_9584,N_4121,N_1006);
xnor U9585 (N_9585,N_3580,N_3498);
xnor U9586 (N_9586,N_3764,N_443);
or U9587 (N_9587,N_2030,N_2725);
and U9588 (N_9588,N_2333,N_3654);
and U9589 (N_9589,N_2116,N_4336);
xor U9590 (N_9590,N_1979,N_434);
and U9591 (N_9591,N_72,N_667);
nor U9592 (N_9592,N_2469,N_2843);
or U9593 (N_9593,N_33,N_4671);
and U9594 (N_9594,N_2970,N_955);
nand U9595 (N_9595,N_4470,N_1490);
nand U9596 (N_9596,N_4971,N_1825);
nand U9597 (N_9597,N_2357,N_4706);
nor U9598 (N_9598,N_3920,N_2725);
nor U9599 (N_9599,N_4471,N_1049);
nand U9600 (N_9600,N_1432,N_620);
xnor U9601 (N_9601,N_2366,N_3945);
xor U9602 (N_9602,N_3045,N_3086);
nor U9603 (N_9603,N_1767,N_1501);
or U9604 (N_9604,N_2346,N_4990);
or U9605 (N_9605,N_2020,N_2192);
xnor U9606 (N_9606,N_1881,N_4389);
and U9607 (N_9607,N_1971,N_1479);
nor U9608 (N_9608,N_3216,N_4968);
nand U9609 (N_9609,N_588,N_3729);
nand U9610 (N_9610,N_4579,N_260);
or U9611 (N_9611,N_2569,N_1692);
nand U9612 (N_9612,N_111,N_1737);
nor U9613 (N_9613,N_2747,N_686);
nand U9614 (N_9614,N_92,N_3392);
nor U9615 (N_9615,N_3300,N_3822);
nor U9616 (N_9616,N_4445,N_92);
xnor U9617 (N_9617,N_4808,N_1299);
nand U9618 (N_9618,N_2525,N_868);
nor U9619 (N_9619,N_2140,N_96);
or U9620 (N_9620,N_70,N_4767);
and U9621 (N_9621,N_1842,N_1658);
and U9622 (N_9622,N_2594,N_1343);
or U9623 (N_9623,N_947,N_2369);
and U9624 (N_9624,N_4499,N_797);
xnor U9625 (N_9625,N_1773,N_200);
xor U9626 (N_9626,N_1138,N_4688);
nor U9627 (N_9627,N_4944,N_161);
nor U9628 (N_9628,N_3858,N_3130);
and U9629 (N_9629,N_4153,N_2373);
xor U9630 (N_9630,N_1020,N_3198);
and U9631 (N_9631,N_2247,N_4482);
nand U9632 (N_9632,N_1124,N_708);
xnor U9633 (N_9633,N_3050,N_2381);
nor U9634 (N_9634,N_4666,N_4102);
nor U9635 (N_9635,N_1080,N_3312);
nand U9636 (N_9636,N_2500,N_2847);
nor U9637 (N_9637,N_3229,N_4205);
or U9638 (N_9638,N_700,N_2098);
or U9639 (N_9639,N_2839,N_936);
nand U9640 (N_9640,N_3318,N_3846);
nor U9641 (N_9641,N_3569,N_1311);
nand U9642 (N_9642,N_4324,N_4223);
nand U9643 (N_9643,N_2956,N_1494);
nand U9644 (N_9644,N_2498,N_2335);
xor U9645 (N_9645,N_2231,N_1523);
or U9646 (N_9646,N_243,N_480);
xor U9647 (N_9647,N_2273,N_4482);
xnor U9648 (N_9648,N_375,N_3178);
or U9649 (N_9649,N_2351,N_2171);
xnor U9650 (N_9650,N_895,N_4862);
nor U9651 (N_9651,N_3619,N_718);
nand U9652 (N_9652,N_2573,N_2978);
or U9653 (N_9653,N_292,N_4457);
xor U9654 (N_9654,N_3386,N_3728);
or U9655 (N_9655,N_2691,N_4372);
and U9656 (N_9656,N_4967,N_137);
or U9657 (N_9657,N_1800,N_692);
nor U9658 (N_9658,N_4078,N_4522);
xnor U9659 (N_9659,N_996,N_1390);
nor U9660 (N_9660,N_3862,N_3278);
nor U9661 (N_9661,N_1576,N_1425);
and U9662 (N_9662,N_512,N_2436);
and U9663 (N_9663,N_4933,N_1292);
or U9664 (N_9664,N_2989,N_2431);
nand U9665 (N_9665,N_4554,N_1386);
or U9666 (N_9666,N_2952,N_1043);
xor U9667 (N_9667,N_404,N_231);
and U9668 (N_9668,N_522,N_2154);
and U9669 (N_9669,N_4671,N_2975);
nand U9670 (N_9670,N_3019,N_2269);
xnor U9671 (N_9671,N_4877,N_3451);
or U9672 (N_9672,N_2657,N_1735);
and U9673 (N_9673,N_3077,N_1701);
nor U9674 (N_9674,N_2546,N_194);
nand U9675 (N_9675,N_4244,N_4463);
and U9676 (N_9676,N_1129,N_3062);
or U9677 (N_9677,N_297,N_261);
xor U9678 (N_9678,N_2332,N_1893);
xor U9679 (N_9679,N_4431,N_1173);
xnor U9680 (N_9680,N_2104,N_4032);
nand U9681 (N_9681,N_3049,N_3604);
nand U9682 (N_9682,N_4692,N_83);
nand U9683 (N_9683,N_3426,N_3144);
nor U9684 (N_9684,N_4982,N_4830);
xnor U9685 (N_9685,N_1992,N_3837);
nand U9686 (N_9686,N_2018,N_4758);
and U9687 (N_9687,N_814,N_938);
nand U9688 (N_9688,N_3637,N_1152);
xnor U9689 (N_9689,N_1334,N_4565);
or U9690 (N_9690,N_4763,N_3926);
or U9691 (N_9691,N_3651,N_1656);
xnor U9692 (N_9692,N_1872,N_1351);
and U9693 (N_9693,N_3466,N_690);
xnor U9694 (N_9694,N_753,N_91);
nand U9695 (N_9695,N_2510,N_1015);
and U9696 (N_9696,N_315,N_3829);
nor U9697 (N_9697,N_3619,N_95);
xor U9698 (N_9698,N_802,N_1840);
nand U9699 (N_9699,N_3476,N_3583);
xor U9700 (N_9700,N_4793,N_1223);
nor U9701 (N_9701,N_3172,N_3246);
and U9702 (N_9702,N_4119,N_3398);
nor U9703 (N_9703,N_1779,N_4221);
nand U9704 (N_9704,N_2296,N_4874);
xnor U9705 (N_9705,N_3316,N_3196);
and U9706 (N_9706,N_1569,N_1069);
and U9707 (N_9707,N_3760,N_4116);
and U9708 (N_9708,N_1661,N_4544);
nand U9709 (N_9709,N_1697,N_280);
and U9710 (N_9710,N_647,N_4642);
or U9711 (N_9711,N_604,N_3462);
nand U9712 (N_9712,N_3688,N_2117);
nor U9713 (N_9713,N_2933,N_1340);
and U9714 (N_9714,N_2758,N_1223);
nor U9715 (N_9715,N_3209,N_3711);
nor U9716 (N_9716,N_2185,N_3379);
and U9717 (N_9717,N_2021,N_3898);
nand U9718 (N_9718,N_2206,N_483);
or U9719 (N_9719,N_1721,N_261);
and U9720 (N_9720,N_2809,N_2792);
or U9721 (N_9721,N_4136,N_4167);
nor U9722 (N_9722,N_3423,N_4591);
or U9723 (N_9723,N_1075,N_3493);
nand U9724 (N_9724,N_1358,N_4542);
nor U9725 (N_9725,N_1614,N_852);
or U9726 (N_9726,N_2955,N_908);
nor U9727 (N_9727,N_109,N_1401);
nor U9728 (N_9728,N_1443,N_2689);
or U9729 (N_9729,N_2259,N_1166);
nand U9730 (N_9730,N_262,N_2097);
and U9731 (N_9731,N_936,N_4562);
nand U9732 (N_9732,N_2067,N_3735);
nand U9733 (N_9733,N_4732,N_3649);
and U9734 (N_9734,N_4846,N_4440);
nand U9735 (N_9735,N_2890,N_4563);
nand U9736 (N_9736,N_3544,N_2491);
nand U9737 (N_9737,N_2333,N_433);
nand U9738 (N_9738,N_4293,N_2136);
xnor U9739 (N_9739,N_2109,N_1544);
nor U9740 (N_9740,N_4221,N_2394);
or U9741 (N_9741,N_3468,N_915);
or U9742 (N_9742,N_2747,N_3072);
or U9743 (N_9743,N_2941,N_3231);
nor U9744 (N_9744,N_994,N_1805);
nor U9745 (N_9745,N_3774,N_4929);
nor U9746 (N_9746,N_1879,N_4157);
xor U9747 (N_9747,N_3172,N_4911);
xnor U9748 (N_9748,N_4800,N_220);
or U9749 (N_9749,N_134,N_2010);
xor U9750 (N_9750,N_2611,N_3245);
nand U9751 (N_9751,N_1560,N_1883);
nand U9752 (N_9752,N_3197,N_3017);
nor U9753 (N_9753,N_1312,N_315);
nand U9754 (N_9754,N_970,N_2898);
nor U9755 (N_9755,N_390,N_937);
nand U9756 (N_9756,N_2415,N_3469);
nor U9757 (N_9757,N_4250,N_4293);
nor U9758 (N_9758,N_2486,N_2365);
nor U9759 (N_9759,N_2556,N_2432);
nor U9760 (N_9760,N_768,N_1521);
xor U9761 (N_9761,N_4698,N_4533);
and U9762 (N_9762,N_3913,N_3638);
nand U9763 (N_9763,N_3526,N_4929);
nor U9764 (N_9764,N_2318,N_4579);
xor U9765 (N_9765,N_1594,N_849);
nor U9766 (N_9766,N_2362,N_4185);
or U9767 (N_9767,N_3074,N_3481);
and U9768 (N_9768,N_1031,N_2273);
xnor U9769 (N_9769,N_4857,N_4449);
nand U9770 (N_9770,N_3749,N_4516);
xnor U9771 (N_9771,N_1621,N_1646);
xnor U9772 (N_9772,N_4859,N_4810);
nor U9773 (N_9773,N_321,N_1376);
nand U9774 (N_9774,N_3682,N_2476);
xnor U9775 (N_9775,N_1020,N_940);
and U9776 (N_9776,N_3904,N_784);
and U9777 (N_9777,N_583,N_4812);
xor U9778 (N_9778,N_3191,N_551);
xnor U9779 (N_9779,N_3116,N_1420);
or U9780 (N_9780,N_4389,N_329);
nand U9781 (N_9781,N_1782,N_4296);
and U9782 (N_9782,N_459,N_1344);
xnor U9783 (N_9783,N_1522,N_4240);
nand U9784 (N_9784,N_2233,N_2092);
nor U9785 (N_9785,N_2066,N_4643);
xor U9786 (N_9786,N_2164,N_1618);
nand U9787 (N_9787,N_3918,N_531);
nand U9788 (N_9788,N_4830,N_2748);
or U9789 (N_9789,N_3214,N_2451);
xor U9790 (N_9790,N_1572,N_4670);
or U9791 (N_9791,N_4752,N_1099);
and U9792 (N_9792,N_892,N_478);
xor U9793 (N_9793,N_3604,N_2839);
xnor U9794 (N_9794,N_2782,N_4182);
nand U9795 (N_9795,N_2764,N_2448);
nor U9796 (N_9796,N_3946,N_3858);
nor U9797 (N_9797,N_1870,N_4985);
or U9798 (N_9798,N_3590,N_1562);
xor U9799 (N_9799,N_1300,N_2484);
nand U9800 (N_9800,N_933,N_2999);
nand U9801 (N_9801,N_1339,N_2679);
or U9802 (N_9802,N_413,N_1157);
nor U9803 (N_9803,N_4559,N_2725);
xor U9804 (N_9804,N_2681,N_1834);
and U9805 (N_9805,N_4036,N_2124);
nand U9806 (N_9806,N_1251,N_2295);
or U9807 (N_9807,N_1977,N_4654);
nand U9808 (N_9808,N_3421,N_4642);
xnor U9809 (N_9809,N_4115,N_1369);
and U9810 (N_9810,N_4796,N_579);
or U9811 (N_9811,N_1423,N_1802);
and U9812 (N_9812,N_463,N_4482);
or U9813 (N_9813,N_3764,N_3105);
nand U9814 (N_9814,N_1179,N_652);
nand U9815 (N_9815,N_811,N_2915);
xor U9816 (N_9816,N_874,N_675);
or U9817 (N_9817,N_980,N_787);
xnor U9818 (N_9818,N_4772,N_3970);
or U9819 (N_9819,N_2937,N_386);
xor U9820 (N_9820,N_2334,N_4965);
or U9821 (N_9821,N_4520,N_3969);
and U9822 (N_9822,N_4824,N_706);
and U9823 (N_9823,N_3674,N_1707);
xor U9824 (N_9824,N_2634,N_3137);
nand U9825 (N_9825,N_3472,N_328);
xor U9826 (N_9826,N_2995,N_4918);
and U9827 (N_9827,N_168,N_1949);
nand U9828 (N_9828,N_4950,N_2023);
or U9829 (N_9829,N_4872,N_2343);
and U9830 (N_9830,N_2717,N_314);
xor U9831 (N_9831,N_941,N_4385);
and U9832 (N_9832,N_4455,N_4335);
nor U9833 (N_9833,N_3862,N_1154);
nand U9834 (N_9834,N_2717,N_1344);
and U9835 (N_9835,N_2884,N_1611);
nand U9836 (N_9836,N_4469,N_1233);
nand U9837 (N_9837,N_1607,N_4304);
nor U9838 (N_9838,N_59,N_4858);
and U9839 (N_9839,N_4134,N_942);
or U9840 (N_9840,N_4472,N_4414);
nand U9841 (N_9841,N_4409,N_3337);
or U9842 (N_9842,N_2533,N_2130);
xor U9843 (N_9843,N_4808,N_1627);
nor U9844 (N_9844,N_1328,N_4699);
or U9845 (N_9845,N_2012,N_409);
or U9846 (N_9846,N_1832,N_3361);
nor U9847 (N_9847,N_371,N_1583);
and U9848 (N_9848,N_2884,N_4803);
nand U9849 (N_9849,N_4736,N_4720);
and U9850 (N_9850,N_2302,N_112);
xnor U9851 (N_9851,N_4739,N_2466);
and U9852 (N_9852,N_3597,N_2011);
and U9853 (N_9853,N_2047,N_312);
nor U9854 (N_9854,N_337,N_344);
nand U9855 (N_9855,N_4484,N_3194);
and U9856 (N_9856,N_2401,N_3466);
xor U9857 (N_9857,N_951,N_3526);
or U9858 (N_9858,N_4846,N_4173);
nor U9859 (N_9859,N_3302,N_681);
xor U9860 (N_9860,N_2584,N_2399);
or U9861 (N_9861,N_614,N_1797);
nand U9862 (N_9862,N_2387,N_3179);
or U9863 (N_9863,N_600,N_2033);
xor U9864 (N_9864,N_4050,N_863);
and U9865 (N_9865,N_4273,N_2627);
xor U9866 (N_9866,N_836,N_2451);
and U9867 (N_9867,N_4134,N_513);
and U9868 (N_9868,N_4840,N_2368);
and U9869 (N_9869,N_2731,N_2529);
and U9870 (N_9870,N_2291,N_2146);
xnor U9871 (N_9871,N_3834,N_4521);
nand U9872 (N_9872,N_609,N_1861);
nor U9873 (N_9873,N_3276,N_956);
xor U9874 (N_9874,N_3180,N_4501);
or U9875 (N_9875,N_989,N_4121);
and U9876 (N_9876,N_540,N_1045);
nor U9877 (N_9877,N_4070,N_3156);
and U9878 (N_9878,N_3275,N_3729);
and U9879 (N_9879,N_1412,N_205);
nor U9880 (N_9880,N_2971,N_2096);
nor U9881 (N_9881,N_3253,N_994);
and U9882 (N_9882,N_2763,N_3458);
xnor U9883 (N_9883,N_491,N_1694);
nand U9884 (N_9884,N_380,N_4338);
and U9885 (N_9885,N_4901,N_1965);
nand U9886 (N_9886,N_1320,N_2625);
or U9887 (N_9887,N_963,N_4183);
nand U9888 (N_9888,N_3927,N_3349);
and U9889 (N_9889,N_3829,N_3988);
and U9890 (N_9890,N_4176,N_407);
nor U9891 (N_9891,N_1816,N_4697);
xnor U9892 (N_9892,N_1374,N_362);
or U9893 (N_9893,N_3371,N_1178);
and U9894 (N_9894,N_2053,N_4411);
nand U9895 (N_9895,N_1476,N_4492);
nand U9896 (N_9896,N_2482,N_3938);
xor U9897 (N_9897,N_3563,N_1961);
and U9898 (N_9898,N_4589,N_4688);
nand U9899 (N_9899,N_2508,N_2496);
or U9900 (N_9900,N_2123,N_4041);
and U9901 (N_9901,N_4754,N_2492);
nor U9902 (N_9902,N_4845,N_2436);
and U9903 (N_9903,N_1001,N_1122);
and U9904 (N_9904,N_2222,N_229);
or U9905 (N_9905,N_2980,N_4764);
nor U9906 (N_9906,N_198,N_2790);
nor U9907 (N_9907,N_3989,N_3583);
or U9908 (N_9908,N_3892,N_943);
xor U9909 (N_9909,N_987,N_3097);
or U9910 (N_9910,N_1030,N_2122);
or U9911 (N_9911,N_307,N_2273);
nor U9912 (N_9912,N_4645,N_1328);
or U9913 (N_9913,N_833,N_3244);
and U9914 (N_9914,N_1419,N_695);
nand U9915 (N_9915,N_3729,N_576);
xor U9916 (N_9916,N_3326,N_1398);
nand U9917 (N_9917,N_3961,N_4774);
nand U9918 (N_9918,N_1844,N_3127);
or U9919 (N_9919,N_2518,N_2200);
nand U9920 (N_9920,N_1381,N_3871);
and U9921 (N_9921,N_3182,N_3114);
nand U9922 (N_9922,N_2537,N_249);
nand U9923 (N_9923,N_3923,N_491);
nand U9924 (N_9924,N_2054,N_1948);
or U9925 (N_9925,N_3874,N_1204);
or U9926 (N_9926,N_3757,N_424);
xor U9927 (N_9927,N_4558,N_1179);
nand U9928 (N_9928,N_4378,N_3403);
nor U9929 (N_9929,N_1200,N_805);
nor U9930 (N_9930,N_3189,N_1629);
nor U9931 (N_9931,N_4948,N_298);
xnor U9932 (N_9932,N_4535,N_860);
nor U9933 (N_9933,N_4807,N_2535);
nand U9934 (N_9934,N_2430,N_4434);
and U9935 (N_9935,N_3138,N_1299);
xor U9936 (N_9936,N_2119,N_1865);
or U9937 (N_9937,N_3087,N_4256);
nand U9938 (N_9938,N_3963,N_3205);
nor U9939 (N_9939,N_3963,N_1630);
and U9940 (N_9940,N_2627,N_4314);
nand U9941 (N_9941,N_2154,N_2237);
nor U9942 (N_9942,N_3179,N_2808);
nor U9943 (N_9943,N_2724,N_4902);
nand U9944 (N_9944,N_4325,N_84);
xnor U9945 (N_9945,N_2901,N_3177);
nand U9946 (N_9946,N_4684,N_3989);
nor U9947 (N_9947,N_1448,N_3728);
nand U9948 (N_9948,N_4200,N_3779);
nand U9949 (N_9949,N_3858,N_4412);
and U9950 (N_9950,N_570,N_292);
and U9951 (N_9951,N_217,N_1619);
xor U9952 (N_9952,N_2722,N_1770);
or U9953 (N_9953,N_3038,N_1732);
xnor U9954 (N_9954,N_1965,N_1392);
or U9955 (N_9955,N_1540,N_2750);
and U9956 (N_9956,N_2313,N_600);
nand U9957 (N_9957,N_2596,N_430);
or U9958 (N_9958,N_1632,N_4433);
nand U9959 (N_9959,N_3978,N_1931);
nand U9960 (N_9960,N_2084,N_702);
nor U9961 (N_9961,N_1447,N_10);
and U9962 (N_9962,N_1985,N_3482);
or U9963 (N_9963,N_3532,N_1854);
nor U9964 (N_9964,N_4913,N_4453);
xnor U9965 (N_9965,N_2221,N_2830);
and U9966 (N_9966,N_2941,N_438);
or U9967 (N_9967,N_1837,N_1091);
and U9968 (N_9968,N_4041,N_1967);
nand U9969 (N_9969,N_2758,N_3300);
nor U9970 (N_9970,N_3518,N_4997);
or U9971 (N_9971,N_3934,N_2842);
and U9972 (N_9972,N_1861,N_3587);
nor U9973 (N_9973,N_2249,N_4338);
nor U9974 (N_9974,N_1526,N_3461);
and U9975 (N_9975,N_2277,N_2741);
nor U9976 (N_9976,N_2461,N_776);
or U9977 (N_9977,N_3850,N_1872);
and U9978 (N_9978,N_1706,N_1256);
and U9979 (N_9979,N_2980,N_4819);
nor U9980 (N_9980,N_1005,N_2484);
nand U9981 (N_9981,N_3299,N_283);
or U9982 (N_9982,N_4300,N_906);
nor U9983 (N_9983,N_818,N_3857);
nor U9984 (N_9984,N_2941,N_4026);
or U9985 (N_9985,N_3521,N_1752);
xor U9986 (N_9986,N_2034,N_817);
or U9987 (N_9987,N_4037,N_2554);
or U9988 (N_9988,N_1799,N_1652);
nor U9989 (N_9989,N_4434,N_3881);
and U9990 (N_9990,N_4767,N_1436);
nand U9991 (N_9991,N_924,N_2329);
and U9992 (N_9992,N_2341,N_2487);
or U9993 (N_9993,N_3130,N_4356);
and U9994 (N_9994,N_36,N_1774);
xnor U9995 (N_9995,N_450,N_3105);
xor U9996 (N_9996,N_3973,N_2640);
nor U9997 (N_9997,N_3929,N_4114);
or U9998 (N_9998,N_2323,N_2225);
and U9999 (N_9999,N_3982,N_2557);
xor U10000 (N_10000,N_9044,N_9198);
and U10001 (N_10001,N_6371,N_9048);
or U10002 (N_10002,N_9689,N_5008);
and U10003 (N_10003,N_9249,N_9751);
and U10004 (N_10004,N_8570,N_5469);
nand U10005 (N_10005,N_9371,N_9327);
nand U10006 (N_10006,N_9428,N_7681);
and U10007 (N_10007,N_7096,N_5012);
and U10008 (N_10008,N_5103,N_5989);
and U10009 (N_10009,N_9370,N_8354);
and U10010 (N_10010,N_8390,N_6117);
or U10011 (N_10011,N_6504,N_7936);
or U10012 (N_10012,N_6287,N_9638);
and U10013 (N_10013,N_9779,N_8759);
xor U10014 (N_10014,N_7359,N_9684);
or U10015 (N_10015,N_7308,N_6307);
nand U10016 (N_10016,N_7849,N_9499);
and U10017 (N_10017,N_5742,N_6116);
and U10018 (N_10018,N_5621,N_8542);
nand U10019 (N_10019,N_9448,N_7589);
and U10020 (N_10020,N_6545,N_7387);
nor U10021 (N_10021,N_9395,N_5860);
nor U10022 (N_10022,N_6482,N_5306);
nand U10023 (N_10023,N_8822,N_8079);
and U10024 (N_10024,N_5874,N_8655);
nor U10025 (N_10025,N_7874,N_8018);
xor U10026 (N_10026,N_8474,N_5245);
xor U10027 (N_10027,N_6831,N_9136);
or U10028 (N_10028,N_6904,N_6212);
nand U10029 (N_10029,N_8497,N_5142);
xnor U10030 (N_10030,N_6632,N_6842);
xor U10031 (N_10031,N_5633,N_7323);
xor U10032 (N_10032,N_8604,N_9899);
and U10033 (N_10033,N_7048,N_6011);
and U10034 (N_10034,N_8836,N_8156);
or U10035 (N_10035,N_6685,N_6568);
or U10036 (N_10036,N_7971,N_6706);
or U10037 (N_10037,N_7859,N_9995);
xor U10038 (N_10038,N_8954,N_6666);
xnor U10039 (N_10039,N_6923,N_7367);
nor U10040 (N_10040,N_8033,N_7126);
nor U10041 (N_10041,N_7315,N_6939);
xnor U10042 (N_10042,N_9766,N_9404);
and U10043 (N_10043,N_8064,N_5506);
nor U10044 (N_10044,N_5180,N_8870);
and U10045 (N_10045,N_5525,N_8402);
nor U10046 (N_10046,N_9208,N_5852);
nand U10047 (N_10047,N_5848,N_8324);
xor U10048 (N_10048,N_7947,N_7610);
nor U10049 (N_10049,N_8806,N_7366);
nor U10050 (N_10050,N_7214,N_5992);
or U10051 (N_10051,N_5945,N_5671);
or U10052 (N_10052,N_7811,N_6674);
xor U10053 (N_10053,N_6669,N_8588);
nor U10054 (N_10054,N_7292,N_6910);
xnor U10055 (N_10055,N_8971,N_5831);
or U10056 (N_10056,N_6898,N_5734);
nand U10057 (N_10057,N_6886,N_6094);
and U10058 (N_10058,N_5825,N_6384);
nor U10059 (N_10059,N_5712,N_9469);
nor U10060 (N_10060,N_5604,N_5272);
or U10061 (N_10061,N_9944,N_6259);
nand U10062 (N_10062,N_7021,N_9292);
and U10063 (N_10063,N_6266,N_8353);
or U10064 (N_10064,N_7817,N_9719);
nand U10065 (N_10065,N_7412,N_5805);
nor U10066 (N_10066,N_7599,N_9980);
or U10067 (N_10067,N_8272,N_6804);
or U10068 (N_10068,N_9966,N_5169);
xor U10069 (N_10069,N_5987,N_9456);
nor U10070 (N_10070,N_5079,N_5188);
nor U10071 (N_10071,N_9425,N_6148);
nand U10072 (N_10072,N_8919,N_5045);
and U10073 (N_10073,N_6986,N_9098);
and U10074 (N_10074,N_6142,N_6090);
xnor U10075 (N_10075,N_5637,N_9118);
nand U10076 (N_10076,N_9313,N_9608);
nor U10077 (N_10077,N_6678,N_8879);
nor U10078 (N_10078,N_7889,N_9884);
xnor U10079 (N_10079,N_5190,N_9713);
and U10080 (N_10080,N_9837,N_8608);
and U10081 (N_10081,N_6047,N_7683);
and U10082 (N_10082,N_8916,N_5206);
or U10083 (N_10083,N_7511,N_7954);
nor U10084 (N_10084,N_6022,N_5819);
xor U10085 (N_10085,N_6583,N_7437);
nor U10086 (N_10086,N_5226,N_7180);
nor U10087 (N_10087,N_9345,N_8055);
xor U10088 (N_10088,N_6314,N_6777);
xnor U10089 (N_10089,N_8467,N_9380);
or U10090 (N_10090,N_6593,N_7747);
and U10091 (N_10091,N_8847,N_8125);
nand U10092 (N_10092,N_9527,N_5127);
and U10093 (N_10093,N_7446,N_7306);
nand U10094 (N_10094,N_5870,N_9673);
or U10095 (N_10095,N_9969,N_8465);
or U10096 (N_10096,N_9300,N_5577);
or U10097 (N_10097,N_6869,N_5539);
nor U10098 (N_10098,N_9488,N_8789);
nand U10099 (N_10099,N_8453,N_6378);
nor U10100 (N_10100,N_7415,N_9374);
nor U10101 (N_10101,N_6549,N_6636);
xor U10102 (N_10102,N_7627,N_7647);
nand U10103 (N_10103,N_8974,N_6942);
nor U10104 (N_10104,N_5751,N_8152);
or U10105 (N_10105,N_6346,N_7503);
or U10106 (N_10106,N_6931,N_7582);
and U10107 (N_10107,N_6229,N_6269);
nor U10108 (N_10108,N_7287,N_9815);
or U10109 (N_10109,N_6106,N_7790);
or U10110 (N_10110,N_5010,N_5707);
or U10111 (N_10111,N_6386,N_5051);
xor U10112 (N_10112,N_7901,N_5849);
and U10113 (N_10113,N_5919,N_7029);
and U10114 (N_10114,N_8449,N_8308);
or U10115 (N_10115,N_7091,N_7536);
or U10116 (N_10116,N_8020,N_9343);
nand U10117 (N_10117,N_6780,N_7893);
nand U10118 (N_10118,N_9976,N_7602);
and U10119 (N_10119,N_6885,N_7429);
nor U10120 (N_10120,N_7320,N_5823);
xor U10121 (N_10121,N_9341,N_6256);
nor U10122 (N_10122,N_9549,N_5954);
and U10123 (N_10123,N_5075,N_6396);
xor U10124 (N_10124,N_7912,N_9872);
or U10125 (N_10125,N_5981,N_5664);
nor U10126 (N_10126,N_9493,N_9718);
and U10127 (N_10127,N_9591,N_5465);
and U10128 (N_10128,N_7679,N_8809);
or U10129 (N_10129,N_9619,N_9737);
or U10130 (N_10130,N_8006,N_9229);
and U10131 (N_10131,N_6498,N_8294);
and U10132 (N_10132,N_7127,N_8635);
xor U10133 (N_10133,N_8163,N_8984);
and U10134 (N_10134,N_5474,N_8735);
xor U10135 (N_10135,N_5351,N_6121);
xnor U10136 (N_10136,N_8729,N_8948);
xnor U10137 (N_10137,N_7239,N_8365);
or U10138 (N_10138,N_5162,N_8179);
nor U10139 (N_10139,N_7333,N_8867);
or U10140 (N_10140,N_8382,N_8446);
nand U10141 (N_10141,N_5027,N_9741);
xnor U10142 (N_10142,N_7550,N_6155);
xnor U10143 (N_10143,N_6356,N_6213);
nand U10144 (N_10144,N_5126,N_6963);
or U10145 (N_10145,N_7656,N_5341);
or U10146 (N_10146,N_9419,N_7077);
nand U10147 (N_10147,N_5523,N_7364);
nand U10148 (N_10148,N_8337,N_8910);
nand U10149 (N_10149,N_5962,N_8469);
nand U10150 (N_10150,N_8917,N_7116);
and U10151 (N_10151,N_6203,N_5387);
and U10152 (N_10152,N_7153,N_9631);
xor U10153 (N_10153,N_6895,N_5236);
xor U10154 (N_10154,N_7355,N_6354);
or U10155 (N_10155,N_9334,N_8464);
nand U10156 (N_10156,N_8201,N_7211);
xor U10157 (N_10157,N_6349,N_9784);
nor U10158 (N_10158,N_8439,N_5301);
or U10159 (N_10159,N_5266,N_9353);
or U10160 (N_10160,N_6751,N_5533);
nor U10161 (N_10161,N_6360,N_7275);
or U10162 (N_10162,N_6451,N_7813);
nor U10163 (N_10163,N_5456,N_9150);
nand U10164 (N_10164,N_5723,N_7965);
nor U10165 (N_10165,N_7402,N_8805);
nor U10166 (N_10166,N_5388,N_6063);
or U10167 (N_10167,N_5367,N_9926);
nor U10168 (N_10168,N_6864,N_6889);
xor U10169 (N_10169,N_5099,N_6393);
nand U10170 (N_10170,N_6171,N_7770);
nand U10171 (N_10171,N_7278,N_6702);
xor U10172 (N_10172,N_5448,N_5714);
xnor U10173 (N_10173,N_9546,N_7809);
or U10174 (N_10174,N_9935,N_8673);
xnor U10175 (N_10175,N_8621,N_9536);
nor U10176 (N_10176,N_5885,N_7959);
xnor U10177 (N_10177,N_7869,N_6459);
xor U10178 (N_10178,N_9145,N_8719);
xor U10179 (N_10179,N_5338,N_7976);
or U10180 (N_10180,N_8244,N_6007);
or U10181 (N_10181,N_9955,N_9682);
nand U10182 (N_10182,N_7798,N_9242);
or U10183 (N_10183,N_6855,N_6736);
nor U10184 (N_10184,N_9207,N_9644);
nor U10185 (N_10185,N_9927,N_7110);
or U10186 (N_10186,N_9250,N_5763);
or U10187 (N_10187,N_8320,N_5078);
nand U10188 (N_10188,N_6437,N_5749);
nor U10189 (N_10189,N_9683,N_6714);
xor U10190 (N_10190,N_6773,N_9418);
nor U10191 (N_10191,N_9595,N_9728);
xor U10192 (N_10192,N_6873,N_9765);
or U10193 (N_10193,N_9530,N_6529);
or U10194 (N_10194,N_8059,N_9480);
or U10195 (N_10195,N_7439,N_7873);
nand U10196 (N_10196,N_5537,N_7265);
nand U10197 (N_10197,N_7114,N_7611);
or U10198 (N_10198,N_5186,N_7777);
nand U10199 (N_10199,N_9964,N_9065);
nor U10200 (N_10200,N_5313,N_7184);
and U10201 (N_10201,N_9059,N_7396);
nand U10202 (N_10202,N_9584,N_7062);
nand U10203 (N_10203,N_6077,N_7067);
nand U10204 (N_10204,N_6132,N_8685);
nor U10205 (N_10205,N_5554,N_5513);
and U10206 (N_10206,N_5166,N_5106);
xor U10207 (N_10207,N_6660,N_9285);
xnor U10208 (N_10208,N_5959,N_7187);
or U10209 (N_10209,N_6173,N_9729);
nor U10210 (N_10210,N_8060,N_7887);
or U10211 (N_10211,N_7150,N_9568);
nand U10212 (N_10212,N_7090,N_6536);
or U10213 (N_10213,N_8691,N_7102);
nor U10214 (N_10214,N_5298,N_7175);
or U10215 (N_10215,N_9951,N_7023);
nor U10216 (N_10216,N_9756,N_6818);
nor U10217 (N_10217,N_9175,N_5251);
nor U10218 (N_10218,N_6357,N_5558);
nor U10219 (N_10219,N_9110,N_8263);
and U10220 (N_10220,N_6958,N_5455);
and U10221 (N_10221,N_6561,N_6535);
nand U10222 (N_10222,N_5982,N_6774);
and U10223 (N_10223,N_6065,N_6091);
or U10224 (N_10224,N_8733,N_6084);
nor U10225 (N_10225,N_6646,N_5678);
and U10226 (N_10226,N_9047,N_8275);
nand U10227 (N_10227,N_8702,N_9776);
xnor U10228 (N_10228,N_5071,N_9852);
or U10229 (N_10229,N_9318,N_7016);
or U10230 (N_10230,N_7216,N_7092);
and U10231 (N_10231,N_5591,N_6581);
xor U10232 (N_10232,N_6595,N_5203);
nand U10233 (N_10233,N_8025,N_6806);
nand U10234 (N_10234,N_9535,N_6683);
nand U10235 (N_10235,N_5667,N_5917);
and U10236 (N_10236,N_7422,N_9795);
and U10237 (N_10237,N_5590,N_5691);
nand U10238 (N_10238,N_8440,N_7009);
xor U10239 (N_10239,N_9213,N_5787);
and U10240 (N_10240,N_9898,N_8953);
xnor U10241 (N_10241,N_9303,N_6093);
nor U10242 (N_10242,N_9339,N_8569);
or U10243 (N_10243,N_5312,N_8958);
and U10244 (N_10244,N_7946,N_6402);
nand U10245 (N_10245,N_9509,N_6273);
nand U10246 (N_10246,N_7693,N_8622);
nand U10247 (N_10247,N_7833,N_8577);
or U10248 (N_10248,N_7558,N_8098);
nor U10249 (N_10249,N_6756,N_6737);
or U10250 (N_10250,N_6596,N_8716);
and U10251 (N_10251,N_9062,N_6291);
nor U10252 (N_10252,N_6537,N_5391);
nand U10253 (N_10253,N_9986,N_7230);
nor U10254 (N_10254,N_7407,N_8457);
nor U10255 (N_10255,N_5655,N_5960);
xor U10256 (N_10256,N_5949,N_9476);
nor U10257 (N_10257,N_5891,N_9262);
nor U10258 (N_10258,N_9900,N_6060);
xor U10259 (N_10259,N_7988,N_9632);
nand U10260 (N_10260,N_5610,N_6410);
nor U10261 (N_10261,N_9650,N_7049);
and U10262 (N_10262,N_7913,N_8739);
nor U10263 (N_10263,N_5555,N_7725);
or U10264 (N_10264,N_8319,N_5116);
nor U10265 (N_10265,N_6005,N_5969);
nor U10266 (N_10266,N_5845,N_8146);
nand U10267 (N_10267,N_5973,N_9954);
nand U10268 (N_10268,N_5517,N_9794);
nand U10269 (N_10269,N_6779,N_6131);
nor U10270 (N_10270,N_9646,N_8034);
or U10271 (N_10271,N_6486,N_7181);
or U10272 (N_10272,N_7806,N_8723);
nor U10273 (N_10273,N_6692,N_6882);
or U10274 (N_10274,N_6210,N_5185);
nand U10275 (N_10275,N_9426,N_6358);
nor U10276 (N_10276,N_5725,N_5606);
nor U10277 (N_10277,N_7515,N_8500);
xor U10278 (N_10278,N_7152,N_8232);
nand U10279 (N_10279,N_6485,N_5735);
nand U10280 (N_10280,N_8782,N_5508);
and U10281 (N_10281,N_5481,N_7842);
nand U10282 (N_10282,N_5853,N_5473);
xor U10283 (N_10283,N_8835,N_6381);
and U10284 (N_10284,N_6871,N_9486);
and U10285 (N_10285,N_7236,N_6071);
and U10286 (N_10286,N_7022,N_5627);
or U10287 (N_10287,N_9227,N_5977);
nand U10288 (N_10288,N_6341,N_5109);
nand U10289 (N_10289,N_7424,N_9709);
and U10290 (N_10290,N_8221,N_9373);
nand U10291 (N_10291,N_9305,N_6681);
nand U10292 (N_10292,N_6829,N_7937);
nand U10293 (N_10293,N_5899,N_9037);
nand U10294 (N_10294,N_5785,N_7970);
xor U10295 (N_10295,N_5731,N_8385);
nand U10296 (N_10296,N_8398,N_9447);
xnor U10297 (N_10297,N_6503,N_8821);
xnor U10298 (N_10298,N_9063,N_6709);
nand U10299 (N_10299,N_6096,N_5929);
nand U10300 (N_10300,N_5175,N_7232);
xor U10301 (N_10301,N_8321,N_6230);
xnor U10302 (N_10302,N_6563,N_6987);
xor U10303 (N_10303,N_9093,N_8498);
nor U10304 (N_10304,N_9695,N_9721);
and U10305 (N_10305,N_8829,N_6530);
xnor U10306 (N_10306,N_8371,N_8892);
or U10307 (N_10307,N_5578,N_9272);
or U10308 (N_10308,N_7358,N_5457);
nor U10309 (N_10309,N_9519,N_5529);
xnor U10310 (N_10310,N_6363,N_7768);
and U10311 (N_10311,N_6615,N_5068);
nor U10312 (N_10312,N_9687,N_8734);
or U10313 (N_10313,N_8259,N_5327);
and U10314 (N_10314,N_6419,N_7646);
xnor U10315 (N_10315,N_5824,N_8400);
or U10316 (N_10316,N_7784,N_6231);
nor U10317 (N_10317,N_5613,N_9026);
nor U10318 (N_10318,N_5993,N_9775);
nor U10319 (N_10319,N_9844,N_9102);
and U10320 (N_10320,N_9886,N_6604);
or U10321 (N_10321,N_9885,N_5470);
nor U10322 (N_10322,N_8462,N_6207);
or U10323 (N_10323,N_9176,N_5101);
xor U10324 (N_10324,N_6334,N_9203);
nor U10325 (N_10325,N_9551,N_5946);
xnor U10326 (N_10326,N_6150,N_5693);
or U10327 (N_10327,N_6279,N_7303);
nand U10328 (N_10328,N_9726,N_5161);
or U10329 (N_10329,N_8786,N_8514);
and U10330 (N_10330,N_8965,N_9321);
nand U10331 (N_10331,N_8743,N_6425);
and U10332 (N_10332,N_6301,N_9114);
nor U10333 (N_10333,N_7998,N_5717);
nor U10334 (N_10334,N_7186,N_8442);
nand U10335 (N_10335,N_5672,N_6978);
xor U10336 (N_10336,N_6754,N_6560);
nor U10337 (N_10337,N_7860,N_8862);
xor U10338 (N_10338,N_8959,N_9479);
and U10339 (N_10339,N_6226,N_6708);
and U10340 (N_10340,N_9335,N_5400);
xor U10341 (N_10341,N_9280,N_5365);
xor U10342 (N_10342,N_5795,N_7399);
nor U10343 (N_10343,N_5278,N_9802);
xor U10344 (N_10344,N_6211,N_7888);
nor U10345 (N_10345,N_9574,N_8136);
and U10346 (N_10346,N_7018,N_7989);
or U10347 (N_10347,N_6523,N_6282);
nand U10348 (N_10348,N_6555,N_6032);
nor U10349 (N_10349,N_7587,N_5141);
nand U10350 (N_10350,N_6979,N_8425);
and U10351 (N_10351,N_5256,N_6786);
nand U10352 (N_10352,N_5253,N_5938);
or U10353 (N_10353,N_9130,N_5786);
nand U10354 (N_10354,N_7196,N_6748);
nand U10355 (N_10355,N_5440,N_7072);
xnor U10356 (N_10356,N_6020,N_8317);
xor U10357 (N_10357,N_9829,N_5883);
nor U10358 (N_10358,N_9609,N_9391);
and U10359 (N_10359,N_8128,N_7204);
nor U10360 (N_10360,N_5348,N_5738);
nor U10361 (N_10361,N_7548,N_8812);
or U10362 (N_10362,N_7256,N_5295);
or U10363 (N_10363,N_9038,N_9538);
or U10364 (N_10364,N_8900,N_8150);
and U10365 (N_10365,N_6329,N_9874);
nand U10366 (N_10366,N_8473,N_8127);
and U10367 (N_10367,N_8920,N_7138);
or U10368 (N_10368,N_6033,N_6470);
and U10369 (N_10369,N_7738,N_7604);
xnor U10370 (N_10370,N_5893,N_8857);
or U10371 (N_10371,N_6543,N_6006);
and U10372 (N_10372,N_6479,N_9274);
or U10373 (N_10373,N_5096,N_8684);
nand U10374 (N_10374,N_8423,N_6608);
and U10375 (N_10375,N_9032,N_9464);
xor U10376 (N_10376,N_5050,N_6924);
and U10377 (N_10377,N_5730,N_8672);
nand U10378 (N_10378,N_7815,N_6696);
xor U10379 (N_10379,N_7793,N_9139);
and U10380 (N_10380,N_8504,N_5417);
xor U10381 (N_10381,N_9733,N_9645);
nor U10382 (N_10382,N_5896,N_7735);
nand U10383 (N_10383,N_6526,N_9006);
nand U10384 (N_10384,N_7246,N_9155);
nand U10385 (N_10385,N_6981,N_7782);
nor U10386 (N_10386,N_6614,N_7004);
nor U10387 (N_10387,N_7455,N_6110);
and U10388 (N_10388,N_8662,N_5361);
nand U10389 (N_10389,N_8468,N_7146);
nand U10390 (N_10390,N_6176,N_5368);
or U10391 (N_10391,N_9873,N_6083);
or U10392 (N_10392,N_9381,N_9581);
nand U10393 (N_10393,N_7339,N_6455);
xor U10394 (N_10394,N_8051,N_5472);
or U10395 (N_10395,N_6388,N_7019);
xor U10396 (N_10396,N_7791,N_9501);
or U10397 (N_10397,N_6687,N_6477);
or U10398 (N_10398,N_6799,N_9841);
nor U10399 (N_10399,N_9972,N_5005);
xnor U10400 (N_10400,N_8676,N_7002);
xnor U10401 (N_10401,N_5724,N_8709);
nand U10402 (N_10402,N_8798,N_5399);
and U10403 (N_10403,N_8488,N_8929);
nand U10404 (N_10404,N_8600,N_6122);
xor U10405 (N_10405,N_6901,N_6613);
nor U10406 (N_10406,N_6957,N_8664);
nor U10407 (N_10407,N_6832,N_9366);
nor U10408 (N_10408,N_9553,N_8630);
xnor U10409 (N_10409,N_8566,N_8036);
xnor U10410 (N_10410,N_9962,N_9012);
nor U10411 (N_10411,N_7933,N_5176);
and U10412 (N_10412,N_8800,N_7968);
and U10413 (N_10413,N_8188,N_9291);
nand U10414 (N_10414,N_8346,N_6299);
xor U10415 (N_10415,N_6438,N_9836);
nor U10416 (N_10416,N_9035,N_9563);
and U10417 (N_10417,N_8381,N_7923);
or U10418 (N_10418,N_7928,N_7173);
nand U10419 (N_10419,N_8027,N_7567);
or U10420 (N_10420,N_7089,N_9758);
or U10421 (N_10421,N_6571,N_7969);
nor U10422 (N_10422,N_8582,N_5225);
xnor U10423 (N_10423,N_9314,N_8225);
nand U10424 (N_10424,N_8138,N_9813);
xnor U10425 (N_10425,N_6190,N_8489);
and U10426 (N_10426,N_8891,N_7519);
or U10427 (N_10427,N_6265,N_9902);
nor U10428 (N_10428,N_9140,N_7420);
xor U10429 (N_10429,N_7578,N_5854);
or U10430 (N_10430,N_5665,N_8979);
or U10431 (N_10431,N_5733,N_7373);
nand U10432 (N_10432,N_7159,N_6056);
or U10433 (N_10433,N_8070,N_6919);
nor U10434 (N_10434,N_7122,N_9624);
and U10435 (N_10435,N_9611,N_7316);
nand U10436 (N_10436,N_6625,N_9316);
and U10437 (N_10437,N_7348,N_9671);
or U10438 (N_10438,N_9296,N_5028);
xor U10439 (N_10439,N_5252,N_5450);
or U10440 (N_10440,N_6463,N_7994);
nor U10441 (N_10441,N_8993,N_8174);
nor U10442 (N_10442,N_6174,N_5489);
or U10443 (N_10443,N_7561,N_5437);
nor U10444 (N_10444,N_9070,N_9166);
nand U10445 (N_10445,N_5454,N_8625);
nand U10446 (N_10446,N_6713,N_9491);
or U10447 (N_10447,N_5970,N_7244);
nand U10448 (N_10448,N_5697,N_8714);
nand U10449 (N_10449,N_6562,N_7631);
nor U10450 (N_10450,N_7950,N_6186);
nand U10451 (N_10451,N_6264,N_6735);
nand U10452 (N_10452,N_6680,N_8196);
and U10453 (N_10453,N_6544,N_9512);
nor U10454 (N_10454,N_6743,N_9979);
xnor U10455 (N_10455,N_7593,N_5641);
or U10456 (N_10456,N_8115,N_8192);
nand U10457 (N_10457,N_5422,N_7496);
or U10458 (N_10458,N_7450,N_6701);
nand U10459 (N_10459,N_7466,N_6344);
and U10460 (N_10460,N_9803,N_7207);
or U10461 (N_10461,N_7592,N_8161);
and U10462 (N_10462,N_6461,N_5828);
and U10463 (N_10463,N_7565,N_9005);
or U10464 (N_10464,N_6192,N_7034);
xor U10465 (N_10465,N_8536,N_7288);
nor U10466 (N_10466,N_5014,N_7046);
nor U10467 (N_10467,N_5102,N_6817);
nand U10468 (N_10468,N_5215,N_8640);
and U10469 (N_10469,N_8022,N_5342);
nor U10470 (N_10470,N_6100,N_5385);
xor U10471 (N_10471,N_8191,N_7866);
xor U10472 (N_10472,N_6631,N_8532);
nand U10473 (N_10473,N_7036,N_7013);
or U10474 (N_10474,N_8545,N_7231);
and U10475 (N_10475,N_9503,N_5560);
xnor U10476 (N_10476,N_9889,N_7635);
nand U10477 (N_10477,N_9787,N_6087);
and U10478 (N_10478,N_5031,N_7545);
xnor U10479 (N_10479,N_7774,N_6932);
and U10480 (N_10480,N_9311,N_8853);
or U10481 (N_10481,N_5497,N_9903);
nand U10482 (N_10482,N_6367,N_8361);
xnor U10483 (N_10483,N_5940,N_8763);
and U10484 (N_10484,N_7573,N_8963);
and U10485 (N_10485,N_6390,N_7751);
nand U10486 (N_10486,N_5413,N_6682);
nand U10487 (N_10487,N_9210,N_6883);
nor U10488 (N_10488,N_7063,N_5006);
xor U10489 (N_10489,N_8922,N_6950);
nor U10490 (N_10490,N_9801,N_5895);
nor U10491 (N_10491,N_8384,N_6913);
and U10492 (N_10492,N_7020,N_9994);
nor U10493 (N_10493,N_7840,N_6172);
nand U10494 (N_10494,N_9736,N_5543);
xnor U10495 (N_10495,N_8680,N_5189);
xor U10496 (N_10496,N_5131,N_5813);
nand U10497 (N_10497,N_6689,N_5906);
or U10498 (N_10498,N_7961,N_6618);
nand U10499 (N_10499,N_5257,N_5685);
or U10500 (N_10500,N_7890,N_7271);
or U10501 (N_10501,N_5722,N_8396);
nor U10502 (N_10502,N_9061,N_6741);
nand U10503 (N_10503,N_9759,N_5330);
xor U10504 (N_10504,N_5952,N_8037);
or U10505 (N_10505,N_9298,N_8675);
nor U10506 (N_10506,N_5037,N_9372);
nand U10507 (N_10507,N_7277,N_7942);
xor U10508 (N_10508,N_7403,N_6415);
or U10509 (N_10509,N_6428,N_6602);
xor U10510 (N_10510,N_8681,N_5409);
nand U10511 (N_10511,N_5441,N_7780);
xnor U10512 (N_10512,N_5767,N_6721);
or U10513 (N_10513,N_6490,N_8135);
or U10514 (N_10514,N_5300,N_8978);
and U10515 (N_10515,N_5663,N_5198);
or U10516 (N_10516,N_9990,N_7796);
nand U10517 (N_10517,N_7480,N_5652);
and U10518 (N_10518,N_7907,N_5863);
nand U10519 (N_10519,N_8141,N_7397);
nor U10520 (N_10520,N_7224,N_9664);
or U10521 (N_10521,N_8615,N_6216);
or U10522 (N_10522,N_7234,N_7058);
nor U10523 (N_10523,N_5237,N_8073);
nor U10524 (N_10524,N_5337,N_5262);
or U10525 (N_10525,N_7624,N_8243);
nor U10526 (N_10526,N_9606,N_8181);
nor U10527 (N_10527,N_6487,N_7956);
and U10528 (N_10528,N_5748,N_9573);
nor U10529 (N_10529,N_6260,N_9982);
nor U10530 (N_10530,N_7017,N_7409);
or U10531 (N_10531,N_8831,N_8246);
or U10532 (N_10532,N_8200,N_8775);
xor U10533 (N_10533,N_6025,N_9396);
nor U10534 (N_10534,N_6383,N_7434);
xor U10535 (N_10535,N_9961,N_5442);
nor U10536 (N_10536,N_7293,N_6409);
xor U10537 (N_10537,N_5137,N_6058);
nor U10538 (N_10538,N_5283,N_8871);
nand U10539 (N_10539,N_6235,N_8745);
or U10540 (N_10540,N_8634,N_5231);
nor U10541 (N_10541,N_8052,N_9394);
or U10542 (N_10542,N_6611,N_9403);
nor U10543 (N_10543,N_6232,N_7761);
nor U10544 (N_10544,N_5168,N_7031);
xnor U10545 (N_10545,N_7896,N_5209);
or U10546 (N_10546,N_7283,N_9830);
nand U10547 (N_10547,N_8911,N_7705);
and U10548 (N_10548,N_8233,N_7324);
and U10549 (N_10549,N_9919,N_6915);
nand U10550 (N_10550,N_9875,N_6520);
and U10551 (N_10551,N_9120,N_9984);
nand U10552 (N_10552,N_7894,N_7351);
or U10553 (N_10553,N_9622,N_5098);
nor U10554 (N_10554,N_7839,N_8895);
and U10555 (N_10555,N_8944,N_7975);
nand U10556 (N_10556,N_5774,N_5926);
nand U10557 (N_10557,N_6377,N_8293);
nor U10558 (N_10558,N_9217,N_7084);
nand U10559 (N_10559,N_7949,N_6276);
or U10560 (N_10560,N_9185,N_5942);
xor U10561 (N_10561,N_5307,N_6964);
nand U10562 (N_10562,N_5144,N_5356);
nand U10563 (N_10563,N_6342,N_9757);
xor U10564 (N_10564,N_5053,N_5648);
nand U10565 (N_10565,N_9045,N_5043);
or U10566 (N_10566,N_5953,N_8103);
and U10567 (N_10567,N_7273,N_6204);
nand U10568 (N_10568,N_5549,N_6290);
nor U10569 (N_10569,N_8413,N_9705);
and U10570 (N_10570,N_7448,N_8661);
xor U10571 (N_10571,N_6813,N_9168);
or U10572 (N_10572,N_5129,N_6993);
xor U10573 (N_10573,N_7616,N_5377);
or U10574 (N_10574,N_6489,N_5939);
nand U10575 (N_10575,N_5635,N_7922);
or U10576 (N_10576,N_7335,N_5532);
xnor U10577 (N_10577,N_5761,N_8299);
and U10578 (N_10578,N_9735,N_9723);
and U10579 (N_10579,N_6308,N_6202);
nor U10580 (N_10580,N_5898,N_6564);
or U10581 (N_10581,N_6694,N_8864);
xnor U10582 (N_10582,N_5004,N_9011);
or U10583 (N_10583,N_5308,N_8069);
and U10584 (N_10584,N_9111,N_9287);
nor U10585 (N_10585,N_8985,N_7368);
nand U10586 (N_10586,N_6665,N_9599);
xnor U10587 (N_10587,N_6875,N_8747);
or U10588 (N_10588,N_5755,N_8066);
and U10589 (N_10589,N_5158,N_9839);
nand U10590 (N_10590,N_7703,N_6195);
or U10591 (N_10591,N_8392,N_9235);
nand U10592 (N_10592,N_8491,N_6720);
and U10593 (N_10593,N_6297,N_6044);
and U10594 (N_10594,N_8043,N_6826);
and U10595 (N_10595,N_8377,N_9807);
nand U10596 (N_10596,N_9798,N_6182);
or U10597 (N_10597,N_7195,N_5023);
xor U10598 (N_10598,N_7787,N_8517);
nor U10599 (N_10599,N_6123,N_7026);
and U10600 (N_10600,N_5692,N_9251);
nand U10601 (N_10601,N_6413,N_7483);
or U10602 (N_10602,N_6343,N_8254);
nor U10603 (N_10603,N_6900,N_7371);
nand U10604 (N_10604,N_8050,N_8696);
xor U10605 (N_10605,N_8215,N_9420);
and U10606 (N_10606,N_9429,N_9430);
nand U10607 (N_10607,N_5069,N_5526);
or U10608 (N_10608,N_5222,N_7997);
nor U10609 (N_10609,N_7032,N_8652);
or U10610 (N_10610,N_7279,N_9782);
nand U10611 (N_10611,N_8785,N_7132);
nor U10612 (N_10612,N_5013,N_5647);
nor U10613 (N_10613,N_8774,N_5897);
nor U10614 (N_10614,N_7290,N_8715);
nor U10615 (N_10615,N_5115,N_9558);
nand U10616 (N_10616,N_8725,N_8017);
or U10617 (N_10617,N_8303,N_8562);
and U10618 (N_10618,N_6597,N_8445);
nor U10619 (N_10619,N_8405,N_8389);
xnor U10620 (N_10620,N_6234,N_6153);
or U10621 (N_10621,N_8594,N_9556);
and U10622 (N_10622,N_6746,N_7820);
xnor U10623 (N_10623,N_7886,N_6552);
or U10624 (N_10624,N_6816,N_7752);
nor U10625 (N_10625,N_6277,N_9771);
or U10626 (N_10626,N_9620,N_5816);
nand U10627 (N_10627,N_8967,N_5067);
xor U10628 (N_10628,N_7447,N_8162);
and U10629 (N_10629,N_5411,N_6136);
xor U10630 (N_10630,N_9967,N_6368);
and U10631 (N_10631,N_9234,N_7245);
nand U10632 (N_10632,N_9616,N_8679);
xnor U10633 (N_10633,N_7326,N_8996);
and U10634 (N_10634,N_6313,N_6288);
or U10635 (N_10635,N_9522,N_9950);
nor U10636 (N_10636,N_8650,N_5553);
and U10637 (N_10637,N_5458,N_8297);
and U10638 (N_10638,N_5837,N_6532);
nor U10639 (N_10639,N_6464,N_7608);
xnor U10640 (N_10640,N_6000,N_9422);
and U10641 (N_10641,N_8648,N_9744);
nor U10642 (N_10642,N_8779,N_8872);
nand U10643 (N_10643,N_6601,N_9148);
nor U10644 (N_10644,N_9710,N_7743);
xor U10645 (N_10645,N_5081,N_5636);
or U10646 (N_10646,N_8708,N_7711);
and U10647 (N_10647,N_7532,N_5263);
nor U10648 (N_10648,N_9016,N_6525);
and U10649 (N_10649,N_8801,N_8274);
nand U10650 (N_10650,N_7488,N_8370);
and U10651 (N_10651,N_6292,N_7304);
nand U10652 (N_10652,N_8960,N_6655);
or U10653 (N_10653,N_9119,N_7382);
xnor U10654 (N_10654,N_5401,N_6306);
xor U10655 (N_10655,N_7490,N_7615);
xor U10656 (N_10656,N_9040,N_5587);
nand U10657 (N_10657,N_9596,N_6519);
or U10658 (N_10658,N_6651,N_8626);
and U10659 (N_10659,N_5183,N_5502);
xnor U10660 (N_10660,N_7603,N_8632);
and U10661 (N_10661,N_7492,N_8359);
and U10662 (N_10662,N_8599,N_5614);
nor U10663 (N_10663,N_8842,N_7882);
and U10664 (N_10664,N_7107,N_9487);
xor U10665 (N_10665,N_9386,N_6324);
or U10666 (N_10666,N_6730,N_9109);
or U10667 (N_10667,N_7562,N_8595);
nor U10668 (N_10668,N_6350,N_6661);
or U10669 (N_10669,N_8823,N_9490);
xor U10670 (N_10670,N_7826,N_6506);
and U10671 (N_10671,N_9223,N_8781);
nor U10672 (N_10672,N_5381,N_5117);
or U10673 (N_10673,N_5628,N_5971);
xor U10674 (N_10674,N_7870,N_5515);
or U10675 (N_10675,N_5750,N_7540);
nand U10676 (N_10676,N_7139,N_5546);
and U10677 (N_10677,N_6196,N_5133);
or U10678 (N_10678,N_8534,N_8926);
nor U10679 (N_10679,N_5446,N_8342);
xor U10680 (N_10680,N_5376,N_6278);
or U10681 (N_10681,N_9834,N_9892);
nor U10682 (N_10682,N_7479,N_9197);
nor U10683 (N_10683,N_5410,N_8077);
xor U10684 (N_10684,N_7255,N_8989);
or U10685 (N_10685,N_9652,N_7383);
xor U10686 (N_10686,N_8816,N_8572);
or U10687 (N_10687,N_6541,N_7648);
nor U10688 (N_10688,N_6639,N_5623);
nor U10689 (N_10689,N_7321,N_9455);
and U10690 (N_10690,N_8350,N_6421);
xor U10691 (N_10691,N_8799,N_6994);
and U10692 (N_10692,N_9375,N_9764);
or U10693 (N_10693,N_7755,N_6640);
nand U10694 (N_10694,N_6513,N_9135);
and U10695 (N_10695,N_9257,N_5643);
nor U10696 (N_10696,N_7133,N_6125);
nand U10697 (N_10697,N_6243,N_8004);
or U10698 (N_10698,N_8040,N_6586);
or U10699 (N_10699,N_8833,N_7476);
or U10700 (N_10700,N_8825,N_5044);
nor U10701 (N_10701,N_8700,N_9561);
or U10702 (N_10702,N_7141,N_6380);
and U10703 (N_10703,N_7469,N_7411);
xor U10704 (N_10704,N_6382,N_7079);
and U10705 (N_10705,N_8845,N_9400);
or U10706 (N_10706,N_6985,N_9914);
nand U10707 (N_10707,N_7680,N_6331);
xnor U10708 (N_10708,N_8997,N_7374);
or U10709 (N_10709,N_8082,N_5220);
and U10710 (N_10710,N_6258,N_6339);
nand U10711 (N_10711,N_6936,N_5421);
xor U10712 (N_10712,N_8116,N_9157);
or U10713 (N_10713,N_5475,N_5398);
nand U10714 (N_10714,N_8455,N_8969);
nor U10715 (N_10715,N_7783,N_5644);
nand U10716 (N_10716,N_9009,N_7987);
and U10717 (N_10717,N_6101,N_9471);
or U10718 (N_10718,N_7066,N_7272);
and U10719 (N_10719,N_8452,N_9812);
xor U10720 (N_10720,N_8357,N_7846);
nand U10721 (N_10721,N_8435,N_7865);
nand U10722 (N_10722,N_8726,N_6145);
xor U10723 (N_10723,N_8424,N_8591);
nor U10724 (N_10724,N_7549,N_5963);
or U10725 (N_10725,N_9957,N_9390);
or U10726 (N_10726,N_5988,N_7188);
xor U10727 (N_10727,N_8287,N_8245);
nand U10728 (N_10728,N_7675,N_6671);
nor U10729 (N_10729,N_8038,N_8584);
or U10730 (N_10730,N_7691,N_9542);
nand U10731 (N_10731,N_5662,N_6704);
and U10732 (N_10732,N_7852,N_7872);
nand U10733 (N_10733,N_9289,N_8941);
or U10734 (N_10734,N_8508,N_9162);
nand U10735 (N_10735,N_6778,N_7955);
and U10736 (N_10736,N_5916,N_8167);
nand U10737 (N_10737,N_7213,N_9651);
xor U10738 (N_10738,N_5466,N_5034);
nor U10739 (N_10739,N_5187,N_9338);
nand U10740 (N_10740,N_5850,N_8893);
and U10741 (N_10741,N_7125,N_9918);
or U10742 (N_10742,N_5932,N_6637);
xor U10743 (N_10743,N_6473,N_9554);
nand U10744 (N_10744,N_6242,N_6365);
nand U10745 (N_10745,N_7721,N_5646);
nor U10746 (N_10746,N_7291,N_8081);
nand U10747 (N_10747,N_9362,N_8404);
nor U10748 (N_10748,N_8031,N_7581);
nand U10749 (N_10749,N_5232,N_5482);
nor U10750 (N_10750,N_5706,N_9075);
and U10751 (N_10751,N_9594,N_9932);
or U10752 (N_10752,N_7903,N_8977);
nand U10753 (N_10753,N_7818,N_6548);
nand U10754 (N_10754,N_7590,N_6867);
or U10755 (N_10755,N_6134,N_7767);
xnor U10756 (N_10756,N_8056,N_7242);
nor U10757 (N_10757,N_9674,N_5317);
nor U10758 (N_10758,N_7528,N_6099);
nand U10759 (N_10759,N_7510,N_5700);
xor U10760 (N_10760,N_6580,N_6821);
or U10761 (N_10761,N_7398,N_8432);
nor U10762 (N_10762,N_6317,N_9186);
or U10763 (N_10763,N_8928,N_9068);
xnor U10764 (N_10764,N_5924,N_6239);
or U10765 (N_10765,N_7376,N_9661);
nand U10766 (N_10766,N_7974,N_7461);
and U10767 (N_10767,N_7671,N_6879);
nand U10768 (N_10768,N_7193,N_6036);
nand U10769 (N_10769,N_9923,N_7047);
nand U10770 (N_10770,N_7135,N_8148);
xnor U10771 (N_10771,N_6024,N_6967);
nand U10772 (N_10772,N_6547,N_9492);
xor U10773 (N_10773,N_6417,N_8818);
nor U10774 (N_10774,N_6285,N_9211);
nor U10775 (N_10775,N_6824,N_8654);
nand U10776 (N_10776,N_9697,N_8126);
nor U10777 (N_10777,N_7553,N_5156);
and U10778 (N_10778,N_9122,N_5255);
nand U10779 (N_10779,N_5210,N_6184);
nor U10780 (N_10780,N_9029,N_9707);
nor U10781 (N_10781,N_5122,N_7908);
xor U10782 (N_10782,N_8257,N_9701);
nand U10783 (N_10783,N_7557,N_6760);
xor U10784 (N_10784,N_9507,N_6159);
nand U10785 (N_10785,N_7281,N_5592);
nand U10786 (N_10786,N_8197,N_9003);
xor U10787 (N_10787,N_7045,N_8688);
nor U10788 (N_10788,N_5100,N_5803);
nand U10789 (N_10789,N_6129,N_6610);
or U10790 (N_10790,N_6820,N_7667);
or U10791 (N_10791,N_7832,N_7816);
xor U10792 (N_10792,N_7007,N_8757);
nand U10793 (N_10793,N_7972,N_8415);
or U10794 (N_10794,N_5178,N_6359);
or U10795 (N_10795,N_5990,N_6629);
or U10796 (N_10796,N_7560,N_7240);
or U10797 (N_10797,N_9474,N_5908);
nor U10798 (N_10798,N_5192,N_7343);
or U10799 (N_10799,N_7507,N_5181);
nor U10800 (N_10800,N_5806,N_8373);
nor U10801 (N_10801,N_8002,N_9747);
and U10802 (N_10802,N_9416,N_6059);
nor U10803 (N_10803,N_6933,N_6941);
nand U10804 (N_10804,N_6484,N_8277);
xor U10805 (N_10805,N_7554,N_8088);
xor U10806 (N_10806,N_5776,N_7370);
or U10807 (N_10807,N_7812,N_9989);
nor U10808 (N_10808,N_5500,N_9930);
xnor U10809 (N_10809,N_9877,N_8241);
nand U10810 (N_10810,N_5243,N_8195);
or U10811 (N_10811,N_7268,N_7140);
xor U10812 (N_10812,N_6642,N_7719);
nand U10813 (N_10813,N_6189,N_9271);
and U10814 (N_10814,N_6983,N_6079);
nand U10815 (N_10815,N_7622,N_8076);
nor U10816 (N_10816,N_6483,N_7850);
and U10817 (N_10817,N_6999,N_6250);
and U10818 (N_10818,N_8395,N_6905);
or U10819 (N_10819,N_8991,N_8065);
and U10820 (N_10820,N_5135,N_9461);
nand U10821 (N_10821,N_7229,N_8930);
nand U10822 (N_10822,N_8873,N_5451);
nand U10823 (N_10823,N_6335,N_5911);
nor U10824 (N_10824,N_6897,N_5265);
nand U10825 (N_10825,N_8938,N_5682);
or U10826 (N_10826,N_9742,N_7394);
or U10827 (N_10827,N_9301,N_6556);
and U10828 (N_10828,N_8543,N_6995);
or U10829 (N_10829,N_6828,N_5207);
nand U10830 (N_10830,N_8428,N_6594);
and U10831 (N_10831,N_5490,N_8703);
nand U10832 (N_10832,N_7637,N_9617);
nand U10833 (N_10833,N_7551,N_5273);
and U10834 (N_10834,N_9295,N_6514);
nor U10835 (N_10835,N_8165,N_7630);
nand U10836 (N_10836,N_9402,N_6876);
nor U10837 (N_10837,N_8142,N_7861);
xor U10838 (N_10838,N_8436,N_9663);
nor U10839 (N_10839,N_7215,N_6781);
or U10840 (N_10840,N_6268,N_6330);
or U10841 (N_10841,N_6061,N_8698);
or U10842 (N_10842,N_7346,N_5857);
xnor U10843 (N_10843,N_9190,N_6238);
or U10844 (N_10844,N_8788,N_7964);
and U10845 (N_10845,N_5927,N_6109);
nor U10846 (N_10846,N_5113,N_6376);
nand U10847 (N_10847,N_8868,N_5710);
or U10848 (N_10848,N_6952,N_8597);
or U10849 (N_10849,N_8659,N_9840);
nor U10850 (N_10850,N_6430,N_6742);
and U10851 (N_10851,N_7843,N_5097);
xnor U10852 (N_10852,N_8236,N_8151);
or U10853 (N_10853,N_5564,N_9768);
or U10854 (N_10854,N_8669,N_7512);
nand U10855 (N_10855,N_5947,N_8752);
nor U10856 (N_10856,N_8952,N_7082);
and U10857 (N_10857,N_6471,N_6416);
nor U10858 (N_10858,N_5910,N_7413);
nor U10859 (N_10859,N_9393,N_5571);
or U10860 (N_10860,N_8607,N_5056);
and U10861 (N_10861,N_5221,N_6768);
and U10862 (N_10862,N_9096,N_9857);
and U10863 (N_10863,N_9237,N_9694);
nor U10864 (N_10864,N_6734,N_5881);
or U10865 (N_10865,N_5783,N_6045);
or U10866 (N_10866,N_8107,N_6890);
and U10867 (N_10867,N_5673,N_5443);
nand U10868 (N_10868,N_6352,N_8521);
nor U10869 (N_10869,N_8015,N_8623);
and U10870 (N_10870,N_7919,N_9799);
or U10871 (N_10871,N_5716,N_5721);
xor U10872 (N_10872,N_5866,N_5416);
nand U10873 (N_10873,N_8947,N_6578);
nand U10874 (N_10874,N_9212,N_7405);
xor U10875 (N_10875,N_8333,N_5090);
nand U10876 (N_10876,N_6982,N_5271);
nand U10877 (N_10877,N_5656,N_7166);
nand U10878 (N_10878,N_9825,N_5842);
and U10879 (N_10879,N_7655,N_6135);
xnor U10880 (N_10880,N_8108,N_8269);
nor U10881 (N_10881,N_7453,N_7482);
nand U10882 (N_10882,N_9113,N_6955);
or U10883 (N_10883,N_8787,N_8061);
or U10884 (N_10884,N_8166,N_8754);
nor U10885 (N_10885,N_5758,N_9000);
nor U10886 (N_10886,N_9597,N_6572);
or U10887 (N_10887,N_5867,N_6884);
and U10888 (N_10888,N_8838,N_7070);
xor U10889 (N_10889,N_9911,N_5340);
xor U10890 (N_10890,N_9243,N_7855);
or U10891 (N_10891,N_6719,N_8433);
nand U10892 (N_10892,N_6156,N_6494);
and U10893 (N_10893,N_9247,N_8981);
xor U10894 (N_10894,N_6253,N_9843);
nor U10895 (N_10895,N_7720,N_6797);
or U10896 (N_10896,N_7924,N_9389);
and U10897 (N_10897,N_8186,N_8252);
or U10898 (N_10898,N_9676,N_5382);
and U10899 (N_10899,N_5581,N_6337);
nor U10900 (N_10900,N_5923,N_9297);
or U10901 (N_10901,N_5322,N_6075);
or U10902 (N_10902,N_6012,N_7322);
nor U10903 (N_10903,N_5847,N_8067);
nor U10904 (N_10904,N_6454,N_5948);
xor U10905 (N_10905,N_7033,N_9115);
nor U10906 (N_10906,N_6943,N_7329);
and U10907 (N_10907,N_8129,N_8329);
nand U10908 (N_10908,N_7269,N_8466);
nor U10909 (N_10909,N_8100,N_6800);
nor U10910 (N_10910,N_6662,N_7172);
and U10911 (N_10911,N_6902,N_6643);
xor U10912 (N_10912,N_6868,N_8843);
and U10913 (N_10913,N_7877,N_6550);
xnor U10914 (N_10914,N_5600,N_9929);
nand U10915 (N_10915,N_5093,N_6622);
nor U10916 (N_10916,N_7867,N_7620);
nand U10917 (N_10917,N_9680,N_9600);
xor U10918 (N_10918,N_7210,N_6953);
nor U10919 (N_10919,N_5608,N_9022);
or U10920 (N_10920,N_7494,N_5261);
nor U10921 (N_10921,N_6178,N_9625);
and U10922 (N_10922,N_8813,N_9613);
and U10923 (N_10923,N_8638,N_6435);
and U10924 (N_10924,N_7459,N_9189);
nor U10925 (N_10925,N_5402,N_5760);
nand U10926 (N_10926,N_6971,N_5868);
xor U10927 (N_10927,N_7164,N_9174);
xnor U10928 (N_10928,N_8590,N_8705);
xor U10929 (N_10929,N_5522,N_6711);
nor U10930 (N_10930,N_6534,N_8417);
nor U10931 (N_10931,N_6257,N_9806);
and U10932 (N_10932,N_6300,N_6609);
or U10933 (N_10933,N_9948,N_8431);
nand U10934 (N_10934,N_9072,N_8642);
xnor U10935 (N_10935,N_9936,N_5715);
nand U10936 (N_10936,N_9863,N_8372);
xnor U10937 (N_10937,N_8444,N_5229);
xnor U10938 (N_10938,N_5764,N_7564);
and U10939 (N_10939,N_9916,N_7563);
or U10940 (N_10940,N_7996,N_9255);
nand U10941 (N_10941,N_8118,N_7056);
nand U10942 (N_10942,N_7119,N_6794);
or U10943 (N_10943,N_8177,N_5638);
or U10944 (N_10944,N_5629,N_7830);
and U10945 (N_10945,N_5160,N_6798);
nor U10946 (N_10946,N_9412,N_8556);
nand U10947 (N_10947,N_5258,N_7661);
or U10948 (N_10948,N_9376,N_5711);
xnor U10949 (N_10949,N_9355,N_8769);
xor U10950 (N_10950,N_6731,N_8624);
nand U10951 (N_10951,N_5775,N_7500);
nor U10952 (N_10952,N_5218,N_5759);
xnor U10953 (N_10953,N_9824,N_6723);
nand U10954 (N_10954,N_6283,N_8001);
or U10955 (N_10955,N_5070,N_7538);
nand U10956 (N_10956,N_9283,N_7837);
or U10957 (N_10957,N_8578,N_5452);
or U10958 (N_10958,N_8360,N_5002);
nor U10959 (N_10959,N_8886,N_8362);
or U10960 (N_10960,N_9937,N_8183);
xnor U10961 (N_10961,N_8539,N_9725);
xnor U10962 (N_10962,N_8102,N_8629);
nand U10963 (N_10963,N_6406,N_7426);
nand U10964 (N_10964,N_8214,N_7902);
and U10965 (N_10965,N_7199,N_8987);
nor U10966 (N_10966,N_7991,N_5986);
nand U10967 (N_10967,N_8075,N_5380);
nor U10968 (N_10968,N_5812,N_5285);
and U10969 (N_10969,N_5579,N_8768);
and U10970 (N_10970,N_8940,N_9438);
or U10971 (N_10971,N_8327,N_7513);
xor U10972 (N_10972,N_7131,N_5370);
nor U10973 (N_10973,N_8182,N_6115);
and U10974 (N_10974,N_6830,N_5512);
xor U10975 (N_10975,N_9991,N_5167);
or U10976 (N_10976,N_6456,N_6361);
nor U10977 (N_10977,N_5339,N_7744);
or U10978 (N_10978,N_5305,N_6938);
nand U10979 (N_10979,N_9592,N_8841);
nor U10980 (N_10980,N_5260,N_6918);
and U10981 (N_10981,N_8771,N_9562);
nand U10982 (N_10982,N_7470,N_8567);
nor U10983 (N_10983,N_8528,N_8470);
xor U10984 (N_10984,N_9912,N_7803);
nor U10985 (N_10985,N_5912,N_9809);
and U10986 (N_10986,N_8341,N_7905);
nand U10987 (N_10987,N_9028,N_6961);
and U10988 (N_10988,N_5744,N_8885);
nand U10989 (N_10989,N_8982,N_9529);
and U10990 (N_10990,N_7495,N_7802);
nor U10991 (N_10991,N_7904,N_7733);
or U10992 (N_10992,N_6351,N_6480);
xnor U10993 (N_10993,N_9586,N_6654);
and U10994 (N_10994,N_8811,N_7658);
or U10995 (N_10995,N_6841,N_6236);
xor U10996 (N_10996,N_5875,N_9649);
nor U10997 (N_10997,N_6750,N_5435);
nand U10998 (N_10998,N_9041,N_6198);
xnor U10999 (N_10999,N_8220,N_6718);
or U11000 (N_11000,N_9337,N_6509);
nor U11001 (N_11001,N_5274,N_8345);
or U11002 (N_11002,N_5384,N_6744);
nand U11003 (N_11003,N_6551,N_8335);
and U11004 (N_11004,N_8686,N_6894);
nor U11005 (N_11005,N_8352,N_5228);
nor U11006 (N_11006,N_5904,N_9895);
nor U11007 (N_11007,N_5681,N_7775);
nor U11008 (N_11008,N_8194,N_5829);
or U11009 (N_11009,N_7435,N_5279);
or U11010 (N_11010,N_6697,N_6098);
xnor U11011 (N_11011,N_7443,N_6411);
nor U11012 (N_11012,N_9952,N_7300);
nand U11013 (N_11013,N_7088,N_6772);
or U11014 (N_11014,N_9576,N_8349);
nor U11015 (N_11015,N_7644,N_6521);
and U11016 (N_11016,N_8741,N_8495);
xnor U11017 (N_11017,N_8096,N_7660);
xor U11018 (N_11018,N_8946,N_5695);
nand U11019 (N_11019,N_5389,N_7375);
or U11020 (N_11020,N_8094,N_6167);
and U11021 (N_11021,N_6575,N_9773);
nor U11022 (N_11022,N_8531,N_5650);
or U11023 (N_11023,N_9890,N_7785);
or U11024 (N_11024,N_9221,N_6139);
and U11025 (N_11025,N_8784,N_8229);
nand U11026 (N_11026,N_9220,N_8193);
xnor U11027 (N_11027,N_6998,N_8348);
and U11028 (N_11028,N_8512,N_9238);
or U11029 (N_11029,N_5661,N_9934);
xnor U11030 (N_11030,N_5699,N_7189);
nor U11031 (N_11031,N_7591,N_6398);
and U11032 (N_11032,N_8695,N_8249);
and U11033 (N_11033,N_8558,N_7325);
and U11034 (N_11034,N_6074,N_5799);
xor U11035 (N_11035,N_7571,N_6240);
xor U11036 (N_11036,N_8513,N_6431);
xor U11037 (N_11037,N_6107,N_7336);
or U11038 (N_11038,N_5363,N_5882);
xor U11039 (N_11039,N_7337,N_5861);
nor U11040 (N_11040,N_6119,N_9205);
and U11041 (N_11041,N_6001,N_8820);
or U11042 (N_11042,N_9672,N_9069);
nand U11043 (N_11043,N_6850,N_6453);
or U11044 (N_11044,N_5548,N_6427);
xnor U11045 (N_11045,N_7151,N_8932);
or U11046 (N_11046,N_6951,N_7313);
xnor U11047 (N_11047,N_6974,N_5462);
or U11048 (N_11048,N_7280,N_9261);
and U11049 (N_11049,N_5670,N_8202);
xnor U11050 (N_11050,N_8666,N_9502);
and U11051 (N_11051,N_7884,N_7786);
nand U11052 (N_11052,N_5880,N_8364);
and U11053 (N_11053,N_8231,N_9308);
and U11054 (N_11054,N_9017,N_5696);
xor U11055 (N_11055,N_9164,N_5194);
xor U11056 (N_11056,N_5689,N_8486);
nor U11057 (N_11057,N_6653,N_6929);
or U11058 (N_11058,N_9046,N_8248);
xnor U11059 (N_11059,N_9347,N_6980);
or U11060 (N_11060,N_6457,N_8817);
nand U11061 (N_11061,N_6505,N_9330);
xnor U11062 (N_11062,N_6163,N_5483);
nand U11063 (N_11063,N_7633,N_5371);
or U11064 (N_11064,N_8326,N_7692);
nor U11065 (N_11065,N_8019,N_5035);
and U11066 (N_11066,N_8883,N_7178);
xnor U11067 (N_11067,N_5892,N_7701);
nand U11068 (N_11068,N_9567,N_9481);
and U11069 (N_11069,N_7094,N_7400);
and U11070 (N_11070,N_7795,N_7161);
nand U11071 (N_11071,N_7319,N_5640);
nand U11072 (N_11072,N_8706,N_7249);
or U11073 (N_11073,N_8933,N_6124);
or U11074 (N_11074,N_5492,N_6603);
or U11075 (N_11075,N_5504,N_9407);
or U11076 (N_11076,N_9432,N_8427);
xor U11077 (N_11077,N_5172,N_9971);
xnor U11078 (N_11078,N_6403,N_9128);
xor U11079 (N_11079,N_9931,N_6762);
or U11080 (N_11080,N_7298,N_6327);
and U11081 (N_11081,N_5765,N_8238);
nand U11082 (N_11082,N_7778,N_9662);
xnor U11083 (N_11083,N_5843,N_9206);
xor U11084 (N_11084,N_5570,N_8574);
and U11085 (N_11085,N_8261,N_5598);
xor U11086 (N_11086,N_9515,N_6600);
nand U11087 (N_11087,N_5121,N_6881);
xor U11088 (N_11088,N_9322,N_7819);
xnor U11089 (N_11089,N_8516,N_7674);
nand U11090 (N_11090,N_6870,N_5844);
xnor U11091 (N_11091,N_7586,N_9392);
and U11092 (N_11092,N_5568,N_8753);
xnor U11093 (N_11093,N_8909,N_5531);
or U11094 (N_11094,N_8544,N_7228);
nand U11095 (N_11095,N_7638,N_9214);
xnor U11096 (N_11096,N_6332,N_6623);
nor U11097 (N_11097,N_6927,N_8401);
and U11098 (N_11098,N_5567,N_8258);
xor U11099 (N_11099,N_5651,N_8645);
nand U11100 (N_11100,N_5164,N_9959);
and U11101 (N_11101,N_6157,N_6996);
and U11102 (N_11102,N_5174,N_6789);
or U11103 (N_11103,N_5373,N_9089);
and U11104 (N_11104,N_6793,N_9575);
or U11105 (N_11105,N_9405,N_8583);
nand U11106 (N_11106,N_8898,N_9359);
or U11107 (N_11107,N_9385,N_5914);
nor U11108 (N_11108,N_6345,N_9654);
or U11109 (N_11109,N_6859,N_8085);
and U11110 (N_11110,N_6289,N_7087);
nand U11111 (N_11111,N_8717,N_8605);
nor U11112 (N_11112,N_7030,N_9466);
nor U11113 (N_11113,N_6727,N_5838);
nor U11114 (N_11114,N_8901,N_6576);
nand U11115 (N_11115,N_8224,N_6787);
nor U11116 (N_11116,N_9540,N_6758);
and U11117 (N_11117,N_5660,N_7035);
or U11118 (N_11118,N_7220,N_7254);
and U11119 (N_11119,N_9383,N_9557);
nor U11120 (N_11120,N_8222,N_6899);
xnor U11121 (N_11121,N_7636,N_9910);
nor U11122 (N_11122,N_5493,N_7042);
nor U11123 (N_11123,N_5701,N_5021);
nand U11124 (N_11124,N_6179,N_9354);
xor U11125 (N_11125,N_6546,N_6215);
and U11126 (N_11126,N_5374,N_6073);
or U11127 (N_11127,N_7814,N_6251);
or U11128 (N_11128,N_8732,N_6921);
nor U11129 (N_11129,N_6527,N_5352);
and U11130 (N_11130,N_9023,N_8931);
and U11131 (N_11131,N_6270,N_7144);
or U11132 (N_11132,N_9087,N_6040);
and U11133 (N_11133,N_9960,N_7427);
nor U11134 (N_11134,N_8701,N_7442);
or U11135 (N_11135,N_8683,N_6838);
nand U11136 (N_11136,N_8481,N_5372);
nor U11137 (N_11137,N_8581,N_6776);
or U11138 (N_11138,N_5781,N_5128);
nand U11139 (N_11139,N_6940,N_8131);
xnor U11140 (N_11140,N_6018,N_5015);
nor U11141 (N_11141,N_5772,N_8234);
and U11142 (N_11142,N_5718,N_9537);
and U11143 (N_11143,N_9855,N_6825);
nand U11144 (N_11144,N_8783,N_9437);
nand U11145 (N_11145,N_6755,N_5040);
or U11146 (N_11146,N_5392,N_8028);
and U11147 (N_11147,N_5439,N_8777);
xnor U11148 (N_11148,N_5431,N_9078);
nor U11149 (N_11149,N_9941,N_5326);
nor U11150 (N_11150,N_9630,N_7666);
xnor U11151 (N_11151,N_5396,N_7579);
and U11152 (N_11152,N_8561,N_8748);
xor U11153 (N_11153,N_7659,N_8858);
nor U11154 (N_11154,N_9410,N_6990);
xnor U11155 (N_11155,N_8035,N_9473);
xnor U11156 (N_11156,N_7417,N_8211);
nor U11157 (N_11157,N_9459,N_9439);
nor U11158 (N_11158,N_9328,N_7722);
nor U11159 (N_11159,N_8399,N_7569);
and U11160 (N_11160,N_8730,N_6478);
nand U11161 (N_11161,N_5154,N_6510);
or U11162 (N_11162,N_9252,N_5740);
xor U11163 (N_11163,N_9132,N_7357);
nand U11164 (N_11164,N_9077,N_9692);
nor U11165 (N_11165,N_5336,N_5246);
nand U11166 (N_11166,N_8378,N_5003);
or U11167 (N_11167,N_6621,N_5620);
nand U11168 (N_11168,N_8690,N_9058);
or U11169 (N_11169,N_5905,N_7527);
xnor U11170 (N_11170,N_6488,N_5547);
nor U11171 (N_11171,N_7043,N_8839);
nor U11172 (N_11172,N_7709,N_6309);
xor U11173 (N_11173,N_5872,N_6836);
nor U11174 (N_11174,N_9015,N_9559);
nor U11175 (N_11175,N_9879,N_5199);
and U11176 (N_11176,N_6511,N_9225);
or U11177 (N_11177,N_6218,N_6326);
nand U11178 (N_11178,N_9401,N_6861);
nor U11179 (N_11179,N_8687,N_7012);
nor U11180 (N_11180,N_8312,N_9677);
nand U11181 (N_11181,N_5527,N_7221);
or U11182 (N_11182,N_6703,N_7626);
nor U11183 (N_11183,N_5347,N_7794);
or U11184 (N_11184,N_6089,N_6263);
or U11185 (N_11185,N_5609,N_6338);
xor U11186 (N_11186,N_9643,N_7698);
nand U11187 (N_11187,N_7748,N_8461);
or U11188 (N_11188,N_6598,N_9288);
or U11189 (N_11189,N_7686,N_5683);
nor U11190 (N_11190,N_5935,N_6854);
nor U11191 (N_11191,N_6019,N_7664);
nor U11192 (N_11192,N_6589,N_8397);
xor U11193 (N_11193,N_7612,N_7732);
nor U11194 (N_11194,N_8658,N_5728);
nand U11195 (N_11195,N_7311,N_6810);
or U11196 (N_11196,N_6034,N_9463);
and U11197 (N_11197,N_5165,N_6221);
xnor U11198 (N_11198,N_6557,N_5211);
and U11199 (N_11199,N_8124,N_8144);
and U11200 (N_11200,N_5163,N_5922);
nor U11201 (N_11201,N_5593,N_6466);
nand U11202 (N_11202,N_8039,N_6181);
xnor U11203 (N_11203,N_6989,N_5107);
nor U11204 (N_11204,N_5645,N_5259);
or U11205 (N_11205,N_7362,N_6008);
and U11206 (N_11206,N_5420,N_8589);
nand U11207 (N_11207,N_9703,N_8596);
xor U11208 (N_11208,N_9827,N_5807);
nor U11209 (N_11209,N_6400,N_8204);
or U11210 (N_11210,N_5534,N_8964);
xor U11211 (N_11211,N_8366,N_8828);
or U11212 (N_11212,N_6114,N_9781);
nor U11213 (N_11213,N_7753,N_6764);
nor U11214 (N_11214,N_6194,N_6219);
nor U11215 (N_11215,N_7895,N_6877);
or U11216 (N_11216,N_8861,N_8707);
or U11217 (N_11217,N_8057,N_5049);
nand U11218 (N_11218,N_7576,N_6657);
and U11219 (N_11219,N_9973,N_6146);
or U11220 (N_11220,N_7756,N_5197);
xor U11221 (N_11221,N_9882,N_5999);
or U11222 (N_11222,N_6010,N_8689);
nor U11223 (N_11223,N_7718,N_8737);
xnor U11224 (N_11224,N_7572,N_5955);
nor U11225 (N_11225,N_5752,N_8744);
nor U11226 (N_11226,N_8888,N_7401);
and U11227 (N_11227,N_6969,N_8130);
and U11228 (N_11228,N_9382,N_8260);
or U11229 (N_11229,N_9310,N_5020);
nand U11230 (N_11230,N_7100,N_7714);
or U11231 (N_11231,N_8117,N_9178);
nand U11232 (N_11232,N_9014,N_8656);
and U11233 (N_11233,N_9209,N_5393);
nor U11234 (N_11234,N_5444,N_7606);
xnor U11235 (N_11235,N_9025,N_9539);
xor U11236 (N_11236,N_6049,N_6429);
and U11237 (N_11237,N_8347,N_5205);
xor U11238 (N_11238,N_6028,N_7892);
nor U11239 (N_11239,N_6379,N_7663);
xnor U11240 (N_11240,N_6745,N_8157);
and U11241 (N_11241,N_6408,N_6081);
or U11242 (N_11242,N_5994,N_9269);
and U11243 (N_11243,N_8855,N_6851);
nor U11244 (N_11244,N_5332,N_6567);
and U11245 (N_11245,N_6935,N_7580);
nor U11246 (N_11246,N_9714,N_6807);
xor U11247 (N_11247,N_9517,N_8164);
nor U11248 (N_11248,N_9856,N_8894);
xnor U11249 (N_11249,N_5132,N_6591);
and U11250 (N_11250,N_5479,N_8502);
nand U11251 (N_11251,N_8718,N_8463);
nor U11252 (N_11252,N_5052,N_5708);
and U11253 (N_11253,N_5887,N_6648);
and U11254 (N_11254,N_7537,N_5290);
nand U11255 (N_11255,N_6222,N_8998);
nand U11256 (N_11256,N_7248,N_5862);
xnor U11257 (N_11257,N_9350,N_6197);
xor U11258 (N_11258,N_8990,N_5335);
xor U11259 (N_11259,N_7838,N_8863);
nor U11260 (N_11260,N_8208,N_7117);
and U11261 (N_11261,N_5634,N_9086);
or U11262 (N_11262,N_7509,N_5907);
xor U11263 (N_11263,N_9368,N_7025);
nand U11264 (N_11264,N_8080,N_9870);
nand U11265 (N_11265,N_8280,N_6042);
nor U11266 (N_11266,N_8494,N_5865);
and U11267 (N_11267,N_8315,N_9458);
nor U11268 (N_11268,N_7771,N_9548);
xnor U11269 (N_11269,N_6612,N_8550);
and U11270 (N_11270,N_7001,N_5536);
xnor U11271 (N_11271,N_8313,N_9607);
xor U11272 (N_11272,N_8564,N_5414);
nand U11273 (N_11273,N_6185,N_7174);
xor U11274 (N_11274,N_6617,N_9156);
nor U11275 (N_11275,N_8256,N_7990);
nor U11276 (N_11276,N_9179,N_7360);
nor U11277 (N_11277,N_8764,N_5702);
and U11278 (N_11278,N_5777,N_8153);
xor U11279 (N_11279,N_6726,N_5626);
and U11280 (N_11280,N_6628,N_9054);
nand U11281 (N_11281,N_8198,N_8927);
nor U11282 (N_11282,N_6364,N_8158);
nor U11283 (N_11283,N_7983,N_5603);
and U11284 (N_11284,N_9324,N_9699);
or U11285 (N_11285,N_5110,N_8419);
or U11286 (N_11286,N_9302,N_7085);
nand U11287 (N_11287,N_7212,N_6347);
xnor U11288 (N_11288,N_7502,N_9760);
nor U11289 (N_11289,N_9435,N_6670);
and U11290 (N_11290,N_5191,N_9188);
nand U11291 (N_11291,N_6275,N_9832);
and U11292 (N_11292,N_7717,N_6770);
or U11293 (N_11293,N_9260,N_5559);
nor U11294 (N_11294,N_7341,N_5913);
nand U11295 (N_11295,N_5467,N_9408);
xnor U11296 (N_11296,N_8024,N_8850);
xor U11297 (N_11297,N_6909,N_9307);
nor U11298 (N_11298,N_8956,N_9266);
or U11299 (N_11299,N_9163,N_5653);
or U11300 (N_11300,N_6080,N_6097);
nor U11301 (N_11301,N_9279,N_5436);
or U11302 (N_11302,N_5528,N_7190);
or U11303 (N_11303,N_9745,N_7741);
or U11304 (N_11304,N_5510,N_5111);
xor U11305 (N_11305,N_8936,N_5179);
nor U11306 (N_11306,N_6418,N_9284);
xor U11307 (N_11307,N_8851,N_6321);
nor U11308 (N_11308,N_5562,N_6858);
and U11309 (N_11309,N_7713,N_7372);
or U11310 (N_11310,N_8123,N_8134);
and U11311 (N_11311,N_7243,N_5858);
nor U11312 (N_11312,N_9896,N_6029);
or U11313 (N_11313,N_8694,N_8860);
xnor U11314 (N_11314,N_9789,N_5412);
and U11315 (N_11315,N_6143,N_5476);
nor U11316 (N_11316,N_5321,N_8235);
nor U11317 (N_11317,N_9655,N_9013);
and U11318 (N_11318,N_6272,N_8602);
nand U11319 (N_11319,N_5611,N_6261);
nor U11320 (N_11320,N_8915,N_9092);
xor U11321 (N_11321,N_5499,N_9634);
or U11322 (N_11322,N_6554,N_5944);
nand U11323 (N_11323,N_6893,N_5856);
nor U11324 (N_11324,N_5280,N_8456);
nor U11325 (N_11325,N_7433,N_6495);
xor U11326 (N_11326,N_9161,N_5619);
nand U11327 (N_11327,N_8009,N_7217);
and U11328 (N_11328,N_8242,N_5048);
or U11329 (N_11329,N_9500,N_6164);
nand U11330 (N_11330,N_5463,N_8643);
nand U11331 (N_11331,N_9253,N_6515);
and U11332 (N_11332,N_6064,N_8983);
or U11333 (N_11333,N_6039,N_8289);
nand U11334 (N_11334,N_9706,N_9194);
nand U11335 (N_11335,N_8114,N_7958);
xor U11336 (N_11336,N_5541,N_6803);
or U11337 (N_11337,N_5516,N_7309);
and U11338 (N_11338,N_5552,N_6659);
and U11339 (N_11339,N_5605,N_8441);
nand U11340 (N_11340,N_9528,N_5802);
and U11341 (N_11341,N_6707,N_7829);
or U11342 (N_11342,N_6312,N_9647);
and U11343 (N_11343,N_7925,N_7168);
nor U11344 (N_11344,N_6319,N_8253);
xor U11345 (N_11345,N_8286,N_5449);
nand U11346 (N_11346,N_8145,N_6206);
xor U11347 (N_11347,N_5713,N_6245);
xnor U11348 (N_11348,N_9052,N_9888);
and U11349 (N_11349,N_7169,N_8565);
or U11350 (N_11350,N_6699,N_5784);
and U11351 (N_11351,N_5425,N_7708);
nor U11352 (N_11352,N_6053,N_7727);
xor U11353 (N_11353,N_6385,N_5429);
and U11354 (N_11354,N_7520,N_5242);
nand U11355 (N_11355,N_6475,N_7525);
nor U11356 (N_11356,N_8961,N_7052);
nor U11357 (N_11357,N_8178,N_5622);
nor U11358 (N_11358,N_8159,N_9722);
and U11359 (N_11359,N_5216,N_8807);
nand U11360 (N_11360,N_7652,N_8637);
nor U11361 (N_11361,N_8667,N_9055);
or U11362 (N_11362,N_9138,N_8560);
and U11363 (N_11363,N_7261,N_6149);
and U11364 (N_11364,N_7206,N_7318);
nor U11365 (N_11365,N_9640,N_7506);
or U11366 (N_11366,N_9498,N_9133);
xor U11367 (N_11367,N_8773,N_6391);
nand U11368 (N_11368,N_6280,N_6805);
xnor U11369 (N_11369,N_6968,N_5796);
nand U11370 (N_11370,N_6784,N_6630);
xnor U11371 (N_11371,N_9336,N_8301);
xor U11372 (N_11372,N_9602,N_7327);
or U11373 (N_11373,N_9504,N_5360);
nor U11374 (N_11374,N_8758,N_8674);
and U11375 (N_11375,N_5666,N_7010);
nand U11376 (N_11376,N_9066,N_7543);
and U11377 (N_11377,N_7868,N_8547);
and U11378 (N_11378,N_6038,N_7694);
xnor U11379 (N_11379,N_9659,N_7726);
and U11380 (N_11380,N_9081,N_5859);
nor U11381 (N_11381,N_9743,N_6241);
or U11382 (N_11382,N_6860,N_7641);
xor U11383 (N_11383,N_5088,N_6833);
nor U11384 (N_11384,N_9793,N_9196);
nor U11385 (N_11385,N_7332,N_5460);
xor U11386 (N_11386,N_6003,N_7931);
or U11387 (N_11387,N_7377,N_5974);
xor U11388 (N_11388,N_7444,N_9691);
and U11389 (N_11389,N_6170,N_8649);
nor U11390 (N_11390,N_6224,N_9170);
or U11391 (N_11391,N_9593,N_6023);
xor U11392 (N_11392,N_7369,N_9446);
and U11393 (N_11393,N_6469,N_6244);
and U11394 (N_11394,N_6853,N_9853);
or U11395 (N_11395,N_5746,N_8554);
and U11396 (N_11396,N_7406,N_9906);
and U11397 (N_11397,N_6686,N_9987);
nand U11398 (N_11398,N_8408,N_6700);
nand U11399 (N_11399,N_8980,N_9732);
nand U11400 (N_11400,N_7781,N_8992);
and U11401 (N_11401,N_5408,N_5369);
nor U11402 (N_11402,N_9785,N_6688);
and U11403 (N_11403,N_9245,N_6644);
or U11404 (N_11404,N_5518,N_8973);
nor U11405 (N_11405,N_7822,N_8943);
and U11406 (N_11406,N_5315,N_5676);
or U11407 (N_11407,N_8203,N_9614);
and U11408 (N_11408,N_5879,N_8736);
or U11409 (N_11409,N_6016,N_5140);
nor U11410 (N_11410,N_6501,N_6362);
nand U11411 (N_11411,N_8905,N_9865);
and U11412 (N_11412,N_6656,N_5991);
nand U11413 (N_11413,N_6127,N_5778);
xnor U11414 (N_11414,N_5589,N_5659);
or U11415 (N_11415,N_5501,N_9901);
and U11416 (N_11416,N_8328,N_7128);
xor U11417 (N_11417,N_8538,N_8505);
nand U11418 (N_11418,N_7123,N_5404);
nand U11419 (N_11419,N_8772,N_5119);
xor U11420 (N_11420,N_8380,N_9804);
nand U11421 (N_11421,N_6021,N_6284);
nand U11422 (N_11422,N_6072,N_6310);
nand U11423 (N_11423,N_7736,N_8187);
xnor U11424 (N_11424,N_9508,N_9746);
and U11425 (N_11425,N_9137,N_8368);
nor U11426 (N_11426,N_8790,N_6988);
xor U11427 (N_11427,N_8749,N_6796);
or U11428 (N_11428,N_8288,N_6769);
and U11429 (N_11429,N_9173,N_8804);
nand U11430 (N_11430,N_9494,N_7516);
and U11431 (N_11431,N_6423,N_7621);
nor U11432 (N_11432,N_6009,N_7766);
and U11433 (N_11433,N_6752,N_8154);
and U11434 (N_11434,N_6333,N_9204);
nor U11435 (N_11435,N_9810,N_5649);
and U11436 (N_11436,N_7883,N_7805);
and U11437 (N_11437,N_7699,N_9201);
or U11438 (N_11438,N_6626,N_9010);
xor U11439 (N_11439,N_5432,N_8762);
or U11440 (N_11440,N_8112,N_5966);
or U11441 (N_11441,N_8994,N_7162);
or U11442 (N_11442,N_7619,N_9108);
xor U11443 (N_11443,N_6137,N_6966);
or U11444 (N_11444,N_9845,N_5148);
or U11445 (N_11445,N_9555,N_9358);
nor U11446 (N_11446,N_5826,N_7746);
nor U11447 (N_11447,N_9183,N_8032);
xnor U11448 (N_11448,N_7282,N_8485);
nor U11449 (N_11449,N_6078,N_8021);
or U11450 (N_11450,N_5997,N_7864);
or U11451 (N_11451,N_7881,N_8237);
xnor U11452 (N_11452,N_6676,N_7584);
nor U11453 (N_11453,N_7739,N_6638);
nand U11454 (N_11454,N_6570,N_6992);
or U11455 (N_11455,N_9050,N_9277);
nand U11456 (N_11456,N_9998,N_5430);
and U11457 (N_11457,N_6606,N_6499);
nor U11458 (N_11458,N_9018,N_8330);
xor U11459 (N_11459,N_8986,N_7825);
xnor U11460 (N_11460,N_6738,N_9158);
or U11461 (N_11461,N_5250,N_6538);
nand U11462 (N_11462,N_5461,N_8306);
nand U11463 (N_11463,N_8618,N_5686);
nor U11464 (N_11464,N_9083,N_5022);
xor U11465 (N_11465,N_7334,N_8087);
nor U11466 (N_11466,N_7064,N_9770);
nor U11467 (N_11467,N_6492,N_7534);
and U11468 (N_11468,N_7081,N_9417);
xor U11469 (N_11469,N_8434,N_9142);
and U11470 (N_11470,N_5544,N_6067);
nand U11471 (N_11471,N_7992,N_8665);
or U11472 (N_11472,N_7486,N_5505);
and U11473 (N_11473,N_5299,N_5630);
and U11474 (N_11474,N_5834,N_8344);
xnor U11475 (N_11475,N_7885,N_5241);
or U11476 (N_11476,N_9866,N_9811);
xor U11477 (N_11477,N_5089,N_9195);
nand U11478 (N_11478,N_8641,N_6474);
xor U11479 (N_11479,N_8934,N_8972);
and U11480 (N_11480,N_6026,N_8606);
or U11481 (N_11481,N_6843,N_8506);
nand U11482 (N_11482,N_9397,N_7848);
nor U11483 (N_11483,N_9933,N_9254);
nor U11484 (N_11484,N_7951,N_8580);
or U11485 (N_11485,N_7845,N_7050);
and U11486 (N_11486,N_9248,N_5602);
nor U11487 (N_11487,N_5318,N_6712);
nand U11488 (N_11488,N_6811,N_5958);
nand U11489 (N_11489,N_8227,N_5320);
and U11490 (N_11490,N_7218,N_5230);
xnor U11491 (N_11491,N_6847,N_6973);
xnor U11492 (N_11492,N_8814,N_6399);
nand U11493 (N_11493,N_6318,N_5530);
or U11494 (N_11494,N_9002,N_6553);
and U11495 (N_11495,N_6340,N_9566);
nand U11496 (N_11496,N_7891,N_8351);
xor U11497 (N_11497,N_8478,N_6316);
or U11498 (N_11498,N_5804,N_9997);
nor U11499 (N_11499,N_7008,N_7006);
nand U11500 (N_11500,N_6705,N_8023);
nor U11501 (N_11501,N_5601,N_8484);
xnor U11502 (N_11502,N_6217,N_7185);
nand U11503 (N_11503,N_6959,N_6507);
nor U11504 (N_11504,N_9094,N_7760);
xnor U11505 (N_11505,N_5538,N_7957);
and U11506 (N_11506,N_9033,N_5720);
nor U11507 (N_11507,N_6468,N_7451);
xnor U11508 (N_11508,N_7312,N_5698);
nor U11509 (N_11509,N_8827,N_9883);
and U11510 (N_11510,N_9369,N_7932);
nand U11511 (N_11511,N_9579,N_7715);
or U11512 (N_11512,N_8731,N_5200);
xnor U11513 (N_11513,N_7863,N_9547);
nor U11514 (N_11514,N_7799,N_8526);
xnor U11515 (N_11515,N_7856,N_7706);
xnor U11516 (N_11516,N_7927,N_9975);
and U11517 (N_11517,N_5514,N_5269);
and U11518 (N_11518,N_8840,N_5471);
xor U11519 (N_11519,N_9306,N_9409);
xor U11520 (N_11520,N_7742,N_7834);
or U11521 (N_11521,N_9352,N_9398);
and U11522 (N_11522,N_9199,N_5217);
and U11523 (N_11523,N_6633,N_7807);
xnor U11524 (N_11524,N_7523,N_6728);
nand U11525 (N_11525,N_8720,N_6452);
xnor U11526 (N_11526,N_5276,N_7285);
xor U11527 (N_11527,N_7772,N_6389);
xnor U11528 (N_11528,N_5395,N_8099);
or U11529 (N_11529,N_7728,N_5433);
and U11530 (N_11530,N_6446,N_9887);
or U11531 (N_11531,N_7750,N_5153);
xnor U11532 (N_11532,N_9378,N_7328);
and U11533 (N_11533,N_5573,N_6320);
nor U11534 (N_11534,N_6849,N_6812);
or U11535 (N_11535,N_8511,N_8409);
and U11536 (N_11536,N_5967,N_7643);
and U11537 (N_11537,N_7456,N_5087);
xor U11538 (N_11538,N_8011,N_7365);
or U11539 (N_11539,N_7758,N_7918);
and U11540 (N_11540,N_6667,N_9134);
xor U11541 (N_11541,N_6848,N_9774);
nor U11542 (N_11542,N_5000,N_6180);
or U11543 (N_11543,N_7202,N_7574);
and U11544 (N_11544,N_5836,N_7299);
xor U11545 (N_11545,N_9981,N_8877);
xnor U11546 (N_11546,N_6237,N_9526);
or U11547 (N_11547,N_9963,N_8660);
or U11548 (N_11548,N_6641,N_5125);
and U11549 (N_11549,N_6533,N_5350);
or U11550 (N_11550,N_5428,N_7294);
nand U11551 (N_11551,N_5818,N_8598);
xor U11552 (N_11552,N_8054,N_7526);
nor U11553 (N_11553,N_7508,N_5797);
nor U11554 (N_11554,N_6903,N_6518);
xnor U11555 (N_11555,N_8169,N_7389);
and U11556 (N_11556,N_7392,N_7745);
xnor U11557 (N_11557,N_8437,N_5943);
or U11558 (N_11558,N_7121,N_5238);
xor U11559 (N_11559,N_7361,N_8902);
nand U11560 (N_11560,N_6118,N_7342);
nor U11561 (N_11561,N_6102,N_8728);
and U11562 (N_11562,N_8651,N_8290);
xor U11563 (N_11563,N_8180,N_5086);
and U11564 (N_11564,N_9091,N_9532);
nand U11565 (N_11565,N_9230,N_5484);
nor U11566 (N_11566,N_5346,N_7054);
nor U11567 (N_11567,N_5223,N_8267);
nand U11568 (N_11568,N_7546,N_5354);
nand U11569 (N_11569,N_7404,N_9543);
xnor U11570 (N_11570,N_9363,N_5809);
xor U11571 (N_11571,N_5771,N_9281);
and U11572 (N_11572,N_5201,N_9051);
nor U11573 (N_11573,N_9893,N_9333);
and U11574 (N_11574,N_5509,N_6857);
xor U11575 (N_11575,N_5800,N_5957);
and U11576 (N_11576,N_9379,N_8546);
nor U11577 (N_11577,N_6649,N_6108);
xnor U11578 (N_11578,N_5468,N_8939);
xnor U11579 (N_11579,N_5085,N_8585);
nor U11580 (N_11580,N_7514,N_8537);
and U11581 (N_11581,N_9187,N_7134);
or U11582 (N_11582,N_9273,N_9583);
xnor U11583 (N_11583,N_8044,N_7645);
xor U11584 (N_11584,N_8697,N_6920);
or U11585 (N_11585,N_9079,N_9847);
or U11586 (N_11586,N_5282,N_9064);
and U11587 (N_11587,N_6566,N_9505);
nor U11588 (N_11588,N_5753,N_9043);
or U11589 (N_11589,N_9193,N_9531);
xor U11590 (N_11590,N_6775,N_6449);
nor U11591 (N_11591,N_8304,N_8375);
nand U11592 (N_11592,N_7120,N_9326);
nand U11593 (N_11593,N_5739,N_7734);
nand U11594 (N_11594,N_9008,N_7157);
or U11595 (N_11595,N_6126,N_5903);
nor U11596 (N_11596,N_8896,N_9457);
nor U11597 (N_11597,N_5001,N_8899);
nor U11598 (N_11598,N_7363,N_9112);
nor U11599 (N_11599,N_6569,N_7276);
nand U11600 (N_11600,N_9653,N_8420);
and U11601 (N_11601,N_6908,N_9585);
or U11602 (N_11602,N_7065,N_6926);
or U11603 (N_11603,N_7295,N_5047);
and U11604 (N_11604,N_9240,N_6878);
xor U11605 (N_11605,N_5170,N_9657);
and U11606 (N_11606,N_8318,N_5674);
nor U11607 (N_11607,N_7899,N_7529);
nor U11608 (N_11608,N_9228,N_6158);
and U11609 (N_11609,N_6369,N_5762);
xnor U11610 (N_11610,N_7491,N_8058);
nor U11611 (N_11611,N_7263,N_6844);
xnor U11612 (N_11612,N_7963,N_5061);
nor U11613 (N_11613,N_8406,N_6255);
and U11614 (N_11614,N_8480,N_9104);
and U11615 (N_11615,N_7763,N_6205);
and U11616 (N_11616,N_6433,N_5542);
nor U11617 (N_11617,N_9367,N_9922);
nor U11618 (N_11618,N_8746,N_9323);
or U11619 (N_11619,N_7614,N_8239);
nor U11620 (N_11620,N_9805,N_7251);
and U11621 (N_11621,N_9329,N_8824);
and U11622 (N_11622,N_8738,N_9424);
or U11623 (N_11623,N_9769,N_8575);
xnor U11624 (N_11624,N_8949,N_5995);
and U11625 (N_11625,N_5690,N_5642);
and U11626 (N_11626,N_5030,N_8751);
or U11627 (N_11627,N_9472,N_8323);
or U11628 (N_11628,N_8859,N_8975);
and U11629 (N_11629,N_7875,N_9823);
xnor U11630 (N_11630,N_9315,N_7871);
or U11631 (N_11631,N_6891,N_8906);
and U11632 (N_11632,N_8137,N_5677);
nor U11633 (N_11633,N_5572,N_7177);
nor U11634 (N_11634,N_8808,N_7634);
and U11635 (N_11635,N_7835,N_8761);
or U11636 (N_11636,N_5036,N_8358);
and U11637 (N_11637,N_9478,N_6862);
nand U11638 (N_11638,N_5851,N_6315);
and U11639 (N_11639,N_8393,N_8219);
xnor U11640 (N_11640,N_9678,N_5596);
and U11641 (N_11641,N_6112,N_9482);
and U11642 (N_11642,N_8525,N_8000);
and U11643 (N_11643,N_9564,N_9450);
nor U11644 (N_11644,N_6765,N_7460);
and U11645 (N_11645,N_7350,N_6782);
and U11646 (N_11646,N_7851,N_9715);
nor U11647 (N_11647,N_5485,N_5104);
or U11648 (N_11648,N_7487,N_7934);
nand U11649 (N_11649,N_7194,N_7380);
or U11650 (N_11650,N_7900,N_8722);
xnor U11651 (N_11651,N_6802,N_7391);
and U11652 (N_11652,N_8325,N_8795);
nand U11653 (N_11653,N_8549,N_8876);
xor U11654 (N_11654,N_7689,N_7555);
nor U11655 (N_11655,N_7386,N_9124);
nand U11656 (N_11656,N_9095,N_6187);
xnor U11657 (N_11657,N_6286,N_7307);
xnor U11658 (N_11658,N_6620,N_8379);
xnor U11659 (N_11659,N_9848,N_8012);
or U11660 (N_11660,N_5403,N_7544);
or U11661 (N_11661,N_9690,N_5768);
and U11662 (N_11662,N_6209,N_5878);
or U11663 (N_11663,N_9360,N_8533);
or U11664 (N_11664,N_7051,N_5405);
and U11665 (N_11665,N_8639,N_8175);
xnor U11666 (N_11666,N_9704,N_8155);
and U11667 (N_11667,N_9231,N_7978);
xnor U11668 (N_11668,N_9790,N_7310);
nand U11669 (N_11669,N_7238,N_7640);
nor U11670 (N_11670,N_9842,N_9603);
and U11671 (N_11671,N_9039,N_9965);
xor U11672 (N_11672,N_8217,N_5329);
or U11673 (N_11673,N_7789,N_6795);
xnor U11674 (N_11674,N_7129,N_9496);
xor U11675 (N_11675,N_8865,N_6481);
or U11676 (N_11676,N_5227,N_8522);
nor U11677 (N_11677,N_5846,N_8573);
and U11678 (N_11678,N_8619,N_9103);
nor U11679 (N_11679,N_6733,N_6766);
xnor U11680 (N_11680,N_7935,N_9818);
or U11681 (N_11681,N_9406,N_7731);
nand U11682 (N_11682,N_5811,N_5091);
nand U11683 (N_11683,N_8499,N_5780);
and U11684 (N_11684,N_6070,N_6055);
nor U11685 (N_11685,N_6582,N_8053);
or U11686 (N_11686,N_6930,N_5268);
nand U11687 (N_11687,N_5134,N_7260);
nand U11688 (N_11688,N_6267,N_5193);
and U11689 (N_11689,N_5309,N_9153);
xnor U11690 (N_11690,N_8755,N_8356);
and U11691 (N_11691,N_9421,N_6945);
nand U11692 (N_11692,N_8247,N_5915);
xor U11693 (N_11693,N_6972,N_6710);
and U11694 (N_11694,N_9031,N_6169);
xor U11695 (N_11695,N_6962,N_7779);
nor U11696 (N_11696,N_9477,N_8265);
xnor U11697 (N_11697,N_6984,N_7639);
nand U11698 (N_11698,N_9258,N_6465);
nand U11699 (N_11699,N_9717,N_9497);
or U11700 (N_11700,N_6249,N_9730);
or U11701 (N_11701,N_7075,N_8493);
and U11702 (N_11702,N_6138,N_5928);
and U11703 (N_11703,N_6274,N_6162);
or U11704 (N_11704,N_7147,N_6645);
nor U11705 (N_11705,N_6722,N_9545);
xnor U11706 (N_11706,N_9915,N_9780);
xnor U11707 (N_11707,N_9817,N_7015);
and U11708 (N_11708,N_8120,N_6761);
and U11709 (N_11709,N_5415,N_7583);
nand U11710 (N_11710,N_5139,N_7252);
xnor U11711 (N_11711,N_6303,N_5876);
nand U11712 (N_11712,N_6225,N_5719);
nor U11713 (N_11713,N_5841,N_7101);
xor U11714 (N_11714,N_7044,N_9667);
nor U11715 (N_11715,N_7191,N_5612);
or U11716 (N_11716,N_9348,N_7609);
and U11717 (N_11717,N_6922,N_6305);
nand U11718 (N_11718,N_8518,N_8903);
and U11719 (N_11719,N_9905,N_5364);
xnor U11720 (N_11720,N_8475,N_6373);
or U11721 (N_11721,N_7788,N_8147);
nand U11722 (N_11722,N_9518,N_8770);
and U11723 (N_11723,N_9182,N_8918);
nor U11724 (N_11724,N_9881,N_8951);
nand U11725 (N_11725,N_8369,N_8199);
nor U11726 (N_11726,N_8837,N_7876);
nor U11727 (N_11727,N_8047,N_6865);
nor U11728 (N_11728,N_7962,N_9668);
nor U11729 (N_11729,N_9117,N_6584);
or U11730 (N_11730,N_8520,N_7824);
nor U11731 (N_11731,N_7493,N_8592);
xor U11732 (N_11732,N_8563,N_8416);
nand U11733 (N_11733,N_9514,N_5833);
nand U11734 (N_11734,N_7898,N_9126);
and U11735 (N_11735,N_8760,N_7700);
nand U11736 (N_11736,N_9988,N_6976);
xor U11737 (N_11737,N_7163,N_9423);
nand U11738 (N_11738,N_9468,N_8767);
nor U11739 (N_11739,N_5930,N_9001);
nand U11740 (N_11740,N_7474,N_9154);
nand U11741 (N_11741,N_9191,N_9610);
nand U11742 (N_11742,N_7003,N_8995);
nand U11743 (N_11743,N_9454,N_9891);
xnor U11744 (N_11744,N_9996,N_8309);
xnor U11745 (N_11745,N_6104,N_7841);
and U11746 (N_11746,N_9444,N_8086);
or U11747 (N_11747,N_9993,N_9783);
nor U11748 (N_11748,N_9485,N_6017);
and U11749 (N_11749,N_5464,N_6763);
and U11750 (N_11750,N_6739,N_9151);
xor U11751 (N_11751,N_8907,N_5798);
or U11752 (N_11752,N_7737,N_7941);
nor U11753 (N_11753,N_7179,N_8527);
and U11754 (N_11754,N_8810,N_5108);
nor U11755 (N_11755,N_6647,N_8612);
and U11756 (N_11756,N_9938,N_7160);
nand U11757 (N_11757,N_9861,N_8476);
nand U11758 (N_11758,N_9057,N_9445);
and U11759 (N_11759,N_8776,N_9414);
and U11760 (N_11760,N_8962,N_6311);
xor U11761 (N_11761,N_7481,N_9686);
and U11762 (N_11762,N_7945,N_6916);
nor U11763 (N_11763,N_5669,N_8653);
nor U11764 (N_11764,N_8887,N_5507);
or U11765 (N_11765,N_9534,N_7097);
and U11766 (N_11766,N_7171,N_9521);
nor U11767 (N_11767,N_8097,N_9222);
and U11768 (N_11768,N_9265,N_5576);
nand U11769 (N_11769,N_6880,N_6160);
nor U11770 (N_11770,N_9236,N_8548);
and U11771 (N_11771,N_9850,N_6151);
or U11772 (N_11772,N_9580,N_8160);
nor U11773 (N_11773,N_5511,N_9660);
or U11774 (N_11774,N_7831,N_8613);
nand U11775 (N_11775,N_7098,N_6392);
nor U11776 (N_11776,N_9939,N_7136);
nor U11777 (N_11777,N_9346,N_8881);
or U11778 (N_11778,N_6852,N_7952);
or U11779 (N_11779,N_7650,N_9786);
nand U11780 (N_11780,N_5143,N_8355);
or U11781 (N_11781,N_9777,N_7595);
nor U11782 (N_11782,N_7897,N_5933);
and U11783 (N_11783,N_8968,N_9740);
or U11784 (N_11784,N_9833,N_9312);
nor U11785 (N_11785,N_5334,N_8693);
nor U11786 (N_11786,N_8677,N_8443);
nand U11787 (N_11787,N_5688,N_5704);
nand U11788 (N_11788,N_5146,N_9388);
and U11789 (N_11789,N_7473,N_5808);
nor U11790 (N_11790,N_5830,N_7143);
and U11791 (N_11791,N_7093,N_7201);
or U11792 (N_11792,N_9071,N_7673);
nand U11793 (N_11793,N_6663,N_7467);
or U11794 (N_11794,N_9452,N_6874);
or U11795 (N_11795,N_9867,N_6624);
xnor U11796 (N_11796,N_7687,N_6302);
nand U11797 (N_11797,N_6147,N_8016);
xnor U11798 (N_11798,N_7522,N_6223);
xnor U11799 (N_11799,N_7690,N_9772);
xor U11800 (N_11800,N_9411,N_7156);
nand U11801 (N_11801,N_8988,N_5105);
nand U11802 (N_11802,N_7192,N_7597);
or U11803 (N_11803,N_9816,N_8276);
nor U11804 (N_11804,N_5212,N_5054);
nand U11805 (N_11805,N_9325,N_5331);
nand U11806 (N_11806,N_9604,N_5277);
and U11807 (N_11807,N_5017,N_8848);
nor U11808 (N_11808,N_6027,N_5736);
xnor U11809 (N_11809,N_6907,N_7836);
nand U11810 (N_11810,N_5072,N_6054);
and U11811 (N_11811,N_5394,N_5325);
xnor U11812 (N_11812,N_5041,N_6493);
nand U11813 (N_11813,N_6050,N_5147);
xnor U11814 (N_11814,N_9200,N_8271);
and U11815 (N_11815,N_5018,N_9256);
and U11816 (N_11816,N_9460,N_9637);
nor U11817 (N_11817,N_6426,N_6592);
and U11818 (N_11818,N_5679,N_6422);
and U11819 (N_11819,N_6827,N_8336);
and U11820 (N_11820,N_7197,N_8228);
nand U11821 (N_11821,N_7078,N_7632);
nor U11822 (N_11822,N_9056,N_5585);
xnor U11823 (N_11823,N_8213,N_7804);
nand U11824 (N_11824,N_7103,N_5419);
and U11825 (N_11825,N_6046,N_6652);
or U11826 (N_11826,N_6144,N_5445);
or U11827 (N_11827,N_5064,N_7948);
nor U11828 (N_11828,N_6111,N_8282);
or U11829 (N_11829,N_9105,N_7302);
nor U11830 (N_11830,N_9656,N_8579);
nor U11831 (N_11831,N_7354,N_6808);
and U11832 (N_11832,N_7517,N_7879);
xnor U11833 (N_11833,N_7533,N_6444);
nor U11834 (N_11834,N_5065,N_7594);
xor U11835 (N_11835,N_5597,N_9754);
nor U11836 (N_11836,N_6066,N_9483);
or U11837 (N_11837,N_9513,N_9299);
nor U11838 (N_11838,N_7485,N_7475);
nand U11839 (N_11839,N_7792,N_9716);
and U11840 (N_11840,N_5453,N_8106);
nand U11841 (N_11841,N_9082,N_6460);
nor U11842 (N_11842,N_9449,N_5617);
xor U11843 (N_11843,N_9908,N_8924);
nand U11844 (N_11844,N_7148,N_7440);
xor U11845 (N_11845,N_6030,N_8657);
nor U11846 (N_11846,N_7600,N_9181);
nand U11847 (N_11847,N_6271,N_7827);
xor U11848 (N_11848,N_5333,N_7235);
nand U11849 (N_11849,N_7225,N_8796);
xor U11850 (N_11850,N_8529,N_8923);
and U11851 (N_11851,N_9849,N_6691);
and U11852 (N_11852,N_7458,N_6724);
nand U11853 (N_11853,N_9320,N_9475);
and U11854 (N_11854,N_7685,N_7716);
xor U11855 (N_11855,N_7613,N_9088);
nor U11856 (N_11856,N_5920,N_8310);
xnor U11857 (N_11857,N_8171,N_7823);
nor U11858 (N_11858,N_8490,N_5118);
and U11859 (N_11859,N_8240,N_5025);
nor U11860 (N_11860,N_9642,N_5042);
or U11861 (N_11861,N_5607,N_8403);
xnor U11862 (N_11862,N_8074,N_6528);
nand U11863 (N_11863,N_6954,N_6788);
or U11864 (N_11864,N_9763,N_9970);
nor U11865 (N_11865,N_6082,N_6809);
nor U11866 (N_11866,N_9020,N_6387);
or U11867 (N_11867,N_8105,N_5328);
and U11868 (N_11868,N_6370,N_8343);
and U11869 (N_11869,N_8819,N_5732);
xor U11870 (N_11870,N_5747,N_9361);
or U11871 (N_11871,N_8908,N_8937);
nand U11872 (N_11872,N_5046,N_8407);
and U11873 (N_11873,N_7678,N_8176);
nor U11874 (N_11874,N_6944,N_7418);
xnor U11875 (N_11875,N_8866,N_9838);
or U11876 (N_11876,N_9180,N_5871);
nor U11877 (N_11877,N_9192,N_9293);
xor U11878 (N_11878,N_8852,N_5016);
and U11879 (N_11879,N_7233,N_5984);
and U11880 (N_11880,N_6559,N_7080);
and U11881 (N_11881,N_7472,N_6771);
xor U11882 (N_11882,N_5311,N_6193);
and U11883 (N_11883,N_5029,N_8644);
nand U11884 (N_11884,N_8451,N_7800);
nor U11885 (N_11885,N_5032,N_6434);
nand U11886 (N_11886,N_6937,N_9821);
and U11887 (N_11887,N_7628,N_5909);
nor U11888 (N_11888,N_5668,N_9074);
or U11889 (N_11889,N_9904,N_8185);
or U11890 (N_11890,N_6051,N_6103);
nor U11891 (N_11891,N_9720,N_6183);
nand U11892 (N_11892,N_9924,N_9968);
xor U11893 (N_11893,N_8571,N_5545);
nor U11894 (N_11894,N_7981,N_6587);
nor U11895 (N_11895,N_8139,N_9294);
xor U11896 (N_11896,N_7979,N_7729);
nand U11897 (N_11897,N_6839,N_7757);
xor U11898 (N_11898,N_5980,N_6684);
nand U11899 (N_11899,N_9434,N_8844);
or U11900 (N_11900,N_7095,N_7940);
or U11901 (N_11901,N_7797,N_8882);
xor U11902 (N_11902,N_6914,N_5491);
and U11903 (N_11903,N_9943,N_7999);
and U11904 (N_11904,N_8460,N_8331);
or U11905 (N_11905,N_6997,N_5951);
and U11906 (N_11906,N_6068,N_8846);
nor U11907 (N_11907,N_8740,N_9524);
xor U11908 (N_11908,N_9007,N_8889);
xor U11909 (N_11909,N_9004,N_5011);
xor U11910 (N_11910,N_7916,N_7542);
and U11911 (N_11911,N_5789,N_5832);
nand U11912 (N_11912,N_9615,N_7227);
and U11913 (N_11913,N_9060,N_7465);
nand U11914 (N_11914,N_7038,N_8230);
xnor U11915 (N_11915,N_8668,N_9978);
xnor U11916 (N_11916,N_5563,N_9956);
nand U11917 (N_11917,N_9862,N_9331);
xor U11918 (N_11918,N_7222,N_7618);
nor U11919 (N_11919,N_8307,N_5756);
nor U11920 (N_11920,N_9101,N_8049);
or U11921 (N_11921,N_9090,N_9748);
nor U11922 (N_11922,N_6092,N_6355);
or U11923 (N_11923,N_6658,N_8942);
xnor U11924 (N_11924,N_7556,N_5817);
or U11925 (N_11925,N_6031,N_7137);
nand U11926 (N_11926,N_8524,N_9232);
nand U11927 (N_11927,N_9489,N_6500);
nor U11928 (N_11928,N_9107,N_5487);
nor U11929 (N_11929,N_5741,N_9076);
nor U11930 (N_11930,N_5983,N_8122);
xor U11931 (N_11931,N_6792,N_9658);
nand U11932 (N_11932,N_6588,N_6130);
nor U11933 (N_11933,N_5934,N_8897);
xnor U11934 (N_11934,N_7688,N_8084);
and U11935 (N_11935,N_9541,N_5889);
nand U11936 (N_11936,N_8914,N_6395);
or U11937 (N_11937,N_8830,N_5434);
and U11938 (N_11938,N_5319,N_5900);
and U11939 (N_11939,N_5979,N_8832);
nand U11940 (N_11940,N_8611,N_8095);
and U11941 (N_11941,N_9544,N_5985);
nor U11942 (N_11942,N_6856,N_7266);
and U11943 (N_11943,N_6531,N_7258);
xnor U11944 (N_11944,N_8190,N_9565);
and U11945 (N_11945,N_5297,N_9909);
nor U11946 (N_11946,N_9202,N_5358);
xnor U11947 (N_11947,N_6467,N_9340);
or U11948 (N_11948,N_6439,N_7911);
nor U11949 (N_11949,N_7740,N_8093);
and U11950 (N_11950,N_8472,N_8904);
xnor U11951 (N_11951,N_6759,N_8976);
and U11952 (N_11952,N_8586,N_7108);
xor U11953 (N_11953,N_6177,N_5540);
and U11954 (N_11954,N_5080,N_9106);
and U11955 (N_11955,N_5477,N_8834);
nand U11956 (N_11956,N_9239,N_5729);
nor U11957 (N_11957,N_5145,N_6970);
nand U11958 (N_11958,N_7662,N_5810);
nor U11959 (N_11959,N_9639,N_5737);
or U11960 (N_11960,N_9042,N_7000);
and U11961 (N_11961,N_7055,N_9121);
and U11962 (N_11962,N_8091,N_9167);
nand U11963 (N_11963,N_7649,N_6917);
xor U11964 (N_11964,N_7109,N_5901);
or U11965 (N_11965,N_7953,N_6281);
xnor U11966 (N_11966,N_6729,N_5624);
nand U11967 (N_11967,N_9983,N_6447);
and U11968 (N_11968,N_8756,N_5884);
nor U11969 (N_11969,N_7130,N_8386);
nor U11970 (N_11970,N_7041,N_8880);
or U11971 (N_11971,N_9085,N_7980);
nand U11972 (N_11972,N_5343,N_9828);
nor U11973 (N_11973,N_5058,N_8268);
nand U11974 (N_11974,N_8671,N_5902);
xnor U11975 (N_11975,N_7457,N_8008);
xor U11976 (N_11976,N_8945,N_8367);
nor U11977 (N_11977,N_5822,N_7106);
nor U11978 (N_11978,N_7384,N_7601);
xnor U11979 (N_11979,N_6835,N_5521);
or U11980 (N_11980,N_8042,N_5888);
and U11981 (N_11981,N_7854,N_6491);
xor U11982 (N_11982,N_6462,N_9752);
nor U11983 (N_11983,N_7414,N_6128);
nand U11984 (N_11984,N_6295,N_7821);
and U11985 (N_11985,N_8559,N_7118);
nand U11986 (N_11986,N_8950,N_8912);
nand U11987 (N_11987,N_7463,N_8133);
nor U11988 (N_11988,N_9820,N_8616);
nand U11989 (N_11989,N_7005,N_8957);
and U11990 (N_11990,N_8966,N_6141);
xnor U11991 (N_11991,N_7264,N_5565);
nor U11992 (N_11992,N_7521,N_9860);
and U11993 (N_11993,N_9125,N_7441);
and U11994 (N_11994,N_8210,N_5112);
nor U11995 (N_11995,N_6394,N_5956);
nand U11996 (N_11996,N_8283,N_9925);
nand U11997 (N_11997,N_8633,N_6599);
xor U11998 (N_11998,N_7598,N_9387);
or U11999 (N_11999,N_9344,N_6840);
nor U12000 (N_12000,N_6590,N_5950);
xor U12001 (N_12001,N_5438,N_6925);
nand U12002 (N_12002,N_6294,N_7449);
nand U12003 (N_12003,N_5076,N_9958);
nand U12004 (N_12004,N_5657,N_7145);
and U12005 (N_12005,N_7198,N_5743);
nor U12006 (N_12006,N_7808,N_7677);
nor U12007 (N_12007,N_7559,N_9357);
nand U12008 (N_12008,N_9084,N_6191);
and U12009 (N_12009,N_5582,N_6846);
and U12010 (N_12010,N_5583,N_6823);
nor U12011 (N_12011,N_5349,N_9858);
nand U12012 (N_12012,N_7149,N_9099);
nand U12013 (N_12013,N_6497,N_5520);
and U12014 (N_12014,N_7566,N_7617);
nand U12015 (N_12015,N_5009,N_7208);
nor U12016 (N_12016,N_8072,N_8285);
nor U12017 (N_12017,N_9286,N_8316);
xor U12018 (N_12018,N_7286,N_9724);
or U12019 (N_12019,N_7844,N_9027);
nand U12020 (N_12020,N_9342,N_9588);
or U12021 (N_12021,N_9572,N_8048);
nor U12022 (N_12022,N_9097,N_7274);
xor U12023 (N_12023,N_9750,N_5864);
nor U12024 (N_12024,N_6015,N_7596);
nor U12025 (N_12025,N_9160,N_8078);
and U12026 (N_12026,N_8387,N_6757);
nor U12027 (N_12027,N_9523,N_9700);
or U12028 (N_12028,N_8631,N_9589);
or U12029 (N_12029,N_9143,N_7665);
and U12030 (N_12030,N_9184,N_7105);
and U12031 (N_12031,N_9123,N_9263);
or U12032 (N_12032,N_7445,N_5066);
or U12033 (N_12033,N_5355,N_6912);
xnor U12034 (N_12034,N_6069,N_7378);
nand U12035 (N_12035,N_9569,N_6872);
and U12036 (N_12036,N_5323,N_6348);
nand U12037 (N_12037,N_5996,N_7338);
or U12038 (N_12038,N_8791,N_9431);
and U12039 (N_12039,N_8429,N_7524);
nand U12040 (N_12040,N_9633,N_7651);
and U12041 (N_12041,N_5486,N_8298);
xnor U12042 (N_12042,N_6906,N_9907);
and U12043 (N_12043,N_8856,N_9894);
xor U12044 (N_12044,N_7464,N_8869);
nor U12045 (N_12045,N_9427,N_9693);
and U12046 (N_12046,N_8119,N_7759);
nor U12047 (N_12047,N_5976,N_5063);
or U12048 (N_12048,N_9605,N_5291);
nor U12049 (N_12049,N_8483,N_9147);
and U12050 (N_12050,N_6516,N_6441);
and U12051 (N_12051,N_9224,N_7452);
and U12052 (N_12052,N_6577,N_6672);
or U12053 (N_12053,N_8101,N_5182);
nor U12054 (N_12054,N_8374,N_9244);
or U12055 (N_12055,N_7535,N_5535);
or U12056 (N_12056,N_6168,N_9259);
nor U12057 (N_12057,N_7702,N_8496);
and U12058 (N_12058,N_8712,N_9749);
nor U12059 (N_12059,N_9626,N_8913);
xnor U12060 (N_12060,N_8780,N_6573);
and U12061 (N_12061,N_9442,N_8262);
nor U12062 (N_12062,N_9275,N_7253);
and U12063 (N_12063,N_7390,N_5694);
nor U12064 (N_12064,N_9219,N_9159);
nand U12065 (N_12065,N_6819,N_7477);
xnor U12066 (N_12066,N_8711,N_5556);
xor U12067 (N_12067,N_7568,N_6165);
and U12068 (N_12068,N_6767,N_9399);
xnor U12069 (N_12069,N_6522,N_6161);
and U12070 (N_12070,N_5840,N_5213);
or U12071 (N_12071,N_7423,N_6965);
or U12072 (N_12072,N_7518,N_7724);
xnor U12073 (N_12073,N_8218,N_6668);
xor U12074 (N_12074,N_5770,N_5978);
or U12075 (N_12075,N_7462,N_6679);
nand U12076 (N_12076,N_6732,N_7730);
or U12077 (N_12077,N_7762,N_7914);
xnor U12078 (N_12078,N_5316,N_6740);
and U12079 (N_12079,N_9977,N_7430);
nor U12080 (N_12080,N_5886,N_8089);
xnor U12081 (N_12081,N_6246,N_8255);
or U12082 (N_12082,N_5921,N_6085);
nand U12083 (N_12083,N_5204,N_6323);
nor U12084 (N_12084,N_6888,N_6814);
nand U12085 (N_12085,N_5353,N_9131);
nand U12086 (N_12086,N_6673,N_5379);
nand U12087 (N_12087,N_5595,N_6747);
xnor U12088 (N_12088,N_5057,N_5195);
nor U12089 (N_12089,N_6512,N_8482);
nand U12090 (N_12090,N_8849,N_5423);
nor U12091 (N_12091,N_6716,N_6227);
nand U12092 (N_12092,N_6304,N_9629);
nor U12093 (N_12093,N_5918,N_8206);
or U12094 (N_12094,N_6887,N_6414);
xnor U12095 (N_12095,N_8721,N_8503);
or U12096 (N_12096,N_7349,N_6105);
xor U12097 (N_12097,N_5793,N_9808);
xnor U12098 (N_12098,N_7113,N_6405);
nor U12099 (N_12099,N_5157,N_5240);
or U12100 (N_12100,N_9871,N_6062);
xnor U12101 (N_12101,N_9920,N_7468);
nand U12102 (N_12102,N_8430,N_9550);
or U12103 (N_12103,N_8279,N_5234);
or U12104 (N_12104,N_9739,N_7176);
and U12105 (N_12105,N_9636,N_7154);
nor U12106 (N_12106,N_7099,N_7028);
and U12107 (N_12107,N_5424,N_8610);
nand U12108 (N_12108,N_5390,N_9712);
and U12109 (N_12109,N_7880,N_6175);
and U12110 (N_12110,N_7489,N_6565);
xnor U12111 (N_12111,N_9698,N_5615);
or U12112 (N_12112,N_7498,N_9152);
or U12113 (N_12113,N_8925,N_7575);
xor U12114 (N_12114,N_5726,N_8426);
and U12115 (N_12115,N_7083,N_9484);
xnor U12116 (N_12116,N_6048,N_7115);
nor U12117 (N_12117,N_9172,N_9510);
and U12118 (N_12118,N_9731,N_9755);
xnor U12119 (N_12119,N_8884,N_7014);
nand U12120 (N_12120,N_5375,N_7167);
or U12121 (N_12121,N_9800,N_5254);
nand U12122 (N_12122,N_8890,N_8045);
or U12123 (N_12123,N_9560,N_5873);
or U12124 (N_12124,N_8647,N_9030);
nand U12125 (N_12125,N_6254,N_6397);
xnor U12126 (N_12126,N_8226,N_9669);
and U12127 (N_12127,N_7289,N_8284);
nand U12128 (N_12128,N_6948,N_8541);
and U12129 (N_12129,N_8110,N_7920);
nor U12130 (N_12130,N_5095,N_6448);
or U12131 (N_12131,N_5965,N_5304);
and U12132 (N_12132,N_8501,N_8170);
nor U12133 (N_12133,N_9309,N_9218);
nand U12134 (N_12134,N_6041,N_7906);
and U12135 (N_12135,N_5639,N_8376);
nand U12136 (N_12136,N_6442,N_9467);
and U12137 (N_12137,N_8727,N_5357);
xor U12138 (N_12138,N_5801,N_5177);
xnor U12139 (N_12139,N_7270,N_7973);
nand U12140 (N_12140,N_9688,N_7381);
or U12141 (N_12141,N_6052,N_8477);
xor U12142 (N_12142,N_7060,N_7428);
nor U12143 (N_12143,N_5094,N_6690);
xor U12144 (N_12144,N_7262,N_8140);
or U12145 (N_12145,N_5488,N_7810);
or U12146 (N_12146,N_6353,N_5303);
xor U12147 (N_12147,N_9679,N_9436);
xor U12148 (N_12148,N_9506,N_5975);
xor U12149 (N_12149,N_8273,N_9767);
xnor U12150 (N_12150,N_9864,N_7317);
or U12151 (N_12151,N_6791,N_9598);
nor U12152 (N_12152,N_7670,N_9945);
and U12153 (N_12153,N_9846,N_6863);
nand U12154 (N_12154,N_9953,N_7223);
and U12155 (N_12155,N_6252,N_6166);
or U12156 (N_12156,N_5821,N_6154);
nand U12157 (N_12157,N_7977,N_9946);
xor U12158 (N_12158,N_5184,N_8535);
or U12159 (N_12159,N_5407,N_7629);
and U12160 (N_12160,N_5114,N_5293);
nor U12161 (N_12161,N_5687,N_7284);
and U12162 (N_12162,N_7669,N_8509);
and U12163 (N_12163,N_5575,N_8090);
and U12164 (N_12164,N_5270,N_5171);
nor U12165 (N_12165,N_8471,N_8792);
xnor U12166 (N_12166,N_8184,N_8617);
nand U12167 (N_12167,N_7497,N_7345);
nor U12168 (N_12168,N_5794,N_5286);
and U12169 (N_12169,N_5855,N_6004);
or U12170 (N_12170,N_8062,N_9641);
and U12171 (N_12171,N_6664,N_7395);
and U12172 (N_12172,N_8793,N_5378);
xnor U12173 (N_12173,N_6374,N_9520);
nor U12174 (N_12174,N_7061,N_6113);
and U12175 (N_12175,N_8999,N_9917);
xor U12176 (N_12176,N_5007,N_5244);
nor U12177 (N_12177,N_5839,N_9648);
xor U12178 (N_12178,N_9665,N_6977);
nor U12179 (N_12179,N_5998,N_8029);
xnor U12180 (N_12180,N_9601,N_7158);
and U12181 (N_12181,N_8207,N_6013);
xor U12182 (N_12182,N_6928,N_8092);
xor U12183 (N_12183,N_9814,N_9443);
nor U12184 (N_12184,N_7219,N_9578);
or U12185 (N_12185,N_5754,N_8875);
nor U12186 (N_12186,N_9073,N_6783);
or U12187 (N_12187,N_5820,N_6450);
nor U12188 (N_12188,N_7926,N_7340);
nor U12189 (N_12189,N_6293,N_7057);
nand U12190 (N_12190,N_5296,N_8970);
and U12191 (N_12191,N_8292,N_6605);
and U12192 (N_12192,N_8007,N_6717);
nor U12193 (N_12193,N_8251,N_6956);
nand U12194 (N_12194,N_6785,N_5073);
nor U12195 (N_12195,N_8519,N_5239);
nand U12196 (N_12196,N_8874,N_8593);
xor U12197 (N_12197,N_7570,N_5557);
nand U12198 (N_12198,N_6911,N_9049);
nor U12199 (N_12199,N_7259,N_6801);
and U12200 (N_12200,N_9675,N_7625);
xnor U12201 (N_12201,N_5150,N_6037);
xor U12202 (N_12202,N_6579,N_7074);
or U12203 (N_12203,N_9792,N_9451);
or U12204 (N_12204,N_8205,N_5877);
nor U12205 (N_12205,N_6296,N_6975);
and U12206 (N_12206,N_7237,N_7301);
nor U12207 (N_12207,N_5788,N_9974);
nand U12208 (N_12208,N_5292,N_7471);
and U12209 (N_12209,N_9796,N_7393);
and U12210 (N_12210,N_9696,N_9233);
nor U12211 (N_12211,N_9034,N_7499);
or U12212 (N_12212,N_5202,N_7344);
xnor U12213 (N_12213,N_8305,N_8334);
xnor U12214 (N_12214,N_8778,N_6088);
xor U12215 (N_12215,N_8551,N_7086);
nand U12216 (N_12216,N_8281,N_6627);
and U12217 (N_12217,N_5972,N_5397);
and U12218 (N_12218,N_7069,N_8149);
nand U12219 (N_12219,N_5968,N_5705);
and U12220 (N_12220,N_5757,N_9495);
or U12221 (N_12221,N_5675,N_7421);
xor U12222 (N_12222,N_6607,N_6524);
or U12223 (N_12223,N_8438,N_5782);
nand U12224 (N_12224,N_7037,N_7484);
nor U12225 (N_12225,N_6140,N_6585);
or U12226 (N_12226,N_5159,N_6404);
and U12227 (N_12227,N_5890,N_7966);
xnor U12228 (N_12228,N_5149,N_5120);
or U12229 (N_12229,N_6420,N_8340);
nor U12230 (N_12230,N_6035,N_5447);
xnor U12231 (N_12231,N_9868,N_8339);
xnor U12232 (N_12232,N_6866,N_7943);
or U12233 (N_12233,N_7250,N_8026);
nand U12234 (N_12234,N_5344,N_5302);
and U12235 (N_12235,N_8921,N_8935);
or U12236 (N_12236,N_7939,N_5684);
and U12237 (N_12237,N_7967,N_8005);
nand U12238 (N_12238,N_5519,N_8314);
and U12239 (N_12239,N_7111,N_5427);
or U12240 (N_12240,N_6325,N_6650);
nand U12241 (N_12241,N_9618,N_5152);
nor U12242 (N_12242,N_9878,N_7432);
and U12243 (N_12243,N_7165,N_9317);
and U12244 (N_12244,N_9913,N_8510);
nor U12245 (N_12245,N_9949,N_8338);
nor U12246 (N_12246,N_9080,N_5294);
nand U12247 (N_12247,N_9365,N_8223);
or U12248 (N_12248,N_8003,N_6133);
nor U12249 (N_12249,N_9278,N_9441);
nor U12250 (N_12250,N_7541,N_7296);
nand U12251 (N_12251,N_6539,N_8614);
xnor U12252 (N_12252,N_5124,N_8663);
nand U12253 (N_12253,N_9552,N_5478);
nand U12254 (N_12254,N_5233,N_8794);
xor U12255 (N_12255,N_5498,N_7226);
or U12256 (N_12256,N_8414,N_5616);
xnor U12257 (N_12257,N_8410,N_6220);
nand U12258 (N_12258,N_7909,N_5033);
and U12259 (N_12259,N_9819,N_6574);
xor U12260 (N_12260,N_9268,N_9666);
nand U12261 (N_12261,N_6336,N_5566);
and U12262 (N_12262,N_9623,N_8704);
nor U12263 (N_12263,N_9141,N_6372);
and U12264 (N_12264,N_5287,N_5247);
nand U12265 (N_12265,N_6247,N_8557);
xnor U12266 (N_12266,N_9144,N_6715);
and U12267 (N_12267,N_6960,N_7995);
xor U12268 (N_12268,N_8459,N_7828);
xnor U12269 (N_12269,N_8955,N_9067);
nor U12270 (N_12270,N_8332,N_9702);
and U12271 (N_12271,N_8109,N_9921);
and U12272 (N_12272,N_8815,N_5092);
nand U12273 (N_12273,N_7353,N_7454);
nand U12274 (N_12274,N_8412,N_8553);
and U12275 (N_12275,N_5618,N_6407);
and U12276 (N_12276,N_7531,N_8168);
nand U12277 (N_12277,N_6375,N_9149);
xnor U12278 (N_12278,N_7039,N_7684);
nor U12279 (N_12279,N_8250,N_6057);
and U12280 (N_12280,N_9053,N_5459);
xor U12281 (N_12281,N_8394,N_8750);
or U12282 (N_12282,N_9876,N_7205);
xor U12283 (N_12283,N_5925,N_6542);
and U12284 (N_12284,N_5964,N_8724);
and U12285 (N_12285,N_8216,N_8765);
xnor U12286 (N_12286,N_5281,N_9711);
nor U12287 (N_12287,N_7416,N_9577);
or U12288 (N_12288,N_8013,N_5588);
xor U12289 (N_12289,N_5815,N_5288);
nor U12290 (N_12290,N_7347,N_5586);
nor U12291 (N_12291,N_6476,N_7438);
nor U12292 (N_12292,N_9788,N_5632);
nor U12293 (N_12293,N_6152,N_5625);
and U12294 (N_12294,N_7209,N_7200);
nor U12295 (N_12295,N_8803,N_7203);
and U12296 (N_12296,N_9246,N_7929);
nor U12297 (N_12297,N_9582,N_8189);
and U12298 (N_12298,N_6233,N_8030);
or U12299 (N_12299,N_6298,N_7588);
and U12300 (N_12300,N_8742,N_7436);
nand U12301 (N_12301,N_6695,N_9127);
xnor U12302 (N_12302,N_5039,N_7984);
nor U12303 (N_12303,N_5792,N_5345);
nand U12304 (N_12304,N_8113,N_9835);
or U12305 (N_12305,N_8555,N_8826);
xor U12306 (N_12306,N_9859,N_5703);
or U12307 (N_12307,N_9897,N_9734);
or U12308 (N_12308,N_9177,N_9869);
nor U12309 (N_12309,N_8802,N_6043);
xor U12310 (N_12310,N_6616,N_9171);
or U12311 (N_12311,N_9826,N_9628);
nand U12312 (N_12312,N_8878,N_5155);
xor U12313 (N_12313,N_6322,N_8636);
nor U12314 (N_12314,N_9169,N_9364);
nand U12315 (N_12315,N_6496,N_7754);
nor U12316 (N_12316,N_8540,N_6790);
xnor U12317 (N_12317,N_9511,N_7944);
nand U12318 (N_12318,N_5208,N_9992);
and U12319 (N_12319,N_5366,N_5275);
and U12320 (N_12320,N_5426,N_9384);
nor U12321 (N_12321,N_6401,N_5062);
xnor U12322 (N_12322,N_9267,N_8458);
nor U12323 (N_12323,N_6540,N_8270);
or U12324 (N_12324,N_5136,N_5138);
xor U12325 (N_12325,N_7068,N_7552);
or U12326 (N_12326,N_7539,N_7765);
nor U12327 (N_12327,N_9940,N_8552);
or U12328 (N_12328,N_9453,N_8311);
or U12329 (N_12329,N_5599,N_5219);
nor U12330 (N_12330,N_7547,N_8172);
xor U12331 (N_12331,N_6949,N_9226);
nand U12332 (N_12332,N_7769,N_9727);
nand U12333 (N_12333,N_6677,N_6214);
nand U12334 (N_12334,N_8300,N_8143);
and U12335 (N_12335,N_9349,N_5680);
nor U12336 (N_12336,N_7305,N_8601);
or U12337 (N_12337,N_7668,N_7408);
xnor U12338 (N_12338,N_5494,N_7331);
nand U12339 (N_12339,N_9433,N_8713);
or U12340 (N_12340,N_9440,N_6845);
nand U12341 (N_12341,N_7059,N_5038);
and U12342 (N_12342,N_5123,N_5937);
and U12343 (N_12343,N_8487,N_7431);
xnor U12344 (N_12344,N_8391,N_5931);
nand U12345 (N_12345,N_9851,N_7410);
and U12346 (N_12346,N_6749,N_8212);
and U12347 (N_12347,N_5480,N_9019);
nand U12348 (N_12348,N_7993,N_9778);
xor U12349 (N_12349,N_9738,N_9377);
and U12350 (N_12350,N_7682,N_7672);
or U12351 (N_12351,N_6086,N_5173);
and U12352 (N_12352,N_9570,N_5561);
or U12353 (N_12353,N_9129,N_7170);
and U12354 (N_12354,N_5267,N_8173);
nand U12355 (N_12355,N_5827,N_5495);
xor U12356 (N_12356,N_8678,N_7040);
nand U12357 (N_12357,N_7938,N_9264);
nand U12358 (N_12358,N_9928,N_5835);
nand U12359 (N_12359,N_6896,N_5779);
xnor U12360 (N_12360,N_9304,N_9525);
nand U12361 (N_12361,N_6508,N_9413);
or U12362 (N_12362,N_8291,N_9241);
xnor U12363 (N_12363,N_6328,N_7847);
nor U12364 (N_12364,N_6837,N_7024);
nor U12365 (N_12365,N_8507,N_6076);
nor U12366 (N_12366,N_6412,N_9761);
nor U12367 (N_12367,N_6946,N_6834);
or U12368 (N_12368,N_6619,N_5019);
or U12369 (N_12369,N_5631,N_6201);
xor U12370 (N_12370,N_9290,N_9947);
or U12371 (N_12371,N_8797,N_7985);
xor U12372 (N_12372,N_7982,N_8278);
nor U12373 (N_12373,N_5055,N_7182);
nor U12374 (N_12374,N_6120,N_5264);
and U12375 (N_12375,N_6002,N_7073);
nor U12376 (N_12376,N_9215,N_9985);
xor U12377 (N_12377,N_8454,N_6095);
or U12378 (N_12378,N_9670,N_6502);
nor U12379 (N_12379,N_6517,N_6635);
nand U12380 (N_12380,N_9753,N_9762);
or U12381 (N_12381,N_9356,N_5224);
or U12382 (N_12382,N_6208,N_9685);
or U12383 (N_12383,N_5658,N_7696);
xnor U12384 (N_12384,N_8104,N_5214);
xnor U12385 (N_12385,N_8447,N_7577);
xor U12386 (N_12386,N_5936,N_7853);
xnor U12387 (N_12387,N_7314,N_9332);
or U12388 (N_12388,N_5766,N_5584);
nor U12389 (N_12389,N_8083,N_6014);
nand U12390 (N_12390,N_9635,N_8266);
and U12391 (N_12391,N_8121,N_6248);
nand U12392 (N_12392,N_7707,N_7356);
nand U12393 (N_12393,N_7857,N_8411);
and U12394 (N_12394,N_8295,N_8710);
and U12395 (N_12395,N_7773,N_7878);
or U12396 (N_12396,N_6228,N_8854);
and U12397 (N_12397,N_9708,N_7801);
nand U12398 (N_12398,N_9621,N_7124);
xnor U12399 (N_12399,N_5383,N_8448);
xor U12400 (N_12400,N_9999,N_7388);
and U12401 (N_12401,N_6445,N_7858);
nand U12402 (N_12402,N_6472,N_9021);
xnor U12403 (N_12403,N_7425,N_5894);
or U12404 (N_12404,N_7257,N_8014);
and U12405 (N_12405,N_7710,N_8132);
nor U12406 (N_12406,N_9587,N_5773);
or U12407 (N_12407,N_5151,N_7653);
and U12408 (N_12408,N_6199,N_7917);
or U12409 (N_12409,N_9797,N_7697);
and U12410 (N_12410,N_5524,N_9612);
and U12411 (N_12411,N_5083,N_7505);
nand U12412 (N_12412,N_9165,N_5082);
nor U12413 (N_12413,N_9942,N_7501);
nor U12414 (N_12414,N_9681,N_8609);
or U12415 (N_12415,N_6424,N_7712);
or U12416 (N_12416,N_7267,N_7053);
and U12417 (N_12417,N_7585,N_9627);
nor U12418 (N_12418,N_5418,N_8576);
nand U12419 (N_12419,N_7241,N_5961);
xor U12420 (N_12420,N_6892,N_9465);
nand U12421 (N_12421,N_8603,N_9854);
and U12422 (N_12422,N_5790,N_8628);
nand U12423 (N_12423,N_6436,N_8383);
nor U12424 (N_12424,N_8418,N_5026);
nor U12425 (N_12425,N_5580,N_9831);
or U12426 (N_12426,N_6432,N_8046);
and U12427 (N_12427,N_7419,N_7657);
nand U12428 (N_12428,N_8627,N_7986);
xnor U12429 (N_12429,N_7071,N_6753);
xor U12430 (N_12430,N_7478,N_7385);
or U12431 (N_12431,N_9880,N_6440);
nand U12432 (N_12432,N_5727,N_5769);
nor U12433 (N_12433,N_7749,N_8063);
or U12434 (N_12434,N_5359,N_8302);
and U12435 (N_12435,N_8068,N_5084);
and U12436 (N_12436,N_9462,N_5059);
nand U12437 (N_12437,N_6693,N_5406);
nor U12438 (N_12438,N_8450,N_7155);
nor U12439 (N_12439,N_5551,N_6200);
or U12440 (N_12440,N_8010,N_7183);
nand U12441 (N_12441,N_7112,N_7930);
nand U12442 (N_12442,N_5284,N_9516);
or U12443 (N_12443,N_5574,N_6991);
xnor U12444 (N_12444,N_6262,N_9216);
or U12445 (N_12445,N_7504,N_8587);
xnor U12446 (N_12446,N_5248,N_9276);
nand U12447 (N_12447,N_5024,N_7027);
nand U12448 (N_12448,N_7915,N_8363);
or U12449 (N_12449,N_9100,N_5249);
and U12450 (N_12450,N_5235,N_7776);
and U12451 (N_12451,N_8682,N_8620);
xor U12452 (N_12452,N_9415,N_7921);
or U12453 (N_12453,N_8530,N_7764);
or U12454 (N_12454,N_8646,N_5709);
or U12455 (N_12455,N_5074,N_9024);
nor U12456 (N_12456,N_8111,N_5362);
nor U12457 (N_12457,N_5310,N_7605);
or U12458 (N_12458,N_7642,N_9533);
or U12459 (N_12459,N_5496,N_7142);
xor U12460 (N_12460,N_5550,N_7330);
and U12461 (N_12461,N_5077,N_7623);
or U12462 (N_12462,N_6675,N_9282);
and U12463 (N_12463,N_9036,N_8422);
xnor U12464 (N_12464,N_7676,N_7910);
nand U12465 (N_12465,N_7076,N_5594);
nand U12466 (N_12466,N_7704,N_5745);
or U12467 (N_12467,N_9319,N_9590);
or U12468 (N_12468,N_7723,N_8322);
nor U12469 (N_12469,N_6443,N_5324);
nor U12470 (N_12470,N_8296,N_7352);
and U12471 (N_12471,N_8766,N_6725);
nand U12472 (N_12472,N_5196,N_7530);
xor U12473 (N_12473,N_7862,N_9146);
and U12474 (N_12474,N_9822,N_5654);
or U12475 (N_12475,N_7607,N_5289);
xor U12476 (N_12476,N_7247,N_7654);
and U12477 (N_12477,N_6947,N_8071);
nor U12478 (N_12478,N_7297,N_8523);
or U12479 (N_12479,N_6188,N_6822);
and U12480 (N_12480,N_6634,N_7379);
xor U12481 (N_12481,N_5314,N_6366);
and U12482 (N_12482,N_9470,N_5869);
nand U12483 (N_12483,N_8264,N_8515);
xnor U12484 (N_12484,N_8568,N_5130);
nor U12485 (N_12485,N_5060,N_8041);
or U12486 (N_12486,N_5814,N_9571);
nand U12487 (N_12487,N_6934,N_8388);
nand U12488 (N_12488,N_5791,N_7104);
nor U12489 (N_12489,N_8699,N_6815);
nor U12490 (N_12490,N_8421,N_6558);
and U12491 (N_12491,N_8479,N_6698);
nand U12492 (N_12492,N_8492,N_9351);
or U12493 (N_12493,N_5569,N_5386);
xor U12494 (N_12494,N_7011,N_9270);
nand U12495 (N_12495,N_6458,N_5503);
and U12496 (N_12496,N_8692,N_5941);
nand U12497 (N_12497,N_8670,N_7960);
nor U12498 (N_12498,N_9791,N_7695);
nand U12499 (N_12499,N_8209,N_9116);
nor U12500 (N_12500,N_7473,N_8580);
or U12501 (N_12501,N_5534,N_9368);
xor U12502 (N_12502,N_7524,N_6631);
xnor U12503 (N_12503,N_9467,N_8423);
nand U12504 (N_12504,N_6326,N_5429);
or U12505 (N_12505,N_8090,N_9431);
and U12506 (N_12506,N_5267,N_6734);
and U12507 (N_12507,N_7408,N_6722);
nand U12508 (N_12508,N_7113,N_5368);
or U12509 (N_12509,N_5937,N_9304);
and U12510 (N_12510,N_5067,N_5522);
and U12511 (N_12511,N_9621,N_9415);
or U12512 (N_12512,N_9600,N_5230);
nor U12513 (N_12513,N_9388,N_5490);
or U12514 (N_12514,N_5612,N_6428);
and U12515 (N_12515,N_5426,N_6285);
and U12516 (N_12516,N_8377,N_6831);
or U12517 (N_12517,N_8285,N_5276);
or U12518 (N_12518,N_8846,N_6172);
xor U12519 (N_12519,N_8808,N_6856);
or U12520 (N_12520,N_5950,N_5643);
and U12521 (N_12521,N_7258,N_6886);
and U12522 (N_12522,N_9853,N_8596);
xor U12523 (N_12523,N_7370,N_7906);
or U12524 (N_12524,N_6897,N_6783);
and U12525 (N_12525,N_7741,N_8734);
nand U12526 (N_12526,N_6162,N_9924);
nand U12527 (N_12527,N_6528,N_7159);
or U12528 (N_12528,N_7658,N_8904);
nand U12529 (N_12529,N_9703,N_6512);
or U12530 (N_12530,N_6594,N_5938);
or U12531 (N_12531,N_9167,N_7923);
nand U12532 (N_12532,N_6376,N_5630);
nand U12533 (N_12533,N_5278,N_7368);
nand U12534 (N_12534,N_6321,N_5839);
xor U12535 (N_12535,N_5190,N_8335);
and U12536 (N_12536,N_9907,N_8935);
and U12537 (N_12537,N_6802,N_9381);
and U12538 (N_12538,N_8643,N_5317);
nor U12539 (N_12539,N_6640,N_8135);
nor U12540 (N_12540,N_7521,N_5840);
nand U12541 (N_12541,N_8016,N_6709);
nand U12542 (N_12542,N_9180,N_8999);
and U12543 (N_12543,N_9325,N_5997);
or U12544 (N_12544,N_7713,N_5842);
nand U12545 (N_12545,N_9501,N_6256);
or U12546 (N_12546,N_5451,N_6760);
nor U12547 (N_12547,N_7401,N_9783);
or U12548 (N_12548,N_6271,N_8438);
xor U12549 (N_12549,N_5699,N_6744);
nor U12550 (N_12550,N_8015,N_8934);
xnor U12551 (N_12551,N_6235,N_5131);
nand U12552 (N_12552,N_5035,N_6180);
or U12553 (N_12553,N_7279,N_9117);
nand U12554 (N_12554,N_7656,N_7817);
nor U12555 (N_12555,N_9038,N_7874);
nand U12556 (N_12556,N_8863,N_8550);
and U12557 (N_12557,N_8399,N_8707);
and U12558 (N_12558,N_6476,N_5419);
and U12559 (N_12559,N_9008,N_5826);
xnor U12560 (N_12560,N_7599,N_9111);
and U12561 (N_12561,N_7222,N_7610);
nand U12562 (N_12562,N_7264,N_6627);
or U12563 (N_12563,N_7531,N_5642);
or U12564 (N_12564,N_6016,N_6051);
nand U12565 (N_12565,N_6699,N_5948);
or U12566 (N_12566,N_7549,N_9296);
xnor U12567 (N_12567,N_8226,N_7609);
and U12568 (N_12568,N_9273,N_6292);
nor U12569 (N_12569,N_9782,N_6726);
nor U12570 (N_12570,N_6333,N_8360);
nand U12571 (N_12571,N_7910,N_7886);
and U12572 (N_12572,N_8589,N_5060);
and U12573 (N_12573,N_7738,N_5447);
nand U12574 (N_12574,N_6100,N_6004);
and U12575 (N_12575,N_5796,N_6888);
xor U12576 (N_12576,N_9651,N_5436);
xnor U12577 (N_12577,N_5504,N_9876);
nor U12578 (N_12578,N_6515,N_9082);
xnor U12579 (N_12579,N_8552,N_7948);
xor U12580 (N_12580,N_5357,N_8289);
and U12581 (N_12581,N_7025,N_5511);
and U12582 (N_12582,N_5274,N_5044);
xor U12583 (N_12583,N_9661,N_6235);
and U12584 (N_12584,N_7995,N_7304);
xor U12585 (N_12585,N_5800,N_9671);
nand U12586 (N_12586,N_7589,N_8209);
nor U12587 (N_12587,N_7766,N_7490);
or U12588 (N_12588,N_7574,N_8782);
and U12589 (N_12589,N_7504,N_9313);
xor U12590 (N_12590,N_5042,N_5079);
nand U12591 (N_12591,N_9952,N_9731);
xor U12592 (N_12592,N_6400,N_8254);
xor U12593 (N_12593,N_7891,N_5411);
nand U12594 (N_12594,N_5975,N_9667);
or U12595 (N_12595,N_5687,N_6745);
xor U12596 (N_12596,N_6034,N_6932);
nand U12597 (N_12597,N_9590,N_6329);
xor U12598 (N_12598,N_5935,N_5509);
and U12599 (N_12599,N_6262,N_5553);
and U12600 (N_12600,N_6490,N_8290);
xnor U12601 (N_12601,N_6516,N_8186);
xnor U12602 (N_12602,N_5227,N_8732);
or U12603 (N_12603,N_8906,N_8107);
nor U12604 (N_12604,N_5479,N_9068);
xnor U12605 (N_12605,N_7206,N_6283);
or U12606 (N_12606,N_6723,N_5815);
and U12607 (N_12607,N_6062,N_6698);
nand U12608 (N_12608,N_9416,N_6979);
or U12609 (N_12609,N_7695,N_6917);
nor U12610 (N_12610,N_6532,N_8903);
nor U12611 (N_12611,N_9342,N_9785);
nor U12612 (N_12612,N_7221,N_8586);
nand U12613 (N_12613,N_9610,N_8308);
nand U12614 (N_12614,N_6991,N_9015);
xnor U12615 (N_12615,N_5203,N_8669);
or U12616 (N_12616,N_6757,N_7723);
and U12617 (N_12617,N_5843,N_8838);
and U12618 (N_12618,N_6695,N_6611);
nand U12619 (N_12619,N_8433,N_8520);
xnor U12620 (N_12620,N_8924,N_7212);
and U12621 (N_12621,N_6479,N_8048);
nor U12622 (N_12622,N_9688,N_6086);
nor U12623 (N_12623,N_9517,N_6457);
nor U12624 (N_12624,N_5151,N_5814);
and U12625 (N_12625,N_5759,N_8868);
xnor U12626 (N_12626,N_7828,N_8914);
or U12627 (N_12627,N_9818,N_5718);
or U12628 (N_12628,N_5069,N_9210);
nand U12629 (N_12629,N_9490,N_5087);
nor U12630 (N_12630,N_9727,N_6066);
and U12631 (N_12631,N_9996,N_9928);
or U12632 (N_12632,N_6827,N_8268);
and U12633 (N_12633,N_6134,N_8524);
nand U12634 (N_12634,N_6582,N_8071);
nand U12635 (N_12635,N_6475,N_5995);
nand U12636 (N_12636,N_8205,N_7772);
nand U12637 (N_12637,N_9521,N_9843);
xor U12638 (N_12638,N_5884,N_9441);
or U12639 (N_12639,N_8681,N_8455);
nor U12640 (N_12640,N_5786,N_6462);
and U12641 (N_12641,N_5355,N_8278);
or U12642 (N_12642,N_9587,N_6679);
nor U12643 (N_12643,N_5142,N_8136);
or U12644 (N_12644,N_9171,N_8600);
nand U12645 (N_12645,N_7721,N_5467);
and U12646 (N_12646,N_6849,N_8549);
and U12647 (N_12647,N_9412,N_8372);
and U12648 (N_12648,N_7827,N_8081);
nand U12649 (N_12649,N_8533,N_8311);
nand U12650 (N_12650,N_8739,N_8654);
nor U12651 (N_12651,N_8790,N_8045);
nor U12652 (N_12652,N_5048,N_8215);
nor U12653 (N_12653,N_8973,N_8941);
nor U12654 (N_12654,N_5728,N_7985);
nand U12655 (N_12655,N_6881,N_7635);
and U12656 (N_12656,N_8789,N_9882);
nor U12657 (N_12657,N_9317,N_9682);
and U12658 (N_12658,N_7174,N_6518);
nor U12659 (N_12659,N_9402,N_7952);
xor U12660 (N_12660,N_9225,N_8365);
nor U12661 (N_12661,N_7940,N_9123);
xor U12662 (N_12662,N_9887,N_6977);
nor U12663 (N_12663,N_7301,N_6843);
nand U12664 (N_12664,N_7781,N_5632);
and U12665 (N_12665,N_5718,N_5350);
and U12666 (N_12666,N_5800,N_5484);
xor U12667 (N_12667,N_8426,N_9143);
and U12668 (N_12668,N_5211,N_6107);
and U12669 (N_12669,N_5853,N_5705);
nor U12670 (N_12670,N_7732,N_8128);
nor U12671 (N_12671,N_9721,N_8816);
or U12672 (N_12672,N_7645,N_6570);
xor U12673 (N_12673,N_9933,N_9961);
nor U12674 (N_12674,N_8495,N_6470);
nor U12675 (N_12675,N_9724,N_5016);
xnor U12676 (N_12676,N_6973,N_7569);
or U12677 (N_12677,N_8131,N_8518);
nand U12678 (N_12678,N_6835,N_9393);
nand U12679 (N_12679,N_8893,N_5606);
nor U12680 (N_12680,N_9524,N_7251);
nor U12681 (N_12681,N_8582,N_9678);
nor U12682 (N_12682,N_9063,N_7123);
nand U12683 (N_12683,N_6330,N_5998);
nand U12684 (N_12684,N_8182,N_8581);
nor U12685 (N_12685,N_7001,N_8426);
and U12686 (N_12686,N_7412,N_6382);
or U12687 (N_12687,N_7109,N_9887);
or U12688 (N_12688,N_6375,N_5538);
nor U12689 (N_12689,N_5688,N_5217);
or U12690 (N_12690,N_5229,N_5376);
nand U12691 (N_12691,N_5387,N_6367);
xor U12692 (N_12692,N_9298,N_9586);
and U12693 (N_12693,N_8895,N_5713);
xor U12694 (N_12694,N_6981,N_7503);
xnor U12695 (N_12695,N_8663,N_6953);
and U12696 (N_12696,N_5361,N_8297);
xor U12697 (N_12697,N_9411,N_7869);
xor U12698 (N_12698,N_6736,N_7727);
nand U12699 (N_12699,N_7564,N_8119);
or U12700 (N_12700,N_8224,N_7615);
and U12701 (N_12701,N_9439,N_9727);
nor U12702 (N_12702,N_8243,N_5192);
nand U12703 (N_12703,N_8547,N_6169);
nand U12704 (N_12704,N_6765,N_8035);
or U12705 (N_12705,N_9476,N_9037);
and U12706 (N_12706,N_5008,N_8328);
and U12707 (N_12707,N_5247,N_7403);
xnor U12708 (N_12708,N_7025,N_9405);
and U12709 (N_12709,N_9294,N_9651);
nand U12710 (N_12710,N_5848,N_9142);
or U12711 (N_12711,N_8307,N_9700);
nand U12712 (N_12712,N_8042,N_8940);
or U12713 (N_12713,N_8806,N_6929);
nor U12714 (N_12714,N_9022,N_5307);
nand U12715 (N_12715,N_6479,N_7810);
and U12716 (N_12716,N_5918,N_7482);
and U12717 (N_12717,N_8602,N_6840);
or U12718 (N_12718,N_5161,N_8117);
nand U12719 (N_12719,N_5219,N_8451);
or U12720 (N_12720,N_6662,N_9751);
xnor U12721 (N_12721,N_7863,N_9488);
or U12722 (N_12722,N_5604,N_7815);
or U12723 (N_12723,N_8214,N_6052);
or U12724 (N_12724,N_9737,N_5160);
and U12725 (N_12725,N_7213,N_9206);
nor U12726 (N_12726,N_8296,N_6648);
and U12727 (N_12727,N_8395,N_9802);
xor U12728 (N_12728,N_6769,N_5400);
or U12729 (N_12729,N_6355,N_6071);
xor U12730 (N_12730,N_5482,N_5639);
nand U12731 (N_12731,N_8845,N_6539);
xnor U12732 (N_12732,N_7119,N_9135);
xor U12733 (N_12733,N_6566,N_8898);
nor U12734 (N_12734,N_9726,N_9345);
xnor U12735 (N_12735,N_5838,N_9882);
xor U12736 (N_12736,N_9413,N_5418);
and U12737 (N_12737,N_9975,N_9245);
xor U12738 (N_12738,N_8807,N_9729);
xor U12739 (N_12739,N_6453,N_8496);
or U12740 (N_12740,N_8649,N_8176);
xor U12741 (N_12741,N_5493,N_8100);
xor U12742 (N_12742,N_7288,N_8962);
nor U12743 (N_12743,N_6837,N_8173);
nand U12744 (N_12744,N_5332,N_7712);
or U12745 (N_12745,N_8808,N_9431);
nand U12746 (N_12746,N_9579,N_7924);
or U12747 (N_12747,N_6089,N_6879);
nor U12748 (N_12748,N_5439,N_7065);
nand U12749 (N_12749,N_7321,N_6356);
nand U12750 (N_12750,N_8313,N_8941);
xnor U12751 (N_12751,N_9593,N_7239);
nor U12752 (N_12752,N_6958,N_9593);
or U12753 (N_12753,N_6521,N_6492);
xnor U12754 (N_12754,N_6145,N_9661);
xor U12755 (N_12755,N_7762,N_8825);
nand U12756 (N_12756,N_8633,N_7373);
xnor U12757 (N_12757,N_6945,N_6685);
nand U12758 (N_12758,N_6685,N_6026);
xor U12759 (N_12759,N_6873,N_6950);
nor U12760 (N_12760,N_9342,N_8642);
and U12761 (N_12761,N_7365,N_5373);
or U12762 (N_12762,N_8101,N_8453);
and U12763 (N_12763,N_8172,N_7356);
nor U12764 (N_12764,N_8645,N_6731);
and U12765 (N_12765,N_7581,N_9533);
nor U12766 (N_12766,N_7385,N_6900);
xnor U12767 (N_12767,N_6839,N_9878);
nor U12768 (N_12768,N_5901,N_7189);
nor U12769 (N_12769,N_5717,N_9318);
nand U12770 (N_12770,N_9705,N_6406);
or U12771 (N_12771,N_6687,N_8596);
nor U12772 (N_12772,N_5852,N_7161);
and U12773 (N_12773,N_5790,N_9804);
or U12774 (N_12774,N_7416,N_6271);
nor U12775 (N_12775,N_8978,N_9383);
nand U12776 (N_12776,N_7152,N_6237);
xor U12777 (N_12777,N_9591,N_7549);
nand U12778 (N_12778,N_9001,N_7626);
and U12779 (N_12779,N_9098,N_9269);
xnor U12780 (N_12780,N_8299,N_8061);
nor U12781 (N_12781,N_6912,N_6901);
xor U12782 (N_12782,N_5589,N_6512);
or U12783 (N_12783,N_9930,N_7387);
nor U12784 (N_12784,N_9931,N_8637);
nand U12785 (N_12785,N_5752,N_9417);
nand U12786 (N_12786,N_8845,N_8207);
nand U12787 (N_12787,N_8107,N_6940);
or U12788 (N_12788,N_6874,N_9864);
or U12789 (N_12789,N_6363,N_9246);
nor U12790 (N_12790,N_6376,N_7394);
xnor U12791 (N_12791,N_5356,N_9377);
xnor U12792 (N_12792,N_5713,N_5304);
nand U12793 (N_12793,N_6754,N_5562);
and U12794 (N_12794,N_7535,N_9511);
or U12795 (N_12795,N_8623,N_6122);
or U12796 (N_12796,N_6003,N_6305);
nor U12797 (N_12797,N_5748,N_5146);
and U12798 (N_12798,N_7254,N_5868);
and U12799 (N_12799,N_9653,N_8026);
nand U12800 (N_12800,N_8242,N_8065);
or U12801 (N_12801,N_9319,N_9777);
and U12802 (N_12802,N_9878,N_8164);
xnor U12803 (N_12803,N_5118,N_7785);
or U12804 (N_12804,N_6626,N_9902);
nand U12805 (N_12805,N_7832,N_7697);
nor U12806 (N_12806,N_8938,N_5500);
nor U12807 (N_12807,N_8987,N_6381);
and U12808 (N_12808,N_6511,N_8944);
nand U12809 (N_12809,N_7120,N_5876);
or U12810 (N_12810,N_5690,N_9296);
nand U12811 (N_12811,N_6934,N_8945);
and U12812 (N_12812,N_7438,N_9891);
and U12813 (N_12813,N_6970,N_5050);
and U12814 (N_12814,N_5650,N_7541);
nor U12815 (N_12815,N_6049,N_9512);
or U12816 (N_12816,N_7605,N_8986);
or U12817 (N_12817,N_6028,N_7362);
nor U12818 (N_12818,N_7144,N_6161);
nand U12819 (N_12819,N_9466,N_5009);
nand U12820 (N_12820,N_7022,N_9650);
xor U12821 (N_12821,N_7561,N_8599);
or U12822 (N_12822,N_7472,N_8640);
nand U12823 (N_12823,N_7578,N_5800);
and U12824 (N_12824,N_7629,N_8301);
nand U12825 (N_12825,N_6813,N_7585);
nor U12826 (N_12826,N_8891,N_7334);
and U12827 (N_12827,N_9824,N_7681);
nand U12828 (N_12828,N_5995,N_7573);
xnor U12829 (N_12829,N_8091,N_8033);
and U12830 (N_12830,N_9912,N_8835);
and U12831 (N_12831,N_9775,N_9095);
and U12832 (N_12832,N_8248,N_6243);
nand U12833 (N_12833,N_5681,N_8405);
nor U12834 (N_12834,N_9818,N_9443);
xnor U12835 (N_12835,N_7531,N_9055);
or U12836 (N_12836,N_5010,N_7293);
nor U12837 (N_12837,N_9976,N_8489);
or U12838 (N_12838,N_6066,N_6598);
nor U12839 (N_12839,N_7791,N_9314);
nand U12840 (N_12840,N_8267,N_7340);
nand U12841 (N_12841,N_9240,N_8166);
nor U12842 (N_12842,N_7837,N_9321);
and U12843 (N_12843,N_8120,N_9783);
xnor U12844 (N_12844,N_6879,N_7971);
nor U12845 (N_12845,N_8541,N_5382);
or U12846 (N_12846,N_8696,N_8944);
nor U12847 (N_12847,N_8107,N_5360);
or U12848 (N_12848,N_5964,N_6891);
nor U12849 (N_12849,N_8603,N_9028);
xor U12850 (N_12850,N_6257,N_5935);
or U12851 (N_12851,N_5937,N_8447);
xnor U12852 (N_12852,N_9532,N_5920);
and U12853 (N_12853,N_6047,N_7636);
nand U12854 (N_12854,N_7885,N_9607);
or U12855 (N_12855,N_8074,N_9114);
nand U12856 (N_12856,N_8678,N_6391);
nand U12857 (N_12857,N_8425,N_5548);
or U12858 (N_12858,N_9751,N_8913);
nand U12859 (N_12859,N_7429,N_9872);
nand U12860 (N_12860,N_7585,N_5672);
xnor U12861 (N_12861,N_5648,N_8754);
nand U12862 (N_12862,N_6720,N_7600);
nand U12863 (N_12863,N_5838,N_7703);
nor U12864 (N_12864,N_5556,N_5626);
nor U12865 (N_12865,N_8213,N_7797);
nor U12866 (N_12866,N_6536,N_7038);
nor U12867 (N_12867,N_7621,N_6763);
and U12868 (N_12868,N_7239,N_9821);
and U12869 (N_12869,N_6068,N_7137);
or U12870 (N_12870,N_6516,N_5286);
nor U12871 (N_12871,N_9207,N_7457);
or U12872 (N_12872,N_5365,N_8707);
xnor U12873 (N_12873,N_6536,N_8178);
or U12874 (N_12874,N_8330,N_8685);
and U12875 (N_12875,N_9264,N_6683);
nand U12876 (N_12876,N_5241,N_5772);
nor U12877 (N_12877,N_7002,N_9411);
and U12878 (N_12878,N_6797,N_8057);
nand U12879 (N_12879,N_5042,N_6376);
xnor U12880 (N_12880,N_8153,N_6818);
and U12881 (N_12881,N_9659,N_8428);
nor U12882 (N_12882,N_5057,N_9997);
and U12883 (N_12883,N_8105,N_7344);
and U12884 (N_12884,N_9514,N_8187);
and U12885 (N_12885,N_8740,N_8077);
nand U12886 (N_12886,N_8220,N_6386);
or U12887 (N_12887,N_9995,N_6319);
and U12888 (N_12888,N_5783,N_8529);
nor U12889 (N_12889,N_9084,N_9247);
or U12890 (N_12890,N_7334,N_7150);
xor U12891 (N_12891,N_6877,N_5549);
xnor U12892 (N_12892,N_6644,N_9722);
nand U12893 (N_12893,N_7738,N_7172);
nor U12894 (N_12894,N_9550,N_6041);
xor U12895 (N_12895,N_6377,N_8664);
nand U12896 (N_12896,N_9713,N_9201);
xor U12897 (N_12897,N_9337,N_8392);
nand U12898 (N_12898,N_5441,N_9376);
or U12899 (N_12899,N_9658,N_6023);
nand U12900 (N_12900,N_5947,N_5871);
xnor U12901 (N_12901,N_9919,N_9684);
or U12902 (N_12902,N_6521,N_6496);
nor U12903 (N_12903,N_5742,N_7311);
and U12904 (N_12904,N_5518,N_6251);
xnor U12905 (N_12905,N_9992,N_5823);
and U12906 (N_12906,N_5781,N_5901);
nor U12907 (N_12907,N_9910,N_7753);
or U12908 (N_12908,N_8185,N_8560);
xor U12909 (N_12909,N_8307,N_8148);
and U12910 (N_12910,N_7851,N_7007);
nor U12911 (N_12911,N_8660,N_9865);
xor U12912 (N_12912,N_8270,N_7519);
nand U12913 (N_12913,N_7591,N_9579);
nand U12914 (N_12914,N_5528,N_8280);
and U12915 (N_12915,N_8010,N_8591);
xnor U12916 (N_12916,N_6232,N_8838);
or U12917 (N_12917,N_5979,N_8148);
nand U12918 (N_12918,N_6966,N_8520);
and U12919 (N_12919,N_7300,N_6565);
or U12920 (N_12920,N_9182,N_9215);
xnor U12921 (N_12921,N_8206,N_9484);
or U12922 (N_12922,N_5735,N_7676);
xnor U12923 (N_12923,N_7736,N_5134);
or U12924 (N_12924,N_6635,N_7215);
nand U12925 (N_12925,N_5831,N_8423);
nand U12926 (N_12926,N_5327,N_9589);
and U12927 (N_12927,N_6975,N_7760);
nor U12928 (N_12928,N_6606,N_6253);
nand U12929 (N_12929,N_5207,N_5088);
and U12930 (N_12930,N_6515,N_7498);
nand U12931 (N_12931,N_6776,N_9130);
or U12932 (N_12932,N_8757,N_6602);
and U12933 (N_12933,N_5584,N_5947);
or U12934 (N_12934,N_6617,N_7392);
and U12935 (N_12935,N_5272,N_5755);
nand U12936 (N_12936,N_9095,N_8149);
and U12937 (N_12937,N_7865,N_6804);
nor U12938 (N_12938,N_5435,N_9484);
or U12939 (N_12939,N_7279,N_7049);
nand U12940 (N_12940,N_9790,N_8561);
nand U12941 (N_12941,N_9338,N_8424);
or U12942 (N_12942,N_8571,N_8572);
and U12943 (N_12943,N_9977,N_8217);
or U12944 (N_12944,N_6987,N_6726);
xnor U12945 (N_12945,N_9219,N_9456);
nor U12946 (N_12946,N_9253,N_5558);
and U12947 (N_12947,N_6305,N_6975);
or U12948 (N_12948,N_5287,N_8111);
nor U12949 (N_12949,N_6343,N_5901);
and U12950 (N_12950,N_5523,N_6125);
and U12951 (N_12951,N_7010,N_6291);
xor U12952 (N_12952,N_5963,N_7481);
and U12953 (N_12953,N_9661,N_9927);
or U12954 (N_12954,N_6104,N_5620);
and U12955 (N_12955,N_7911,N_8647);
or U12956 (N_12956,N_5142,N_8773);
nor U12957 (N_12957,N_6264,N_8035);
nand U12958 (N_12958,N_5720,N_8399);
nor U12959 (N_12959,N_6449,N_7390);
nand U12960 (N_12960,N_9896,N_7621);
nand U12961 (N_12961,N_7670,N_6460);
nand U12962 (N_12962,N_6132,N_5395);
xnor U12963 (N_12963,N_6478,N_6914);
xnor U12964 (N_12964,N_5418,N_6653);
or U12965 (N_12965,N_5648,N_5417);
or U12966 (N_12966,N_7715,N_9821);
and U12967 (N_12967,N_9850,N_6139);
nor U12968 (N_12968,N_8882,N_6706);
and U12969 (N_12969,N_6293,N_5608);
nand U12970 (N_12970,N_9960,N_9776);
nor U12971 (N_12971,N_5527,N_6662);
nand U12972 (N_12972,N_6246,N_8733);
or U12973 (N_12973,N_5839,N_7681);
nand U12974 (N_12974,N_6391,N_9583);
and U12975 (N_12975,N_5694,N_9997);
nand U12976 (N_12976,N_8168,N_7087);
or U12977 (N_12977,N_8190,N_5163);
nand U12978 (N_12978,N_6373,N_6838);
nand U12979 (N_12979,N_6125,N_6679);
or U12980 (N_12980,N_7753,N_6865);
and U12981 (N_12981,N_8264,N_5767);
or U12982 (N_12982,N_6176,N_8137);
nor U12983 (N_12983,N_9184,N_9747);
xor U12984 (N_12984,N_9937,N_6307);
xnor U12985 (N_12985,N_9064,N_9991);
and U12986 (N_12986,N_9070,N_6655);
and U12987 (N_12987,N_8318,N_5322);
xor U12988 (N_12988,N_9691,N_5206);
or U12989 (N_12989,N_5461,N_5974);
or U12990 (N_12990,N_7766,N_7465);
xnor U12991 (N_12991,N_8272,N_9704);
nand U12992 (N_12992,N_8594,N_7668);
xor U12993 (N_12993,N_5464,N_7639);
xnor U12994 (N_12994,N_7555,N_5474);
nand U12995 (N_12995,N_8523,N_5848);
and U12996 (N_12996,N_9866,N_9663);
nand U12997 (N_12997,N_7033,N_9380);
or U12998 (N_12998,N_5987,N_8971);
xor U12999 (N_12999,N_5946,N_7959);
nor U13000 (N_13000,N_6524,N_8921);
or U13001 (N_13001,N_5918,N_5051);
nand U13002 (N_13002,N_9159,N_9143);
and U13003 (N_13003,N_7985,N_9366);
xor U13004 (N_13004,N_9907,N_6212);
nand U13005 (N_13005,N_8658,N_6736);
or U13006 (N_13006,N_6796,N_5186);
xor U13007 (N_13007,N_7236,N_7319);
and U13008 (N_13008,N_5509,N_6916);
nand U13009 (N_13009,N_7385,N_8268);
nor U13010 (N_13010,N_6162,N_5325);
and U13011 (N_13011,N_6907,N_9569);
and U13012 (N_13012,N_7266,N_8186);
or U13013 (N_13013,N_7402,N_7723);
nand U13014 (N_13014,N_9144,N_8297);
nor U13015 (N_13015,N_7533,N_7231);
nor U13016 (N_13016,N_9061,N_7380);
and U13017 (N_13017,N_6610,N_6876);
or U13018 (N_13018,N_6647,N_8671);
xnor U13019 (N_13019,N_8520,N_9825);
or U13020 (N_13020,N_6800,N_7688);
nor U13021 (N_13021,N_9341,N_6949);
xnor U13022 (N_13022,N_8325,N_8761);
xnor U13023 (N_13023,N_5073,N_8448);
or U13024 (N_13024,N_7811,N_6004);
nor U13025 (N_13025,N_6728,N_8555);
nor U13026 (N_13026,N_7681,N_8054);
nor U13027 (N_13027,N_8749,N_5425);
nor U13028 (N_13028,N_6572,N_5858);
nand U13029 (N_13029,N_6376,N_6118);
nor U13030 (N_13030,N_6920,N_7782);
xnor U13031 (N_13031,N_5709,N_8307);
nand U13032 (N_13032,N_5674,N_9316);
or U13033 (N_13033,N_8950,N_8542);
or U13034 (N_13034,N_6198,N_7294);
nor U13035 (N_13035,N_5689,N_9796);
and U13036 (N_13036,N_8911,N_7488);
and U13037 (N_13037,N_7220,N_7365);
nand U13038 (N_13038,N_6150,N_8367);
or U13039 (N_13039,N_5091,N_8635);
xor U13040 (N_13040,N_7392,N_5054);
or U13041 (N_13041,N_5033,N_6208);
and U13042 (N_13042,N_5168,N_5093);
nor U13043 (N_13043,N_8417,N_5245);
nor U13044 (N_13044,N_9976,N_7995);
and U13045 (N_13045,N_8606,N_5395);
xnor U13046 (N_13046,N_9854,N_9647);
nor U13047 (N_13047,N_6839,N_6709);
nor U13048 (N_13048,N_6320,N_5435);
xor U13049 (N_13049,N_8000,N_9385);
and U13050 (N_13050,N_8245,N_7671);
nand U13051 (N_13051,N_5440,N_9207);
xor U13052 (N_13052,N_9359,N_9365);
nand U13053 (N_13053,N_6368,N_9399);
and U13054 (N_13054,N_8248,N_7134);
and U13055 (N_13055,N_8880,N_7360);
or U13056 (N_13056,N_8750,N_6165);
nor U13057 (N_13057,N_8521,N_5277);
or U13058 (N_13058,N_6867,N_5095);
xnor U13059 (N_13059,N_7215,N_9408);
and U13060 (N_13060,N_8591,N_9441);
xor U13061 (N_13061,N_9036,N_5466);
nor U13062 (N_13062,N_5598,N_9376);
or U13063 (N_13063,N_9862,N_5582);
nand U13064 (N_13064,N_7873,N_8930);
and U13065 (N_13065,N_9645,N_7697);
and U13066 (N_13066,N_6334,N_8194);
nor U13067 (N_13067,N_7248,N_7792);
nand U13068 (N_13068,N_7977,N_9290);
nand U13069 (N_13069,N_5313,N_9922);
xnor U13070 (N_13070,N_5667,N_9860);
and U13071 (N_13071,N_9819,N_7091);
nand U13072 (N_13072,N_8197,N_8113);
and U13073 (N_13073,N_6490,N_5030);
nor U13074 (N_13074,N_5020,N_8533);
nor U13075 (N_13075,N_7923,N_7596);
nand U13076 (N_13076,N_5749,N_6363);
or U13077 (N_13077,N_7271,N_6977);
and U13078 (N_13078,N_5235,N_6740);
nor U13079 (N_13079,N_7117,N_8299);
nand U13080 (N_13080,N_6375,N_5138);
and U13081 (N_13081,N_5676,N_8291);
or U13082 (N_13082,N_6020,N_8335);
xor U13083 (N_13083,N_6503,N_5196);
nor U13084 (N_13084,N_5445,N_7986);
xor U13085 (N_13085,N_5750,N_5136);
or U13086 (N_13086,N_6674,N_7702);
nand U13087 (N_13087,N_8836,N_9503);
xnor U13088 (N_13088,N_8950,N_8040);
nand U13089 (N_13089,N_7885,N_6417);
nor U13090 (N_13090,N_5757,N_6758);
or U13091 (N_13091,N_6469,N_7062);
nor U13092 (N_13092,N_7288,N_6794);
and U13093 (N_13093,N_5897,N_7937);
nor U13094 (N_13094,N_8510,N_5800);
xnor U13095 (N_13095,N_5811,N_9816);
xnor U13096 (N_13096,N_8347,N_9507);
nand U13097 (N_13097,N_9128,N_8204);
and U13098 (N_13098,N_6016,N_6138);
and U13099 (N_13099,N_8525,N_8239);
and U13100 (N_13100,N_7769,N_8005);
xor U13101 (N_13101,N_5912,N_5061);
or U13102 (N_13102,N_7942,N_7958);
and U13103 (N_13103,N_5896,N_7574);
or U13104 (N_13104,N_5330,N_6380);
xor U13105 (N_13105,N_9560,N_6183);
nand U13106 (N_13106,N_9228,N_9211);
and U13107 (N_13107,N_7924,N_9014);
and U13108 (N_13108,N_6688,N_7808);
xnor U13109 (N_13109,N_6505,N_9239);
nor U13110 (N_13110,N_8342,N_7266);
nor U13111 (N_13111,N_6798,N_5702);
xor U13112 (N_13112,N_8358,N_5578);
xor U13113 (N_13113,N_8012,N_5119);
xor U13114 (N_13114,N_7087,N_7100);
nor U13115 (N_13115,N_6800,N_7408);
or U13116 (N_13116,N_8858,N_7157);
and U13117 (N_13117,N_9109,N_7953);
xnor U13118 (N_13118,N_6331,N_5470);
nor U13119 (N_13119,N_7375,N_5369);
and U13120 (N_13120,N_5215,N_6923);
or U13121 (N_13121,N_8573,N_8630);
or U13122 (N_13122,N_5564,N_7012);
xnor U13123 (N_13123,N_5978,N_8329);
and U13124 (N_13124,N_5559,N_9386);
xor U13125 (N_13125,N_5453,N_7630);
nor U13126 (N_13126,N_7315,N_5902);
xnor U13127 (N_13127,N_8111,N_8334);
or U13128 (N_13128,N_7977,N_8579);
nand U13129 (N_13129,N_6900,N_6147);
and U13130 (N_13130,N_5175,N_5720);
xor U13131 (N_13131,N_8483,N_5487);
nor U13132 (N_13132,N_7753,N_5979);
or U13133 (N_13133,N_6116,N_9798);
nor U13134 (N_13134,N_8521,N_5502);
or U13135 (N_13135,N_7480,N_5887);
nor U13136 (N_13136,N_9822,N_6341);
nor U13137 (N_13137,N_7562,N_9352);
xnor U13138 (N_13138,N_9989,N_9888);
nor U13139 (N_13139,N_8111,N_5560);
nand U13140 (N_13140,N_6347,N_8934);
nor U13141 (N_13141,N_7499,N_6526);
nand U13142 (N_13142,N_9839,N_7190);
xnor U13143 (N_13143,N_6046,N_9241);
or U13144 (N_13144,N_6022,N_9596);
or U13145 (N_13145,N_8246,N_6147);
nand U13146 (N_13146,N_6278,N_6194);
xor U13147 (N_13147,N_8720,N_6527);
and U13148 (N_13148,N_7980,N_6630);
nor U13149 (N_13149,N_5799,N_9453);
and U13150 (N_13150,N_9471,N_9738);
and U13151 (N_13151,N_9180,N_9504);
nor U13152 (N_13152,N_6024,N_7491);
xnor U13153 (N_13153,N_5794,N_6372);
nor U13154 (N_13154,N_9072,N_6160);
xnor U13155 (N_13155,N_6698,N_9494);
and U13156 (N_13156,N_5521,N_5949);
xor U13157 (N_13157,N_7972,N_8936);
nand U13158 (N_13158,N_7653,N_7289);
nand U13159 (N_13159,N_6326,N_6366);
xnor U13160 (N_13160,N_7631,N_5307);
nand U13161 (N_13161,N_5142,N_8711);
nand U13162 (N_13162,N_7432,N_5811);
and U13163 (N_13163,N_5153,N_7798);
nand U13164 (N_13164,N_8417,N_7722);
and U13165 (N_13165,N_6014,N_5157);
nor U13166 (N_13166,N_5340,N_6416);
nor U13167 (N_13167,N_5949,N_9475);
or U13168 (N_13168,N_5203,N_5117);
nor U13169 (N_13169,N_6327,N_9410);
nor U13170 (N_13170,N_9670,N_7368);
xnor U13171 (N_13171,N_7755,N_6204);
and U13172 (N_13172,N_5145,N_7223);
nand U13173 (N_13173,N_8268,N_6313);
nor U13174 (N_13174,N_7320,N_8059);
or U13175 (N_13175,N_8541,N_8222);
or U13176 (N_13176,N_6557,N_5218);
or U13177 (N_13177,N_7816,N_9536);
and U13178 (N_13178,N_6752,N_7307);
or U13179 (N_13179,N_6525,N_7836);
or U13180 (N_13180,N_6741,N_7200);
and U13181 (N_13181,N_9560,N_9701);
xor U13182 (N_13182,N_6587,N_5125);
xor U13183 (N_13183,N_5548,N_5952);
nor U13184 (N_13184,N_6792,N_9027);
xnor U13185 (N_13185,N_5808,N_9684);
and U13186 (N_13186,N_8564,N_6822);
and U13187 (N_13187,N_9099,N_8095);
xnor U13188 (N_13188,N_7349,N_5559);
nor U13189 (N_13189,N_6086,N_9236);
nand U13190 (N_13190,N_5309,N_7616);
or U13191 (N_13191,N_9718,N_8612);
and U13192 (N_13192,N_7588,N_5782);
nor U13193 (N_13193,N_7717,N_8198);
nor U13194 (N_13194,N_6439,N_5870);
nor U13195 (N_13195,N_7184,N_6963);
nor U13196 (N_13196,N_7285,N_5908);
nor U13197 (N_13197,N_7953,N_7472);
nand U13198 (N_13198,N_8817,N_5386);
nand U13199 (N_13199,N_6045,N_9468);
and U13200 (N_13200,N_7073,N_6268);
or U13201 (N_13201,N_5750,N_6727);
nand U13202 (N_13202,N_6458,N_8658);
nand U13203 (N_13203,N_7786,N_7672);
nand U13204 (N_13204,N_8533,N_7427);
and U13205 (N_13205,N_8925,N_8587);
or U13206 (N_13206,N_6285,N_5182);
nor U13207 (N_13207,N_7337,N_7235);
or U13208 (N_13208,N_7835,N_8590);
nand U13209 (N_13209,N_9173,N_7215);
or U13210 (N_13210,N_6717,N_9493);
nor U13211 (N_13211,N_9143,N_7757);
or U13212 (N_13212,N_8191,N_6125);
or U13213 (N_13213,N_7038,N_6654);
or U13214 (N_13214,N_6906,N_8406);
or U13215 (N_13215,N_5362,N_5292);
nand U13216 (N_13216,N_7616,N_5051);
nor U13217 (N_13217,N_9531,N_7848);
xor U13218 (N_13218,N_7653,N_6268);
nand U13219 (N_13219,N_8319,N_9583);
and U13220 (N_13220,N_7104,N_5940);
nor U13221 (N_13221,N_7279,N_9539);
and U13222 (N_13222,N_7024,N_7921);
or U13223 (N_13223,N_6332,N_8672);
and U13224 (N_13224,N_8561,N_6503);
or U13225 (N_13225,N_8752,N_9652);
or U13226 (N_13226,N_6791,N_7988);
or U13227 (N_13227,N_8304,N_7817);
nand U13228 (N_13228,N_5108,N_7861);
nor U13229 (N_13229,N_6297,N_7434);
nand U13230 (N_13230,N_5729,N_5845);
nor U13231 (N_13231,N_5205,N_6975);
nor U13232 (N_13232,N_6173,N_6685);
xor U13233 (N_13233,N_8604,N_7283);
nand U13234 (N_13234,N_5622,N_8941);
or U13235 (N_13235,N_8718,N_7110);
and U13236 (N_13236,N_5074,N_9970);
or U13237 (N_13237,N_5031,N_9060);
and U13238 (N_13238,N_5037,N_6983);
nand U13239 (N_13239,N_9302,N_9604);
nand U13240 (N_13240,N_8708,N_7659);
nor U13241 (N_13241,N_8685,N_6626);
nor U13242 (N_13242,N_6368,N_6705);
xnor U13243 (N_13243,N_5395,N_7345);
xor U13244 (N_13244,N_9335,N_6264);
nor U13245 (N_13245,N_7597,N_7331);
and U13246 (N_13246,N_6739,N_7104);
nor U13247 (N_13247,N_5388,N_6420);
and U13248 (N_13248,N_7114,N_8800);
or U13249 (N_13249,N_9029,N_7049);
xor U13250 (N_13250,N_9200,N_9328);
and U13251 (N_13251,N_8322,N_8187);
nand U13252 (N_13252,N_5144,N_7474);
or U13253 (N_13253,N_5804,N_5113);
or U13254 (N_13254,N_6513,N_5128);
nor U13255 (N_13255,N_5764,N_9400);
xor U13256 (N_13256,N_6621,N_7535);
nor U13257 (N_13257,N_9283,N_8266);
nor U13258 (N_13258,N_9533,N_8490);
or U13259 (N_13259,N_9583,N_7814);
nand U13260 (N_13260,N_7788,N_8635);
xor U13261 (N_13261,N_6702,N_7895);
or U13262 (N_13262,N_8467,N_8810);
nor U13263 (N_13263,N_9793,N_8668);
nand U13264 (N_13264,N_6929,N_9506);
nand U13265 (N_13265,N_5455,N_7518);
or U13266 (N_13266,N_8521,N_6693);
nor U13267 (N_13267,N_5435,N_9017);
and U13268 (N_13268,N_5974,N_9336);
nand U13269 (N_13269,N_7532,N_8454);
or U13270 (N_13270,N_7907,N_9459);
xor U13271 (N_13271,N_8268,N_6908);
or U13272 (N_13272,N_6679,N_9199);
or U13273 (N_13273,N_6836,N_9367);
or U13274 (N_13274,N_5233,N_9620);
xnor U13275 (N_13275,N_6624,N_8863);
or U13276 (N_13276,N_8505,N_7642);
xor U13277 (N_13277,N_7592,N_5049);
nor U13278 (N_13278,N_7542,N_5665);
nor U13279 (N_13279,N_5799,N_5318);
nand U13280 (N_13280,N_8574,N_5289);
xor U13281 (N_13281,N_6269,N_8152);
nand U13282 (N_13282,N_5183,N_8519);
nor U13283 (N_13283,N_6354,N_9951);
and U13284 (N_13284,N_5739,N_6899);
and U13285 (N_13285,N_6490,N_8854);
or U13286 (N_13286,N_5258,N_5131);
nor U13287 (N_13287,N_7631,N_6851);
and U13288 (N_13288,N_8591,N_8595);
or U13289 (N_13289,N_6203,N_9911);
nor U13290 (N_13290,N_7080,N_5632);
xnor U13291 (N_13291,N_6155,N_6592);
or U13292 (N_13292,N_8407,N_8347);
and U13293 (N_13293,N_8665,N_8922);
or U13294 (N_13294,N_5714,N_7502);
xor U13295 (N_13295,N_8769,N_7050);
nand U13296 (N_13296,N_9948,N_8455);
nor U13297 (N_13297,N_5510,N_7909);
xor U13298 (N_13298,N_6501,N_8392);
or U13299 (N_13299,N_5803,N_7139);
xnor U13300 (N_13300,N_5074,N_9974);
and U13301 (N_13301,N_5765,N_6463);
or U13302 (N_13302,N_8079,N_9905);
and U13303 (N_13303,N_5809,N_5582);
or U13304 (N_13304,N_6356,N_5539);
nor U13305 (N_13305,N_8494,N_5561);
or U13306 (N_13306,N_5735,N_5732);
nand U13307 (N_13307,N_7242,N_8219);
or U13308 (N_13308,N_5527,N_9897);
xnor U13309 (N_13309,N_8340,N_5656);
and U13310 (N_13310,N_9169,N_7674);
xnor U13311 (N_13311,N_6707,N_8192);
xor U13312 (N_13312,N_9109,N_9454);
nand U13313 (N_13313,N_8193,N_5596);
nand U13314 (N_13314,N_9395,N_6602);
or U13315 (N_13315,N_8383,N_7283);
xnor U13316 (N_13316,N_8040,N_9690);
and U13317 (N_13317,N_7105,N_6585);
or U13318 (N_13318,N_6465,N_8011);
nand U13319 (N_13319,N_8951,N_8427);
and U13320 (N_13320,N_9523,N_7099);
nor U13321 (N_13321,N_8624,N_8848);
xor U13322 (N_13322,N_7890,N_6256);
and U13323 (N_13323,N_6292,N_8925);
and U13324 (N_13324,N_6006,N_5099);
or U13325 (N_13325,N_8042,N_8821);
or U13326 (N_13326,N_5520,N_5439);
nor U13327 (N_13327,N_9554,N_6280);
xor U13328 (N_13328,N_5516,N_8446);
nor U13329 (N_13329,N_9835,N_5751);
or U13330 (N_13330,N_8066,N_7180);
or U13331 (N_13331,N_6898,N_7830);
xor U13332 (N_13332,N_6945,N_8358);
xor U13333 (N_13333,N_8279,N_6678);
xor U13334 (N_13334,N_8019,N_6696);
or U13335 (N_13335,N_8476,N_5635);
nand U13336 (N_13336,N_6167,N_8975);
or U13337 (N_13337,N_9644,N_9744);
nor U13338 (N_13338,N_6609,N_7027);
and U13339 (N_13339,N_6212,N_8271);
nor U13340 (N_13340,N_9790,N_9842);
xnor U13341 (N_13341,N_5262,N_8477);
nand U13342 (N_13342,N_8171,N_6276);
nand U13343 (N_13343,N_9860,N_8046);
xor U13344 (N_13344,N_8076,N_8578);
or U13345 (N_13345,N_8410,N_6886);
xnor U13346 (N_13346,N_7543,N_6217);
and U13347 (N_13347,N_7976,N_9863);
xor U13348 (N_13348,N_9896,N_9529);
and U13349 (N_13349,N_6423,N_8604);
or U13350 (N_13350,N_9411,N_9501);
and U13351 (N_13351,N_9712,N_7543);
nand U13352 (N_13352,N_8735,N_8626);
nand U13353 (N_13353,N_5968,N_5069);
or U13354 (N_13354,N_8234,N_7612);
nand U13355 (N_13355,N_8132,N_6252);
or U13356 (N_13356,N_8365,N_5118);
nand U13357 (N_13357,N_7891,N_6860);
or U13358 (N_13358,N_7194,N_9588);
xor U13359 (N_13359,N_5523,N_5414);
nor U13360 (N_13360,N_5872,N_9604);
nand U13361 (N_13361,N_5698,N_9748);
nand U13362 (N_13362,N_6894,N_8378);
and U13363 (N_13363,N_9679,N_8711);
xnor U13364 (N_13364,N_5602,N_5188);
nand U13365 (N_13365,N_5162,N_5710);
or U13366 (N_13366,N_5202,N_5295);
nor U13367 (N_13367,N_5171,N_6472);
or U13368 (N_13368,N_5560,N_9875);
and U13369 (N_13369,N_7830,N_6144);
or U13370 (N_13370,N_7835,N_7713);
or U13371 (N_13371,N_6982,N_9200);
or U13372 (N_13372,N_5514,N_9616);
xor U13373 (N_13373,N_6475,N_7896);
xnor U13374 (N_13374,N_6155,N_9423);
and U13375 (N_13375,N_8172,N_5260);
and U13376 (N_13376,N_8499,N_5951);
or U13377 (N_13377,N_8930,N_6497);
nor U13378 (N_13378,N_9214,N_9933);
nand U13379 (N_13379,N_7230,N_9824);
xor U13380 (N_13380,N_6358,N_5586);
or U13381 (N_13381,N_6959,N_9812);
xor U13382 (N_13382,N_9419,N_6201);
xor U13383 (N_13383,N_5538,N_7287);
nor U13384 (N_13384,N_6184,N_8758);
and U13385 (N_13385,N_6962,N_6137);
xor U13386 (N_13386,N_5634,N_8716);
nor U13387 (N_13387,N_7510,N_5118);
or U13388 (N_13388,N_8067,N_5331);
xor U13389 (N_13389,N_6466,N_9991);
and U13390 (N_13390,N_8763,N_9276);
nand U13391 (N_13391,N_8593,N_9790);
or U13392 (N_13392,N_7061,N_7166);
or U13393 (N_13393,N_6210,N_6498);
and U13394 (N_13394,N_6756,N_6735);
xor U13395 (N_13395,N_5000,N_6070);
xor U13396 (N_13396,N_7701,N_5621);
nand U13397 (N_13397,N_5380,N_5643);
or U13398 (N_13398,N_9036,N_5518);
or U13399 (N_13399,N_6965,N_6828);
nand U13400 (N_13400,N_5824,N_6612);
nor U13401 (N_13401,N_5012,N_6180);
nor U13402 (N_13402,N_5175,N_9808);
and U13403 (N_13403,N_6039,N_9310);
xor U13404 (N_13404,N_6929,N_6347);
xor U13405 (N_13405,N_8683,N_9234);
nand U13406 (N_13406,N_7961,N_5190);
or U13407 (N_13407,N_9089,N_6602);
xor U13408 (N_13408,N_6727,N_7445);
nand U13409 (N_13409,N_6161,N_6834);
xor U13410 (N_13410,N_7569,N_9963);
nor U13411 (N_13411,N_5464,N_8351);
and U13412 (N_13412,N_7327,N_6172);
xor U13413 (N_13413,N_9998,N_6383);
or U13414 (N_13414,N_8951,N_6122);
nand U13415 (N_13415,N_9679,N_9759);
nor U13416 (N_13416,N_5913,N_8386);
xnor U13417 (N_13417,N_6069,N_5465);
nor U13418 (N_13418,N_6794,N_6920);
and U13419 (N_13419,N_5015,N_6284);
nor U13420 (N_13420,N_9778,N_5008);
xnor U13421 (N_13421,N_7181,N_5359);
or U13422 (N_13422,N_5660,N_5705);
or U13423 (N_13423,N_8437,N_9684);
nor U13424 (N_13424,N_7077,N_6907);
nand U13425 (N_13425,N_7490,N_5753);
nand U13426 (N_13426,N_6672,N_5797);
nand U13427 (N_13427,N_7576,N_7160);
nor U13428 (N_13428,N_7873,N_8058);
or U13429 (N_13429,N_6239,N_6488);
nor U13430 (N_13430,N_7849,N_8955);
nor U13431 (N_13431,N_7983,N_7078);
and U13432 (N_13432,N_9531,N_7942);
nor U13433 (N_13433,N_9353,N_8066);
nor U13434 (N_13434,N_7311,N_7833);
nand U13435 (N_13435,N_6509,N_8895);
xnor U13436 (N_13436,N_9687,N_8612);
xor U13437 (N_13437,N_5297,N_7429);
or U13438 (N_13438,N_7624,N_7558);
xnor U13439 (N_13439,N_5164,N_5823);
nand U13440 (N_13440,N_7988,N_7991);
nor U13441 (N_13441,N_8398,N_5078);
nand U13442 (N_13442,N_5703,N_8847);
or U13443 (N_13443,N_5704,N_5296);
xor U13444 (N_13444,N_8606,N_6358);
nand U13445 (N_13445,N_8648,N_6570);
xor U13446 (N_13446,N_5681,N_8460);
nor U13447 (N_13447,N_7190,N_8743);
or U13448 (N_13448,N_8396,N_5674);
nor U13449 (N_13449,N_9561,N_6522);
xnor U13450 (N_13450,N_5235,N_6050);
and U13451 (N_13451,N_7996,N_5765);
nor U13452 (N_13452,N_8918,N_6030);
and U13453 (N_13453,N_9822,N_8209);
nand U13454 (N_13454,N_8562,N_9277);
and U13455 (N_13455,N_6827,N_9106);
nand U13456 (N_13456,N_7620,N_7729);
nor U13457 (N_13457,N_5229,N_9368);
xnor U13458 (N_13458,N_5024,N_5120);
and U13459 (N_13459,N_6435,N_9735);
and U13460 (N_13460,N_6910,N_5015);
or U13461 (N_13461,N_7250,N_8526);
and U13462 (N_13462,N_9821,N_5041);
xnor U13463 (N_13463,N_6667,N_6340);
and U13464 (N_13464,N_6876,N_8008);
or U13465 (N_13465,N_8340,N_5681);
nand U13466 (N_13466,N_6677,N_7977);
nand U13467 (N_13467,N_6673,N_9882);
nand U13468 (N_13468,N_9422,N_7741);
and U13469 (N_13469,N_6373,N_7503);
or U13470 (N_13470,N_9439,N_5457);
and U13471 (N_13471,N_8931,N_5647);
nand U13472 (N_13472,N_7183,N_6742);
nand U13473 (N_13473,N_6557,N_8070);
or U13474 (N_13474,N_6994,N_6430);
and U13475 (N_13475,N_8003,N_8902);
nand U13476 (N_13476,N_6707,N_8657);
and U13477 (N_13477,N_7530,N_6592);
or U13478 (N_13478,N_5245,N_7910);
nand U13479 (N_13479,N_5263,N_6808);
xor U13480 (N_13480,N_8439,N_8278);
or U13481 (N_13481,N_6427,N_5488);
nor U13482 (N_13482,N_7062,N_6020);
and U13483 (N_13483,N_9440,N_7804);
nor U13484 (N_13484,N_7551,N_5953);
xnor U13485 (N_13485,N_5327,N_6401);
or U13486 (N_13486,N_6343,N_7942);
or U13487 (N_13487,N_5703,N_9028);
nand U13488 (N_13488,N_6012,N_5795);
nor U13489 (N_13489,N_9176,N_9863);
nor U13490 (N_13490,N_5648,N_5364);
nor U13491 (N_13491,N_8125,N_8855);
xor U13492 (N_13492,N_5606,N_6030);
nor U13493 (N_13493,N_6594,N_7734);
xnor U13494 (N_13494,N_6273,N_8559);
nor U13495 (N_13495,N_5099,N_9072);
xor U13496 (N_13496,N_6529,N_7923);
xnor U13497 (N_13497,N_5952,N_8026);
nor U13498 (N_13498,N_9528,N_9142);
and U13499 (N_13499,N_8685,N_5454);
and U13500 (N_13500,N_7666,N_7565);
nor U13501 (N_13501,N_8616,N_5014);
nor U13502 (N_13502,N_9105,N_5554);
nand U13503 (N_13503,N_5255,N_6699);
or U13504 (N_13504,N_8148,N_5308);
and U13505 (N_13505,N_5070,N_8459);
and U13506 (N_13506,N_9704,N_6669);
xor U13507 (N_13507,N_9282,N_5605);
xnor U13508 (N_13508,N_6104,N_9635);
or U13509 (N_13509,N_5507,N_9838);
nand U13510 (N_13510,N_8598,N_6507);
nor U13511 (N_13511,N_8394,N_5579);
nor U13512 (N_13512,N_8996,N_9978);
or U13513 (N_13513,N_8476,N_9643);
nand U13514 (N_13514,N_5353,N_6715);
nor U13515 (N_13515,N_8623,N_5163);
and U13516 (N_13516,N_7832,N_9382);
xnor U13517 (N_13517,N_9637,N_5549);
nor U13518 (N_13518,N_9271,N_7552);
and U13519 (N_13519,N_6779,N_6232);
or U13520 (N_13520,N_9948,N_7968);
and U13521 (N_13521,N_7163,N_6308);
xnor U13522 (N_13522,N_7420,N_7898);
xnor U13523 (N_13523,N_6334,N_8227);
xnor U13524 (N_13524,N_8957,N_7090);
nor U13525 (N_13525,N_8380,N_5707);
and U13526 (N_13526,N_8070,N_8394);
nand U13527 (N_13527,N_8413,N_8465);
nand U13528 (N_13528,N_5487,N_9339);
or U13529 (N_13529,N_6384,N_7897);
nand U13530 (N_13530,N_9056,N_7674);
xnor U13531 (N_13531,N_9589,N_5934);
nand U13532 (N_13532,N_5744,N_6480);
nand U13533 (N_13533,N_9643,N_7183);
or U13534 (N_13534,N_6784,N_6862);
or U13535 (N_13535,N_5867,N_6062);
nor U13536 (N_13536,N_8648,N_5189);
xor U13537 (N_13537,N_6840,N_5032);
xnor U13538 (N_13538,N_5486,N_9845);
or U13539 (N_13539,N_9773,N_8587);
nor U13540 (N_13540,N_9592,N_8630);
nor U13541 (N_13541,N_7452,N_5744);
or U13542 (N_13542,N_8168,N_8398);
nor U13543 (N_13543,N_8134,N_5616);
xor U13544 (N_13544,N_8722,N_6407);
nand U13545 (N_13545,N_8194,N_8300);
xor U13546 (N_13546,N_8823,N_5961);
nand U13547 (N_13547,N_5604,N_8992);
nor U13548 (N_13548,N_8377,N_5485);
xor U13549 (N_13549,N_8428,N_7115);
nor U13550 (N_13550,N_7840,N_6528);
nor U13551 (N_13551,N_6494,N_9041);
or U13552 (N_13552,N_5896,N_7312);
and U13553 (N_13553,N_9479,N_5698);
or U13554 (N_13554,N_6770,N_8186);
xnor U13555 (N_13555,N_9605,N_9484);
xor U13556 (N_13556,N_9488,N_7875);
or U13557 (N_13557,N_9552,N_5579);
and U13558 (N_13558,N_7164,N_7771);
and U13559 (N_13559,N_5588,N_5997);
or U13560 (N_13560,N_6400,N_5438);
and U13561 (N_13561,N_7423,N_7390);
nor U13562 (N_13562,N_5072,N_5280);
or U13563 (N_13563,N_7976,N_7827);
nand U13564 (N_13564,N_5085,N_7640);
and U13565 (N_13565,N_6359,N_6395);
and U13566 (N_13566,N_9126,N_8707);
nor U13567 (N_13567,N_8733,N_5042);
nor U13568 (N_13568,N_8974,N_6038);
nand U13569 (N_13569,N_8691,N_9441);
and U13570 (N_13570,N_6659,N_8603);
nor U13571 (N_13571,N_8233,N_6553);
or U13572 (N_13572,N_9237,N_5323);
or U13573 (N_13573,N_8695,N_8241);
and U13574 (N_13574,N_9114,N_8187);
nand U13575 (N_13575,N_5481,N_6778);
and U13576 (N_13576,N_6122,N_7250);
xnor U13577 (N_13577,N_9553,N_9811);
nor U13578 (N_13578,N_6815,N_7900);
xnor U13579 (N_13579,N_9539,N_6513);
or U13580 (N_13580,N_7070,N_7325);
or U13581 (N_13581,N_5158,N_7501);
nand U13582 (N_13582,N_7270,N_6532);
and U13583 (N_13583,N_7665,N_6091);
nor U13584 (N_13584,N_9148,N_6867);
and U13585 (N_13585,N_5683,N_9124);
xnor U13586 (N_13586,N_5580,N_8117);
and U13587 (N_13587,N_6812,N_7643);
nor U13588 (N_13588,N_5332,N_6269);
or U13589 (N_13589,N_6252,N_8309);
nor U13590 (N_13590,N_7711,N_5098);
nand U13591 (N_13591,N_5835,N_6993);
and U13592 (N_13592,N_7840,N_8704);
and U13593 (N_13593,N_7658,N_6757);
nand U13594 (N_13594,N_8462,N_7943);
and U13595 (N_13595,N_5575,N_6635);
and U13596 (N_13596,N_8150,N_7984);
or U13597 (N_13597,N_7703,N_6000);
nor U13598 (N_13598,N_7205,N_6056);
nor U13599 (N_13599,N_8241,N_9338);
xor U13600 (N_13600,N_6570,N_6255);
nor U13601 (N_13601,N_9668,N_7147);
nand U13602 (N_13602,N_5504,N_8377);
nand U13603 (N_13603,N_9309,N_7691);
or U13604 (N_13604,N_9998,N_9595);
or U13605 (N_13605,N_8340,N_6846);
and U13606 (N_13606,N_6236,N_8818);
nor U13607 (N_13607,N_8208,N_5588);
or U13608 (N_13608,N_9427,N_6199);
and U13609 (N_13609,N_5037,N_9654);
nand U13610 (N_13610,N_9129,N_9319);
or U13611 (N_13611,N_9548,N_5219);
nand U13612 (N_13612,N_5672,N_6628);
nor U13613 (N_13613,N_7949,N_7646);
or U13614 (N_13614,N_6910,N_6150);
nand U13615 (N_13615,N_9653,N_9851);
xnor U13616 (N_13616,N_9805,N_6149);
and U13617 (N_13617,N_7903,N_5800);
and U13618 (N_13618,N_8988,N_8418);
xor U13619 (N_13619,N_6454,N_9307);
xnor U13620 (N_13620,N_7970,N_5983);
and U13621 (N_13621,N_9505,N_8823);
nand U13622 (N_13622,N_9743,N_7940);
or U13623 (N_13623,N_7541,N_9758);
and U13624 (N_13624,N_8364,N_5625);
nand U13625 (N_13625,N_6705,N_7834);
and U13626 (N_13626,N_8900,N_8575);
and U13627 (N_13627,N_8403,N_8072);
xor U13628 (N_13628,N_8480,N_5902);
nor U13629 (N_13629,N_8625,N_9253);
nand U13630 (N_13630,N_5424,N_9670);
nand U13631 (N_13631,N_8072,N_6241);
and U13632 (N_13632,N_7639,N_5175);
xor U13633 (N_13633,N_8219,N_8805);
or U13634 (N_13634,N_6471,N_9313);
nand U13635 (N_13635,N_5548,N_9599);
nor U13636 (N_13636,N_5061,N_5995);
or U13637 (N_13637,N_9571,N_9050);
xnor U13638 (N_13638,N_6972,N_6999);
and U13639 (N_13639,N_5527,N_7726);
nor U13640 (N_13640,N_6138,N_7541);
xor U13641 (N_13641,N_5860,N_7213);
or U13642 (N_13642,N_5153,N_8302);
or U13643 (N_13643,N_6392,N_9895);
and U13644 (N_13644,N_8776,N_7618);
and U13645 (N_13645,N_5933,N_7499);
nor U13646 (N_13646,N_6100,N_6077);
xnor U13647 (N_13647,N_8733,N_9342);
nand U13648 (N_13648,N_8283,N_6516);
nand U13649 (N_13649,N_5906,N_6685);
xnor U13650 (N_13650,N_9314,N_6225);
nand U13651 (N_13651,N_9772,N_6273);
xor U13652 (N_13652,N_7926,N_9864);
nor U13653 (N_13653,N_6929,N_5504);
xnor U13654 (N_13654,N_6546,N_5166);
and U13655 (N_13655,N_8056,N_7966);
nand U13656 (N_13656,N_7554,N_8229);
nand U13657 (N_13657,N_5328,N_6541);
nand U13658 (N_13658,N_9335,N_5380);
and U13659 (N_13659,N_5353,N_9606);
xor U13660 (N_13660,N_5769,N_6927);
and U13661 (N_13661,N_7923,N_8235);
xor U13662 (N_13662,N_7303,N_6912);
xnor U13663 (N_13663,N_9046,N_8718);
nor U13664 (N_13664,N_8721,N_5190);
and U13665 (N_13665,N_7212,N_7304);
xnor U13666 (N_13666,N_5861,N_9310);
xor U13667 (N_13667,N_7312,N_5721);
or U13668 (N_13668,N_6685,N_6109);
xor U13669 (N_13669,N_7089,N_7505);
or U13670 (N_13670,N_8126,N_9420);
and U13671 (N_13671,N_6493,N_5916);
or U13672 (N_13672,N_9976,N_9570);
or U13673 (N_13673,N_7965,N_9427);
nand U13674 (N_13674,N_9062,N_7924);
or U13675 (N_13675,N_8032,N_9983);
xnor U13676 (N_13676,N_7761,N_8691);
xnor U13677 (N_13677,N_6857,N_8801);
and U13678 (N_13678,N_9219,N_8483);
and U13679 (N_13679,N_8294,N_7384);
xnor U13680 (N_13680,N_7247,N_9859);
or U13681 (N_13681,N_6857,N_8271);
nand U13682 (N_13682,N_7965,N_9148);
or U13683 (N_13683,N_9181,N_7671);
and U13684 (N_13684,N_7384,N_5208);
nor U13685 (N_13685,N_7038,N_7726);
nor U13686 (N_13686,N_8497,N_8029);
nand U13687 (N_13687,N_5762,N_5639);
nor U13688 (N_13688,N_6331,N_6285);
nor U13689 (N_13689,N_8247,N_8221);
and U13690 (N_13690,N_6001,N_8611);
xnor U13691 (N_13691,N_8352,N_5043);
and U13692 (N_13692,N_7503,N_6995);
nand U13693 (N_13693,N_6156,N_8547);
nor U13694 (N_13694,N_5786,N_9470);
xnor U13695 (N_13695,N_6923,N_7942);
xor U13696 (N_13696,N_8754,N_8805);
or U13697 (N_13697,N_9702,N_7123);
nand U13698 (N_13698,N_9426,N_7541);
or U13699 (N_13699,N_6072,N_9168);
nor U13700 (N_13700,N_7351,N_7237);
and U13701 (N_13701,N_8636,N_5741);
nand U13702 (N_13702,N_5013,N_5505);
and U13703 (N_13703,N_6074,N_7863);
or U13704 (N_13704,N_8481,N_8524);
nand U13705 (N_13705,N_7498,N_5004);
xnor U13706 (N_13706,N_9935,N_8811);
and U13707 (N_13707,N_8581,N_6781);
nor U13708 (N_13708,N_5311,N_6100);
nand U13709 (N_13709,N_9098,N_6901);
xor U13710 (N_13710,N_8757,N_9999);
nand U13711 (N_13711,N_5942,N_8553);
and U13712 (N_13712,N_7615,N_9196);
or U13713 (N_13713,N_9288,N_6137);
or U13714 (N_13714,N_9163,N_9259);
and U13715 (N_13715,N_9615,N_5264);
and U13716 (N_13716,N_6647,N_7853);
nor U13717 (N_13717,N_6622,N_7205);
nand U13718 (N_13718,N_9116,N_6055);
nand U13719 (N_13719,N_9601,N_5886);
xnor U13720 (N_13720,N_8450,N_5238);
xnor U13721 (N_13721,N_5047,N_8432);
nor U13722 (N_13722,N_5462,N_6330);
xnor U13723 (N_13723,N_9121,N_6750);
nor U13724 (N_13724,N_9975,N_8605);
nand U13725 (N_13725,N_5676,N_9993);
or U13726 (N_13726,N_5437,N_8362);
xnor U13727 (N_13727,N_9376,N_6701);
nor U13728 (N_13728,N_7678,N_9278);
xor U13729 (N_13729,N_9695,N_6568);
nor U13730 (N_13730,N_9692,N_7791);
or U13731 (N_13731,N_8026,N_6834);
or U13732 (N_13732,N_5780,N_8623);
xnor U13733 (N_13733,N_7154,N_8909);
or U13734 (N_13734,N_9160,N_6226);
and U13735 (N_13735,N_8066,N_6543);
xnor U13736 (N_13736,N_5987,N_7957);
xnor U13737 (N_13737,N_8810,N_8972);
nand U13738 (N_13738,N_6421,N_5278);
nand U13739 (N_13739,N_6418,N_8612);
and U13740 (N_13740,N_6157,N_8255);
or U13741 (N_13741,N_5095,N_7122);
or U13742 (N_13742,N_9127,N_5779);
or U13743 (N_13743,N_6860,N_7342);
xnor U13744 (N_13744,N_5736,N_9122);
nor U13745 (N_13745,N_8876,N_9749);
nor U13746 (N_13746,N_7500,N_9687);
nand U13747 (N_13747,N_8698,N_8747);
nand U13748 (N_13748,N_8436,N_8348);
xor U13749 (N_13749,N_6696,N_6363);
nand U13750 (N_13750,N_5888,N_9699);
or U13751 (N_13751,N_5073,N_7629);
or U13752 (N_13752,N_5624,N_7279);
and U13753 (N_13753,N_5027,N_8442);
nor U13754 (N_13754,N_9514,N_7114);
nor U13755 (N_13755,N_8763,N_6357);
and U13756 (N_13756,N_5617,N_6381);
nand U13757 (N_13757,N_6783,N_7786);
nor U13758 (N_13758,N_9674,N_6493);
nand U13759 (N_13759,N_6726,N_8807);
or U13760 (N_13760,N_9092,N_8064);
nor U13761 (N_13761,N_5103,N_9250);
nor U13762 (N_13762,N_5799,N_5897);
and U13763 (N_13763,N_7175,N_5422);
xor U13764 (N_13764,N_8686,N_8714);
or U13765 (N_13765,N_9813,N_7247);
xnor U13766 (N_13766,N_9069,N_7961);
or U13767 (N_13767,N_8997,N_5631);
and U13768 (N_13768,N_5247,N_5407);
nand U13769 (N_13769,N_5240,N_6781);
nand U13770 (N_13770,N_9739,N_9135);
and U13771 (N_13771,N_7142,N_9665);
xnor U13772 (N_13772,N_5965,N_6498);
nor U13773 (N_13773,N_9374,N_9462);
xor U13774 (N_13774,N_6359,N_7958);
nand U13775 (N_13775,N_6926,N_5709);
or U13776 (N_13776,N_9918,N_9186);
nand U13777 (N_13777,N_5286,N_7862);
xnor U13778 (N_13778,N_8076,N_7850);
xor U13779 (N_13779,N_8378,N_8494);
nand U13780 (N_13780,N_6242,N_5131);
or U13781 (N_13781,N_6593,N_9342);
nand U13782 (N_13782,N_5846,N_6344);
xnor U13783 (N_13783,N_8250,N_5305);
nor U13784 (N_13784,N_5040,N_7535);
or U13785 (N_13785,N_5709,N_5509);
or U13786 (N_13786,N_8068,N_8948);
and U13787 (N_13787,N_5742,N_9817);
nor U13788 (N_13788,N_5430,N_9553);
nand U13789 (N_13789,N_9288,N_6718);
and U13790 (N_13790,N_7715,N_7409);
nand U13791 (N_13791,N_8214,N_5862);
nand U13792 (N_13792,N_9513,N_6935);
and U13793 (N_13793,N_5150,N_9404);
xor U13794 (N_13794,N_8706,N_9090);
nand U13795 (N_13795,N_6284,N_7215);
or U13796 (N_13796,N_8058,N_9149);
or U13797 (N_13797,N_9119,N_6416);
nand U13798 (N_13798,N_5128,N_6850);
nand U13799 (N_13799,N_6303,N_9634);
xnor U13800 (N_13800,N_8327,N_6291);
or U13801 (N_13801,N_5691,N_8635);
or U13802 (N_13802,N_9673,N_6315);
xor U13803 (N_13803,N_5260,N_6685);
nor U13804 (N_13804,N_6591,N_9858);
xor U13805 (N_13805,N_8356,N_6551);
nor U13806 (N_13806,N_5809,N_9867);
xnor U13807 (N_13807,N_5152,N_6842);
and U13808 (N_13808,N_6897,N_5081);
or U13809 (N_13809,N_5757,N_6222);
nor U13810 (N_13810,N_6094,N_9471);
or U13811 (N_13811,N_9340,N_9414);
nand U13812 (N_13812,N_9907,N_5541);
nor U13813 (N_13813,N_8488,N_9612);
nand U13814 (N_13814,N_6279,N_6072);
nand U13815 (N_13815,N_5472,N_8172);
and U13816 (N_13816,N_9839,N_9810);
and U13817 (N_13817,N_6256,N_7925);
nand U13818 (N_13818,N_5751,N_5825);
and U13819 (N_13819,N_8292,N_9478);
nand U13820 (N_13820,N_7006,N_8396);
and U13821 (N_13821,N_6267,N_8123);
xnor U13822 (N_13822,N_6028,N_9238);
nor U13823 (N_13823,N_6098,N_8046);
nor U13824 (N_13824,N_6957,N_8621);
xnor U13825 (N_13825,N_9846,N_5102);
and U13826 (N_13826,N_6858,N_9781);
nor U13827 (N_13827,N_6525,N_9334);
or U13828 (N_13828,N_5462,N_8486);
xnor U13829 (N_13829,N_7864,N_7436);
nor U13830 (N_13830,N_5691,N_6660);
and U13831 (N_13831,N_8777,N_8291);
and U13832 (N_13832,N_8754,N_9501);
or U13833 (N_13833,N_6635,N_7198);
and U13834 (N_13834,N_5073,N_8659);
nand U13835 (N_13835,N_5571,N_9080);
and U13836 (N_13836,N_9376,N_7837);
and U13837 (N_13837,N_9324,N_6035);
and U13838 (N_13838,N_8987,N_6101);
and U13839 (N_13839,N_8578,N_7665);
nand U13840 (N_13840,N_6398,N_8679);
and U13841 (N_13841,N_7046,N_7145);
xor U13842 (N_13842,N_6428,N_8466);
nor U13843 (N_13843,N_5693,N_8335);
nor U13844 (N_13844,N_6740,N_9174);
nand U13845 (N_13845,N_8870,N_7814);
nand U13846 (N_13846,N_5443,N_6534);
and U13847 (N_13847,N_8981,N_7412);
xor U13848 (N_13848,N_5715,N_5179);
nor U13849 (N_13849,N_8844,N_8778);
nand U13850 (N_13850,N_7657,N_9726);
and U13851 (N_13851,N_7044,N_9765);
xnor U13852 (N_13852,N_6968,N_6439);
nor U13853 (N_13853,N_5853,N_7149);
xnor U13854 (N_13854,N_6534,N_9425);
nor U13855 (N_13855,N_5256,N_9025);
and U13856 (N_13856,N_7893,N_5728);
or U13857 (N_13857,N_5924,N_8575);
nor U13858 (N_13858,N_9676,N_8914);
xor U13859 (N_13859,N_8520,N_8282);
nand U13860 (N_13860,N_8169,N_8458);
xnor U13861 (N_13861,N_5893,N_7405);
nor U13862 (N_13862,N_6363,N_9248);
xnor U13863 (N_13863,N_9480,N_5980);
or U13864 (N_13864,N_6275,N_8213);
xnor U13865 (N_13865,N_6261,N_8000);
nand U13866 (N_13866,N_8882,N_9245);
nand U13867 (N_13867,N_9091,N_6179);
and U13868 (N_13868,N_7858,N_9392);
and U13869 (N_13869,N_9092,N_7843);
or U13870 (N_13870,N_6002,N_7160);
nor U13871 (N_13871,N_5600,N_6532);
and U13872 (N_13872,N_9955,N_5819);
or U13873 (N_13873,N_7164,N_8868);
xor U13874 (N_13874,N_6591,N_7238);
nor U13875 (N_13875,N_6645,N_7544);
or U13876 (N_13876,N_7063,N_9991);
or U13877 (N_13877,N_7414,N_6596);
nand U13878 (N_13878,N_6600,N_5637);
nor U13879 (N_13879,N_7161,N_9663);
or U13880 (N_13880,N_7201,N_8474);
nor U13881 (N_13881,N_5076,N_8202);
xnor U13882 (N_13882,N_7987,N_6674);
xnor U13883 (N_13883,N_5307,N_9419);
nor U13884 (N_13884,N_6400,N_5874);
xnor U13885 (N_13885,N_9155,N_7888);
xor U13886 (N_13886,N_8912,N_8314);
nand U13887 (N_13887,N_6510,N_8721);
nand U13888 (N_13888,N_8070,N_9789);
or U13889 (N_13889,N_6138,N_8461);
nand U13890 (N_13890,N_7626,N_5764);
nor U13891 (N_13891,N_7723,N_7489);
or U13892 (N_13892,N_5492,N_5983);
nand U13893 (N_13893,N_6144,N_5534);
nand U13894 (N_13894,N_5692,N_9693);
or U13895 (N_13895,N_9159,N_5149);
and U13896 (N_13896,N_9231,N_6097);
and U13897 (N_13897,N_9758,N_5808);
and U13898 (N_13898,N_5874,N_5810);
or U13899 (N_13899,N_6064,N_7397);
xor U13900 (N_13900,N_7267,N_6095);
and U13901 (N_13901,N_9236,N_5824);
xor U13902 (N_13902,N_9925,N_5312);
nor U13903 (N_13903,N_9916,N_9081);
xor U13904 (N_13904,N_9109,N_6855);
nand U13905 (N_13905,N_6888,N_8310);
and U13906 (N_13906,N_6521,N_9483);
or U13907 (N_13907,N_9587,N_6092);
nand U13908 (N_13908,N_7844,N_5545);
xor U13909 (N_13909,N_6319,N_7701);
or U13910 (N_13910,N_7326,N_7440);
nand U13911 (N_13911,N_9590,N_6582);
xnor U13912 (N_13912,N_7939,N_9493);
xor U13913 (N_13913,N_6100,N_6635);
xor U13914 (N_13914,N_8769,N_5587);
nor U13915 (N_13915,N_5493,N_7937);
or U13916 (N_13916,N_8909,N_9604);
and U13917 (N_13917,N_8899,N_5165);
nand U13918 (N_13918,N_8906,N_9213);
or U13919 (N_13919,N_8688,N_9961);
nand U13920 (N_13920,N_5118,N_9269);
or U13921 (N_13921,N_6218,N_5778);
nor U13922 (N_13922,N_9812,N_7723);
and U13923 (N_13923,N_7546,N_8739);
nand U13924 (N_13924,N_5168,N_5027);
nand U13925 (N_13925,N_9362,N_8058);
nor U13926 (N_13926,N_5316,N_8132);
and U13927 (N_13927,N_9901,N_5970);
or U13928 (N_13928,N_9408,N_6903);
and U13929 (N_13929,N_8092,N_9756);
and U13930 (N_13930,N_5944,N_9905);
or U13931 (N_13931,N_6536,N_9951);
and U13932 (N_13932,N_9373,N_5186);
nand U13933 (N_13933,N_8932,N_9746);
nand U13934 (N_13934,N_8314,N_8680);
xor U13935 (N_13935,N_6757,N_7051);
and U13936 (N_13936,N_6253,N_6800);
or U13937 (N_13937,N_6116,N_9115);
nor U13938 (N_13938,N_7053,N_8705);
nand U13939 (N_13939,N_8764,N_6329);
or U13940 (N_13940,N_5596,N_9825);
nand U13941 (N_13941,N_7117,N_8602);
or U13942 (N_13942,N_9656,N_6592);
nor U13943 (N_13943,N_7949,N_7632);
or U13944 (N_13944,N_9591,N_9876);
and U13945 (N_13945,N_7274,N_8296);
or U13946 (N_13946,N_5195,N_9467);
nand U13947 (N_13947,N_5399,N_6807);
xor U13948 (N_13948,N_8416,N_6631);
xnor U13949 (N_13949,N_8121,N_8596);
xor U13950 (N_13950,N_5269,N_6332);
or U13951 (N_13951,N_8390,N_6958);
xor U13952 (N_13952,N_8044,N_7288);
xnor U13953 (N_13953,N_9228,N_7530);
nand U13954 (N_13954,N_5814,N_5145);
nand U13955 (N_13955,N_8033,N_8292);
nor U13956 (N_13956,N_8916,N_9641);
nor U13957 (N_13957,N_6060,N_9255);
and U13958 (N_13958,N_5332,N_7311);
and U13959 (N_13959,N_8215,N_6471);
and U13960 (N_13960,N_9734,N_7921);
and U13961 (N_13961,N_7063,N_7855);
xor U13962 (N_13962,N_6437,N_7246);
nand U13963 (N_13963,N_8862,N_7470);
or U13964 (N_13964,N_8960,N_5426);
or U13965 (N_13965,N_9127,N_7455);
nand U13966 (N_13966,N_6385,N_9689);
xnor U13967 (N_13967,N_5324,N_6534);
xor U13968 (N_13968,N_5705,N_5508);
nor U13969 (N_13969,N_8577,N_7288);
xnor U13970 (N_13970,N_5427,N_9276);
or U13971 (N_13971,N_9049,N_5380);
nand U13972 (N_13972,N_6410,N_8327);
nand U13973 (N_13973,N_7750,N_7538);
nor U13974 (N_13974,N_6439,N_6128);
or U13975 (N_13975,N_7835,N_9039);
or U13976 (N_13976,N_7309,N_6809);
and U13977 (N_13977,N_7195,N_8408);
or U13978 (N_13978,N_6944,N_8028);
or U13979 (N_13979,N_5395,N_7530);
xnor U13980 (N_13980,N_5507,N_6966);
or U13981 (N_13981,N_8642,N_8426);
and U13982 (N_13982,N_9924,N_9419);
nand U13983 (N_13983,N_5703,N_5627);
and U13984 (N_13984,N_7732,N_8351);
nor U13985 (N_13985,N_5185,N_8135);
or U13986 (N_13986,N_8142,N_7190);
or U13987 (N_13987,N_9149,N_8293);
nand U13988 (N_13988,N_8671,N_8971);
nand U13989 (N_13989,N_9200,N_5527);
nor U13990 (N_13990,N_6239,N_6622);
or U13991 (N_13991,N_7810,N_8443);
nand U13992 (N_13992,N_8323,N_7267);
nand U13993 (N_13993,N_7479,N_6264);
xor U13994 (N_13994,N_6324,N_8717);
xnor U13995 (N_13995,N_5704,N_5941);
nor U13996 (N_13996,N_8076,N_8163);
xor U13997 (N_13997,N_5030,N_6525);
nor U13998 (N_13998,N_7030,N_5261);
nor U13999 (N_13999,N_5603,N_6419);
or U14000 (N_14000,N_8681,N_9553);
nand U14001 (N_14001,N_7616,N_5550);
or U14002 (N_14002,N_8591,N_9553);
and U14003 (N_14003,N_8238,N_8040);
and U14004 (N_14004,N_7351,N_5615);
or U14005 (N_14005,N_9137,N_9393);
and U14006 (N_14006,N_7349,N_6349);
nand U14007 (N_14007,N_8105,N_5561);
or U14008 (N_14008,N_7493,N_9325);
xor U14009 (N_14009,N_5498,N_6549);
xor U14010 (N_14010,N_7800,N_6990);
nand U14011 (N_14011,N_5845,N_5462);
nor U14012 (N_14012,N_7534,N_9767);
nand U14013 (N_14013,N_8876,N_8667);
nand U14014 (N_14014,N_7175,N_6425);
nand U14015 (N_14015,N_9700,N_8114);
nand U14016 (N_14016,N_9840,N_7306);
and U14017 (N_14017,N_7606,N_7013);
nor U14018 (N_14018,N_7439,N_8124);
or U14019 (N_14019,N_7355,N_5326);
xor U14020 (N_14020,N_6640,N_9416);
or U14021 (N_14021,N_5811,N_6011);
nor U14022 (N_14022,N_8460,N_6320);
and U14023 (N_14023,N_7198,N_9906);
and U14024 (N_14024,N_6963,N_7573);
nand U14025 (N_14025,N_7656,N_8129);
and U14026 (N_14026,N_8336,N_5784);
nor U14027 (N_14027,N_9577,N_9875);
and U14028 (N_14028,N_6340,N_9415);
or U14029 (N_14029,N_7161,N_7921);
and U14030 (N_14030,N_7342,N_7242);
or U14031 (N_14031,N_5308,N_7198);
or U14032 (N_14032,N_5370,N_5149);
xor U14033 (N_14033,N_5046,N_6556);
nand U14034 (N_14034,N_7820,N_5545);
or U14035 (N_14035,N_8103,N_7361);
xnor U14036 (N_14036,N_8671,N_9798);
nand U14037 (N_14037,N_9861,N_9628);
and U14038 (N_14038,N_6776,N_8458);
xnor U14039 (N_14039,N_7548,N_7364);
nor U14040 (N_14040,N_9309,N_9907);
xor U14041 (N_14041,N_6481,N_6076);
nand U14042 (N_14042,N_9481,N_8467);
nor U14043 (N_14043,N_7792,N_5187);
or U14044 (N_14044,N_9342,N_8829);
or U14045 (N_14045,N_7678,N_6464);
xnor U14046 (N_14046,N_7310,N_6912);
nor U14047 (N_14047,N_8094,N_6047);
and U14048 (N_14048,N_7716,N_5109);
nor U14049 (N_14049,N_9280,N_7982);
and U14050 (N_14050,N_9405,N_9069);
xor U14051 (N_14051,N_8873,N_9071);
nor U14052 (N_14052,N_7693,N_7488);
nand U14053 (N_14053,N_8548,N_5114);
and U14054 (N_14054,N_6454,N_6509);
nand U14055 (N_14055,N_8859,N_6387);
or U14056 (N_14056,N_9468,N_8056);
or U14057 (N_14057,N_5612,N_6292);
nand U14058 (N_14058,N_6860,N_7440);
xnor U14059 (N_14059,N_5800,N_7303);
nand U14060 (N_14060,N_7104,N_9137);
xnor U14061 (N_14061,N_5690,N_5912);
and U14062 (N_14062,N_9457,N_8277);
nor U14063 (N_14063,N_9869,N_5011);
and U14064 (N_14064,N_5699,N_8230);
nor U14065 (N_14065,N_5228,N_6392);
and U14066 (N_14066,N_7346,N_7646);
and U14067 (N_14067,N_6826,N_9870);
or U14068 (N_14068,N_7814,N_6440);
nand U14069 (N_14069,N_5175,N_7828);
xnor U14070 (N_14070,N_8387,N_7955);
and U14071 (N_14071,N_8967,N_5565);
xnor U14072 (N_14072,N_7625,N_6726);
and U14073 (N_14073,N_6072,N_9406);
xor U14074 (N_14074,N_6730,N_8128);
nand U14075 (N_14075,N_8706,N_6698);
nand U14076 (N_14076,N_8931,N_9489);
xnor U14077 (N_14077,N_6863,N_9661);
or U14078 (N_14078,N_5251,N_5357);
and U14079 (N_14079,N_8500,N_6095);
nor U14080 (N_14080,N_8903,N_8946);
nand U14081 (N_14081,N_8726,N_8969);
nand U14082 (N_14082,N_5813,N_5796);
nor U14083 (N_14083,N_9112,N_8507);
nand U14084 (N_14084,N_6474,N_7269);
and U14085 (N_14085,N_6515,N_8038);
and U14086 (N_14086,N_7682,N_7994);
nor U14087 (N_14087,N_6951,N_9312);
and U14088 (N_14088,N_5422,N_6168);
nor U14089 (N_14089,N_6373,N_8611);
nor U14090 (N_14090,N_6416,N_5158);
nand U14091 (N_14091,N_5890,N_8762);
nand U14092 (N_14092,N_9257,N_6715);
and U14093 (N_14093,N_9505,N_9007);
xor U14094 (N_14094,N_9867,N_8499);
nand U14095 (N_14095,N_5410,N_6026);
or U14096 (N_14096,N_6237,N_5564);
and U14097 (N_14097,N_7797,N_6731);
and U14098 (N_14098,N_8503,N_5600);
or U14099 (N_14099,N_5258,N_9054);
or U14100 (N_14100,N_5306,N_6430);
nand U14101 (N_14101,N_8505,N_7610);
nand U14102 (N_14102,N_7873,N_9461);
xnor U14103 (N_14103,N_5878,N_5336);
nand U14104 (N_14104,N_9959,N_6502);
and U14105 (N_14105,N_8982,N_6480);
or U14106 (N_14106,N_9918,N_9303);
nand U14107 (N_14107,N_7699,N_8249);
nor U14108 (N_14108,N_5304,N_6014);
nor U14109 (N_14109,N_6881,N_9762);
nor U14110 (N_14110,N_7754,N_5194);
nand U14111 (N_14111,N_5030,N_7320);
nor U14112 (N_14112,N_6509,N_9519);
and U14113 (N_14113,N_9385,N_5658);
nor U14114 (N_14114,N_6836,N_6814);
xor U14115 (N_14115,N_6573,N_7735);
and U14116 (N_14116,N_6120,N_7298);
or U14117 (N_14117,N_8754,N_9102);
or U14118 (N_14118,N_8748,N_9527);
and U14119 (N_14119,N_7023,N_8102);
nor U14120 (N_14120,N_8212,N_9465);
nand U14121 (N_14121,N_9683,N_6677);
nor U14122 (N_14122,N_9786,N_7478);
xor U14123 (N_14123,N_5128,N_9369);
nand U14124 (N_14124,N_8782,N_8930);
nor U14125 (N_14125,N_8144,N_5684);
nor U14126 (N_14126,N_5570,N_6829);
xor U14127 (N_14127,N_8644,N_7333);
nor U14128 (N_14128,N_9012,N_7155);
and U14129 (N_14129,N_7957,N_9957);
or U14130 (N_14130,N_9817,N_7736);
nand U14131 (N_14131,N_6776,N_8046);
xnor U14132 (N_14132,N_6116,N_9424);
nor U14133 (N_14133,N_7018,N_8563);
xor U14134 (N_14134,N_6864,N_9148);
or U14135 (N_14135,N_7172,N_7125);
or U14136 (N_14136,N_6412,N_9391);
nand U14137 (N_14137,N_8610,N_9284);
or U14138 (N_14138,N_7519,N_9317);
or U14139 (N_14139,N_6396,N_7696);
and U14140 (N_14140,N_8351,N_7674);
xnor U14141 (N_14141,N_7333,N_7645);
or U14142 (N_14142,N_9258,N_5416);
or U14143 (N_14143,N_7716,N_5841);
and U14144 (N_14144,N_8732,N_9769);
or U14145 (N_14145,N_8110,N_9056);
xnor U14146 (N_14146,N_8136,N_8386);
nand U14147 (N_14147,N_8731,N_7327);
xor U14148 (N_14148,N_9351,N_5765);
and U14149 (N_14149,N_9672,N_8976);
xnor U14150 (N_14150,N_5115,N_5255);
or U14151 (N_14151,N_5659,N_5685);
xnor U14152 (N_14152,N_9345,N_6855);
nor U14153 (N_14153,N_6800,N_6465);
or U14154 (N_14154,N_5850,N_9223);
nand U14155 (N_14155,N_8870,N_9597);
nor U14156 (N_14156,N_7642,N_5374);
nand U14157 (N_14157,N_5536,N_6185);
nand U14158 (N_14158,N_8499,N_6306);
and U14159 (N_14159,N_7392,N_7149);
nand U14160 (N_14160,N_6793,N_6493);
xor U14161 (N_14161,N_5020,N_6454);
and U14162 (N_14162,N_8220,N_6445);
or U14163 (N_14163,N_5334,N_9774);
nand U14164 (N_14164,N_9162,N_6652);
and U14165 (N_14165,N_8588,N_6102);
nor U14166 (N_14166,N_7198,N_6047);
and U14167 (N_14167,N_6531,N_8179);
xnor U14168 (N_14168,N_8324,N_6214);
nor U14169 (N_14169,N_6085,N_9995);
nand U14170 (N_14170,N_6367,N_5788);
nand U14171 (N_14171,N_7565,N_8360);
nand U14172 (N_14172,N_6191,N_7523);
and U14173 (N_14173,N_9080,N_6308);
or U14174 (N_14174,N_9428,N_9128);
xnor U14175 (N_14175,N_7330,N_5449);
nand U14176 (N_14176,N_5548,N_9381);
or U14177 (N_14177,N_9142,N_6407);
nand U14178 (N_14178,N_6709,N_8820);
nand U14179 (N_14179,N_6465,N_9753);
nand U14180 (N_14180,N_9320,N_5867);
or U14181 (N_14181,N_5125,N_5854);
nor U14182 (N_14182,N_9839,N_8454);
xnor U14183 (N_14183,N_8223,N_8700);
nor U14184 (N_14184,N_6974,N_8269);
nand U14185 (N_14185,N_9623,N_7979);
nand U14186 (N_14186,N_5263,N_6163);
nand U14187 (N_14187,N_9528,N_9789);
nand U14188 (N_14188,N_7444,N_8363);
nand U14189 (N_14189,N_9605,N_5319);
and U14190 (N_14190,N_8810,N_5950);
or U14191 (N_14191,N_5189,N_9499);
nor U14192 (N_14192,N_7880,N_7599);
nor U14193 (N_14193,N_6516,N_8217);
or U14194 (N_14194,N_7142,N_7609);
and U14195 (N_14195,N_6181,N_7894);
and U14196 (N_14196,N_9864,N_7996);
xnor U14197 (N_14197,N_5298,N_8237);
or U14198 (N_14198,N_8890,N_5677);
xor U14199 (N_14199,N_5008,N_5932);
nand U14200 (N_14200,N_7874,N_6583);
nand U14201 (N_14201,N_6936,N_6649);
or U14202 (N_14202,N_5422,N_7243);
xor U14203 (N_14203,N_7391,N_6787);
xor U14204 (N_14204,N_9608,N_7941);
and U14205 (N_14205,N_6208,N_8724);
or U14206 (N_14206,N_9591,N_6014);
and U14207 (N_14207,N_6405,N_6963);
and U14208 (N_14208,N_8802,N_8732);
and U14209 (N_14209,N_8997,N_7478);
nor U14210 (N_14210,N_7857,N_6381);
nand U14211 (N_14211,N_6125,N_8670);
or U14212 (N_14212,N_9043,N_8416);
xnor U14213 (N_14213,N_9408,N_8004);
xnor U14214 (N_14214,N_6755,N_6159);
nand U14215 (N_14215,N_9731,N_9306);
nor U14216 (N_14216,N_7848,N_9186);
and U14217 (N_14217,N_5952,N_8678);
nor U14218 (N_14218,N_8297,N_6542);
and U14219 (N_14219,N_7850,N_8886);
nor U14220 (N_14220,N_8119,N_7212);
nand U14221 (N_14221,N_5244,N_8756);
or U14222 (N_14222,N_7907,N_6190);
nand U14223 (N_14223,N_5724,N_5406);
nand U14224 (N_14224,N_6184,N_8007);
nor U14225 (N_14225,N_8375,N_8335);
nand U14226 (N_14226,N_8128,N_5539);
nor U14227 (N_14227,N_6541,N_5990);
or U14228 (N_14228,N_5350,N_8209);
nor U14229 (N_14229,N_5562,N_9682);
or U14230 (N_14230,N_6618,N_6257);
and U14231 (N_14231,N_7700,N_8480);
or U14232 (N_14232,N_7153,N_5439);
nand U14233 (N_14233,N_7419,N_6491);
and U14234 (N_14234,N_5080,N_9990);
nand U14235 (N_14235,N_6548,N_5052);
and U14236 (N_14236,N_8728,N_5789);
and U14237 (N_14237,N_9268,N_7631);
xnor U14238 (N_14238,N_7613,N_7748);
and U14239 (N_14239,N_6838,N_9844);
nor U14240 (N_14240,N_8538,N_8940);
nand U14241 (N_14241,N_6333,N_8722);
nor U14242 (N_14242,N_8638,N_8501);
or U14243 (N_14243,N_9335,N_8445);
nand U14244 (N_14244,N_8065,N_5509);
nand U14245 (N_14245,N_5709,N_6729);
nand U14246 (N_14246,N_7122,N_5030);
and U14247 (N_14247,N_9211,N_6522);
xnor U14248 (N_14248,N_5473,N_8764);
or U14249 (N_14249,N_6973,N_7000);
nand U14250 (N_14250,N_9325,N_6522);
nor U14251 (N_14251,N_9305,N_8271);
nor U14252 (N_14252,N_6614,N_6544);
xor U14253 (N_14253,N_8350,N_7943);
xnor U14254 (N_14254,N_9904,N_9437);
nand U14255 (N_14255,N_8286,N_8935);
or U14256 (N_14256,N_8920,N_9649);
and U14257 (N_14257,N_9290,N_9611);
nand U14258 (N_14258,N_7515,N_6799);
or U14259 (N_14259,N_5773,N_6346);
or U14260 (N_14260,N_8649,N_5848);
xor U14261 (N_14261,N_8157,N_8694);
nor U14262 (N_14262,N_7322,N_8970);
xnor U14263 (N_14263,N_6996,N_6510);
nor U14264 (N_14264,N_7953,N_6767);
xnor U14265 (N_14265,N_6501,N_5520);
or U14266 (N_14266,N_7643,N_8427);
xor U14267 (N_14267,N_9822,N_6822);
xnor U14268 (N_14268,N_9323,N_5630);
nand U14269 (N_14269,N_8076,N_9040);
or U14270 (N_14270,N_6603,N_5968);
or U14271 (N_14271,N_7148,N_9672);
nand U14272 (N_14272,N_5638,N_6803);
and U14273 (N_14273,N_7081,N_8215);
and U14274 (N_14274,N_9336,N_7578);
or U14275 (N_14275,N_7481,N_6418);
and U14276 (N_14276,N_5158,N_8325);
or U14277 (N_14277,N_6018,N_7390);
or U14278 (N_14278,N_6623,N_9975);
nand U14279 (N_14279,N_8493,N_8746);
xor U14280 (N_14280,N_9656,N_5479);
or U14281 (N_14281,N_6085,N_5506);
xor U14282 (N_14282,N_9451,N_6145);
or U14283 (N_14283,N_5680,N_8084);
or U14284 (N_14284,N_8032,N_5786);
nor U14285 (N_14285,N_8263,N_7901);
xnor U14286 (N_14286,N_6932,N_5816);
nor U14287 (N_14287,N_6722,N_6833);
and U14288 (N_14288,N_6869,N_6043);
and U14289 (N_14289,N_9320,N_7781);
and U14290 (N_14290,N_6030,N_8791);
nor U14291 (N_14291,N_8622,N_7427);
nand U14292 (N_14292,N_6412,N_6844);
nand U14293 (N_14293,N_8100,N_6243);
xnor U14294 (N_14294,N_7804,N_9483);
nand U14295 (N_14295,N_8702,N_9128);
and U14296 (N_14296,N_5712,N_7203);
or U14297 (N_14297,N_5264,N_9144);
nor U14298 (N_14298,N_6024,N_6894);
nor U14299 (N_14299,N_5085,N_7412);
xnor U14300 (N_14300,N_9075,N_5283);
or U14301 (N_14301,N_6054,N_7142);
nand U14302 (N_14302,N_8503,N_7926);
xor U14303 (N_14303,N_7481,N_5209);
and U14304 (N_14304,N_9604,N_5653);
xor U14305 (N_14305,N_5120,N_8420);
nor U14306 (N_14306,N_8901,N_5459);
and U14307 (N_14307,N_8582,N_9512);
nand U14308 (N_14308,N_7185,N_9756);
or U14309 (N_14309,N_6738,N_5465);
xor U14310 (N_14310,N_7865,N_7569);
nand U14311 (N_14311,N_6835,N_8250);
nand U14312 (N_14312,N_9530,N_6910);
xnor U14313 (N_14313,N_5071,N_8120);
nand U14314 (N_14314,N_8348,N_8362);
or U14315 (N_14315,N_7712,N_6621);
or U14316 (N_14316,N_5710,N_9674);
nand U14317 (N_14317,N_9669,N_8529);
and U14318 (N_14318,N_9522,N_5239);
or U14319 (N_14319,N_5631,N_6613);
or U14320 (N_14320,N_7003,N_7006);
or U14321 (N_14321,N_5570,N_6479);
and U14322 (N_14322,N_7622,N_5133);
nor U14323 (N_14323,N_5783,N_6100);
or U14324 (N_14324,N_8932,N_7145);
nand U14325 (N_14325,N_8068,N_7385);
xor U14326 (N_14326,N_9942,N_5747);
nand U14327 (N_14327,N_5279,N_6382);
and U14328 (N_14328,N_6743,N_9374);
nand U14329 (N_14329,N_9633,N_5248);
or U14330 (N_14330,N_8182,N_9064);
nand U14331 (N_14331,N_9749,N_9298);
and U14332 (N_14332,N_7938,N_5371);
or U14333 (N_14333,N_7938,N_6818);
nand U14334 (N_14334,N_5165,N_7716);
nor U14335 (N_14335,N_5223,N_7956);
nand U14336 (N_14336,N_5730,N_9692);
nor U14337 (N_14337,N_8607,N_7418);
and U14338 (N_14338,N_6038,N_5264);
xor U14339 (N_14339,N_7757,N_8351);
and U14340 (N_14340,N_8263,N_8140);
nor U14341 (N_14341,N_9307,N_5306);
and U14342 (N_14342,N_7467,N_8646);
nor U14343 (N_14343,N_7963,N_9020);
or U14344 (N_14344,N_8459,N_8583);
or U14345 (N_14345,N_5167,N_6487);
nor U14346 (N_14346,N_5396,N_6482);
xnor U14347 (N_14347,N_9312,N_9904);
xor U14348 (N_14348,N_5823,N_7596);
nor U14349 (N_14349,N_5299,N_5862);
and U14350 (N_14350,N_7423,N_6232);
nor U14351 (N_14351,N_6819,N_5692);
and U14352 (N_14352,N_6418,N_7783);
xnor U14353 (N_14353,N_9187,N_5636);
nand U14354 (N_14354,N_5116,N_9410);
or U14355 (N_14355,N_7309,N_6416);
nand U14356 (N_14356,N_5225,N_5310);
xnor U14357 (N_14357,N_6296,N_9268);
xor U14358 (N_14358,N_5370,N_7826);
nand U14359 (N_14359,N_8742,N_9149);
and U14360 (N_14360,N_9233,N_7879);
nor U14361 (N_14361,N_6364,N_9295);
nor U14362 (N_14362,N_6431,N_9994);
nor U14363 (N_14363,N_9897,N_7394);
and U14364 (N_14364,N_5404,N_5510);
and U14365 (N_14365,N_6656,N_7549);
nand U14366 (N_14366,N_7735,N_6140);
and U14367 (N_14367,N_8613,N_6913);
or U14368 (N_14368,N_8320,N_5850);
and U14369 (N_14369,N_6864,N_5772);
nand U14370 (N_14370,N_8264,N_9397);
or U14371 (N_14371,N_8991,N_5906);
nand U14372 (N_14372,N_5188,N_6113);
xor U14373 (N_14373,N_8313,N_5183);
or U14374 (N_14374,N_8779,N_5626);
nor U14375 (N_14375,N_5515,N_7848);
xnor U14376 (N_14376,N_8607,N_8224);
nor U14377 (N_14377,N_9516,N_8735);
nor U14378 (N_14378,N_5022,N_6719);
xor U14379 (N_14379,N_6791,N_9410);
and U14380 (N_14380,N_6483,N_7600);
xor U14381 (N_14381,N_6113,N_7454);
and U14382 (N_14382,N_7859,N_8328);
xor U14383 (N_14383,N_8951,N_9957);
nor U14384 (N_14384,N_7640,N_6374);
and U14385 (N_14385,N_5256,N_9567);
nor U14386 (N_14386,N_8327,N_9507);
xnor U14387 (N_14387,N_5160,N_9246);
and U14388 (N_14388,N_8185,N_5357);
or U14389 (N_14389,N_5807,N_9310);
and U14390 (N_14390,N_7573,N_9228);
or U14391 (N_14391,N_9475,N_6323);
nand U14392 (N_14392,N_7515,N_5495);
or U14393 (N_14393,N_9236,N_7500);
nand U14394 (N_14394,N_5671,N_6463);
nor U14395 (N_14395,N_5643,N_5679);
and U14396 (N_14396,N_6735,N_6037);
nand U14397 (N_14397,N_8753,N_9779);
or U14398 (N_14398,N_5015,N_6968);
xor U14399 (N_14399,N_7275,N_5851);
nor U14400 (N_14400,N_6766,N_9807);
xor U14401 (N_14401,N_6608,N_8624);
nor U14402 (N_14402,N_8026,N_6882);
nor U14403 (N_14403,N_9568,N_6383);
and U14404 (N_14404,N_5223,N_8611);
or U14405 (N_14405,N_9827,N_9433);
xor U14406 (N_14406,N_6724,N_6813);
or U14407 (N_14407,N_7792,N_7771);
nor U14408 (N_14408,N_8123,N_8885);
or U14409 (N_14409,N_6032,N_5523);
and U14410 (N_14410,N_8026,N_7001);
and U14411 (N_14411,N_5044,N_9311);
and U14412 (N_14412,N_7448,N_6308);
or U14413 (N_14413,N_7935,N_7644);
nor U14414 (N_14414,N_7677,N_8149);
nand U14415 (N_14415,N_8413,N_7853);
or U14416 (N_14416,N_6703,N_6875);
or U14417 (N_14417,N_9286,N_9204);
nor U14418 (N_14418,N_6536,N_9145);
nor U14419 (N_14419,N_6651,N_5950);
xnor U14420 (N_14420,N_8411,N_7826);
nand U14421 (N_14421,N_5004,N_5890);
or U14422 (N_14422,N_9816,N_8280);
and U14423 (N_14423,N_8302,N_9460);
nor U14424 (N_14424,N_8646,N_6031);
xnor U14425 (N_14425,N_6693,N_7601);
xnor U14426 (N_14426,N_7380,N_7116);
or U14427 (N_14427,N_6884,N_6173);
xor U14428 (N_14428,N_9306,N_7376);
or U14429 (N_14429,N_8371,N_7696);
and U14430 (N_14430,N_8296,N_9005);
nand U14431 (N_14431,N_9118,N_8402);
or U14432 (N_14432,N_6864,N_6527);
nand U14433 (N_14433,N_9699,N_9208);
xor U14434 (N_14434,N_6023,N_7365);
and U14435 (N_14435,N_5102,N_9967);
xor U14436 (N_14436,N_8259,N_6025);
and U14437 (N_14437,N_7366,N_9996);
and U14438 (N_14438,N_5199,N_8369);
and U14439 (N_14439,N_6664,N_8537);
and U14440 (N_14440,N_5682,N_6985);
and U14441 (N_14441,N_9976,N_5196);
xor U14442 (N_14442,N_8144,N_8085);
and U14443 (N_14443,N_5413,N_6401);
nor U14444 (N_14444,N_7641,N_5143);
nor U14445 (N_14445,N_9324,N_9689);
xnor U14446 (N_14446,N_6577,N_7747);
nor U14447 (N_14447,N_5449,N_7482);
and U14448 (N_14448,N_9391,N_7160);
nor U14449 (N_14449,N_8808,N_8474);
nor U14450 (N_14450,N_5156,N_5444);
nor U14451 (N_14451,N_9463,N_8385);
xnor U14452 (N_14452,N_8128,N_8948);
xor U14453 (N_14453,N_5494,N_7459);
nand U14454 (N_14454,N_9572,N_9983);
xnor U14455 (N_14455,N_9877,N_6061);
nand U14456 (N_14456,N_6009,N_6962);
and U14457 (N_14457,N_7037,N_6243);
or U14458 (N_14458,N_6580,N_7857);
nor U14459 (N_14459,N_9014,N_8239);
and U14460 (N_14460,N_7199,N_5090);
or U14461 (N_14461,N_8443,N_8751);
or U14462 (N_14462,N_6072,N_5167);
nor U14463 (N_14463,N_8174,N_6424);
xor U14464 (N_14464,N_6607,N_5665);
and U14465 (N_14465,N_6428,N_8764);
nand U14466 (N_14466,N_5298,N_9235);
nand U14467 (N_14467,N_6690,N_6789);
nand U14468 (N_14468,N_6432,N_7970);
nor U14469 (N_14469,N_7128,N_7941);
and U14470 (N_14470,N_5341,N_6637);
nor U14471 (N_14471,N_9311,N_8653);
nand U14472 (N_14472,N_6799,N_9437);
or U14473 (N_14473,N_9840,N_6374);
nand U14474 (N_14474,N_7418,N_6774);
and U14475 (N_14475,N_6481,N_5360);
or U14476 (N_14476,N_6002,N_8595);
and U14477 (N_14477,N_7906,N_6812);
or U14478 (N_14478,N_5733,N_5262);
nor U14479 (N_14479,N_5458,N_7958);
nor U14480 (N_14480,N_8676,N_7878);
and U14481 (N_14481,N_8077,N_5245);
nor U14482 (N_14482,N_8137,N_8811);
nor U14483 (N_14483,N_5298,N_5596);
xnor U14484 (N_14484,N_5250,N_5119);
and U14485 (N_14485,N_5711,N_9992);
nor U14486 (N_14486,N_7745,N_7610);
or U14487 (N_14487,N_7112,N_6604);
xnor U14488 (N_14488,N_9065,N_9922);
nor U14489 (N_14489,N_9639,N_5114);
nor U14490 (N_14490,N_7832,N_6258);
xnor U14491 (N_14491,N_6797,N_8570);
nor U14492 (N_14492,N_6456,N_6072);
nand U14493 (N_14493,N_6825,N_7816);
or U14494 (N_14494,N_6337,N_7066);
nand U14495 (N_14495,N_9276,N_8184);
xnor U14496 (N_14496,N_6166,N_7520);
and U14497 (N_14497,N_6848,N_7122);
nand U14498 (N_14498,N_9756,N_7462);
or U14499 (N_14499,N_7901,N_8872);
nand U14500 (N_14500,N_5793,N_7143);
nand U14501 (N_14501,N_8720,N_6403);
xor U14502 (N_14502,N_5026,N_9497);
and U14503 (N_14503,N_9222,N_8898);
and U14504 (N_14504,N_5096,N_5612);
nand U14505 (N_14505,N_9797,N_5186);
and U14506 (N_14506,N_6424,N_5885);
or U14507 (N_14507,N_5587,N_8218);
xnor U14508 (N_14508,N_8873,N_8652);
nand U14509 (N_14509,N_6349,N_5895);
nand U14510 (N_14510,N_9695,N_8917);
xnor U14511 (N_14511,N_5403,N_5961);
nor U14512 (N_14512,N_8467,N_9417);
nand U14513 (N_14513,N_5576,N_9777);
or U14514 (N_14514,N_8249,N_5609);
nor U14515 (N_14515,N_8668,N_8113);
or U14516 (N_14516,N_7478,N_7602);
and U14517 (N_14517,N_6672,N_9916);
xnor U14518 (N_14518,N_5642,N_8992);
xor U14519 (N_14519,N_7433,N_9549);
nand U14520 (N_14520,N_9925,N_7185);
and U14521 (N_14521,N_7135,N_7575);
and U14522 (N_14522,N_9292,N_6497);
and U14523 (N_14523,N_6761,N_5430);
and U14524 (N_14524,N_7365,N_7480);
or U14525 (N_14525,N_6002,N_9268);
xnor U14526 (N_14526,N_9387,N_9267);
and U14527 (N_14527,N_9950,N_5413);
or U14528 (N_14528,N_8274,N_6224);
xor U14529 (N_14529,N_5364,N_5184);
nor U14530 (N_14530,N_7386,N_7366);
and U14531 (N_14531,N_8695,N_8039);
or U14532 (N_14532,N_9238,N_8981);
nor U14533 (N_14533,N_9367,N_7410);
nand U14534 (N_14534,N_8024,N_9670);
and U14535 (N_14535,N_8411,N_7943);
xor U14536 (N_14536,N_7870,N_7418);
nand U14537 (N_14537,N_6355,N_6647);
and U14538 (N_14538,N_5808,N_7863);
nor U14539 (N_14539,N_9690,N_7366);
or U14540 (N_14540,N_5339,N_7097);
nand U14541 (N_14541,N_9906,N_9027);
or U14542 (N_14542,N_8183,N_6297);
nand U14543 (N_14543,N_5694,N_9422);
xor U14544 (N_14544,N_5213,N_6547);
or U14545 (N_14545,N_6502,N_7911);
nor U14546 (N_14546,N_8172,N_8878);
or U14547 (N_14547,N_7976,N_5679);
or U14548 (N_14548,N_8265,N_7701);
or U14549 (N_14549,N_9104,N_6448);
nand U14550 (N_14550,N_8976,N_9971);
or U14551 (N_14551,N_5305,N_8175);
or U14552 (N_14552,N_5489,N_8640);
xor U14553 (N_14553,N_7309,N_7022);
xor U14554 (N_14554,N_9792,N_6518);
nor U14555 (N_14555,N_6153,N_6844);
xor U14556 (N_14556,N_9997,N_9818);
or U14557 (N_14557,N_9507,N_7380);
or U14558 (N_14558,N_5211,N_9201);
xor U14559 (N_14559,N_9489,N_5277);
xnor U14560 (N_14560,N_5227,N_6497);
nand U14561 (N_14561,N_7227,N_5126);
nand U14562 (N_14562,N_7953,N_7785);
or U14563 (N_14563,N_9844,N_5953);
or U14564 (N_14564,N_7849,N_6378);
and U14565 (N_14565,N_9005,N_5238);
and U14566 (N_14566,N_9163,N_5958);
nor U14567 (N_14567,N_6800,N_7386);
and U14568 (N_14568,N_8055,N_6263);
or U14569 (N_14569,N_5074,N_8593);
and U14570 (N_14570,N_7995,N_8431);
xnor U14571 (N_14571,N_8473,N_7303);
xor U14572 (N_14572,N_6940,N_6727);
nor U14573 (N_14573,N_5329,N_6317);
or U14574 (N_14574,N_9209,N_5713);
nor U14575 (N_14575,N_5801,N_6311);
nand U14576 (N_14576,N_6797,N_9437);
xnor U14577 (N_14577,N_9160,N_6723);
nand U14578 (N_14578,N_6633,N_7508);
xnor U14579 (N_14579,N_6089,N_7565);
or U14580 (N_14580,N_7340,N_7796);
or U14581 (N_14581,N_6290,N_8087);
or U14582 (N_14582,N_9376,N_6569);
or U14583 (N_14583,N_5541,N_5267);
nand U14584 (N_14584,N_5171,N_8901);
xnor U14585 (N_14585,N_6658,N_5009);
xnor U14586 (N_14586,N_7265,N_9915);
nor U14587 (N_14587,N_6279,N_6359);
nor U14588 (N_14588,N_5365,N_5838);
xor U14589 (N_14589,N_7496,N_7939);
nor U14590 (N_14590,N_7393,N_7667);
nor U14591 (N_14591,N_5145,N_5505);
nor U14592 (N_14592,N_8279,N_9945);
nor U14593 (N_14593,N_8168,N_5753);
nor U14594 (N_14594,N_9140,N_7902);
or U14595 (N_14595,N_7744,N_6375);
nor U14596 (N_14596,N_9671,N_5652);
or U14597 (N_14597,N_5254,N_8123);
xnor U14598 (N_14598,N_8188,N_6174);
and U14599 (N_14599,N_8135,N_6307);
nand U14600 (N_14600,N_6776,N_7245);
or U14601 (N_14601,N_9377,N_5128);
or U14602 (N_14602,N_7456,N_9716);
nand U14603 (N_14603,N_6528,N_6070);
and U14604 (N_14604,N_9366,N_8837);
and U14605 (N_14605,N_5191,N_8479);
and U14606 (N_14606,N_7247,N_9538);
nor U14607 (N_14607,N_8526,N_5972);
nand U14608 (N_14608,N_9375,N_8033);
and U14609 (N_14609,N_8210,N_9098);
nor U14610 (N_14610,N_8909,N_5956);
and U14611 (N_14611,N_8809,N_8864);
or U14612 (N_14612,N_7929,N_7875);
or U14613 (N_14613,N_5271,N_7443);
or U14614 (N_14614,N_6964,N_9109);
nand U14615 (N_14615,N_7468,N_6564);
nor U14616 (N_14616,N_7454,N_7922);
or U14617 (N_14617,N_7254,N_8468);
or U14618 (N_14618,N_9872,N_9770);
nand U14619 (N_14619,N_5115,N_6071);
and U14620 (N_14620,N_8084,N_5931);
nand U14621 (N_14621,N_8487,N_9425);
nand U14622 (N_14622,N_9231,N_7163);
xor U14623 (N_14623,N_9549,N_8968);
xnor U14624 (N_14624,N_9629,N_8991);
nand U14625 (N_14625,N_5008,N_5678);
xor U14626 (N_14626,N_7727,N_8651);
nand U14627 (N_14627,N_9867,N_7935);
nand U14628 (N_14628,N_6465,N_9420);
nand U14629 (N_14629,N_9657,N_6695);
nor U14630 (N_14630,N_5304,N_5135);
nor U14631 (N_14631,N_6904,N_9530);
xor U14632 (N_14632,N_8377,N_7723);
nor U14633 (N_14633,N_5395,N_9693);
and U14634 (N_14634,N_6195,N_6184);
and U14635 (N_14635,N_7145,N_9536);
xor U14636 (N_14636,N_8557,N_5544);
xnor U14637 (N_14637,N_6054,N_9251);
or U14638 (N_14638,N_6412,N_5505);
xnor U14639 (N_14639,N_8808,N_5927);
or U14640 (N_14640,N_9665,N_9713);
or U14641 (N_14641,N_7217,N_6292);
or U14642 (N_14642,N_6981,N_8628);
xor U14643 (N_14643,N_9475,N_5607);
xnor U14644 (N_14644,N_9299,N_5379);
or U14645 (N_14645,N_8182,N_7318);
nor U14646 (N_14646,N_8915,N_8427);
or U14647 (N_14647,N_7971,N_9873);
or U14648 (N_14648,N_5675,N_9365);
xor U14649 (N_14649,N_6847,N_7120);
and U14650 (N_14650,N_8631,N_6645);
and U14651 (N_14651,N_5248,N_7942);
nor U14652 (N_14652,N_6777,N_6806);
nor U14653 (N_14653,N_5581,N_6188);
or U14654 (N_14654,N_6079,N_5475);
xor U14655 (N_14655,N_8415,N_6119);
or U14656 (N_14656,N_9627,N_7662);
xnor U14657 (N_14657,N_5937,N_6237);
and U14658 (N_14658,N_5437,N_6086);
nand U14659 (N_14659,N_6083,N_5749);
or U14660 (N_14660,N_6625,N_9493);
and U14661 (N_14661,N_6793,N_6668);
and U14662 (N_14662,N_8808,N_9303);
or U14663 (N_14663,N_7719,N_5960);
xnor U14664 (N_14664,N_8906,N_9318);
nand U14665 (N_14665,N_7079,N_6640);
and U14666 (N_14666,N_5105,N_6896);
nand U14667 (N_14667,N_6784,N_8260);
and U14668 (N_14668,N_7356,N_5749);
and U14669 (N_14669,N_9225,N_7922);
xnor U14670 (N_14670,N_7316,N_6080);
and U14671 (N_14671,N_9245,N_6445);
and U14672 (N_14672,N_5483,N_7560);
nand U14673 (N_14673,N_7672,N_5545);
nand U14674 (N_14674,N_5435,N_5371);
nand U14675 (N_14675,N_6146,N_9174);
nor U14676 (N_14676,N_5267,N_6378);
and U14677 (N_14677,N_5623,N_8405);
nand U14678 (N_14678,N_6808,N_8398);
or U14679 (N_14679,N_6967,N_8608);
nor U14680 (N_14680,N_7204,N_7247);
nand U14681 (N_14681,N_6246,N_5340);
xnor U14682 (N_14682,N_7645,N_6712);
or U14683 (N_14683,N_5945,N_5087);
xor U14684 (N_14684,N_8799,N_7524);
nor U14685 (N_14685,N_5717,N_7989);
nor U14686 (N_14686,N_8088,N_6384);
nand U14687 (N_14687,N_9927,N_5419);
nand U14688 (N_14688,N_7663,N_9837);
nand U14689 (N_14689,N_9803,N_8955);
and U14690 (N_14690,N_6355,N_9519);
nand U14691 (N_14691,N_6162,N_8262);
and U14692 (N_14692,N_5953,N_8106);
and U14693 (N_14693,N_9661,N_9797);
nor U14694 (N_14694,N_6812,N_6211);
nand U14695 (N_14695,N_6487,N_7955);
nand U14696 (N_14696,N_6152,N_9465);
xor U14697 (N_14697,N_5056,N_5905);
nor U14698 (N_14698,N_5686,N_7729);
xnor U14699 (N_14699,N_5631,N_9899);
and U14700 (N_14700,N_6207,N_8356);
or U14701 (N_14701,N_5406,N_9127);
xnor U14702 (N_14702,N_9287,N_6756);
or U14703 (N_14703,N_5450,N_9941);
xnor U14704 (N_14704,N_9992,N_7623);
nand U14705 (N_14705,N_6548,N_5528);
xor U14706 (N_14706,N_5030,N_5112);
and U14707 (N_14707,N_5051,N_9379);
nand U14708 (N_14708,N_8617,N_6214);
or U14709 (N_14709,N_9096,N_8042);
nand U14710 (N_14710,N_8728,N_8297);
nor U14711 (N_14711,N_9758,N_6197);
and U14712 (N_14712,N_6798,N_5255);
or U14713 (N_14713,N_7493,N_6005);
or U14714 (N_14714,N_6232,N_5461);
xor U14715 (N_14715,N_6426,N_9660);
or U14716 (N_14716,N_5896,N_7125);
or U14717 (N_14717,N_8196,N_7029);
xnor U14718 (N_14718,N_6263,N_7697);
xor U14719 (N_14719,N_8601,N_6041);
or U14720 (N_14720,N_7766,N_5819);
and U14721 (N_14721,N_7774,N_6667);
and U14722 (N_14722,N_9743,N_8655);
xnor U14723 (N_14723,N_5168,N_7691);
or U14724 (N_14724,N_9655,N_9054);
nor U14725 (N_14725,N_6759,N_8275);
xor U14726 (N_14726,N_6036,N_7519);
or U14727 (N_14727,N_9431,N_7754);
xor U14728 (N_14728,N_5013,N_7717);
and U14729 (N_14729,N_8836,N_5714);
nor U14730 (N_14730,N_5227,N_6924);
nand U14731 (N_14731,N_7734,N_9525);
nand U14732 (N_14732,N_5977,N_9852);
and U14733 (N_14733,N_8453,N_5869);
and U14734 (N_14734,N_6407,N_8487);
and U14735 (N_14735,N_8262,N_5100);
and U14736 (N_14736,N_8574,N_7498);
or U14737 (N_14737,N_5380,N_5893);
xnor U14738 (N_14738,N_5671,N_9421);
xnor U14739 (N_14739,N_6117,N_7235);
nand U14740 (N_14740,N_8120,N_9900);
nand U14741 (N_14741,N_7559,N_8332);
nor U14742 (N_14742,N_7991,N_6670);
nand U14743 (N_14743,N_6903,N_7436);
nand U14744 (N_14744,N_8875,N_5853);
xnor U14745 (N_14745,N_6883,N_6851);
nand U14746 (N_14746,N_5621,N_7211);
xnor U14747 (N_14747,N_9311,N_7769);
nor U14748 (N_14748,N_5047,N_5799);
xor U14749 (N_14749,N_6835,N_8417);
nand U14750 (N_14750,N_9969,N_8478);
xnor U14751 (N_14751,N_9700,N_9998);
or U14752 (N_14752,N_6559,N_8366);
xnor U14753 (N_14753,N_5769,N_6610);
xnor U14754 (N_14754,N_7214,N_7266);
and U14755 (N_14755,N_5112,N_6484);
nor U14756 (N_14756,N_6201,N_5617);
nor U14757 (N_14757,N_5608,N_9647);
nand U14758 (N_14758,N_7721,N_6557);
nand U14759 (N_14759,N_5941,N_7107);
or U14760 (N_14760,N_6734,N_5343);
nor U14761 (N_14761,N_7022,N_7395);
nand U14762 (N_14762,N_9110,N_5574);
nand U14763 (N_14763,N_5404,N_6831);
xnor U14764 (N_14764,N_5052,N_7145);
nor U14765 (N_14765,N_7395,N_8325);
nor U14766 (N_14766,N_6153,N_8198);
xor U14767 (N_14767,N_8903,N_6780);
and U14768 (N_14768,N_5675,N_5285);
nand U14769 (N_14769,N_7565,N_8038);
nor U14770 (N_14770,N_8985,N_9596);
nand U14771 (N_14771,N_6567,N_9420);
or U14772 (N_14772,N_9754,N_6129);
nor U14773 (N_14773,N_7009,N_6173);
nor U14774 (N_14774,N_7717,N_6538);
nor U14775 (N_14775,N_8944,N_8562);
or U14776 (N_14776,N_5646,N_6016);
and U14777 (N_14777,N_8705,N_9014);
xor U14778 (N_14778,N_8182,N_6404);
xnor U14779 (N_14779,N_7318,N_6769);
xnor U14780 (N_14780,N_7865,N_8935);
nor U14781 (N_14781,N_5918,N_8846);
and U14782 (N_14782,N_8788,N_7227);
nand U14783 (N_14783,N_5675,N_6891);
xnor U14784 (N_14784,N_5167,N_8100);
or U14785 (N_14785,N_8374,N_5917);
nand U14786 (N_14786,N_8890,N_6018);
nand U14787 (N_14787,N_7976,N_5951);
or U14788 (N_14788,N_9167,N_8257);
xor U14789 (N_14789,N_7778,N_6774);
or U14790 (N_14790,N_8781,N_8900);
nand U14791 (N_14791,N_8513,N_7708);
nand U14792 (N_14792,N_8209,N_5068);
xnor U14793 (N_14793,N_5373,N_6339);
nor U14794 (N_14794,N_8646,N_9595);
or U14795 (N_14795,N_6290,N_8327);
nand U14796 (N_14796,N_6282,N_7388);
nand U14797 (N_14797,N_7658,N_8125);
and U14798 (N_14798,N_7549,N_8427);
xnor U14799 (N_14799,N_9270,N_5976);
nand U14800 (N_14800,N_8415,N_9681);
nand U14801 (N_14801,N_7592,N_5124);
nor U14802 (N_14802,N_9902,N_6772);
and U14803 (N_14803,N_9332,N_9899);
and U14804 (N_14804,N_9349,N_6201);
and U14805 (N_14805,N_7367,N_5757);
or U14806 (N_14806,N_5745,N_6917);
xnor U14807 (N_14807,N_8585,N_6250);
nand U14808 (N_14808,N_9831,N_6634);
or U14809 (N_14809,N_8860,N_7573);
nor U14810 (N_14810,N_8362,N_7724);
nor U14811 (N_14811,N_8550,N_9120);
nor U14812 (N_14812,N_9333,N_5854);
or U14813 (N_14813,N_8934,N_8678);
xor U14814 (N_14814,N_6057,N_8770);
nor U14815 (N_14815,N_5766,N_5045);
and U14816 (N_14816,N_8379,N_6059);
xnor U14817 (N_14817,N_5217,N_7935);
and U14818 (N_14818,N_6944,N_7616);
or U14819 (N_14819,N_5577,N_9892);
and U14820 (N_14820,N_7958,N_6021);
or U14821 (N_14821,N_7132,N_6312);
and U14822 (N_14822,N_7089,N_7552);
nand U14823 (N_14823,N_6796,N_8540);
or U14824 (N_14824,N_6473,N_5284);
or U14825 (N_14825,N_9231,N_6256);
xor U14826 (N_14826,N_9688,N_7487);
xor U14827 (N_14827,N_8175,N_8896);
nand U14828 (N_14828,N_5368,N_8525);
and U14829 (N_14829,N_6011,N_6478);
and U14830 (N_14830,N_6442,N_8463);
or U14831 (N_14831,N_9988,N_9894);
nor U14832 (N_14832,N_5243,N_8243);
or U14833 (N_14833,N_8352,N_7513);
nand U14834 (N_14834,N_7241,N_7830);
nand U14835 (N_14835,N_9399,N_9140);
nand U14836 (N_14836,N_6774,N_9235);
and U14837 (N_14837,N_9413,N_9042);
nand U14838 (N_14838,N_6353,N_6760);
xnor U14839 (N_14839,N_7491,N_6831);
nor U14840 (N_14840,N_5763,N_7302);
nor U14841 (N_14841,N_8226,N_7782);
and U14842 (N_14842,N_9475,N_8798);
xor U14843 (N_14843,N_5780,N_8702);
and U14844 (N_14844,N_5720,N_9204);
nor U14845 (N_14845,N_7891,N_7808);
and U14846 (N_14846,N_6291,N_6591);
nor U14847 (N_14847,N_5647,N_5796);
xnor U14848 (N_14848,N_6125,N_9487);
nor U14849 (N_14849,N_9274,N_7309);
and U14850 (N_14850,N_5288,N_9094);
xor U14851 (N_14851,N_5680,N_7407);
and U14852 (N_14852,N_7796,N_6806);
and U14853 (N_14853,N_6948,N_9410);
nand U14854 (N_14854,N_8362,N_7712);
nand U14855 (N_14855,N_9823,N_7231);
or U14856 (N_14856,N_9679,N_8371);
or U14857 (N_14857,N_7199,N_5816);
and U14858 (N_14858,N_5370,N_6340);
nor U14859 (N_14859,N_5596,N_5204);
xnor U14860 (N_14860,N_8105,N_6590);
nor U14861 (N_14861,N_6955,N_5545);
and U14862 (N_14862,N_7740,N_8745);
nor U14863 (N_14863,N_9236,N_9725);
or U14864 (N_14864,N_8172,N_6969);
or U14865 (N_14865,N_5531,N_9388);
and U14866 (N_14866,N_7053,N_5571);
nand U14867 (N_14867,N_9178,N_5936);
nand U14868 (N_14868,N_9794,N_7869);
or U14869 (N_14869,N_9775,N_5090);
and U14870 (N_14870,N_8922,N_7501);
xnor U14871 (N_14871,N_8024,N_5979);
nor U14872 (N_14872,N_8187,N_9174);
nand U14873 (N_14873,N_8594,N_7633);
nor U14874 (N_14874,N_8714,N_6228);
and U14875 (N_14875,N_5405,N_8646);
nand U14876 (N_14876,N_6119,N_5738);
or U14877 (N_14877,N_9938,N_9773);
nor U14878 (N_14878,N_7293,N_6044);
and U14879 (N_14879,N_7249,N_9501);
nor U14880 (N_14880,N_5634,N_7668);
nand U14881 (N_14881,N_6274,N_6158);
and U14882 (N_14882,N_9681,N_7440);
or U14883 (N_14883,N_8361,N_8537);
and U14884 (N_14884,N_5699,N_8316);
and U14885 (N_14885,N_9858,N_6927);
and U14886 (N_14886,N_7286,N_5183);
nor U14887 (N_14887,N_7312,N_7331);
and U14888 (N_14888,N_5577,N_6803);
and U14889 (N_14889,N_9116,N_5719);
or U14890 (N_14890,N_8729,N_8428);
or U14891 (N_14891,N_5843,N_8149);
nor U14892 (N_14892,N_8806,N_6792);
xnor U14893 (N_14893,N_7866,N_8282);
and U14894 (N_14894,N_6497,N_9939);
nor U14895 (N_14895,N_5379,N_8123);
or U14896 (N_14896,N_6888,N_7950);
xor U14897 (N_14897,N_9629,N_9644);
or U14898 (N_14898,N_6915,N_7965);
nor U14899 (N_14899,N_7375,N_8100);
xnor U14900 (N_14900,N_6989,N_8370);
nor U14901 (N_14901,N_9801,N_9092);
nand U14902 (N_14902,N_9414,N_7073);
nand U14903 (N_14903,N_6776,N_7184);
nor U14904 (N_14904,N_7576,N_9351);
or U14905 (N_14905,N_5272,N_6080);
xor U14906 (N_14906,N_7560,N_9198);
nand U14907 (N_14907,N_6957,N_9790);
xor U14908 (N_14908,N_8747,N_6508);
nor U14909 (N_14909,N_9280,N_6701);
or U14910 (N_14910,N_5925,N_6606);
nand U14911 (N_14911,N_5005,N_5864);
and U14912 (N_14912,N_5283,N_9635);
and U14913 (N_14913,N_6936,N_5109);
nor U14914 (N_14914,N_5048,N_9123);
or U14915 (N_14915,N_7336,N_7365);
xnor U14916 (N_14916,N_9704,N_6178);
and U14917 (N_14917,N_9525,N_9832);
nand U14918 (N_14918,N_7263,N_9553);
nand U14919 (N_14919,N_5439,N_7563);
and U14920 (N_14920,N_9020,N_7020);
nor U14921 (N_14921,N_8195,N_5239);
nor U14922 (N_14922,N_9479,N_7078);
and U14923 (N_14923,N_9267,N_6490);
nand U14924 (N_14924,N_5409,N_5110);
or U14925 (N_14925,N_6774,N_8216);
and U14926 (N_14926,N_7273,N_7173);
and U14927 (N_14927,N_9577,N_6354);
or U14928 (N_14928,N_5693,N_6493);
nand U14929 (N_14929,N_7824,N_9519);
nor U14930 (N_14930,N_6009,N_6270);
and U14931 (N_14931,N_6015,N_9647);
or U14932 (N_14932,N_8909,N_6256);
nand U14933 (N_14933,N_8121,N_6888);
or U14934 (N_14934,N_6952,N_7313);
nand U14935 (N_14935,N_6199,N_5898);
xor U14936 (N_14936,N_8553,N_5883);
xnor U14937 (N_14937,N_8916,N_6905);
xnor U14938 (N_14938,N_6203,N_5788);
and U14939 (N_14939,N_6046,N_7832);
or U14940 (N_14940,N_8851,N_6539);
or U14941 (N_14941,N_6915,N_7427);
and U14942 (N_14942,N_7984,N_9525);
nand U14943 (N_14943,N_8984,N_9418);
and U14944 (N_14944,N_6889,N_7983);
nor U14945 (N_14945,N_8975,N_5321);
xnor U14946 (N_14946,N_6292,N_8579);
nor U14947 (N_14947,N_7079,N_9736);
or U14948 (N_14948,N_8996,N_7884);
xnor U14949 (N_14949,N_6723,N_5335);
and U14950 (N_14950,N_6584,N_7643);
or U14951 (N_14951,N_7236,N_8503);
nand U14952 (N_14952,N_8426,N_5380);
nor U14953 (N_14953,N_7872,N_6675);
xor U14954 (N_14954,N_8296,N_9247);
nand U14955 (N_14955,N_6471,N_7583);
xor U14956 (N_14956,N_7583,N_9992);
and U14957 (N_14957,N_8041,N_8833);
xnor U14958 (N_14958,N_7225,N_8547);
and U14959 (N_14959,N_6484,N_7252);
and U14960 (N_14960,N_7471,N_6137);
xor U14961 (N_14961,N_6069,N_8573);
nand U14962 (N_14962,N_9581,N_7571);
nor U14963 (N_14963,N_8628,N_6834);
xnor U14964 (N_14964,N_6367,N_5486);
nand U14965 (N_14965,N_7074,N_7307);
nand U14966 (N_14966,N_8679,N_6570);
and U14967 (N_14967,N_8144,N_9623);
and U14968 (N_14968,N_5639,N_5088);
or U14969 (N_14969,N_8998,N_7312);
and U14970 (N_14970,N_9625,N_8030);
xor U14971 (N_14971,N_9831,N_7498);
nor U14972 (N_14972,N_9731,N_6644);
xor U14973 (N_14973,N_9758,N_5184);
and U14974 (N_14974,N_6144,N_8653);
xor U14975 (N_14975,N_8103,N_6849);
and U14976 (N_14976,N_9829,N_9867);
nor U14977 (N_14977,N_9672,N_5010);
nand U14978 (N_14978,N_6188,N_9829);
and U14979 (N_14979,N_5071,N_6159);
and U14980 (N_14980,N_6250,N_9142);
xnor U14981 (N_14981,N_8092,N_5083);
nand U14982 (N_14982,N_9285,N_5049);
or U14983 (N_14983,N_7781,N_8059);
xor U14984 (N_14984,N_7315,N_6265);
nand U14985 (N_14985,N_8787,N_9981);
xnor U14986 (N_14986,N_9103,N_5221);
nand U14987 (N_14987,N_9057,N_6209);
nand U14988 (N_14988,N_9530,N_9938);
xor U14989 (N_14989,N_5794,N_5944);
nand U14990 (N_14990,N_6796,N_5372);
and U14991 (N_14991,N_6170,N_9390);
nand U14992 (N_14992,N_5984,N_9944);
and U14993 (N_14993,N_7170,N_9998);
and U14994 (N_14994,N_5281,N_8851);
and U14995 (N_14995,N_6579,N_6876);
nor U14996 (N_14996,N_9112,N_6337);
nand U14997 (N_14997,N_6449,N_8920);
or U14998 (N_14998,N_8651,N_5250);
xor U14999 (N_14999,N_7765,N_8400);
or U15000 (N_15000,N_13847,N_10551);
or U15001 (N_15001,N_13177,N_11097);
xnor U15002 (N_15002,N_14034,N_12937);
xnor U15003 (N_15003,N_11840,N_14432);
nor U15004 (N_15004,N_10250,N_13829);
or U15005 (N_15005,N_10308,N_11508);
or U15006 (N_15006,N_12384,N_14231);
nor U15007 (N_15007,N_13542,N_14512);
or U15008 (N_15008,N_13752,N_12736);
xor U15009 (N_15009,N_13511,N_13367);
nand U15010 (N_15010,N_14038,N_10450);
xnor U15011 (N_15011,N_13644,N_12274);
nand U15012 (N_15012,N_10651,N_14307);
nor U15013 (N_15013,N_14398,N_14255);
and U15014 (N_15014,N_10330,N_14373);
or U15015 (N_15015,N_14205,N_14568);
xnor U15016 (N_15016,N_11115,N_14549);
or U15017 (N_15017,N_14771,N_13759);
xnor U15018 (N_15018,N_13486,N_11376);
nand U15019 (N_15019,N_14413,N_10861);
or U15020 (N_15020,N_12462,N_13495);
nor U15021 (N_15021,N_11882,N_13278);
xor U15022 (N_15022,N_14901,N_11237);
and U15023 (N_15023,N_10119,N_14260);
nor U15024 (N_15024,N_11394,N_14388);
or U15025 (N_15025,N_10801,N_11706);
nor U15026 (N_15026,N_14378,N_10632);
nand U15027 (N_15027,N_14759,N_10735);
and U15028 (N_15028,N_11675,N_12538);
or U15029 (N_15029,N_14560,N_13352);
xor U15030 (N_15030,N_12821,N_10769);
or U15031 (N_15031,N_10665,N_11952);
or U15032 (N_15032,N_13794,N_12555);
xnor U15033 (N_15033,N_14139,N_11057);
and U15034 (N_15034,N_10822,N_11514);
and U15035 (N_15035,N_10678,N_10664);
nor U15036 (N_15036,N_11728,N_12119);
and U15037 (N_15037,N_11737,N_13476);
nand U15038 (N_15038,N_10655,N_14000);
nor U15039 (N_15039,N_10724,N_11272);
or U15040 (N_15040,N_14003,N_11784);
nand U15041 (N_15041,N_12654,N_11761);
and U15042 (N_15042,N_14698,N_12929);
xnor U15043 (N_15043,N_10509,N_13425);
nor U15044 (N_15044,N_11933,N_11162);
nand U15045 (N_15045,N_11816,N_10054);
or U15046 (N_15046,N_13297,N_11183);
nand U15047 (N_15047,N_13749,N_13030);
and U15048 (N_15048,N_10370,N_10685);
and U15049 (N_15049,N_12469,N_10560);
and U15050 (N_15050,N_12315,N_12557);
nor U15051 (N_15051,N_11461,N_11854);
and U15052 (N_15052,N_11165,N_11665);
nor U15053 (N_15053,N_14739,N_10668);
or U15054 (N_15054,N_10725,N_11850);
and U15055 (N_15055,N_10599,N_13783);
nand U15056 (N_15056,N_11651,N_11253);
xnor U15057 (N_15057,N_13593,N_13727);
or U15058 (N_15058,N_13139,N_12710);
xnor U15059 (N_15059,N_12218,N_10025);
xnor U15060 (N_15060,N_12897,N_13731);
or U15061 (N_15061,N_12322,N_10072);
nor U15062 (N_15062,N_13600,N_12797);
nor U15063 (N_15063,N_11060,N_13518);
and U15064 (N_15064,N_10293,N_11821);
nor U15065 (N_15065,N_11179,N_12790);
xor U15066 (N_15066,N_12443,N_10000);
and U15067 (N_15067,N_13011,N_10647);
and U15068 (N_15068,N_12446,N_11871);
nand U15069 (N_15069,N_12418,N_10006);
and U15070 (N_15070,N_10985,N_14132);
nor U15071 (N_15071,N_10317,N_12985);
xor U15072 (N_15072,N_10302,N_11746);
nor U15073 (N_15073,N_10439,N_13268);
or U15074 (N_15074,N_10579,N_14480);
nand U15075 (N_15075,N_14304,N_12295);
nand U15076 (N_15076,N_12019,N_11388);
nor U15077 (N_15077,N_12109,N_14521);
nor U15078 (N_15078,N_10559,N_12297);
xor U15079 (N_15079,N_10583,N_13730);
nor U15080 (N_15080,N_10398,N_10197);
nor U15081 (N_15081,N_11369,N_10917);
nor U15082 (N_15082,N_14658,N_13928);
nor U15083 (N_15083,N_10311,N_14915);
and U15084 (N_15084,N_12740,N_10991);
nor U15085 (N_15085,N_13843,N_14696);
or U15086 (N_15086,N_10109,N_14562);
nand U15087 (N_15087,N_13360,N_11013);
nand U15088 (N_15088,N_12166,N_12636);
xor U15089 (N_15089,N_10972,N_14939);
and U15090 (N_15090,N_11507,N_13611);
nand U15091 (N_15091,N_10561,N_12073);
and U15092 (N_15092,N_10737,N_13299);
nor U15093 (N_15093,N_11039,N_10835);
xnor U15094 (N_15094,N_12831,N_11009);
nand U15095 (N_15095,N_11061,N_11075);
xor U15096 (N_15096,N_10783,N_10211);
nor U15097 (N_15097,N_13499,N_11518);
and U15098 (N_15098,N_10037,N_12035);
nand U15099 (N_15099,N_12076,N_14914);
xor U15100 (N_15100,N_12270,N_14389);
nor U15101 (N_15101,N_14297,N_14588);
and U15102 (N_15102,N_14346,N_14923);
or U15103 (N_15103,N_10891,N_10521);
nor U15104 (N_15104,N_11926,N_13899);
and U15105 (N_15105,N_14174,N_10947);
or U15106 (N_15106,N_11741,N_10981);
nor U15107 (N_15107,N_13066,N_14835);
and U15108 (N_15108,N_12352,N_10837);
and U15109 (N_15109,N_12974,N_14276);
nand U15110 (N_15110,N_13019,N_11722);
or U15111 (N_15111,N_10849,N_14285);
or U15112 (N_15112,N_11723,N_10076);
and U15113 (N_15113,N_13962,N_14965);
and U15114 (N_15114,N_10720,N_13646);
xnor U15115 (N_15115,N_11607,N_13159);
xor U15116 (N_15116,N_12908,N_13024);
xor U15117 (N_15117,N_12771,N_14671);
and U15118 (N_15118,N_13801,N_11585);
nor U15119 (N_15119,N_12904,N_14456);
nand U15120 (N_15120,N_12133,N_13116);
nand U15121 (N_15121,N_14317,N_11537);
xnor U15122 (N_15122,N_12602,N_12940);
or U15123 (N_15123,N_13036,N_12379);
nand U15124 (N_15124,N_11591,N_10553);
and U15125 (N_15125,N_14256,N_13756);
nor U15126 (N_15126,N_14274,N_12359);
nand U15127 (N_15127,N_12021,N_12521);
and U15128 (N_15128,N_12578,N_14889);
nor U15129 (N_15129,N_13525,N_10797);
nor U15130 (N_15130,N_14640,N_14214);
nand U15131 (N_15131,N_10018,N_10320);
or U15132 (N_15132,N_12962,N_12535);
or U15133 (N_15133,N_12098,N_13723);
nor U15134 (N_15134,N_14689,N_12241);
nand U15135 (N_15135,N_13325,N_12249);
xnor U15136 (N_15136,N_10518,N_13535);
or U15137 (N_15137,N_14870,N_12999);
nand U15138 (N_15138,N_12504,N_11666);
and U15139 (N_15139,N_11993,N_11225);
or U15140 (N_15140,N_11469,N_13197);
nand U15141 (N_15141,N_10762,N_12139);
nand U15142 (N_15142,N_14200,N_10192);
nor U15143 (N_15143,N_13844,N_12769);
xor U15144 (N_15144,N_11181,N_14970);
xnor U15145 (N_15145,N_10160,N_11407);
or U15146 (N_15146,N_12991,N_13787);
xor U15147 (N_15147,N_13185,N_12095);
or U15148 (N_15148,N_14576,N_12012);
or U15149 (N_15149,N_14111,N_11863);
or U15150 (N_15150,N_11405,N_13414);
or U15151 (N_15151,N_10003,N_14728);
nand U15152 (N_15152,N_12569,N_12230);
xor U15153 (N_15153,N_13991,N_13242);
nor U15154 (N_15154,N_11466,N_13208);
or U15155 (N_15155,N_14077,N_13869);
and U15156 (N_15156,N_13624,N_14185);
and U15157 (N_15157,N_11564,N_11359);
or U15158 (N_15158,N_10992,N_10306);
nand U15159 (N_15159,N_14156,N_12993);
or U15160 (N_15160,N_13097,N_10613);
xor U15161 (N_15161,N_11476,N_10814);
and U15162 (N_15162,N_11966,N_14451);
and U15163 (N_15163,N_12575,N_14999);
xor U15164 (N_15164,N_10777,N_10935);
nand U15165 (N_15165,N_11468,N_12090);
or U15166 (N_15166,N_11202,N_10152);
and U15167 (N_15167,N_13851,N_12630);
or U15168 (N_15168,N_14046,N_13101);
or U15169 (N_15169,N_11453,N_11358);
or U15170 (N_15170,N_11963,N_14873);
and U15171 (N_15171,N_10221,N_11629);
and U15172 (N_15172,N_14426,N_10683);
nor U15173 (N_15173,N_14005,N_13539);
nand U15174 (N_15174,N_10957,N_14263);
and U15175 (N_15175,N_12552,N_10879);
nor U15176 (N_15176,N_13190,N_12977);
or U15177 (N_15177,N_10968,N_12323);
or U15178 (N_15178,N_12163,N_10165);
nand U15179 (N_15179,N_10434,N_13063);
xor U15180 (N_15180,N_13547,N_14164);
or U15181 (N_15181,N_11941,N_10130);
or U15182 (N_15182,N_14750,N_10421);
or U15183 (N_15183,N_14172,N_11605);
nand U15184 (N_15184,N_10209,N_14711);
nor U15185 (N_15185,N_11983,N_12261);
and U15186 (N_15186,N_13983,N_13893);
or U15187 (N_15187,N_10066,N_14395);
nor U15188 (N_15188,N_14673,N_14392);
xnor U15189 (N_15189,N_11556,N_11553);
nand U15190 (N_15190,N_10527,N_11008);
nand U15191 (N_15191,N_10078,N_14128);
nor U15192 (N_15192,N_10349,N_14613);
or U15193 (N_15193,N_10299,N_11891);
nor U15194 (N_15194,N_12312,N_13709);
or U15195 (N_15195,N_12416,N_11695);
nand U15196 (N_15196,N_11119,N_10490);
nor U15197 (N_15197,N_10718,N_12406);
nor U15198 (N_15198,N_11943,N_10823);
nand U15199 (N_15199,N_11472,N_14683);
nand U15200 (N_15200,N_10813,N_12096);
nand U15201 (N_15201,N_11163,N_14848);
nor U15202 (N_15202,N_10229,N_14208);
or U15203 (N_15203,N_14025,N_11562);
nand U15204 (N_15204,N_14887,N_12455);
nor U15205 (N_15205,N_14226,N_12470);
and U15206 (N_15206,N_14367,N_10011);
and U15207 (N_15207,N_13627,N_13722);
or U15208 (N_15208,N_14353,N_14736);
or U15209 (N_15209,N_14031,N_12373);
or U15210 (N_15210,N_14802,N_14151);
xnor U15211 (N_15211,N_10112,N_14840);
xnor U15212 (N_15212,N_12219,N_13519);
nor U15213 (N_15213,N_10864,N_13815);
nor U15214 (N_15214,N_10913,N_10510);
nand U15215 (N_15215,N_10501,N_12318);
and U15216 (N_15216,N_10923,N_12757);
xor U15217 (N_15217,N_12795,N_10567);
nand U15218 (N_15218,N_10044,N_12804);
xnor U15219 (N_15219,N_14384,N_11501);
or U15220 (N_15220,N_10485,N_10322);
nand U15221 (N_15221,N_12078,N_10889);
nand U15222 (N_15222,N_10540,N_14559);
nand U15223 (N_15223,N_14827,N_11631);
xnor U15224 (N_15224,N_13091,N_13803);
and U15225 (N_15225,N_13006,N_11839);
nor U15226 (N_15226,N_11245,N_10051);
and U15227 (N_15227,N_12498,N_10164);
or U15228 (N_15228,N_13427,N_10159);
nor U15229 (N_15229,N_14183,N_13599);
xor U15230 (N_15230,N_12070,N_13174);
nand U15231 (N_15231,N_10691,N_12687);
and U15232 (N_15232,N_11226,N_11826);
and U15233 (N_15233,N_13253,N_10815);
nor U15234 (N_15234,N_12217,N_13065);
and U15235 (N_15235,N_14067,N_13919);
and U15236 (N_15236,N_14474,N_13305);
or U15237 (N_15237,N_10385,N_10832);
and U15238 (N_15238,N_12492,N_10145);
and U15239 (N_15239,N_14533,N_13175);
xor U15240 (N_15240,N_11798,N_13937);
and U15241 (N_15241,N_11547,N_14851);
and U15242 (N_15242,N_13092,N_10852);
or U15243 (N_15243,N_12099,N_10682);
and U15244 (N_15244,N_13656,N_14819);
and U15245 (N_15245,N_11534,N_11528);
nor U15246 (N_15246,N_12001,N_13114);
and U15247 (N_15247,N_13343,N_14041);
nor U15248 (N_15248,N_14730,N_10939);
nand U15249 (N_15249,N_13864,N_12881);
or U15250 (N_15250,N_13469,N_14141);
xnor U15251 (N_15251,N_12648,N_14268);
nand U15252 (N_15252,N_13573,N_13357);
nor U15253 (N_15253,N_11146,N_11221);
and U15254 (N_15254,N_10220,N_14403);
and U15255 (N_15255,N_13306,N_12817);
nor U15256 (N_15256,N_11938,N_14047);
nor U15257 (N_15257,N_11417,N_13247);
nand U15258 (N_15258,N_13659,N_11979);
nor U15259 (N_15259,N_12606,N_11834);
xor U15260 (N_15260,N_13123,N_12588);
or U15261 (N_15261,N_14845,N_12420);
xor U15262 (N_15262,N_13396,N_12190);
nor U15263 (N_15263,N_11747,N_10589);
xnor U15264 (N_15264,N_11457,N_12043);
xnor U15265 (N_15265,N_11026,N_12691);
nand U15266 (N_15266,N_11006,N_12425);
xnor U15267 (N_15267,N_14023,N_13854);
nor U15268 (N_15268,N_10824,N_13583);
nand U15269 (N_15269,N_10378,N_14675);
nand U15270 (N_15270,N_10663,N_14612);
xnor U15271 (N_15271,N_11445,N_10848);
or U15272 (N_15272,N_10169,N_11076);
xnor U15273 (N_15273,N_14587,N_11596);
or U15274 (N_15274,N_13826,N_11392);
or U15275 (N_15275,N_12942,N_11649);
nand U15276 (N_15276,N_13321,N_14997);
and U15277 (N_15277,N_10318,N_13812);
or U15278 (N_15278,N_14291,N_10042);
xnor U15279 (N_15279,N_14905,N_14390);
nor U15280 (N_15280,N_10883,N_11645);
nor U15281 (N_15281,N_14407,N_12149);
and U15282 (N_15282,N_13680,N_13497);
and U15283 (N_15283,N_13737,N_14891);
xor U15284 (N_15284,N_10836,N_12450);
and U15285 (N_15285,N_14779,N_14108);
or U15286 (N_15286,N_10468,N_10043);
or U15287 (N_15287,N_13913,N_10695);
nor U15288 (N_15288,N_12135,N_13809);
xor U15289 (N_15289,N_13914,N_12819);
xor U15290 (N_15290,N_13412,N_12642);
nor U15291 (N_15291,N_11016,N_13956);
and U15292 (N_15292,N_14314,N_11180);
and U15293 (N_15293,N_14780,N_13523);
nor U15294 (N_15294,N_11391,N_10107);
nor U15295 (N_15295,N_14859,N_14712);
and U15296 (N_15296,N_13086,N_12176);
or U15297 (N_15297,N_10892,N_14188);
nor U15298 (N_15298,N_14941,N_10873);
and U15299 (N_15299,N_10020,N_13977);
nor U15300 (N_15300,N_13835,N_12826);
and U15301 (N_15301,N_13373,N_12242);
and U15302 (N_15302,N_14095,N_11311);
nor U15303 (N_15303,N_10175,N_10854);
nor U15304 (N_15304,N_10733,N_10807);
nor U15305 (N_15305,N_10536,N_12240);
nor U15306 (N_15306,N_12433,N_14189);
or U15307 (N_15307,N_13700,N_12961);
nand U15308 (N_15308,N_13952,N_11250);
and U15309 (N_15309,N_14785,N_13435);
xnor U15310 (N_15310,N_12540,N_14322);
nor U15311 (N_15311,N_10362,N_12692);
nand U15312 (N_15312,N_12998,N_13182);
nand U15313 (N_15313,N_11024,N_12832);
nor U15314 (N_15314,N_10471,N_14947);
nor U15315 (N_15315,N_13963,N_10336);
nor U15316 (N_15316,N_14879,N_11962);
xor U15317 (N_15317,N_14610,N_14366);
nor U15318 (N_15318,N_12252,N_10853);
or U15319 (N_15319,N_13852,N_10996);
xnor U15320 (N_15320,N_13764,N_12104);
and U15321 (N_15321,N_13686,N_13503);
or U15322 (N_15322,N_14142,N_10467);
nor U15323 (N_15323,N_13781,N_10893);
or U15324 (N_15324,N_14862,N_14433);
nand U15325 (N_15325,N_14977,N_14863);
nand U15326 (N_15326,N_14381,N_11458);
xnor U15327 (N_15327,N_12667,N_14415);
xnor U15328 (N_15328,N_12143,N_11708);
xor U15329 (N_15329,N_11851,N_11827);
nand U15330 (N_15330,N_12150,N_13702);
xor U15331 (N_15331,N_14394,N_13432);
or U15332 (N_15332,N_14742,N_14198);
nor U15333 (N_15333,N_13566,N_12660);
nand U15334 (N_15334,N_10126,N_13084);
nor U15335 (N_15335,N_11557,N_11340);
xnor U15336 (N_15336,N_14738,N_12476);
xor U15337 (N_15337,N_14931,N_11716);
or U15338 (N_15338,N_13556,N_14455);
xnor U15339 (N_15339,N_10260,N_11561);
nand U15340 (N_15340,N_11520,N_11378);
or U15341 (N_15341,N_11140,N_10137);
and U15342 (N_15342,N_12449,N_10565);
and U15343 (N_15343,N_14306,N_10995);
nand U15344 (N_15344,N_13677,N_12199);
nand U15345 (N_15345,N_11465,N_13415);
nor U15346 (N_15346,N_10062,N_10028);
xor U15347 (N_15347,N_14216,N_14973);
xnor U15348 (N_15348,N_12356,N_13560);
or U15349 (N_15349,N_14438,N_12522);
nor U15350 (N_15350,N_12807,N_14133);
or U15351 (N_15351,N_14801,N_12197);
or U15352 (N_15352,N_11931,N_11361);
nand U15353 (N_15353,N_14747,N_13155);
xnor U15354 (N_15354,N_12286,N_11693);
nor U15355 (N_15355,N_14158,N_10396);
nand U15356 (N_15356,N_12011,N_14866);
xor U15357 (N_15357,N_10546,N_13342);
xor U15358 (N_15358,N_14335,N_11733);
nand U15359 (N_15359,N_12571,N_12992);
xor U15360 (N_15360,N_10369,N_14545);
xor U15361 (N_15361,N_14962,N_12623);
nor U15362 (N_15362,N_11604,N_14769);
and U15363 (N_15363,N_14875,N_11364);
nor U15364 (N_15364,N_10834,N_12553);
xnor U15365 (N_15365,N_10156,N_12127);
or U15366 (N_15366,N_10556,N_10931);
and U15367 (N_15367,N_14792,N_12823);
xnor U15368 (N_15368,N_13958,N_12800);
and U15369 (N_15369,N_12672,N_11449);
nand U15370 (N_15370,N_14953,N_12935);
or U15371 (N_15371,N_10674,N_13302);
xnor U15372 (N_15372,N_10158,N_11948);
nor U15373 (N_15373,N_14918,N_12594);
nor U15374 (N_15374,N_10381,N_14656);
xor U15375 (N_15375,N_13034,N_13642);
nand U15376 (N_15376,N_10870,N_10268);
xnor U15377 (N_15377,N_14277,N_12305);
or U15378 (N_15378,N_11262,N_11434);
and U15379 (N_15379,N_10089,N_12256);
or U15380 (N_15380,N_10980,N_12296);
or U15381 (N_15381,N_10606,N_14577);
nor U15382 (N_15382,N_11421,N_12385);
nor U15383 (N_15383,N_13178,N_14502);
xor U15384 (N_15384,N_10614,N_13742);
nand U15385 (N_15385,N_12953,N_14607);
xnor U15386 (N_15386,N_14760,N_11273);
nand U15387 (N_15387,N_11815,N_13046);
and U15388 (N_15388,N_10855,N_13459);
or U15389 (N_15389,N_14352,N_12188);
xnor U15390 (N_15390,N_12888,N_10590);
and U15391 (N_15391,N_12709,N_10754);
and U15392 (N_15392,N_10358,N_11859);
xnor U15393 (N_15393,N_14626,N_11397);
xnor U15394 (N_15394,N_14572,N_10217);
nand U15395 (N_15395,N_12234,N_10438);
or U15396 (N_15396,N_10756,N_14147);
or U15397 (N_15397,N_12387,N_13072);
and U15398 (N_15398,N_12747,N_12154);
xor U15399 (N_15399,N_11430,N_13716);
nand U15400 (N_15400,N_12331,N_12868);
or U15401 (N_15401,N_10462,N_12120);
or U15402 (N_15402,N_10454,N_12034);
nor U15403 (N_15403,N_10281,N_11806);
and U15404 (N_15404,N_10266,N_11320);
or U15405 (N_15405,N_13870,N_13681);
nor U15406 (N_15406,N_11310,N_14539);
or U15407 (N_15407,N_13473,N_13558);
nor U15408 (N_15408,N_12457,N_11612);
nor U15409 (N_15409,N_11847,N_11803);
or U15410 (N_15410,N_11251,N_13865);
nor U15411 (N_15411,N_13521,N_11531);
and U15412 (N_15412,N_14908,N_12894);
nor U15413 (N_15413,N_14064,N_10451);
and U15414 (N_15414,N_14452,N_14429);
nor U15415 (N_15415,N_11809,N_13438);
nor U15416 (N_15416,N_12415,N_13944);
nand U15417 (N_15417,N_13385,N_11935);
nand U15418 (N_15418,N_14496,N_14987);
nand U15419 (N_15419,N_11523,N_14471);
and U15420 (N_15420,N_14595,N_14217);
and U15421 (N_15421,N_13064,N_13203);
or U15422 (N_15422,N_11099,N_13222);
nor U15423 (N_15423,N_13947,N_14633);
nor U15424 (N_15424,N_11240,N_10914);
or U15425 (N_15425,N_14431,N_10908);
or U15426 (N_15426,N_13721,N_10932);
xnor U15427 (N_15427,N_13652,N_11744);
or U15428 (N_15428,N_13274,N_11450);
xor U15429 (N_15429,N_10831,N_10272);
and U15430 (N_15430,N_12262,N_13776);
or U15431 (N_15431,N_13340,N_10920);
xor U15432 (N_15432,N_12517,N_13200);
xnor U15433 (N_15433,N_13632,N_10446);
nand U15434 (N_15434,N_11663,N_12341);
or U15435 (N_15435,N_14240,N_14167);
or U15436 (N_15436,N_14877,N_14150);
and U15437 (N_15437,N_11515,N_11735);
nor U15438 (N_15438,N_11877,N_13773);
or U15439 (N_15439,N_10727,N_11265);
xor U15440 (N_15440,N_12701,N_10186);
nor U15441 (N_15441,N_11495,N_13201);
or U15442 (N_15442,N_14547,N_11322);
nor U15443 (N_15443,N_11589,N_10496);
xnor U15444 (N_15444,N_12276,N_10595);
nor U15445 (N_15445,N_14755,N_14227);
nand U15446 (N_15446,N_12547,N_10752);
nor U15447 (N_15447,N_12475,N_10646);
xor U15448 (N_15448,N_10515,N_14491);
xnor U15449 (N_15449,N_14063,N_10731);
nor U15450 (N_15450,N_11902,N_11467);
and U15451 (N_15451,N_10817,N_10472);
and U15452 (N_15452,N_11498,N_13233);
nor U15453 (N_15453,N_10424,N_11486);
or U15454 (N_15454,N_11263,N_11090);
nand U15455 (N_15455,N_12015,N_10170);
nor U15456 (N_15456,N_10729,N_12563);
or U15457 (N_15457,N_11415,N_11185);
xnor U15458 (N_15458,N_10403,N_14110);
xor U15459 (N_15459,N_13027,N_10508);
and U15460 (N_15460,N_13935,N_14505);
xnor U15461 (N_15461,N_10693,N_14513);
xnor U15462 (N_15462,N_10397,N_10466);
nor U15463 (N_15463,N_11156,N_14551);
nor U15464 (N_15464,N_14045,N_10662);
and U15465 (N_15465,N_14791,N_11572);
and U15466 (N_15466,N_14334,N_13649);
xor U15467 (N_15467,N_12577,N_12306);
nor U15468 (N_15468,N_13619,N_11113);
nand U15469 (N_15469,N_12485,N_11010);
xor U15470 (N_15470,N_13366,N_10484);
and U15471 (N_15471,N_10481,N_10327);
nor U15472 (N_15472,N_10440,N_13337);
nand U15473 (N_15473,N_13874,N_14404);
nor U15474 (N_15474,N_12003,N_11046);
or U15475 (N_15475,N_11177,N_14466);
nand U15476 (N_15476,N_14035,N_12766);
nand U15477 (N_15477,N_10200,N_13315);
and U15478 (N_15478,N_11872,N_12941);
nor U15479 (N_15479,N_14036,N_11890);
xor U15480 (N_15480,N_11802,N_14855);
or U15481 (N_15481,N_13882,N_12558);
or U15482 (N_15482,N_13471,N_13607);
xor U15483 (N_15483,N_13949,N_11095);
nor U15484 (N_15484,N_12027,N_12607);
nor U15485 (N_15485,N_10698,N_14437);
and U15486 (N_15486,N_14218,N_11647);
and U15487 (N_15487,N_11883,N_11576);
nand U15488 (N_15488,N_14103,N_10304);
or U15489 (N_15489,N_10649,N_13615);
and U15490 (N_15490,N_12928,N_12040);
or U15491 (N_15491,N_10643,N_10263);
nand U15492 (N_15492,N_10912,N_10065);
nor U15493 (N_15493,N_13285,N_13160);
nand U15494 (N_15494,N_12069,N_13141);
or U15495 (N_15495,N_14190,N_12292);
nand U15496 (N_15496,N_10759,N_14872);
nand U15497 (N_15497,N_13095,N_12417);
nand U15498 (N_15498,N_14184,N_14186);
nor U15499 (N_15499,N_12271,N_10463);
or U15500 (N_15500,N_12264,N_10081);
nor U15501 (N_15501,N_11930,N_11644);
nor U15502 (N_15502,N_12789,N_11223);
xor U15503 (N_15503,N_12468,N_13822);
or U15504 (N_15504,N_11153,N_10641);
nand U15505 (N_15505,N_12390,N_13805);
nor U15506 (N_15506,N_14768,N_13501);
or U15507 (N_15507,N_12678,N_13117);
xnor U15508 (N_15508,N_12793,N_14702);
and U15509 (N_15509,N_13127,N_13698);
nand U15510 (N_15510,N_11351,N_12228);
xor U15511 (N_15511,N_11951,N_13405);
nor U15512 (N_15512,N_10477,N_14477);
nor U15513 (N_15513,N_12082,N_10488);
nand U15514 (N_15514,N_13930,N_11081);
nor U15515 (N_15515,N_13591,N_10504);
nand U15516 (N_15516,N_13746,N_14800);
or U15517 (N_15517,N_12722,N_13969);
nor U15518 (N_15518,N_11538,N_14101);
and U15519 (N_15519,N_11636,N_10886);
xnor U15520 (N_15520,N_13484,N_13666);
and U15521 (N_15521,N_10257,N_11494);
or U15522 (N_15522,N_13966,N_11985);
xor U15523 (N_15523,N_14749,N_10291);
nand U15524 (N_15524,N_11116,N_10978);
xor U15525 (N_15525,N_12750,N_10804);
xnor U15526 (N_15526,N_10790,N_12730);
nor U15527 (N_15527,N_13853,N_14567);
nor U15528 (N_15528,N_11268,N_12626);
and U15529 (N_15529,N_13398,N_13610);
nand U15530 (N_15530,N_10743,N_12556);
nor U15531 (N_15531,N_13265,N_10778);
or U15532 (N_15532,N_13061,N_12964);
nor U15533 (N_15533,N_10057,N_13586);
xor U15534 (N_15534,N_14333,N_12032);
nand U15535 (N_15535,N_14236,N_11797);
or U15536 (N_15536,N_13785,N_12645);
nand U15537 (N_15537,N_13628,N_14365);
xnor U15538 (N_15538,N_12837,N_11373);
or U15539 (N_15539,N_11148,N_10416);
and U15540 (N_15540,N_10627,N_10513);
xor U15541 (N_15541,N_13363,N_11750);
and U15542 (N_15542,N_10184,N_14649);
and U15543 (N_15543,N_11438,N_10194);
nand U15544 (N_15544,N_12774,N_14912);
or U15545 (N_15545,N_13808,N_12644);
nand U15546 (N_15546,N_11627,N_13636);
and U15547 (N_15547,N_14523,N_13837);
or U15548 (N_15548,N_10658,N_14648);
or U15549 (N_15549,N_12957,N_14124);
nor U15550 (N_15550,N_14832,N_14645);
nand U15551 (N_15551,N_10681,N_10452);
nor U15552 (N_15552,N_11937,N_12805);
or U15553 (N_15553,N_12978,N_11974);
or U15554 (N_15554,N_10620,N_14717);
nor U15555 (N_15555,N_10826,N_10784);
xnor U15556 (N_15556,N_13219,N_14405);
and U15557 (N_15557,N_12748,N_13020);
nor U15558 (N_15558,N_10392,N_14359);
xor U15559 (N_15559,N_11955,N_10189);
nand U15560 (N_15560,N_10616,N_11726);
and U15561 (N_15561,N_12816,N_13049);
or U15562 (N_15562,N_10634,N_11048);
xor U15563 (N_15563,N_11389,N_10265);
nor U15564 (N_15564,N_13633,N_13401);
nor U15565 (N_15565,N_13238,N_11206);
xor U15566 (N_15566,N_14278,N_12378);
or U15567 (N_15567,N_12560,N_12212);
xor U15568 (N_15568,N_14642,N_12050);
nor U15569 (N_15569,N_12208,N_13051);
or U15570 (N_15570,N_10168,N_10228);
nand U15571 (N_15571,N_10247,N_14289);
xnor U15572 (N_15572,N_12062,N_13453);
xor U15573 (N_15573,N_13597,N_13841);
nor U15574 (N_15574,N_12346,N_14082);
xnor U15575 (N_15575,N_13392,N_11831);
or U15576 (N_15576,N_12971,N_10728);
or U15577 (N_15577,N_10203,N_12214);
nor U15578 (N_15578,N_12089,N_13070);
or U15579 (N_15579,N_11677,N_11137);
xor U15580 (N_15580,N_10445,N_14148);
nand U15581 (N_15581,N_12587,N_14004);
xnor U15582 (N_15582,N_14127,N_10079);
xnor U15583 (N_15583,N_10802,N_14168);
or U15584 (N_15584,N_13007,N_11764);
xor U15585 (N_15585,N_11682,N_12369);
or U15586 (N_15586,N_14628,N_12625);
and U15587 (N_15587,N_11356,N_14892);
nand U15588 (N_15588,N_14228,N_14542);
and U15589 (N_15589,N_13867,N_10603);
or U15590 (N_15590,N_11654,N_11947);
or U15591 (N_15591,N_13529,N_13555);
and U15592 (N_15592,N_14955,N_12243);
nand U15593 (N_15593,N_11174,N_12951);
or U15594 (N_15594,N_10584,N_10190);
xor U15595 (N_15595,N_10514,N_13456);
and U15596 (N_15596,N_11243,N_11404);
nor U15597 (N_15597,N_13713,N_11106);
xnor U15598 (N_15598,N_12511,N_13210);
nor U15599 (N_15599,N_13033,N_11044);
and U15600 (N_15600,N_12007,N_11968);
or U15601 (N_15601,N_12137,N_10208);
nand U15602 (N_15602,N_14788,N_10290);
nor U15603 (N_15603,N_13215,N_14860);
and U15604 (N_15604,N_10218,N_13338);
nor U15605 (N_15605,N_13488,N_13729);
nor U15606 (N_15606,N_10755,N_11012);
xnor U15607 (N_15607,N_14015,N_14275);
nor U15608 (N_15608,N_12700,N_11939);
nand U15609 (N_15609,N_13187,N_10375);
or U15610 (N_15610,N_13192,N_12334);
nand U15611 (N_15611,N_14789,N_10986);
xor U15612 (N_15612,N_13603,N_12798);
nand U15613 (N_15613,N_10697,N_13477);
nor U15614 (N_15614,N_14326,N_12435);
nor U15615 (N_15615,N_10899,N_13961);
and U15616 (N_15616,N_12308,N_13403);
and U15617 (N_15617,N_13779,N_13145);
nand U15618 (N_15618,N_14420,N_12952);
or U15619 (N_15619,N_11889,N_11056);
and U15620 (N_15620,N_14514,N_14329);
xnor U15621 (N_15621,N_14657,N_12434);
xor U15622 (N_15622,N_12885,N_14160);
xor U15623 (N_15623,N_11390,N_12266);
nor U15624 (N_15624,N_12486,N_10897);
nand U15625 (N_15625,N_14529,N_14777);
nor U15626 (N_15626,N_14593,N_11343);
xor U15627 (N_15627,N_12734,N_13055);
nand U15628 (N_15628,N_11641,N_14380);
and U15629 (N_15629,N_10470,N_12091);
nor U15630 (N_15630,N_10708,N_13504);
and U15631 (N_15631,N_13587,N_11448);
nor U15632 (N_15632,N_14569,N_14387);
nand U15633 (N_15633,N_10487,N_13202);
nor U15634 (N_15634,N_10095,N_13158);
nor U15635 (N_15635,N_13653,N_13353);
xnor U15636 (N_15636,N_10748,N_12355);
and U15637 (N_15637,N_11403,N_10111);
and U15638 (N_15638,N_12088,N_13134);
nand U15639 (N_15639,N_12102,N_11530);
nand U15640 (N_15640,N_11005,N_11089);
nand U15641 (N_15641,N_12756,N_11517);
and U15642 (N_15642,N_13188,N_13310);
and U15643 (N_15643,N_10343,N_11942);
and U15644 (N_15644,N_10846,N_13371);
nor U15645 (N_15645,N_14500,N_14293);
or U15646 (N_15646,N_11642,N_11584);
nor U15647 (N_15647,N_11995,N_11608);
and U15648 (N_15648,N_11611,N_10001);
nand U15649 (N_15649,N_12713,N_10702);
nor U15650 (N_15650,N_13189,N_11578);
or U15651 (N_15651,N_10064,N_11248);
or U15652 (N_15652,N_11984,N_12056);
nand U15653 (N_15653,N_12613,N_14638);
xor U15654 (N_15654,N_14558,N_10934);
xor U15655 (N_15655,N_11961,N_11662);
nor U15656 (N_15656,N_14804,N_13047);
nand U15657 (N_15657,N_12589,N_13520);
nand U15658 (N_15658,N_10312,N_12400);
nand U15659 (N_15659,N_10185,N_10365);
nor U15660 (N_15660,N_12852,N_13120);
and U15661 (N_15661,N_12140,N_11600);
and U15662 (N_15662,N_11017,N_11505);
or U15663 (N_15663,N_13099,N_12367);
xnor U15664 (N_15664,N_10511,N_11903);
nand U15665 (N_15665,N_13395,N_11102);
xor U15666 (N_15666,N_13062,N_10422);
xnor U15667 (N_15667,N_12158,N_10564);
nor U15668 (N_15668,N_13465,N_14273);
nor U15669 (N_15669,N_14831,N_14836);
nor U15670 (N_15670,N_11759,N_13236);
xnor U15671 (N_15671,N_13059,N_12554);
nand U15672 (N_15672,N_10659,N_11497);
xor U15673 (N_15673,N_10071,N_10377);
xor U15674 (N_15674,N_12924,N_14068);
and U15675 (N_15675,N_14668,N_12437);
and U15676 (N_15676,N_13993,N_12177);
and U15677 (N_15677,N_14494,N_10456);
nand U15678 (N_15678,N_12488,N_12403);
and U15679 (N_15679,N_13674,N_12000);
nand U15680 (N_15680,N_13506,N_14355);
nor U15681 (N_15681,N_14974,N_14504);
and U15682 (N_15682,N_10004,N_14267);
xor U15683 (N_15683,N_10319,N_14421);
nor U15684 (N_15684,N_10407,N_14393);
nor U15685 (N_15685,N_14828,N_14968);
xor U15686 (N_15686,N_11957,N_10520);
nand U15687 (N_15687,N_12044,N_14153);
nor U15688 (N_15688,N_11845,N_11650);
nor U15689 (N_15689,N_10585,N_10171);
or U15690 (N_15690,N_10115,N_11131);
nand U15691 (N_15691,N_13252,N_14309);
or U15692 (N_15692,N_11126,N_10254);
nand U15693 (N_15693,N_12688,N_13689);
and U15694 (N_15694,N_10038,N_10793);
nor U15695 (N_15695,N_10325,N_10328);
and U15696 (N_15696,N_13281,N_10460);
xor U15697 (N_15697,N_10214,N_12629);
xor U15698 (N_15698,N_14741,N_12338);
and U15699 (N_15699,N_12399,N_12482);
xnor U15700 (N_15700,N_12921,N_13129);
nor U15701 (N_15701,N_10872,N_12772);
nand U15702 (N_15702,N_11594,N_13298);
nor U15703 (N_15703,N_10050,N_11464);
nand U15704 (N_15704,N_13150,N_11217);
nand U15705 (N_15705,N_12111,N_11541);
and U15706 (N_15706,N_11701,N_11242);
xnor U15707 (N_15707,N_10024,N_10672);
nor U15708 (N_15708,N_11965,N_13037);
or U15709 (N_15709,N_10997,N_11194);
nand U15710 (N_15710,N_11078,N_14473);
or U15711 (N_15711,N_14422,N_11401);
and U15712 (N_15712,N_11493,N_12045);
nand U15713 (N_15713,N_13549,N_11380);
or U15714 (N_15714,N_14767,N_12591);
nand U15715 (N_15715,N_14620,N_13318);
nand U15716 (N_15716,N_14938,N_10287);
xor U15717 (N_15717,N_12164,N_10785);
and U15718 (N_15718,N_14181,N_12787);
nand U15719 (N_15719,N_10833,N_11583);
nand U15720 (N_15720,N_10337,N_14902);
and U15721 (N_15721,N_14706,N_14729);
or U15722 (N_15722,N_11302,N_12812);
xnor U15723 (N_15723,N_12124,N_13541);
and U15724 (N_15724,N_13058,N_11953);
and U15725 (N_15725,N_12849,N_14439);
and U15726 (N_15726,N_11027,N_10367);
nor U15727 (N_15727,N_13850,N_10789);
nand U15728 (N_15728,N_14252,N_12366);
nor U15729 (N_15729,N_11339,N_13548);
nand U15730 (N_15730,N_10402,N_11568);
and U15731 (N_15731,N_13657,N_10573);
xor U15732 (N_15732,N_11857,N_12524);
xor U15733 (N_15733,N_10340,N_11103);
nand U15734 (N_15734,N_13960,N_12316);
nor U15735 (N_15735,N_13409,N_10142);
nor U15736 (N_15736,N_14936,N_13216);
or U15737 (N_15737,N_13819,N_12423);
or U15738 (N_15738,N_12408,N_14113);
nor U15739 (N_15739,N_11959,N_11368);
nand U15740 (N_15740,N_12646,N_12549);
nor U15741 (N_15741,N_14992,N_10608);
or U15742 (N_15742,N_11213,N_11460);
xor U15743 (N_15743,N_14903,N_14564);
nand U15744 (N_15744,N_13211,N_14517);
or U15745 (N_15745,N_13795,N_14805);
or U15746 (N_15746,N_12085,N_10246);
or U15747 (N_15747,N_12103,N_10014);
nand U15748 (N_15748,N_14809,N_14586);
nor U15749 (N_15749,N_14748,N_13711);
nand U15750 (N_15750,N_10180,N_14245);
nor U15751 (N_15751,N_13282,N_11544);
and U15752 (N_15752,N_10118,N_13354);
and U15753 (N_15753,N_11613,N_13981);
nand U15754 (N_15754,N_12767,N_13817);
nor U15755 (N_15755,N_11218,N_13972);
or U15756 (N_15756,N_11760,N_14821);
or U15757 (N_15757,N_14166,N_14945);
and U15758 (N_15758,N_11789,N_13088);
nor U15759 (N_15759,N_12884,N_11835);
xnor U15760 (N_15760,N_13575,N_10143);
or U15761 (N_15761,N_10224,N_12441);
or U15762 (N_15762,N_11618,N_13695);
or U15763 (N_15763,N_12684,N_13384);
nand U15764 (N_15764,N_11971,N_14435);
xnor U15765 (N_15765,N_10486,N_11428);
nor U15766 (N_15766,N_11098,N_12345);
nor U15767 (N_15767,N_11241,N_13266);
or U15768 (N_15768,N_12743,N_10545);
xnor U15769 (N_15769,N_12186,N_13658);
nor U15770 (N_15770,N_12586,N_12600);
nor U15771 (N_15771,N_10636,N_11870);
nor U15772 (N_15772,N_12010,N_14904);
and U15773 (N_15773,N_12920,N_12806);
nand U15774 (N_15774,N_13369,N_12200);
xor U15775 (N_15775,N_10036,N_12751);
xnor U15776 (N_15776,N_13660,N_12530);
xnor U15777 (N_15777,N_11192,N_14540);
nor U15778 (N_15778,N_14907,N_11989);
xnor U15779 (N_15779,N_11166,N_14112);
or U15780 (N_15780,N_11640,N_11276);
nand U15781 (N_15781,N_14206,N_14961);
or U15782 (N_15782,N_12083,N_14199);
xnor U15783 (N_15783,N_12365,N_11066);
and U15784 (N_15784,N_10537,N_12307);
and U15785 (N_15785,N_13481,N_14723);
nor U15786 (N_15786,N_10415,N_10761);
nor U15787 (N_15787,N_14091,N_12674);
nand U15788 (N_15788,N_14727,N_12321);
and U15789 (N_15789,N_10973,N_13613);
xnor U15790 (N_15790,N_14434,N_13146);
nor U15791 (N_15791,N_10667,N_11988);
or U15792 (N_15792,N_13426,N_11712);
or U15793 (N_15793,N_14909,N_12136);
nand U15794 (N_15794,N_11793,N_11291);
xor U15795 (N_15795,N_14104,N_13916);
nand U15796 (N_15796,N_12236,N_14118);
nand U15797 (N_15797,N_14731,N_11145);
xor U15798 (N_15798,N_10811,N_11021);
xnor U15799 (N_15799,N_13534,N_11704);
xor U15800 (N_15800,N_11279,N_11205);
nor U15801 (N_15801,N_11545,N_11503);
xor U15802 (N_15802,N_12231,N_10629);
or U15803 (N_15803,N_11780,N_13482);
nand U15804 (N_15804,N_12758,N_10630);
or U15805 (N_15805,N_14495,N_11306);
or U15806 (N_15806,N_14618,N_14195);
and U15807 (N_15807,N_11696,N_12782);
nand U15808 (N_15808,N_13154,N_14964);
and U15809 (N_15809,N_12580,N_13267);
or U15810 (N_15810,N_10300,N_11195);
or U15811 (N_15811,N_13810,N_13183);
xor U15812 (N_15812,N_12715,N_14138);
nor U15813 (N_15813,N_11483,N_11986);
or U15814 (N_15814,N_13478,N_11309);
nor U15815 (N_15815,N_11521,N_14507);
nand U15816 (N_15816,N_13225,N_12042);
nand U15817 (N_15817,N_10586,N_13212);
and U15818 (N_15818,N_10138,N_10140);
nand U15819 (N_15819,N_14795,N_12814);
and U15820 (N_15820,N_10245,N_13314);
xor U15821 (N_15821,N_11396,N_13733);
xnor U15822 (N_15822,N_10773,N_14981);
nor U15823 (N_15823,N_14092,N_11286);
nand U15824 (N_15824,N_12944,N_12075);
xnor U15825 (N_15825,N_12376,N_10715);
nor U15826 (N_15826,N_11379,N_13563);
nor U15827 (N_15827,N_11581,N_13406);
nor U15828 (N_15828,N_14520,N_11147);
or U15829 (N_15829,N_10178,N_11207);
nand U15830 (N_15830,N_11598,N_12773);
or U15831 (N_15831,N_12855,N_13172);
or U15832 (N_15832,N_14475,N_12651);
xnor U15833 (N_15833,N_13662,N_10141);
and U15834 (N_15834,N_14204,N_12661);
nand U15835 (N_15835,N_13386,N_11510);
nand U15836 (N_15836,N_14994,N_13455);
nor U15837 (N_15837,N_11810,N_11739);
xor U15838 (N_15838,N_14175,N_10827);
and U15839 (N_15839,N_12633,N_13138);
and U15840 (N_15840,N_12932,N_14510);
nand U15841 (N_15841,N_14084,N_14342);
nand U15842 (N_15842,N_12967,N_14989);
or U15843 (N_15843,N_11330,N_13988);
or U15844 (N_15844,N_13544,N_12317);
xnor U15845 (N_15845,N_10721,N_14448);
nor U15846 (N_15846,N_11065,N_12159);
and U15847 (N_15847,N_10882,N_14525);
nor U15848 (N_15848,N_14834,N_14592);
nand U15849 (N_15849,N_13553,N_11282);
or U15850 (N_15850,N_14173,N_14051);
xor U15851 (N_15851,N_11341,N_13261);
nor U15852 (N_15852,N_14370,N_12609);
nor U15853 (N_15853,N_13319,N_11779);
nand U15854 (N_15854,N_12248,N_13094);
xnor U15855 (N_15855,N_10116,N_13474);
xnor U15856 (N_15856,N_12142,N_12529);
nor U15857 (N_15857,N_14709,N_14756);
and U15858 (N_15858,N_12057,N_13358);
and U15859 (N_15859,N_11617,N_12728);
xnor U15860 (N_15860,N_12041,N_10825);
or U15861 (N_15861,N_13673,N_14581);
or U15862 (N_15862,N_11173,N_11371);
xnor U15863 (N_15863,N_13965,N_10026);
xor U15864 (N_15864,N_11463,N_14298);
nand U15865 (N_15865,N_14006,N_11656);
nand U15866 (N_15866,N_12059,N_14679);
nor U15867 (N_15867,N_10099,N_14582);
or U15868 (N_15868,N_11208,N_14934);
nand U15869 (N_15869,N_13209,N_11577);
nor U15870 (N_15870,N_11419,N_13341);
nor U15871 (N_15871,N_14557,N_11958);
nand U15872 (N_15872,N_14114,N_11529);
or U15873 (N_15873,N_12279,N_12179);
and U15874 (N_15874,N_14258,N_10075);
nor U15875 (N_15875,N_14776,N_12289);
or U15876 (N_15876,N_14627,N_11400);
or U15877 (N_15877,N_14881,N_11399);
nand U15878 (N_15878,N_11900,N_10859);
or U15879 (N_15879,N_13031,N_11825);
nand U15880 (N_15880,N_14270,N_12335);
and U15881 (N_15881,N_13757,N_10408);
xor U15882 (N_15882,N_13490,N_10706);
nand U15883 (N_15883,N_10017,N_12551);
nor U15884 (N_15884,N_11638,N_10943);
or U15885 (N_15885,N_12786,N_14489);
xor U15886 (N_15886,N_13206,N_10427);
nand U15887 (N_15887,N_10710,N_12749);
nand U15888 (N_15888,N_11763,N_12216);
and U15889 (N_15889,N_13171,N_14056);
and U15890 (N_15890,N_12386,N_12426);
xor U15891 (N_15891,N_13362,N_13090);
nor U15892 (N_15892,N_13348,N_13612);
nor U15893 (N_15893,N_12304,N_13934);
nand U15894 (N_15894,N_14462,N_12047);
or U15895 (N_15895,N_10905,N_14279);
and U15896 (N_15896,N_11786,N_13741);
nand U15897 (N_15897,N_14585,N_11543);
nand U15898 (N_15898,N_14686,N_10491);
nor U15899 (N_15899,N_12838,N_10524);
xor U15900 (N_15900,N_12620,N_11822);
nor U15901 (N_15901,N_13317,N_13601);
nand U15902 (N_15902,N_11856,N_11011);
nor U15903 (N_15903,N_13235,N_10803);
or U15904 (N_15904,N_10661,N_13943);
or U15905 (N_15905,N_13257,N_12452);
nand U15906 (N_15906,N_11755,N_14358);
and U15907 (N_15907,N_12794,N_10856);
nor U15908 (N_15908,N_13634,N_12875);
xor U15909 (N_15909,N_12975,N_14096);
nand U15910 (N_15910,N_14022,N_14080);
and U15911 (N_15911,N_11260,N_10181);
nor U15912 (N_15912,N_12347,N_14674);
nor U15913 (N_15913,N_10948,N_10894);
xor U15914 (N_15914,N_12324,N_14315);
or U15915 (N_15915,N_10371,N_12063);
and U15916 (N_15916,N_14843,N_12196);
xor U15917 (N_15917,N_12340,N_11072);
nand U15918 (N_15918,N_13571,N_11881);
nand U15919 (N_15919,N_11289,N_14251);
nand U15920 (N_15920,N_11837,N_10711);
nor U15921 (N_15921,N_11383,N_10104);
xnor U15922 (N_15922,N_13110,N_12914);
nor U15923 (N_15923,N_11684,N_12430);
nand U15924 (N_15924,N_13858,N_12708);
nand U15925 (N_15925,N_11259,N_13333);
or U15926 (N_15926,N_12900,N_13402);
and U15927 (N_15927,N_13585,N_12493);
xor U15928 (N_15928,N_13389,N_11533);
xnor U15929 (N_15929,N_10578,N_11982);
nand U15930 (N_15930,N_13942,N_13582);
nand U15931 (N_15931,N_13714,N_13692);
nand U15932 (N_15932,N_13468,N_12172);
or U15933 (N_15933,N_14993,N_12055);
nor U15934 (N_15934,N_14425,N_10951);
nand U15935 (N_15935,N_14050,N_10863);
or U15936 (N_15936,N_14272,N_10763);
xnor U15937 (N_15937,N_12255,N_13028);
and U15938 (N_15938,N_10073,N_10714);
nor U15939 (N_15939,N_11470,N_14929);
nor U15940 (N_15940,N_11830,N_10444);
xor U15941 (N_15941,N_14976,N_14710);
nand U15942 (N_15942,N_14119,N_12635);
nand U15943 (N_15943,N_10019,N_10162);
nand U15944 (N_15944,N_14900,N_12979);
xor U15945 (N_15945,N_10455,N_10713);
nand U15946 (N_15946,N_13806,N_12525);
and U15947 (N_15947,N_10604,N_10557);
and U15948 (N_15948,N_10136,N_11657);
nand U15949 (N_15949,N_11074,N_11833);
or U15950 (N_15950,N_11278,N_13945);
nand U15951 (N_15951,N_12948,N_13434);
nor U15952 (N_15952,N_12815,N_10033);
nor U15953 (N_15953,N_12505,N_11197);
nor U15954 (N_15954,N_13264,N_14813);
and U15955 (N_15955,N_14890,N_13286);
xnor U15956 (N_15956,N_14376,N_12016);
and U15957 (N_15957,N_14120,N_10106);
and U15958 (N_15958,N_13221,N_14100);
or U15959 (N_15959,N_12976,N_11301);
xnor U15960 (N_15960,N_10259,N_11655);
nand U15961 (N_15961,N_13507,N_11688);
or U15962 (N_15962,N_11484,N_12776);
xor U15963 (N_15963,N_10906,N_12401);
nor U15964 (N_15964,N_12939,N_11292);
nor U15965 (N_15965,N_12851,N_14328);
and U15966 (N_15966,N_14720,N_12861);
or U15967 (N_15967,N_12719,N_14363);
nand U15968 (N_15968,N_11047,N_12247);
nand U15969 (N_15969,N_14937,N_13772);
xnor U15970 (N_15970,N_11481,N_10357);
and U15971 (N_15971,N_13245,N_12299);
nand U15972 (N_15972,N_14311,N_11519);
nor U15973 (N_15973,N_13388,N_10149);
and U15974 (N_15974,N_14616,N_12389);
and U15975 (N_15975,N_14959,N_10828);
or U15976 (N_15976,N_14316,N_14606);
nand U15977 (N_15977,N_12657,N_11711);
nand U15978 (N_15978,N_14069,N_14097);
nor U15979 (N_15979,N_14296,N_11773);
nand U15980 (N_15980,N_14179,N_12539);
or U15981 (N_15981,N_13015,N_13606);
nand U15982 (N_15982,N_11865,N_10437);
or U15983 (N_15983,N_14599,N_11283);
nand U15984 (N_15984,N_12550,N_11795);
nand U15985 (N_15985,N_13880,N_10944);
xnor U15986 (N_15986,N_10503,N_11949);
nand U15987 (N_15987,N_12585,N_14565);
xnor U15988 (N_15988,N_12429,N_12046);
and U15989 (N_15989,N_14677,N_14522);
and U15990 (N_15990,N_11522,N_12640);
or U15991 (N_15991,N_14782,N_11920);
nor U15992 (N_15992,N_13838,N_10150);
and U15993 (N_15993,N_13905,N_14220);
xnor U15994 (N_15994,N_11621,N_10591);
nor U15995 (N_15995,N_12122,N_14928);
nor U15996 (N_15996,N_11504,N_10391);
or U15997 (N_15997,N_11042,N_14664);
and U15998 (N_15998,N_14154,N_10410);
xor U15999 (N_15999,N_10120,N_12546);
or U16000 (N_16000,N_11201,N_14519);
or U16001 (N_16001,N_14288,N_12427);
nand U16002 (N_16002,N_14060,N_10354);
or U16003 (N_16003,N_10177,N_14632);
nor U16004 (N_16004,N_13609,N_14654);
nor U16005 (N_16005,N_12107,N_11409);
nor U16006 (N_16006,N_13622,N_12167);
and U16007 (N_16007,N_10157,N_12374);
and U16008 (N_16008,N_10666,N_14238);
and U16009 (N_16009,N_13130,N_12744);
xnor U16010 (N_16010,N_14692,N_12453);
nor U16011 (N_16011,N_12272,N_11169);
or U16012 (N_16012,N_14746,N_14833);
xor U16013 (N_16013,N_10525,N_11603);
xor U16014 (N_16014,N_12988,N_13294);
and U16015 (N_16015,N_11349,N_14849);
nor U16016 (N_16016,N_10628,N_12981);
xnor U16017 (N_16017,N_11477,N_11969);
nand U16018 (N_16018,N_12336,N_10473);
or U16019 (N_16019,N_14623,N_10027);
and U16020 (N_16020,N_13820,N_10173);
xnor U16021 (N_16021,N_10380,N_10497);
nand U16022 (N_16022,N_11142,N_14484);
nand U16023 (N_16023,N_14044,N_11471);
nand U16024 (N_16024,N_10350,N_12650);
xnor U16025 (N_16025,N_13532,N_11717);
or U16026 (N_16026,N_12958,N_11144);
nor U16027 (N_16027,N_12596,N_11168);
nor U16028 (N_16028,N_14672,N_10592);
and U16029 (N_16029,N_12969,N_10423);
or U16030 (N_16030,N_13375,N_12514);
or U16031 (N_16031,N_11615,N_14770);
nand U16032 (N_16032,N_14797,N_11817);
nor U16033 (N_16033,N_12801,N_10770);
nor U16034 (N_16034,N_12380,N_12680);
nor U16035 (N_16035,N_13641,N_14895);
nand U16036 (N_16036,N_13246,N_14397);
and U16037 (N_16037,N_13280,N_11807);
or U16038 (N_16038,N_10924,N_11509);
nor U16039 (N_16039,N_10363,N_11255);
or U16040 (N_16040,N_13463,N_11055);
and U16041 (N_16041,N_14414,N_14467);
and U16042 (N_16042,N_10742,N_14803);
or U16043 (N_16043,N_10007,N_11030);
and U16044 (N_16044,N_14117,N_12354);
and U16045 (N_16045,N_12388,N_10352);
or U16046 (N_16046,N_11751,N_13010);
nand U16047 (N_16047,N_11406,N_11768);
nor U16048 (N_16048,N_14563,N_13023);
nand U16049 (N_16049,N_14758,N_13048);
or U16050 (N_16050,N_10840,N_10990);
nor U16051 (N_16051,N_12965,N_13813);
or U16052 (N_16052,N_10096,N_10401);
nand U16053 (N_16053,N_12716,N_10867);
xor U16054 (N_16054,N_11297,N_11922);
nor U16055 (N_16055,N_14643,N_13071);
nand U16056 (N_16056,N_13604,N_14259);
or U16057 (N_16057,N_10040,N_11412);
or U16058 (N_16058,N_14318,N_12464);
nor U16059 (N_16059,N_13074,N_12984);
nor U16060 (N_16060,N_13915,N_12170);
nand U16061 (N_16061,N_12829,N_12548);
or U16062 (N_16062,N_13693,N_11824);
and U16063 (N_16063,N_11164,N_13744);
xnor U16064 (N_16064,N_12785,N_13244);
or U16065 (N_16065,N_11811,N_14634);
and U16066 (N_16066,N_14703,N_10283);
or U16067 (N_16067,N_12235,N_14253);
or U16068 (N_16068,N_12968,N_11710);
or U16069 (N_16069,N_14820,N_11155);
or U16070 (N_16070,N_14016,N_14145);
or U16071 (N_16071,N_12503,N_10374);
or U16072 (N_16072,N_10903,N_12298);
or U16073 (N_16073,N_12178,N_10278);
nor U16074 (N_16074,N_10750,N_13324);
nand U16075 (N_16075,N_12204,N_10230);
or U16076 (N_16076,N_14330,N_11370);
nor U16077 (N_16077,N_11625,N_10097);
xor U16078 (N_16078,N_12959,N_13466);
nand U16079 (N_16079,N_11490,N_11643);
nand U16080 (N_16080,N_13941,N_11014);
or U16081 (N_16081,N_12973,N_13891);
nor U16082 (N_16082,N_11068,N_10176);
or U16083 (N_16083,N_13361,N_10901);
and U16084 (N_16084,N_11002,N_13830);
nor U16085 (N_16085,N_13672,N_12496);
nand U16086 (N_16086,N_13763,N_13440);
nor U16087 (N_16087,N_13906,N_13884);
nor U16088 (N_16088,N_13875,N_10240);
xnor U16089 (N_16089,N_11678,N_14670);
or U16090 (N_16090,N_13043,N_14209);
and U16091 (N_16091,N_12564,N_14830);
or U16092 (N_16092,N_13703,N_10687);
or U16093 (N_16093,N_11327,N_14262);
nor U16094 (N_16094,N_10210,N_12206);
nor U16095 (N_16095,N_14011,N_13797);
nor U16096 (N_16096,N_14629,N_12329);
xor U16097 (N_16097,N_12668,N_14611);
and U16098 (N_16098,N_11064,N_10505);
and U16099 (N_16099,N_12444,N_12567);
or U16100 (N_16100,N_14946,N_10324);
or U16101 (N_16101,N_12145,N_10689);
xnor U16102 (N_16102,N_10705,N_10215);
nor U16103 (N_16103,N_13647,N_11132);
and U16104 (N_16104,N_13978,N_13052);
xnor U16105 (N_16105,N_14436,N_11134);
xor U16106 (N_16106,N_10030,N_11893);
nand U16107 (N_16107,N_13998,N_11374);
and U16108 (N_16108,N_10610,N_10023);
xnor U16109 (N_16109,N_12512,N_11777);
or U16110 (N_16110,N_11908,N_13115);
or U16111 (N_16111,N_13704,N_10009);
nand U16112 (N_16112,N_11120,N_10390);
and U16113 (N_16113,N_10798,N_12545);
xnor U16114 (N_16114,N_14498,N_14219);
nand U16115 (N_16115,N_13424,N_12775);
or U16116 (N_16116,N_11754,N_12822);
nand U16117 (N_16117,N_10393,N_14009);
nor U16118 (N_16118,N_13640,N_14445);
and U16119 (N_16119,N_13614,N_10132);
nor U16120 (N_16120,N_14008,N_14350);
or U16121 (N_16121,N_14053,N_11018);
or U16122 (N_16122,N_11506,N_11653);
xnor U16123 (N_16123,N_11190,N_12465);
xor U16124 (N_16124,N_12173,N_14858);
nand U16125 (N_16125,N_10844,N_10795);
nand U16126 (N_16126,N_11424,N_13578);
xor U16127 (N_16127,N_12081,N_14300);
nand U16128 (N_16128,N_13199,N_11727);
nor U16129 (N_16129,N_12871,N_12487);
or U16130 (N_16130,N_11905,N_13445);
nor U16131 (N_16131,N_14461,N_13546);
or U16132 (N_16132,N_11679,N_12497);
or U16133 (N_16133,N_10722,N_13309);
xnor U16134 (N_16134,N_11848,N_12666);
and U16135 (N_16135,N_10298,N_14192);
nand U16136 (N_16136,N_11353,N_14385);
nand U16137 (N_16137,N_10133,N_11234);
and U16138 (N_16138,N_12788,N_14615);
nand U16139 (N_16139,N_12802,N_12281);
nor U16140 (N_16140,N_11692,N_11694);
nor U16141 (N_16141,N_12238,N_12839);
nand U16142 (N_16142,N_10558,N_11999);
and U16143 (N_16143,N_11787,N_11158);
nor U16144 (N_16144,N_10223,N_12291);
and U16145 (N_16145,N_10041,N_10128);
and U16146 (N_16146,N_13081,N_10767);
and U16147 (N_16147,N_11020,N_10074);
or U16148 (N_16148,N_13355,N_14837);
or U16149 (N_16149,N_10155,N_11336);
or U16150 (N_16150,N_12854,N_10239);
xnor U16151 (N_16151,N_11593,N_10273);
xor U16152 (N_16152,N_12080,N_13831);
or U16153 (N_16153,N_10786,N_14485);
or U16154 (N_16154,N_12277,N_13924);
or U16155 (N_16155,N_12368,N_10808);
and U16156 (N_16156,N_12647,N_13527);
and U16157 (N_16157,N_13376,N_14086);
xor U16158 (N_16158,N_11705,N_14465);
or U16159 (N_16159,N_10090,N_13347);
nand U16160 (N_16160,N_11159,N_10232);
nand U16161 (N_16161,N_13311,N_12603);
xnor U16162 (N_16162,N_11841,N_14497);
or U16163 (N_16163,N_13234,N_12725);
xnor U16164 (N_16164,N_13528,N_12130);
nor U16165 (N_16165,N_14135,N_10499);
and U16166 (N_16166,N_13137,N_10430);
nor U16167 (N_16167,N_13408,N_14418);
and U16168 (N_16168,N_14597,N_12123);
or U16169 (N_16169,N_10946,N_13009);
nand U16170 (N_16170,N_14536,N_12931);
or U16171 (N_16171,N_14978,N_10941);
xor U16172 (N_16172,N_13418,N_14303);
or U16173 (N_16173,N_11567,N_13971);
and U16174 (N_16174,N_12824,N_14071);
nand U16175 (N_16175,N_12381,N_14472);
xor U16176 (N_16176,N_11138,N_11725);
nor U16177 (N_16177,N_11911,N_13767);
nor U16178 (N_16178,N_10332,N_12519);
and U16179 (N_16179,N_10639,N_14428);
or U16180 (N_16180,N_11944,N_13411);
or U16181 (N_16181,N_11480,N_10942);
and U16182 (N_16182,N_11702,N_14054);
xor U16183 (N_16183,N_14469,N_12148);
or U16184 (N_16184,N_11288,N_14048);
nand U16185 (N_16185,N_13032,N_14088);
nor U16186 (N_16186,N_10342,N_13754);
nand U16187 (N_16187,N_14721,N_14637);
or U16188 (N_16188,N_13365,N_14604);
nand U16189 (N_16189,N_12641,N_14772);
and U16190 (N_16190,N_10012,N_14583);
nor U16191 (N_16191,N_12803,N_14956);
or U16192 (N_16192,N_14301,N_10202);
nor U16193 (N_16193,N_14794,N_11334);
xor U16194 (N_16194,N_11123,N_11660);
nor U16195 (N_16195,N_14261,N_14687);
nand U16196 (N_16196,N_10962,N_10640);
or U16197 (N_16197,N_11070,N_14302);
nand U16198 (N_16198,N_14018,N_11774);
and U16199 (N_16199,N_13734,N_13413);
nand U16200 (N_16200,N_14235,N_11762);
xor U16201 (N_16201,N_14850,N_14952);
xnor U16202 (N_16202,N_10866,N_10723);
xnor U16203 (N_16203,N_11776,N_11130);
xnor U16204 (N_16204,N_13788,N_14823);
nor U16205 (N_16205,N_14320,N_13277);
nand U16206 (N_16206,N_10061,N_11664);
and U16207 (N_16207,N_11454,N_11233);
nand U16208 (N_16208,N_10871,N_11767);
nand U16209 (N_16209,N_10961,N_10800);
nor U16210 (N_16210,N_13502,N_14074);
xnor U16211 (N_16211,N_14971,N_11812);
nand U16212 (N_16212,N_12697,N_13255);
xor U16213 (N_16213,N_11609,N_13075);
nand U16214 (N_16214,N_12333,N_12656);
nor U16215 (N_16215,N_10085,N_13269);
and U16216 (N_16216,N_14499,N_13491);
nand U16217 (N_16217,N_14131,N_13428);
or U16218 (N_16218,N_14774,N_13564);
or U16219 (N_16219,N_14661,N_10372);
nor U16220 (N_16220,N_12584,N_13017);
or U16221 (N_16221,N_11104,N_12224);
nand U16222 (N_16222,N_13696,N_12768);
xnor U16223 (N_16223,N_11347,N_12087);
xor U16224 (N_16224,N_14685,N_14682);
and U16225 (N_16225,N_13262,N_11676);
xor U16226 (N_16226,N_14020,N_14085);
xnor U16227 (N_16227,N_10654,N_13250);
xor U16228 (N_16228,N_11254,N_14134);
xnor U16229 (N_16229,N_11934,N_12405);
nor U16230 (N_16230,N_13946,N_11410);
and U16231 (N_16231,N_13483,N_12419);
nor U16232 (N_16232,N_14663,N_14130);
or U16233 (N_16233,N_12472,N_13878);
xor U16234 (N_16234,N_13577,N_10083);
xor U16235 (N_16235,N_12483,N_11601);
nor U16236 (N_16236,N_11752,N_14765);
or U16237 (N_16237,N_11632,N_12223);
nor U16238 (N_16238,N_13931,N_12404);
or U16239 (N_16239,N_12054,N_11885);
or U16240 (N_16240,N_10820,N_14733);
or U16241 (N_16241,N_10425,N_13537);
or U16242 (N_16242,N_13454,N_10500);
xor U16243 (N_16243,N_10008,N_12791);
or U16244 (N_16244,N_10125,N_11766);
xor U16245 (N_16245,N_11513,N_13926);
nand U16246 (N_16246,N_10878,N_12877);
nand U16247 (N_16247,N_12431,N_12614);
and U16248 (N_16248,N_11778,N_14988);
and U16249 (N_16249,N_10387,N_14922);
or U16250 (N_16250,N_14651,N_13876);
nand U16251 (N_16251,N_12923,N_14450);
nand U16252 (N_16252,N_13040,N_11211);
nand U16253 (N_16253,N_11143,N_14061);
and U16254 (N_16254,N_12006,N_11118);
and U16255 (N_16255,N_12211,N_11122);
and U16256 (N_16256,N_11718,N_11269);
xnor U16257 (N_16257,N_13917,N_12943);
or U16258 (N_16258,N_11973,N_13957);
xnor U16259 (N_16259,N_14364,N_13868);
nor U16260 (N_16260,N_11794,N_10084);
or U16261 (N_16261,N_13896,N_10707);
nor U16262 (N_16262,N_10032,N_13740);
nor U16263 (N_16263,N_11887,N_14773);
nand U16264 (N_16264,N_11753,N_11133);
and U16265 (N_16265,N_11023,N_10348);
xor U16266 (N_16266,N_14039,N_14694);
or U16267 (N_16267,N_12963,N_13761);
or U16268 (N_16268,N_12014,N_14876);
xnor U16269 (N_16269,N_14995,N_10569);
xnor U16270 (N_16270,N_12162,N_13472);
nand U16271 (N_16271,N_14786,N_12541);
xor U16272 (N_16272,N_14571,N_13224);
xnor U16273 (N_16273,N_14234,N_13557);
and U16274 (N_16274,N_13728,N_11687);
and U16275 (N_16275,N_10574,N_13416);
nand U16276 (N_16276,N_12870,N_11783);
and U16277 (N_16277,N_14345,N_10301);
xnor U16278 (N_16278,N_10738,N_10829);
or U16279 (N_16279,N_10648,N_14409);
nand U16280 (N_16280,N_11571,N_13706);
nand U16281 (N_16281,N_10288,N_10812);
or U16282 (N_16282,N_14202,N_12590);
or U16283 (N_16283,N_13654,N_11161);
nand U16284 (N_16284,N_12887,N_12949);
nor U16285 (N_16285,N_12926,N_14579);
or U16286 (N_16286,N_11198,N_10276);
nand U16287 (N_16287,N_10989,N_14182);
nor U16288 (N_16288,N_14715,N_13069);
nor U16289 (N_16289,N_12265,N_10799);
nor U16290 (N_16290,N_14191,N_11285);
and U16291 (N_16291,N_13999,N_14998);
xor U16292 (N_16292,N_13845,N_10612);
nor U16293 (N_16293,N_13629,N_11386);
nor U16294 (N_16294,N_14470,N_12421);
nor U16295 (N_16295,N_10954,N_10275);
or U16296 (N_16296,N_12899,N_10679);
or U16297 (N_16297,N_10843,N_10351);
xor U16298 (N_16298,N_14996,N_14899);
or U16299 (N_16299,N_13165,N_11141);
or U16300 (N_16300,N_11898,N_12402);
nand U16301 (N_16301,N_10680,N_13648);
xnor U16302 (N_16302,N_10673,N_14290);
or U16303 (N_16303,N_10055,N_11796);
nor U16304 (N_16304,N_10749,N_11829);
nand U16305 (N_16305,N_11117,N_11086);
nand U16306 (N_16306,N_10794,N_10015);
and U16307 (N_16307,N_14481,N_11091);
xor U16308 (N_16308,N_13790,N_11964);
xor U16309 (N_16309,N_12876,N_10252);
nor U16310 (N_16310,N_13718,N_11154);
xor U16311 (N_16311,N_12936,N_12909);
or U16312 (N_16312,N_12808,N_11788);
xor U16313 (N_16313,N_10052,N_14194);
nand U16314 (N_16314,N_10219,N_13857);
or U16315 (N_16315,N_14402,N_12445);
nand U16316 (N_16316,N_12160,N_14636);
nand U16317 (N_16317,N_14816,N_14969);
and U16318 (N_16318,N_12731,N_12699);
and U16319 (N_16319,N_12439,N_12448);
nand U16320 (N_16320,N_13743,N_11402);
or U16321 (N_16321,N_14281,N_11331);
and U16322 (N_16322,N_14178,N_14449);
xor U16323 (N_16323,N_13973,N_12986);
or U16324 (N_16324,N_11479,N_11775);
nand U16325 (N_16325,N_10547,N_12721);
nor U16326 (N_16326,N_11022,N_10045);
nor U16327 (N_16327,N_13559,N_11843);
nand U16328 (N_16328,N_10346,N_12720);
or U16329 (N_16329,N_12193,N_14327);
and U16330 (N_16330,N_13708,N_12706);
and U16331 (N_16331,N_14951,N_11321);
and U16332 (N_16332,N_11894,N_12879);
xnor U16333 (N_16333,N_14921,N_13531);
nand U16334 (N_16334,N_11945,N_10135);
nand U16335 (N_16335,N_10936,N_14874);
nand U16336 (N_16336,N_10179,N_12631);
nor U16337 (N_16337,N_12663,N_14340);
nand U16338 (N_16338,N_13974,N_11004);
or U16339 (N_16339,N_12129,N_14935);
nor U16340 (N_16340,N_14596,N_11620);
xnor U16341 (N_16341,N_11323,N_11674);
or U16342 (N_16342,N_10571,N_11036);
xnor U16343 (N_16343,N_13379,N_14443);
nand U16344 (N_16344,N_10237,N_12513);
nor U16345 (N_16345,N_12225,N_12105);
nor U16346 (N_16346,N_11559,N_12820);
or U16347 (N_16347,N_13568,N_12765);
or U16348 (N_16348,N_14090,N_14897);
nor U16349 (N_16349,N_11035,N_11992);
or U16350 (N_16350,N_11149,N_12886);
xnor U16351 (N_16351,N_13391,N_11398);
xnor U16352 (N_16352,N_13762,N_14600);
or U16353 (N_16353,N_12739,N_13060);
xor U16354 (N_16354,N_13798,N_10816);
nor U16355 (N_16355,N_13562,N_13661);
nand U16356 (N_16356,N_12649,N_14690);
or U16357 (N_16357,N_13707,N_14550);
nor U16358 (N_16358,N_14377,N_14716);
xor U16359 (N_16359,N_10395,N_14109);
xnor U16360 (N_16360,N_14829,N_10459);
and U16361 (N_16361,N_12363,N_12499);
nor U16362 (N_16362,N_11203,N_13894);
xnor U16363 (N_16363,N_13320,N_12005);
xor U16364 (N_16364,N_12072,N_12778);
nand U16365 (N_16365,N_10703,N_13131);
xor U16366 (N_16366,N_10994,N_13457);
or U16367 (N_16367,N_13699,N_11423);
or U16368 (N_16368,N_13832,N_14552);
nor U16369 (N_16369,N_11425,N_11478);
or U16370 (N_16370,N_10782,N_10732);
nand U16371 (N_16371,N_10002,N_12213);
nand U16372 (N_16372,N_10144,N_10568);
and U16373 (N_16373,N_12398,N_12106);
or U16374 (N_16374,N_12872,N_13530);
or U16375 (N_16375,N_14408,N_13113);
or U16376 (N_16376,N_10344,N_10366);
or U16377 (N_16377,N_13554,N_13576);
xor U16378 (N_16378,N_10898,N_11667);
and U16379 (N_16379,N_14241,N_14882);
nand U16380 (N_16380,N_13903,N_14348);
or U16381 (N_16381,N_10059,N_12741);
or U16382 (N_16382,N_12830,N_11925);
or U16383 (N_16383,N_12658,N_13237);
and U16384 (N_16384,N_14372,N_13118);
or U16385 (N_16385,N_11312,N_10838);
nor U16386 (N_16386,N_11686,N_14223);
nor U16387 (N_16387,N_12724,N_10495);
and U16388 (N_16388,N_11630,N_14239);
nor U16389 (N_16389,N_13122,N_11277);
xnor U16390 (N_16390,N_13818,N_12121);
and U16391 (N_16391,N_14906,N_14503);
xnor U16392 (N_16392,N_11878,N_13016);
xor U16393 (N_16393,N_11897,N_11626);
or U16394 (N_16394,N_12246,N_10161);
or U16395 (N_16395,N_12038,N_14066);
and U16396 (N_16396,N_14927,N_11182);
or U16397 (N_16397,N_14699,N_12424);
nand U16398 (N_16398,N_14246,N_11298);
and U16399 (N_16399,N_13364,N_10338);
xor U16400 (N_16400,N_10587,N_11319);
or U16401 (N_16401,N_13569,N_10196);
xor U16402 (N_16402,N_14014,N_13227);
or U16403 (N_16403,N_14655,N_13987);
xnor U16404 (N_16404,N_10326,N_10926);
and U16405 (N_16405,N_11456,N_14424);
or U16406 (N_16406,N_11691,N_10690);
xor U16407 (N_16407,N_10945,N_13990);
nor U16408 (N_16408,N_12290,N_12917);
and U16409 (N_16409,N_14313,N_12138);
xor U16410 (N_16410,N_14757,N_13448);
nor U16411 (N_16411,N_14920,N_13335);
nor U16412 (N_16412,N_12818,N_11542);
xnor U16413 (N_16413,N_13751,N_10333);
or U16414 (N_16414,N_14667,N_12049);
nor U16415 (N_16415,N_12349,N_13735);
and U16416 (N_16416,N_11440,N_12518);
and U16417 (N_16417,N_11196,N_11869);
xor U16418 (N_16418,N_13551,N_13923);
nor U16419 (N_16419,N_13166,N_11936);
nor U16420 (N_16420,N_10068,N_10105);
and U16421 (N_16421,N_10433,N_11222);
nor U16422 (N_16422,N_11668,N_14856);
or U16423 (N_16423,N_10124,N_12194);
nor U16424 (N_16424,N_11548,N_10172);
nor U16425 (N_16425,N_11284,N_13561);
nand U16426 (N_16426,N_11646,N_12263);
nand U16427 (N_16427,N_10929,N_12632);
and U16428 (N_16428,N_13552,N_12559);
and U16429 (N_16429,N_10809,N_13119);
nand U16430 (N_16430,N_11906,N_12393);
xor U16431 (N_16431,N_10086,N_11413);
nand U16432 (N_16432,N_12624,N_10361);
or U16433 (N_16433,N_14556,N_14037);
nor U16434 (N_16434,N_10238,N_13780);
nand U16435 (N_16435,N_14693,N_11730);
or U16436 (N_16436,N_13802,N_14295);
and U16437 (N_16437,N_11912,N_14482);
and U16438 (N_16438,N_11790,N_13460);
or U16439 (N_16439,N_14926,N_13442);
nand U16440 (N_16440,N_12972,N_11923);
or U16441 (N_16441,N_14724,N_11838);
nand U16442 (N_16442,N_14073,N_12890);
and U16443 (N_16443,N_13897,N_11587);
xor U16444 (N_16444,N_12114,N_14594);
xnor U16445 (N_16445,N_14919,N_14237);
nand U16446 (N_16446,N_10726,N_11551);
xor U16447 (N_16447,N_13039,N_11462);
nor U16448 (N_16448,N_10094,N_11069);
xor U16449 (N_16449,N_10285,N_12409);
and U16450 (N_16450,N_12174,N_14146);
nor U16451 (N_16451,N_10880,N_10598);
nand U16452 (N_16452,N_13284,N_11300);
xnor U16453 (N_16453,N_10475,N_13643);
or U16454 (N_16454,N_11540,N_13296);
or U16455 (N_16455,N_10469,N_14410);
and U16456 (N_16456,N_11536,N_14282);
or U16457 (N_16457,N_12947,N_13449);
nand U16458 (N_16458,N_10282,N_11681);
and U16459 (N_16459,N_13898,N_12008);
xor U16460 (N_16460,N_13035,N_11431);
nor U16461 (N_16461,N_11565,N_12746);
nor U16462 (N_16462,N_12639,N_10373);
nor U16463 (N_16463,N_10271,N_11511);
xor U16464 (N_16464,N_12735,N_11801);
nand U16465 (N_16465,N_10607,N_12842);
nand U16466 (N_16466,N_14324,N_14338);
xor U16467 (N_16467,N_11092,N_11003);
or U16468 (N_16468,N_14704,N_14886);
or U16469 (N_16469,N_13232,N_13461);
xnor U16470 (N_16470,N_12414,N_10413);
xor U16471 (N_16471,N_13994,N_13650);
nor U16472 (N_16472,N_11967,N_12481);
nand U16473 (N_16473,N_12397,N_14659);
nor U16474 (N_16474,N_10928,N_13475);
nor U16475 (N_16475,N_13429,N_10625);
or U16476 (N_16476,N_10134,N_12966);
xnor U16477 (N_16477,N_10963,N_10675);
nor U16478 (N_16478,N_11844,N_13493);
nor U16479 (N_16479,N_12460,N_11875);
nor U16480 (N_16480,N_14531,N_11648);
nor U16481 (N_16481,N_10865,N_13617);
or U16482 (N_16482,N_10046,N_12637);
xor U16483 (N_16483,N_14745,N_11015);
xor U16484 (N_16484,N_12579,N_12048);
and U16485 (N_16485,N_13100,N_13230);
and U16486 (N_16486,N_13512,N_10787);
xnor U16487 (N_16487,N_13243,N_10131);
and U16488 (N_16488,N_14639,N_14808);
xnor U16489 (N_16489,N_12703,N_12471);
and U16490 (N_16490,N_11160,N_13909);
nand U16491 (N_16491,N_13933,N_14412);
or U16492 (N_16492,N_13207,N_12407);
xor U16493 (N_16493,N_13068,N_14924);
nand U16494 (N_16494,N_11303,N_10958);
nor U16495 (N_16495,N_12339,N_12693);
nor U16496 (N_16496,N_11034,N_11427);
xor U16497 (N_16497,N_12422,N_12994);
nor U16498 (N_16498,N_11488,N_13667);
and U16499 (N_16499,N_14029,N_11873);
nor U16500 (N_16500,N_12244,N_10316);
nor U16501 (N_16501,N_13390,N_14806);
or U16502 (N_16502,N_14098,N_12125);
nand U16503 (N_16503,N_11997,N_12303);
nand U16504 (N_16504,N_12565,N_10909);
xnor U16505 (N_16505,N_10771,N_10432);
nor U16506 (N_16506,N_10359,N_13056);
nor U16507 (N_16507,N_13900,N_12844);
and U16508 (N_16508,N_10657,N_13193);
or U16509 (N_16509,N_10765,N_10256);
or U16510 (N_16510,N_12561,N_14888);
or U16511 (N_16511,N_10183,N_13515);
xor U16512 (N_16512,N_11348,N_14040);
nand U16513 (N_16513,N_11381,N_10182);
or U16514 (N_16514,N_14310,N_13886);
nor U16515 (N_16515,N_10615,N_12846);
xor U16516 (N_16516,N_13786,N_10594);
xnor U16517 (N_16517,N_11152,N_10198);
or U16518 (N_16518,N_13968,N_14932);
nor U16519 (N_16519,N_12101,N_13524);
nand U16520 (N_16520,N_10479,N_12325);
xor U16521 (N_16521,N_11088,N_13758);
or U16522 (N_16522,N_10644,N_14894);
nand U16523 (N_16523,N_14123,N_14817);
nor U16524 (N_16524,N_12752,N_10353);
nand U16525 (N_16525,N_14028,N_12500);
nand U16526 (N_16526,N_10744,N_12755);
nand U16527 (N_16527,N_10876,N_10575);
xor U16528 (N_16528,N_10242,N_12610);
nand U16529 (N_16529,N_13920,N_13979);
and U16530 (N_16530,N_12473,N_10758);
nand U16531 (N_16531,N_12617,N_12220);
nor U16532 (N_16532,N_13682,N_12337);
xnor U16533 (N_16533,N_11532,N_12918);
or U16534 (N_16534,N_13431,N_11913);
or U16535 (N_16535,N_13516,N_10243);
nor U16536 (N_16536,N_14049,N_12302);
nor U16537 (N_16537,N_10930,N_12619);
xnor U16538 (N_16538,N_12911,N_13167);
or U16539 (N_16539,N_11749,N_12980);
or U16540 (N_16540,N_13678,N_12501);
or U16541 (N_16541,N_12079,N_10522);
or U16542 (N_16542,N_13301,N_13816);
nor U16543 (N_16543,N_13769,N_10478);
nand U16544 (N_16544,N_10146,N_10562);
nor U16545 (N_16545,N_14810,N_13125);
or U16546 (N_16546,N_14884,N_12301);
nand U16547 (N_16547,N_13104,N_11385);
nor U16548 (N_16548,N_10602,N_14966);
nand U16549 (N_16549,N_11239,N_13618);
nor U16550 (N_16550,N_12621,N_11892);
xor U16551 (N_16551,N_11879,N_11109);
nor U16552 (N_16552,N_11112,N_11907);
or U16553 (N_16553,N_13005,N_10949);
or U16554 (N_16554,N_11855,N_14854);
or U16555 (N_16555,N_14584,N_14537);
or U16556 (N_16556,N_12229,N_11724);
and U16557 (N_16557,N_10335,N_13128);
nand U16558 (N_16558,N_10147,N_14162);
or U16559 (N_16559,N_11355,N_13825);
or U16560 (N_16560,N_13925,N_11365);
or U16561 (N_16561,N_10818,N_14319);
or U16562 (N_16562,N_11852,N_13345);
or U16563 (N_16563,N_11367,N_10461);
nor U16564 (N_16564,N_13044,N_10310);
nor U16565 (N_16565,N_10166,N_10884);
xor U16566 (N_16566,N_14751,N_12850);
xor U16567 (N_16567,N_13736,N_10717);
and U16568 (N_16568,N_10868,N_11324);
and U16569 (N_16569,N_11734,N_11007);
or U16570 (N_16570,N_13050,N_14598);
and U16571 (N_16571,N_14601,N_10067);
xnor U16572 (N_16572,N_14043,N_12634);
and U16573 (N_16573,N_10966,N_14360);
nor U16574 (N_16574,N_14508,N_13383);
and U16575 (N_16575,N_11516,N_10597);
xnor U16576 (N_16576,N_14878,N_13651);
and U16577 (N_16577,N_14229,N_10516);
or U16578 (N_16578,N_14081,N_14269);
or U16579 (N_16579,N_10269,N_13590);
nand U16580 (N_16580,N_14713,N_10810);
nand U16581 (N_16581,N_10264,N_13588);
nand U16582 (N_16582,N_12169,N_12847);
and U16583 (N_16583,N_10999,N_12938);
nor U16584 (N_16584,N_11443,N_14284);
and U16585 (N_16585,N_11293,N_14538);
xor U16586 (N_16586,N_14222,N_12253);
nand U16587 (N_16587,N_10507,N_10549);
nand U16588 (N_16588,N_10082,N_12836);
and U16589 (N_16589,N_12686,N_13498);
nor U16590 (N_16590,N_12202,N_10900);
nand U16591 (N_16591,N_10781,N_10670);
or U16592 (N_16592,N_10669,N_10294);
and U16593 (N_16593,N_11209,N_10922);
or U16594 (N_16594,N_11001,N_11876);
xor U16595 (N_16595,N_14453,N_14299);
xor U16596 (N_16596,N_12117,N_11031);
and U16597 (N_16597,N_14561,N_11582);
xnor U16598 (N_16598,N_14544,N_11436);
or U16599 (N_16599,N_12796,N_12183);
nand U16600 (N_16600,N_12859,N_12950);
nor U16601 (N_16601,N_13229,N_10191);
and U16602 (N_16602,N_11828,N_14244);
xnor U16603 (N_16603,N_14811,N_11698);
or U16604 (N_16604,N_11442,N_12726);
nor U16605 (N_16605,N_12698,N_12037);
and U16606 (N_16606,N_10619,N_10464);
xnor U16607 (N_16607,N_12313,N_12825);
xnor U16608 (N_16608,N_13147,N_12477);
nor U16609 (N_16609,N_10635,N_13344);
nand U16610 (N_16610,N_12679,N_11991);
and U16611 (N_16611,N_12705,N_10049);
and U16612 (N_16612,N_10154,N_14526);
xnor U16613 (N_16613,N_12029,N_13505);
and U16614 (N_16614,N_13877,N_11418);
xor U16615 (N_16615,N_10971,N_13771);
xnor U16616 (N_16616,N_11318,N_13002);
or U16617 (N_16617,N_12273,N_10341);
xnor U16618 (N_16618,N_13378,N_11212);
nor U16619 (N_16619,N_14399,N_12287);
nand U16620 (N_16620,N_12536,N_11858);
or U16621 (N_16621,N_11050,N_14737);
xor U16622 (N_16622,N_14865,N_11080);
nor U16623 (N_16623,N_12461,N_13811);
xnor U16624 (N_16624,N_12294,N_14719);
nand U16625 (N_16625,N_10577,N_10772);
xor U16626 (N_16626,N_12601,N_14635);
nand U16627 (N_16627,N_10005,N_13540);
and U16628 (N_16628,N_11683,N_13669);
nand U16629 (N_16629,N_14885,N_10417);
nand U16630 (N_16630,N_13142,N_12702);
nand U16631 (N_16631,N_14210,N_11193);
xor U16632 (N_16632,N_10122,N_12071);
or U16633 (N_16633,N_13316,N_12280);
nand U16634 (N_16634,N_11899,N_14250);
and U16635 (N_16635,N_10542,N_12689);
nor U16636 (N_16636,N_11700,N_13196);
and U16637 (N_16637,N_12983,N_14501);
nand U16638 (N_16638,N_13430,N_10552);
xnor U16639 (N_16639,N_12898,N_10910);
xor U16640 (N_16640,N_10386,N_11738);
nor U16641 (N_16641,N_10887,N_10845);
and U16642 (N_16642,N_10696,N_10489);
nand U16643 (N_16643,N_10530,N_12652);
nand U16644 (N_16644,N_11492,N_10297);
nand U16645 (N_16645,N_12945,N_10029);
or U16646 (N_16646,N_12922,N_14763);
xor U16647 (N_16647,N_10100,N_12182);
or U16648 (N_16648,N_13712,N_14506);
nand U16649 (N_16649,N_12100,N_11673);
xnor U16650 (N_16650,N_12913,N_13467);
and U16651 (N_16651,N_10235,N_12413);
nand U16652 (N_16652,N_10321,N_10686);
nand U16653 (N_16653,N_14487,N_14516);
or U16654 (N_16654,N_12763,N_10435);
or U16655 (N_16655,N_14893,N_13638);
nor U16656 (N_16656,N_14722,N_11362);
xor U16657 (N_16657,N_12257,N_10360);
and U16658 (N_16658,N_12987,N_13975);
or U16659 (N_16659,N_13012,N_10492);
xnor U16660 (N_16660,N_10775,N_14554);
xor U16661 (N_16661,N_13279,N_11670);
nand U16662 (N_16662,N_10409,N_10376);
nand U16663 (N_16663,N_12023,N_11157);
and U16664 (N_16664,N_12066,N_13784);
or U16665 (N_16665,N_13814,N_14735);
xnor U16666 (N_16666,N_10548,N_12282);
or U16667 (N_16667,N_12732,N_11554);
nand U16668 (N_16668,N_12683,N_11981);
nor U16669 (N_16669,N_12597,N_13492);
or U16670 (N_16670,N_12576,N_10611);
or U16671 (N_16671,N_12989,N_11732);
nand U16672 (N_16672,N_12675,N_12669);
or U16673 (N_16673,N_12841,N_14725);
nor U16674 (N_16674,N_12022,N_13630);
and U16675 (N_16675,N_14033,N_10692);
nor U16676 (N_16676,N_13276,N_10907);
nand U16677 (N_16677,N_12665,N_13997);
or U16678 (N_16678,N_11077,N_10631);
and U16679 (N_16679,N_10851,N_13918);
xor U16680 (N_16680,N_13143,N_12867);
nand U16681 (N_16681,N_13148,N_14605);
or U16682 (N_16682,N_13258,N_14991);
and U16683 (N_16683,N_10988,N_14541);
nand U16684 (N_16684,N_13833,N_11860);
xor U16685 (N_16685,N_10289,N_12251);
xnor U16686 (N_16686,N_13205,N_14933);
or U16687 (N_16687,N_14171,N_14401);
xor U16688 (N_16688,N_11441,N_14447);
nor U16689 (N_16689,N_10123,N_13307);
and U16690 (N_16690,N_11377,N_10457);
or U16691 (N_16691,N_14072,N_13513);
or U16692 (N_16692,N_12351,N_11256);
nor U16693 (N_16693,N_14666,N_14249);
nor U16694 (N_16694,N_12144,N_10103);
nor U16695 (N_16695,N_12995,N_11290);
nor U16696 (N_16696,N_10952,N_10712);
or U16697 (N_16697,N_14957,N_10576);
nand U16698 (N_16698,N_14527,N_14578);
and U16699 (N_16699,N_14010,N_12061);
and U16700 (N_16700,N_14911,N_13251);
nand U16701 (N_16701,N_11019,N_10959);
nor U16702 (N_16702,N_13346,N_12933);
nor U16703 (N_16703,N_14726,N_13789);
or U16704 (N_16704,N_14940,N_12064);
and U16705 (N_16705,N_12892,N_11745);
xor U16706 (N_16706,N_10474,N_13133);
xor U16707 (N_16707,N_10389,N_11563);
and U16708 (N_16708,N_10975,N_13792);
and U16709 (N_16709,N_10447,N_13655);
nand U16710 (N_16710,N_12311,N_14336);
nand U16711 (N_16711,N_11110,N_11191);
nor U16712 (N_16712,N_13275,N_12221);
xor U16713 (N_16713,N_11690,N_10309);
nor U16714 (N_16714,N_14055,N_13288);
nand U16715 (N_16715,N_12428,N_11555);
xor U16716 (N_16716,N_13901,N_12478);
and U16717 (N_16717,N_11199,N_12284);
and U16718 (N_16718,N_14339,N_12618);
or U16719 (N_16719,N_12907,N_10580);
nor U16720 (N_16720,N_11634,N_10405);
nand U16721 (N_16721,N_14026,N_12655);
xor U16722 (N_16722,N_14963,N_13102);
nor U16723 (N_16723,N_12682,N_14490);
nand U16724 (N_16724,N_11836,N_10915);
or U16725 (N_16725,N_11295,N_10420);
xor U16726 (N_16726,N_12009,N_13986);
nand U16727 (N_16727,N_10225,N_14917);
and U16728 (N_16728,N_14930,N_14580);
nand U16729 (N_16729,N_14176,N_12896);
nand U16730 (N_16730,N_13980,N_12531);
or U16731 (N_16731,N_11244,N_13022);
and U16732 (N_16732,N_13887,N_13126);
nand U16733 (N_16733,N_14024,N_14705);
nor U16734 (N_16734,N_10633,N_14524);
xnor U16735 (N_16735,N_12004,N_11216);
nor U16736 (N_16736,N_13195,N_14852);
nor U16737 (N_16737,N_12611,N_13124);
or U16738 (N_16738,N_13085,N_14264);
or U16739 (N_16739,N_14027,N_11975);
and U16740 (N_16740,N_11491,N_11868);
and U16741 (N_16741,N_10480,N_13904);
and U16742 (N_16742,N_10745,N_14530);
or U16743 (N_16743,N_13665,N_10600);
nor U16744 (N_16744,N_11446,N_14292);
or U16745 (N_16745,N_12544,N_12930);
nor U16746 (N_16746,N_14391,N_14644);
nor U16747 (N_16747,N_14743,N_13579);
and U16748 (N_16748,N_11994,N_10976);
and U16749 (N_16749,N_12002,N_10850);
xor U16750 (N_16750,N_10601,N_14621);
xor U16751 (N_16751,N_11874,N_10933);
and U16752 (N_16752,N_11271,N_14243);
xor U16753 (N_16753,N_14106,N_13970);
nor U16754 (N_16754,N_13270,N_14761);
nor U16755 (N_16755,N_12878,N_11669);
xnor U16756 (N_16756,N_11307,N_11267);
and U16757 (N_16757,N_12479,N_11326);
or U16758 (N_16758,N_14799,N_13290);
xnor U16759 (N_16759,N_14775,N_14841);
or U16760 (N_16760,N_10193,N_10098);
and U16761 (N_16761,N_11045,N_10329);
nor U16762 (N_16762,N_11862,N_13157);
xnor U16763 (N_16763,N_11111,N_13782);
xnor U16764 (N_16764,N_12516,N_10412);
xor U16765 (N_16765,N_12543,N_12411);
nand U16766 (N_16766,N_11214,N_11703);
or U16767 (N_16767,N_13259,N_11366);
nand U16768 (N_16768,N_14954,N_12960);
and U16769 (N_16769,N_13804,N_14896);
and U16770 (N_16770,N_10993,N_12853);
nand U16771 (N_16771,N_14603,N_12466);
nand U16772 (N_16772,N_14144,N_13760);
nor U16773 (N_16773,N_10222,N_11896);
or U16774 (N_16774,N_10069,N_14515);
nand U16775 (N_16775,N_14630,N_12328);
xor U16776 (N_16776,N_13420,N_14784);
or U16777 (N_16777,N_12156,N_11338);
nand U16778 (N_16778,N_14371,N_12131);
nand U16779 (N_16779,N_14265,N_13929);
nand U16780 (N_16780,N_13073,N_13217);
nand U16781 (N_16781,N_10113,N_14707);
xor U16782 (N_16782,N_10127,N_13625);
or U16783 (N_16783,N_11257,N_11482);
nor U16784 (N_16784,N_14382,N_14574);
nand U16785 (N_16785,N_13964,N_11188);
xor U16786 (N_16786,N_12110,N_12738);
and U16787 (N_16787,N_12467,N_12562);
and U16788 (N_16788,N_14159,N_12777);
nor U16789 (N_16789,N_11512,N_13855);
nor U16790 (N_16790,N_12840,N_14369);
nand U16791 (N_16791,N_12259,N_14349);
nor U16792 (N_16792,N_11315,N_13984);
nor U16793 (N_16793,N_14701,N_13907);
xnor U16794 (N_16794,N_14441,N_12394);
and U16795 (N_16795,N_13889,N_11287);
xnor U16796 (N_16796,N_10642,N_14203);
nor U16797 (N_16797,N_13029,N_12712);
xnor U16798 (N_16798,N_11073,N_12067);
nor U16799 (N_16799,N_10624,N_14868);
nor U16800 (N_16800,N_11977,N_11329);
nand U16801 (N_16801,N_13292,N_10916);
or U16802 (N_16802,N_11569,N_10519);
and U16803 (N_16803,N_12526,N_10776);
nand U16804 (N_16804,N_14695,N_12310);
and U16805 (N_16805,N_14864,N_12615);
nor U16806 (N_16806,N_11792,N_14853);
nand U16807 (N_16807,N_13834,N_13750);
or U16808 (N_16808,N_10847,N_11085);
xor U16809 (N_16809,N_11200,N_12955);
nand U16810 (N_16810,N_10506,N_13107);
nand U16811 (N_16811,N_10384,N_12175);
and U16812 (N_16812,N_11884,N_14357);
nand U16813 (N_16813,N_12833,N_13014);
nand U16814 (N_16814,N_12326,N_14960);
xnor U16815 (N_16815,N_14566,N_11124);
and U16816 (N_16816,N_10965,N_14099);
nor U16817 (N_16817,N_13748,N_11032);
and U16818 (N_16818,N_11697,N_14136);
or U16819 (N_16819,N_14718,N_14871);
nand U16820 (N_16820,N_12946,N_13719);
and U16821 (N_16821,N_12436,N_14778);
nor U16822 (N_16822,N_13824,N_14325);
and U16823 (N_16823,N_10442,N_12783);
nand U16824 (N_16824,N_13271,N_13694);
and U16825 (N_16825,N_14948,N_12084);
nor U16826 (N_16826,N_12205,N_13976);
or U16827 (N_16827,N_10418,N_14396);
or U16828 (N_16828,N_14440,N_13581);
nor U16829 (N_16829,N_13169,N_12198);
and U16830 (N_16830,N_11619,N_10623);
or U16831 (N_16831,N_10582,N_10167);
nor U16832 (N_16832,N_11231,N_14105);
nor U16833 (N_16833,N_11429,N_12447);
or U16834 (N_16834,N_10458,N_13397);
nor U16835 (N_16835,N_13093,N_13380);
or U16836 (N_16836,N_10532,N_10960);
nand U16837 (N_16837,N_11500,N_13995);
nor U16838 (N_16838,N_11087,N_14790);
xnor U16839 (N_16839,N_13112,N_12677);
and U16840 (N_16840,N_10779,N_14575);
and U16841 (N_16841,N_10139,N_11393);
nand U16842 (N_16842,N_12523,N_11333);
and U16843 (N_16843,N_13076,N_10429);
and U16844 (N_16844,N_10187,N_13186);
nand U16845 (N_16845,N_10274,N_11661);
or U16846 (N_16846,N_11659,N_12593);
nand U16847 (N_16847,N_10482,N_13967);
xor U16848 (N_16848,N_12168,N_14116);
nand U16849 (N_16849,N_13620,N_13911);
or U16850 (N_16850,N_11422,N_14126);
nand U16851 (N_16851,N_10676,N_11426);
or U16852 (N_16852,N_10987,N_10768);
xor U16853 (N_16853,N_10857,N_11595);
nor U16854 (N_16854,N_11972,N_11866);
xnor U16855 (N_16855,N_12132,N_14857);
nand U16856 (N_16856,N_11474,N_13248);
or U16857 (N_16857,N_11411,N_12300);
or U16858 (N_16858,N_14221,N_13359);
and U16859 (N_16859,N_12377,N_13000);
nor U16860 (N_16860,N_10806,N_12115);
nor U16861 (N_16861,N_13859,N_12714);
nand U16862 (N_16862,N_14714,N_13334);
and U16863 (N_16863,N_12086,N_13462);
xor U16864 (N_16864,N_11819,N_11597);
nor U16865 (N_16865,N_10671,N_13953);
and U16866 (N_16866,N_12759,N_10199);
xor U16867 (N_16867,N_12574,N_12874);
nand U16868 (N_16868,N_14617,N_13594);
nor U16869 (N_16869,N_11176,N_13170);
xnor U16870 (N_16870,N_10736,N_11170);
nor U16871 (N_16871,N_13393,N_10888);
nand U16872 (N_16872,N_12118,N_12927);
and U16873 (N_16873,N_14427,N_11917);
xor U16874 (N_16874,N_11433,N_11910);
nor U16875 (N_16875,N_13326,N_14624);
nor U16876 (N_16876,N_14419,N_14430);
or U16877 (N_16877,N_13922,N_11408);
nor U16878 (N_16878,N_11455,N_10528);
or U16879 (N_16879,N_14163,N_13885);
nor U16880 (N_16880,N_14416,N_13616);
or U16881 (N_16881,N_11880,N_13149);
xor U16882 (N_16882,N_13194,N_10431);
nand U16883 (N_16883,N_13892,N_11184);
xnor U16884 (N_16884,N_10830,N_12532);
xor U16885 (N_16885,N_14949,N_10531);
nor U16886 (N_16886,N_13675,N_12509);
nor U16887 (N_16887,N_10760,N_12970);
xor U16888 (N_16888,N_10244,N_13451);
or U16889 (N_16889,N_12659,N_12025);
xor U16890 (N_16890,N_13840,N_12717);
nand U16891 (N_16891,N_12809,N_14869);
and U16892 (N_16892,N_14535,N_12954);
nand U16893 (N_16893,N_11731,N_10307);
and U16894 (N_16894,N_13705,N_14652);
or U16895 (N_16895,N_14680,N_12753);
nor U16896 (N_16896,N_14361,N_12275);
nor U16897 (N_16897,N_10034,N_10093);
or U16898 (N_16898,N_12155,N_11420);
or U16899 (N_16899,N_13770,N_10121);
nor U16900 (N_16900,N_11929,N_10313);
nor U16901 (N_16901,N_14312,N_10719);
xor U16902 (N_16902,N_14193,N_13807);
or U16903 (N_16903,N_11579,N_14684);
and U16904 (N_16904,N_12662,N_10751);
nor U16905 (N_16905,N_10339,N_14764);
nand U16906 (N_16906,N_10315,N_13881);
nand U16907 (N_16907,N_11264,N_12996);
and U16908 (N_16908,N_11187,N_11395);
nor U16909 (N_16909,N_13220,N_10529);
xnor U16910 (N_16910,N_13053,N_13018);
and U16911 (N_16911,N_13683,N_11685);
and U16912 (N_16912,N_10056,N_13105);
nor U16913 (N_16913,N_14898,N_12451);
xor U16914 (N_16914,N_13985,N_12828);
or U16915 (N_16915,N_14076,N_14913);
xor U16916 (N_16916,N_13021,N_10048);
nand U16917 (N_16917,N_14573,N_13738);
nand U16918 (N_16918,N_14444,N_12489);
or U16919 (N_16919,N_11524,N_14647);
nor U16920 (N_16920,N_13382,N_11713);
xor U16921 (N_16921,N_11606,N_11384);
and U16922 (N_16922,N_10734,N_12215);
nor U16923 (N_16923,N_13589,N_12226);
nand U16924 (N_16924,N_11041,N_10918);
xor U16925 (N_16925,N_12910,N_13921);
xor U16926 (N_16926,N_11987,N_10875);
and U16927 (N_16927,N_14990,N_13109);
nor U16928 (N_16928,N_11864,N_12134);
or U16929 (N_16929,N_11709,N_12254);
nand U16930 (N_16930,N_13080,N_12030);
or U16931 (N_16931,N_14553,N_12616);
and U16932 (N_16932,N_11610,N_11940);
xnor U16933 (N_16933,N_13374,N_13862);
or U16934 (N_16934,N_13273,N_10406);
and U16935 (N_16935,N_11204,N_11853);
and U16936 (N_16936,N_11136,N_13992);
nor U16937 (N_16937,N_11452,N_12092);
nor U16938 (N_16938,N_11946,N_11025);
xnor U16939 (N_16939,N_13635,N_14814);
and U16940 (N_16940,N_14017,N_11238);
nand U16941 (N_16941,N_13910,N_13938);
xnor U16942 (N_16942,N_14555,N_13240);
xor U16943 (N_16943,N_14688,N_14867);
or U16944 (N_16944,N_13067,N_10684);
xnor U16945 (N_16945,N_12901,N_13959);
nand U16946 (N_16946,N_13372,N_14248);
xor U16947 (N_16947,N_10334,N_11560);
and U16948 (N_16948,N_13715,N_13001);
and U16949 (N_16949,N_10063,N_14294);
xor U16950 (N_16950,N_11040,N_12232);
xnor U16951 (N_16951,N_12780,N_13514);
nand U16952 (N_16952,N_10270,N_10021);
xnor U16953 (N_16953,N_14007,N_10163);
xor U16954 (N_16954,N_13184,N_10974);
or U16955 (N_16955,N_13008,N_13421);
nor U16956 (N_16956,N_14232,N_12627);
and U16957 (N_16957,N_12141,N_10581);
nor U16958 (N_16958,N_11489,N_10709);
nand U16959 (N_16959,N_10047,N_13312);
nand U16960 (N_16960,N_14660,N_14344);
or U16961 (N_16961,N_12161,N_13545);
and U16962 (N_16962,N_14042,N_11914);
and U16963 (N_16963,N_12784,N_10596);
nand U16964 (N_16964,N_12906,N_10117);
nor U16965 (N_16965,N_10251,N_12919);
nor U16966 (N_16966,N_10101,N_11178);
and U16967 (N_16967,N_11616,N_11270);
nand U16968 (N_16968,N_11093,N_12392);
xnor U16969 (N_16969,N_10241,N_11861);
or U16970 (N_16970,N_13890,N_11671);
nor U16971 (N_16971,N_11129,N_12915);
xor U16972 (N_16972,N_13848,N_12382);
nor U16973 (N_16973,N_11574,N_14589);
and U16974 (N_16974,N_10701,N_14822);
nand U16975 (N_16975,N_13955,N_14681);
xnor U16976 (N_16976,N_10950,N_11904);
nand U16977 (N_16977,N_11439,N_14197);
or U16978 (N_16978,N_11680,N_10414);
and U16979 (N_16979,N_14591,N_13856);
xor U16980 (N_16980,N_11459,N_11051);
and U16981 (N_16981,N_14152,N_13688);
xnor U16982 (N_16982,N_10092,N_13464);
nand U16983 (N_16983,N_14224,N_14075);
nand U16984 (N_16984,N_11558,N_10740);
and U16985 (N_16985,N_14844,N_12827);
nand U16986 (N_16986,N_12595,N_11748);
xnor U16987 (N_16987,N_11038,N_10766);
xor U16988 (N_16988,N_14509,N_13485);
nor U16989 (N_16989,N_10153,N_11927);
nand U16990 (N_16990,N_11252,N_13447);
or U16991 (N_16991,N_12116,N_13487);
nand U16992 (N_16992,N_14492,N_11352);
or U16993 (N_16993,N_11304,N_12598);
xor U16994 (N_16994,N_11229,N_11499);
or U16995 (N_16995,N_13697,N_12694);
and U16996 (N_16996,N_10984,N_10448);
xnor U16997 (N_16997,N_12834,N_12581);
xor U16998 (N_16998,N_14807,N_14102);
and U16999 (N_16999,N_12320,N_11575);
xor U17000 (N_17000,N_11672,N_14646);
nand U17001 (N_17001,N_11950,N_14463);
and U17002 (N_17002,N_11071,N_10453);
xor U17003 (N_17003,N_14343,N_14057);
or U17004 (N_17004,N_10091,N_14177);
nand U17005 (N_17005,N_11128,N_10885);
nor U17006 (N_17006,N_14406,N_11781);
or U17007 (N_17007,N_14986,N_12742);
or U17008 (N_17008,N_10279,N_13570);
xor U17009 (N_17009,N_13300,N_14910);
or U17010 (N_17010,N_12707,N_10526);
nand U17011 (N_17011,N_10035,N_13679);
xor U17012 (N_17012,N_11108,N_14356);
or U17013 (N_17013,N_13778,N_14676);
xor U17014 (N_17014,N_10102,N_11094);
nor U17015 (N_17015,N_12891,N_12268);
or U17016 (N_17016,N_10249,N_10539);
nor U17017 (N_17017,N_11623,N_10356);
xor U17018 (N_17018,N_12573,N_13198);
nor U17019 (N_17019,N_13331,N_13078);
nor U17020 (N_17020,N_10593,N_14678);
xnor U17021 (N_17021,N_12572,N_12696);
and U17022 (N_17022,N_13419,N_11832);
or U17023 (N_17023,N_13256,N_10979);
xnor U17024 (N_17024,N_10399,N_13725);
or U17025 (N_17025,N_10213,N_13437);
xor U17026 (N_17026,N_11823,N_13079);
nor U17027 (N_17027,N_12902,N_11916);
xor U17028 (N_17028,N_13690,N_10236);
xor U17029 (N_17029,N_13685,N_10588);
or U17030 (N_17030,N_11689,N_12053);
and U17031 (N_17031,N_14532,N_14983);
and U17032 (N_17032,N_13846,N_10938);
nor U17033 (N_17033,N_11332,N_13565);
and U17034 (N_17034,N_10258,N_13796);
and U17035 (N_17035,N_12956,N_11886);
xnor U17036 (N_17036,N_13239,N_10967);
nor U17037 (N_17037,N_12599,N_13543);
nor U17038 (N_17038,N_14883,N_14347);
or U17039 (N_17039,N_10688,N_12189);
xnor U17040 (N_17040,N_10566,N_14783);
nand U17041 (N_17041,N_12474,N_11928);
and U17042 (N_17042,N_11699,N_11345);
and U17043 (N_17043,N_13872,N_11100);
nor U17044 (N_17044,N_10148,N_11602);
or U17045 (N_17045,N_10195,N_11043);
nor U17046 (N_17046,N_12210,N_13866);
or U17047 (N_17047,N_13272,N_11052);
or U17048 (N_17048,N_12934,N_12592);
nor U17049 (N_17049,N_11818,N_10368);
and U17050 (N_17050,N_10660,N_10956);
nor U17051 (N_17051,N_12113,N_11350);
xnor U17052 (N_17052,N_10626,N_12065);
or U17053 (N_17053,N_12201,N_11437);
xnor U17054 (N_17054,N_13883,N_11151);
xnor U17055 (N_17055,N_11757,N_11360);
nor U17056 (N_17056,N_13013,N_12185);
xor U17057 (N_17057,N_12146,N_12077);
nor U17058 (N_17058,N_11590,N_13098);
nand U17059 (N_17059,N_13350,N_11354);
or U17060 (N_17060,N_12643,N_14058);
nor U17061 (N_17061,N_13181,N_10206);
nand U17062 (N_17062,N_12233,N_11771);
xor U17063 (N_17063,N_13228,N_13839);
xor U17064 (N_17064,N_12612,N_13422);
xnor U17065 (N_17065,N_10937,N_10379);
or U17066 (N_17066,N_12350,N_14734);
and U17067 (N_17067,N_11549,N_10494);
nor U17068 (N_17068,N_12745,N_14766);
and U17069 (N_17069,N_12391,N_10788);
or U17070 (N_17070,N_12372,N_10534);
nand U17071 (N_17071,N_12395,N_14846);
nor U17072 (N_17072,N_11658,N_14442);
and U17073 (N_17073,N_14121,N_11624);
nor U17074 (N_17074,N_12018,N_13496);
or U17075 (N_17075,N_12288,N_12704);
xor U17076 (N_17076,N_10860,N_12997);
xor U17077 (N_17077,N_11758,N_14212);
nor U17078 (N_17078,N_13436,N_14411);
nor U17079 (N_17079,N_12060,N_11299);
or U17080 (N_17080,N_11247,N_10443);
nand U17081 (N_17081,N_11266,N_11313);
nand U17082 (N_17082,N_11736,N_14079);
xnor U17083 (N_17083,N_13176,N_14984);
nand U17084 (N_17084,N_13517,N_10970);
xor U17085 (N_17085,N_11552,N_14201);
and U17086 (N_17086,N_10757,N_14464);
or U17087 (N_17087,N_11059,N_12028);
and U17088 (N_17088,N_10207,N_10286);
and U17089 (N_17089,N_13218,N_11296);
and U17090 (N_17090,N_10617,N_11772);
or U17091 (N_17091,N_13336,N_14107);
or U17092 (N_17092,N_13550,N_13982);
xor U17093 (N_17093,N_11219,N_10498);
or U17094 (N_17094,N_10881,N_10212);
xnor U17095 (N_17095,N_14362,N_11909);
nor U17096 (N_17096,N_11135,N_12285);
nor U17097 (N_17097,N_13450,N_13766);
or U17098 (N_17098,N_13863,N_14483);
or U17099 (N_17099,N_13410,N_12024);
and U17100 (N_17100,N_11375,N_14225);
and U17101 (N_17101,N_12835,N_14942);
and U17102 (N_17102,N_14161,N_12332);
and U17103 (N_17103,N_11539,N_10533);
or U17104 (N_17104,N_14781,N_11715);
xnor U17105 (N_17105,N_11924,N_12357);
xnor U17106 (N_17106,N_12533,N_13873);
or U17107 (N_17107,N_14143,N_11062);
nand U17108 (N_17108,N_10753,N_10428);
xnor U17109 (N_17109,N_12813,N_10652);
and U17110 (N_17110,N_14215,N_11079);
xnor U17111 (N_17111,N_11842,N_14266);
and U17112 (N_17112,N_12039,N_12074);
xor U17113 (N_17113,N_13038,N_11614);
and U17114 (N_17114,N_12628,N_14012);
nand U17115 (N_17115,N_14062,N_14762);
or U17116 (N_17116,N_12604,N_14196);
and U17117 (N_17117,N_14459,N_11101);
nor U17118 (N_17118,N_11475,N_12528);
nand U17119 (N_17119,N_14543,N_10039);
nand U17120 (N_17120,N_14323,N_11502);
and U17121 (N_17121,N_11220,N_12319);
nor U17122 (N_17122,N_13108,N_12494);
xor U17123 (N_17123,N_12348,N_12454);
nand U17124 (N_17124,N_13330,N_12410);
or U17125 (N_17125,N_12582,N_13684);
nand U17126 (N_17126,N_11049,N_13574);
and U17127 (N_17127,N_14287,N_12358);
or U17128 (N_17128,N_14337,N_10292);
xor U17129 (N_17129,N_14967,N_11227);
nor U17130 (N_17130,N_13793,N_13026);
and U17131 (N_17131,N_13339,N_13132);
and U17132 (N_17132,N_12608,N_13592);
or U17133 (N_17133,N_13939,N_10261);
nand U17134 (N_17134,N_14083,N_13584);
xnor U17135 (N_17135,N_14486,N_10284);
nor U17136 (N_17136,N_11236,N_12711);
or U17137 (N_17137,N_10205,N_13861);
nor U17138 (N_17138,N_14925,N_13254);
nor U17139 (N_17139,N_12982,N_12396);
and U17140 (N_17140,N_14943,N_12191);
or U17141 (N_17141,N_11485,N_14818);
xor U17142 (N_17142,N_11867,N_10890);
xnor U17143 (N_17143,N_13161,N_12239);
xor U17144 (N_17144,N_10622,N_10262);
nor U17145 (N_17145,N_13223,N_12309);
or U17146 (N_17146,N_14115,N_10267);
nor U17147 (N_17147,N_11573,N_11639);
and U17148 (N_17148,N_12779,N_10016);
nor U17149 (N_17149,N_10404,N_11294);
and U17150 (N_17150,N_12260,N_10741);
nand U17151 (N_17151,N_11357,N_13888);
nand U17152 (N_17152,N_14631,N_12327);
or U17153 (N_17153,N_14271,N_11189);
and U17154 (N_17154,N_11114,N_11635);
and U17155 (N_17155,N_12278,N_12685);
nor U17156 (N_17156,N_10216,N_13387);
nand U17157 (N_17157,N_14744,N_10998);
nor U17158 (N_17158,N_11918,N_10394);
and U17159 (N_17159,N_14622,N_14094);
xnor U17160 (N_17160,N_11586,N_12375);
nor U17161 (N_17161,N_10572,N_14478);
xnor U17162 (N_17162,N_11337,N_10411);
nand U17163 (N_17163,N_13621,N_14379);
and U17164 (N_17164,N_12681,N_10869);
and U17165 (N_17165,N_13263,N_13452);
or U17166 (N_17166,N_13775,N_12353);
or U17167 (N_17167,N_10874,N_11258);
and U17168 (N_17168,N_14169,N_13394);
nor U17169 (N_17169,N_14351,N_11172);
xnor U17170 (N_17170,N_11084,N_13828);
nand U17171 (N_17171,N_12051,N_12258);
nor U17172 (N_17172,N_11328,N_13598);
and U17173 (N_17173,N_12097,N_11546);
nand U17174 (N_17174,N_12653,N_14798);
xor U17175 (N_17175,N_11280,N_13580);
or U17176 (N_17176,N_11566,N_11622);
or U17177 (N_17177,N_13249,N_13356);
and U17178 (N_17178,N_12903,N_14368);
xnor U17179 (N_17179,N_10449,N_13293);
nand U17180 (N_17180,N_11127,N_11382);
nor U17181 (N_17181,N_12180,N_13687);
xnor U17182 (N_17182,N_13291,N_14708);
nand U17183 (N_17183,N_13327,N_14247);
or U17184 (N_17184,N_14602,N_12737);
or U17185 (N_17185,N_12209,N_13289);
nand U17186 (N_17186,N_14880,N_14982);
or U17187 (N_17187,N_13140,N_13645);
nand U17188 (N_17188,N_12013,N_14155);
nand U17189 (N_17189,N_11526,N_13400);
or U17190 (N_17190,N_14950,N_10618);
xor U17191 (N_17191,N_12727,N_12733);
and U17192 (N_17192,N_11344,N_10493);
and U17193 (N_17193,N_10465,N_13308);
and U17194 (N_17194,N_10383,N_14308);
nand U17195 (N_17195,N_12799,N_10983);
xor U17196 (N_17196,N_12364,N_14165);
and U17197 (N_17197,N_12153,N_11063);
nor U17198 (N_17198,N_14958,N_10700);
and U17199 (N_17199,N_12108,N_10476);
nand U17200 (N_17200,N_10774,N_12495);
xnor U17201 (N_17201,N_12542,N_10255);
nor U17202 (N_17202,N_12181,N_13313);
nor U17203 (N_17203,N_10621,N_12764);
and U17204 (N_17204,N_14460,N_13025);
xor U17205 (N_17205,N_13626,N_12052);
and U17206 (N_17206,N_10554,N_14662);
nor U17207 (N_17207,N_10077,N_14125);
or U17208 (N_17208,N_13087,N_13226);
nor U17209 (N_17209,N_14825,N_12227);
xnor U17210 (N_17210,N_13368,N_13404);
and U17211 (N_17211,N_14787,N_14826);
xnor U17212 (N_17212,N_11525,N_13003);
xor U17213 (N_17213,N_14838,N_13089);
and U17214 (N_17214,N_10895,N_14242);
and U17215 (N_17215,N_11281,N_12203);
and U17216 (N_17216,N_11729,N_12293);
nand U17217 (N_17217,N_10382,N_10791);
nor U17218 (N_17218,N_10314,N_12865);
and U17219 (N_17219,N_10555,N_12344);
nand U17220 (N_17220,N_14065,N_10296);
xor U17221 (N_17221,N_10129,N_13381);
and U17222 (N_17222,N_13096,N_10277);
or U17223 (N_17223,N_12893,N_11714);
or U17224 (N_17224,N_10550,N_11996);
and U17225 (N_17225,N_10911,N_13407);
xor U17226 (N_17226,N_11316,N_14021);
xor U17227 (N_17227,N_13755,N_12026);
nand U17228 (N_17228,N_11230,N_13538);
nor U17229 (N_17229,N_13596,N_12184);
nor U17230 (N_17230,N_13351,N_13180);
xor U17231 (N_17231,N_14793,N_11235);
nand U17232 (N_17232,N_11342,N_13676);
xor U17233 (N_17233,N_11215,N_12781);
or U17234 (N_17234,N_14423,N_12860);
xnor U17235 (N_17235,N_11414,N_13443);
nand U17236 (N_17236,N_11186,N_11756);
nand U17237 (N_17237,N_12502,N_11805);
and U17238 (N_17238,N_14528,N_14641);
xnor U17239 (N_17239,N_13799,N_13470);
nand U17240 (N_17240,N_10541,N_10638);
nand U17241 (N_17241,N_10925,N_10108);
xor U17242 (N_17242,N_11274,N_13572);
and U17243 (N_17243,N_11720,N_14032);
nand U17244 (N_17244,N_14609,N_13168);
nor U17245 (N_17245,N_13329,N_12520);
or U17246 (N_17246,N_12147,N_11785);
xnor U17247 (N_17247,N_14137,N_12342);
nand U17248 (N_17248,N_12848,N_13849);
and U17249 (N_17249,N_10436,N_11167);
nand U17250 (N_17250,N_10730,N_10819);
nand U17251 (N_17251,N_10204,N_10280);
nand U17252 (N_17252,N_13595,N_13623);
xor U17253 (N_17253,N_12695,N_10483);
nor U17254 (N_17254,N_12880,N_13800);
nor U17255 (N_17255,N_11954,N_14233);
and U17256 (N_17256,N_12638,N_14341);
nand U17257 (N_17257,N_13827,N_13753);
or U17258 (N_17258,N_11998,N_12187);
nor U17259 (N_17259,N_12566,N_11058);
nor U17260 (N_17260,N_10400,N_12664);
xnor U17261 (N_17261,N_13508,N_11849);
or U17262 (N_17262,N_13668,N_10523);
nor U17263 (N_17263,N_13717,N_10331);
and U17264 (N_17264,N_11980,N_12491);
and U17265 (N_17265,N_13479,N_12033);
nand U17266 (N_17266,N_11037,N_14625);
nand U17267 (N_17267,N_10704,N_11473);
nand U17268 (N_17268,N_12370,N_11083);
and U17269 (N_17269,N_11432,N_13260);
or U17270 (N_17270,N_11029,N_10839);
xnor U17271 (N_17271,N_14815,N_10796);
and U17272 (N_17272,N_12484,N_10650);
nand U17273 (N_17273,N_14332,N_14570);
and U17274 (N_17274,N_10502,N_13509);
or U17275 (N_17275,N_14518,N_10904);
and U17276 (N_17276,N_11314,N_14254);
xor U17277 (N_17277,N_12863,N_11960);
xnor U17278 (N_17278,N_11372,N_13153);
or U17279 (N_17279,N_12762,N_10637);
nand U17280 (N_17280,N_12676,N_13895);
and U17281 (N_17281,N_13103,N_13136);
and U17282 (N_17282,N_12583,N_10858);
nor U17283 (N_17283,N_10087,N_11765);
or U17284 (N_17284,N_13152,N_12811);
nand U17285 (N_17285,N_13439,N_13567);
nor U17286 (N_17286,N_11028,N_13500);
nor U17287 (N_17287,N_14170,N_11895);
or U17288 (N_17288,N_13720,N_13399);
and U17289 (N_17289,N_13605,N_10080);
or U17290 (N_17290,N_10902,N_13304);
nand U17291 (N_17291,N_13151,N_14697);
nor U17292 (N_17292,N_14052,N_13701);
nor U17293 (N_17293,N_14944,N_10821);
nand U17294 (N_17294,N_11435,N_10896);
or U17295 (N_17295,N_10060,N_10070);
or U17296 (N_17296,N_13823,N_10538);
nor U17297 (N_17297,N_10535,N_12990);
or U17298 (N_17298,N_13480,N_11317);
xor U17299 (N_17299,N_12506,N_13241);
nand U17300 (N_17300,N_11550,N_12250);
and U17301 (N_17301,N_14842,N_12770);
and U17302 (N_17302,N_11305,N_11652);
and U17303 (N_17303,N_12237,N_11105);
or U17304 (N_17304,N_11451,N_10645);
or U17305 (N_17305,N_14213,N_10151);
xnor U17306 (N_17306,N_12442,N_14740);
xnor U17307 (N_17307,N_12537,N_12510);
nand U17308 (N_17308,N_13732,N_12690);
nand U17309 (N_17309,N_10780,N_11782);
and U17310 (N_17310,N_11121,N_13441);
or U17311 (N_17311,N_14129,N_12126);
or U17312 (N_17312,N_13664,N_14753);
and U17313 (N_17313,N_13936,N_11416);
nand U17314 (N_17314,N_14059,N_13446);
nor U17315 (N_17315,N_10841,N_14972);
xor U17316 (N_17316,N_14650,N_11261);
nand U17317 (N_17317,N_12031,N_13004);
or U17318 (N_17318,N_12856,N_13522);
xnor U17319 (N_17319,N_10231,N_14614);
nor U17320 (N_17320,N_12192,N_14847);
and U17321 (N_17321,N_13077,N_10969);
and U17322 (N_17322,N_10114,N_13940);
xor U17323 (N_17323,N_12058,N_14980);
or U17324 (N_17324,N_11820,N_12864);
nand U17325 (N_17325,N_11175,N_13821);
and U17326 (N_17326,N_11808,N_12151);
or U17327 (N_17327,N_14752,N_10919);
xor U17328 (N_17328,N_13836,N_11496);
and U17329 (N_17329,N_10716,N_10388);
nor U17330 (N_17330,N_10877,N_14030);
and U17331 (N_17331,N_11743,N_11535);
or U17332 (N_17332,N_13191,N_10013);
xnor U17333 (N_17333,N_14458,N_13444);
and U17334 (N_17334,N_14207,N_13323);
nand U17335 (N_17335,N_12527,N_12605);
nand U17336 (N_17336,N_10248,N_10234);
and U17337 (N_17337,N_11742,N_10609);
xnor U17338 (N_17338,N_14002,N_10792);
and U17339 (N_17339,N_14383,N_12314);
nor U17340 (N_17340,N_10419,N_11721);
or U17341 (N_17341,N_13739,N_12207);
nand U17342 (N_17342,N_13774,N_13710);
nand U17343 (N_17343,N_13996,N_11970);
xnor U17344 (N_17344,N_11527,N_14511);
nor U17345 (N_17345,N_13458,N_13173);
nor U17346 (N_17346,N_13745,N_12480);
xor U17347 (N_17347,N_11444,N_11633);
and U17348 (N_17348,N_11224,N_11978);
and U17349 (N_17349,N_10512,N_14187);
nand U17350 (N_17350,N_14653,N_13927);
and U17351 (N_17351,N_14331,N_13179);
nand U17352 (N_17352,N_11580,N_14700);
and U17353 (N_17353,N_10964,N_12440);
xor U17354 (N_17354,N_13948,N_10031);
or U17355 (N_17355,N_11791,N_14454);
nor U17356 (N_17356,N_12570,N_12889);
nor U17357 (N_17357,N_12036,N_10739);
nor U17358 (N_17358,N_14979,N_12267);
nand U17359 (N_17359,N_12112,N_11033);
xor U17360 (N_17360,N_10842,N_12869);
nand U17361 (N_17361,N_12845,N_13908);
or U17362 (N_17362,N_11956,N_13691);
or U17363 (N_17363,N_10927,N_14089);
nand U17364 (N_17364,N_13777,N_13842);
nand U17365 (N_17365,N_10303,N_13526);
or U17366 (N_17366,N_13631,N_10226);
nor U17367 (N_17367,N_13671,N_14608);
or U17368 (N_17368,N_14493,N_11054);
and U17369 (N_17369,N_14861,N_10699);
xor U17370 (N_17370,N_13726,N_13111);
xnor U17371 (N_17371,N_12438,N_11171);
and U17372 (N_17372,N_11570,N_10088);
nor U17373 (N_17373,N_12670,N_10953);
or U17374 (N_17374,N_10955,N_12094);
xnor U17375 (N_17375,N_13041,N_10746);
and U17376 (N_17376,N_11990,N_10764);
nand U17377 (N_17377,N_10233,N_13950);
xor U17378 (N_17378,N_12245,N_13860);
or U17379 (N_17379,N_14732,N_13433);
or U17380 (N_17380,N_13747,N_14691);
xor U17381 (N_17381,N_11325,N_13213);
xnor U17382 (N_17382,N_10201,N_10010);
xor U17383 (N_17383,N_11335,N_13328);
nor U17384 (N_17384,N_14374,N_10694);
or U17385 (N_17385,N_11932,N_13082);
xnor U17386 (N_17386,N_10977,N_14796);
or U17387 (N_17387,N_11588,N_13423);
nand U17388 (N_17388,N_11799,N_12508);
and U17389 (N_17389,N_11637,N_13156);
xnor U17390 (N_17390,N_10544,N_13989);
xnor U17391 (N_17391,N_11363,N_12729);
nor U17392 (N_17392,N_13670,N_14286);
nor U17393 (N_17393,N_12916,N_12673);
xnor U17394 (N_17394,N_11813,N_12171);
nand U17395 (N_17395,N_10188,N_11096);
or U17396 (N_17396,N_13214,N_10563);
or U17397 (N_17397,N_10426,N_12361);
xor U17398 (N_17398,N_14354,N_12862);
or U17399 (N_17399,N_12362,N_11387);
and U17400 (N_17400,N_14590,N_12412);
xor U17401 (N_17401,N_13637,N_14280);
or U17402 (N_17402,N_11308,N_10747);
xnor U17403 (N_17403,N_13283,N_11888);
and U17404 (N_17404,N_14975,N_14211);
and U17405 (N_17405,N_12017,N_13932);
nand U17406 (N_17406,N_13417,N_10805);
and U17407 (N_17407,N_12458,N_14669);
or U17408 (N_17408,N_12754,N_10570);
and U17409 (N_17409,N_13231,N_14548);
and U17410 (N_17410,N_12905,N_11249);
and U17411 (N_17411,N_13370,N_12718);
or U17412 (N_17412,N_14070,N_11707);
xor U17413 (N_17413,N_11740,N_12128);
nand U17414 (N_17414,N_10253,N_10862);
and U17415 (N_17415,N_12843,N_11921);
nand U17416 (N_17416,N_12068,N_11228);
and U17417 (N_17417,N_13163,N_10921);
and U17418 (N_17418,N_14754,N_10364);
nor U17419 (N_17419,N_13639,N_10345);
or U17420 (N_17420,N_12330,N_12507);
and U17421 (N_17421,N_12269,N_12343);
xnor U17422 (N_17422,N_12157,N_14093);
nand U17423 (N_17423,N_14140,N_14476);
or U17424 (N_17424,N_14321,N_11976);
xor U17425 (N_17425,N_11719,N_11846);
nand U17426 (N_17426,N_13879,N_11770);
and U17427 (N_17427,N_10355,N_12383);
and U17428 (N_17428,N_14305,N_11125);
nor U17429 (N_17429,N_13871,N_10110);
or U17430 (N_17430,N_14534,N_11053);
nand U17431 (N_17431,N_11346,N_12761);
nand U17432 (N_17432,N_12858,N_10323);
or U17433 (N_17433,N_14230,N_13954);
xnor U17434 (N_17434,N_13724,N_13533);
nand U17435 (N_17435,N_12810,N_13768);
or U17436 (N_17436,N_11800,N_11804);
nand U17437 (N_17437,N_14468,N_13144);
nor U17438 (N_17438,N_12671,N_14019);
nor U17439 (N_17439,N_14446,N_14417);
nand U17440 (N_17440,N_14839,N_13322);
xnor U17441 (N_17441,N_13057,N_11599);
and U17442 (N_17442,N_11067,N_13106);
nand U17443 (N_17443,N_11210,N_11814);
and U17444 (N_17444,N_12456,N_12883);
nor U17445 (N_17445,N_14180,N_12020);
nor U17446 (N_17446,N_12360,N_11628);
nor U17447 (N_17447,N_13536,N_13135);
nand U17448 (N_17448,N_13608,N_10305);
nand U17449 (N_17449,N_13045,N_12723);
and U17450 (N_17450,N_12882,N_12873);
nand U17451 (N_17451,N_13204,N_13510);
and U17452 (N_17452,N_14824,N_13663);
or U17453 (N_17453,N_13912,N_12432);
nor U17454 (N_17454,N_12459,N_12165);
or U17455 (N_17455,N_12857,N_11901);
or U17456 (N_17456,N_13349,N_14283);
nor U17457 (N_17457,N_14001,N_14457);
nor U17458 (N_17458,N_11919,N_11139);
nand U17459 (N_17459,N_12895,N_10656);
nand U17460 (N_17460,N_13303,N_10022);
or U17461 (N_17461,N_11915,N_14812);
nand U17462 (N_17462,N_11232,N_14619);
nor U17463 (N_17463,N_13602,N_13951);
and U17464 (N_17464,N_10605,N_13494);
nor U17465 (N_17465,N_14087,N_11000);
nor U17466 (N_17466,N_12568,N_14386);
xnor U17467 (N_17467,N_14078,N_13162);
xor U17468 (N_17468,N_13083,N_12093);
xor U17469 (N_17469,N_11592,N_12760);
nand U17470 (N_17470,N_10174,N_13902);
nand U17471 (N_17471,N_12283,N_12622);
xnor U17472 (N_17472,N_14157,N_11487);
or U17473 (N_17473,N_13054,N_14546);
xnor U17474 (N_17474,N_12222,N_13121);
nand U17475 (N_17475,N_10347,N_10982);
or U17476 (N_17476,N_11246,N_13377);
and U17477 (N_17477,N_11275,N_13287);
xor U17478 (N_17478,N_10653,N_14665);
or U17479 (N_17479,N_12195,N_13489);
and U17480 (N_17480,N_10295,N_14985);
and U17481 (N_17481,N_14479,N_13332);
xor U17482 (N_17482,N_12912,N_14400);
xnor U17483 (N_17483,N_14916,N_10543);
xor U17484 (N_17484,N_12534,N_11769);
nor U17485 (N_17485,N_10940,N_13791);
and U17486 (N_17486,N_13765,N_12463);
and U17487 (N_17487,N_10227,N_11447);
or U17488 (N_17488,N_10677,N_14257);
nand U17489 (N_17489,N_13164,N_14122);
or U17490 (N_17490,N_12866,N_12490);
and U17491 (N_17491,N_12371,N_14375);
xor U17492 (N_17492,N_12515,N_13042);
or U17493 (N_17493,N_12152,N_10517);
nor U17494 (N_17494,N_10441,N_10058);
nor U17495 (N_17495,N_14149,N_13295);
xnor U17496 (N_17496,N_14488,N_14013);
nor U17497 (N_17497,N_11150,N_11107);
xor U17498 (N_17498,N_11082,N_12792);
xor U17499 (N_17499,N_10053,N_12925);
xnor U17500 (N_17500,N_14911,N_13893);
and U17501 (N_17501,N_12317,N_10656);
and U17502 (N_17502,N_12798,N_13441);
or U17503 (N_17503,N_11367,N_13236);
nand U17504 (N_17504,N_14737,N_10307);
nand U17505 (N_17505,N_13186,N_10987);
and U17506 (N_17506,N_13027,N_10452);
xor U17507 (N_17507,N_10278,N_12896);
nor U17508 (N_17508,N_12447,N_10837);
nor U17509 (N_17509,N_11065,N_13734);
nor U17510 (N_17510,N_10897,N_11575);
xnor U17511 (N_17511,N_14608,N_12273);
nor U17512 (N_17512,N_12033,N_10566);
xnor U17513 (N_17513,N_12033,N_14020);
and U17514 (N_17514,N_10043,N_10306);
nand U17515 (N_17515,N_12106,N_11327);
or U17516 (N_17516,N_14569,N_11788);
and U17517 (N_17517,N_13202,N_12114);
and U17518 (N_17518,N_12221,N_12690);
xor U17519 (N_17519,N_11622,N_10130);
xor U17520 (N_17520,N_10671,N_13845);
nor U17521 (N_17521,N_10412,N_11622);
and U17522 (N_17522,N_12390,N_10453);
xor U17523 (N_17523,N_14565,N_10553);
nand U17524 (N_17524,N_12323,N_11474);
xor U17525 (N_17525,N_14635,N_13469);
nand U17526 (N_17526,N_10957,N_12094);
nor U17527 (N_17527,N_12171,N_13244);
nand U17528 (N_17528,N_11291,N_12270);
and U17529 (N_17529,N_14032,N_11282);
xnor U17530 (N_17530,N_12920,N_14992);
and U17531 (N_17531,N_11238,N_12392);
nor U17532 (N_17532,N_12970,N_12633);
nor U17533 (N_17533,N_12600,N_11071);
nor U17534 (N_17534,N_10371,N_14443);
nor U17535 (N_17535,N_14736,N_14633);
and U17536 (N_17536,N_11989,N_14649);
xor U17537 (N_17537,N_11938,N_11029);
nand U17538 (N_17538,N_11450,N_11014);
or U17539 (N_17539,N_11972,N_12716);
xnor U17540 (N_17540,N_10802,N_14624);
xor U17541 (N_17541,N_13507,N_14468);
nor U17542 (N_17542,N_12222,N_13158);
nand U17543 (N_17543,N_11149,N_11127);
or U17544 (N_17544,N_12976,N_14756);
or U17545 (N_17545,N_13651,N_14830);
nand U17546 (N_17546,N_11476,N_10131);
nand U17547 (N_17547,N_12987,N_11735);
xor U17548 (N_17548,N_10854,N_12550);
or U17549 (N_17549,N_10728,N_10713);
and U17550 (N_17550,N_11399,N_10442);
nand U17551 (N_17551,N_14833,N_14636);
and U17552 (N_17552,N_13160,N_12062);
or U17553 (N_17553,N_12851,N_13458);
xor U17554 (N_17554,N_10091,N_10214);
or U17555 (N_17555,N_10248,N_14132);
nor U17556 (N_17556,N_11806,N_12336);
xor U17557 (N_17557,N_14090,N_14934);
xor U17558 (N_17558,N_12477,N_10055);
xnor U17559 (N_17559,N_14522,N_11389);
nand U17560 (N_17560,N_10659,N_12521);
nand U17561 (N_17561,N_13633,N_13868);
nand U17562 (N_17562,N_12883,N_11151);
nand U17563 (N_17563,N_14736,N_13377);
nand U17564 (N_17564,N_10973,N_13880);
or U17565 (N_17565,N_13089,N_11292);
xnor U17566 (N_17566,N_11730,N_11209);
or U17567 (N_17567,N_11528,N_13948);
and U17568 (N_17568,N_13551,N_12050);
and U17569 (N_17569,N_12053,N_10067);
or U17570 (N_17570,N_12642,N_12626);
and U17571 (N_17571,N_13138,N_12565);
nand U17572 (N_17572,N_14993,N_12121);
xnor U17573 (N_17573,N_12365,N_14827);
nand U17574 (N_17574,N_12381,N_14901);
nand U17575 (N_17575,N_14158,N_13034);
nor U17576 (N_17576,N_10749,N_13359);
nor U17577 (N_17577,N_11468,N_10456);
nor U17578 (N_17578,N_13556,N_14413);
or U17579 (N_17579,N_14323,N_11893);
and U17580 (N_17580,N_10449,N_13698);
and U17581 (N_17581,N_13787,N_12366);
or U17582 (N_17582,N_12260,N_10869);
and U17583 (N_17583,N_11539,N_11288);
and U17584 (N_17584,N_10810,N_10350);
nand U17585 (N_17585,N_11411,N_10697);
or U17586 (N_17586,N_11501,N_10003);
nor U17587 (N_17587,N_11327,N_14202);
xnor U17588 (N_17588,N_13676,N_12325);
nand U17589 (N_17589,N_14433,N_13764);
xor U17590 (N_17590,N_11683,N_11982);
nand U17591 (N_17591,N_12858,N_10070);
nand U17592 (N_17592,N_10761,N_13001);
nor U17593 (N_17593,N_11357,N_14409);
nor U17594 (N_17594,N_14964,N_14725);
xnor U17595 (N_17595,N_14643,N_13208);
xor U17596 (N_17596,N_11200,N_10465);
nand U17597 (N_17597,N_12096,N_14199);
nor U17598 (N_17598,N_12123,N_10612);
xnor U17599 (N_17599,N_13869,N_14464);
nand U17600 (N_17600,N_10618,N_10944);
nand U17601 (N_17601,N_11981,N_14720);
xnor U17602 (N_17602,N_11633,N_10857);
xor U17603 (N_17603,N_11834,N_13061);
nor U17604 (N_17604,N_11272,N_11935);
nor U17605 (N_17605,N_13837,N_12389);
nand U17606 (N_17606,N_11185,N_14459);
and U17607 (N_17607,N_13627,N_11009);
xnor U17608 (N_17608,N_11207,N_14324);
nand U17609 (N_17609,N_10618,N_10437);
xor U17610 (N_17610,N_11483,N_10044);
nand U17611 (N_17611,N_13481,N_10336);
and U17612 (N_17612,N_12777,N_10955);
or U17613 (N_17613,N_12365,N_14816);
or U17614 (N_17614,N_13936,N_14262);
xnor U17615 (N_17615,N_14510,N_10112);
xnor U17616 (N_17616,N_12746,N_10642);
xnor U17617 (N_17617,N_14729,N_13135);
or U17618 (N_17618,N_10960,N_13895);
nand U17619 (N_17619,N_14905,N_14536);
xnor U17620 (N_17620,N_11459,N_13562);
xor U17621 (N_17621,N_11772,N_10222);
nand U17622 (N_17622,N_11692,N_11867);
nand U17623 (N_17623,N_10502,N_14744);
or U17624 (N_17624,N_11456,N_10615);
nand U17625 (N_17625,N_13783,N_11501);
xor U17626 (N_17626,N_13777,N_11479);
or U17627 (N_17627,N_11016,N_13598);
xor U17628 (N_17628,N_10749,N_13205);
nand U17629 (N_17629,N_12628,N_11208);
or U17630 (N_17630,N_10175,N_14817);
xor U17631 (N_17631,N_13304,N_12389);
xnor U17632 (N_17632,N_12131,N_11818);
nor U17633 (N_17633,N_13229,N_12179);
nand U17634 (N_17634,N_14685,N_12379);
nor U17635 (N_17635,N_13154,N_13254);
xnor U17636 (N_17636,N_12865,N_14200);
or U17637 (N_17637,N_11406,N_13828);
and U17638 (N_17638,N_14308,N_13272);
nor U17639 (N_17639,N_13421,N_14697);
xor U17640 (N_17640,N_14800,N_14566);
nand U17641 (N_17641,N_12665,N_14327);
or U17642 (N_17642,N_14077,N_12402);
xnor U17643 (N_17643,N_13386,N_10054);
and U17644 (N_17644,N_10451,N_14982);
nor U17645 (N_17645,N_14036,N_12990);
nor U17646 (N_17646,N_13682,N_10287);
nor U17647 (N_17647,N_14301,N_11956);
and U17648 (N_17648,N_14773,N_14960);
nand U17649 (N_17649,N_11472,N_13307);
or U17650 (N_17650,N_10062,N_12604);
nor U17651 (N_17651,N_10429,N_14455);
xnor U17652 (N_17652,N_11836,N_11902);
nor U17653 (N_17653,N_13272,N_14108);
nand U17654 (N_17654,N_11939,N_14909);
nand U17655 (N_17655,N_14005,N_11756);
nor U17656 (N_17656,N_14834,N_10528);
and U17657 (N_17657,N_12243,N_13558);
nor U17658 (N_17658,N_14017,N_10239);
xnor U17659 (N_17659,N_12009,N_11109);
nand U17660 (N_17660,N_13636,N_13839);
and U17661 (N_17661,N_10394,N_11521);
xnor U17662 (N_17662,N_12073,N_11175);
or U17663 (N_17663,N_14880,N_13432);
and U17664 (N_17664,N_13171,N_13726);
nor U17665 (N_17665,N_13717,N_11105);
nor U17666 (N_17666,N_11958,N_13854);
and U17667 (N_17667,N_12982,N_13988);
and U17668 (N_17668,N_13116,N_12087);
nor U17669 (N_17669,N_11982,N_10171);
nand U17670 (N_17670,N_12249,N_14948);
xnor U17671 (N_17671,N_12765,N_12106);
nor U17672 (N_17672,N_13015,N_10562);
nor U17673 (N_17673,N_10159,N_11550);
nor U17674 (N_17674,N_10706,N_14916);
or U17675 (N_17675,N_12966,N_14787);
nand U17676 (N_17676,N_10768,N_11056);
and U17677 (N_17677,N_13260,N_12443);
or U17678 (N_17678,N_13009,N_14922);
and U17679 (N_17679,N_10494,N_12108);
nor U17680 (N_17680,N_12263,N_13691);
nand U17681 (N_17681,N_12290,N_13959);
or U17682 (N_17682,N_10742,N_13885);
and U17683 (N_17683,N_11130,N_13753);
nand U17684 (N_17684,N_11106,N_12540);
or U17685 (N_17685,N_10103,N_12104);
nand U17686 (N_17686,N_14092,N_12495);
nand U17687 (N_17687,N_11971,N_13386);
or U17688 (N_17688,N_10331,N_14811);
nand U17689 (N_17689,N_13823,N_10127);
xnor U17690 (N_17690,N_13516,N_12628);
nand U17691 (N_17691,N_11429,N_12406);
or U17692 (N_17692,N_10876,N_13450);
nor U17693 (N_17693,N_11959,N_10549);
nand U17694 (N_17694,N_14967,N_14497);
and U17695 (N_17695,N_12005,N_14307);
nor U17696 (N_17696,N_10974,N_13240);
xnor U17697 (N_17697,N_11738,N_14941);
and U17698 (N_17698,N_10474,N_14118);
xor U17699 (N_17699,N_13897,N_10177);
nor U17700 (N_17700,N_14072,N_14834);
nor U17701 (N_17701,N_12201,N_10030);
nor U17702 (N_17702,N_10530,N_11718);
xnor U17703 (N_17703,N_14748,N_11273);
nor U17704 (N_17704,N_11649,N_10044);
xnor U17705 (N_17705,N_13120,N_13694);
nor U17706 (N_17706,N_10393,N_10811);
and U17707 (N_17707,N_10919,N_13601);
xor U17708 (N_17708,N_11580,N_13193);
and U17709 (N_17709,N_11835,N_10195);
nand U17710 (N_17710,N_13796,N_12850);
nand U17711 (N_17711,N_14798,N_10217);
and U17712 (N_17712,N_11738,N_10349);
nand U17713 (N_17713,N_10445,N_12178);
nor U17714 (N_17714,N_13446,N_13588);
and U17715 (N_17715,N_11908,N_13298);
or U17716 (N_17716,N_13212,N_12885);
nand U17717 (N_17717,N_10920,N_14541);
nor U17718 (N_17718,N_11612,N_10993);
xor U17719 (N_17719,N_12777,N_10167);
and U17720 (N_17720,N_11666,N_10667);
or U17721 (N_17721,N_12819,N_12126);
and U17722 (N_17722,N_14575,N_14065);
nor U17723 (N_17723,N_10281,N_11330);
xor U17724 (N_17724,N_11082,N_11162);
nor U17725 (N_17725,N_10690,N_13544);
or U17726 (N_17726,N_13054,N_10283);
and U17727 (N_17727,N_10263,N_10310);
or U17728 (N_17728,N_11654,N_14886);
nand U17729 (N_17729,N_10597,N_13393);
nor U17730 (N_17730,N_10875,N_12988);
nor U17731 (N_17731,N_13384,N_12638);
nand U17732 (N_17732,N_10174,N_14824);
or U17733 (N_17733,N_10988,N_11358);
or U17734 (N_17734,N_12106,N_10401);
nand U17735 (N_17735,N_14581,N_11833);
xor U17736 (N_17736,N_12368,N_14318);
nor U17737 (N_17737,N_14842,N_14191);
and U17738 (N_17738,N_10181,N_10107);
nor U17739 (N_17739,N_11056,N_10132);
and U17740 (N_17740,N_11718,N_10727);
nand U17741 (N_17741,N_12940,N_13611);
nor U17742 (N_17742,N_11244,N_14282);
nand U17743 (N_17743,N_11978,N_10442);
xor U17744 (N_17744,N_13968,N_14410);
or U17745 (N_17745,N_13176,N_11285);
nand U17746 (N_17746,N_12231,N_14155);
nand U17747 (N_17747,N_12729,N_11467);
and U17748 (N_17748,N_11774,N_14287);
nor U17749 (N_17749,N_13943,N_14890);
xnor U17750 (N_17750,N_10707,N_12957);
nor U17751 (N_17751,N_11227,N_14167);
nand U17752 (N_17752,N_10981,N_13448);
or U17753 (N_17753,N_13361,N_11984);
and U17754 (N_17754,N_14535,N_10104);
xnor U17755 (N_17755,N_10844,N_10517);
or U17756 (N_17756,N_11834,N_13687);
xor U17757 (N_17757,N_11946,N_11986);
or U17758 (N_17758,N_12105,N_14034);
nor U17759 (N_17759,N_11069,N_11482);
nor U17760 (N_17760,N_10208,N_14540);
nor U17761 (N_17761,N_13695,N_11532);
and U17762 (N_17762,N_13396,N_12091);
and U17763 (N_17763,N_13048,N_13506);
nor U17764 (N_17764,N_14206,N_10993);
and U17765 (N_17765,N_11711,N_14370);
xor U17766 (N_17766,N_12068,N_11953);
xor U17767 (N_17767,N_10542,N_10096);
nand U17768 (N_17768,N_14866,N_11290);
or U17769 (N_17769,N_14437,N_14168);
nor U17770 (N_17770,N_12085,N_11575);
and U17771 (N_17771,N_13565,N_10231);
xor U17772 (N_17772,N_10870,N_14980);
and U17773 (N_17773,N_10401,N_14384);
and U17774 (N_17774,N_12551,N_11516);
nand U17775 (N_17775,N_12296,N_11521);
and U17776 (N_17776,N_13048,N_11423);
nor U17777 (N_17777,N_11426,N_13847);
or U17778 (N_17778,N_14919,N_12757);
and U17779 (N_17779,N_12459,N_11684);
nand U17780 (N_17780,N_12366,N_13509);
nor U17781 (N_17781,N_13123,N_13671);
or U17782 (N_17782,N_13276,N_10999);
nand U17783 (N_17783,N_10255,N_13591);
xnor U17784 (N_17784,N_12534,N_13639);
xnor U17785 (N_17785,N_12174,N_12754);
nand U17786 (N_17786,N_12798,N_11543);
nand U17787 (N_17787,N_11224,N_12108);
nand U17788 (N_17788,N_13420,N_12822);
xnor U17789 (N_17789,N_13572,N_10488);
nor U17790 (N_17790,N_13306,N_13016);
nand U17791 (N_17791,N_13603,N_12310);
or U17792 (N_17792,N_12693,N_11218);
or U17793 (N_17793,N_13851,N_13976);
nand U17794 (N_17794,N_10992,N_10516);
nor U17795 (N_17795,N_10291,N_13848);
xor U17796 (N_17796,N_14797,N_11499);
xnor U17797 (N_17797,N_14248,N_14093);
and U17798 (N_17798,N_13411,N_10704);
and U17799 (N_17799,N_12878,N_10026);
nor U17800 (N_17800,N_11452,N_12882);
and U17801 (N_17801,N_12607,N_13129);
and U17802 (N_17802,N_10254,N_11195);
xnor U17803 (N_17803,N_14687,N_13617);
or U17804 (N_17804,N_13775,N_14561);
and U17805 (N_17805,N_13350,N_10848);
and U17806 (N_17806,N_11658,N_10799);
nand U17807 (N_17807,N_12504,N_10379);
and U17808 (N_17808,N_11224,N_10606);
or U17809 (N_17809,N_11888,N_10275);
and U17810 (N_17810,N_14361,N_12307);
nand U17811 (N_17811,N_12196,N_13199);
or U17812 (N_17812,N_11362,N_10439);
xor U17813 (N_17813,N_12614,N_11552);
nor U17814 (N_17814,N_10944,N_14185);
and U17815 (N_17815,N_11040,N_13260);
nand U17816 (N_17816,N_12782,N_12584);
and U17817 (N_17817,N_13252,N_11402);
and U17818 (N_17818,N_14032,N_14377);
nand U17819 (N_17819,N_10027,N_10786);
nor U17820 (N_17820,N_12187,N_10033);
and U17821 (N_17821,N_14786,N_14549);
xnor U17822 (N_17822,N_13418,N_13564);
nor U17823 (N_17823,N_11935,N_13012);
xnor U17824 (N_17824,N_11680,N_12045);
and U17825 (N_17825,N_11753,N_12672);
or U17826 (N_17826,N_12269,N_10751);
and U17827 (N_17827,N_14267,N_12081);
nor U17828 (N_17828,N_10632,N_14330);
nor U17829 (N_17829,N_12326,N_12415);
xnor U17830 (N_17830,N_11058,N_14706);
xor U17831 (N_17831,N_13344,N_13166);
nand U17832 (N_17832,N_12493,N_12437);
and U17833 (N_17833,N_13559,N_14281);
nand U17834 (N_17834,N_10568,N_14204);
xor U17835 (N_17835,N_13546,N_11565);
nor U17836 (N_17836,N_12905,N_11562);
nor U17837 (N_17837,N_14638,N_13676);
nor U17838 (N_17838,N_13135,N_13764);
nor U17839 (N_17839,N_11018,N_12070);
nor U17840 (N_17840,N_13112,N_14865);
or U17841 (N_17841,N_13565,N_13550);
xnor U17842 (N_17842,N_12304,N_10981);
nand U17843 (N_17843,N_13047,N_13267);
or U17844 (N_17844,N_10656,N_12343);
and U17845 (N_17845,N_12479,N_14652);
xor U17846 (N_17846,N_14031,N_10090);
or U17847 (N_17847,N_12599,N_11876);
or U17848 (N_17848,N_12319,N_14333);
nor U17849 (N_17849,N_11840,N_13654);
nand U17850 (N_17850,N_13802,N_12065);
nand U17851 (N_17851,N_13198,N_13352);
and U17852 (N_17852,N_14399,N_13162);
or U17853 (N_17853,N_11034,N_12060);
nor U17854 (N_17854,N_12560,N_11195);
xor U17855 (N_17855,N_10256,N_10935);
or U17856 (N_17856,N_14245,N_12440);
nand U17857 (N_17857,N_10987,N_11606);
xnor U17858 (N_17858,N_13322,N_12614);
xor U17859 (N_17859,N_12822,N_12188);
nand U17860 (N_17860,N_13270,N_10494);
xor U17861 (N_17861,N_10768,N_11952);
or U17862 (N_17862,N_14395,N_13886);
and U17863 (N_17863,N_11003,N_14844);
or U17864 (N_17864,N_14526,N_13440);
nand U17865 (N_17865,N_12850,N_10684);
nand U17866 (N_17866,N_11228,N_13222);
nand U17867 (N_17867,N_12241,N_11009);
or U17868 (N_17868,N_11200,N_12070);
nand U17869 (N_17869,N_12115,N_14247);
or U17870 (N_17870,N_11896,N_14297);
nor U17871 (N_17871,N_11731,N_13936);
xor U17872 (N_17872,N_14010,N_10454);
and U17873 (N_17873,N_12118,N_13300);
nand U17874 (N_17874,N_12185,N_13902);
nand U17875 (N_17875,N_10165,N_11409);
or U17876 (N_17876,N_11430,N_10885);
nand U17877 (N_17877,N_10416,N_14079);
nor U17878 (N_17878,N_14559,N_14031);
and U17879 (N_17879,N_14306,N_14921);
nand U17880 (N_17880,N_13654,N_11402);
nor U17881 (N_17881,N_12952,N_14225);
or U17882 (N_17882,N_14872,N_13454);
and U17883 (N_17883,N_13558,N_10495);
xor U17884 (N_17884,N_12354,N_11955);
xor U17885 (N_17885,N_12688,N_10047);
or U17886 (N_17886,N_10392,N_10286);
nor U17887 (N_17887,N_13944,N_12762);
nor U17888 (N_17888,N_14048,N_12474);
or U17889 (N_17889,N_12532,N_10504);
and U17890 (N_17890,N_12379,N_13808);
nand U17891 (N_17891,N_11265,N_11522);
nor U17892 (N_17892,N_12011,N_12659);
or U17893 (N_17893,N_12117,N_10212);
or U17894 (N_17894,N_11867,N_10354);
or U17895 (N_17895,N_13794,N_14890);
or U17896 (N_17896,N_12276,N_11893);
or U17897 (N_17897,N_11641,N_14042);
nand U17898 (N_17898,N_11422,N_10525);
xor U17899 (N_17899,N_10815,N_11013);
or U17900 (N_17900,N_14066,N_14937);
nor U17901 (N_17901,N_10489,N_13264);
and U17902 (N_17902,N_10669,N_14120);
and U17903 (N_17903,N_14694,N_11341);
nor U17904 (N_17904,N_12248,N_14118);
and U17905 (N_17905,N_14956,N_10299);
and U17906 (N_17906,N_14902,N_12748);
nand U17907 (N_17907,N_14714,N_10667);
nor U17908 (N_17908,N_11988,N_10984);
and U17909 (N_17909,N_11823,N_11589);
or U17910 (N_17910,N_13229,N_12151);
nor U17911 (N_17911,N_13046,N_13495);
and U17912 (N_17912,N_10633,N_11154);
nand U17913 (N_17913,N_12936,N_11394);
nand U17914 (N_17914,N_10986,N_14784);
and U17915 (N_17915,N_12480,N_11352);
and U17916 (N_17916,N_12855,N_11026);
nor U17917 (N_17917,N_12093,N_12403);
or U17918 (N_17918,N_12096,N_11392);
xnor U17919 (N_17919,N_14383,N_10187);
or U17920 (N_17920,N_10550,N_14173);
and U17921 (N_17921,N_13470,N_10258);
or U17922 (N_17922,N_10410,N_13226);
nand U17923 (N_17923,N_11438,N_13965);
or U17924 (N_17924,N_12960,N_11639);
xor U17925 (N_17925,N_10940,N_13647);
xor U17926 (N_17926,N_13181,N_13911);
and U17927 (N_17927,N_10148,N_12470);
and U17928 (N_17928,N_11964,N_14183);
nand U17929 (N_17929,N_12450,N_10538);
and U17930 (N_17930,N_12322,N_10750);
or U17931 (N_17931,N_10943,N_11796);
or U17932 (N_17932,N_10900,N_11594);
nand U17933 (N_17933,N_11780,N_10093);
or U17934 (N_17934,N_10396,N_10942);
or U17935 (N_17935,N_13710,N_12636);
and U17936 (N_17936,N_10321,N_12437);
nor U17937 (N_17937,N_12208,N_10655);
nor U17938 (N_17938,N_12144,N_10834);
nand U17939 (N_17939,N_14823,N_14542);
and U17940 (N_17940,N_10221,N_14683);
and U17941 (N_17941,N_11053,N_14287);
nand U17942 (N_17942,N_11908,N_13614);
nor U17943 (N_17943,N_12468,N_13019);
xnor U17944 (N_17944,N_13664,N_14958);
nor U17945 (N_17945,N_13116,N_12784);
xnor U17946 (N_17946,N_13845,N_14089);
xnor U17947 (N_17947,N_13986,N_10423);
nor U17948 (N_17948,N_11597,N_10761);
and U17949 (N_17949,N_12553,N_11146);
nor U17950 (N_17950,N_13825,N_13580);
or U17951 (N_17951,N_14676,N_14912);
nor U17952 (N_17952,N_11961,N_10940);
xnor U17953 (N_17953,N_11834,N_10724);
or U17954 (N_17954,N_11280,N_12739);
xnor U17955 (N_17955,N_14295,N_14816);
or U17956 (N_17956,N_14464,N_10935);
xor U17957 (N_17957,N_13077,N_13656);
nand U17958 (N_17958,N_14444,N_14999);
and U17959 (N_17959,N_10201,N_10848);
and U17960 (N_17960,N_11003,N_10993);
nor U17961 (N_17961,N_10725,N_14561);
and U17962 (N_17962,N_11279,N_11026);
nand U17963 (N_17963,N_14093,N_12261);
or U17964 (N_17964,N_12154,N_10882);
nand U17965 (N_17965,N_14759,N_11599);
xnor U17966 (N_17966,N_13640,N_13529);
or U17967 (N_17967,N_13639,N_14909);
and U17968 (N_17968,N_14404,N_10341);
or U17969 (N_17969,N_12811,N_12987);
xnor U17970 (N_17970,N_12045,N_14556);
xor U17971 (N_17971,N_12843,N_10830);
nand U17972 (N_17972,N_14694,N_12365);
nand U17973 (N_17973,N_14894,N_13324);
or U17974 (N_17974,N_12541,N_11665);
nor U17975 (N_17975,N_12716,N_13348);
or U17976 (N_17976,N_11007,N_10300);
nor U17977 (N_17977,N_14288,N_10521);
nand U17978 (N_17978,N_12045,N_11629);
nor U17979 (N_17979,N_13749,N_14048);
nor U17980 (N_17980,N_14096,N_12803);
and U17981 (N_17981,N_12489,N_13999);
nand U17982 (N_17982,N_13193,N_10449);
nor U17983 (N_17983,N_11041,N_14698);
xor U17984 (N_17984,N_13548,N_12656);
nand U17985 (N_17985,N_14878,N_13105);
nand U17986 (N_17986,N_14976,N_13941);
xnor U17987 (N_17987,N_12851,N_12975);
nand U17988 (N_17988,N_11225,N_10358);
nand U17989 (N_17989,N_10225,N_14695);
nand U17990 (N_17990,N_12465,N_10303);
nor U17991 (N_17991,N_12408,N_14799);
nor U17992 (N_17992,N_11379,N_10970);
nor U17993 (N_17993,N_10158,N_10501);
nor U17994 (N_17994,N_12916,N_11369);
nand U17995 (N_17995,N_10170,N_12926);
nand U17996 (N_17996,N_13267,N_12981);
xnor U17997 (N_17997,N_11411,N_10514);
xor U17998 (N_17998,N_13362,N_12053);
xnor U17999 (N_17999,N_10992,N_11385);
nor U18000 (N_18000,N_11159,N_13528);
xor U18001 (N_18001,N_10457,N_12288);
and U18002 (N_18002,N_10727,N_13402);
xnor U18003 (N_18003,N_13536,N_10152);
or U18004 (N_18004,N_13609,N_12903);
or U18005 (N_18005,N_12462,N_14164);
xnor U18006 (N_18006,N_10496,N_13292);
nand U18007 (N_18007,N_10928,N_10932);
nor U18008 (N_18008,N_10334,N_11833);
nor U18009 (N_18009,N_14082,N_13822);
nor U18010 (N_18010,N_10314,N_14699);
nor U18011 (N_18011,N_12837,N_14409);
and U18012 (N_18012,N_14084,N_10224);
and U18013 (N_18013,N_13227,N_12633);
xor U18014 (N_18014,N_11578,N_13762);
nand U18015 (N_18015,N_11098,N_11413);
or U18016 (N_18016,N_13919,N_12361);
nor U18017 (N_18017,N_10267,N_12237);
and U18018 (N_18018,N_14846,N_10467);
nand U18019 (N_18019,N_14924,N_13285);
or U18020 (N_18020,N_11131,N_11843);
nor U18021 (N_18021,N_12081,N_13211);
or U18022 (N_18022,N_13504,N_10536);
or U18023 (N_18023,N_10945,N_10266);
nor U18024 (N_18024,N_11531,N_14679);
nor U18025 (N_18025,N_14569,N_13161);
nor U18026 (N_18026,N_13962,N_13884);
nand U18027 (N_18027,N_13446,N_14114);
xnor U18028 (N_18028,N_12216,N_10560);
or U18029 (N_18029,N_10524,N_10975);
xor U18030 (N_18030,N_12074,N_10356);
and U18031 (N_18031,N_10128,N_14991);
or U18032 (N_18032,N_12621,N_10552);
and U18033 (N_18033,N_10697,N_10242);
and U18034 (N_18034,N_13568,N_11676);
nand U18035 (N_18035,N_10248,N_12201);
xnor U18036 (N_18036,N_14921,N_10509);
and U18037 (N_18037,N_10954,N_10350);
nand U18038 (N_18038,N_14616,N_12502);
nor U18039 (N_18039,N_10675,N_10169);
nor U18040 (N_18040,N_11067,N_12884);
and U18041 (N_18041,N_14236,N_11687);
or U18042 (N_18042,N_14694,N_10576);
nor U18043 (N_18043,N_10628,N_14824);
nand U18044 (N_18044,N_13316,N_14744);
or U18045 (N_18045,N_10455,N_10525);
xnor U18046 (N_18046,N_13915,N_14119);
and U18047 (N_18047,N_10532,N_10658);
xnor U18048 (N_18048,N_10129,N_14568);
nor U18049 (N_18049,N_12533,N_11354);
nor U18050 (N_18050,N_11814,N_10436);
and U18051 (N_18051,N_12448,N_10717);
nor U18052 (N_18052,N_12379,N_10414);
and U18053 (N_18053,N_13205,N_12065);
or U18054 (N_18054,N_13965,N_13469);
nor U18055 (N_18055,N_14628,N_11713);
nand U18056 (N_18056,N_14098,N_10263);
and U18057 (N_18057,N_11544,N_12427);
nor U18058 (N_18058,N_14975,N_14478);
xnor U18059 (N_18059,N_11043,N_11590);
xor U18060 (N_18060,N_11595,N_10277);
and U18061 (N_18061,N_12201,N_13758);
and U18062 (N_18062,N_13650,N_13567);
nand U18063 (N_18063,N_12064,N_10774);
nor U18064 (N_18064,N_13331,N_14079);
nand U18065 (N_18065,N_10115,N_14196);
nand U18066 (N_18066,N_11803,N_13831);
and U18067 (N_18067,N_14435,N_10303);
nor U18068 (N_18068,N_11825,N_11315);
nor U18069 (N_18069,N_14945,N_13879);
nand U18070 (N_18070,N_12914,N_11861);
and U18071 (N_18071,N_13363,N_11426);
nand U18072 (N_18072,N_10789,N_13554);
nor U18073 (N_18073,N_12652,N_14729);
or U18074 (N_18074,N_13221,N_13537);
nor U18075 (N_18075,N_14495,N_10837);
nor U18076 (N_18076,N_12948,N_12924);
xor U18077 (N_18077,N_14133,N_11006);
nor U18078 (N_18078,N_14552,N_10236);
xnor U18079 (N_18079,N_10894,N_11232);
or U18080 (N_18080,N_14891,N_10491);
nor U18081 (N_18081,N_13132,N_13836);
xor U18082 (N_18082,N_11096,N_10508);
nor U18083 (N_18083,N_13722,N_13303);
and U18084 (N_18084,N_12945,N_12030);
nor U18085 (N_18085,N_11331,N_12547);
nand U18086 (N_18086,N_11748,N_13845);
nor U18087 (N_18087,N_13236,N_12830);
or U18088 (N_18088,N_10245,N_13685);
nor U18089 (N_18089,N_13040,N_12467);
or U18090 (N_18090,N_12597,N_10218);
xor U18091 (N_18091,N_12851,N_14833);
or U18092 (N_18092,N_14631,N_11152);
nand U18093 (N_18093,N_11532,N_10187);
and U18094 (N_18094,N_12743,N_14276);
nor U18095 (N_18095,N_12059,N_12313);
nor U18096 (N_18096,N_12206,N_12081);
xor U18097 (N_18097,N_14622,N_12848);
xnor U18098 (N_18098,N_11868,N_11953);
xor U18099 (N_18099,N_11971,N_14493);
and U18100 (N_18100,N_14185,N_14327);
or U18101 (N_18101,N_14427,N_10488);
and U18102 (N_18102,N_10777,N_14488);
xnor U18103 (N_18103,N_12141,N_13871);
nor U18104 (N_18104,N_12597,N_11709);
and U18105 (N_18105,N_11216,N_11888);
xnor U18106 (N_18106,N_11238,N_12172);
xnor U18107 (N_18107,N_14459,N_11112);
and U18108 (N_18108,N_13886,N_10478);
xor U18109 (N_18109,N_11479,N_11545);
xor U18110 (N_18110,N_12602,N_12919);
xor U18111 (N_18111,N_12190,N_11172);
and U18112 (N_18112,N_11382,N_10109);
or U18113 (N_18113,N_12259,N_11275);
nand U18114 (N_18114,N_13229,N_11075);
xnor U18115 (N_18115,N_13246,N_14133);
nand U18116 (N_18116,N_12117,N_14143);
or U18117 (N_18117,N_12879,N_13432);
and U18118 (N_18118,N_12434,N_14024);
and U18119 (N_18119,N_14609,N_12524);
nand U18120 (N_18120,N_14214,N_13208);
nor U18121 (N_18121,N_12859,N_11440);
nor U18122 (N_18122,N_14149,N_10298);
xor U18123 (N_18123,N_11139,N_12485);
nand U18124 (N_18124,N_14291,N_13297);
or U18125 (N_18125,N_11375,N_13044);
nand U18126 (N_18126,N_11379,N_13052);
nand U18127 (N_18127,N_11257,N_10235);
or U18128 (N_18128,N_10883,N_13857);
nor U18129 (N_18129,N_13862,N_12365);
nand U18130 (N_18130,N_13877,N_11633);
nand U18131 (N_18131,N_10327,N_12557);
nor U18132 (N_18132,N_10000,N_14522);
or U18133 (N_18133,N_11251,N_13937);
nand U18134 (N_18134,N_10831,N_11654);
and U18135 (N_18135,N_14844,N_14994);
nor U18136 (N_18136,N_13776,N_11572);
xnor U18137 (N_18137,N_12898,N_10929);
nand U18138 (N_18138,N_12703,N_14771);
nor U18139 (N_18139,N_13370,N_11191);
or U18140 (N_18140,N_13498,N_14581);
or U18141 (N_18141,N_13202,N_10733);
nand U18142 (N_18142,N_11355,N_12506);
nand U18143 (N_18143,N_14829,N_12383);
and U18144 (N_18144,N_10585,N_10638);
xor U18145 (N_18145,N_12187,N_13839);
nor U18146 (N_18146,N_13253,N_10905);
and U18147 (N_18147,N_12463,N_14273);
nand U18148 (N_18148,N_12806,N_10849);
nand U18149 (N_18149,N_10357,N_10125);
or U18150 (N_18150,N_10132,N_14973);
nor U18151 (N_18151,N_13308,N_12185);
and U18152 (N_18152,N_11458,N_14781);
or U18153 (N_18153,N_14224,N_11823);
nand U18154 (N_18154,N_14428,N_12405);
or U18155 (N_18155,N_10920,N_14977);
and U18156 (N_18156,N_10412,N_12949);
nor U18157 (N_18157,N_14154,N_14711);
or U18158 (N_18158,N_13373,N_10969);
nor U18159 (N_18159,N_11015,N_13689);
or U18160 (N_18160,N_12860,N_12983);
xnor U18161 (N_18161,N_13365,N_10258);
xor U18162 (N_18162,N_12128,N_11668);
xor U18163 (N_18163,N_11224,N_14967);
nor U18164 (N_18164,N_14003,N_14481);
nand U18165 (N_18165,N_10157,N_12363);
and U18166 (N_18166,N_11769,N_13866);
and U18167 (N_18167,N_10435,N_10574);
or U18168 (N_18168,N_14818,N_14638);
nand U18169 (N_18169,N_10114,N_13872);
nand U18170 (N_18170,N_10886,N_14817);
and U18171 (N_18171,N_10600,N_11346);
nand U18172 (N_18172,N_10204,N_10603);
and U18173 (N_18173,N_11586,N_14479);
nand U18174 (N_18174,N_12779,N_13520);
xor U18175 (N_18175,N_14116,N_10107);
xnor U18176 (N_18176,N_13416,N_14964);
nand U18177 (N_18177,N_14315,N_13795);
and U18178 (N_18178,N_12491,N_13783);
xnor U18179 (N_18179,N_12497,N_12890);
xor U18180 (N_18180,N_11010,N_14880);
and U18181 (N_18181,N_10511,N_12080);
nand U18182 (N_18182,N_14239,N_12864);
nand U18183 (N_18183,N_14557,N_14752);
nor U18184 (N_18184,N_10493,N_14021);
nor U18185 (N_18185,N_10929,N_12450);
and U18186 (N_18186,N_13061,N_14829);
xnor U18187 (N_18187,N_13782,N_10718);
xor U18188 (N_18188,N_13286,N_14082);
nor U18189 (N_18189,N_11100,N_10080);
and U18190 (N_18190,N_12926,N_13917);
nand U18191 (N_18191,N_12262,N_10417);
xor U18192 (N_18192,N_11354,N_13317);
xor U18193 (N_18193,N_13312,N_12276);
nand U18194 (N_18194,N_10006,N_10259);
nor U18195 (N_18195,N_10336,N_10408);
nand U18196 (N_18196,N_12286,N_10590);
and U18197 (N_18197,N_12877,N_12263);
xnor U18198 (N_18198,N_11523,N_14795);
nor U18199 (N_18199,N_14033,N_14049);
and U18200 (N_18200,N_12355,N_13179);
or U18201 (N_18201,N_12802,N_14830);
nor U18202 (N_18202,N_12043,N_11569);
and U18203 (N_18203,N_14921,N_10785);
and U18204 (N_18204,N_10254,N_12847);
and U18205 (N_18205,N_13037,N_10985);
xor U18206 (N_18206,N_13877,N_11648);
xor U18207 (N_18207,N_13527,N_13781);
or U18208 (N_18208,N_10474,N_12352);
nand U18209 (N_18209,N_13882,N_13628);
xnor U18210 (N_18210,N_10131,N_10893);
xnor U18211 (N_18211,N_10621,N_10618);
xnor U18212 (N_18212,N_10016,N_10401);
nand U18213 (N_18213,N_13692,N_14630);
xnor U18214 (N_18214,N_12294,N_11731);
xnor U18215 (N_18215,N_11319,N_12137);
or U18216 (N_18216,N_14466,N_14177);
xor U18217 (N_18217,N_12950,N_12129);
nand U18218 (N_18218,N_10477,N_14687);
and U18219 (N_18219,N_12077,N_13102);
nand U18220 (N_18220,N_13425,N_13444);
or U18221 (N_18221,N_11968,N_14527);
or U18222 (N_18222,N_10176,N_12504);
and U18223 (N_18223,N_11621,N_13836);
nor U18224 (N_18224,N_11467,N_13530);
xnor U18225 (N_18225,N_14934,N_13557);
xor U18226 (N_18226,N_14817,N_10584);
xnor U18227 (N_18227,N_14389,N_13330);
and U18228 (N_18228,N_14242,N_12332);
and U18229 (N_18229,N_12819,N_10922);
and U18230 (N_18230,N_11082,N_13061);
or U18231 (N_18231,N_12329,N_10203);
and U18232 (N_18232,N_12261,N_12446);
nor U18233 (N_18233,N_12535,N_11331);
nor U18234 (N_18234,N_10021,N_13036);
nor U18235 (N_18235,N_13898,N_10441);
and U18236 (N_18236,N_12410,N_13263);
and U18237 (N_18237,N_11788,N_13463);
or U18238 (N_18238,N_11003,N_14359);
xnor U18239 (N_18239,N_12205,N_13668);
nand U18240 (N_18240,N_10874,N_10488);
nand U18241 (N_18241,N_12655,N_10113);
nand U18242 (N_18242,N_14495,N_12606);
nor U18243 (N_18243,N_14176,N_13881);
nand U18244 (N_18244,N_13550,N_14964);
or U18245 (N_18245,N_13715,N_13826);
and U18246 (N_18246,N_14987,N_10167);
nor U18247 (N_18247,N_12775,N_13793);
or U18248 (N_18248,N_13629,N_13252);
nand U18249 (N_18249,N_14002,N_14485);
xor U18250 (N_18250,N_13731,N_13185);
xnor U18251 (N_18251,N_13852,N_14123);
nor U18252 (N_18252,N_14789,N_14731);
xor U18253 (N_18253,N_10071,N_11669);
nor U18254 (N_18254,N_11090,N_14324);
xor U18255 (N_18255,N_12503,N_13703);
or U18256 (N_18256,N_11569,N_11338);
xor U18257 (N_18257,N_14076,N_13585);
xnor U18258 (N_18258,N_13164,N_14480);
or U18259 (N_18259,N_11809,N_14217);
nand U18260 (N_18260,N_10660,N_12996);
xnor U18261 (N_18261,N_10337,N_14558);
or U18262 (N_18262,N_14204,N_10729);
nand U18263 (N_18263,N_14911,N_11504);
or U18264 (N_18264,N_14664,N_13961);
nor U18265 (N_18265,N_12699,N_14275);
nor U18266 (N_18266,N_11960,N_10939);
or U18267 (N_18267,N_13867,N_10073);
xor U18268 (N_18268,N_13264,N_13025);
xnor U18269 (N_18269,N_14752,N_12931);
nor U18270 (N_18270,N_14432,N_13909);
nand U18271 (N_18271,N_12755,N_10146);
xor U18272 (N_18272,N_14263,N_14622);
nand U18273 (N_18273,N_14603,N_10686);
nand U18274 (N_18274,N_12238,N_11119);
xor U18275 (N_18275,N_11219,N_13415);
or U18276 (N_18276,N_14614,N_13396);
xor U18277 (N_18277,N_10335,N_10539);
nor U18278 (N_18278,N_12869,N_11417);
and U18279 (N_18279,N_14214,N_12703);
xor U18280 (N_18280,N_14294,N_12249);
xor U18281 (N_18281,N_10195,N_11832);
and U18282 (N_18282,N_13972,N_11768);
nand U18283 (N_18283,N_11514,N_12918);
xnor U18284 (N_18284,N_10535,N_10976);
nor U18285 (N_18285,N_12871,N_13983);
nand U18286 (N_18286,N_13972,N_13902);
nand U18287 (N_18287,N_13804,N_12720);
or U18288 (N_18288,N_12457,N_14909);
xnor U18289 (N_18289,N_10311,N_14343);
or U18290 (N_18290,N_14975,N_13336);
xor U18291 (N_18291,N_10244,N_10565);
nor U18292 (N_18292,N_10465,N_14110);
nand U18293 (N_18293,N_13451,N_14431);
xor U18294 (N_18294,N_13924,N_14460);
and U18295 (N_18295,N_10367,N_13159);
and U18296 (N_18296,N_11869,N_11143);
and U18297 (N_18297,N_10588,N_12342);
nor U18298 (N_18298,N_11964,N_13518);
and U18299 (N_18299,N_12801,N_14061);
or U18300 (N_18300,N_13213,N_13206);
and U18301 (N_18301,N_12968,N_11846);
or U18302 (N_18302,N_14648,N_10150);
nor U18303 (N_18303,N_12973,N_10009);
xor U18304 (N_18304,N_11933,N_12235);
nor U18305 (N_18305,N_13340,N_14138);
nor U18306 (N_18306,N_11428,N_11757);
or U18307 (N_18307,N_13022,N_14767);
nor U18308 (N_18308,N_11770,N_12063);
and U18309 (N_18309,N_10667,N_10854);
nand U18310 (N_18310,N_13745,N_14596);
and U18311 (N_18311,N_12322,N_13612);
nor U18312 (N_18312,N_10838,N_10707);
or U18313 (N_18313,N_12502,N_14764);
and U18314 (N_18314,N_14888,N_10319);
or U18315 (N_18315,N_14748,N_14880);
or U18316 (N_18316,N_12530,N_10198);
nor U18317 (N_18317,N_14884,N_14283);
nor U18318 (N_18318,N_14626,N_12166);
xnor U18319 (N_18319,N_13428,N_12135);
and U18320 (N_18320,N_13300,N_14509);
or U18321 (N_18321,N_10489,N_14512);
and U18322 (N_18322,N_11490,N_14677);
xnor U18323 (N_18323,N_11168,N_12399);
and U18324 (N_18324,N_11978,N_14915);
xnor U18325 (N_18325,N_11814,N_11772);
nor U18326 (N_18326,N_13961,N_13262);
and U18327 (N_18327,N_10510,N_12901);
and U18328 (N_18328,N_10110,N_11947);
or U18329 (N_18329,N_13026,N_10994);
nand U18330 (N_18330,N_13019,N_10132);
nor U18331 (N_18331,N_12755,N_13069);
and U18332 (N_18332,N_10323,N_11809);
nand U18333 (N_18333,N_13244,N_13600);
xor U18334 (N_18334,N_11526,N_12068);
and U18335 (N_18335,N_11259,N_12991);
nand U18336 (N_18336,N_12014,N_13762);
or U18337 (N_18337,N_13862,N_14509);
and U18338 (N_18338,N_14623,N_13365);
nor U18339 (N_18339,N_10505,N_11766);
and U18340 (N_18340,N_10966,N_10340);
nand U18341 (N_18341,N_14225,N_10908);
nor U18342 (N_18342,N_10642,N_13876);
or U18343 (N_18343,N_12286,N_13383);
or U18344 (N_18344,N_11596,N_11723);
and U18345 (N_18345,N_11809,N_11379);
nand U18346 (N_18346,N_11432,N_10820);
or U18347 (N_18347,N_10431,N_10667);
and U18348 (N_18348,N_14756,N_11119);
nor U18349 (N_18349,N_10190,N_13915);
or U18350 (N_18350,N_12646,N_14411);
and U18351 (N_18351,N_11799,N_13499);
nand U18352 (N_18352,N_14315,N_14967);
and U18353 (N_18353,N_10912,N_12804);
and U18354 (N_18354,N_10990,N_13349);
nand U18355 (N_18355,N_12490,N_11974);
nand U18356 (N_18356,N_12925,N_10174);
or U18357 (N_18357,N_14656,N_14351);
xnor U18358 (N_18358,N_13499,N_11890);
nand U18359 (N_18359,N_13117,N_11600);
nand U18360 (N_18360,N_11844,N_12054);
nor U18361 (N_18361,N_13605,N_14348);
nand U18362 (N_18362,N_11882,N_13274);
nand U18363 (N_18363,N_12648,N_13489);
nand U18364 (N_18364,N_12085,N_13816);
and U18365 (N_18365,N_11227,N_11298);
or U18366 (N_18366,N_11972,N_10768);
nand U18367 (N_18367,N_11259,N_11155);
nand U18368 (N_18368,N_11970,N_13952);
and U18369 (N_18369,N_13932,N_11620);
nand U18370 (N_18370,N_10493,N_13481);
nand U18371 (N_18371,N_10374,N_14618);
xnor U18372 (N_18372,N_14982,N_14472);
xnor U18373 (N_18373,N_14058,N_12765);
nor U18374 (N_18374,N_13274,N_12933);
nor U18375 (N_18375,N_14557,N_12134);
xnor U18376 (N_18376,N_10699,N_11933);
xnor U18377 (N_18377,N_10091,N_14451);
and U18378 (N_18378,N_13889,N_10114);
and U18379 (N_18379,N_12922,N_12733);
or U18380 (N_18380,N_10914,N_12693);
and U18381 (N_18381,N_13512,N_10308);
nor U18382 (N_18382,N_13603,N_14385);
or U18383 (N_18383,N_12221,N_11606);
and U18384 (N_18384,N_11655,N_10250);
nor U18385 (N_18385,N_12552,N_13215);
nand U18386 (N_18386,N_10684,N_10670);
nand U18387 (N_18387,N_12887,N_10705);
or U18388 (N_18388,N_10560,N_10774);
and U18389 (N_18389,N_12263,N_10964);
nor U18390 (N_18390,N_10240,N_12880);
nor U18391 (N_18391,N_14899,N_10951);
nand U18392 (N_18392,N_14810,N_14151);
nor U18393 (N_18393,N_11780,N_14289);
or U18394 (N_18394,N_12280,N_13518);
or U18395 (N_18395,N_11802,N_10653);
or U18396 (N_18396,N_12123,N_10223);
or U18397 (N_18397,N_11150,N_11118);
and U18398 (N_18398,N_11085,N_10639);
nand U18399 (N_18399,N_13966,N_11828);
and U18400 (N_18400,N_14972,N_13804);
nor U18401 (N_18401,N_14820,N_13090);
and U18402 (N_18402,N_10772,N_13526);
or U18403 (N_18403,N_10232,N_13076);
nor U18404 (N_18404,N_10253,N_14743);
nor U18405 (N_18405,N_13920,N_11160);
xor U18406 (N_18406,N_10406,N_12358);
and U18407 (N_18407,N_10185,N_13839);
or U18408 (N_18408,N_11863,N_13209);
and U18409 (N_18409,N_10915,N_10282);
or U18410 (N_18410,N_11484,N_13679);
nor U18411 (N_18411,N_13556,N_10694);
xor U18412 (N_18412,N_14128,N_13864);
xnor U18413 (N_18413,N_12366,N_13364);
nand U18414 (N_18414,N_14697,N_10140);
nand U18415 (N_18415,N_12012,N_14678);
nand U18416 (N_18416,N_11211,N_13194);
and U18417 (N_18417,N_10898,N_12012);
nand U18418 (N_18418,N_11171,N_10217);
and U18419 (N_18419,N_13617,N_12497);
or U18420 (N_18420,N_11761,N_11028);
and U18421 (N_18421,N_12215,N_11607);
nand U18422 (N_18422,N_11938,N_12260);
or U18423 (N_18423,N_10119,N_12926);
nor U18424 (N_18424,N_14458,N_10150);
nor U18425 (N_18425,N_14429,N_12231);
and U18426 (N_18426,N_14042,N_14918);
nor U18427 (N_18427,N_13227,N_10738);
and U18428 (N_18428,N_10569,N_14120);
nor U18429 (N_18429,N_14451,N_10046);
xnor U18430 (N_18430,N_13151,N_13350);
or U18431 (N_18431,N_12737,N_13217);
or U18432 (N_18432,N_11772,N_10084);
and U18433 (N_18433,N_12933,N_13184);
or U18434 (N_18434,N_12822,N_13002);
nor U18435 (N_18435,N_12670,N_12596);
or U18436 (N_18436,N_11315,N_10867);
or U18437 (N_18437,N_13002,N_11510);
or U18438 (N_18438,N_11344,N_12413);
nand U18439 (N_18439,N_11218,N_13723);
or U18440 (N_18440,N_14817,N_12026);
nand U18441 (N_18441,N_14338,N_10182);
or U18442 (N_18442,N_11133,N_11327);
nor U18443 (N_18443,N_10144,N_11695);
nor U18444 (N_18444,N_10932,N_13486);
or U18445 (N_18445,N_13391,N_13052);
nor U18446 (N_18446,N_10990,N_14926);
or U18447 (N_18447,N_14461,N_10135);
nor U18448 (N_18448,N_10467,N_10103);
or U18449 (N_18449,N_14867,N_11614);
xor U18450 (N_18450,N_12433,N_14450);
or U18451 (N_18451,N_14818,N_12643);
nand U18452 (N_18452,N_10550,N_12820);
or U18453 (N_18453,N_10137,N_11440);
nor U18454 (N_18454,N_13845,N_14636);
or U18455 (N_18455,N_12878,N_10485);
and U18456 (N_18456,N_12091,N_11493);
xor U18457 (N_18457,N_12733,N_13041);
or U18458 (N_18458,N_13833,N_12287);
or U18459 (N_18459,N_14326,N_13870);
xnor U18460 (N_18460,N_10157,N_13364);
nor U18461 (N_18461,N_10836,N_12802);
or U18462 (N_18462,N_10605,N_10989);
and U18463 (N_18463,N_10643,N_12986);
or U18464 (N_18464,N_13572,N_12048);
nand U18465 (N_18465,N_13074,N_11332);
xor U18466 (N_18466,N_10432,N_11029);
nand U18467 (N_18467,N_11753,N_12380);
nand U18468 (N_18468,N_14397,N_12522);
or U18469 (N_18469,N_13419,N_14617);
nand U18470 (N_18470,N_11225,N_14555);
nand U18471 (N_18471,N_11409,N_12101);
xor U18472 (N_18472,N_10966,N_11001);
or U18473 (N_18473,N_10689,N_13600);
xnor U18474 (N_18474,N_14351,N_14517);
nor U18475 (N_18475,N_12831,N_10074);
and U18476 (N_18476,N_10220,N_11202);
nor U18477 (N_18477,N_11026,N_12225);
nand U18478 (N_18478,N_14153,N_11183);
nor U18479 (N_18479,N_10150,N_11332);
and U18480 (N_18480,N_12542,N_11009);
nor U18481 (N_18481,N_10238,N_12664);
or U18482 (N_18482,N_14760,N_10356);
or U18483 (N_18483,N_11544,N_11381);
nand U18484 (N_18484,N_13206,N_11752);
and U18485 (N_18485,N_10520,N_10538);
nand U18486 (N_18486,N_11286,N_11104);
nor U18487 (N_18487,N_11015,N_10879);
nand U18488 (N_18488,N_14652,N_11638);
xnor U18489 (N_18489,N_13062,N_14175);
nor U18490 (N_18490,N_11874,N_10537);
nand U18491 (N_18491,N_11933,N_10995);
nor U18492 (N_18492,N_13635,N_12459);
nor U18493 (N_18493,N_11738,N_10639);
and U18494 (N_18494,N_10948,N_14458);
nor U18495 (N_18495,N_14469,N_14856);
and U18496 (N_18496,N_12442,N_12566);
xnor U18497 (N_18497,N_12138,N_10403);
and U18498 (N_18498,N_12061,N_11329);
nor U18499 (N_18499,N_12808,N_10629);
nand U18500 (N_18500,N_10804,N_13708);
or U18501 (N_18501,N_10871,N_14736);
nor U18502 (N_18502,N_12288,N_13719);
and U18503 (N_18503,N_12567,N_10736);
and U18504 (N_18504,N_12268,N_10724);
xor U18505 (N_18505,N_10546,N_14179);
xor U18506 (N_18506,N_11085,N_13286);
nand U18507 (N_18507,N_11992,N_12515);
nand U18508 (N_18508,N_11114,N_10299);
nand U18509 (N_18509,N_13452,N_10253);
or U18510 (N_18510,N_10507,N_12126);
nor U18511 (N_18511,N_11823,N_11161);
xnor U18512 (N_18512,N_12370,N_12768);
nand U18513 (N_18513,N_10175,N_14026);
nand U18514 (N_18514,N_12575,N_13592);
and U18515 (N_18515,N_10479,N_13727);
nand U18516 (N_18516,N_10588,N_10715);
nand U18517 (N_18517,N_11941,N_10970);
nand U18518 (N_18518,N_13113,N_13449);
nor U18519 (N_18519,N_10232,N_10242);
or U18520 (N_18520,N_12717,N_12076);
xor U18521 (N_18521,N_10563,N_13333);
or U18522 (N_18522,N_11439,N_14362);
or U18523 (N_18523,N_13387,N_12541);
xnor U18524 (N_18524,N_13595,N_14609);
nor U18525 (N_18525,N_14049,N_10857);
and U18526 (N_18526,N_11395,N_13399);
or U18527 (N_18527,N_11975,N_14783);
and U18528 (N_18528,N_12468,N_13232);
or U18529 (N_18529,N_11177,N_11593);
or U18530 (N_18530,N_12753,N_14811);
xnor U18531 (N_18531,N_10354,N_13449);
and U18532 (N_18532,N_12010,N_13308);
nand U18533 (N_18533,N_12431,N_12101);
or U18534 (N_18534,N_10386,N_13026);
or U18535 (N_18535,N_12047,N_11349);
or U18536 (N_18536,N_13031,N_14432);
or U18537 (N_18537,N_13429,N_11678);
and U18538 (N_18538,N_14961,N_11133);
or U18539 (N_18539,N_14518,N_13550);
and U18540 (N_18540,N_10232,N_11873);
nand U18541 (N_18541,N_13691,N_11481);
or U18542 (N_18542,N_12766,N_13451);
and U18543 (N_18543,N_11677,N_14364);
xor U18544 (N_18544,N_14470,N_14806);
and U18545 (N_18545,N_12594,N_10173);
xnor U18546 (N_18546,N_14118,N_12457);
or U18547 (N_18547,N_11635,N_12947);
and U18548 (N_18548,N_13857,N_12195);
nor U18549 (N_18549,N_10196,N_11255);
nand U18550 (N_18550,N_12086,N_14888);
nand U18551 (N_18551,N_10458,N_13759);
or U18552 (N_18552,N_13115,N_13291);
xor U18553 (N_18553,N_12192,N_14052);
nand U18554 (N_18554,N_13185,N_11765);
nand U18555 (N_18555,N_12125,N_11538);
and U18556 (N_18556,N_10086,N_13558);
xnor U18557 (N_18557,N_10832,N_13560);
and U18558 (N_18558,N_11699,N_13583);
and U18559 (N_18559,N_10835,N_14960);
xnor U18560 (N_18560,N_11303,N_14908);
nand U18561 (N_18561,N_14342,N_11149);
nand U18562 (N_18562,N_13239,N_14214);
nand U18563 (N_18563,N_11446,N_12085);
nand U18564 (N_18564,N_11912,N_13970);
or U18565 (N_18565,N_10749,N_14417);
nand U18566 (N_18566,N_11786,N_12830);
nor U18567 (N_18567,N_14572,N_13117);
or U18568 (N_18568,N_13748,N_10671);
nand U18569 (N_18569,N_12495,N_10869);
nor U18570 (N_18570,N_11398,N_13765);
or U18571 (N_18571,N_13702,N_14536);
nand U18572 (N_18572,N_13436,N_12960);
xor U18573 (N_18573,N_12752,N_11692);
xnor U18574 (N_18574,N_13947,N_12478);
nor U18575 (N_18575,N_13951,N_14158);
and U18576 (N_18576,N_10597,N_10394);
or U18577 (N_18577,N_10048,N_14231);
nand U18578 (N_18578,N_10846,N_14660);
and U18579 (N_18579,N_11605,N_12440);
nor U18580 (N_18580,N_11472,N_10622);
xor U18581 (N_18581,N_10239,N_13129);
and U18582 (N_18582,N_12934,N_13535);
nor U18583 (N_18583,N_13103,N_12372);
nand U18584 (N_18584,N_13229,N_14765);
or U18585 (N_18585,N_10355,N_11170);
or U18586 (N_18586,N_12887,N_10723);
nor U18587 (N_18587,N_13531,N_10643);
nand U18588 (N_18588,N_11558,N_11996);
and U18589 (N_18589,N_14867,N_11387);
nor U18590 (N_18590,N_14719,N_10072);
nor U18591 (N_18591,N_10174,N_13528);
and U18592 (N_18592,N_10573,N_12001);
and U18593 (N_18593,N_14813,N_13860);
and U18594 (N_18594,N_10644,N_10801);
nand U18595 (N_18595,N_11271,N_10121);
and U18596 (N_18596,N_12875,N_12186);
nor U18597 (N_18597,N_12609,N_13434);
and U18598 (N_18598,N_14385,N_11754);
nand U18599 (N_18599,N_13034,N_10134);
xnor U18600 (N_18600,N_10366,N_13424);
xnor U18601 (N_18601,N_10920,N_11881);
and U18602 (N_18602,N_11325,N_10826);
nand U18603 (N_18603,N_10604,N_13254);
nand U18604 (N_18604,N_11618,N_12449);
nand U18605 (N_18605,N_13604,N_10795);
or U18606 (N_18606,N_12651,N_12429);
nand U18607 (N_18607,N_12100,N_12418);
xor U18608 (N_18608,N_12640,N_10879);
and U18609 (N_18609,N_11648,N_11121);
or U18610 (N_18610,N_13096,N_14678);
nor U18611 (N_18611,N_10856,N_10032);
and U18612 (N_18612,N_13060,N_14743);
xnor U18613 (N_18613,N_10966,N_12288);
nand U18614 (N_18614,N_10867,N_11888);
xnor U18615 (N_18615,N_14227,N_14666);
or U18616 (N_18616,N_14252,N_11123);
nand U18617 (N_18617,N_14018,N_14790);
or U18618 (N_18618,N_11558,N_12692);
nor U18619 (N_18619,N_13005,N_12905);
nor U18620 (N_18620,N_11728,N_12673);
xnor U18621 (N_18621,N_14446,N_14986);
xor U18622 (N_18622,N_11994,N_10827);
and U18623 (N_18623,N_14250,N_11713);
nand U18624 (N_18624,N_10238,N_12010);
nor U18625 (N_18625,N_13038,N_12516);
nor U18626 (N_18626,N_11702,N_12066);
nor U18627 (N_18627,N_11523,N_11107);
or U18628 (N_18628,N_10488,N_11810);
xor U18629 (N_18629,N_11602,N_11819);
or U18630 (N_18630,N_11490,N_12956);
nand U18631 (N_18631,N_10555,N_13497);
nor U18632 (N_18632,N_10625,N_10646);
nor U18633 (N_18633,N_14136,N_11076);
or U18634 (N_18634,N_10289,N_13160);
nor U18635 (N_18635,N_10384,N_12555);
and U18636 (N_18636,N_10197,N_11835);
xnor U18637 (N_18637,N_12317,N_11707);
or U18638 (N_18638,N_11220,N_10727);
nor U18639 (N_18639,N_13519,N_11078);
nand U18640 (N_18640,N_13124,N_10246);
or U18641 (N_18641,N_13798,N_13368);
nor U18642 (N_18642,N_14422,N_14953);
nor U18643 (N_18643,N_13476,N_14963);
or U18644 (N_18644,N_14255,N_11718);
nor U18645 (N_18645,N_13528,N_12405);
xor U18646 (N_18646,N_11704,N_13720);
or U18647 (N_18647,N_14013,N_11841);
nor U18648 (N_18648,N_10632,N_12938);
xor U18649 (N_18649,N_10108,N_11431);
nor U18650 (N_18650,N_13482,N_14947);
and U18651 (N_18651,N_10960,N_13181);
xor U18652 (N_18652,N_13812,N_11066);
nor U18653 (N_18653,N_10813,N_11687);
xor U18654 (N_18654,N_10159,N_11899);
and U18655 (N_18655,N_11979,N_12313);
or U18656 (N_18656,N_13028,N_13426);
xor U18657 (N_18657,N_14868,N_10347);
and U18658 (N_18658,N_11567,N_10143);
xnor U18659 (N_18659,N_11041,N_11874);
nor U18660 (N_18660,N_13027,N_14264);
or U18661 (N_18661,N_10163,N_11807);
nand U18662 (N_18662,N_10050,N_11684);
nand U18663 (N_18663,N_14261,N_13332);
nor U18664 (N_18664,N_11556,N_11840);
xnor U18665 (N_18665,N_12617,N_12929);
nor U18666 (N_18666,N_14238,N_13587);
nand U18667 (N_18667,N_13358,N_14875);
xor U18668 (N_18668,N_14403,N_13526);
xnor U18669 (N_18669,N_10162,N_14132);
or U18670 (N_18670,N_12455,N_12003);
or U18671 (N_18671,N_13484,N_13840);
nand U18672 (N_18672,N_12724,N_12147);
nand U18673 (N_18673,N_12654,N_11527);
nand U18674 (N_18674,N_11348,N_14195);
nand U18675 (N_18675,N_13984,N_11425);
xnor U18676 (N_18676,N_10173,N_12476);
and U18677 (N_18677,N_11824,N_10157);
nand U18678 (N_18678,N_10539,N_11601);
or U18679 (N_18679,N_12503,N_14789);
or U18680 (N_18680,N_11496,N_11695);
xnor U18681 (N_18681,N_11217,N_14691);
nor U18682 (N_18682,N_14301,N_12124);
or U18683 (N_18683,N_12925,N_14957);
nor U18684 (N_18684,N_13433,N_12205);
and U18685 (N_18685,N_13294,N_14880);
xor U18686 (N_18686,N_10936,N_14158);
nand U18687 (N_18687,N_10465,N_14784);
nand U18688 (N_18688,N_14517,N_14623);
or U18689 (N_18689,N_12686,N_11692);
or U18690 (N_18690,N_13674,N_12878);
nor U18691 (N_18691,N_14400,N_13182);
xnor U18692 (N_18692,N_13433,N_13764);
nand U18693 (N_18693,N_14640,N_13814);
or U18694 (N_18694,N_13115,N_13434);
nor U18695 (N_18695,N_11743,N_14792);
xor U18696 (N_18696,N_12825,N_14014);
xor U18697 (N_18697,N_10530,N_11020);
or U18698 (N_18698,N_12146,N_12771);
nor U18699 (N_18699,N_13404,N_10586);
nand U18700 (N_18700,N_13684,N_14628);
nor U18701 (N_18701,N_13016,N_10894);
nand U18702 (N_18702,N_13636,N_13093);
or U18703 (N_18703,N_10083,N_12825);
xnor U18704 (N_18704,N_14255,N_12387);
nand U18705 (N_18705,N_11518,N_14313);
nor U18706 (N_18706,N_14901,N_10018);
and U18707 (N_18707,N_12599,N_11485);
xor U18708 (N_18708,N_10116,N_10814);
nor U18709 (N_18709,N_11021,N_11323);
and U18710 (N_18710,N_10199,N_12201);
nor U18711 (N_18711,N_12738,N_11792);
xnor U18712 (N_18712,N_11186,N_10949);
and U18713 (N_18713,N_14282,N_14177);
or U18714 (N_18714,N_11398,N_13510);
nor U18715 (N_18715,N_12286,N_13888);
nand U18716 (N_18716,N_13414,N_13434);
nor U18717 (N_18717,N_13134,N_14395);
or U18718 (N_18718,N_14455,N_10444);
nor U18719 (N_18719,N_13954,N_11600);
xor U18720 (N_18720,N_12499,N_14298);
and U18721 (N_18721,N_12208,N_13753);
nand U18722 (N_18722,N_11639,N_10173);
and U18723 (N_18723,N_11011,N_10067);
xor U18724 (N_18724,N_10148,N_14573);
or U18725 (N_18725,N_11576,N_11535);
or U18726 (N_18726,N_11548,N_14574);
xor U18727 (N_18727,N_14971,N_14849);
xor U18728 (N_18728,N_11215,N_14721);
or U18729 (N_18729,N_12047,N_13955);
nor U18730 (N_18730,N_13817,N_13366);
nand U18731 (N_18731,N_13171,N_12126);
nand U18732 (N_18732,N_12294,N_12359);
nand U18733 (N_18733,N_11423,N_14243);
and U18734 (N_18734,N_13137,N_14913);
nor U18735 (N_18735,N_14058,N_10692);
or U18736 (N_18736,N_13185,N_13747);
and U18737 (N_18737,N_12755,N_13283);
or U18738 (N_18738,N_11104,N_12784);
nor U18739 (N_18739,N_10917,N_12627);
xnor U18740 (N_18740,N_10069,N_10941);
nor U18741 (N_18741,N_10977,N_13200);
nor U18742 (N_18742,N_12810,N_13927);
and U18743 (N_18743,N_11402,N_13169);
and U18744 (N_18744,N_14166,N_11661);
and U18745 (N_18745,N_10884,N_14879);
nor U18746 (N_18746,N_12650,N_10132);
nor U18747 (N_18747,N_10166,N_13555);
and U18748 (N_18748,N_10422,N_14633);
xor U18749 (N_18749,N_13962,N_12213);
or U18750 (N_18750,N_13168,N_11155);
xor U18751 (N_18751,N_10821,N_10914);
nand U18752 (N_18752,N_13508,N_10615);
nand U18753 (N_18753,N_12102,N_14696);
and U18754 (N_18754,N_11341,N_14851);
and U18755 (N_18755,N_13232,N_12703);
xnor U18756 (N_18756,N_13826,N_14274);
nand U18757 (N_18757,N_14305,N_10320);
nand U18758 (N_18758,N_13011,N_12662);
or U18759 (N_18759,N_13551,N_14361);
and U18760 (N_18760,N_10773,N_10705);
xor U18761 (N_18761,N_10904,N_12882);
or U18762 (N_18762,N_14834,N_13463);
nor U18763 (N_18763,N_10019,N_10226);
nor U18764 (N_18764,N_11244,N_10251);
nor U18765 (N_18765,N_12647,N_13320);
or U18766 (N_18766,N_14249,N_10118);
xnor U18767 (N_18767,N_10957,N_11064);
or U18768 (N_18768,N_11180,N_12933);
nor U18769 (N_18769,N_12307,N_11169);
and U18770 (N_18770,N_10488,N_14896);
nor U18771 (N_18771,N_10205,N_13088);
or U18772 (N_18772,N_11899,N_12800);
xor U18773 (N_18773,N_10290,N_13430);
nand U18774 (N_18774,N_11991,N_11612);
or U18775 (N_18775,N_13672,N_10368);
or U18776 (N_18776,N_10965,N_14803);
or U18777 (N_18777,N_12355,N_12457);
and U18778 (N_18778,N_13590,N_11911);
and U18779 (N_18779,N_11504,N_14913);
xnor U18780 (N_18780,N_10482,N_14861);
xnor U18781 (N_18781,N_10934,N_13812);
xnor U18782 (N_18782,N_12725,N_11722);
xor U18783 (N_18783,N_10760,N_13321);
xor U18784 (N_18784,N_14044,N_10391);
xor U18785 (N_18785,N_14418,N_13412);
nand U18786 (N_18786,N_14350,N_14147);
and U18787 (N_18787,N_11710,N_11001);
xor U18788 (N_18788,N_10641,N_10136);
xnor U18789 (N_18789,N_13338,N_13006);
and U18790 (N_18790,N_11443,N_11136);
xor U18791 (N_18791,N_13698,N_14617);
nand U18792 (N_18792,N_12250,N_10072);
or U18793 (N_18793,N_12470,N_14640);
and U18794 (N_18794,N_11175,N_13264);
and U18795 (N_18795,N_10004,N_11988);
nor U18796 (N_18796,N_13722,N_12231);
or U18797 (N_18797,N_11484,N_10602);
or U18798 (N_18798,N_10216,N_11671);
or U18799 (N_18799,N_13016,N_10724);
and U18800 (N_18800,N_12388,N_13739);
and U18801 (N_18801,N_12243,N_11510);
xnor U18802 (N_18802,N_10316,N_14547);
and U18803 (N_18803,N_10772,N_12143);
or U18804 (N_18804,N_12222,N_10037);
and U18805 (N_18805,N_11611,N_10655);
and U18806 (N_18806,N_10653,N_14399);
or U18807 (N_18807,N_12556,N_12481);
nor U18808 (N_18808,N_11815,N_14338);
and U18809 (N_18809,N_13017,N_14467);
or U18810 (N_18810,N_10605,N_12857);
or U18811 (N_18811,N_11180,N_11416);
nand U18812 (N_18812,N_10499,N_13715);
nand U18813 (N_18813,N_11550,N_11754);
nand U18814 (N_18814,N_10617,N_11346);
and U18815 (N_18815,N_14824,N_10330);
nand U18816 (N_18816,N_10765,N_10512);
nor U18817 (N_18817,N_14500,N_13478);
nor U18818 (N_18818,N_14771,N_12016);
nor U18819 (N_18819,N_11778,N_10556);
xnor U18820 (N_18820,N_10332,N_14811);
nand U18821 (N_18821,N_13994,N_11176);
nand U18822 (N_18822,N_13497,N_12939);
or U18823 (N_18823,N_11378,N_13961);
xor U18824 (N_18824,N_11792,N_13994);
xnor U18825 (N_18825,N_14746,N_12615);
and U18826 (N_18826,N_10964,N_12810);
xnor U18827 (N_18827,N_12249,N_11258);
nand U18828 (N_18828,N_12341,N_10300);
xnor U18829 (N_18829,N_13415,N_13229);
nor U18830 (N_18830,N_11761,N_10916);
or U18831 (N_18831,N_14846,N_14019);
and U18832 (N_18832,N_13549,N_11651);
nand U18833 (N_18833,N_11236,N_13661);
nor U18834 (N_18834,N_11652,N_11831);
nand U18835 (N_18835,N_12699,N_11675);
nor U18836 (N_18836,N_14925,N_11234);
and U18837 (N_18837,N_13123,N_10960);
and U18838 (N_18838,N_14711,N_14407);
and U18839 (N_18839,N_12805,N_11857);
or U18840 (N_18840,N_13483,N_12999);
and U18841 (N_18841,N_13206,N_13998);
nand U18842 (N_18842,N_14830,N_11995);
nand U18843 (N_18843,N_14244,N_12177);
xnor U18844 (N_18844,N_13053,N_13874);
nor U18845 (N_18845,N_13050,N_14361);
xnor U18846 (N_18846,N_11431,N_14839);
xor U18847 (N_18847,N_14249,N_12574);
and U18848 (N_18848,N_12779,N_13922);
nand U18849 (N_18849,N_14386,N_12728);
nor U18850 (N_18850,N_10336,N_11728);
and U18851 (N_18851,N_13581,N_12912);
nand U18852 (N_18852,N_11677,N_14777);
nor U18853 (N_18853,N_13331,N_11712);
nor U18854 (N_18854,N_12779,N_10962);
nand U18855 (N_18855,N_14113,N_11018);
and U18856 (N_18856,N_14170,N_10138);
or U18857 (N_18857,N_10424,N_13542);
xor U18858 (N_18858,N_13149,N_10383);
or U18859 (N_18859,N_12635,N_10787);
or U18860 (N_18860,N_12221,N_12054);
nand U18861 (N_18861,N_10586,N_12117);
nor U18862 (N_18862,N_14326,N_12306);
xor U18863 (N_18863,N_13452,N_14498);
and U18864 (N_18864,N_11614,N_10522);
or U18865 (N_18865,N_14406,N_12937);
and U18866 (N_18866,N_10660,N_13084);
nand U18867 (N_18867,N_12214,N_11403);
nor U18868 (N_18868,N_13833,N_11023);
or U18869 (N_18869,N_10685,N_10940);
and U18870 (N_18870,N_11531,N_14574);
nand U18871 (N_18871,N_11911,N_13017);
and U18872 (N_18872,N_11620,N_10428);
xnor U18873 (N_18873,N_13900,N_14217);
and U18874 (N_18874,N_14095,N_10556);
or U18875 (N_18875,N_10535,N_12951);
or U18876 (N_18876,N_12344,N_14252);
nand U18877 (N_18877,N_13379,N_10686);
or U18878 (N_18878,N_12715,N_11787);
or U18879 (N_18879,N_13708,N_11552);
and U18880 (N_18880,N_10638,N_14729);
nor U18881 (N_18881,N_11506,N_11444);
and U18882 (N_18882,N_10710,N_10553);
nor U18883 (N_18883,N_10122,N_11451);
nor U18884 (N_18884,N_10819,N_14687);
xnor U18885 (N_18885,N_13533,N_13049);
nor U18886 (N_18886,N_11893,N_11913);
nor U18887 (N_18887,N_11092,N_10530);
nor U18888 (N_18888,N_14139,N_11126);
xor U18889 (N_18889,N_13904,N_14717);
and U18890 (N_18890,N_13919,N_11347);
nand U18891 (N_18891,N_14383,N_13071);
nor U18892 (N_18892,N_12938,N_12212);
nand U18893 (N_18893,N_12701,N_12652);
nand U18894 (N_18894,N_10446,N_13444);
nor U18895 (N_18895,N_14665,N_13860);
or U18896 (N_18896,N_14387,N_10280);
nand U18897 (N_18897,N_10657,N_13983);
or U18898 (N_18898,N_10683,N_10273);
nor U18899 (N_18899,N_13829,N_10397);
and U18900 (N_18900,N_11045,N_14262);
nor U18901 (N_18901,N_12019,N_12344);
nand U18902 (N_18902,N_11681,N_11626);
nor U18903 (N_18903,N_12484,N_13408);
nor U18904 (N_18904,N_10881,N_14152);
nor U18905 (N_18905,N_11137,N_12805);
and U18906 (N_18906,N_13200,N_14369);
xor U18907 (N_18907,N_13948,N_13357);
nand U18908 (N_18908,N_11552,N_14271);
and U18909 (N_18909,N_14809,N_10851);
xnor U18910 (N_18910,N_12523,N_12109);
nand U18911 (N_18911,N_11457,N_12474);
nor U18912 (N_18912,N_13156,N_12140);
or U18913 (N_18913,N_11178,N_13525);
nand U18914 (N_18914,N_14159,N_10868);
xor U18915 (N_18915,N_10906,N_14810);
nor U18916 (N_18916,N_11452,N_11776);
nor U18917 (N_18917,N_11267,N_14924);
xor U18918 (N_18918,N_12432,N_13859);
and U18919 (N_18919,N_10914,N_13674);
nand U18920 (N_18920,N_12320,N_10964);
xor U18921 (N_18921,N_10111,N_13451);
or U18922 (N_18922,N_12344,N_11061);
and U18923 (N_18923,N_14569,N_13685);
nand U18924 (N_18924,N_12301,N_14083);
nor U18925 (N_18925,N_10817,N_13681);
nand U18926 (N_18926,N_13413,N_12543);
xnor U18927 (N_18927,N_11362,N_10674);
nor U18928 (N_18928,N_14206,N_13719);
and U18929 (N_18929,N_11461,N_10044);
nor U18930 (N_18930,N_14468,N_11830);
nor U18931 (N_18931,N_12870,N_10618);
nand U18932 (N_18932,N_10003,N_13610);
or U18933 (N_18933,N_11149,N_13341);
xor U18934 (N_18934,N_14161,N_10832);
nand U18935 (N_18935,N_12878,N_10736);
nand U18936 (N_18936,N_12702,N_11285);
nor U18937 (N_18937,N_10395,N_12798);
nor U18938 (N_18938,N_11358,N_13841);
or U18939 (N_18939,N_14797,N_11755);
or U18940 (N_18940,N_11373,N_12832);
nand U18941 (N_18941,N_10635,N_12282);
nor U18942 (N_18942,N_12661,N_14477);
and U18943 (N_18943,N_12684,N_11293);
nor U18944 (N_18944,N_11103,N_12661);
nand U18945 (N_18945,N_10383,N_13824);
or U18946 (N_18946,N_13705,N_14166);
xor U18947 (N_18947,N_13261,N_10511);
or U18948 (N_18948,N_10074,N_14029);
or U18949 (N_18949,N_11215,N_11073);
or U18950 (N_18950,N_14005,N_11058);
nand U18951 (N_18951,N_11026,N_10185);
nor U18952 (N_18952,N_13972,N_13755);
or U18953 (N_18953,N_13556,N_14572);
nand U18954 (N_18954,N_12853,N_10797);
xnor U18955 (N_18955,N_14515,N_12279);
xnor U18956 (N_18956,N_12122,N_10286);
or U18957 (N_18957,N_13079,N_14906);
nor U18958 (N_18958,N_11876,N_11488);
nand U18959 (N_18959,N_10655,N_14056);
xnor U18960 (N_18960,N_14734,N_10049);
nand U18961 (N_18961,N_10549,N_13029);
nand U18962 (N_18962,N_11416,N_13800);
and U18963 (N_18963,N_14561,N_14582);
and U18964 (N_18964,N_12195,N_13858);
and U18965 (N_18965,N_14432,N_13413);
and U18966 (N_18966,N_11210,N_10726);
xor U18967 (N_18967,N_13497,N_12410);
xor U18968 (N_18968,N_11292,N_11855);
xnor U18969 (N_18969,N_11927,N_10679);
nand U18970 (N_18970,N_13780,N_12512);
xor U18971 (N_18971,N_13251,N_11313);
or U18972 (N_18972,N_12353,N_10513);
and U18973 (N_18973,N_13331,N_10621);
nor U18974 (N_18974,N_10798,N_12328);
and U18975 (N_18975,N_11768,N_14781);
nand U18976 (N_18976,N_11731,N_13174);
nand U18977 (N_18977,N_13059,N_13202);
nor U18978 (N_18978,N_13338,N_14972);
nand U18979 (N_18979,N_10895,N_11528);
or U18980 (N_18980,N_11653,N_11096);
and U18981 (N_18981,N_10489,N_10156);
nand U18982 (N_18982,N_10856,N_13544);
or U18983 (N_18983,N_10720,N_12577);
nor U18984 (N_18984,N_13523,N_14266);
or U18985 (N_18985,N_11746,N_12836);
or U18986 (N_18986,N_14070,N_10921);
or U18987 (N_18987,N_14378,N_10835);
or U18988 (N_18988,N_13211,N_12564);
nand U18989 (N_18989,N_14644,N_12752);
or U18990 (N_18990,N_12201,N_10019);
nor U18991 (N_18991,N_10600,N_12778);
xnor U18992 (N_18992,N_11440,N_12527);
xnor U18993 (N_18993,N_12857,N_14445);
xnor U18994 (N_18994,N_13992,N_13455);
nand U18995 (N_18995,N_12156,N_12701);
xnor U18996 (N_18996,N_14917,N_11846);
and U18997 (N_18997,N_10396,N_14977);
xor U18998 (N_18998,N_13890,N_13520);
nand U18999 (N_18999,N_10675,N_12287);
or U19000 (N_19000,N_13330,N_12975);
nand U19001 (N_19001,N_12110,N_13588);
nor U19002 (N_19002,N_11143,N_14847);
and U19003 (N_19003,N_10560,N_10922);
nand U19004 (N_19004,N_10714,N_12619);
nor U19005 (N_19005,N_14325,N_10248);
and U19006 (N_19006,N_14998,N_10885);
or U19007 (N_19007,N_13991,N_13868);
xor U19008 (N_19008,N_11842,N_12382);
or U19009 (N_19009,N_11124,N_14294);
nand U19010 (N_19010,N_12371,N_11888);
or U19011 (N_19011,N_10153,N_13394);
and U19012 (N_19012,N_10282,N_13368);
or U19013 (N_19013,N_12107,N_12278);
nand U19014 (N_19014,N_12414,N_14167);
and U19015 (N_19015,N_11176,N_10478);
and U19016 (N_19016,N_14051,N_12083);
nor U19017 (N_19017,N_10197,N_13373);
or U19018 (N_19018,N_14772,N_13247);
and U19019 (N_19019,N_14948,N_11163);
and U19020 (N_19020,N_13630,N_12213);
nand U19021 (N_19021,N_10044,N_12264);
or U19022 (N_19022,N_13327,N_10116);
nand U19023 (N_19023,N_11879,N_13214);
and U19024 (N_19024,N_14053,N_13391);
nor U19025 (N_19025,N_10137,N_13793);
or U19026 (N_19026,N_10015,N_11162);
nor U19027 (N_19027,N_13427,N_10519);
or U19028 (N_19028,N_14161,N_13918);
nor U19029 (N_19029,N_11685,N_14273);
xor U19030 (N_19030,N_13577,N_10947);
and U19031 (N_19031,N_12860,N_10560);
and U19032 (N_19032,N_11862,N_14836);
or U19033 (N_19033,N_13798,N_11688);
xnor U19034 (N_19034,N_11768,N_14536);
nand U19035 (N_19035,N_13058,N_11838);
and U19036 (N_19036,N_11502,N_12230);
xor U19037 (N_19037,N_13628,N_12964);
or U19038 (N_19038,N_12209,N_12213);
nand U19039 (N_19039,N_10018,N_13863);
or U19040 (N_19040,N_14658,N_13509);
or U19041 (N_19041,N_14567,N_14202);
nand U19042 (N_19042,N_10234,N_11380);
nand U19043 (N_19043,N_14668,N_14049);
and U19044 (N_19044,N_10455,N_14500);
or U19045 (N_19045,N_11658,N_11662);
or U19046 (N_19046,N_10719,N_11350);
nand U19047 (N_19047,N_12708,N_13293);
nand U19048 (N_19048,N_11082,N_14068);
and U19049 (N_19049,N_10987,N_14874);
or U19050 (N_19050,N_11584,N_12647);
or U19051 (N_19051,N_14204,N_14218);
nand U19052 (N_19052,N_13663,N_12751);
nand U19053 (N_19053,N_12928,N_14781);
nor U19054 (N_19054,N_10702,N_14446);
xnor U19055 (N_19055,N_11258,N_13751);
and U19056 (N_19056,N_11303,N_13897);
or U19057 (N_19057,N_11119,N_14971);
xor U19058 (N_19058,N_14371,N_14471);
nand U19059 (N_19059,N_10228,N_13279);
and U19060 (N_19060,N_10114,N_11942);
or U19061 (N_19061,N_14421,N_11668);
and U19062 (N_19062,N_12135,N_11956);
nand U19063 (N_19063,N_10370,N_11945);
nor U19064 (N_19064,N_13788,N_11057);
and U19065 (N_19065,N_12820,N_11420);
xor U19066 (N_19066,N_12937,N_14616);
or U19067 (N_19067,N_14128,N_14112);
nand U19068 (N_19068,N_11722,N_14070);
nand U19069 (N_19069,N_12853,N_11102);
and U19070 (N_19070,N_11606,N_13720);
xor U19071 (N_19071,N_11329,N_13912);
xnor U19072 (N_19072,N_11483,N_10938);
xnor U19073 (N_19073,N_12370,N_12512);
nor U19074 (N_19074,N_10779,N_14681);
nand U19075 (N_19075,N_11253,N_10429);
nor U19076 (N_19076,N_10731,N_13787);
nand U19077 (N_19077,N_10388,N_11629);
and U19078 (N_19078,N_12282,N_11462);
xnor U19079 (N_19079,N_10859,N_13461);
and U19080 (N_19080,N_10719,N_13648);
and U19081 (N_19081,N_11070,N_14955);
or U19082 (N_19082,N_12376,N_14412);
or U19083 (N_19083,N_11047,N_10266);
xor U19084 (N_19084,N_14855,N_14640);
nor U19085 (N_19085,N_14145,N_14524);
nor U19086 (N_19086,N_13776,N_11203);
nor U19087 (N_19087,N_11908,N_11749);
and U19088 (N_19088,N_10090,N_10401);
nand U19089 (N_19089,N_13302,N_13355);
and U19090 (N_19090,N_10620,N_13517);
and U19091 (N_19091,N_14688,N_13178);
nand U19092 (N_19092,N_13872,N_13808);
nor U19093 (N_19093,N_14836,N_14719);
nand U19094 (N_19094,N_11548,N_13667);
nand U19095 (N_19095,N_13737,N_10723);
nor U19096 (N_19096,N_13507,N_10053);
nor U19097 (N_19097,N_14084,N_14458);
nand U19098 (N_19098,N_12430,N_13064);
xor U19099 (N_19099,N_13058,N_14663);
and U19100 (N_19100,N_11886,N_12066);
nand U19101 (N_19101,N_10956,N_11700);
xnor U19102 (N_19102,N_12345,N_13823);
or U19103 (N_19103,N_12615,N_10310);
nor U19104 (N_19104,N_11118,N_11981);
and U19105 (N_19105,N_10239,N_12882);
nor U19106 (N_19106,N_13970,N_14524);
or U19107 (N_19107,N_11129,N_14695);
nand U19108 (N_19108,N_12769,N_13444);
and U19109 (N_19109,N_10508,N_10073);
and U19110 (N_19110,N_13701,N_14485);
nor U19111 (N_19111,N_10627,N_14286);
nand U19112 (N_19112,N_13545,N_14470);
nand U19113 (N_19113,N_12972,N_11472);
nor U19114 (N_19114,N_13283,N_12327);
nand U19115 (N_19115,N_11253,N_14965);
nor U19116 (N_19116,N_14103,N_13587);
nor U19117 (N_19117,N_12882,N_12780);
and U19118 (N_19118,N_11330,N_11397);
nor U19119 (N_19119,N_10689,N_11208);
nor U19120 (N_19120,N_14805,N_14968);
nand U19121 (N_19121,N_12290,N_10950);
or U19122 (N_19122,N_10711,N_11383);
xor U19123 (N_19123,N_14026,N_12080);
nand U19124 (N_19124,N_11341,N_10903);
nand U19125 (N_19125,N_10889,N_14126);
nand U19126 (N_19126,N_14768,N_11223);
nor U19127 (N_19127,N_13009,N_13604);
nor U19128 (N_19128,N_11340,N_10797);
xor U19129 (N_19129,N_13189,N_14755);
nand U19130 (N_19130,N_13162,N_11425);
and U19131 (N_19131,N_14552,N_13517);
or U19132 (N_19132,N_11354,N_12481);
or U19133 (N_19133,N_12951,N_12736);
and U19134 (N_19134,N_10958,N_11976);
nor U19135 (N_19135,N_10880,N_11143);
nand U19136 (N_19136,N_12257,N_14591);
nand U19137 (N_19137,N_13270,N_12069);
xnor U19138 (N_19138,N_10894,N_13570);
and U19139 (N_19139,N_12244,N_10495);
nand U19140 (N_19140,N_11712,N_11744);
and U19141 (N_19141,N_10810,N_14791);
or U19142 (N_19142,N_10946,N_10913);
xor U19143 (N_19143,N_12761,N_14970);
xnor U19144 (N_19144,N_12967,N_11788);
nor U19145 (N_19145,N_10806,N_12879);
or U19146 (N_19146,N_11164,N_10157);
nor U19147 (N_19147,N_13361,N_11276);
nor U19148 (N_19148,N_12120,N_12244);
or U19149 (N_19149,N_10151,N_12730);
or U19150 (N_19150,N_14976,N_10220);
and U19151 (N_19151,N_14199,N_12666);
or U19152 (N_19152,N_13989,N_14407);
nor U19153 (N_19153,N_13637,N_13044);
or U19154 (N_19154,N_12896,N_13276);
nand U19155 (N_19155,N_12349,N_13781);
or U19156 (N_19156,N_12914,N_13568);
and U19157 (N_19157,N_12913,N_10706);
xnor U19158 (N_19158,N_13011,N_12697);
and U19159 (N_19159,N_10122,N_13890);
or U19160 (N_19160,N_13179,N_14958);
xor U19161 (N_19161,N_12498,N_13019);
or U19162 (N_19162,N_11689,N_12244);
or U19163 (N_19163,N_12852,N_11411);
and U19164 (N_19164,N_12942,N_12683);
nor U19165 (N_19165,N_10884,N_14186);
nor U19166 (N_19166,N_11162,N_14080);
nor U19167 (N_19167,N_14228,N_11947);
or U19168 (N_19168,N_13093,N_12229);
nor U19169 (N_19169,N_13862,N_12982);
and U19170 (N_19170,N_10883,N_10228);
nand U19171 (N_19171,N_11274,N_10736);
or U19172 (N_19172,N_11294,N_14599);
and U19173 (N_19173,N_14341,N_12942);
and U19174 (N_19174,N_10037,N_11398);
nor U19175 (N_19175,N_10864,N_10371);
or U19176 (N_19176,N_11281,N_12050);
and U19177 (N_19177,N_14983,N_14677);
nor U19178 (N_19178,N_10671,N_10796);
nor U19179 (N_19179,N_13928,N_11491);
nand U19180 (N_19180,N_11055,N_11128);
or U19181 (N_19181,N_12219,N_11755);
nor U19182 (N_19182,N_10513,N_13133);
nor U19183 (N_19183,N_12738,N_13650);
or U19184 (N_19184,N_12467,N_10223);
or U19185 (N_19185,N_11299,N_14424);
nand U19186 (N_19186,N_13916,N_14657);
or U19187 (N_19187,N_11553,N_12337);
nor U19188 (N_19188,N_14483,N_12297);
or U19189 (N_19189,N_12235,N_14173);
or U19190 (N_19190,N_11732,N_13597);
nor U19191 (N_19191,N_13010,N_11021);
or U19192 (N_19192,N_14025,N_10103);
or U19193 (N_19193,N_11669,N_11988);
and U19194 (N_19194,N_10855,N_13598);
xnor U19195 (N_19195,N_14179,N_14599);
xor U19196 (N_19196,N_13983,N_13279);
nand U19197 (N_19197,N_12569,N_10498);
xor U19198 (N_19198,N_13951,N_14047);
nand U19199 (N_19199,N_14453,N_12683);
nor U19200 (N_19200,N_11373,N_12713);
or U19201 (N_19201,N_14153,N_13961);
nand U19202 (N_19202,N_12341,N_14612);
nand U19203 (N_19203,N_12352,N_10939);
nand U19204 (N_19204,N_13314,N_13342);
or U19205 (N_19205,N_11486,N_12830);
or U19206 (N_19206,N_11965,N_11596);
nand U19207 (N_19207,N_12118,N_14400);
xnor U19208 (N_19208,N_13371,N_11312);
nor U19209 (N_19209,N_14126,N_14686);
nand U19210 (N_19210,N_11498,N_13110);
nand U19211 (N_19211,N_12639,N_14583);
or U19212 (N_19212,N_12011,N_10024);
nand U19213 (N_19213,N_13631,N_11844);
xor U19214 (N_19214,N_11804,N_11988);
and U19215 (N_19215,N_11912,N_14302);
or U19216 (N_19216,N_14333,N_14549);
xnor U19217 (N_19217,N_13726,N_12287);
nand U19218 (N_19218,N_10819,N_12798);
nand U19219 (N_19219,N_13532,N_11935);
or U19220 (N_19220,N_11596,N_14847);
or U19221 (N_19221,N_13795,N_12271);
and U19222 (N_19222,N_10979,N_12013);
and U19223 (N_19223,N_14044,N_12888);
nand U19224 (N_19224,N_10335,N_11353);
nand U19225 (N_19225,N_13706,N_12674);
xor U19226 (N_19226,N_12183,N_14768);
xnor U19227 (N_19227,N_13450,N_11915);
nor U19228 (N_19228,N_14070,N_13951);
nor U19229 (N_19229,N_13057,N_14560);
xor U19230 (N_19230,N_12544,N_10420);
xor U19231 (N_19231,N_10310,N_11255);
nor U19232 (N_19232,N_14978,N_14195);
nand U19233 (N_19233,N_10061,N_14290);
nand U19234 (N_19234,N_12504,N_14651);
xor U19235 (N_19235,N_13338,N_13371);
nand U19236 (N_19236,N_10205,N_10871);
nor U19237 (N_19237,N_10885,N_14105);
nand U19238 (N_19238,N_10434,N_12361);
nor U19239 (N_19239,N_14905,N_12900);
or U19240 (N_19240,N_11228,N_11370);
and U19241 (N_19241,N_13404,N_14171);
and U19242 (N_19242,N_11598,N_11159);
or U19243 (N_19243,N_11165,N_10401);
xnor U19244 (N_19244,N_12497,N_11829);
xor U19245 (N_19245,N_12613,N_11194);
nand U19246 (N_19246,N_13863,N_10101);
nor U19247 (N_19247,N_12573,N_12013);
or U19248 (N_19248,N_13447,N_14696);
and U19249 (N_19249,N_10036,N_13615);
xor U19250 (N_19250,N_14693,N_14165);
nor U19251 (N_19251,N_10963,N_12429);
and U19252 (N_19252,N_11794,N_14212);
nor U19253 (N_19253,N_11043,N_14617);
or U19254 (N_19254,N_12217,N_10666);
or U19255 (N_19255,N_11706,N_10482);
nor U19256 (N_19256,N_14849,N_10860);
nand U19257 (N_19257,N_13911,N_13499);
nand U19258 (N_19258,N_13237,N_12268);
nand U19259 (N_19259,N_10466,N_13904);
xnor U19260 (N_19260,N_10394,N_13403);
or U19261 (N_19261,N_11338,N_10524);
and U19262 (N_19262,N_10140,N_10050);
nand U19263 (N_19263,N_13127,N_11066);
nor U19264 (N_19264,N_13151,N_10254);
and U19265 (N_19265,N_12980,N_10048);
nor U19266 (N_19266,N_13735,N_12750);
xnor U19267 (N_19267,N_12789,N_12247);
xor U19268 (N_19268,N_14546,N_13775);
nor U19269 (N_19269,N_12773,N_13932);
xor U19270 (N_19270,N_12546,N_10159);
or U19271 (N_19271,N_10980,N_12827);
xor U19272 (N_19272,N_10342,N_10898);
or U19273 (N_19273,N_12232,N_11197);
nand U19274 (N_19274,N_10936,N_14943);
and U19275 (N_19275,N_12110,N_12924);
nor U19276 (N_19276,N_11148,N_13309);
nor U19277 (N_19277,N_12084,N_10436);
and U19278 (N_19278,N_11869,N_13154);
xnor U19279 (N_19279,N_13801,N_12085);
or U19280 (N_19280,N_11117,N_11474);
or U19281 (N_19281,N_13816,N_14306);
or U19282 (N_19282,N_12869,N_12348);
nand U19283 (N_19283,N_11820,N_12478);
nand U19284 (N_19284,N_11942,N_14575);
nor U19285 (N_19285,N_10990,N_10778);
and U19286 (N_19286,N_13591,N_14026);
nor U19287 (N_19287,N_11167,N_14871);
nor U19288 (N_19288,N_11133,N_10164);
nand U19289 (N_19289,N_10729,N_14370);
nor U19290 (N_19290,N_14836,N_12190);
nand U19291 (N_19291,N_12869,N_10222);
and U19292 (N_19292,N_10275,N_14749);
nand U19293 (N_19293,N_12842,N_14398);
xor U19294 (N_19294,N_10311,N_12528);
and U19295 (N_19295,N_10378,N_13235);
or U19296 (N_19296,N_13722,N_11389);
xnor U19297 (N_19297,N_11491,N_14729);
nand U19298 (N_19298,N_12820,N_14634);
and U19299 (N_19299,N_11851,N_13907);
xor U19300 (N_19300,N_11717,N_12275);
and U19301 (N_19301,N_10685,N_12107);
nor U19302 (N_19302,N_13468,N_14461);
nand U19303 (N_19303,N_13159,N_14830);
nand U19304 (N_19304,N_11736,N_13391);
nor U19305 (N_19305,N_12398,N_14144);
nand U19306 (N_19306,N_12663,N_12920);
or U19307 (N_19307,N_13681,N_12635);
nor U19308 (N_19308,N_14994,N_11677);
xnor U19309 (N_19309,N_13120,N_13383);
nand U19310 (N_19310,N_12341,N_14584);
or U19311 (N_19311,N_14786,N_12680);
nor U19312 (N_19312,N_12521,N_13758);
nor U19313 (N_19313,N_12026,N_10718);
nand U19314 (N_19314,N_13823,N_13167);
nor U19315 (N_19315,N_11288,N_12213);
nand U19316 (N_19316,N_11457,N_11684);
nor U19317 (N_19317,N_14801,N_11664);
and U19318 (N_19318,N_13664,N_13179);
or U19319 (N_19319,N_10944,N_11614);
xor U19320 (N_19320,N_13661,N_12240);
and U19321 (N_19321,N_11478,N_12829);
nand U19322 (N_19322,N_12500,N_12256);
xnor U19323 (N_19323,N_10503,N_10386);
nand U19324 (N_19324,N_11564,N_12533);
nand U19325 (N_19325,N_10788,N_10061);
or U19326 (N_19326,N_11942,N_14403);
nand U19327 (N_19327,N_11165,N_12674);
and U19328 (N_19328,N_12878,N_14249);
nand U19329 (N_19329,N_12317,N_10413);
and U19330 (N_19330,N_12877,N_11126);
or U19331 (N_19331,N_10461,N_14808);
nand U19332 (N_19332,N_14891,N_12794);
nand U19333 (N_19333,N_12553,N_12343);
nand U19334 (N_19334,N_12405,N_12510);
and U19335 (N_19335,N_11837,N_10524);
and U19336 (N_19336,N_14485,N_10309);
nor U19337 (N_19337,N_11623,N_10540);
and U19338 (N_19338,N_11629,N_12133);
nand U19339 (N_19339,N_13122,N_12277);
xnor U19340 (N_19340,N_11700,N_10868);
xnor U19341 (N_19341,N_11388,N_14307);
and U19342 (N_19342,N_13423,N_12730);
xnor U19343 (N_19343,N_11653,N_14202);
nor U19344 (N_19344,N_12506,N_10975);
nand U19345 (N_19345,N_12433,N_11402);
or U19346 (N_19346,N_10238,N_12288);
nor U19347 (N_19347,N_11042,N_10230);
and U19348 (N_19348,N_12591,N_12082);
and U19349 (N_19349,N_10697,N_11038);
nor U19350 (N_19350,N_11812,N_10659);
or U19351 (N_19351,N_14980,N_12718);
xor U19352 (N_19352,N_13082,N_11038);
nand U19353 (N_19353,N_14030,N_13808);
nand U19354 (N_19354,N_11646,N_12626);
xnor U19355 (N_19355,N_11509,N_13912);
nor U19356 (N_19356,N_12003,N_14748);
and U19357 (N_19357,N_13828,N_14024);
nand U19358 (N_19358,N_10164,N_14661);
or U19359 (N_19359,N_13932,N_11227);
nand U19360 (N_19360,N_13456,N_13787);
nor U19361 (N_19361,N_12450,N_11408);
and U19362 (N_19362,N_11770,N_11033);
nand U19363 (N_19363,N_10906,N_10426);
xor U19364 (N_19364,N_12869,N_12890);
xor U19365 (N_19365,N_14335,N_14943);
xnor U19366 (N_19366,N_12177,N_14291);
and U19367 (N_19367,N_11928,N_12952);
xnor U19368 (N_19368,N_12844,N_13349);
xnor U19369 (N_19369,N_13502,N_14534);
nand U19370 (N_19370,N_11551,N_10143);
nor U19371 (N_19371,N_10620,N_11157);
xor U19372 (N_19372,N_13012,N_11009);
nor U19373 (N_19373,N_14332,N_13545);
xnor U19374 (N_19374,N_14237,N_10909);
or U19375 (N_19375,N_14105,N_14656);
nand U19376 (N_19376,N_13602,N_12619);
nor U19377 (N_19377,N_11657,N_10319);
and U19378 (N_19378,N_11874,N_14591);
xnor U19379 (N_19379,N_14283,N_13779);
xnor U19380 (N_19380,N_12720,N_10218);
nand U19381 (N_19381,N_12074,N_14210);
nor U19382 (N_19382,N_14415,N_13545);
and U19383 (N_19383,N_14221,N_13591);
and U19384 (N_19384,N_10125,N_13677);
nor U19385 (N_19385,N_13437,N_10665);
and U19386 (N_19386,N_10060,N_10565);
and U19387 (N_19387,N_13063,N_14558);
or U19388 (N_19388,N_10000,N_11339);
or U19389 (N_19389,N_14412,N_10781);
nand U19390 (N_19390,N_12243,N_10174);
and U19391 (N_19391,N_13966,N_14093);
xnor U19392 (N_19392,N_12020,N_11246);
nor U19393 (N_19393,N_13317,N_12674);
xor U19394 (N_19394,N_10767,N_14730);
and U19395 (N_19395,N_11835,N_12745);
nor U19396 (N_19396,N_10374,N_13186);
nand U19397 (N_19397,N_13277,N_11100);
nor U19398 (N_19398,N_13533,N_11946);
and U19399 (N_19399,N_11829,N_10445);
nor U19400 (N_19400,N_12715,N_11353);
and U19401 (N_19401,N_12929,N_12055);
xor U19402 (N_19402,N_13358,N_13820);
nor U19403 (N_19403,N_10718,N_13759);
and U19404 (N_19404,N_10989,N_13534);
nor U19405 (N_19405,N_10916,N_12785);
or U19406 (N_19406,N_14798,N_11042);
or U19407 (N_19407,N_14515,N_12907);
nand U19408 (N_19408,N_14324,N_10895);
nand U19409 (N_19409,N_13752,N_14902);
or U19410 (N_19410,N_12135,N_12168);
nand U19411 (N_19411,N_14861,N_13224);
xor U19412 (N_19412,N_11392,N_10139);
and U19413 (N_19413,N_12273,N_10954);
nand U19414 (N_19414,N_14944,N_13176);
and U19415 (N_19415,N_13317,N_10912);
or U19416 (N_19416,N_10870,N_11554);
xor U19417 (N_19417,N_14378,N_13736);
or U19418 (N_19418,N_12804,N_11030);
or U19419 (N_19419,N_13682,N_13363);
nor U19420 (N_19420,N_10471,N_13617);
nand U19421 (N_19421,N_14144,N_14098);
or U19422 (N_19422,N_13277,N_10330);
nor U19423 (N_19423,N_13579,N_11653);
and U19424 (N_19424,N_10697,N_14330);
and U19425 (N_19425,N_14694,N_14616);
and U19426 (N_19426,N_13760,N_12782);
nand U19427 (N_19427,N_11458,N_12593);
nand U19428 (N_19428,N_12058,N_14128);
nand U19429 (N_19429,N_13592,N_13706);
xnor U19430 (N_19430,N_13180,N_11990);
or U19431 (N_19431,N_13245,N_11501);
or U19432 (N_19432,N_14435,N_10007);
nor U19433 (N_19433,N_11993,N_10641);
or U19434 (N_19434,N_11539,N_14710);
and U19435 (N_19435,N_11736,N_13680);
nand U19436 (N_19436,N_10283,N_10900);
xor U19437 (N_19437,N_12150,N_10635);
nor U19438 (N_19438,N_12174,N_10318);
nand U19439 (N_19439,N_14925,N_13832);
nand U19440 (N_19440,N_13053,N_11685);
nand U19441 (N_19441,N_12273,N_10538);
nand U19442 (N_19442,N_14800,N_13919);
nand U19443 (N_19443,N_11999,N_13254);
nand U19444 (N_19444,N_13111,N_11093);
nand U19445 (N_19445,N_11388,N_13848);
nand U19446 (N_19446,N_12700,N_13064);
or U19447 (N_19447,N_13256,N_10960);
nor U19448 (N_19448,N_12173,N_10810);
nand U19449 (N_19449,N_11170,N_11845);
and U19450 (N_19450,N_10183,N_14583);
or U19451 (N_19451,N_10980,N_14525);
or U19452 (N_19452,N_10299,N_13509);
xor U19453 (N_19453,N_13376,N_14386);
or U19454 (N_19454,N_12875,N_10899);
nand U19455 (N_19455,N_13877,N_13862);
nand U19456 (N_19456,N_13478,N_13093);
nand U19457 (N_19457,N_12448,N_10320);
nand U19458 (N_19458,N_12395,N_12720);
and U19459 (N_19459,N_10223,N_12853);
nand U19460 (N_19460,N_10722,N_13037);
nor U19461 (N_19461,N_11823,N_11950);
nor U19462 (N_19462,N_11469,N_10722);
or U19463 (N_19463,N_13555,N_10843);
nor U19464 (N_19464,N_10995,N_10609);
or U19465 (N_19465,N_12118,N_13485);
nor U19466 (N_19466,N_14159,N_14707);
nand U19467 (N_19467,N_12561,N_12145);
nor U19468 (N_19468,N_11994,N_13691);
or U19469 (N_19469,N_14601,N_12754);
or U19470 (N_19470,N_11843,N_11772);
nor U19471 (N_19471,N_10182,N_13786);
nand U19472 (N_19472,N_12582,N_14302);
or U19473 (N_19473,N_14638,N_13926);
xnor U19474 (N_19474,N_14325,N_12108);
xnor U19475 (N_19475,N_13853,N_12784);
and U19476 (N_19476,N_14260,N_14827);
nor U19477 (N_19477,N_10634,N_10982);
xnor U19478 (N_19478,N_13894,N_13354);
nand U19479 (N_19479,N_14004,N_10846);
xor U19480 (N_19480,N_10763,N_14007);
nand U19481 (N_19481,N_12265,N_12728);
and U19482 (N_19482,N_14212,N_10928);
or U19483 (N_19483,N_10895,N_11265);
and U19484 (N_19484,N_13767,N_12514);
or U19485 (N_19485,N_10536,N_12971);
or U19486 (N_19486,N_10644,N_10203);
nand U19487 (N_19487,N_12283,N_10204);
and U19488 (N_19488,N_13293,N_13816);
xnor U19489 (N_19489,N_12928,N_14471);
or U19490 (N_19490,N_13461,N_11363);
xor U19491 (N_19491,N_11784,N_14053);
nor U19492 (N_19492,N_12148,N_10443);
nand U19493 (N_19493,N_11991,N_13554);
nor U19494 (N_19494,N_11554,N_14695);
nor U19495 (N_19495,N_11951,N_14213);
or U19496 (N_19496,N_14259,N_12726);
nor U19497 (N_19497,N_10553,N_13553);
nor U19498 (N_19498,N_14278,N_13196);
xor U19499 (N_19499,N_10543,N_11089);
xor U19500 (N_19500,N_14470,N_11266);
xor U19501 (N_19501,N_11495,N_12150);
nand U19502 (N_19502,N_12460,N_14338);
and U19503 (N_19503,N_12714,N_10254);
nor U19504 (N_19504,N_12149,N_11926);
nor U19505 (N_19505,N_14360,N_10693);
nand U19506 (N_19506,N_12389,N_13472);
nand U19507 (N_19507,N_14540,N_14887);
xnor U19508 (N_19508,N_10609,N_13414);
nand U19509 (N_19509,N_14711,N_11646);
and U19510 (N_19510,N_14080,N_14009);
nor U19511 (N_19511,N_12539,N_12772);
nand U19512 (N_19512,N_10711,N_11315);
or U19513 (N_19513,N_10566,N_13205);
nand U19514 (N_19514,N_11613,N_12210);
or U19515 (N_19515,N_11871,N_11558);
nand U19516 (N_19516,N_12218,N_10357);
nand U19517 (N_19517,N_10591,N_13837);
nand U19518 (N_19518,N_12154,N_14686);
or U19519 (N_19519,N_12083,N_10374);
xnor U19520 (N_19520,N_13153,N_10056);
xor U19521 (N_19521,N_14627,N_12663);
or U19522 (N_19522,N_11609,N_12642);
and U19523 (N_19523,N_13763,N_13352);
xor U19524 (N_19524,N_10543,N_11333);
nor U19525 (N_19525,N_13150,N_10364);
xor U19526 (N_19526,N_12364,N_11484);
xor U19527 (N_19527,N_10111,N_10011);
nand U19528 (N_19528,N_11556,N_13874);
or U19529 (N_19529,N_10901,N_11980);
xor U19530 (N_19530,N_14906,N_10476);
and U19531 (N_19531,N_14062,N_14126);
xor U19532 (N_19532,N_11522,N_10373);
nor U19533 (N_19533,N_14913,N_11779);
xor U19534 (N_19534,N_14953,N_12812);
or U19535 (N_19535,N_12968,N_12534);
nor U19536 (N_19536,N_14395,N_11853);
or U19537 (N_19537,N_10597,N_11195);
nand U19538 (N_19538,N_13404,N_11058);
or U19539 (N_19539,N_12349,N_14380);
xor U19540 (N_19540,N_13902,N_14203);
xor U19541 (N_19541,N_10612,N_10809);
and U19542 (N_19542,N_10496,N_13771);
nor U19543 (N_19543,N_11654,N_11154);
and U19544 (N_19544,N_13777,N_10207);
and U19545 (N_19545,N_14609,N_13490);
nor U19546 (N_19546,N_10513,N_12694);
and U19547 (N_19547,N_13261,N_14430);
xnor U19548 (N_19548,N_11495,N_10989);
or U19549 (N_19549,N_10000,N_13120);
nand U19550 (N_19550,N_11829,N_13724);
xnor U19551 (N_19551,N_11437,N_13420);
and U19552 (N_19552,N_12937,N_11149);
and U19553 (N_19553,N_13056,N_10061);
and U19554 (N_19554,N_14853,N_14801);
or U19555 (N_19555,N_13663,N_12306);
or U19556 (N_19556,N_13278,N_14704);
and U19557 (N_19557,N_10968,N_14441);
and U19558 (N_19558,N_11204,N_13867);
or U19559 (N_19559,N_10364,N_13065);
and U19560 (N_19560,N_14500,N_13904);
xnor U19561 (N_19561,N_13792,N_10650);
and U19562 (N_19562,N_14262,N_13811);
and U19563 (N_19563,N_13259,N_11263);
nand U19564 (N_19564,N_11463,N_13907);
and U19565 (N_19565,N_11550,N_13018);
or U19566 (N_19566,N_14633,N_10450);
or U19567 (N_19567,N_14816,N_13474);
or U19568 (N_19568,N_13564,N_12731);
xnor U19569 (N_19569,N_14483,N_14202);
xor U19570 (N_19570,N_13082,N_13481);
nor U19571 (N_19571,N_13269,N_10237);
nor U19572 (N_19572,N_12263,N_13326);
and U19573 (N_19573,N_13888,N_12659);
nor U19574 (N_19574,N_14266,N_13712);
nand U19575 (N_19575,N_13724,N_11923);
and U19576 (N_19576,N_12696,N_13569);
nand U19577 (N_19577,N_14870,N_14756);
xnor U19578 (N_19578,N_10665,N_10937);
or U19579 (N_19579,N_14210,N_12672);
and U19580 (N_19580,N_12646,N_10941);
nand U19581 (N_19581,N_13666,N_11870);
or U19582 (N_19582,N_11207,N_14396);
or U19583 (N_19583,N_10862,N_14888);
nor U19584 (N_19584,N_12998,N_11256);
nor U19585 (N_19585,N_10102,N_11572);
nand U19586 (N_19586,N_14284,N_11357);
xnor U19587 (N_19587,N_11288,N_13867);
nand U19588 (N_19588,N_11356,N_12529);
and U19589 (N_19589,N_12727,N_10571);
nand U19590 (N_19590,N_12097,N_10353);
and U19591 (N_19591,N_14817,N_13906);
or U19592 (N_19592,N_13320,N_13420);
nand U19593 (N_19593,N_14777,N_11908);
xor U19594 (N_19594,N_13656,N_12364);
xnor U19595 (N_19595,N_13332,N_12235);
or U19596 (N_19596,N_14756,N_13332);
nor U19597 (N_19597,N_13531,N_13082);
and U19598 (N_19598,N_11969,N_12020);
nand U19599 (N_19599,N_13088,N_13505);
or U19600 (N_19600,N_14836,N_10901);
and U19601 (N_19601,N_11931,N_14700);
and U19602 (N_19602,N_10939,N_12186);
nand U19603 (N_19603,N_13013,N_11162);
nand U19604 (N_19604,N_14603,N_11993);
and U19605 (N_19605,N_10407,N_12519);
xor U19606 (N_19606,N_10785,N_13049);
nand U19607 (N_19607,N_14507,N_12781);
nand U19608 (N_19608,N_14962,N_12811);
nor U19609 (N_19609,N_10981,N_11259);
nand U19610 (N_19610,N_13659,N_13744);
xor U19611 (N_19611,N_11440,N_14909);
nor U19612 (N_19612,N_13614,N_12221);
xor U19613 (N_19613,N_12626,N_10803);
nand U19614 (N_19614,N_11213,N_12401);
or U19615 (N_19615,N_11455,N_12440);
or U19616 (N_19616,N_13627,N_10991);
and U19617 (N_19617,N_10741,N_13936);
or U19618 (N_19618,N_13444,N_14155);
and U19619 (N_19619,N_12342,N_14481);
and U19620 (N_19620,N_14635,N_11786);
xnor U19621 (N_19621,N_14275,N_13616);
and U19622 (N_19622,N_13433,N_14395);
xor U19623 (N_19623,N_11792,N_14136);
nor U19624 (N_19624,N_12968,N_13825);
nor U19625 (N_19625,N_12844,N_12489);
nand U19626 (N_19626,N_14235,N_13881);
or U19627 (N_19627,N_12398,N_11494);
or U19628 (N_19628,N_10472,N_14675);
and U19629 (N_19629,N_14403,N_11425);
or U19630 (N_19630,N_12333,N_10531);
nor U19631 (N_19631,N_12788,N_12537);
or U19632 (N_19632,N_14159,N_11928);
xnor U19633 (N_19633,N_11699,N_12865);
xnor U19634 (N_19634,N_11291,N_11053);
nor U19635 (N_19635,N_12454,N_12243);
nor U19636 (N_19636,N_13512,N_12112);
and U19637 (N_19637,N_10273,N_11365);
xor U19638 (N_19638,N_14025,N_10366);
nor U19639 (N_19639,N_13587,N_14329);
or U19640 (N_19640,N_11165,N_12017);
nor U19641 (N_19641,N_11204,N_12539);
nor U19642 (N_19642,N_10864,N_11174);
or U19643 (N_19643,N_14769,N_13751);
xor U19644 (N_19644,N_11586,N_13779);
xor U19645 (N_19645,N_10124,N_13515);
xor U19646 (N_19646,N_13103,N_10136);
and U19647 (N_19647,N_14737,N_10339);
nand U19648 (N_19648,N_10677,N_13897);
or U19649 (N_19649,N_10901,N_13954);
xnor U19650 (N_19650,N_12341,N_12929);
and U19651 (N_19651,N_12227,N_14399);
nand U19652 (N_19652,N_10463,N_10438);
nor U19653 (N_19653,N_12782,N_11051);
and U19654 (N_19654,N_14413,N_13921);
and U19655 (N_19655,N_13973,N_14636);
xnor U19656 (N_19656,N_14199,N_14013);
nand U19657 (N_19657,N_14335,N_11587);
nor U19658 (N_19658,N_14172,N_13232);
nand U19659 (N_19659,N_14853,N_13843);
xnor U19660 (N_19660,N_13636,N_14765);
xor U19661 (N_19661,N_10806,N_11280);
or U19662 (N_19662,N_13985,N_11475);
and U19663 (N_19663,N_11431,N_12245);
or U19664 (N_19664,N_14227,N_11878);
nor U19665 (N_19665,N_12269,N_10578);
and U19666 (N_19666,N_12792,N_11893);
and U19667 (N_19667,N_13816,N_11562);
xor U19668 (N_19668,N_13998,N_10853);
and U19669 (N_19669,N_11651,N_10456);
and U19670 (N_19670,N_10009,N_13857);
xor U19671 (N_19671,N_13490,N_14502);
nor U19672 (N_19672,N_10672,N_13719);
nand U19673 (N_19673,N_13945,N_13160);
nand U19674 (N_19674,N_12745,N_10977);
and U19675 (N_19675,N_12017,N_11696);
nor U19676 (N_19676,N_11134,N_12987);
nor U19677 (N_19677,N_10056,N_10526);
nand U19678 (N_19678,N_10170,N_12967);
nor U19679 (N_19679,N_10589,N_12258);
and U19680 (N_19680,N_10706,N_12622);
nand U19681 (N_19681,N_12279,N_14032);
nand U19682 (N_19682,N_11631,N_14562);
xor U19683 (N_19683,N_13660,N_13437);
and U19684 (N_19684,N_10944,N_10354);
nor U19685 (N_19685,N_14495,N_14889);
nor U19686 (N_19686,N_12863,N_12385);
nor U19687 (N_19687,N_12494,N_13703);
xor U19688 (N_19688,N_13944,N_14033);
and U19689 (N_19689,N_13950,N_12341);
and U19690 (N_19690,N_13081,N_14285);
xor U19691 (N_19691,N_11091,N_11411);
or U19692 (N_19692,N_14671,N_14407);
xnor U19693 (N_19693,N_14749,N_11347);
nor U19694 (N_19694,N_13564,N_12923);
and U19695 (N_19695,N_11069,N_14691);
or U19696 (N_19696,N_13007,N_13821);
nor U19697 (N_19697,N_10767,N_12279);
nor U19698 (N_19698,N_12977,N_13263);
nand U19699 (N_19699,N_14142,N_12043);
nand U19700 (N_19700,N_11254,N_14559);
or U19701 (N_19701,N_12360,N_10032);
nor U19702 (N_19702,N_10060,N_12245);
and U19703 (N_19703,N_14642,N_14821);
or U19704 (N_19704,N_11481,N_13665);
or U19705 (N_19705,N_12405,N_11347);
nand U19706 (N_19706,N_10127,N_10619);
nand U19707 (N_19707,N_11237,N_12113);
nand U19708 (N_19708,N_12316,N_11794);
nand U19709 (N_19709,N_14190,N_13544);
or U19710 (N_19710,N_14562,N_11797);
xnor U19711 (N_19711,N_14934,N_14779);
xor U19712 (N_19712,N_14660,N_12994);
nor U19713 (N_19713,N_11146,N_10268);
nand U19714 (N_19714,N_14656,N_11603);
xnor U19715 (N_19715,N_13104,N_13454);
nor U19716 (N_19716,N_10801,N_13315);
nor U19717 (N_19717,N_12585,N_12793);
xnor U19718 (N_19718,N_13887,N_14482);
or U19719 (N_19719,N_10525,N_13613);
nand U19720 (N_19720,N_14821,N_13966);
nor U19721 (N_19721,N_13383,N_10990);
and U19722 (N_19722,N_11300,N_11628);
nor U19723 (N_19723,N_12258,N_10365);
and U19724 (N_19724,N_11408,N_14767);
nor U19725 (N_19725,N_14299,N_13449);
nand U19726 (N_19726,N_12416,N_12625);
nor U19727 (N_19727,N_14187,N_12755);
or U19728 (N_19728,N_12244,N_14837);
and U19729 (N_19729,N_10746,N_12782);
xor U19730 (N_19730,N_12741,N_11767);
or U19731 (N_19731,N_13193,N_14695);
nor U19732 (N_19732,N_11003,N_13174);
nand U19733 (N_19733,N_13441,N_12873);
nand U19734 (N_19734,N_14986,N_12002);
nor U19735 (N_19735,N_10007,N_13462);
xor U19736 (N_19736,N_12111,N_11745);
xnor U19737 (N_19737,N_12474,N_13245);
xor U19738 (N_19738,N_12218,N_11660);
nor U19739 (N_19739,N_14126,N_14777);
and U19740 (N_19740,N_11085,N_13132);
xor U19741 (N_19741,N_10457,N_14486);
xnor U19742 (N_19742,N_14417,N_11764);
nor U19743 (N_19743,N_12686,N_11907);
or U19744 (N_19744,N_11626,N_13099);
nand U19745 (N_19745,N_12540,N_11480);
nand U19746 (N_19746,N_11570,N_12509);
and U19747 (N_19747,N_13358,N_13500);
xor U19748 (N_19748,N_14545,N_10214);
and U19749 (N_19749,N_12890,N_14945);
or U19750 (N_19750,N_12315,N_13612);
xor U19751 (N_19751,N_13521,N_13419);
or U19752 (N_19752,N_12411,N_10084);
xnor U19753 (N_19753,N_13740,N_11737);
or U19754 (N_19754,N_12423,N_11752);
nor U19755 (N_19755,N_14130,N_12789);
nor U19756 (N_19756,N_13305,N_11550);
and U19757 (N_19757,N_14609,N_13205);
or U19758 (N_19758,N_14266,N_13085);
nand U19759 (N_19759,N_13768,N_12603);
xor U19760 (N_19760,N_14864,N_14078);
xor U19761 (N_19761,N_11348,N_13826);
nand U19762 (N_19762,N_13887,N_13339);
nand U19763 (N_19763,N_12851,N_14052);
and U19764 (N_19764,N_11002,N_13678);
nand U19765 (N_19765,N_13741,N_10864);
nand U19766 (N_19766,N_11102,N_13717);
or U19767 (N_19767,N_13275,N_11227);
and U19768 (N_19768,N_11484,N_11042);
and U19769 (N_19769,N_12638,N_12070);
or U19770 (N_19770,N_14874,N_11690);
or U19771 (N_19771,N_12957,N_12430);
or U19772 (N_19772,N_12732,N_13681);
and U19773 (N_19773,N_12121,N_11927);
nor U19774 (N_19774,N_10466,N_12095);
nor U19775 (N_19775,N_14643,N_10900);
and U19776 (N_19776,N_11964,N_14162);
or U19777 (N_19777,N_13223,N_11976);
xor U19778 (N_19778,N_11184,N_12669);
and U19779 (N_19779,N_10837,N_14017);
and U19780 (N_19780,N_13376,N_14177);
or U19781 (N_19781,N_12509,N_14092);
nand U19782 (N_19782,N_14792,N_12221);
and U19783 (N_19783,N_10224,N_11665);
xor U19784 (N_19784,N_11586,N_14445);
xor U19785 (N_19785,N_11944,N_14654);
xnor U19786 (N_19786,N_10568,N_13150);
or U19787 (N_19787,N_11072,N_13958);
xor U19788 (N_19788,N_14813,N_13674);
nand U19789 (N_19789,N_10449,N_14692);
or U19790 (N_19790,N_11751,N_11124);
and U19791 (N_19791,N_13564,N_12279);
nand U19792 (N_19792,N_11701,N_13952);
nand U19793 (N_19793,N_11752,N_10901);
and U19794 (N_19794,N_14613,N_13777);
nand U19795 (N_19795,N_13085,N_12542);
nand U19796 (N_19796,N_13104,N_12298);
nand U19797 (N_19797,N_12433,N_10856);
nand U19798 (N_19798,N_13305,N_11463);
and U19799 (N_19799,N_11026,N_10476);
xor U19800 (N_19800,N_13180,N_11275);
and U19801 (N_19801,N_10532,N_11466);
nand U19802 (N_19802,N_12222,N_11141);
nor U19803 (N_19803,N_13926,N_11740);
xnor U19804 (N_19804,N_12623,N_11560);
and U19805 (N_19805,N_11557,N_13640);
nand U19806 (N_19806,N_11077,N_13282);
nor U19807 (N_19807,N_11610,N_14516);
xor U19808 (N_19808,N_14891,N_13483);
or U19809 (N_19809,N_12734,N_14564);
nand U19810 (N_19810,N_14371,N_13873);
nand U19811 (N_19811,N_13688,N_11215);
nand U19812 (N_19812,N_12427,N_14486);
nand U19813 (N_19813,N_14178,N_12559);
xnor U19814 (N_19814,N_14896,N_13680);
and U19815 (N_19815,N_10209,N_12961);
or U19816 (N_19816,N_14380,N_12970);
xor U19817 (N_19817,N_14241,N_12814);
and U19818 (N_19818,N_12022,N_13085);
nor U19819 (N_19819,N_13075,N_10329);
nor U19820 (N_19820,N_13301,N_11326);
nand U19821 (N_19821,N_12308,N_11632);
or U19822 (N_19822,N_14145,N_14724);
nand U19823 (N_19823,N_13432,N_10744);
and U19824 (N_19824,N_12984,N_14738);
nor U19825 (N_19825,N_12106,N_14278);
and U19826 (N_19826,N_11085,N_12111);
nand U19827 (N_19827,N_11005,N_11945);
nand U19828 (N_19828,N_14900,N_12750);
or U19829 (N_19829,N_11842,N_13717);
and U19830 (N_19830,N_11986,N_14259);
or U19831 (N_19831,N_10382,N_13730);
xor U19832 (N_19832,N_11194,N_11011);
nor U19833 (N_19833,N_10012,N_12966);
nand U19834 (N_19834,N_13274,N_10327);
xor U19835 (N_19835,N_11185,N_11713);
xor U19836 (N_19836,N_14297,N_13981);
xor U19837 (N_19837,N_11025,N_10783);
xor U19838 (N_19838,N_10164,N_14412);
nor U19839 (N_19839,N_12520,N_14987);
and U19840 (N_19840,N_14848,N_10643);
nor U19841 (N_19841,N_10575,N_13519);
and U19842 (N_19842,N_13945,N_13260);
nor U19843 (N_19843,N_10317,N_12130);
nor U19844 (N_19844,N_11360,N_13296);
nor U19845 (N_19845,N_12406,N_11141);
or U19846 (N_19846,N_11272,N_13158);
nor U19847 (N_19847,N_10446,N_11407);
nor U19848 (N_19848,N_11373,N_13771);
xor U19849 (N_19849,N_14080,N_12031);
nor U19850 (N_19850,N_11850,N_10844);
or U19851 (N_19851,N_12813,N_14676);
xor U19852 (N_19852,N_13335,N_11781);
and U19853 (N_19853,N_11030,N_10208);
nor U19854 (N_19854,N_14126,N_13065);
xnor U19855 (N_19855,N_10583,N_14662);
and U19856 (N_19856,N_11747,N_13723);
or U19857 (N_19857,N_14482,N_11132);
xnor U19858 (N_19858,N_14910,N_14173);
nor U19859 (N_19859,N_14953,N_14845);
and U19860 (N_19860,N_13364,N_13388);
xor U19861 (N_19861,N_11022,N_11206);
nor U19862 (N_19862,N_12068,N_10827);
xnor U19863 (N_19863,N_12636,N_12646);
xnor U19864 (N_19864,N_14816,N_11060);
nand U19865 (N_19865,N_10266,N_13839);
nand U19866 (N_19866,N_13072,N_13465);
nand U19867 (N_19867,N_11473,N_11873);
nand U19868 (N_19868,N_11012,N_11466);
nor U19869 (N_19869,N_14574,N_14444);
xnor U19870 (N_19870,N_11218,N_12338);
nor U19871 (N_19871,N_10394,N_11163);
xor U19872 (N_19872,N_11374,N_11555);
and U19873 (N_19873,N_10585,N_14933);
xnor U19874 (N_19874,N_12247,N_13495);
or U19875 (N_19875,N_14935,N_13171);
nor U19876 (N_19876,N_11866,N_13972);
and U19877 (N_19877,N_10410,N_13826);
nand U19878 (N_19878,N_11578,N_11319);
nor U19879 (N_19879,N_11637,N_11349);
and U19880 (N_19880,N_10540,N_10644);
nor U19881 (N_19881,N_14436,N_11814);
xnor U19882 (N_19882,N_14735,N_10236);
and U19883 (N_19883,N_13502,N_10126);
xor U19884 (N_19884,N_13852,N_10371);
nand U19885 (N_19885,N_14056,N_10321);
xnor U19886 (N_19886,N_12453,N_11425);
and U19887 (N_19887,N_10255,N_12105);
nor U19888 (N_19888,N_12325,N_10554);
nor U19889 (N_19889,N_14171,N_11982);
xor U19890 (N_19890,N_13057,N_12307);
and U19891 (N_19891,N_14557,N_11462);
xor U19892 (N_19892,N_12790,N_10366);
xnor U19893 (N_19893,N_12572,N_12838);
or U19894 (N_19894,N_13119,N_12780);
nor U19895 (N_19895,N_10687,N_14195);
nor U19896 (N_19896,N_12993,N_12664);
and U19897 (N_19897,N_10875,N_13487);
nand U19898 (N_19898,N_13840,N_14684);
and U19899 (N_19899,N_14476,N_12852);
nand U19900 (N_19900,N_10268,N_12992);
nand U19901 (N_19901,N_12838,N_14965);
nor U19902 (N_19902,N_11595,N_11699);
xnor U19903 (N_19903,N_14481,N_10725);
xnor U19904 (N_19904,N_14221,N_10308);
and U19905 (N_19905,N_12883,N_11700);
and U19906 (N_19906,N_12388,N_10859);
nand U19907 (N_19907,N_13262,N_14611);
nor U19908 (N_19908,N_12860,N_14597);
nor U19909 (N_19909,N_11212,N_10486);
xor U19910 (N_19910,N_12472,N_12355);
and U19911 (N_19911,N_10909,N_10857);
xor U19912 (N_19912,N_12332,N_10222);
and U19913 (N_19913,N_12912,N_12755);
or U19914 (N_19914,N_10106,N_12039);
nor U19915 (N_19915,N_10642,N_12633);
and U19916 (N_19916,N_10829,N_11455);
nor U19917 (N_19917,N_12270,N_10792);
nor U19918 (N_19918,N_13948,N_12000);
or U19919 (N_19919,N_12561,N_11187);
and U19920 (N_19920,N_10249,N_11792);
and U19921 (N_19921,N_10797,N_14454);
or U19922 (N_19922,N_12129,N_13476);
or U19923 (N_19923,N_11993,N_13358);
nor U19924 (N_19924,N_11923,N_13898);
nor U19925 (N_19925,N_13372,N_14271);
nand U19926 (N_19926,N_14984,N_14940);
nor U19927 (N_19927,N_14811,N_10367);
nor U19928 (N_19928,N_13193,N_14132);
xor U19929 (N_19929,N_13380,N_13718);
nor U19930 (N_19930,N_10639,N_12396);
or U19931 (N_19931,N_10550,N_10208);
xnor U19932 (N_19932,N_12906,N_10216);
or U19933 (N_19933,N_14721,N_13574);
or U19934 (N_19934,N_14546,N_12479);
or U19935 (N_19935,N_11087,N_10282);
xnor U19936 (N_19936,N_14747,N_10050);
and U19937 (N_19937,N_14449,N_14277);
nor U19938 (N_19938,N_14849,N_14656);
or U19939 (N_19939,N_10498,N_11012);
xor U19940 (N_19940,N_11398,N_12449);
nand U19941 (N_19941,N_12830,N_14000);
and U19942 (N_19942,N_14725,N_14163);
xor U19943 (N_19943,N_13879,N_13446);
or U19944 (N_19944,N_11814,N_13609);
nor U19945 (N_19945,N_14144,N_12025);
or U19946 (N_19946,N_14914,N_12220);
nor U19947 (N_19947,N_13086,N_12584);
xnor U19948 (N_19948,N_10698,N_11635);
and U19949 (N_19949,N_10590,N_12065);
and U19950 (N_19950,N_13377,N_13904);
nor U19951 (N_19951,N_11223,N_13665);
nor U19952 (N_19952,N_10206,N_14467);
nor U19953 (N_19953,N_13985,N_10643);
or U19954 (N_19954,N_11633,N_14356);
or U19955 (N_19955,N_11726,N_13639);
xnor U19956 (N_19956,N_12036,N_14426);
or U19957 (N_19957,N_14215,N_11318);
and U19958 (N_19958,N_12275,N_11564);
and U19959 (N_19959,N_12405,N_13369);
or U19960 (N_19960,N_11320,N_13649);
or U19961 (N_19961,N_12077,N_12712);
and U19962 (N_19962,N_13068,N_12784);
nor U19963 (N_19963,N_14965,N_13006);
and U19964 (N_19964,N_12087,N_11566);
or U19965 (N_19965,N_12959,N_14850);
and U19966 (N_19966,N_13206,N_13862);
or U19967 (N_19967,N_13897,N_10118);
nand U19968 (N_19968,N_11545,N_13700);
and U19969 (N_19969,N_11784,N_13715);
xor U19970 (N_19970,N_13381,N_13314);
and U19971 (N_19971,N_13385,N_11853);
nand U19972 (N_19972,N_10112,N_10990);
and U19973 (N_19973,N_14754,N_13613);
and U19974 (N_19974,N_14006,N_14418);
xor U19975 (N_19975,N_10296,N_13105);
and U19976 (N_19976,N_11439,N_14598);
and U19977 (N_19977,N_10685,N_10903);
nand U19978 (N_19978,N_11231,N_14469);
nor U19979 (N_19979,N_10167,N_12937);
xor U19980 (N_19980,N_14818,N_14396);
xnor U19981 (N_19981,N_14055,N_14887);
and U19982 (N_19982,N_12925,N_13728);
or U19983 (N_19983,N_13637,N_10160);
or U19984 (N_19984,N_13998,N_10915);
nor U19985 (N_19985,N_14950,N_11069);
nand U19986 (N_19986,N_13247,N_12438);
nand U19987 (N_19987,N_12241,N_14000);
nand U19988 (N_19988,N_10077,N_14822);
or U19989 (N_19989,N_10683,N_14635);
and U19990 (N_19990,N_10155,N_12598);
or U19991 (N_19991,N_11745,N_10741);
xnor U19992 (N_19992,N_11371,N_12305);
or U19993 (N_19993,N_13973,N_13054);
nor U19994 (N_19994,N_10724,N_10835);
nor U19995 (N_19995,N_14478,N_12995);
and U19996 (N_19996,N_10725,N_10664);
nand U19997 (N_19997,N_11762,N_12950);
or U19998 (N_19998,N_10015,N_11800);
and U19999 (N_19999,N_14136,N_10083);
or U20000 (N_20000,N_15899,N_18838);
xnor U20001 (N_20001,N_16164,N_18476);
and U20002 (N_20002,N_15265,N_19369);
nand U20003 (N_20003,N_15811,N_16532);
or U20004 (N_20004,N_18416,N_18169);
and U20005 (N_20005,N_17449,N_17645);
and U20006 (N_20006,N_19639,N_17287);
xor U20007 (N_20007,N_16698,N_18814);
nand U20008 (N_20008,N_19073,N_16271);
nand U20009 (N_20009,N_18508,N_19642);
nand U20010 (N_20010,N_19196,N_15962);
xnor U20011 (N_20011,N_16097,N_17982);
nor U20012 (N_20012,N_19388,N_16963);
nor U20013 (N_20013,N_15306,N_19247);
nor U20014 (N_20014,N_18804,N_15398);
and U20015 (N_20015,N_17588,N_17097);
xor U20016 (N_20016,N_19270,N_16380);
and U20017 (N_20017,N_16582,N_18865);
xnor U20018 (N_20018,N_18408,N_16086);
and U20019 (N_20019,N_15296,N_19605);
xnor U20020 (N_20020,N_17635,N_15388);
xnor U20021 (N_20021,N_19376,N_19028);
or U20022 (N_20022,N_17275,N_15600);
and U20023 (N_20023,N_18253,N_15708);
and U20024 (N_20024,N_18751,N_17986);
nand U20025 (N_20025,N_19184,N_16798);
and U20026 (N_20026,N_17028,N_15444);
nor U20027 (N_20027,N_19865,N_18199);
and U20028 (N_20028,N_15266,N_17554);
nor U20029 (N_20029,N_18525,N_19870);
or U20030 (N_20030,N_19275,N_16146);
nand U20031 (N_20031,N_15127,N_15924);
or U20032 (N_20032,N_18321,N_17571);
and U20033 (N_20033,N_19987,N_16690);
and U20034 (N_20034,N_16827,N_16722);
nor U20035 (N_20035,N_19451,N_19128);
and U20036 (N_20036,N_19613,N_19000);
or U20037 (N_20037,N_15568,N_17556);
nor U20038 (N_20038,N_18504,N_15264);
or U20039 (N_20039,N_16976,N_16083);
nand U20040 (N_20040,N_15246,N_18615);
nor U20041 (N_20041,N_15474,N_17011);
xnor U20042 (N_20042,N_18337,N_15299);
nand U20043 (N_20043,N_17881,N_16280);
and U20044 (N_20044,N_17203,N_18786);
nor U20045 (N_20045,N_16784,N_17467);
nor U20046 (N_20046,N_19330,N_19201);
xnor U20047 (N_20047,N_16904,N_19039);
xnor U20048 (N_20048,N_18203,N_15091);
and U20049 (N_20049,N_16687,N_19589);
or U20050 (N_20050,N_16006,N_15241);
nand U20051 (N_20051,N_18839,N_18820);
and U20052 (N_20052,N_16936,N_16817);
xor U20053 (N_20053,N_16064,N_16286);
nand U20054 (N_20054,N_17950,N_18904);
xor U20055 (N_20055,N_18585,N_19161);
nand U20056 (N_20056,N_18538,N_15820);
and U20057 (N_20057,N_19017,N_15861);
xnor U20058 (N_20058,N_17922,N_18734);
or U20059 (N_20059,N_18836,N_18540);
and U20060 (N_20060,N_15448,N_18876);
nand U20061 (N_20061,N_17395,N_19291);
nand U20062 (N_20062,N_16121,N_19647);
or U20063 (N_20063,N_17808,N_16292);
xor U20064 (N_20064,N_17562,N_17494);
or U20065 (N_20065,N_19868,N_16719);
and U20066 (N_20066,N_17811,N_19090);
and U20067 (N_20067,N_16569,N_18668);
nor U20068 (N_20068,N_19449,N_19322);
nand U20069 (N_20069,N_15124,N_16291);
nor U20070 (N_20070,N_18269,N_17429);
nand U20071 (N_20071,N_18545,N_17767);
nand U20072 (N_20072,N_15068,N_17921);
nor U20073 (N_20073,N_18143,N_17594);
and U20074 (N_20074,N_18148,N_16246);
nor U20075 (N_20075,N_16033,N_16343);
nor U20076 (N_20076,N_17798,N_17244);
and U20077 (N_20077,N_16853,N_16010);
xor U20078 (N_20078,N_16840,N_15669);
xnor U20079 (N_20079,N_15193,N_19095);
and U20080 (N_20080,N_17785,N_18149);
nor U20081 (N_20081,N_18139,N_18825);
and U20082 (N_20082,N_17729,N_15510);
or U20083 (N_20083,N_18479,N_18796);
or U20084 (N_20084,N_19816,N_15289);
or U20085 (N_20085,N_16617,N_18245);
or U20086 (N_20086,N_19357,N_16733);
nand U20087 (N_20087,N_16516,N_17602);
or U20088 (N_20088,N_17587,N_15523);
xor U20089 (N_20089,N_15786,N_15873);
or U20090 (N_20090,N_19818,N_17001);
nor U20091 (N_20091,N_16412,N_17697);
nor U20092 (N_20092,N_16908,N_18872);
xor U20093 (N_20093,N_19611,N_18834);
nand U20094 (N_20094,N_18835,N_17178);
or U20095 (N_20095,N_16074,N_17291);
and U20096 (N_20096,N_17955,N_18644);
nor U20097 (N_20097,N_16767,N_18889);
and U20098 (N_20098,N_15944,N_16008);
nor U20099 (N_20099,N_17276,N_16873);
and U20100 (N_20100,N_18930,N_19918);
xor U20101 (N_20101,N_18772,N_17730);
xnor U20102 (N_20102,N_17096,N_17476);
xor U20103 (N_20103,N_18767,N_18600);
xor U20104 (N_20104,N_15544,N_16273);
xnor U20105 (N_20105,N_16051,N_15982);
or U20106 (N_20106,N_18141,N_19525);
nand U20107 (N_20107,N_17719,N_18992);
nor U20108 (N_20108,N_15485,N_17755);
nand U20109 (N_20109,N_16196,N_18305);
nand U20110 (N_20110,N_16552,N_17833);
or U20111 (N_20111,N_18465,N_16169);
and U20112 (N_20112,N_16547,N_19846);
and U20113 (N_20113,N_19656,N_15908);
and U20114 (N_20114,N_16539,N_15524);
nand U20115 (N_20115,N_17609,N_19541);
or U20116 (N_20116,N_15905,N_16180);
nor U20117 (N_20117,N_16898,N_16250);
xnor U20118 (N_20118,N_15431,N_18312);
and U20119 (N_20119,N_16630,N_19547);
nor U20120 (N_20120,N_18156,N_19381);
xnor U20121 (N_20121,N_17453,N_15890);
nor U20122 (N_20122,N_17895,N_15548);
nor U20123 (N_20123,N_17667,N_18678);
nand U20124 (N_20124,N_15619,N_17490);
xnor U20125 (N_20125,N_17945,N_19979);
nand U20126 (N_20126,N_17288,N_15291);
and U20127 (N_20127,N_16759,N_17459);
or U20128 (N_20128,N_19447,N_16805);
nor U20129 (N_20129,N_15043,N_18460);
or U20130 (N_20130,N_19298,N_17089);
xor U20131 (N_20131,N_17825,N_19232);
xnor U20132 (N_20132,N_18415,N_18677);
xor U20133 (N_20133,N_16857,N_17260);
nand U20134 (N_20134,N_17249,N_16483);
nor U20135 (N_20135,N_18639,N_17823);
or U20136 (N_20136,N_19503,N_19934);
and U20137 (N_20137,N_15235,N_16838);
xnor U20138 (N_20138,N_19505,N_15061);
nand U20139 (N_20139,N_19489,N_17427);
xor U20140 (N_20140,N_16761,N_15755);
nor U20141 (N_20141,N_19037,N_17302);
nand U20142 (N_20142,N_15023,N_17295);
nand U20143 (N_20143,N_16636,N_18922);
or U20144 (N_20144,N_18947,N_19137);
or U20145 (N_20145,N_18519,N_15918);
or U20146 (N_20146,N_16392,N_18402);
and U20147 (N_20147,N_19380,N_18941);
or U20148 (N_20148,N_19358,N_15371);
nand U20149 (N_20149,N_19569,N_18687);
xor U20150 (N_20150,N_17840,N_15987);
or U20151 (N_20151,N_17530,N_15116);
xnor U20152 (N_20152,N_17937,N_18469);
nor U20153 (N_20153,N_18628,N_15377);
or U20154 (N_20154,N_18403,N_19335);
xnor U20155 (N_20155,N_19261,N_18393);
nor U20156 (N_20156,N_16365,N_18547);
nand U20157 (N_20157,N_17026,N_18984);
nor U20158 (N_20158,N_17163,N_15624);
xnor U20159 (N_20159,N_15679,N_17149);
and U20160 (N_20160,N_15496,N_16959);
nand U20161 (N_20161,N_19759,N_17054);
or U20162 (N_20162,N_18092,N_18962);
or U20163 (N_20163,N_15034,N_15028);
or U20164 (N_20164,N_17112,N_15693);
nand U20165 (N_20165,N_17100,N_18919);
nor U20166 (N_20166,N_19306,N_19434);
nand U20167 (N_20167,N_15209,N_19096);
xor U20168 (N_20168,N_17417,N_18333);
xor U20169 (N_20169,N_15111,N_17712);
and U20170 (N_20170,N_16803,N_17383);
and U20171 (N_20171,N_18989,N_19431);
and U20172 (N_20172,N_19293,N_15139);
nor U20173 (N_20173,N_16862,N_19627);
xor U20174 (N_20174,N_16682,N_17753);
xnor U20175 (N_20175,N_16608,N_15542);
or U20176 (N_20176,N_16050,N_16397);
or U20177 (N_20177,N_18878,N_19856);
xnor U20178 (N_20178,N_19032,N_15558);
xnor U20179 (N_20179,N_15699,N_18433);
nor U20180 (N_20180,N_17337,N_18349);
and U20181 (N_20181,N_19045,N_16792);
or U20182 (N_20182,N_19114,N_17256);
xnor U20183 (N_20183,N_16821,N_19711);
nand U20184 (N_20184,N_15310,N_15212);
nor U20185 (N_20185,N_19944,N_18478);
xnor U20186 (N_20186,N_18612,N_18590);
nor U20187 (N_20187,N_17359,N_15763);
nand U20188 (N_20188,N_17924,N_17943);
xnor U20189 (N_20189,N_15486,N_17343);
nor U20190 (N_20190,N_18718,N_16334);
or U20191 (N_20191,N_15006,N_19416);
xor U20192 (N_20192,N_17458,N_18944);
and U20193 (N_20193,N_18953,N_19652);
nor U20194 (N_20194,N_17536,N_15706);
nand U20195 (N_20195,N_18068,N_19190);
nor U20196 (N_20196,N_18584,N_18140);
and U20197 (N_20197,N_19477,N_17653);
nor U20198 (N_20198,N_17532,N_19314);
xnor U20199 (N_20199,N_18242,N_16255);
and U20200 (N_20200,N_15141,N_17885);
and U20201 (N_20201,N_17916,N_17122);
nor U20202 (N_20202,N_19708,N_19985);
and U20203 (N_20203,N_17580,N_15260);
nor U20204 (N_20204,N_18692,N_15692);
nor U20205 (N_20205,N_16037,N_16177);
xor U20206 (N_20206,N_18777,N_16345);
nor U20207 (N_20207,N_18499,N_17223);
xnor U20208 (N_20208,N_18917,N_19301);
and U20209 (N_20209,N_16657,N_18495);
xnor U20210 (N_20210,N_15727,N_17118);
and U20211 (N_20211,N_18385,N_19732);
or U20212 (N_20212,N_16409,N_17935);
nand U20213 (N_20213,N_17248,N_15778);
and U20214 (N_20214,N_18029,N_19446);
or U20215 (N_20215,N_17313,N_17592);
or U20216 (N_20216,N_18443,N_18754);
and U20217 (N_20217,N_18317,N_19238);
nor U20218 (N_20218,N_17048,N_15500);
nor U20219 (N_20219,N_17911,N_16531);
and U20220 (N_20220,N_16270,N_17990);
xnor U20221 (N_20221,N_15360,N_19608);
xnor U20222 (N_20222,N_19299,N_18709);
or U20223 (N_20223,N_18188,N_19048);
or U20224 (N_20224,N_16852,N_16410);
and U20225 (N_20225,N_19418,N_17305);
xnor U20226 (N_20226,N_15723,N_19978);
nor U20227 (N_20227,N_18700,N_17187);
nand U20228 (N_20228,N_16455,N_17123);
xnor U20229 (N_20229,N_17761,N_15979);
and U20230 (N_20230,N_16107,N_17726);
xnor U20231 (N_20231,N_15540,N_19784);
and U20232 (N_20232,N_17876,N_18742);
and U20233 (N_20233,N_17322,N_16145);
or U20234 (N_20234,N_18791,N_18789);
or U20235 (N_20235,N_16014,N_15635);
nor U20236 (N_20236,N_17750,N_18232);
and U20237 (N_20237,N_17044,N_19360);
nand U20238 (N_20238,N_17967,N_17548);
and U20239 (N_20239,N_19278,N_18338);
xor U20240 (N_20240,N_19950,N_15914);
nand U20241 (N_20241,N_15741,N_17469);
xnor U20242 (N_20242,N_15971,N_15233);
xor U20243 (N_20243,N_15698,N_19166);
nand U20244 (N_20244,N_19543,N_18708);
xor U20245 (N_20245,N_16741,N_15819);
nor U20246 (N_20246,N_15256,N_17526);
or U20247 (N_20247,N_17963,N_19067);
nor U20248 (N_20248,N_18663,N_17679);
or U20249 (N_20249,N_19373,N_16619);
or U20250 (N_20250,N_16512,N_16937);
or U20251 (N_20251,N_19727,N_15210);
and U20252 (N_20252,N_16829,N_15472);
xnor U20253 (N_20253,N_15365,N_17969);
or U20254 (N_20254,N_19544,N_19635);
or U20255 (N_20255,N_15888,N_15040);
or U20256 (N_20256,N_17831,N_19669);
xnor U20257 (N_20257,N_19375,N_16794);
or U20258 (N_20258,N_19552,N_18304);
nor U20259 (N_20259,N_19926,N_15848);
nand U20260 (N_20260,N_18536,N_16485);
xnor U20261 (N_20261,N_19063,N_18949);
or U20262 (N_20262,N_15695,N_18215);
and U20263 (N_20263,N_16859,N_16379);
or U20264 (N_20264,N_15201,N_18960);
nor U20265 (N_20265,N_15951,N_15508);
xnor U20266 (N_20266,N_17820,N_19676);
nand U20267 (N_20267,N_19404,N_18108);
or U20268 (N_20268,N_15369,N_19205);
or U20269 (N_20269,N_15528,N_19168);
nand U20270 (N_20270,N_19208,N_16167);
nor U20271 (N_20271,N_17629,N_15166);
or U20272 (N_20272,N_19061,N_16766);
nor U20273 (N_20273,N_19966,N_15574);
xnor U20274 (N_20274,N_17403,N_16765);
or U20275 (N_20275,N_17085,N_19530);
and U20276 (N_20276,N_19857,N_19084);
xnor U20277 (N_20277,N_16218,N_15531);
or U20278 (N_20278,N_15064,N_15904);
and U20279 (N_20279,N_17259,N_18522);
and U20280 (N_20280,N_15857,N_15325);
xor U20281 (N_20281,N_15805,N_16093);
xnor U20282 (N_20282,N_15476,N_19125);
and U20283 (N_20283,N_16201,N_16142);
xor U20284 (N_20284,N_17366,N_15037);
or U20285 (N_20285,N_17566,N_19044);
or U20286 (N_20286,N_18111,N_16428);
xnor U20287 (N_20287,N_15866,N_17964);
and U20288 (N_20288,N_15787,N_15419);
or U20289 (N_20289,N_16562,N_18997);
xnor U20290 (N_20290,N_18067,N_16298);
nand U20291 (N_20291,N_15009,N_18886);
nand U20292 (N_20292,N_18081,N_19097);
nand U20293 (N_20293,N_19577,N_19968);
nand U20294 (N_20294,N_15632,N_15222);
nand U20295 (N_20295,N_15469,N_17095);
or U20296 (N_20296,N_15326,N_19562);
xnor U20297 (N_20297,N_18272,N_17647);
nor U20298 (N_20298,N_17827,N_17354);
or U20299 (N_20299,N_17387,N_19283);
and U20300 (N_20300,N_16144,N_19612);
and U20301 (N_20301,N_19210,N_19689);
or U20302 (N_20302,N_16289,N_17764);
nor U20303 (N_20303,N_18358,N_15428);
or U20304 (N_20304,N_17846,N_17977);
and U20305 (N_20305,N_16957,N_17999);
nand U20306 (N_20306,N_19141,N_19911);
and U20307 (N_20307,N_16087,N_15488);
xnor U20308 (N_20308,N_17017,N_15211);
nand U20309 (N_20309,N_16419,N_17909);
nand U20310 (N_20310,N_17781,N_18514);
or U20311 (N_20311,N_18395,N_15909);
or U20312 (N_20312,N_19654,N_17025);
xnor U20313 (N_20313,N_18070,N_18736);
or U20314 (N_20314,N_18714,N_19622);
xnor U20315 (N_20315,N_16236,N_16124);
nor U20316 (N_20316,N_19041,N_18664);
nand U20317 (N_20317,N_18231,N_19406);
nand U20318 (N_20318,N_18940,N_17143);
and U20319 (N_20319,N_16089,N_17076);
and U20320 (N_20320,N_17084,N_16447);
nand U20321 (N_20321,N_17217,N_16955);
xor U20322 (N_20322,N_15162,N_18307);
nand U20323 (N_20323,N_15295,N_15621);
and U20324 (N_20324,N_19377,N_15687);
and U20325 (N_20325,N_15084,N_16187);
xnor U20326 (N_20326,N_15415,N_17830);
nand U20327 (N_20327,N_19571,N_17533);
xor U20328 (N_20328,N_15614,N_16681);
or U20329 (N_20329,N_16028,N_19762);
nor U20330 (N_20330,N_16883,N_18444);
xnor U20331 (N_20331,N_19712,N_18961);
xor U20332 (N_20332,N_17371,N_16257);
nor U20333 (N_20333,N_19550,N_17021);
xor U20334 (N_20334,N_17578,N_19025);
xor U20335 (N_20335,N_16140,N_17329);
nor U20336 (N_20336,N_16889,N_16522);
nor U20337 (N_20337,N_15938,N_16975);
or U20338 (N_20338,N_15153,N_16120);
nand U20339 (N_20339,N_19501,N_17214);
or U20340 (N_20340,N_15172,N_19545);
nand U20341 (N_20341,N_15492,N_17410);
xor U20342 (N_20342,N_17483,N_19217);
xor U20343 (N_20343,N_15102,N_15978);
or U20344 (N_20344,N_17765,N_19456);
and U20345 (N_20345,N_16790,N_17154);
and U20346 (N_20346,N_18711,N_15691);
nor U20347 (N_20347,N_15083,N_17649);
xor U20348 (N_20348,N_16661,N_16101);
or U20349 (N_20349,N_19722,N_19914);
xor U20350 (N_20350,N_15112,N_15389);
or U20351 (N_20351,N_15133,N_17517);
nor U20352 (N_20352,N_15998,N_15839);
and U20353 (N_20353,N_18371,N_17661);
nand U20354 (N_20354,N_16901,N_16019);
or U20355 (N_20355,N_16337,N_16837);
and U20356 (N_20356,N_15581,N_17706);
and U20357 (N_20357,N_16880,N_16247);
nor U20358 (N_20358,N_16530,N_15564);
nand U20359 (N_20359,N_18706,N_18980);
nand U20360 (N_20360,N_15015,N_17774);
nand U20361 (N_20361,N_15593,N_18032);
and U20362 (N_20362,N_16641,N_17793);
nor U20363 (N_20363,N_19139,N_15105);
and U20364 (N_20364,N_16453,N_15590);
xor U20365 (N_20365,N_18244,N_19881);
nor U20366 (N_20366,N_15807,N_17407);
xor U20367 (N_20367,N_15080,N_19703);
nand U20368 (N_20368,N_19551,N_16468);
and U20369 (N_20369,N_18274,N_18320);
xnor U20370 (N_20370,N_16666,N_17603);
nand U20371 (N_20371,N_17158,N_15038);
xor U20372 (N_20372,N_16348,N_15652);
and U20373 (N_20373,N_19399,N_15014);
and U20374 (N_20374,N_15955,N_17065);
or U20375 (N_20375,N_18150,N_18845);
nor U20376 (N_20376,N_18605,N_15364);
xor U20377 (N_20377,N_16094,N_19385);
nand U20378 (N_20378,N_15230,N_17737);
and U20379 (N_20379,N_16882,N_18784);
nor U20380 (N_20380,N_15799,N_16223);
nand U20381 (N_20381,N_16063,N_15526);
nor U20382 (N_20382,N_15946,N_18975);
nor U20383 (N_20383,N_18607,N_19351);
nor U20384 (N_20384,N_16122,N_16336);
or U20385 (N_20385,N_18688,N_15493);
nand U20386 (N_20386,N_17128,N_16671);
or U20387 (N_20387,N_16646,N_17468);
nand U20388 (N_20388,N_15276,N_17870);
or U20389 (N_20389,N_16588,N_16384);
nand U20390 (N_20390,N_16401,N_17621);
nor U20391 (N_20391,N_19806,N_18899);
nand U20392 (N_20392,N_19531,N_19560);
nor U20393 (N_20393,N_18883,N_19255);
or U20394 (N_20394,N_15925,N_18957);
or U20395 (N_20395,N_17917,N_18507);
nor U20396 (N_20396,N_15216,N_17704);
or U20397 (N_20397,N_18228,N_15125);
or U20398 (N_20398,N_15649,N_15020);
nand U20399 (N_20399,N_19221,N_19955);
nand U20400 (N_20400,N_18375,N_15013);
nand U20401 (N_20401,N_15032,N_15719);
or U20402 (N_20402,N_15046,N_15834);
nand U20403 (N_20403,N_17797,N_16287);
xor U20404 (N_20404,N_16043,N_17971);
and U20405 (N_20405,N_16819,N_15279);
nor U20406 (N_20406,N_15069,N_18729);
xor U20407 (N_20407,N_15856,N_16640);
nand U20408 (N_20408,N_18334,N_17082);
xnor U20409 (N_20409,N_15304,N_19587);
nand U20410 (N_20410,N_18740,N_17334);
xor U20411 (N_20411,N_19474,N_16540);
and U20412 (N_20412,N_19638,N_18701);
xnor U20413 (N_20413,N_19743,N_18986);
or U20414 (N_20414,N_15335,N_17722);
nand U20415 (N_20415,N_18048,N_17083);
nor U20416 (N_20416,N_17813,N_18862);
nor U20417 (N_20417,N_17618,N_19862);
or U20418 (N_20418,N_19672,N_16545);
or U20419 (N_20419,N_19593,N_16919);
nor U20420 (N_20420,N_17068,N_18933);
nand U20421 (N_20421,N_16878,N_16263);
or U20422 (N_20422,N_19262,N_15683);
nand U20423 (N_20423,N_18528,N_19930);
nand U20424 (N_20424,N_19415,N_16688);
and U20425 (N_20425,N_17431,N_17799);
and U20426 (N_20426,N_17267,N_16771);
nor U20427 (N_20427,N_17171,N_19737);
and U20428 (N_20428,N_18907,N_15518);
xnor U20429 (N_20429,N_15893,N_18815);
nand U20430 (N_20430,N_17433,N_17420);
nor U20431 (N_20431,N_19425,N_15362);
xor U20432 (N_20432,N_18238,N_19085);
xor U20433 (N_20433,N_15370,N_17607);
and U20434 (N_20434,N_17033,N_15577);
nand U20435 (N_20435,N_15817,N_18945);
or U20436 (N_20436,N_19379,N_15456);
nor U20437 (N_20437,N_17744,N_19332);
nor U20438 (N_20438,N_16351,N_19814);
nor U20439 (N_20439,N_16245,N_16606);
or U20440 (N_20440,N_19256,N_17862);
or U20441 (N_20441,N_16026,N_17292);
xnor U20442 (N_20442,N_17901,N_18347);
nand U20443 (N_20443,N_19014,N_17672);
or U20444 (N_20444,N_16215,N_16222);
or U20445 (N_20445,N_16774,N_18361);
nor U20446 (N_20446,N_17299,N_18824);
xor U20447 (N_20447,N_15840,N_18822);
nor U20448 (N_20448,N_18388,N_15342);
xnor U20449 (N_20449,N_19931,N_18557);
or U20450 (N_20450,N_15425,N_18281);
xor U20451 (N_20451,N_15867,N_17514);
or U20452 (N_20452,N_19591,N_18177);
and U20453 (N_20453,N_16203,N_15302);
nor U20454 (N_20454,N_16420,N_15756);
or U20455 (N_20455,N_16785,N_15413);
or U20456 (N_20456,N_15751,N_19215);
xnor U20457 (N_20457,N_18005,N_18217);
and U20458 (N_20458,N_17720,N_19977);
xor U20459 (N_20459,N_17255,N_17185);
nand U20460 (N_20460,N_16660,N_18830);
nor U20461 (N_20461,N_17683,N_16810);
and U20462 (N_20462,N_19019,N_18775);
or U20463 (N_20463,N_18527,N_18107);
or U20464 (N_20464,N_18474,N_17537);
xnor U20465 (N_20465,N_15721,N_15602);
nand U20466 (N_20466,N_17741,N_19942);
and U20467 (N_20467,N_16021,N_15677);
nand U20468 (N_20468,N_18316,N_16626);
or U20469 (N_20469,N_17480,N_16861);
nand U20470 (N_20470,N_17529,N_15315);
or U20471 (N_20471,N_15976,N_17000);
nand U20472 (N_20472,N_16362,N_15917);
and U20473 (N_20473,N_18223,N_19411);
or U20474 (N_20474,N_17713,N_15989);
nand U20475 (N_20475,N_19159,N_18340);
xnor U20476 (N_20476,N_15464,N_19740);
nor U20477 (N_20477,N_15709,N_18058);
xor U20478 (N_20478,N_16571,N_16584);
nor U20479 (N_20479,N_19428,N_17029);
xor U20480 (N_20480,N_19992,N_17841);
xnor U20481 (N_20481,N_16553,N_17498);
nor U20482 (N_20482,N_16213,N_18524);
nand U20483 (N_20483,N_17794,N_16091);
nor U20484 (N_20484,N_18911,N_19246);
nand U20485 (N_20485,N_18162,N_17333);
or U20486 (N_20486,N_15964,N_15373);
nor U20487 (N_20487,N_15328,N_16160);
xnor U20488 (N_20488,N_17442,N_16372);
or U20489 (N_20489,N_16071,N_18655);
xnor U20490 (N_20490,N_18722,N_16408);
and U20491 (N_20491,N_16333,N_15174);
or U20492 (N_20492,N_16126,N_19288);
and U20493 (N_20493,N_18988,N_19403);
or U20494 (N_20494,N_15354,N_19317);
nand U20495 (N_20495,N_18442,N_16534);
or U20496 (N_20496,N_19362,N_16673);
nor U20497 (N_20497,N_18024,N_15355);
nand U20498 (N_20498,N_18728,N_16519);
and U20499 (N_20499,N_18928,N_17663);
nor U20500 (N_20500,N_15844,N_19223);
and U20501 (N_20501,N_16448,N_18441);
nor U20502 (N_20502,N_16480,N_16635);
xnor U20503 (N_20503,N_16520,N_17397);
and U20504 (N_20504,N_16997,N_19053);
xor U20505 (N_20505,N_19644,N_19609);
or U20506 (N_20506,N_15828,N_15449);
or U20507 (N_20507,N_15086,N_15572);
or U20508 (N_20508,N_18468,N_15674);
nor U20509 (N_20509,N_16020,N_19910);
and U20510 (N_20510,N_15627,N_15999);
or U20511 (N_20511,N_17589,N_17923);
nor U20512 (N_20512,N_15739,N_18932);
nand U20513 (N_20513,N_18534,N_16082);
or U20514 (N_20514,N_17718,N_15483);
nor U20515 (N_20515,N_18895,N_18795);
nand U20516 (N_20516,N_18114,N_19307);
or U20517 (N_20517,N_19580,N_16330);
xnor U20518 (N_20518,N_19269,N_17941);
and U20519 (N_20519,N_17024,N_19570);
and U20520 (N_20520,N_17838,N_18619);
nor U20521 (N_20521,N_16851,N_17912);
and U20522 (N_20522,N_19433,N_19668);
nor U20523 (N_20523,N_15642,N_17369);
nand U20524 (N_20524,N_19876,N_16035);
nand U20525 (N_20525,N_16321,N_16581);
or U20526 (N_20526,N_17008,N_19619);
nor U20527 (N_20527,N_18490,N_18670);
nand U20528 (N_20528,N_17709,N_19675);
xnor U20529 (N_20529,N_17092,N_16320);
and U20530 (N_20530,N_15345,N_15772);
nand U20531 (N_20531,N_15368,N_18915);
xnor U20532 (N_20532,N_15854,N_19236);
and U20533 (N_20533,N_17019,N_17342);
xor U20534 (N_20534,N_15160,N_19495);
nand U20535 (N_20535,N_18273,N_16972);
or U20536 (N_20536,N_19940,N_15482);
nand U20537 (N_20537,N_19202,N_17172);
and U20538 (N_20538,N_19371,N_17543);
or U20539 (N_20539,N_18453,N_15421);
and U20540 (N_20540,N_18247,N_17759);
xor U20541 (N_20541,N_15831,N_18636);
nor U20542 (N_20542,N_17658,N_18401);
xnor U20543 (N_20543,N_19155,N_18996);
or U20544 (N_20544,N_16102,N_15843);
nand U20545 (N_20545,N_17457,N_18938);
nor U20546 (N_20546,N_16993,N_16281);
and U20547 (N_20547,N_15081,N_17063);
nand U20548 (N_20548,N_16238,N_19174);
nor U20549 (N_20549,N_15645,N_19795);
xnor U20550 (N_20550,N_15420,N_15730);
nor U20551 (N_20551,N_15907,N_18650);
or U20552 (N_20552,N_19311,N_19500);
and U20553 (N_20553,N_16796,N_16706);
nand U20554 (N_20554,N_17684,N_16466);
nor U20555 (N_20555,N_19493,N_17221);
nor U20556 (N_20556,N_18952,N_19359);
or U20557 (N_20557,N_17887,N_15737);
or U20558 (N_20558,N_19324,N_16524);
xnor U20559 (N_20559,N_15637,N_15106);
and U20560 (N_20560,N_16157,N_15149);
nand U20561 (N_20561,N_17385,N_17290);
and U20562 (N_20562,N_18012,N_17162);
nand U20563 (N_20563,N_17190,N_19304);
nand U20564 (N_20564,N_16311,N_18912);
and U20565 (N_20565,N_17424,N_16866);
and U20566 (N_20566,N_15594,N_16594);
nor U20567 (N_20567,N_16462,N_16514);
nand U20568 (N_20568,N_19906,N_19507);
xor U20569 (N_20569,N_16268,N_18497);
or U20570 (N_20570,N_17542,N_18112);
and U20571 (N_20571,N_16602,N_15625);
or U20572 (N_20572,N_18175,N_19138);
nor U20573 (N_20573,N_18041,N_19163);
xnor U20574 (N_20574,N_19718,N_15759);
and U20575 (N_20575,N_16529,N_19802);
and U20576 (N_20576,N_16024,N_17555);
xnor U20577 (N_20577,N_15441,N_15514);
nor U20578 (N_20578,N_15261,N_19666);
nor U20579 (N_20579,N_17560,N_16467);
nor U20580 (N_20580,N_16703,N_19329);
or U20581 (N_20581,N_15716,N_17446);
nor U20582 (N_20582,N_18852,N_16678);
xnor U20583 (N_20583,N_18681,N_18021);
or U20584 (N_20584,N_15875,N_19382);
or U20585 (N_20585,N_15314,N_19331);
xnor U20586 (N_20586,N_18298,N_18314);
and U20587 (N_20587,N_19107,N_16069);
or U20588 (N_20588,N_17022,N_15458);
nand U20589 (N_20589,N_15382,N_15825);
nand U20590 (N_20590,N_18324,N_19913);
xnor U20591 (N_20591,N_17805,N_17736);
nand U20592 (N_20592,N_17031,N_18097);
or U20593 (N_20593,N_18500,N_19354);
nand U20594 (N_20594,N_18588,N_19999);
nor U20595 (N_20595,N_19637,N_17985);
nor U20596 (N_20596,N_18682,N_18978);
nand U20597 (N_20597,N_15073,N_18146);
or U20598 (N_20598,N_17182,N_16885);
and U20599 (N_20599,N_18078,N_18475);
nand U20600 (N_20600,N_17637,N_17995);
nor U20601 (N_20601,N_18762,N_17102);
xnor U20602 (N_20602,N_17763,N_17863);
nor U20603 (N_20603,N_15242,N_17742);
and U20604 (N_20604,N_17974,N_19338);
nor U20605 (N_20605,N_19866,N_19022);
and U20606 (N_20606,N_15457,N_17540);
nor U20607 (N_20607,N_19590,N_19528);
nor U20608 (N_20608,N_15079,N_16070);
and U20609 (N_20609,N_18707,N_18543);
nand U20610 (N_20610,N_19834,N_17845);
nand U20611 (N_20611,N_19453,N_15609);
nor U20612 (N_20612,N_16610,N_16129);
xnor U20613 (N_20613,N_15118,N_16172);
nor U20614 (N_20614,N_19043,N_19929);
nor U20615 (N_20615,N_18153,N_15045);
nor U20616 (N_20616,N_17860,N_16072);
nand U20617 (N_20617,N_17743,N_16871);
nand U20618 (N_20618,N_19102,N_19467);
nor U20619 (N_20619,N_18727,N_16017);
or U20620 (N_20620,N_16647,N_15922);
or U20621 (N_20621,N_15808,N_19594);
and U20622 (N_20622,N_17568,N_19280);
nor U20623 (N_20623,N_19951,N_16658);
xnor U20624 (N_20624,N_17996,N_17572);
and U20625 (N_20625,N_16251,N_19129);
and U20626 (N_20626,N_19586,N_18383);
nand U20627 (N_20627,N_18587,N_18343);
or U20628 (N_20628,N_15580,N_18758);
xor U20629 (N_20629,N_16373,N_18119);
nand U20630 (N_20630,N_16381,N_17124);
nor U20631 (N_20631,N_19219,N_19049);
nand U20632 (N_20632,N_17579,N_18440);
and U20633 (N_20633,N_15688,N_18626);
or U20634 (N_20634,N_19312,N_17350);
nand U20635 (N_20635,N_19176,N_16841);
or U20636 (N_20636,N_15936,N_15569);
or U20637 (N_20637,N_16099,N_19869);
or U20638 (N_20638,N_16518,N_19413);
nand U20639 (N_20639,N_18551,N_19981);
or U20640 (N_20640,N_18368,N_17405);
and U20641 (N_20641,N_18176,N_17164);
nor U20642 (N_20642,N_19018,N_16114);
xor U20643 (N_20643,N_15292,N_15277);
xor U20644 (N_20644,N_17900,N_19321);
xor U20645 (N_20645,N_15859,N_18152);
xor U20646 (N_20646,N_17558,N_18843);
and U20647 (N_20647,N_18686,N_16403);
nor U20648 (N_20648,N_15156,N_17202);
or U20649 (N_20649,N_17511,N_19768);
nor U20650 (N_20650,N_16985,N_19191);
and U20651 (N_20651,N_18885,N_19282);
xnor U20652 (N_20652,N_16358,N_19766);
or U20653 (N_20653,N_15416,N_15129);
or U20654 (N_20654,N_16740,N_15654);
xnor U20655 (N_20655,N_19088,N_17792);
nor U20656 (N_20656,N_19794,N_15062);
or U20657 (N_20657,N_18449,N_16935);
and U20658 (N_20658,N_15722,N_19234);
and U20659 (N_20659,N_15475,N_19831);
nor U20660 (N_20660,N_19887,N_16081);
and U20661 (N_20661,N_15108,N_17976);
and U20662 (N_20662,N_16152,N_19807);
nand U20663 (N_20663,N_15317,N_15552);
nor U20664 (N_20664,N_18234,N_18488);
nor U20665 (N_20665,N_19508,N_17373);
xnor U20666 (N_20666,N_17282,N_17199);
or U20667 (N_20667,N_15532,N_19148);
xor U20668 (N_20668,N_16188,N_16476);
xnor U20669 (N_20669,N_17059,N_19209);
and U20670 (N_20670,N_17352,N_15110);
nor U20671 (N_20671,N_19738,N_19736);
nor U20672 (N_20672,N_15331,N_19422);
xor U20673 (N_20673,N_16596,N_17278);
nand U20674 (N_20674,N_16770,N_15868);
or U20675 (N_20675,N_17899,N_16252);
or U20676 (N_20676,N_16367,N_16801);
xor U20677 (N_20677,N_17959,N_18826);
and U20678 (N_20678,N_15170,N_18237);
and U20679 (N_20679,N_16583,N_16618);
nor U20680 (N_20680,N_17049,N_15664);
or U20681 (N_20681,N_16915,N_19402);
nor U20682 (N_20682,N_19751,N_18617);
nor U20683 (N_20683,N_18446,N_17416);
nor U20684 (N_20684,N_15720,N_15615);
xor U20685 (N_20685,N_15308,N_18130);
xnor U20686 (N_20686,N_17628,N_17114);
nor U20687 (N_20687,N_16578,N_15184);
or U20688 (N_20688,N_19878,N_16614);
nor U20689 (N_20689,N_19378,N_17140);
nor U20690 (N_20690,N_19733,N_18896);
xnor U20691 (N_20691,N_16686,N_17698);
nand U20692 (N_20692,N_16624,N_19894);
xor U20693 (N_20693,N_19924,N_17465);
xnor U20694 (N_20694,N_15696,N_16924);
or U20695 (N_20695,N_16922,N_15094);
xnor U20696 (N_20696,N_17283,N_15272);
xor U20697 (N_20697,N_17266,N_15634);
nor U20698 (N_20698,N_17994,N_18101);
or U20699 (N_20699,N_16692,N_19441);
nand U20700 (N_20700,N_15071,N_19030);
nor U20701 (N_20701,N_17748,N_19901);
or U20702 (N_20702,N_19785,N_17108);
and U20703 (N_20703,N_18818,N_17206);
and U20704 (N_20704,N_17330,N_19828);
nand U20705 (N_20705,N_19242,N_15330);
nor U20706 (N_20706,N_19078,N_17866);
nor U20707 (N_20707,N_18897,N_19961);
xor U20708 (N_20708,N_16950,N_15950);
or U20709 (N_20709,N_18489,N_19557);
nand U20710 (N_20710,N_15244,N_18849);
and U20711 (N_20711,N_17073,N_19854);
and U20712 (N_20712,N_19002,N_17495);
nand U20713 (N_20713,N_17988,N_17438);
xor U20714 (N_20714,N_16789,N_18642);
nand U20715 (N_20715,N_15098,N_19631);
xnor U20716 (N_20716,N_17236,N_17473);
nor U20717 (N_20717,N_15985,N_15981);
nor U20718 (N_20718,N_16833,N_16487);
nand U20719 (N_20719,N_16402,N_16181);
xor U20720 (N_20720,N_18136,N_17818);
or U20721 (N_20721,N_17509,N_16005);
nand U20722 (N_20722,N_18491,N_16776);
or U20723 (N_20723,N_19749,N_17471);
nand U20724 (N_20724,N_15851,N_19599);
or U20725 (N_20725,N_15522,N_18185);
and U20726 (N_20726,N_18898,N_15240);
xor U20727 (N_20727,N_19521,N_18693);
and U20728 (N_20728,N_16032,N_19135);
nor U20729 (N_20729,N_19386,N_15378);
nor U20730 (N_20730,N_19258,N_17189);
or U20731 (N_20731,N_19540,N_15407);
nand U20732 (N_20732,N_18486,N_15711);
or U20733 (N_20733,N_19469,N_15021);
nor U20734 (N_20734,N_15749,N_16303);
xnor U20735 (N_20735,N_18183,N_17051);
and U20736 (N_20736,N_19923,N_17847);
or U20737 (N_20737,N_17272,N_19080);
or U20738 (N_20738,N_19170,N_19996);
xnor U20739 (N_20739,N_16643,N_15554);
and U20740 (N_20740,N_18943,N_17328);
and U20741 (N_20741,N_17358,N_18769);
xor U20742 (N_20742,N_18249,N_15417);
xnor U20743 (N_20743,N_18967,N_16217);
and U20744 (N_20744,N_18926,N_18819);
and U20745 (N_20745,N_16426,N_16329);
xnor U20746 (N_20746,N_16016,N_19896);
xor U20747 (N_20747,N_19917,N_19648);
nand U20748 (N_20748,N_18425,N_18336);
nor U20749 (N_20749,N_18792,N_16895);
xor U20750 (N_20750,N_19546,N_17109);
nand U20751 (N_20751,N_17569,N_17979);
and U20752 (N_20752,N_19578,N_19937);
nand U20753 (N_20753,N_19443,N_17740);
xor U20754 (N_20754,N_15322,N_17636);
or U20755 (N_20755,N_19897,N_17598);
nor U20756 (N_20756,N_16314,N_18335);
xor U20757 (N_20757,N_15550,N_18017);
or U20758 (N_20758,N_19734,N_18121);
nand U20759 (N_20759,N_18604,N_18282);
nand U20760 (N_20760,N_15078,N_18060);
and U20761 (N_20761,N_19778,N_16095);
nand U20762 (N_20762,N_17311,N_15048);
xor U20763 (N_20763,N_16103,N_15658);
nand U20764 (N_20764,N_16123,N_16812);
nor U20765 (N_20765,N_16344,N_18799);
and U20766 (N_20766,N_19670,N_16515);
nor U20767 (N_20767,N_16185,N_15366);
or U20768 (N_20768,N_18417,N_18285);
or U20769 (N_20769,N_16675,N_18311);
and U20770 (N_20770,N_19195,N_16214);
nor U20771 (N_20771,N_19840,N_19212);
nor U20772 (N_20772,N_16511,N_18509);
xor U20773 (N_20773,N_19885,N_15093);
and U20774 (N_20774,N_19533,N_17432);
nand U20775 (N_20775,N_18985,N_16727);
xnor U20776 (N_20776,N_18243,N_16084);
xor U20777 (N_20777,N_16921,N_18438);
xor U20778 (N_20778,N_16054,N_18254);
nand U20779 (N_20779,N_18616,N_16450);
and U20780 (N_20780,N_17623,N_16693);
nand U20781 (N_20781,N_16405,N_16754);
xnor U20782 (N_20782,N_16434,N_16128);
nand U20783 (N_20783,N_17832,N_19880);
and U20784 (N_20784,N_15063,N_18829);
or U20785 (N_20785,N_16322,N_19098);
or U20786 (N_20786,N_18106,N_18741);
xnor U20787 (N_20787,N_18637,N_17200);
or U20788 (N_20788,N_15991,N_16756);
nor U20789 (N_20789,N_19848,N_19142);
or U20790 (N_20790,N_19087,N_16777);
nor U20791 (N_20791,N_18155,N_18154);
and U20792 (N_20792,N_15283,N_18516);
xnor U20793 (N_20793,N_19864,N_15150);
xnor U20794 (N_20794,N_15928,N_16456);
or U20795 (N_20795,N_18622,N_16265);
nor U20796 (N_20796,N_15089,N_19250);
nand U20797 (N_20797,N_17141,N_15712);
nand U20798 (N_20798,N_19099,N_18673);
or U20799 (N_20799,N_15423,N_19921);
nand U20800 (N_20800,N_17091,N_15912);
nor U20801 (N_20801,N_17581,N_16780);
xnor U20802 (N_20802,N_17630,N_16067);
and U20803 (N_20803,N_15841,N_17379);
nand U20804 (N_20804,N_16735,N_19364);
nand U20805 (N_20805,N_19459,N_17515);
or U20806 (N_20806,N_17997,N_16987);
nand U20807 (N_20807,N_17522,N_17749);
and U20808 (N_20808,N_15512,N_16749);
nor U20809 (N_20809,N_16556,N_18880);
or U20810 (N_20810,N_15801,N_15744);
nand U20811 (N_20811,N_16432,N_16205);
and U20812 (N_20812,N_19641,N_19437);
nor U20813 (N_20813,N_17531,N_16509);
xnor U20814 (N_20814,N_15099,N_18648);
and U20815 (N_20815,N_15797,N_16546);
and U20816 (N_20816,N_16962,N_19393);
nand U20817 (N_20817,N_15760,N_16056);
nand U20818 (N_20818,N_19847,N_15996);
nor U20819 (N_20819,N_15393,N_16818);
xor U20820 (N_20820,N_16847,N_18568);
or U20821 (N_20821,N_17198,N_17507);
or U20822 (N_20822,N_16105,N_18194);
or U20823 (N_20823,N_19994,N_16791);
xor U20824 (N_20824,N_16865,N_18160);
and U20825 (N_20825,N_19688,N_17281);
nor U20826 (N_20826,N_16537,N_19023);
and U20827 (N_20827,N_16808,N_16758);
xnor U20828 (N_20828,N_18381,N_19352);
or U20829 (N_20829,N_15789,N_19450);
or U20830 (N_20830,N_18946,N_19697);
nand U20831 (N_20831,N_19956,N_16707);
nor U20832 (N_20832,N_19798,N_19919);
nand U20833 (N_20833,N_15408,N_18075);
nor U20834 (N_20834,N_16130,N_19796);
nand U20835 (N_20835,N_19859,N_16709);
xnor U20836 (N_20836,N_16457,N_19891);
or U20837 (N_20837,N_17325,N_19390);
nor U20838 (N_20838,N_19630,N_18589);
and U20839 (N_20839,N_19199,N_19991);
nand U20840 (N_20840,N_18350,N_17673);
or U20841 (N_20841,N_16046,N_16361);
nor U20842 (N_20842,N_18976,N_19384);
xnor U20843 (N_20843,N_18611,N_15019);
nor U20844 (N_20844,N_17908,N_16831);
or U20845 (N_20845,N_19690,N_18501);
and U20846 (N_20846,N_17273,N_19623);
and U20847 (N_20847,N_16654,N_18657);
nand U20848 (N_20848,N_15734,N_18881);
xor U20849 (N_20849,N_19485,N_18454);
nand U20850 (N_20850,N_16676,N_15000);
xor U20851 (N_20851,N_15017,N_16958);
xor U20852 (N_20852,N_18569,N_15123);
xor U20853 (N_20853,N_17245,N_16424);
nor U20854 (N_20854,N_17989,N_15494);
nand U20855 (N_20855,N_18414,N_18131);
nand U20856 (N_20856,N_16267,N_17237);
nand U20857 (N_20857,N_17539,N_18610);
xor U20858 (N_20858,N_19592,N_16283);
xnor U20859 (N_20859,N_16620,N_19513);
nor U20860 (N_20860,N_18660,N_19429);
nand U20861 (N_20861,N_16234,N_18038);
or U20862 (N_20862,N_18613,N_16868);
or U20863 (N_20863,N_16200,N_18566);
and U20864 (N_20864,N_16952,N_15096);
xor U20865 (N_20865,N_19435,N_16404);
and U20866 (N_20866,N_18717,N_17650);
nor U20867 (N_20867,N_18332,N_15249);
nand U20868 (N_20868,N_17317,N_17345);
and U20869 (N_20869,N_19457,N_16049);
xnor U20870 (N_20870,N_19889,N_16151);
or U20871 (N_20871,N_19188,N_15714);
or U20872 (N_20872,N_17788,N_17739);
or U20873 (N_20873,N_15752,N_18023);
nor U20874 (N_20874,N_19092,N_18386);
and U20875 (N_20875,N_17875,N_18964);
and U20876 (N_20876,N_18652,N_17099);
nand U20877 (N_20877,N_18313,N_15132);
nand U20878 (N_20878,N_19713,N_16631);
or U20879 (N_20879,N_16416,N_16585);
nand U20880 (N_20880,N_19251,N_18948);
or U20881 (N_20881,N_15268,N_16629);
and U20882 (N_20882,N_17056,N_18903);
nor U20883 (N_20883,N_17993,N_19072);
nor U20884 (N_20884,N_15847,N_18537);
or U20885 (N_20885,N_16938,N_19497);
or U20886 (N_20886,N_18837,N_18286);
nor U20887 (N_20887,N_17222,N_16806);
or U20888 (N_20888,N_17738,N_15390);
or U20889 (N_20889,N_18410,N_18404);
or U20890 (N_20890,N_18480,N_16459);
nor U20891 (N_20891,N_19819,N_18892);
xnor U20892 (N_20892,N_16797,N_19909);
xnor U20893 (N_20893,N_15729,N_17640);
nand U20894 (N_20894,N_16077,N_15138);
xnor U20895 (N_20895,N_19127,N_19953);
nand U20896 (N_20896,N_19829,N_18656);
xnor U20897 (N_20897,N_18170,N_17745);
nand U20898 (N_20898,N_16132,N_18085);
nor U20899 (N_20899,N_18702,N_18990);
and U20900 (N_20900,N_17181,N_16953);
and U20901 (N_20901,N_17872,N_18439);
nand U20902 (N_20902,N_15830,N_16607);
or U20903 (N_20903,N_17850,N_18257);
or U20904 (N_20904,N_16746,N_17157);
or U20905 (N_20905,N_18698,N_18631);
xor U20906 (N_20906,N_19157,N_15323);
nor U20907 (N_20907,N_19770,N_18515);
xor U20908 (N_20908,N_16932,N_19731);
nor U20909 (N_20909,N_15346,N_17361);
and U20910 (N_20910,N_15736,N_17942);
xnor U20911 (N_20911,N_17053,N_19853);
nor U20912 (N_20912,N_17326,N_17665);
and U20913 (N_20913,N_18430,N_18069);
and U20914 (N_20914,N_15745,N_19774);
nand U20915 (N_20915,N_18591,N_18921);
nand U20916 (N_20916,N_17978,N_16127);
nand U20917 (N_20917,N_19430,N_19813);
or U20918 (N_20918,N_19710,N_18987);
nand U20919 (N_20919,N_16696,N_15519);
nand U20920 (N_20920,N_15117,N_18694);
or U20921 (N_20921,N_18733,N_18206);
xnor U20922 (N_20922,N_17176,N_15489);
nor U20923 (N_20923,N_19473,N_17018);
nor U20924 (N_20924,N_18893,N_18971);
nor U20925 (N_20925,N_18128,N_18325);
or U20926 (N_20926,N_17898,N_16052);
or U20927 (N_20927,N_15316,N_16899);
or U20928 (N_20928,N_17634,N_16171);
nand U20929 (N_20929,N_19319,N_15375);
xor U20930 (N_20930,N_17936,N_17258);
and U20931 (N_20931,N_16363,N_19682);
nand U20932 (N_20932,N_18868,N_17577);
or U20933 (N_20933,N_16282,N_17608);
xor U20934 (N_20934,N_16394,N_15442);
or U20935 (N_20935,N_18265,N_18374);
and U20936 (N_20936,N_18367,N_18745);
nor U20937 (N_20937,N_17254,N_17484);
nand U20938 (N_20938,N_15718,N_16574);
or U20939 (N_20939,N_15027,N_17344);
nor U20940 (N_20940,N_16601,N_16325);
nand U20941 (N_20941,N_17346,N_16042);
xnor U20942 (N_20942,N_19502,N_16034);
and U20943 (N_20943,N_18084,N_15993);
nand U20944 (N_20944,N_18910,N_15056);
nor U20945 (N_20945,N_19316,N_15766);
xor U20946 (N_20946,N_18459,N_17409);
or U20947 (N_20947,N_15974,N_15529);
xor U20948 (N_20948,N_16603,N_18210);
nand U20949 (N_20949,N_17117,N_15969);
xor U20950 (N_20950,N_16820,N_18598);
nand U20951 (N_20951,N_17388,N_17541);
and U20952 (N_20952,N_16458,N_16411);
xor U20953 (N_20953,N_17670,N_18011);
nor U20954 (N_20954,N_15380,N_19786);
nor U20955 (N_20955,N_16443,N_17150);
and U20956 (N_20956,N_17510,N_17130);
and U20957 (N_20957,N_18222,N_18073);
nor U20958 (N_20958,N_16576,N_15740);
or U20959 (N_20959,N_15596,N_15499);
and U20960 (N_20960,N_19588,N_17624);
and U20961 (N_20961,N_18359,N_18362);
nor U20962 (N_20962,N_18665,N_15541);
nor U20963 (N_20963,N_17032,N_16136);
xnor U20964 (N_20964,N_17654,N_16813);
nand U20965 (N_20965,N_17115,N_16825);
and U20966 (N_20966,N_18778,N_16814);
nand U20967 (N_20967,N_16481,N_15057);
xnor U20968 (N_20968,N_16843,N_17575);
or U20969 (N_20969,N_15218,N_15463);
nand U20970 (N_20970,N_18276,N_19972);
nand U20971 (N_20971,N_16340,N_19556);
and U20972 (N_20972,N_18731,N_17148);
or U20973 (N_20973,N_16942,N_17981);
or U20974 (N_20974,N_19065,N_19518);
nor U20975 (N_20975,N_19549,N_16174);
or U20976 (N_20976,N_18137,N_19595);
nor U20977 (N_20977,N_16951,N_18261);
xnor U20978 (N_20978,N_18134,N_15439);
nand U20979 (N_20979,N_16225,N_15746);
nand U20980 (N_20980,N_19498,N_19653);
or U20981 (N_20981,N_17710,N_18120);
nand U20982 (N_20982,N_19220,N_15405);
and U20983 (N_20983,N_17573,N_19468);
xor U20984 (N_20984,N_17478,N_17873);
and U20985 (N_20985,N_17243,N_18260);
nor U20986 (N_20986,N_18396,N_16296);
nand U20987 (N_20987,N_19843,N_15612);
or U20988 (N_20988,N_15948,N_17499);
nor U20989 (N_20989,N_16352,N_19471);
and U20990 (N_20990,N_16243,N_15436);
and U20991 (N_20991,N_17952,N_19939);
xor U20992 (N_20992,N_15821,N_16665);
or U20993 (N_20993,N_15667,N_17757);
xor U20994 (N_20994,N_16726,N_15142);
xor U20995 (N_20995,N_15930,N_17103);
nand U20996 (N_20996,N_18250,N_18118);
nand U20997 (N_20997,N_17079,N_19289);
or U20998 (N_20998,N_15284,N_18192);
xnor U20999 (N_20999,N_15584,N_17520);
or U21000 (N_21000,N_19755,N_15199);
xnor U21001 (N_21001,N_18090,N_15387);
nor U21002 (N_21002,N_15742,N_16659);
and U21003 (N_21003,N_17351,N_15406);
xnor U21004 (N_21004,N_19290,N_16318);
or U21005 (N_21005,N_18297,N_19506);
xnor U21006 (N_21006,N_15795,N_15970);
nor U21007 (N_21007,N_16544,N_17747);
nand U21008 (N_21008,N_18699,N_18034);
nor U21009 (N_21009,N_19758,N_15853);
or U21010 (N_21010,N_18526,N_17796);
and U21011 (N_21011,N_19741,N_19336);
and U21012 (N_21012,N_17300,N_18801);
xor U21013 (N_21013,N_19511,N_17037);
xor U21014 (N_21014,N_17472,N_19721);
xor U21015 (N_21015,N_17843,N_16003);
and U21016 (N_21016,N_17913,N_18394);
or U21017 (N_21017,N_19720,N_18035);
nor U21018 (N_21018,N_18759,N_17659);
xnor U21019 (N_21019,N_17613,N_18970);
and U21020 (N_21020,N_16946,N_15903);
or U21021 (N_21021,N_19106,N_15598);
xor U21022 (N_21022,N_17034,N_17865);
xor U21023 (N_21023,N_19643,N_15497);
or U21024 (N_21024,N_18220,N_19152);
nor U21025 (N_21025,N_18529,N_15270);
xor U21026 (N_21026,N_16926,N_18457);
and U21027 (N_21027,N_17702,N_16566);
or U21028 (N_21028,N_15791,N_16723);
nand U21029 (N_21029,N_16612,N_15101);
or U21030 (N_21030,N_18578,N_16697);
nor U21031 (N_21031,N_18342,N_15761);
nand U21032 (N_21032,N_16712,N_15902);
and U21033 (N_21033,N_17570,N_19193);
and U21034 (N_21034,N_15919,N_16486);
and U21035 (N_21035,N_16664,N_16772);
nor U21036 (N_21036,N_16328,N_16902);
nor U21037 (N_21037,N_15259,N_18001);
or U21038 (N_21038,N_16633,N_19803);
xnor U21039 (N_21039,N_15385,N_18816);
xnor U21040 (N_21040,N_16115,N_19241);
nand U21041 (N_21041,N_19101,N_17691);
nand U21042 (N_21042,N_18634,N_18982);
or U21043 (N_21043,N_16284,N_19007);
nand U21044 (N_21044,N_19013,N_18263);
or U21045 (N_21045,N_15849,N_16536);
and U21046 (N_21046,N_18661,N_15200);
xor U21047 (N_21047,N_19464,N_15185);
nor U21048 (N_21048,N_17606,N_19754);
nand U21049 (N_21049,N_16227,N_17452);
and U21050 (N_21050,N_19004,N_18434);
nand U21051 (N_21051,N_17497,N_19313);
and U21052 (N_21052,N_16523,N_17447);
xnor U21053 (N_21053,N_19294,N_18556);
and U21054 (N_21054,N_16872,N_18853);
and U21055 (N_21055,N_18080,N_18544);
and U21056 (N_21056,N_16316,N_18805);
nand U21057 (N_21057,N_16389,N_17940);
xor U21058 (N_21058,N_16098,N_17252);
nor U21059 (N_21059,N_17926,N_17664);
xor U21060 (N_21060,N_16884,N_19303);
nand U21061 (N_21061,N_17812,N_16914);
or U21062 (N_21062,N_15183,N_18553);
xor U21063 (N_21063,N_16460,N_18241);
nor U21064 (N_21064,N_15363,N_15029);
xnor U21065 (N_21065,N_16048,N_19877);
and U21066 (N_21066,N_19948,N_15173);
nor U21067 (N_21067,N_18780,N_16210);
xor U21068 (N_21068,N_15527,N_19618);
nor U21069 (N_21069,N_18833,N_17893);
xor U21070 (N_21070,N_16961,N_19804);
nor U21071 (N_21071,N_16994,N_16360);
nor U21072 (N_21072,N_17393,N_19198);
nor U21073 (N_21073,N_15384,N_15591);
xnor U21074 (N_21074,N_15576,N_17882);
or U21075 (N_21075,N_18811,N_16826);
and U21076 (N_21076,N_17277,N_19553);
nor U21077 (N_21077,N_17209,N_17894);
nor U21078 (N_21078,N_19395,N_17879);
nand U21079 (N_21079,N_19327,N_16930);
xor U21080 (N_21080,N_17355,N_19213);
nand U21081 (N_21081,N_15780,N_16153);
xor U21082 (N_21082,N_18755,N_16248);
xnor U21083 (N_21083,N_16079,N_18995);
or U21084 (N_21084,N_17968,N_17822);
nor U21085 (N_21085,N_15050,N_18117);
or U21086 (N_21086,N_17586,N_19264);
and U21087 (N_21087,N_17973,N_19691);
nand U21088 (N_21088,N_17688,N_15074);
nor U21089 (N_21089,N_15769,N_16413);
nor U21090 (N_21090,N_19760,N_15329);
xnor U21091 (N_21091,N_17983,N_18575);
and U21092 (N_21092,N_17039,N_18674);
or U21093 (N_21093,N_16637,N_17119);
and U21094 (N_21094,N_19717,N_19822);
and U21095 (N_21095,N_16714,N_16108);
or U21096 (N_21096,N_15517,N_19748);
nor U21097 (N_21097,N_19694,N_18647);
or U21098 (N_21098,N_16751,N_15440);
xor U21099 (N_21099,N_17953,N_18549);
nor U21100 (N_21100,N_16778,N_19621);
xor U21101 (N_21101,N_15700,N_15430);
nand U21102 (N_21102,N_15715,N_16350);
xor U21103 (N_21103,N_15179,N_19118);
or U21104 (N_21104,N_17481,N_19686);
or U21105 (N_21105,N_18047,N_15643);
nand U21106 (N_21106,N_15618,N_19763);
nand U21107 (N_21107,N_16593,N_16541);
and U21108 (N_21108,N_19093,N_15796);
or U21109 (N_21109,N_19852,N_18129);
xnor U21110 (N_21110,N_18638,N_19062);
nor U21111 (N_21111,N_15391,N_19927);
nor U21112 (N_21112,N_15813,N_15725);
nand U21113 (N_21113,N_15359,N_16125);
nor U21114 (N_21114,N_16906,N_17563);
and U21115 (N_21115,N_16449,N_19260);
nor U21116 (N_21116,N_18493,N_17559);
and U21117 (N_21117,N_16141,N_15555);
and U21118 (N_21118,N_15748,N_18171);
nand U21119 (N_21119,N_19325,N_17213);
nor U21120 (N_21120,N_16423,N_16554);
or U21121 (N_21121,N_15135,N_18186);
or U21122 (N_21122,N_17689,N_19350);
xnor U21123 (N_21123,N_15273,N_17724);
and U21124 (N_21124,N_18936,N_16274);
xor U21125 (N_21125,N_17655,N_16053);
nor U21126 (N_21126,N_17837,N_19606);
xnor U21127 (N_21127,N_16807,N_18739);
nand U21128 (N_21128,N_17353,N_18225);
or U21129 (N_21129,N_19308,N_16504);
nor U21130 (N_21130,N_16970,N_15543);
nand U21131 (N_21131,N_16811,N_16431);
nand U21132 (N_21132,N_19861,N_19218);
or U21133 (N_21133,N_17064,N_15243);
or U21134 (N_21134,N_18766,N_19873);
nor U21135 (N_21135,N_18614,N_17151);
nand U21136 (N_21136,N_16580,N_17421);
and U21137 (N_21137,N_19564,N_18969);
or U21138 (N_21138,N_18255,N_18180);
nor U21139 (N_21139,N_16879,N_15303);
xor U21140 (N_21140,N_15100,N_17809);
and U21141 (N_21141,N_17435,N_19216);
xnor U21142 (N_21142,N_17233,N_18562);
xnor U21143 (N_21143,N_17614,N_17619);
nand U21144 (N_21144,N_15412,N_17552);
and U21145 (N_21145,N_16338,N_19488);
xor U21146 (N_21146,N_19009,N_16538);
nor U21147 (N_21147,N_15959,N_16324);
xor U21148 (N_21148,N_16731,N_16104);
xor U21149 (N_21149,N_17104,N_18927);
and U21150 (N_21150,N_16779,N_16651);
nor U21151 (N_21151,N_17732,N_17077);
or U21152 (N_21152,N_16656,N_15686);
xor U21153 (N_21153,N_17676,N_18753);
and U21154 (N_21154,N_16030,N_15109);
xor U21155 (N_21155,N_17551,N_16645);
or U21156 (N_21156,N_19783,N_17521);
and U21157 (N_21157,N_18166,N_16648);
or U21158 (N_21158,N_17886,N_19103);
or U21159 (N_21159,N_17884,N_19971);
or U21160 (N_21160,N_16288,N_18473);
nor U21161 (N_21161,N_17412,N_16204);
nand U21162 (N_21162,N_16277,N_19517);
or U21163 (N_21163,N_18074,N_19936);
xor U21164 (N_21164,N_19108,N_16510);
and U21165 (N_21165,N_15321,N_18296);
and U21166 (N_21166,N_19860,N_17932);
nand U21167 (N_21167,N_19089,N_17284);
xnor U21168 (N_21168,N_18666,N_19120);
and U21169 (N_21169,N_16934,N_17549);
nand U21170 (N_21170,N_18331,N_15865);
xnor U21171 (N_21171,N_17523,N_18003);
nor U21172 (N_21172,N_16356,N_15294);
nor U21173 (N_21173,N_17380,N_19509);
nor U21174 (N_21174,N_19012,N_16567);
and U21175 (N_21175,N_15923,N_19366);
xor U21176 (N_21176,N_16787,N_19844);
nand U21177 (N_21177,N_15535,N_19514);
nand U21178 (N_21178,N_19486,N_18370);
xnor U21179 (N_21179,N_16133,N_19772);
and U21180 (N_21180,N_15913,N_16346);
nand U21181 (N_21181,N_19673,N_16393);
and U21182 (N_21182,N_18810,N_15758);
nor U21183 (N_21183,N_18328,N_19349);
or U21184 (N_21184,N_18472,N_18447);
or U21185 (N_21185,N_16854,N_15608);
nand U21186 (N_21186,N_18082,N_19086);
nand U21187 (N_21187,N_17987,N_19867);
and U21188 (N_21188,N_16835,N_18705);
nand U21189 (N_21189,N_18794,N_18037);
or U21190 (N_21190,N_18303,N_15792);
and U21191 (N_21191,N_15633,N_18869);
nand U21192 (N_21192,N_16701,N_19671);
and U21193 (N_21193,N_16415,N_16399);
xor U21194 (N_21194,N_17565,N_17674);
xor U21195 (N_21195,N_15226,N_15327);
nand U21196 (N_21196,N_15611,N_19879);
nor U21197 (N_21197,N_18322,N_15163);
and U21198 (N_21198,N_16644,N_17828);
and U21199 (N_21199,N_19839,N_19408);
or U21200 (N_21200,N_18574,N_18419);
and U21201 (N_21201,N_19414,N_17666);
nand U21202 (N_21202,N_16669,N_15134);
nor U21203 (N_21203,N_17795,N_18168);
nor U21204 (N_21204,N_16355,N_16390);
and U21205 (N_21205,N_18064,N_15886);
nor U21206 (N_21206,N_15566,N_19235);
and U21207 (N_21207,N_15622,N_15887);
or U21208 (N_21208,N_15977,N_17770);
or U21209 (N_21209,N_18463,N_16725);
and U21210 (N_21210,N_16551,N_16179);
or U21211 (N_21211,N_15300,N_15648);
nand U21212 (N_21212,N_16795,N_16974);
and U21213 (N_21213,N_19496,N_16715);
xnor U21214 (N_21214,N_18972,N_16760);
or U21215 (N_21215,N_15647,N_18218);
nand U21216 (N_21216,N_18184,N_19539);
nor U21217 (N_21217,N_18264,N_18994);
nor U21218 (N_21218,N_15338,N_19692);
and U21219 (N_21219,N_15239,N_16041);
and U21220 (N_21220,N_16183,N_17980);
or U21221 (N_21221,N_18712,N_19983);
nand U21222 (N_21222,N_18420,N_16058);
nor U21223 (N_21223,N_15901,N_15704);
and U21224 (N_21224,N_17878,N_18485);
or U21225 (N_21225,N_18963,N_15773);
nand U21226 (N_21226,N_19837,N_18197);
or U21227 (N_21227,N_17582,N_18028);
nor U21228 (N_21228,N_15767,N_15829);
xnor U21229 (N_21229,N_16897,N_16739);
nand U21230 (N_21230,N_18864,N_15646);
xor U21231 (N_21231,N_18283,N_15251);
nor U21232 (N_21232,N_16143,N_17918);
xor U21233 (N_21233,N_17836,N_15803);
xor U21234 (N_21234,N_18224,N_18863);
xor U21235 (N_21235,N_17907,N_19597);
and U21236 (N_21236,N_18510,N_18608);
xor U21237 (N_21237,N_19566,N_19410);
nand U21238 (N_21238,N_17944,N_18923);
nand U21239 (N_21239,N_19567,N_19144);
and U21240 (N_21240,N_17348,N_18684);
nor U21241 (N_21241,N_19614,N_16166);
nor U21242 (N_21242,N_15182,N_15267);
and U21243 (N_21243,N_16239,N_17247);
nor U21244 (N_21244,N_16729,N_18288);
nor U21245 (N_21245,N_17415,N_15779);
nand U21246 (N_21246,N_19040,N_15202);
nor U21247 (N_21247,N_15775,N_16954);
xor U21248 (N_21248,N_17656,N_17005);
xnor U21249 (N_21249,N_19747,N_18901);
nand U21250 (N_21250,N_15126,N_16500);
xor U21251 (N_21251,N_19730,N_16849);
or U21252 (N_21252,N_17888,N_18013);
xor U21253 (N_21253,N_17365,N_15838);
nor U21254 (N_21254,N_17699,N_17583);
or U21255 (N_21255,N_19178,N_18521);
nor U21256 (N_21256,N_18100,N_18392);
nand U21257 (N_21257,N_15953,N_15257);
nor U21258 (N_21258,N_16175,N_17508);
or U21259 (N_21259,N_18716,N_17853);
nor U21260 (N_21260,N_16689,N_17263);
xnor U21261 (N_21261,N_16649,N_16590);
nor U21262 (N_21262,N_18891,N_16347);
or U21263 (N_21263,N_16369,N_18158);
or U21264 (N_21264,N_16912,N_19699);
and U21265 (N_21265,N_16563,N_17700);
or U21266 (N_21266,N_19679,N_16492);
xnor U21267 (N_21267,N_18095,N_18560);
or U21268 (N_21268,N_16446,N_15290);
xor U21269 (N_21269,N_15781,N_15710);
nand U21270 (N_21270,N_19029,N_19442);
nor U21271 (N_21271,N_17413,N_19902);
and U21272 (N_21272,N_18436,N_18464);
and U21273 (N_21273,N_17806,N_19186);
xnor U21274 (N_21274,N_17576,N_15467);
and U21275 (N_21275,N_16220,N_15626);
and U21276 (N_21276,N_15443,N_16877);
and U21277 (N_21277,N_18126,N_18165);
and U21278 (N_21278,N_18042,N_18550);
xor U21279 (N_21279,N_15404,N_19892);
nand U21280 (N_21280,N_16828,N_18251);
xnor U21281 (N_21281,N_16192,N_16212);
xnor U21282 (N_21282,N_16147,N_16113);
nor U21283 (N_21283,N_16667,N_15639);
or U21284 (N_21284,N_16800,N_19047);
nor U21285 (N_21285,N_17960,N_17192);
nand U21286 (N_21286,N_16368,N_18065);
or U21287 (N_21287,N_17225,N_16096);
nor U21288 (N_21288,N_18823,N_18211);
and U21289 (N_21289,N_19563,N_17129);
nand U21290 (N_21290,N_19982,N_16435);
nand U21291 (N_21291,N_18974,N_19640);
nor U21292 (N_21292,N_18461,N_19077);
nand U21293 (N_21293,N_18513,N_16981);
or U21294 (N_21294,N_16332,N_15818);
and U21295 (N_21295,N_15422,N_17492);
and U21296 (N_21296,N_15793,N_19420);
xnor U21297 (N_21297,N_15035,N_19970);
xor U21298 (N_21298,N_17502,N_17169);
nand U21299 (N_21299,N_15750,N_17675);
and U21300 (N_21300,N_16543,N_18279);
and U21301 (N_21301,N_18159,N_16088);
and U21302 (N_21302,N_16526,N_19387);
xnor U21303 (N_21303,N_19707,N_18429);
or U21304 (N_21304,N_17677,N_19946);
nand U21305 (N_21305,N_16066,N_16743);
or U21306 (N_21306,N_16742,N_15583);
nor U21307 (N_21307,N_18019,N_19001);
nand U21308 (N_21308,N_17687,N_15994);
and U21309 (N_21309,N_19207,N_15501);
or U21310 (N_21310,N_18061,N_16304);
or U21311 (N_21311,N_15935,N_18318);
or U21312 (N_21312,N_19820,N_17047);
nor U21313 (N_21313,N_19069,N_16998);
xnor U21314 (N_21314,N_16262,N_17506);
xnor U21315 (N_21315,N_19346,N_19172);
nand U21316 (N_21316,N_19279,N_17270);
or U21317 (N_21317,N_17301,N_15827);
or U21318 (N_21318,N_15351,N_15332);
xnor U21319 (N_21319,N_18481,N_18561);
or U21320 (N_21320,N_16773,N_16258);
and U21321 (N_21321,N_15336,N_19997);
or U21322 (N_21322,N_15372,N_16984);
nor U21323 (N_21323,N_17814,N_19893);
or U21324 (N_21324,N_16992,N_16652);
nor U21325 (N_21325,N_16573,N_15396);
xnor U21326 (N_21326,N_18675,N_17844);
or U21327 (N_21327,N_19524,N_15490);
and U21328 (N_21328,N_18902,N_16680);
nor U21329 (N_21329,N_15601,N_17078);
nor U21330 (N_21330,N_16916,N_19104);
nand U21331 (N_21331,N_17965,N_15617);
and U21332 (N_21332,N_19800,N_16470);
or U21333 (N_21333,N_17491,N_19162);
and U21334 (N_21334,N_18498,N_17422);
nand U21335 (N_21335,N_19554,N_19601);
xor U21336 (N_21336,N_15140,N_15984);
nor U21337 (N_21337,N_19305,N_18813);
and U21338 (N_21338,N_15675,N_19698);
nand U21339 (N_21339,N_16668,N_16073);
and U21340 (N_21340,N_18422,N_16308);
xnor U21341 (N_21341,N_17610,N_17087);
or U21342 (N_21342,N_19490,N_15656);
or U21343 (N_21343,N_17320,N_15678);
nand U21344 (N_21344,N_15965,N_15707);
nand U21345 (N_21345,N_16684,N_15963);
and U21346 (N_21346,N_19082,N_16031);
and U21347 (N_21347,N_19746,N_19248);
or U21348 (N_21348,N_19164,N_15053);
or U21349 (N_21349,N_17294,N_18918);
nor U21350 (N_21350,N_18246,N_18770);
xor U21351 (N_21351,N_19657,N_15307);
xnor U21352 (N_21352,N_18671,N_15804);
or U21353 (N_21353,N_17121,N_19243);
and U21354 (N_21354,N_15297,N_17902);
nor U21355 (N_21355,N_15816,N_19753);
xor U21356 (N_21356,N_17705,N_15012);
or U21357 (N_21357,N_19079,N_15968);
or U21358 (N_21358,N_15589,N_16297);
xnor U21359 (N_21359,N_17686,N_16254);
nor U21360 (N_21360,N_15783,N_17871);
xnor U21361 (N_21361,N_17324,N_17929);
or U21362 (N_21362,N_15280,N_18840);
xor U21363 (N_21363,N_17246,N_16422);
xor U21364 (N_21364,N_18051,N_17391);
nor U21365 (N_21365,N_17006,N_18292);
and U21366 (N_21366,N_16595,N_19192);
and U21367 (N_21367,N_17928,N_17962);
nor U21368 (N_21368,N_17184,N_17487);
nor U21369 (N_21369,N_18172,N_18103);
and U21370 (N_21370,N_15495,N_18174);
or U21371 (N_21371,N_18055,N_19478);
and U21372 (N_21372,N_15145,N_18581);
or U21373 (N_21373,N_17600,N_19773);
or U21374 (N_21374,N_17451,N_17896);
or U21375 (N_21375,N_18582,N_19651);
or U21376 (N_21376,N_16259,N_16040);
and U21377 (N_21377,N_17167,N_19745);
or U21378 (N_21378,N_18094,N_19634);
xor U21379 (N_21379,N_16059,N_15394);
xor U21380 (N_21380,N_19617,N_19035);
and U21381 (N_21381,N_15399,N_15505);
nor U21382 (N_21382,N_17632,N_15607);
nand U21383 (N_21383,N_15333,N_19660);
nor U21384 (N_21384,N_18800,N_16478);
xnor U21385 (N_21385,N_19576,N_16364);
xnor U21386 (N_21386,N_19832,N_16357);
nand U21387 (N_21387,N_18351,N_16249);
and U21388 (N_21388,N_15672,N_15663);
and U21389 (N_21389,N_16139,N_16893);
nor U21390 (N_21390,N_16496,N_16931);
nor U21391 (N_21391,N_16075,N_19973);
or U21392 (N_21392,N_16822,N_18096);
or U21393 (N_21393,N_17612,N_16359);
and U21394 (N_21394,N_17177,N_17341);
xnor U21395 (N_21395,N_18697,N_16973);
xnor U21396 (N_21396,N_19130,N_19974);
or U21397 (N_21397,N_19412,N_16493);
and U21398 (N_21398,N_18803,N_17821);
and U21399 (N_21399,N_19401,N_16521);
nor U21400 (N_21400,N_19444,N_15087);
or U21401 (N_21401,N_16004,N_16427);
or U21402 (N_21402,N_19884,N_18908);
or U21403 (N_21403,N_19777,N_19151);
or U21404 (N_21404,N_17086,N_18470);
nand U21405 (N_21405,N_15616,N_15361);
nor U21406 (N_21406,N_15433,N_16568);
or U21407 (N_21407,N_15214,N_16015);
and U21408 (N_21408,N_16182,N_19954);
xnor U21409 (N_21409,N_16206,N_17111);
or U21410 (N_21410,N_16023,N_15790);
nor U21411 (N_21411,N_18808,N_17462);
xor U21412 (N_21412,N_18935,N_15731);
nand U21413 (N_21413,N_17193,N_18695);
xnor U21414 (N_21414,N_15228,N_18052);
or U21415 (N_21415,N_16834,N_16783);
or U21416 (N_21416,N_19875,N_19051);
and U21417 (N_21417,N_19050,N_16138);
nor U21418 (N_21418,N_17855,N_18572);
nor U21419 (N_21419,N_19836,N_17553);
nand U21420 (N_21420,N_19726,N_16307);
nor U21421 (N_21421,N_15809,N_17991);
nand U21422 (N_21422,N_19659,N_17790);
nor U21423 (N_21423,N_15255,N_18450);
nor U21424 (N_21424,N_19124,N_19452);
or U21425 (N_21425,N_15954,N_19239);
xor U21426 (N_21426,N_19008,N_18640);
or U21427 (N_21427,N_18142,N_18703);
xor U21428 (N_21428,N_16956,N_18484);
xnor U21429 (N_21429,N_18596,N_16305);
or U21430 (N_21430,N_17466,N_17014);
xor U21431 (N_21431,N_19579,N_15666);
or U21432 (N_21432,N_18683,N_16009);
nand U21433 (N_21433,N_19423,N_18398);
and U21434 (N_21434,N_15312,N_18873);
xnor U21435 (N_21435,N_17477,N_18900);
nand U21436 (N_21436,N_16763,N_19890);
and U21437 (N_21437,N_18586,N_19663);
nor U21438 (N_21438,N_17858,N_15735);
xor U21439 (N_21439,N_17404,N_15681);
or U21440 (N_21440,N_15121,N_16752);
and U21441 (N_21441,N_16158,N_16503);
xor U21442 (N_21442,N_17230,N_17304);
or U21443 (N_21443,N_18879,N_15561);
or U21444 (N_21444,N_19214,N_18452);
and U21445 (N_21445,N_18413,N_17641);
xor U21446 (N_21446,N_15213,N_17003);
nor U21447 (N_21447,N_16736,N_19678);
or U21448 (N_21448,N_17372,N_17402);
and U21449 (N_21449,N_17596,N_17839);
and U21450 (N_21450,N_18266,N_16996);
or U21451 (N_21451,N_17174,N_19821);
and U21452 (N_21452,N_15060,N_18387);
xor U21453 (N_21453,N_16039,N_16339);
and U21454 (N_21454,N_16816,N_16278);
xor U21455 (N_21455,N_19995,N_18423);
nor U21456 (N_21456,N_15154,N_16038);
nor U21457 (N_21457,N_15826,N_17869);
nor U21458 (N_21458,N_17394,N_18993);
and U21459 (N_21459,N_18571,N_16454);
nor U21460 (N_21460,N_19888,N_16474);
nand U21461 (N_21461,N_15534,N_18310);
xor U21462 (N_21462,N_19026,N_17992);
and U21463 (N_21463,N_19295,N_17756);
nand U21464 (N_21464,N_15367,N_18455);
nor U21465 (N_21465,N_16577,N_18007);
and U21466 (N_21466,N_19010,N_15194);
xor U21467 (N_21467,N_16080,N_15895);
and U21468 (N_21468,N_16513,N_15882);
nor U21469 (N_21469,N_16683,N_15395);
and U21470 (N_21470,N_16228,N_15623);
xnor U21471 (N_21471,N_19036,N_18737);
xor U21472 (N_21472,N_15774,N_17377);
nand U21473 (N_21473,N_19582,N_15657);
nand U21474 (N_21474,N_18689,N_16559);
nor U21475 (N_21475,N_15349,N_17310);
nand U21476 (N_21476,N_19598,N_16119);
nand U21477 (N_21477,N_16572,N_17489);
xnor U21478 (N_21478,N_19696,N_17183);
and U21479 (N_21479,N_17877,N_19398);
nand U21480 (N_21480,N_16589,N_17807);
nand U21481 (N_21481,N_19771,N_18913);
nand U21482 (N_21482,N_19858,N_17946);
or U21483 (N_21483,N_17081,N_19274);
or U21484 (N_21484,N_18871,N_19368);
nand U21485 (N_21485,N_16848,N_18558);
nand U21486 (N_21486,N_15613,N_18204);
or U21487 (N_21487,N_15852,N_19254);
or U21488 (N_21488,N_15104,N_16062);
and U21489 (N_21489,N_18851,N_15891);
and U21490 (N_21490,N_16856,N_15281);
or U21491 (N_21491,N_15286,N_19596);
or U21492 (N_21492,N_18909,N_16312);
xor U21493 (N_21493,N_15429,N_16986);
or U21494 (N_21494,N_17966,N_15961);
and U21495 (N_21495,N_15684,N_16202);
or U21496 (N_21496,N_15206,N_15250);
nor U21497 (N_21497,N_15949,N_17286);
xor U21498 (N_21498,N_16623,N_18752);
and U21499 (N_21499,N_19394,N_18022);
or U21500 (N_21500,N_16911,N_17235);
xnor U21501 (N_21501,N_18627,N_15207);
and U21502 (N_21502,N_17842,N_18925);
and U21503 (N_21503,N_17948,N_15085);
nand U21504 (N_21504,N_18301,N_19147);
nor U21505 (N_21505,N_15832,N_18054);
nand U21506 (N_21506,N_19296,N_19801);
and U21507 (N_21507,N_15845,N_15470);
or U21508 (N_21508,N_18623,N_17956);
nand U21509 (N_21509,N_19965,N_18763);
or U21510 (N_21510,N_18641,N_15147);
or U21511 (N_21511,N_19133,N_16090);
and U21512 (N_21512,N_17349,N_18959);
nand U21513 (N_21513,N_17906,N_19226);
or U21514 (N_21514,N_15573,N_15358);
xor U21515 (N_21515,N_19150,N_16317);
nor U21516 (N_21516,N_18620,N_18812);
and U21517 (N_21517,N_18062,N_15659);
xnor U21518 (N_21518,N_16639,N_18426);
nand U21519 (N_21519,N_18161,N_19649);
nor U21520 (N_21520,N_18858,N_18503);
or U21521 (N_21521,N_19328,N_18109);
nand U21522 (N_21522,N_15459,N_15148);
xor U21523 (N_21523,N_17153,N_19175);
or U21524 (N_21524,N_15298,N_17307);
xor U21525 (N_21525,N_19436,N_16479);
nor U21526 (N_21526,N_18793,N_15223);
xor U21527 (N_21527,N_16395,N_16489);
nor U21528 (N_21528,N_18190,N_19607);
and U21529 (N_21529,N_18356,N_15546);
or U21530 (N_21530,N_19729,N_18389);
nand U21531 (N_21531,N_18372,N_16191);
and U21532 (N_21532,N_18715,N_16375);
nor U21533 (N_21533,N_19075,N_15319);
nor U21534 (N_21534,N_17098,N_16632);
and U21535 (N_21535,N_17857,N_17880);
and U21536 (N_21536,N_17625,N_18346);
nor U21537 (N_21537,N_16815,N_19874);
nor U21538 (N_21538,N_18036,N_16517);
xnor U21539 (N_21539,N_19145,N_19074);
or U21540 (N_21540,N_18548,N_16548);
nor U21541 (N_21541,N_16505,N_16604);
nor U21542 (N_21542,N_17834,N_19491);
or U21543 (N_21543,N_17120,N_17824);
or U21544 (N_21544,N_17934,N_18704);
and U21545 (N_21545,N_15414,N_17535);
nor U21546 (N_21546,N_15929,N_19791);
xor U21547 (N_21547,N_18027,N_17644);
or U21548 (N_21548,N_19781,N_16971);
nand U21549 (N_21549,N_17591,N_17728);
xnor U21550 (N_21550,N_18662,N_19265);
and U21551 (N_21551,N_17362,N_15176);
nor U21552 (N_21552,N_16887,N_19735);
or U21553 (N_21553,N_17239,N_16928);
nor U21554 (N_21554,N_17735,N_19244);
xnor U21555 (N_21555,N_19396,N_19683);
nand U21556 (N_21556,N_17685,N_18181);
and U21557 (N_21557,N_17725,N_15835);
or U21558 (N_21558,N_17861,N_16272);
or U21559 (N_21559,N_17933,N_19372);
or U21560 (N_21560,N_15002,N_17766);
nor U21561 (N_21561,N_15238,N_17460);
nand U21562 (N_21562,N_19756,N_17949);
or U21563 (N_21563,N_16007,N_16775);
or U21564 (N_21564,N_18512,N_16118);
nor U21565 (N_21565,N_16747,N_17159);
or U21566 (N_21566,N_18039,N_16720);
or U21567 (N_21567,N_19292,N_16150);
or U21568 (N_21568,N_18817,N_16824);
nand U21569 (N_21569,N_18828,N_16507);
nand U21570 (N_21570,N_18050,N_15641);
nand U21571 (N_21571,N_18059,N_16253);
or U21572 (N_21572,N_17316,N_15137);
and U21573 (N_21573,N_17778,N_17668);
nand U21574 (N_21574,N_17505,N_18212);
xor U21575 (N_21575,N_17547,N_18599);
or U21576 (N_21576,N_15383,N_17220);
and U21577 (N_21577,N_16018,N_17455);
nand U21578 (N_21578,N_16012,N_15788);
or U21579 (N_21579,N_15631,N_15604);
xor U21580 (N_21580,N_19788,N_15171);
nand U21581 (N_21581,N_16170,N_17367);
xnor U21582 (N_21582,N_19916,N_15011);
nand U21583 (N_21583,N_16874,N_16695);
and U21584 (N_21584,N_19005,N_15409);
and U21585 (N_21585,N_18421,N_15452);
or U21586 (N_21586,N_19031,N_19975);
nand U21587 (N_21587,N_16764,N_17651);
or U21588 (N_21588,N_15906,N_15785);
nand U21589 (N_21589,N_17615,N_16910);
nor U21590 (N_21590,N_17016,N_17376);
xnor U21591 (N_21591,N_17802,N_17331);
and U21592 (N_21592,N_19695,N_19483);
nor U21593 (N_21593,N_17067,N_19492);
nor U21594 (N_21594,N_16216,N_18559);
nand U21595 (N_21595,N_17401,N_19076);
nand U21596 (N_21596,N_17595,N_19742);
xnor U21597 (N_21597,N_15466,N_17891);
nor U21598 (N_21598,N_16156,N_18597);
nand U21599 (N_21599,N_17136,N_19990);
nand U21600 (N_21600,N_18797,N_19949);
xor U21601 (N_21601,N_16846,N_17308);
nand U21602 (N_21602,N_18187,N_15599);
and U21603 (N_21603,N_16013,N_17915);
nand U21604 (N_21604,N_15066,N_16382);
or U21605 (N_21605,N_15059,N_15784);
and U21606 (N_21606,N_18760,N_16929);
and U21607 (N_21607,N_17450,N_15794);
or U21608 (N_21608,N_19203,N_15587);
xnor U21609 (N_21609,N_19057,N_19967);
xor U21610 (N_21610,N_17323,N_19083);
xnor U21611 (N_21611,N_19912,N_19400);
or U21612 (N_21612,N_19230,N_19962);
xnor U21613 (N_21613,N_18252,N_16302);
or U21614 (N_21614,N_15511,N_18216);
xnor U21615 (N_21615,N_15426,N_18091);
nand U21616 (N_21616,N_17389,N_17829);
xor U21617 (N_21617,N_17297,N_17229);
and U21618 (N_21618,N_17250,N_16264);
nor U21619 (N_21619,N_17306,N_17485);
or U21620 (N_21620,N_18213,N_17023);
or U21621 (N_21621,N_18127,N_17296);
or U21622 (N_21622,N_15570,N_19194);
nand U21623 (N_21623,N_15247,N_19132);
nand U21624 (N_21624,N_19140,N_18635);
or U21625 (N_21625,N_18290,N_17046);
xor U21626 (N_21626,N_17425,N_16858);
xnor U21627 (N_21627,N_19182,N_15876);
nand U21628 (N_21628,N_16918,N_15288);
nor U21629 (N_21629,N_16186,N_18004);
xor U21630 (N_21630,N_16173,N_16197);
or U21631 (N_21631,N_15916,N_18031);
or U21632 (N_21632,N_17525,N_18046);
nand U21633 (N_21633,N_17007,N_15560);
nand U21634 (N_21634,N_17604,N_18235);
xor U21635 (N_21635,N_19797,N_19504);
and U21636 (N_21636,N_15274,N_15402);
nor U21637 (N_21637,N_16980,N_18412);
xnor U21638 (N_21638,N_19259,N_15130);
nand U21639 (N_21639,N_19714,N_17360);
or U21640 (N_21640,N_17127,N_15597);
or U21641 (N_21641,N_15862,N_18345);
nor U21642 (N_21642,N_16421,N_15559);
nand U21643 (N_21643,N_15567,N_19709);
or U21644 (N_21644,N_17791,N_16293);
xnor U21645 (N_21645,N_16945,N_15640);
nand U21646 (N_21646,N_19842,N_19515);
nand U21647 (N_21647,N_15802,N_15192);
or U21648 (N_21648,N_17464,N_19439);
nor U21649 (N_21649,N_15018,N_15187);
or U21650 (N_21650,N_16705,N_16376);
and U21651 (N_21651,N_18053,N_18546);
and U21652 (N_21652,N_16750,N_18726);
nor U21653 (N_21653,N_16106,N_17390);
nor U21654 (N_21654,N_16242,N_19189);
nand U21655 (N_21655,N_19392,N_18278);
xnor U21656 (N_21656,N_18511,N_17803);
nand U21657 (N_21657,N_18999,N_15227);
nand U21658 (N_21658,N_18646,N_15460);
nand U21659 (N_21659,N_17762,N_19038);
xor U21660 (N_21660,N_15926,N_19581);
or U21661 (N_21661,N_16078,N_19662);
nand U21662 (N_21662,N_19823,N_18219);
nand U21663 (N_21663,N_16148,N_16927);
and U21664 (N_21664,N_18595,N_16528);
or U21665 (N_21665,N_15771,N_17321);
and U21666 (N_21666,N_15481,N_16995);
nand U21667 (N_21667,N_16781,N_17859);
nor U21668 (N_21668,N_17703,N_18300);
and U21669 (N_21669,N_18783,N_19363);
nor U21670 (N_21670,N_18788,N_17071);
and U21671 (N_21671,N_16890,N_18196);
or U21672 (N_21672,N_16045,N_17768);
nor U21673 (N_21673,N_19185,N_17701);
xor U21674 (N_21674,N_19812,N_19165);
nand U21675 (N_21675,N_17036,N_17819);
and U21676 (N_21676,N_15301,N_18806);
and U21677 (N_21677,N_17874,N_19963);
and U21678 (N_21678,N_18723,N_18018);
nand U21679 (N_21679,N_18942,N_15942);
or U21680 (N_21680,N_16441,N_15605);
nor U21681 (N_21681,N_18033,N_18099);
or U21682 (N_21682,N_18776,N_17090);
nor U21683 (N_21683,N_17020,N_19920);
and U21684 (N_21684,N_19684,N_19633);
nand U21685 (N_21685,N_17927,N_16495);
and U21686 (N_21686,N_16949,N_19419);
xnor U21687 (N_21687,N_17168,N_16855);
nand U21688 (N_21688,N_16349,N_18256);
or U21689 (N_21689,N_19761,N_15620);
xnor U21690 (N_21690,N_19448,N_17957);
and U21691 (N_21691,N_15997,N_19286);
or U21692 (N_21692,N_18651,N_15629);
nand U21693 (N_21693,N_19060,N_15842);
nand U21694 (N_21694,N_17984,N_16905);
nor U21695 (N_21695,N_19558,N_17009);
nor U21696 (N_21696,N_15088,N_17868);
and U21697 (N_21697,N_19058,N_15191);
and U21698 (N_21698,N_17197,N_19445);
nand U21699 (N_21699,N_16335,N_18373);
xor U21700 (N_21700,N_17925,N_16990);
or U21701 (N_21701,N_16473,N_15603);
or U21702 (N_21702,N_17338,N_15478);
nor U21703 (N_21703,N_18679,N_18691);
nand U21704 (N_21704,N_17512,N_16135);
nor U21705 (N_21705,N_17226,N_18841);
and U21706 (N_21706,N_16195,N_19700);
nor U21707 (N_21707,N_19267,N_15927);
nand U21708 (N_21708,N_17528,N_17550);
nand U21709 (N_21709,N_17789,N_15934);
and U21710 (N_21710,N_18861,N_17769);
xnor U21711 (N_21711,N_16463,N_19616);
or U21712 (N_21712,N_16702,N_16240);
and U21713 (N_21713,N_17265,N_16306);
and U21714 (N_21714,N_16718,N_15461);
nor U21715 (N_21715,N_18870,N_18040);
or U21716 (N_21716,N_16786,N_17545);
nand U21717 (N_21717,N_19583,N_16211);
nand U21718 (N_21718,N_16839,N_15236);
xnor U21719 (N_21719,N_18291,N_19636);
nor U21720 (N_21720,N_17066,N_19976);
and U21721 (N_21721,N_18732,N_18240);
and U21722 (N_21722,N_16342,N_19285);
nand U21723 (N_21723,N_16616,N_19883);
nor U21724 (N_21724,N_17696,N_17224);
nand U21725 (N_21725,N_17370,N_19600);
xor U21726 (N_21726,N_15575,N_17074);
or U21727 (N_21727,N_15177,N_18044);
or U21728 (N_21728,N_16494,N_18859);
or U21729 (N_21729,N_18144,N_19925);
nand U21730 (N_21730,N_16757,N_18341);
or U21731 (N_21731,N_18000,N_18071);
nand U21732 (N_21732,N_19356,N_18483);
xnor U21733 (N_21733,N_15915,N_18267);
nor U21734 (N_21734,N_19160,N_18323);
and U21735 (N_21735,N_15960,N_15254);
xnor U21736 (N_21736,N_15324,N_16331);
and U21737 (N_21737,N_16414,N_17253);
or U21738 (N_21738,N_19156,N_19932);
nand U21739 (N_21739,N_16881,N_17186);
nand U21740 (N_21740,N_16642,N_15107);
xor U21741 (N_21741,N_19094,N_15262);
and U21742 (N_21742,N_15995,N_16557);
or U21743 (N_21743,N_16670,N_16353);
or U21744 (N_21744,N_19702,N_15956);
and U21745 (N_21745,N_18072,N_16208);
xnor U21746 (N_21746,N_16383,N_17692);
nand U21747 (N_21747,N_18164,N_15313);
and U21748 (N_21748,N_15502,N_19461);
nand U21749 (N_21749,N_17648,N_16983);
nand U21750 (N_21750,N_17179,N_15204);
nand U21751 (N_21751,N_17269,N_18939);
or U21752 (N_21752,N_17817,N_16036);
xnor U21753 (N_21753,N_16804,N_16224);
or U21754 (N_21754,N_19460,N_17386);
xor U21755 (N_21755,N_17890,N_17564);
and U21756 (N_21756,N_17779,N_17524);
or U21757 (N_21757,N_17113,N_19993);
and U21758 (N_21758,N_17597,N_16370);
nand U21759 (N_21759,N_19466,N_17574);
nor U21760 (N_21760,N_15822,N_18353);
nor U21761 (N_21761,N_19225,N_18098);
xor U21762 (N_21762,N_18606,N_15878);
nor U21763 (N_21763,N_15863,N_15539);
nand U21764 (N_21764,N_17428,N_18214);
and U21765 (N_21765,N_16968,N_19938);
nor U21766 (N_21766,N_19585,N_15353);
xnor U21767 (N_21767,N_15726,N_19792);
or U21768 (N_21768,N_16967,N_17513);
and U21769 (N_21769,N_15757,N_17475);
xnor U21770 (N_21770,N_17144,N_15049);
and U21771 (N_21771,N_19602,N_16900);
nor U21772 (N_21772,N_16313,N_18554);
xnor U21773 (N_21773,N_16621,N_19811);
and U21774 (N_21774,N_18008,N_18539);
xor U21775 (N_21775,N_15889,N_15724);
and U21776 (N_21776,N_18284,N_17173);
and U21777 (N_21777,N_17867,N_18191);
and U21778 (N_21778,N_15103,N_15471);
or U21779 (N_21779,N_19177,N_17423);
xnor U21780 (N_21780,N_17175,N_17315);
xnor U21781 (N_21781,N_19855,N_16229);
or U21782 (N_21782,N_19233,N_15026);
or U21783 (N_21783,N_15690,N_16860);
and U21784 (N_21784,N_15158,N_19519);
nand U21785 (N_21785,N_16527,N_16011);
nor U21786 (N_21786,N_17646,N_17027);
xor U21787 (N_21787,N_15434,N_18030);
and U21788 (N_21788,N_18832,N_19309);
or U21789 (N_21789,N_17072,N_19933);
and U21790 (N_21790,N_15293,N_16699);
and U21791 (N_21791,N_15520,N_15682);
nand U21792 (N_21792,N_19790,N_16116);
nand U21793 (N_21793,N_16022,N_19417);
nand U21794 (N_21794,N_15453,N_15271);
nand U21795 (N_21795,N_18916,N_15447);
nor U21796 (N_21796,N_18950,N_17914);
xor U21797 (N_21797,N_17101,N_19882);
nand U21798 (N_21798,N_18827,N_16768);
nand U21799 (N_21799,N_17264,N_19715);
or U21800 (N_21800,N_19033,N_17599);
xor U21801 (N_21801,N_18093,N_17211);
nand U21802 (N_21802,N_15445,N_15095);
xnor U21803 (N_21803,N_16315,N_17303);
or U21804 (N_21804,N_19674,N_15973);
or U21805 (N_21805,N_18207,N_19620);
and U21806 (N_21806,N_18725,N_18720);
and U21807 (N_21807,N_15189,N_19628);
or U21808 (N_21808,N_17835,N_19055);
nor U21809 (N_21809,N_15376,N_18929);
or U21810 (N_21810,N_19167,N_17234);
or U21811 (N_21811,N_18230,N_15455);
xor U21812 (N_21812,N_16506,N_17268);
xnor U21813 (N_21813,N_18530,N_17204);
and U21814 (N_21814,N_18006,N_17518);
xnor U21815 (N_21815,N_19300,N_18867);
nand U21816 (N_21816,N_15705,N_18696);
xnor U21817 (N_21817,N_16991,N_19841);
or U21818 (N_21818,N_17501,N_18294);
nand U21819 (N_21819,N_16704,N_18308);
nor U21820 (N_21820,N_16615,N_15920);
or U21821 (N_21821,N_18079,N_18233);
nand U21822 (N_21822,N_15229,N_19988);
nor U21823 (N_21823,N_16002,N_15479);
or U21824 (N_21824,N_15537,N_17207);
xnor U21825 (N_21825,N_18456,N_19481);
or U21826 (N_21826,N_18905,N_19769);
nor U21827 (N_21827,N_16055,N_15305);
nand U21828 (N_21828,N_18193,N_17970);
xor U21829 (N_21829,N_17057,N_18888);
and U21830 (N_21830,N_15258,N_17156);
and U21831 (N_21831,N_18856,N_16782);
nand U21832 (N_21832,N_15454,N_15582);
nor U21833 (N_21833,N_17776,N_19117);
or U21834 (N_21834,N_15877,N_17195);
and U21835 (N_21835,N_15945,N_16235);
nand U21836 (N_21836,N_17445,N_17800);
xor U21837 (N_21837,N_17444,N_15660);
nand U21838 (N_21838,N_18877,N_15670);
xor U21839 (N_21839,N_18083,N_16502);
nor U21840 (N_21840,N_16565,N_17657);
and U21841 (N_21841,N_15717,N_18132);
or U21842 (N_21842,N_15146,N_18309);
nand U21843 (N_21843,N_15855,N_15881);
and U21844 (N_21844,N_19347,N_16625);
nor U21845 (N_21845,N_15165,N_16762);
and U21846 (N_21846,N_15800,N_17419);
and U21847 (N_21847,N_16482,N_18552);
and U21848 (N_21848,N_16194,N_17690);
nor U21849 (N_21849,N_19391,N_18750);
nor U21850 (N_21850,N_16076,N_19059);
xor U21851 (N_21851,N_15571,N_16163);
nor U21852 (N_21852,N_15067,N_16605);
and U21853 (N_21853,N_19158,N_15814);
nand U21854 (N_21854,N_15836,N_19750);
nor U21855 (N_21855,N_19863,N_16586);
and U21856 (N_21856,N_17760,N_18979);
nor U21857 (N_21857,N_16894,N_19757);
or U21858 (N_21858,N_19121,N_15515);
nand U21859 (N_21859,N_16326,N_18914);
nand U21860 (N_21860,N_18874,N_17210);
and U21861 (N_21861,N_16732,N_16917);
or U21862 (N_21862,N_17516,N_18973);
nand U21863 (N_21863,N_18088,N_16845);
or U21864 (N_21864,N_16599,N_15728);
nor U21865 (N_21865,N_16465,N_19752);
nor U21866 (N_21866,N_19021,N_17132);
nor U21867 (N_21867,N_17408,N_19584);
nor U21868 (N_21868,N_17088,N_18189);
or U21869 (N_21869,N_16047,N_19326);
xnor U21870 (N_21870,N_18672,N_17030);
xnor U21871 (N_21871,N_15776,N_19512);
nor U21872 (N_21872,N_17815,N_15513);
nand U21873 (N_21873,N_19424,N_17849);
nor U21874 (N_21874,N_18122,N_17567);
nand U21875 (N_21875,N_17335,N_17638);
or U21876 (N_21876,N_19835,N_19516);
nor U21877 (N_21877,N_15215,N_18680);
or U21878 (N_21878,N_16117,N_18379);
or U21879 (N_21879,N_18110,N_16498);
nor U21880 (N_21880,N_17919,N_19066);
xor U21881 (N_21881,N_16092,N_16295);
and U21882 (N_21882,N_17165,N_16960);
and U21883 (N_21883,N_18659,N_18125);
and U21884 (N_21884,N_16219,N_17616);
nand U21885 (N_21885,N_15347,N_16065);
nand U21886 (N_21886,N_17669,N_16832);
and U21887 (N_21887,N_18746,N_19824);
or U21888 (N_21888,N_19969,N_15530);
xnor U21889 (N_21889,N_18667,N_19146);
and U21890 (N_21890,N_18625,N_17396);
and U21891 (N_21891,N_16226,N_19154);
or U21892 (N_21892,N_16575,N_19003);
and U21893 (N_21893,N_16925,N_19964);
xnor U21894 (N_21894,N_16178,N_17180);
nor U21895 (N_21895,N_15065,N_19134);
nand U21896 (N_21896,N_16560,N_19266);
or U21897 (N_21897,N_15411,N_19465);
and U21898 (N_21898,N_15732,N_16663);
or U21899 (N_21899,N_19898,N_17639);
and U21900 (N_21900,N_15545,N_18924);
or U21901 (N_21901,N_15911,N_18958);
or U21902 (N_21902,N_15551,N_15195);
and U21903 (N_21903,N_17851,N_15665);
nor U21904 (N_21904,N_17931,N_18520);
or U21905 (N_21905,N_16870,N_19340);
or U21906 (N_21906,N_19808,N_18844);
nand U21907 (N_21907,N_17257,N_18363);
nand U21908 (N_21908,N_18565,N_17771);
and U21909 (N_21909,N_15533,N_18151);
or U21910 (N_21910,N_18782,N_15697);
xnor U21911 (N_21911,N_18087,N_19705);
or U21912 (N_21912,N_16939,N_18866);
and U21913 (N_21913,N_17727,N_17356);
and U21914 (N_21914,N_15860,N_15278);
and U21915 (N_21915,N_18104,N_17061);
xnor U21916 (N_21916,N_19484,N_16634);
nor U21917 (N_21917,N_16550,N_17196);
nor U21918 (N_21918,N_17398,N_16199);
and U21919 (N_21919,N_18227,N_15348);
xor U21920 (N_21920,N_15164,N_18790);
or U21921 (N_21921,N_18424,N_19272);
and U21922 (N_21922,N_16940,N_18236);
and U21923 (N_21923,N_16721,N_16134);
xnor U21924 (N_21924,N_17852,N_16525);
xor U21925 (N_21925,N_18629,N_19650);
xor U21926 (N_21926,N_19565,N_16491);
nor U21927 (N_21927,N_15397,N_17660);
nor U21928 (N_21928,N_15487,N_15651);
nor U21929 (N_21929,N_18229,N_18956);
or U21930 (N_21930,N_15864,N_15334);
xnor U21931 (N_21931,N_15713,N_17620);
or U21932 (N_21932,N_18781,N_16627);
nand U21933 (N_21933,N_19111,N_18884);
or U21934 (N_21934,N_16469,N_15673);
xor U21935 (N_21935,N_19815,N_15320);
xor U21936 (N_21936,N_17094,N_18633);
nand U21937 (N_21937,N_16391,N_15004);
nand U21938 (N_21938,N_19827,N_17138);
xor U21939 (N_21939,N_18391,N_17035);
nand U21940 (N_21940,N_18378,N_19810);
nand U21941 (N_21941,N_18609,N_15498);
or U21942 (N_21942,N_19333,N_18135);
or U21943 (N_21943,N_18167,N_17854);
or U21944 (N_21944,N_15992,N_18147);
or U21945 (N_21945,N_19302,N_18771);
or U21946 (N_21946,N_18502,N_17191);
nor U21947 (N_21947,N_18542,N_15547);
nor U21948 (N_21948,N_18275,N_15231);
nor U21949 (N_21949,N_19724,N_15196);
and U21950 (N_21950,N_15628,N_16294);
or U21951 (N_21951,N_16451,N_16230);
xor U21952 (N_21952,N_19181,N_18563);
nand U21953 (N_21953,N_18710,N_17240);
or U21954 (N_21954,N_15972,N_18209);
and U21955 (N_21955,N_16558,N_16162);
and U21956 (N_21956,N_17289,N_17680);
or U21957 (N_21957,N_19908,N_18056);
xnor U21958 (N_21958,N_18966,N_15957);
and U21959 (N_21959,N_19426,N_17784);
nand U21960 (N_21960,N_17070,N_16944);
nor U21961 (N_21961,N_16256,N_18713);
nand U21962 (N_21962,N_16672,N_17414);
nor U21963 (N_21963,N_16655,N_17155);
nand U21964 (N_21964,N_17503,N_19353);
or U21965 (N_21965,N_17319,N_15871);
nor U21966 (N_21966,N_15768,N_19112);
nand U21967 (N_21967,N_15039,N_16716);
or U21968 (N_21968,N_17695,N_19054);
and U21969 (N_21969,N_19680,N_15052);
nand U21970 (N_21970,N_15563,N_18768);
or U21971 (N_21971,N_18965,N_17125);
or U21972 (N_21972,N_19574,N_17170);
nand U21973 (N_21973,N_17069,N_17418);
nor U21974 (N_21974,N_15451,N_15070);
and U21975 (N_21975,N_17188,N_18076);
nor U21976 (N_21976,N_15198,N_17336);
or U21977 (N_21977,N_17519,N_16497);
xor U21978 (N_21978,N_15041,N_16979);
nand U21979 (N_21979,N_17378,N_16864);
nand U21980 (N_21980,N_17961,N_15144);
nand U21981 (N_21981,N_17110,N_17920);
nor U21982 (N_21982,N_15337,N_19725);
nor U21983 (N_21983,N_15743,N_19315);
nor U21984 (N_21984,N_16430,N_18045);
and U21985 (N_21985,N_17775,N_15738);
or U21986 (N_21986,N_15143,N_17904);
and U21987 (N_21987,N_17715,N_18757);
or U21988 (N_21988,N_15753,N_17161);
xnor U21989 (N_21989,N_19542,N_16176);
or U21990 (N_21990,N_18857,N_19661);
or U21991 (N_21991,N_19179,N_17261);
nor U21992 (N_21992,N_15410,N_16638);
xnor U21993 (N_21993,N_16869,N_19572);
nor U21994 (N_21994,N_16738,N_19826);
nor U21995 (N_21995,N_16189,N_19775);
xnor U21996 (N_21996,N_16429,N_17947);
nand U21997 (N_21997,N_17293,N_16948);
nor U21998 (N_21998,N_16982,N_17504);
and U21999 (N_21999,N_19904,N_18523);
nand U22000 (N_22000,N_15356,N_15400);
or U22001 (N_22001,N_18601,N_15869);
or U22002 (N_22002,N_18360,N_19455);
nor U22003 (N_22003,N_18735,N_17052);
nor U22004 (N_22004,N_15381,N_16609);
nor U22005 (N_22005,N_15263,N_16377);
nor U22006 (N_22006,N_18329,N_19529);
xnor U22007 (N_22007,N_17758,N_16261);
nor U22008 (N_22008,N_19603,N_19568);
and U22009 (N_22009,N_17474,N_18487);
nand U22010 (N_22010,N_16748,N_16920);
or U22011 (N_22011,N_16285,N_17939);
nand U22012 (N_22012,N_16060,N_15668);
nor U22013 (N_22013,N_17605,N_16275);
or U22014 (N_22014,N_19900,N_17160);
nor U22015 (N_22015,N_18676,N_18407);
or U22016 (N_22016,N_16159,N_18894);
xnor U22017 (N_22017,N_19928,N_19793);
and U22018 (N_22018,N_15016,N_18645);
nor U22019 (N_22019,N_19472,N_19024);
or U22020 (N_22020,N_15072,N_19136);
nand U22021 (N_22021,N_17496,N_18208);
nand U22022 (N_22022,N_19849,N_16396);
and U22023 (N_22023,N_16154,N_18847);
and U22024 (N_22024,N_17279,N_17786);
or U22025 (N_22025,N_15178,N_17527);
and U22026 (N_22026,N_19952,N_18831);
xnor U22027 (N_22027,N_16110,N_16965);
and U22028 (N_22028,N_16628,N_18427);
and U22029 (N_22029,N_15119,N_19143);
xnor U22030 (N_22030,N_15595,N_18632);
or U22031 (N_22031,N_17848,N_17262);
and U22032 (N_22032,N_15169,N_15644);
nor U22033 (N_22033,N_19537,N_18787);
and U22034 (N_22034,N_17116,N_19169);
and U22035 (N_22035,N_16193,N_19245);
xor U22036 (N_22036,N_15503,N_15113);
xnor U22037 (N_22037,N_17754,N_16737);
nor U22038 (N_22038,N_15823,N_19958);
nor U22039 (N_22039,N_16057,N_15983);
and U22040 (N_22040,N_18773,N_16685);
nand U22041 (N_22041,N_15824,N_19222);
and U22042 (N_22042,N_15638,N_16597);
nor U22043 (N_22043,N_15958,N_18293);
or U22044 (N_22044,N_16799,N_15549);
nor U22045 (N_22045,N_16209,N_16933);
nand U22046 (N_22046,N_19122,N_17045);
and U22047 (N_22047,N_17488,N_15910);
or U22048 (N_22048,N_17215,N_15115);
nor U22049 (N_22049,N_18201,N_15484);
or U22050 (N_22050,N_17437,N_15473);
and U22051 (N_22051,N_16168,N_15030);
nor U22052 (N_22052,N_16549,N_15477);
nand U22053 (N_22053,N_19523,N_19297);
xor U22054 (N_22054,N_15940,N_16310);
and U22055 (N_22055,N_18411,N_19342);
and U22056 (N_22056,N_15092,N_17280);
or U22057 (N_22057,N_15777,N_18178);
and U22058 (N_22058,N_16260,N_18462);
or U22059 (N_22059,N_19229,N_18200);
nor U22060 (N_22060,N_17399,N_19334);
and U22061 (N_22061,N_19510,N_17364);
or U22062 (N_22062,N_17998,N_15898);
nor U22063 (N_22063,N_16989,N_19559);
nand U22064 (N_22064,N_15318,N_15224);
and U22065 (N_22065,N_18380,N_18621);
and U22066 (N_22066,N_18205,N_19817);
or U22067 (N_22067,N_16442,N_16923);
xnor U22068 (N_22068,N_16111,N_15557);
or U22069 (N_22069,N_17152,N_19677);
xor U22070 (N_22070,N_15167,N_16700);
or U22071 (N_22071,N_17434,N_18428);
nor U22072 (N_22072,N_18357,N_19034);
or U22073 (N_22073,N_17892,N_17816);
xnor U22074 (N_22074,N_19240,N_18576);
nor U22075 (N_22075,N_17012,N_15253);
xnor U22076 (N_22076,N_18931,N_19872);
or U22077 (N_22077,N_15671,N_17271);
nand U22078 (N_22078,N_15676,N_16755);
xor U22079 (N_22079,N_19555,N_17080);
and U22080 (N_22080,N_17721,N_16444);
nand U22081 (N_22081,N_15220,N_16488);
and U22082 (N_22082,N_15232,N_17238);
nand U22083 (N_22083,N_16713,N_17470);
and U22084 (N_22084,N_16598,N_19268);
nor U22085 (N_22085,N_17106,N_18458);
or U22086 (N_22086,N_18432,N_18384);
and U22087 (N_22087,N_17137,N_19665);
nor U22088 (N_22088,N_17062,N_17075);
nand U22089 (N_22089,N_16406,N_15418);
nor U22090 (N_22090,N_15694,N_16947);
nand U22091 (N_22091,N_17708,N_15884);
nor U22092 (N_22092,N_18163,N_19180);
and U22093 (N_22093,N_18802,N_19667);
and U22094 (N_22094,N_17642,N_18533);
or U22095 (N_22095,N_17773,N_17456);
or U22096 (N_22096,N_16233,N_19482);
or U22097 (N_22097,N_16386,N_17241);
nor U22098 (N_22098,N_18603,N_15401);
or U22099 (N_22099,N_19632,N_19658);
and U22100 (N_22100,N_18226,N_15427);
or U22101 (N_22101,N_19374,N_17231);
and U22102 (N_22102,N_19011,N_19845);
xor U22103 (N_22103,N_15090,N_15507);
and U22104 (N_22104,N_15506,N_18555);
nand U22105 (N_22105,N_19838,N_16876);
xnor U22106 (N_22106,N_18983,N_19027);
and U22107 (N_22107,N_15610,N_17733);
or U22108 (N_22108,N_15001,N_15556);
nor U22109 (N_22109,N_17903,N_17274);
nand U22110 (N_22110,N_15155,N_19432);
nand U22111 (N_22111,N_19470,N_16276);
nand U22112 (N_22112,N_19499,N_15285);
or U22113 (N_22113,N_16155,N_15900);
and U22114 (N_22114,N_17601,N_18248);
and U22115 (N_22115,N_19716,N_15846);
xnor U22116 (N_22116,N_15190,N_17436);
and U22117 (N_22117,N_18268,N_16149);
or U22118 (N_22118,N_17557,N_19343);
nand U22119 (N_22119,N_17910,N_18202);
or U22120 (N_22120,N_15504,N_15055);
nor U22121 (N_22121,N_17227,N_16319);
xor U22122 (N_22122,N_19886,N_16533);
and U22123 (N_22123,N_18377,N_16068);
xnor U22124 (N_22124,N_17368,N_16978);
or U22125 (N_22125,N_15509,N_17340);
nand U22126 (N_22126,N_15157,N_16591);
or U22127 (N_22127,N_17205,N_19527);
or U22128 (N_22128,N_18577,N_15883);
nor U22129 (N_22129,N_18887,N_17430);
nand U22130 (N_22130,N_16452,N_17500);
and U22131 (N_22131,N_15701,N_15880);
or U22132 (N_22132,N_16941,N_18654);
nor U22133 (N_22133,N_16977,N_15007);
and U22134 (N_22134,N_15175,N_16903);
or U22135 (N_22135,N_17938,N_18418);
xor U22136 (N_22136,N_18920,N_17382);
nor U22137 (N_22137,N_18339,N_19015);
nor U22138 (N_22138,N_15234,N_19532);
nor U22139 (N_22139,N_15131,N_19337);
xnor U22140 (N_22140,N_18355,N_15858);
and U22141 (N_22141,N_19183,N_18649);
or U22142 (N_22142,N_17146,N_15810);
nor U22143 (N_22143,N_18685,N_16907);
and U22144 (N_22144,N_18077,N_17783);
or U22145 (N_22145,N_15680,N_18506);
or U22146 (N_22146,N_19655,N_15188);
nor U22147 (N_22147,N_15650,N_17493);
or U22148 (N_22148,N_15770,N_16279);
nand U22149 (N_22149,N_15025,N_17285);
xnor U22150 (N_22150,N_15606,N_18593);
nor U22151 (N_22151,N_18133,N_18467);
xor U22152 (N_22152,N_15586,N_15128);
or U22153 (N_22153,N_19187,N_15058);
or U22154 (N_22154,N_16385,N_18937);
or U22155 (N_22155,N_18573,N_19536);
xnor U22156 (N_22156,N_16112,N_15437);
nor U22157 (N_22157,N_17826,N_19252);
nor U22158 (N_22158,N_19779,N_18882);
and U22159 (N_22159,N_18602,N_17050);
xnor U22160 (N_22160,N_18492,N_15943);
nand U22161 (N_22161,N_17440,N_15197);
and U22162 (N_22162,N_17216,N_16044);
nor U22163 (N_22163,N_18744,N_15850);
nand U22164 (N_22164,N_17752,N_18471);
xnor U22165 (N_22165,N_15975,N_19348);
or U22166 (N_22166,N_16027,N_15815);
nand U22167 (N_22167,N_15592,N_15762);
nor U22168 (N_22168,N_19809,N_17212);
and U22169 (N_22169,N_19776,N_18798);
nor U22170 (N_22170,N_19383,N_16472);
or U22171 (N_22171,N_16600,N_19463);
and U22172 (N_22172,N_19339,N_15980);
xor U22173 (N_22173,N_18195,N_18066);
nor U22174 (N_22174,N_15521,N_19548);
nand U22175 (N_22175,N_19237,N_19042);
xnor U22176 (N_22176,N_19344,N_15754);
or U22177 (N_22177,N_16886,N_15352);
or U22178 (N_22178,N_15161,N_15047);
nand U22179 (N_22179,N_18239,N_19767);
nand U22180 (N_22180,N_15933,N_15892);
and U22181 (N_22181,N_19475,N_18299);
xor U22182 (N_22182,N_18400,N_15872);
nand U22183 (N_22183,N_15733,N_18977);
nor U22184 (N_22184,N_17714,N_18951);
nand U22185 (N_22185,N_16850,N_16745);
nor U22186 (N_22186,N_17314,N_19895);
or U22187 (N_22187,N_16407,N_15077);
nand U22188 (N_22188,N_17443,N_16085);
or U22189 (N_22189,N_15896,N_15311);
xnor U22190 (N_22190,N_16137,N_18583);
nor U22191 (N_22191,N_15245,N_16388);
and U22192 (N_22192,N_15082,N_15941);
nand U22193 (N_22193,N_18123,N_19739);
and U22194 (N_22194,N_17406,N_17544);
and U22195 (N_22195,N_15988,N_18981);
and U22196 (N_22196,N_15468,N_15661);
and U22197 (N_22197,N_18774,N_19522);
and U22198 (N_22198,N_16241,N_17585);
xor U22199 (N_22199,N_16999,N_15392);
nand U22200 (N_22200,N_19701,N_17662);
nor U22201 (N_22201,N_19764,N_15282);
or U22202 (N_22202,N_16711,N_15287);
nor U22203 (N_22203,N_16653,N_18319);
xnor U22204 (N_22204,N_19421,N_17856);
and U22205 (N_22205,N_15765,N_16445);
nor U22206 (N_22206,N_18535,N_17678);
xor U22207 (N_22207,N_15205,N_15186);
xor U22208 (N_22208,N_18730,N_19986);
nor U22209 (N_22209,N_19284,N_15806);
and U22210 (N_22210,N_19126,N_19625);
or U22211 (N_22211,N_17232,N_16378);
or U22212 (N_22212,N_18807,N_19281);
or U22213 (N_22213,N_19071,N_15221);
nor U22214 (N_22214,N_16184,N_17135);
nor U22215 (N_22215,N_17002,N_18352);
nand U22216 (N_22216,N_16708,N_19850);
and U22217 (N_22217,N_17374,N_18270);
or U22218 (N_22218,N_15403,N_18348);
nand U22219 (N_22219,N_19064,N_17627);
xor U22220 (N_22220,N_17392,N_16677);
nor U22221 (N_22221,N_18326,N_19273);
nor U22222 (N_22222,N_18669,N_19153);
nand U22223 (N_22223,N_18496,N_15022);
and U22224 (N_22224,N_17384,N_17633);
nand U22225 (N_22225,N_16198,N_17043);
nor U22226 (N_22226,N_17055,N_15269);
xor U22227 (N_22227,N_18221,N_19535);
xnor U22228 (N_22228,N_16969,N_17538);
or U22229 (N_22229,N_16564,N_17147);
nand U22230 (N_22230,N_18020,N_16499);
or U22231 (N_22231,N_16896,N_19271);
nor U22232 (N_22232,N_18010,N_18764);
nand U22233 (N_22233,N_18643,N_16611);
or U22234 (N_22234,N_15516,N_19561);
and U22235 (N_22235,N_16366,N_17731);
or U22236 (N_22236,N_15553,N_17060);
nand U22237 (N_22237,N_16371,N_19476);
and U22238 (N_22238,N_17439,N_19915);
xnor U22239 (N_22239,N_15662,N_17131);
nor U22240 (N_22240,N_16484,N_15879);
nand U22241 (N_22241,N_17093,N_16354);
and U22242 (N_22242,N_15343,N_15967);
xnor U22243 (N_22243,N_15181,N_17693);
nand U22244 (N_22244,N_15005,N_19115);
nor U22245 (N_22245,N_18295,N_19487);
nand U22246 (N_22246,N_19109,N_19249);
nor U22247 (N_22247,N_18719,N_18138);
nor U22248 (N_22248,N_19765,N_19318);
and U22249 (N_22249,N_17746,N_18271);
and U22250 (N_22250,N_19462,N_19397);
and U22251 (N_22251,N_18466,N_15008);
or U22252 (N_22252,N_16802,N_19685);
or U22253 (N_22253,N_17448,N_16374);
nand U22254 (N_22254,N_16309,N_15248);
xor U22255 (N_22255,N_15031,N_17864);
or U22256 (N_22256,N_15653,N_19016);
nand U22257 (N_22257,N_16433,N_18157);
nand U22258 (N_22258,N_17707,N_15562);
and U22259 (N_22259,N_16964,N_15536);
nor U22260 (N_22260,N_17694,N_15168);
nor U22261 (N_22261,N_18564,N_15446);
and U22262 (N_22262,N_17546,N_17643);
nand U22263 (N_22263,N_15588,N_17883);
or U22264 (N_22264,N_18761,N_15812);
and U22265 (N_22265,N_15702,N_19957);
nor U22266 (N_22266,N_19744,N_18592);
nand U22267 (N_22267,N_17347,N_15180);
or U22268 (N_22268,N_19131,N_17015);
or U22269 (N_22269,N_18025,N_16579);
xnor U22270 (N_22270,N_19116,N_17357);
nor U22271 (N_22271,N_16301,N_17041);
xor U22272 (N_22272,N_17133,N_18875);
xnor U22273 (N_22273,N_19780,N_19905);
or U22274 (N_22274,N_16830,N_18658);
nand U22275 (N_22275,N_18890,N_19935);
or U22276 (N_22276,N_19277,N_17930);
xnor U22277 (N_22277,N_15340,N_15044);
or U22278 (N_22278,N_17777,N_15114);
and U22279 (N_22279,N_17584,N_17611);
and U22280 (N_22280,N_19534,N_19805);
nand U22281 (N_22281,N_19833,N_18567);
nand U22282 (N_22282,N_18063,N_19228);
xnor U22283 (N_22283,N_15136,N_15036);
or U22284 (N_22284,N_19782,N_19440);
xnor U22285 (N_22285,N_18015,N_18765);
or U22286 (N_22286,N_17804,N_17681);
and U22287 (N_22287,N_17134,N_19355);
and U22288 (N_22288,N_17801,N_19989);
nor U22289 (N_22289,N_19438,N_17400);
xnor U22290 (N_22290,N_17126,N_17780);
or U22291 (N_22291,N_15885,N_15309);
and U22292 (N_22292,N_19789,N_19407);
xnor U22293 (N_22293,N_16587,N_18451);
nor U22294 (N_22294,N_18327,N_18505);
nand U22295 (N_22295,N_15966,N_17897);
and U22296 (N_22296,N_19941,N_15685);
and U22297 (N_22297,N_15565,N_19998);
nor U22298 (N_22298,N_15024,N_18518);
and U22299 (N_22299,N_17905,N_16165);
and U22300 (N_22300,N_16025,N_17810);
xnor U22301 (N_22301,N_15931,N_17716);
nor U22302 (N_22302,N_16844,N_19173);
and U22303 (N_22303,N_17332,N_19361);
and U22304 (N_22304,N_19070,N_19345);
nor U22305 (N_22305,N_19052,N_15538);
nor U22306 (N_22306,N_18364,N_19427);
nand U22307 (N_22307,N_15208,N_16892);
xnor U22308 (N_22308,N_19197,N_19960);
xnor U22309 (N_22309,N_17626,N_18531);
nor U22310 (N_22310,N_15010,N_19263);
or U22311 (N_22311,N_19479,N_15894);
nor U22312 (N_22312,N_15054,N_16542);
nand U22313 (N_22313,N_19871,N_19851);
nor U22314 (N_22314,N_18014,N_18580);
or U22315 (N_22315,N_15655,N_18390);
xnor U22316 (N_22316,N_17318,N_18049);
and U22317 (N_22317,N_16001,N_15921);
and U22318 (N_22318,N_17534,N_19706);
nor U22319 (N_22319,N_17194,N_17590);
and U22320 (N_22320,N_18756,N_16836);
nor U22321 (N_22321,N_17954,N_16888);
and U22322 (N_22322,N_18105,N_16613);
xnor U22323 (N_22323,N_15932,N_15937);
and U22324 (N_22324,N_18855,N_19830);
and U22325 (N_22325,N_18113,N_17208);
and U22326 (N_22326,N_16823,N_16439);
or U22327 (N_22327,N_18954,N_18179);
nand U22328 (N_22328,N_18437,N_15438);
nand U22329 (N_22329,N_19945,N_16679);
xnor U22330 (N_22330,N_18690,N_19204);
xor U22331 (N_22331,N_15424,N_18955);
xor U22332 (N_22332,N_16477,N_16555);
or U22333 (N_22333,N_18906,N_17218);
or U22334 (N_22334,N_17010,N_19646);
xor U22335 (N_22335,N_15379,N_16730);
nor U22336 (N_22336,N_15344,N_15033);
nor U22337 (N_22337,N_19100,N_15225);
or U22338 (N_22338,N_16290,N_18848);
or U22339 (N_22339,N_18009,N_15462);
xor U22340 (N_22340,N_18998,N_19615);
nor U22341 (N_22341,N_16561,N_17561);
nor U22342 (N_22342,N_15747,N_19105);
nand U22343 (N_22343,N_17617,N_18258);
nor U22344 (N_22344,N_18821,N_16387);
xnor U22345 (N_22345,N_15237,N_19367);
nand U22346 (N_22346,N_18406,N_16029);
or U22347 (N_22347,N_15075,N_16674);
xor U22348 (N_22348,N_16650,N_15252);
nand U22349 (N_22349,N_15097,N_15525);
or U22350 (N_22350,N_18198,N_19728);
or U22351 (N_22351,N_18043,N_17751);
nor U22352 (N_22352,N_19211,N_19276);
nand U22353 (N_22353,N_19257,N_16508);
xnor U22354 (N_22354,N_16622,N_18124);
xnor U22355 (N_22355,N_15217,N_17711);
or U22356 (N_22356,N_19799,N_15003);
nor U22357 (N_22357,N_16863,N_19984);
nand U22358 (N_22358,N_18277,N_16231);
xnor U22359 (N_22359,N_18624,N_15764);
nor U22360 (N_22360,N_19056,N_19287);
nor U22361 (N_22361,N_17454,N_19113);
or U22362 (N_22362,N_16570,N_17734);
nand U22363 (N_22363,N_17166,N_19480);
nand U22364 (N_22364,N_15874,N_16398);
nor U22365 (N_22365,N_17042,N_17142);
xor U22366 (N_22366,N_19723,N_18494);
and U22367 (N_22367,N_19389,N_16400);
nor U22368 (N_22368,N_19573,N_18405);
or U22369 (N_22369,N_16909,N_19604);
or U22370 (N_22370,N_16323,N_16207);
nand U22371 (N_22371,N_18968,N_18435);
xnor U22372 (N_22372,N_18382,N_19922);
or U22373 (N_22373,N_19693,N_19526);
xnor U22374 (N_22374,N_19626,N_15480);
nand U22375 (N_22375,N_19320,N_17482);
nor U22376 (N_22376,N_17461,N_18532);
nand U22377 (N_22377,N_17479,N_15837);
and U22378 (N_22378,N_17593,N_18262);
or U22379 (N_22379,N_16437,N_19119);
and U22380 (N_22380,N_18630,N_19947);
xor U22381 (N_22381,N_17038,N_18779);
nand U22382 (N_22382,N_19409,N_19006);
and U22383 (N_22383,N_17787,N_15870);
nand U22384 (N_22384,N_19520,N_18724);
or U22385 (N_22385,N_19629,N_19664);
nor U22386 (N_22386,N_17242,N_17426);
or U22387 (N_22387,N_17375,N_18594);
or U22388 (N_22388,N_19624,N_16300);
and U22389 (N_22389,N_17013,N_19907);
nor U22390 (N_22390,N_15339,N_16694);
and U22391 (N_22391,N_19171,N_15703);
nor U22392 (N_22392,N_17228,N_16161);
nor U22393 (N_22393,N_19538,N_17463);
xor U22394 (N_22394,N_18748,N_15435);
xor U22395 (N_22395,N_16237,N_16341);
nand U22396 (N_22396,N_15151,N_18182);
nor U22397 (N_22397,N_15491,N_15076);
nor U22398 (N_22398,N_19091,N_17486);
nor U22399 (N_22399,N_15798,N_19687);
and U22400 (N_22400,N_18860,N_18445);
xor U22401 (N_22401,N_18259,N_16221);
or U22402 (N_22402,N_17622,N_16501);
nand U22403 (N_22403,N_16966,N_17201);
xnor U22404 (N_22404,N_19206,N_17723);
nor U22405 (N_22405,N_15952,N_17652);
xor U22406 (N_22406,N_17381,N_16461);
xnor U22407 (N_22407,N_18850,N_19365);
nand U22408 (N_22408,N_16232,N_15350);
and U22409 (N_22409,N_19323,N_17671);
and U22410 (N_22410,N_16244,N_18579);
and U22411 (N_22411,N_18315,N_15386);
or U22412 (N_22412,N_16842,N_19494);
or U22413 (N_22413,N_15465,N_15275);
and U22414 (N_22414,N_19231,N_16691);
nand U22415 (N_22415,N_16875,N_17772);
and U22416 (N_22416,N_15122,N_19681);
nor U22417 (N_22417,N_19370,N_17363);
and U22418 (N_22418,N_17782,N_18287);
or U22419 (N_22419,N_15203,N_17251);
xor U22420 (N_22420,N_18541,N_17682);
or U22421 (N_22421,N_16417,N_18738);
or U22422 (N_22422,N_18431,N_16744);
nor U22423 (N_22423,N_17717,N_16425);
and U22424 (N_22424,N_19959,N_18280);
or U22425 (N_22425,N_15585,N_16662);
or U22426 (N_22426,N_17219,N_19980);
nor U22427 (N_22427,N_19068,N_18354);
xor U22428 (N_22428,N_16440,N_19645);
and U22429 (N_22429,N_18517,N_18809);
nor U22430 (N_22430,N_16061,N_16769);
or U22431 (N_22431,N_18330,N_15939);
nand U22432 (N_22432,N_18749,N_16535);
nand U22433 (N_22433,N_18482,N_15833);
and U22434 (N_22434,N_18721,N_17951);
and U22435 (N_22435,N_16891,N_18366);
and U22436 (N_22436,N_18409,N_18016);
nor U22437 (N_22437,N_16131,N_18026);
or U22438 (N_22438,N_15990,N_15630);
or U22439 (N_22439,N_18653,N_16943);
nand U22440 (N_22440,N_18854,N_16728);
nor U22441 (N_22441,N_15986,N_18102);
xor U22442 (N_22442,N_18173,N_15782);
xor U22443 (N_22443,N_16809,N_19787);
xor U22444 (N_22444,N_18369,N_15042);
nor U22445 (N_22445,N_18477,N_19046);
nor U22446 (N_22446,N_17105,N_19704);
nor U22447 (N_22447,N_18570,N_15159);
and U22448 (N_22448,N_16109,N_19200);
xor U22449 (N_22449,N_18448,N_17339);
or U22450 (N_22450,N_16788,N_17975);
xnor U22451 (N_22451,N_17958,N_15897);
nand U22452 (N_22452,N_18785,N_17309);
and U22453 (N_22453,N_17972,N_18289);
or U22454 (N_22454,N_18399,N_19341);
nand U22455 (N_22455,N_17631,N_19081);
and U22456 (N_22456,N_18365,N_19253);
xnor U22457 (N_22457,N_18743,N_19405);
nor U22458 (N_22458,N_19123,N_16592);
or U22459 (N_22459,N_17145,N_17298);
nor U22460 (N_22460,N_19110,N_16490);
nand U22461 (N_22461,N_16475,N_16000);
and U22462 (N_22462,N_15636,N_16100);
and U22463 (N_22463,N_18306,N_17441);
xnor U22464 (N_22464,N_15947,N_16299);
nand U22465 (N_22465,N_16793,N_18145);
and U22466 (N_22466,N_17058,N_16717);
nor U22467 (N_22467,N_16269,N_19575);
or U22468 (N_22468,N_18991,N_16753);
nor U22469 (N_22469,N_18846,N_15450);
xnor U22470 (N_22470,N_19825,N_18618);
nand U22471 (N_22471,N_19224,N_16471);
and U22472 (N_22472,N_15120,N_15152);
nor U22473 (N_22473,N_19020,N_17327);
and U22474 (N_22474,N_19454,N_19899);
nand U22475 (N_22475,N_19610,N_15341);
or U22476 (N_22476,N_18302,N_16438);
and U22477 (N_22477,N_16988,N_16710);
or U22478 (N_22478,N_15578,N_18747);
and U22479 (N_22479,N_16913,N_18376);
xnor U22480 (N_22480,N_19719,N_19310);
and U22481 (N_22481,N_16464,N_16867);
and U22482 (N_22482,N_15051,N_18397);
xnor U22483 (N_22483,N_16327,N_17411);
nand U22484 (N_22484,N_18934,N_15689);
xnor U22485 (N_22485,N_18842,N_18089);
nand U22486 (N_22486,N_17107,N_19149);
or U22487 (N_22487,N_15374,N_16724);
or U22488 (N_22488,N_16436,N_19227);
nand U22489 (N_22489,N_16190,N_16734);
xor U22490 (N_22490,N_19458,N_18344);
or U22491 (N_22491,N_15432,N_18002);
nand U22492 (N_22492,N_15357,N_18115);
xnor U22493 (N_22493,N_15579,N_16418);
or U22494 (N_22494,N_17312,N_16266);
nand U22495 (N_22495,N_17139,N_15219);
or U22496 (N_22496,N_18116,N_17889);
xnor U22497 (N_22497,N_17040,N_17004);
nor U22498 (N_22498,N_18057,N_18086);
xor U22499 (N_22499,N_19943,N_19903);
or U22500 (N_22500,N_17628,N_15115);
nor U22501 (N_22501,N_17305,N_15211);
and U22502 (N_22502,N_18625,N_15585);
nand U22503 (N_22503,N_19296,N_17413);
nand U22504 (N_22504,N_18386,N_19500);
nor U22505 (N_22505,N_17107,N_16052);
xnor U22506 (N_22506,N_17415,N_17323);
xnor U22507 (N_22507,N_19747,N_17332);
xnor U22508 (N_22508,N_16495,N_19411);
and U22509 (N_22509,N_18304,N_15269);
nor U22510 (N_22510,N_17015,N_17201);
xnor U22511 (N_22511,N_15323,N_18407);
xnor U22512 (N_22512,N_17155,N_18927);
nand U22513 (N_22513,N_17162,N_19742);
nor U22514 (N_22514,N_18757,N_19449);
xnor U22515 (N_22515,N_19361,N_19464);
nand U22516 (N_22516,N_19338,N_16065);
nand U22517 (N_22517,N_18976,N_17419);
nand U22518 (N_22518,N_17509,N_18114);
xor U22519 (N_22519,N_17147,N_17087);
xnor U22520 (N_22520,N_16658,N_17805);
nand U22521 (N_22521,N_16036,N_19395);
nor U22522 (N_22522,N_16707,N_19245);
nand U22523 (N_22523,N_19653,N_19649);
nor U22524 (N_22524,N_19281,N_17796);
or U22525 (N_22525,N_17330,N_16724);
nand U22526 (N_22526,N_18370,N_16051);
and U22527 (N_22527,N_19143,N_19867);
nor U22528 (N_22528,N_19612,N_16240);
or U22529 (N_22529,N_17660,N_16532);
and U22530 (N_22530,N_16511,N_16970);
xnor U22531 (N_22531,N_17144,N_17134);
and U22532 (N_22532,N_15224,N_17301);
nand U22533 (N_22533,N_19620,N_17619);
nor U22534 (N_22534,N_19483,N_17595);
and U22535 (N_22535,N_19487,N_15855);
or U22536 (N_22536,N_16445,N_16382);
and U22537 (N_22537,N_19635,N_15088);
nand U22538 (N_22538,N_18606,N_16942);
nor U22539 (N_22539,N_19895,N_18602);
nor U22540 (N_22540,N_15152,N_15593);
and U22541 (N_22541,N_16406,N_16385);
or U22542 (N_22542,N_15953,N_19962);
or U22543 (N_22543,N_18703,N_19115);
or U22544 (N_22544,N_18232,N_17209);
nand U22545 (N_22545,N_19182,N_19753);
nor U22546 (N_22546,N_15062,N_19067);
nor U22547 (N_22547,N_18208,N_18395);
xnor U22548 (N_22548,N_18359,N_16640);
and U22549 (N_22549,N_15294,N_18333);
xnor U22550 (N_22550,N_18390,N_17510);
or U22551 (N_22551,N_15564,N_15247);
xor U22552 (N_22552,N_19418,N_16136);
nor U22553 (N_22553,N_19998,N_15358);
or U22554 (N_22554,N_17132,N_18282);
xnor U22555 (N_22555,N_19277,N_15021);
or U22556 (N_22556,N_18198,N_18836);
nand U22557 (N_22557,N_15572,N_17470);
or U22558 (N_22558,N_15127,N_18202);
nand U22559 (N_22559,N_15105,N_16960);
nand U22560 (N_22560,N_15199,N_17836);
nand U22561 (N_22561,N_19392,N_18637);
and U22562 (N_22562,N_18358,N_19965);
xnor U22563 (N_22563,N_18278,N_16327);
xnor U22564 (N_22564,N_15834,N_18272);
and U22565 (N_22565,N_17129,N_19951);
xor U22566 (N_22566,N_16240,N_19917);
or U22567 (N_22567,N_19977,N_16231);
nand U22568 (N_22568,N_18259,N_17136);
nand U22569 (N_22569,N_15583,N_19471);
or U22570 (N_22570,N_18374,N_19683);
or U22571 (N_22571,N_15117,N_15959);
or U22572 (N_22572,N_17820,N_17493);
xor U22573 (N_22573,N_19836,N_17991);
xnor U22574 (N_22574,N_17201,N_18694);
xnor U22575 (N_22575,N_18416,N_15846);
and U22576 (N_22576,N_17652,N_18094);
or U22577 (N_22577,N_16276,N_15248);
xor U22578 (N_22578,N_15871,N_19700);
or U22579 (N_22579,N_18932,N_19022);
xor U22580 (N_22580,N_15405,N_15465);
or U22581 (N_22581,N_15372,N_17657);
nand U22582 (N_22582,N_17377,N_15015);
nand U22583 (N_22583,N_15248,N_16587);
nor U22584 (N_22584,N_16504,N_15776);
nor U22585 (N_22585,N_18309,N_19075);
or U22586 (N_22586,N_17735,N_19764);
nand U22587 (N_22587,N_19775,N_15241);
xnor U22588 (N_22588,N_18477,N_16357);
nor U22589 (N_22589,N_18381,N_18978);
or U22590 (N_22590,N_18355,N_18831);
xor U22591 (N_22591,N_16137,N_17365);
xnor U22592 (N_22592,N_17594,N_17466);
nand U22593 (N_22593,N_15261,N_15572);
xnor U22594 (N_22594,N_18435,N_16111);
nand U22595 (N_22595,N_15528,N_15062);
or U22596 (N_22596,N_18290,N_18103);
and U22597 (N_22597,N_18964,N_15470);
xnor U22598 (N_22598,N_18690,N_19651);
and U22599 (N_22599,N_15143,N_16862);
nor U22600 (N_22600,N_15120,N_18776);
or U22601 (N_22601,N_16329,N_15801);
nor U22602 (N_22602,N_15332,N_16208);
nor U22603 (N_22603,N_19695,N_17229);
and U22604 (N_22604,N_17500,N_19648);
nor U22605 (N_22605,N_18281,N_16640);
nand U22606 (N_22606,N_19912,N_18921);
or U22607 (N_22607,N_18714,N_17303);
nor U22608 (N_22608,N_18237,N_16929);
or U22609 (N_22609,N_18604,N_18611);
nor U22610 (N_22610,N_17895,N_16292);
nor U22611 (N_22611,N_16151,N_16197);
xor U22612 (N_22612,N_17164,N_19662);
and U22613 (N_22613,N_18239,N_19426);
nand U22614 (N_22614,N_15544,N_19212);
xor U22615 (N_22615,N_16734,N_16375);
and U22616 (N_22616,N_19616,N_15744);
nor U22617 (N_22617,N_15033,N_16106);
nor U22618 (N_22618,N_16137,N_16035);
and U22619 (N_22619,N_19479,N_18526);
and U22620 (N_22620,N_17652,N_19317);
or U22621 (N_22621,N_19616,N_15507);
xnor U22622 (N_22622,N_15914,N_18397);
nand U22623 (N_22623,N_15883,N_19775);
xor U22624 (N_22624,N_18269,N_15022);
nor U22625 (N_22625,N_18721,N_17886);
nor U22626 (N_22626,N_16136,N_18678);
and U22627 (N_22627,N_16269,N_16591);
and U22628 (N_22628,N_16230,N_17363);
or U22629 (N_22629,N_18436,N_15408);
nand U22630 (N_22630,N_17632,N_16632);
xor U22631 (N_22631,N_19928,N_18863);
or U22632 (N_22632,N_17666,N_17946);
or U22633 (N_22633,N_16807,N_15886);
nor U22634 (N_22634,N_19089,N_18848);
and U22635 (N_22635,N_16053,N_18286);
or U22636 (N_22636,N_19588,N_17832);
xor U22637 (N_22637,N_16864,N_19913);
xnor U22638 (N_22638,N_15555,N_17905);
nand U22639 (N_22639,N_17329,N_19211);
or U22640 (N_22640,N_19142,N_19127);
or U22641 (N_22641,N_19546,N_15364);
xnor U22642 (N_22642,N_17385,N_18912);
xor U22643 (N_22643,N_17870,N_15558);
and U22644 (N_22644,N_19643,N_16466);
xor U22645 (N_22645,N_17568,N_19549);
nand U22646 (N_22646,N_19961,N_18239);
and U22647 (N_22647,N_19559,N_15127);
nor U22648 (N_22648,N_16880,N_15426);
and U22649 (N_22649,N_19066,N_17241);
nand U22650 (N_22650,N_19667,N_17357);
nand U22651 (N_22651,N_16051,N_19100);
or U22652 (N_22652,N_19773,N_17072);
nor U22653 (N_22653,N_17738,N_16226);
nand U22654 (N_22654,N_16757,N_18045);
nand U22655 (N_22655,N_16733,N_17736);
and U22656 (N_22656,N_16667,N_16551);
xnor U22657 (N_22657,N_19165,N_16337);
and U22658 (N_22658,N_18729,N_17520);
or U22659 (N_22659,N_17938,N_17029);
nor U22660 (N_22660,N_15405,N_15834);
nand U22661 (N_22661,N_16393,N_19159);
or U22662 (N_22662,N_16341,N_18442);
or U22663 (N_22663,N_19417,N_16540);
or U22664 (N_22664,N_15848,N_16223);
xnor U22665 (N_22665,N_18981,N_17353);
nand U22666 (N_22666,N_15270,N_17198);
nand U22667 (N_22667,N_18161,N_18230);
xnor U22668 (N_22668,N_16379,N_17707);
nand U22669 (N_22669,N_17980,N_19628);
xor U22670 (N_22670,N_18016,N_15022);
or U22671 (N_22671,N_15822,N_19992);
and U22672 (N_22672,N_17551,N_19859);
nand U22673 (N_22673,N_17711,N_18577);
xnor U22674 (N_22674,N_16640,N_17623);
xor U22675 (N_22675,N_15455,N_18647);
and U22676 (N_22676,N_18013,N_19854);
and U22677 (N_22677,N_16658,N_15810);
xnor U22678 (N_22678,N_17722,N_19724);
xnor U22679 (N_22679,N_19008,N_18241);
and U22680 (N_22680,N_18482,N_17121);
xor U22681 (N_22681,N_19208,N_16080);
or U22682 (N_22682,N_15836,N_16754);
or U22683 (N_22683,N_16566,N_19551);
nor U22684 (N_22684,N_15882,N_15923);
nor U22685 (N_22685,N_17845,N_19855);
xor U22686 (N_22686,N_19264,N_16386);
nand U22687 (N_22687,N_17209,N_18325);
nand U22688 (N_22688,N_18943,N_19811);
or U22689 (N_22689,N_15846,N_16620);
xnor U22690 (N_22690,N_16338,N_15539);
and U22691 (N_22691,N_19870,N_15652);
nand U22692 (N_22692,N_16914,N_16152);
nand U22693 (N_22693,N_15908,N_15565);
nand U22694 (N_22694,N_19244,N_16669);
nor U22695 (N_22695,N_17071,N_16098);
nand U22696 (N_22696,N_19414,N_16996);
nor U22697 (N_22697,N_16263,N_15514);
nor U22698 (N_22698,N_18415,N_16658);
nand U22699 (N_22699,N_16147,N_15755);
nor U22700 (N_22700,N_19326,N_18820);
nand U22701 (N_22701,N_19759,N_19286);
nor U22702 (N_22702,N_17069,N_15358);
nand U22703 (N_22703,N_16612,N_19745);
nor U22704 (N_22704,N_19668,N_19600);
xnor U22705 (N_22705,N_16757,N_17310);
or U22706 (N_22706,N_15248,N_17720);
or U22707 (N_22707,N_19856,N_15964);
or U22708 (N_22708,N_17635,N_16506);
nor U22709 (N_22709,N_19411,N_16428);
nand U22710 (N_22710,N_19864,N_19338);
nor U22711 (N_22711,N_15593,N_19785);
nor U22712 (N_22712,N_17105,N_17967);
and U22713 (N_22713,N_17195,N_16871);
nor U22714 (N_22714,N_19366,N_16596);
nor U22715 (N_22715,N_19594,N_17897);
and U22716 (N_22716,N_15445,N_19100);
nor U22717 (N_22717,N_19152,N_18340);
or U22718 (N_22718,N_15780,N_16833);
and U22719 (N_22719,N_15763,N_17877);
and U22720 (N_22720,N_17649,N_19723);
xor U22721 (N_22721,N_16148,N_18666);
nor U22722 (N_22722,N_16514,N_15722);
xnor U22723 (N_22723,N_18910,N_19954);
nand U22724 (N_22724,N_16784,N_15827);
nand U22725 (N_22725,N_17748,N_16694);
and U22726 (N_22726,N_15777,N_19306);
and U22727 (N_22727,N_18729,N_17333);
nand U22728 (N_22728,N_18569,N_16199);
and U22729 (N_22729,N_19486,N_17917);
or U22730 (N_22730,N_17101,N_18008);
nor U22731 (N_22731,N_17881,N_18884);
nand U22732 (N_22732,N_19915,N_16096);
xnor U22733 (N_22733,N_17588,N_18694);
or U22734 (N_22734,N_15533,N_16547);
or U22735 (N_22735,N_15645,N_19179);
nor U22736 (N_22736,N_15743,N_18068);
xor U22737 (N_22737,N_19851,N_17544);
or U22738 (N_22738,N_18962,N_19688);
xor U22739 (N_22739,N_15489,N_15364);
nor U22740 (N_22740,N_17688,N_18662);
or U22741 (N_22741,N_17451,N_18059);
nand U22742 (N_22742,N_19306,N_16143);
and U22743 (N_22743,N_17582,N_19768);
nand U22744 (N_22744,N_19782,N_15361);
nand U22745 (N_22745,N_16416,N_16219);
and U22746 (N_22746,N_16630,N_18262);
nor U22747 (N_22747,N_15042,N_15957);
xnor U22748 (N_22748,N_17540,N_19098);
nand U22749 (N_22749,N_16450,N_15517);
or U22750 (N_22750,N_15246,N_16195);
nor U22751 (N_22751,N_19245,N_19394);
and U22752 (N_22752,N_18832,N_17789);
nand U22753 (N_22753,N_15678,N_19642);
nor U22754 (N_22754,N_15226,N_15822);
xor U22755 (N_22755,N_19253,N_15063);
nor U22756 (N_22756,N_16664,N_16377);
nand U22757 (N_22757,N_15980,N_19203);
and U22758 (N_22758,N_17366,N_18492);
and U22759 (N_22759,N_19432,N_15754);
or U22760 (N_22760,N_18074,N_19910);
nor U22761 (N_22761,N_16892,N_19204);
and U22762 (N_22762,N_16946,N_19388);
nand U22763 (N_22763,N_16087,N_18687);
nand U22764 (N_22764,N_15994,N_17642);
or U22765 (N_22765,N_18530,N_15731);
or U22766 (N_22766,N_15135,N_19942);
and U22767 (N_22767,N_19248,N_19505);
xnor U22768 (N_22768,N_17833,N_19937);
xnor U22769 (N_22769,N_17748,N_15709);
xnor U22770 (N_22770,N_16650,N_19670);
nand U22771 (N_22771,N_17756,N_19375);
nand U22772 (N_22772,N_15152,N_19597);
nor U22773 (N_22773,N_16009,N_17812);
xor U22774 (N_22774,N_18574,N_17358);
nor U22775 (N_22775,N_18690,N_18737);
or U22776 (N_22776,N_17388,N_17757);
and U22777 (N_22777,N_16070,N_15417);
xor U22778 (N_22778,N_19329,N_19835);
nor U22779 (N_22779,N_16546,N_19875);
xnor U22780 (N_22780,N_18648,N_17873);
nor U22781 (N_22781,N_18970,N_15286);
or U22782 (N_22782,N_17276,N_15706);
nor U22783 (N_22783,N_18882,N_19107);
or U22784 (N_22784,N_18381,N_16472);
nand U22785 (N_22785,N_17961,N_16720);
or U22786 (N_22786,N_15006,N_16862);
nor U22787 (N_22787,N_18920,N_15547);
nor U22788 (N_22788,N_17816,N_17284);
nand U22789 (N_22789,N_18595,N_16103);
xnor U22790 (N_22790,N_19070,N_16032);
and U22791 (N_22791,N_19003,N_19844);
nor U22792 (N_22792,N_19778,N_17303);
xnor U22793 (N_22793,N_19807,N_15468);
and U22794 (N_22794,N_17233,N_15955);
nor U22795 (N_22795,N_16419,N_16437);
xnor U22796 (N_22796,N_15544,N_19214);
xnor U22797 (N_22797,N_15427,N_18931);
and U22798 (N_22798,N_15853,N_19011);
nor U22799 (N_22799,N_18168,N_19641);
nand U22800 (N_22800,N_18586,N_16689);
or U22801 (N_22801,N_17838,N_15598);
xor U22802 (N_22802,N_18263,N_16868);
and U22803 (N_22803,N_18630,N_17488);
nand U22804 (N_22804,N_18585,N_18492);
nand U22805 (N_22805,N_18563,N_16040);
xor U22806 (N_22806,N_17420,N_19319);
xnor U22807 (N_22807,N_18253,N_17666);
and U22808 (N_22808,N_17323,N_15741);
or U22809 (N_22809,N_19392,N_19485);
or U22810 (N_22810,N_18528,N_15480);
nor U22811 (N_22811,N_18850,N_17115);
or U22812 (N_22812,N_16607,N_16333);
nand U22813 (N_22813,N_18154,N_15268);
or U22814 (N_22814,N_15190,N_19210);
or U22815 (N_22815,N_15255,N_17916);
or U22816 (N_22816,N_19620,N_16272);
or U22817 (N_22817,N_19197,N_15081);
or U22818 (N_22818,N_15718,N_18735);
xor U22819 (N_22819,N_15335,N_15280);
or U22820 (N_22820,N_18923,N_15275);
and U22821 (N_22821,N_17048,N_18292);
nor U22822 (N_22822,N_15952,N_19314);
or U22823 (N_22823,N_18729,N_18865);
nor U22824 (N_22824,N_15755,N_17240);
xor U22825 (N_22825,N_18349,N_15182);
or U22826 (N_22826,N_19959,N_16845);
nor U22827 (N_22827,N_16140,N_19179);
nor U22828 (N_22828,N_18989,N_17261);
nor U22829 (N_22829,N_19950,N_15260);
nor U22830 (N_22830,N_19505,N_17571);
nand U22831 (N_22831,N_16377,N_17843);
nand U22832 (N_22832,N_17175,N_17186);
and U22833 (N_22833,N_16682,N_18419);
nand U22834 (N_22834,N_16044,N_17785);
nand U22835 (N_22835,N_16829,N_19576);
nor U22836 (N_22836,N_18629,N_15997);
nand U22837 (N_22837,N_17175,N_19956);
xnor U22838 (N_22838,N_19470,N_17995);
xnor U22839 (N_22839,N_16438,N_17210);
nand U22840 (N_22840,N_18172,N_19979);
xnor U22841 (N_22841,N_18738,N_15468);
and U22842 (N_22842,N_19812,N_18807);
nand U22843 (N_22843,N_18795,N_19517);
nand U22844 (N_22844,N_15250,N_16019);
xor U22845 (N_22845,N_19032,N_15776);
or U22846 (N_22846,N_18461,N_18418);
and U22847 (N_22847,N_17244,N_16375);
nand U22848 (N_22848,N_18427,N_16386);
xnor U22849 (N_22849,N_15856,N_18897);
or U22850 (N_22850,N_15172,N_19969);
nor U22851 (N_22851,N_19064,N_15610);
xor U22852 (N_22852,N_17651,N_19239);
and U22853 (N_22853,N_16341,N_15699);
and U22854 (N_22854,N_16100,N_18821);
xor U22855 (N_22855,N_19905,N_16900);
nor U22856 (N_22856,N_18644,N_19674);
and U22857 (N_22857,N_15432,N_18405);
nand U22858 (N_22858,N_19286,N_17082);
and U22859 (N_22859,N_18500,N_18489);
nand U22860 (N_22860,N_17515,N_16763);
nor U22861 (N_22861,N_18217,N_15997);
or U22862 (N_22862,N_19278,N_17778);
nor U22863 (N_22863,N_19583,N_18974);
nor U22864 (N_22864,N_18868,N_18700);
nor U22865 (N_22865,N_18241,N_16245);
or U22866 (N_22866,N_19195,N_19460);
and U22867 (N_22867,N_19641,N_16143);
nor U22868 (N_22868,N_15219,N_18868);
xnor U22869 (N_22869,N_15493,N_19381);
or U22870 (N_22870,N_17429,N_17420);
nor U22871 (N_22871,N_18715,N_19539);
xor U22872 (N_22872,N_18583,N_18850);
and U22873 (N_22873,N_18659,N_17778);
or U22874 (N_22874,N_19070,N_19323);
or U22875 (N_22875,N_15054,N_16785);
xor U22876 (N_22876,N_19506,N_15481);
and U22877 (N_22877,N_15299,N_17192);
nand U22878 (N_22878,N_18898,N_17197);
or U22879 (N_22879,N_16185,N_16587);
or U22880 (N_22880,N_15735,N_17702);
and U22881 (N_22881,N_15021,N_18481);
or U22882 (N_22882,N_16993,N_15922);
nor U22883 (N_22883,N_18066,N_16785);
or U22884 (N_22884,N_18949,N_18067);
xnor U22885 (N_22885,N_15919,N_15956);
or U22886 (N_22886,N_15820,N_17708);
xnor U22887 (N_22887,N_16351,N_19953);
and U22888 (N_22888,N_17277,N_19249);
nand U22889 (N_22889,N_17844,N_15105);
nand U22890 (N_22890,N_16780,N_19040);
xnor U22891 (N_22891,N_15389,N_17420);
nor U22892 (N_22892,N_16137,N_16435);
or U22893 (N_22893,N_19526,N_17605);
or U22894 (N_22894,N_19222,N_19278);
or U22895 (N_22895,N_17758,N_16559);
or U22896 (N_22896,N_15603,N_15693);
or U22897 (N_22897,N_16234,N_17712);
xnor U22898 (N_22898,N_17822,N_18837);
and U22899 (N_22899,N_18531,N_15713);
nand U22900 (N_22900,N_15679,N_17366);
nand U22901 (N_22901,N_15486,N_16874);
and U22902 (N_22902,N_19869,N_18084);
or U22903 (N_22903,N_17939,N_17313);
or U22904 (N_22904,N_17110,N_16033);
or U22905 (N_22905,N_19689,N_18943);
xor U22906 (N_22906,N_17941,N_15012);
nand U22907 (N_22907,N_15018,N_16229);
xnor U22908 (N_22908,N_16362,N_15954);
nor U22909 (N_22909,N_18125,N_18704);
and U22910 (N_22910,N_18827,N_15224);
nor U22911 (N_22911,N_17013,N_16396);
and U22912 (N_22912,N_15714,N_18301);
nand U22913 (N_22913,N_18663,N_15905);
nor U22914 (N_22914,N_16600,N_16531);
or U22915 (N_22915,N_18654,N_17034);
and U22916 (N_22916,N_17355,N_17778);
nand U22917 (N_22917,N_17289,N_15972);
and U22918 (N_22918,N_18207,N_18883);
or U22919 (N_22919,N_19792,N_19235);
and U22920 (N_22920,N_19630,N_17377);
or U22921 (N_22921,N_18577,N_18897);
and U22922 (N_22922,N_15682,N_19738);
and U22923 (N_22923,N_15089,N_17440);
or U22924 (N_22924,N_19326,N_16111);
nor U22925 (N_22925,N_15448,N_15432);
xnor U22926 (N_22926,N_15870,N_19679);
xnor U22927 (N_22927,N_15379,N_17955);
nor U22928 (N_22928,N_19078,N_15183);
nand U22929 (N_22929,N_15322,N_17456);
nor U22930 (N_22930,N_17619,N_18337);
nor U22931 (N_22931,N_15681,N_18536);
nand U22932 (N_22932,N_17776,N_16396);
and U22933 (N_22933,N_17308,N_16947);
and U22934 (N_22934,N_18396,N_18219);
nor U22935 (N_22935,N_15293,N_15469);
nand U22936 (N_22936,N_15007,N_15552);
xnor U22937 (N_22937,N_17026,N_17971);
and U22938 (N_22938,N_17282,N_17296);
xor U22939 (N_22939,N_18514,N_15551);
nor U22940 (N_22940,N_15055,N_19749);
xnor U22941 (N_22941,N_19963,N_15475);
nor U22942 (N_22942,N_18750,N_19129);
nor U22943 (N_22943,N_18937,N_15134);
and U22944 (N_22944,N_16040,N_16566);
nand U22945 (N_22945,N_19945,N_16204);
nor U22946 (N_22946,N_17862,N_19531);
nand U22947 (N_22947,N_16066,N_18007);
xor U22948 (N_22948,N_15199,N_19902);
xnor U22949 (N_22949,N_17919,N_17562);
xor U22950 (N_22950,N_18291,N_15977);
nand U22951 (N_22951,N_15377,N_18759);
nand U22952 (N_22952,N_17071,N_19033);
or U22953 (N_22953,N_19471,N_17248);
and U22954 (N_22954,N_15490,N_15877);
or U22955 (N_22955,N_15673,N_19398);
or U22956 (N_22956,N_19975,N_18362);
nand U22957 (N_22957,N_18778,N_18859);
nand U22958 (N_22958,N_17544,N_19936);
nand U22959 (N_22959,N_19092,N_16990);
xor U22960 (N_22960,N_19859,N_18535);
nand U22961 (N_22961,N_18896,N_18860);
or U22962 (N_22962,N_15320,N_19229);
xor U22963 (N_22963,N_19027,N_18479);
and U22964 (N_22964,N_19590,N_16694);
xor U22965 (N_22965,N_17367,N_15776);
xor U22966 (N_22966,N_19674,N_19857);
or U22967 (N_22967,N_17889,N_16808);
nand U22968 (N_22968,N_15657,N_16406);
xnor U22969 (N_22969,N_15655,N_15862);
or U22970 (N_22970,N_15224,N_19729);
nor U22971 (N_22971,N_18446,N_18097);
xnor U22972 (N_22972,N_17945,N_16108);
nand U22973 (N_22973,N_17055,N_18259);
and U22974 (N_22974,N_19352,N_18388);
nand U22975 (N_22975,N_19916,N_18538);
xnor U22976 (N_22976,N_18259,N_16930);
nand U22977 (N_22977,N_18561,N_18171);
nor U22978 (N_22978,N_18532,N_19040);
nand U22979 (N_22979,N_19570,N_17690);
xnor U22980 (N_22980,N_16531,N_16022);
xnor U22981 (N_22981,N_17346,N_17687);
xnor U22982 (N_22982,N_17337,N_16330);
nand U22983 (N_22983,N_15701,N_16642);
nand U22984 (N_22984,N_17927,N_18264);
xnor U22985 (N_22985,N_18752,N_19910);
or U22986 (N_22986,N_15214,N_16109);
xnor U22987 (N_22987,N_16681,N_15657);
nor U22988 (N_22988,N_18062,N_15764);
and U22989 (N_22989,N_17099,N_15166);
xnor U22990 (N_22990,N_16178,N_15244);
xnor U22991 (N_22991,N_16914,N_15291);
and U22992 (N_22992,N_16902,N_18848);
nand U22993 (N_22993,N_19101,N_17880);
nor U22994 (N_22994,N_19786,N_17868);
nor U22995 (N_22995,N_18041,N_19427);
nor U22996 (N_22996,N_16094,N_16402);
and U22997 (N_22997,N_19277,N_16948);
xnor U22998 (N_22998,N_16014,N_15040);
xnor U22999 (N_22999,N_15851,N_16387);
nor U23000 (N_23000,N_18061,N_15371);
xor U23001 (N_23001,N_18320,N_15284);
nand U23002 (N_23002,N_16577,N_18696);
or U23003 (N_23003,N_15261,N_17571);
nor U23004 (N_23004,N_18780,N_18689);
or U23005 (N_23005,N_16097,N_16836);
or U23006 (N_23006,N_18758,N_16860);
nand U23007 (N_23007,N_18163,N_15352);
nand U23008 (N_23008,N_17839,N_19038);
or U23009 (N_23009,N_16874,N_16396);
xor U23010 (N_23010,N_19898,N_18878);
and U23011 (N_23011,N_19078,N_17685);
or U23012 (N_23012,N_18141,N_16236);
xor U23013 (N_23013,N_19191,N_16782);
xor U23014 (N_23014,N_16406,N_19794);
or U23015 (N_23015,N_17666,N_16810);
nand U23016 (N_23016,N_17186,N_18372);
nor U23017 (N_23017,N_18721,N_19559);
nor U23018 (N_23018,N_16849,N_17883);
or U23019 (N_23019,N_19202,N_17560);
nor U23020 (N_23020,N_15325,N_19155);
or U23021 (N_23021,N_16247,N_16014);
nor U23022 (N_23022,N_18995,N_17590);
nand U23023 (N_23023,N_17734,N_16161);
or U23024 (N_23024,N_19419,N_15278);
or U23025 (N_23025,N_19341,N_16705);
nand U23026 (N_23026,N_15399,N_19207);
nand U23027 (N_23027,N_17985,N_17411);
or U23028 (N_23028,N_15119,N_15710);
or U23029 (N_23029,N_19776,N_15988);
xnor U23030 (N_23030,N_16501,N_17259);
or U23031 (N_23031,N_15255,N_17359);
nand U23032 (N_23032,N_18683,N_17433);
or U23033 (N_23033,N_17235,N_18434);
and U23034 (N_23034,N_19670,N_17009);
or U23035 (N_23035,N_17227,N_16204);
xor U23036 (N_23036,N_17619,N_16041);
xor U23037 (N_23037,N_16058,N_18949);
or U23038 (N_23038,N_18195,N_18290);
or U23039 (N_23039,N_18886,N_17963);
nor U23040 (N_23040,N_15569,N_16947);
or U23041 (N_23041,N_18919,N_18431);
or U23042 (N_23042,N_16295,N_16471);
or U23043 (N_23043,N_15390,N_15078);
nand U23044 (N_23044,N_18144,N_15094);
and U23045 (N_23045,N_16708,N_17764);
nor U23046 (N_23046,N_19741,N_17240);
and U23047 (N_23047,N_18394,N_15103);
nand U23048 (N_23048,N_18718,N_16572);
xor U23049 (N_23049,N_15839,N_15404);
or U23050 (N_23050,N_18484,N_16157);
nor U23051 (N_23051,N_17434,N_15506);
or U23052 (N_23052,N_17944,N_17916);
nor U23053 (N_23053,N_19519,N_17335);
nand U23054 (N_23054,N_17405,N_17590);
or U23055 (N_23055,N_15640,N_18721);
xor U23056 (N_23056,N_15133,N_19882);
nor U23057 (N_23057,N_19332,N_16911);
xor U23058 (N_23058,N_18345,N_18445);
nand U23059 (N_23059,N_16534,N_18082);
nand U23060 (N_23060,N_15353,N_17017);
and U23061 (N_23061,N_15979,N_16209);
or U23062 (N_23062,N_15949,N_16044);
nand U23063 (N_23063,N_19693,N_18551);
nand U23064 (N_23064,N_19999,N_19957);
nand U23065 (N_23065,N_19551,N_15277);
and U23066 (N_23066,N_16088,N_17458);
or U23067 (N_23067,N_15793,N_18294);
nor U23068 (N_23068,N_16901,N_19860);
nand U23069 (N_23069,N_19283,N_16669);
xnor U23070 (N_23070,N_18135,N_18043);
or U23071 (N_23071,N_18147,N_17253);
xnor U23072 (N_23072,N_17504,N_18658);
nor U23073 (N_23073,N_18998,N_18409);
and U23074 (N_23074,N_18733,N_17550);
nor U23075 (N_23075,N_15926,N_15014);
xnor U23076 (N_23076,N_18408,N_15098);
nor U23077 (N_23077,N_18582,N_18614);
nor U23078 (N_23078,N_15255,N_16146);
xnor U23079 (N_23079,N_18568,N_16766);
nor U23080 (N_23080,N_17326,N_17997);
or U23081 (N_23081,N_18535,N_18944);
xnor U23082 (N_23082,N_16132,N_15230);
nand U23083 (N_23083,N_19429,N_17889);
and U23084 (N_23084,N_17904,N_18592);
and U23085 (N_23085,N_17494,N_18799);
nand U23086 (N_23086,N_17918,N_17214);
and U23087 (N_23087,N_17730,N_16231);
xnor U23088 (N_23088,N_19075,N_18812);
and U23089 (N_23089,N_19724,N_17074);
xnor U23090 (N_23090,N_17552,N_15274);
nor U23091 (N_23091,N_18934,N_17523);
and U23092 (N_23092,N_17077,N_17400);
nor U23093 (N_23093,N_18421,N_17854);
xor U23094 (N_23094,N_15883,N_17665);
nor U23095 (N_23095,N_19975,N_15689);
or U23096 (N_23096,N_17336,N_16852);
or U23097 (N_23097,N_19900,N_15374);
nand U23098 (N_23098,N_17694,N_19751);
or U23099 (N_23099,N_18486,N_18321);
or U23100 (N_23100,N_16055,N_19390);
nand U23101 (N_23101,N_18146,N_18984);
nand U23102 (N_23102,N_17204,N_16907);
nand U23103 (N_23103,N_17667,N_18786);
and U23104 (N_23104,N_19469,N_17565);
nor U23105 (N_23105,N_18373,N_16008);
xnor U23106 (N_23106,N_19614,N_18101);
nand U23107 (N_23107,N_16269,N_15901);
and U23108 (N_23108,N_15331,N_16520);
nor U23109 (N_23109,N_19788,N_15863);
nand U23110 (N_23110,N_19986,N_15784);
xor U23111 (N_23111,N_17766,N_16068);
nand U23112 (N_23112,N_16418,N_16333);
xnor U23113 (N_23113,N_16730,N_16812);
nand U23114 (N_23114,N_15599,N_15096);
nand U23115 (N_23115,N_15191,N_19779);
xnor U23116 (N_23116,N_16885,N_19377);
and U23117 (N_23117,N_18721,N_19997);
nor U23118 (N_23118,N_17483,N_15751);
and U23119 (N_23119,N_17752,N_19075);
xnor U23120 (N_23120,N_18388,N_15076);
or U23121 (N_23121,N_19497,N_17816);
nand U23122 (N_23122,N_17447,N_15543);
nor U23123 (N_23123,N_19058,N_16733);
or U23124 (N_23124,N_18413,N_18578);
nand U23125 (N_23125,N_18739,N_19452);
nand U23126 (N_23126,N_15673,N_17389);
nor U23127 (N_23127,N_17526,N_17077);
and U23128 (N_23128,N_15072,N_15863);
or U23129 (N_23129,N_16387,N_19586);
or U23130 (N_23130,N_19387,N_17279);
nand U23131 (N_23131,N_18368,N_16089);
nand U23132 (N_23132,N_16672,N_18146);
nor U23133 (N_23133,N_19301,N_17068);
nand U23134 (N_23134,N_17632,N_18244);
nor U23135 (N_23135,N_17623,N_17842);
nand U23136 (N_23136,N_19078,N_16744);
xor U23137 (N_23137,N_15376,N_16017);
nor U23138 (N_23138,N_16538,N_17765);
nand U23139 (N_23139,N_19032,N_16230);
and U23140 (N_23140,N_18511,N_15611);
and U23141 (N_23141,N_18255,N_17815);
nor U23142 (N_23142,N_15357,N_17657);
xor U23143 (N_23143,N_19789,N_16552);
nor U23144 (N_23144,N_16513,N_19254);
and U23145 (N_23145,N_15090,N_19206);
xnor U23146 (N_23146,N_18194,N_18758);
nor U23147 (N_23147,N_19257,N_18240);
and U23148 (N_23148,N_18889,N_17685);
xnor U23149 (N_23149,N_18181,N_16715);
xor U23150 (N_23150,N_15998,N_19948);
nor U23151 (N_23151,N_16288,N_15937);
nand U23152 (N_23152,N_17858,N_17608);
xor U23153 (N_23153,N_16989,N_19836);
nor U23154 (N_23154,N_18551,N_18664);
xnor U23155 (N_23155,N_17224,N_15390);
nor U23156 (N_23156,N_15038,N_18761);
xor U23157 (N_23157,N_18357,N_15826);
nor U23158 (N_23158,N_18331,N_16508);
nand U23159 (N_23159,N_16119,N_18294);
and U23160 (N_23160,N_17122,N_19616);
nor U23161 (N_23161,N_16440,N_15499);
nand U23162 (N_23162,N_19404,N_17435);
or U23163 (N_23163,N_16543,N_18501);
nand U23164 (N_23164,N_19354,N_17736);
and U23165 (N_23165,N_16238,N_19076);
or U23166 (N_23166,N_16879,N_15845);
nand U23167 (N_23167,N_16739,N_16638);
or U23168 (N_23168,N_17136,N_18367);
and U23169 (N_23169,N_16270,N_18857);
nand U23170 (N_23170,N_16357,N_17624);
nor U23171 (N_23171,N_17443,N_16828);
nor U23172 (N_23172,N_15274,N_16729);
and U23173 (N_23173,N_16266,N_17136);
xor U23174 (N_23174,N_19105,N_18994);
nand U23175 (N_23175,N_17475,N_15403);
nor U23176 (N_23176,N_17122,N_18745);
nand U23177 (N_23177,N_15691,N_18116);
xor U23178 (N_23178,N_17008,N_18489);
nor U23179 (N_23179,N_18078,N_15356);
nor U23180 (N_23180,N_16416,N_15135);
xor U23181 (N_23181,N_16261,N_19328);
nor U23182 (N_23182,N_15444,N_18804);
and U23183 (N_23183,N_16653,N_17088);
nand U23184 (N_23184,N_18552,N_18650);
or U23185 (N_23185,N_19659,N_15999);
and U23186 (N_23186,N_17148,N_18041);
or U23187 (N_23187,N_19070,N_16559);
xor U23188 (N_23188,N_17632,N_18878);
xnor U23189 (N_23189,N_17469,N_18635);
nand U23190 (N_23190,N_17875,N_15917);
xnor U23191 (N_23191,N_18677,N_16942);
and U23192 (N_23192,N_18014,N_15569);
nand U23193 (N_23193,N_17481,N_16028);
xor U23194 (N_23194,N_19893,N_17435);
or U23195 (N_23195,N_18077,N_16552);
or U23196 (N_23196,N_18822,N_19442);
nor U23197 (N_23197,N_19209,N_16782);
nor U23198 (N_23198,N_15214,N_16418);
or U23199 (N_23199,N_17461,N_19809);
and U23200 (N_23200,N_18497,N_15052);
or U23201 (N_23201,N_16642,N_18782);
xnor U23202 (N_23202,N_16600,N_17925);
or U23203 (N_23203,N_16216,N_17272);
nand U23204 (N_23204,N_18323,N_19246);
nand U23205 (N_23205,N_18747,N_16505);
xnor U23206 (N_23206,N_18938,N_19887);
or U23207 (N_23207,N_15270,N_17876);
xnor U23208 (N_23208,N_18175,N_19651);
xor U23209 (N_23209,N_19029,N_18908);
xor U23210 (N_23210,N_16684,N_15536);
nand U23211 (N_23211,N_17845,N_17817);
nand U23212 (N_23212,N_17616,N_19622);
xnor U23213 (N_23213,N_15740,N_15148);
nand U23214 (N_23214,N_15388,N_19447);
or U23215 (N_23215,N_16889,N_19538);
and U23216 (N_23216,N_15018,N_19128);
nand U23217 (N_23217,N_18544,N_16339);
or U23218 (N_23218,N_19137,N_17977);
nand U23219 (N_23219,N_17407,N_18928);
nand U23220 (N_23220,N_19529,N_19630);
or U23221 (N_23221,N_16660,N_15326);
or U23222 (N_23222,N_18777,N_15264);
nand U23223 (N_23223,N_17423,N_16788);
nand U23224 (N_23224,N_17443,N_18717);
nor U23225 (N_23225,N_18645,N_16126);
nand U23226 (N_23226,N_18690,N_15070);
nand U23227 (N_23227,N_16355,N_17669);
nand U23228 (N_23228,N_17324,N_15411);
nor U23229 (N_23229,N_15875,N_18603);
and U23230 (N_23230,N_15132,N_17202);
and U23231 (N_23231,N_19008,N_17477);
or U23232 (N_23232,N_16427,N_16464);
or U23233 (N_23233,N_16533,N_18551);
nor U23234 (N_23234,N_17142,N_18334);
nand U23235 (N_23235,N_17930,N_16078);
xor U23236 (N_23236,N_17998,N_18032);
or U23237 (N_23237,N_16210,N_19104);
or U23238 (N_23238,N_18804,N_19454);
xnor U23239 (N_23239,N_18025,N_19510);
and U23240 (N_23240,N_19774,N_19494);
nand U23241 (N_23241,N_16223,N_19428);
and U23242 (N_23242,N_19397,N_19083);
nor U23243 (N_23243,N_15807,N_17241);
and U23244 (N_23244,N_16584,N_19238);
nand U23245 (N_23245,N_19304,N_17240);
or U23246 (N_23246,N_19070,N_19660);
and U23247 (N_23247,N_15633,N_18410);
and U23248 (N_23248,N_17683,N_17556);
nand U23249 (N_23249,N_19816,N_16030);
nor U23250 (N_23250,N_16193,N_17841);
xor U23251 (N_23251,N_16730,N_15261);
nand U23252 (N_23252,N_15233,N_17759);
xor U23253 (N_23253,N_17657,N_15635);
nor U23254 (N_23254,N_15215,N_17762);
or U23255 (N_23255,N_15068,N_16264);
and U23256 (N_23256,N_18653,N_18641);
and U23257 (N_23257,N_19102,N_18692);
nor U23258 (N_23258,N_16280,N_17680);
and U23259 (N_23259,N_17471,N_16939);
nor U23260 (N_23260,N_17596,N_19563);
xnor U23261 (N_23261,N_19225,N_17099);
nor U23262 (N_23262,N_15868,N_18312);
nor U23263 (N_23263,N_16879,N_17837);
nand U23264 (N_23264,N_19861,N_16807);
nor U23265 (N_23265,N_19953,N_18134);
and U23266 (N_23266,N_17459,N_19524);
and U23267 (N_23267,N_19830,N_16732);
and U23268 (N_23268,N_19309,N_16866);
xor U23269 (N_23269,N_15239,N_17213);
nor U23270 (N_23270,N_15597,N_15523);
xor U23271 (N_23271,N_17057,N_19658);
nor U23272 (N_23272,N_16698,N_15778);
or U23273 (N_23273,N_16420,N_17124);
and U23274 (N_23274,N_16727,N_17685);
nor U23275 (N_23275,N_16803,N_15071);
and U23276 (N_23276,N_18120,N_17392);
xor U23277 (N_23277,N_19752,N_19534);
and U23278 (N_23278,N_18643,N_18001);
and U23279 (N_23279,N_15610,N_17957);
and U23280 (N_23280,N_16403,N_17717);
and U23281 (N_23281,N_17701,N_18849);
or U23282 (N_23282,N_17438,N_17638);
nor U23283 (N_23283,N_19871,N_16908);
nor U23284 (N_23284,N_16707,N_18250);
nand U23285 (N_23285,N_19387,N_18130);
nand U23286 (N_23286,N_16889,N_17125);
nor U23287 (N_23287,N_19483,N_17861);
and U23288 (N_23288,N_15042,N_17553);
nand U23289 (N_23289,N_17614,N_16799);
xor U23290 (N_23290,N_16461,N_19925);
nor U23291 (N_23291,N_17867,N_16898);
xor U23292 (N_23292,N_18526,N_18127);
or U23293 (N_23293,N_17359,N_16946);
xnor U23294 (N_23294,N_16150,N_17416);
or U23295 (N_23295,N_18792,N_17221);
nand U23296 (N_23296,N_17390,N_17610);
or U23297 (N_23297,N_15228,N_16694);
nand U23298 (N_23298,N_17398,N_17425);
or U23299 (N_23299,N_15026,N_18288);
nand U23300 (N_23300,N_16451,N_16056);
or U23301 (N_23301,N_16810,N_15714);
nor U23302 (N_23302,N_15527,N_18879);
nor U23303 (N_23303,N_19511,N_17672);
or U23304 (N_23304,N_17864,N_16392);
xor U23305 (N_23305,N_18997,N_17624);
xnor U23306 (N_23306,N_19393,N_15621);
xor U23307 (N_23307,N_16553,N_19550);
nor U23308 (N_23308,N_16184,N_16840);
xor U23309 (N_23309,N_16957,N_16563);
nor U23310 (N_23310,N_15237,N_17738);
xnor U23311 (N_23311,N_15902,N_18054);
nor U23312 (N_23312,N_18636,N_18311);
nand U23313 (N_23313,N_19976,N_19888);
xnor U23314 (N_23314,N_17794,N_18731);
xnor U23315 (N_23315,N_15767,N_15547);
nand U23316 (N_23316,N_19659,N_17901);
or U23317 (N_23317,N_17378,N_19944);
or U23318 (N_23318,N_16642,N_15544);
and U23319 (N_23319,N_19802,N_15219);
nor U23320 (N_23320,N_18023,N_19399);
nor U23321 (N_23321,N_18668,N_18525);
xnor U23322 (N_23322,N_17806,N_17133);
and U23323 (N_23323,N_16752,N_15751);
or U23324 (N_23324,N_15215,N_16305);
nor U23325 (N_23325,N_19275,N_17463);
or U23326 (N_23326,N_18739,N_15713);
and U23327 (N_23327,N_15581,N_17446);
or U23328 (N_23328,N_19235,N_16831);
and U23329 (N_23329,N_15230,N_17646);
nor U23330 (N_23330,N_16225,N_19435);
and U23331 (N_23331,N_15040,N_19218);
or U23332 (N_23332,N_15190,N_15411);
nor U23333 (N_23333,N_15147,N_17787);
xor U23334 (N_23334,N_17525,N_15158);
and U23335 (N_23335,N_19613,N_16514);
nor U23336 (N_23336,N_18960,N_19326);
xnor U23337 (N_23337,N_15037,N_15740);
nand U23338 (N_23338,N_18056,N_18025);
xnor U23339 (N_23339,N_15807,N_19950);
xnor U23340 (N_23340,N_19298,N_16620);
and U23341 (N_23341,N_16267,N_19080);
or U23342 (N_23342,N_19581,N_16360);
xor U23343 (N_23343,N_18917,N_17429);
nand U23344 (N_23344,N_15434,N_19373);
xor U23345 (N_23345,N_18238,N_18313);
nand U23346 (N_23346,N_16157,N_19159);
nand U23347 (N_23347,N_17765,N_16276);
xnor U23348 (N_23348,N_19461,N_19477);
and U23349 (N_23349,N_18862,N_19991);
xnor U23350 (N_23350,N_16156,N_16574);
and U23351 (N_23351,N_19304,N_17101);
xor U23352 (N_23352,N_19215,N_16053);
and U23353 (N_23353,N_15718,N_19480);
xnor U23354 (N_23354,N_15254,N_19691);
or U23355 (N_23355,N_17493,N_16564);
or U23356 (N_23356,N_17526,N_17413);
xor U23357 (N_23357,N_19156,N_19600);
nand U23358 (N_23358,N_19342,N_18868);
xnor U23359 (N_23359,N_15257,N_17470);
and U23360 (N_23360,N_17815,N_16255);
or U23361 (N_23361,N_18104,N_16602);
xnor U23362 (N_23362,N_16315,N_17652);
nor U23363 (N_23363,N_19948,N_16309);
nand U23364 (N_23364,N_15847,N_18445);
and U23365 (N_23365,N_19295,N_19376);
nand U23366 (N_23366,N_15823,N_15017);
xnor U23367 (N_23367,N_19304,N_18054);
nand U23368 (N_23368,N_15439,N_16510);
nand U23369 (N_23369,N_16577,N_17117);
nand U23370 (N_23370,N_16768,N_15252);
and U23371 (N_23371,N_16930,N_16116);
or U23372 (N_23372,N_17588,N_15988);
or U23373 (N_23373,N_17928,N_16204);
xnor U23374 (N_23374,N_15898,N_15321);
or U23375 (N_23375,N_15766,N_15079);
nand U23376 (N_23376,N_17058,N_17089);
nor U23377 (N_23377,N_17752,N_17888);
nand U23378 (N_23378,N_15023,N_19488);
or U23379 (N_23379,N_17835,N_15553);
and U23380 (N_23380,N_19826,N_15493);
nor U23381 (N_23381,N_15145,N_17406);
and U23382 (N_23382,N_18523,N_15190);
or U23383 (N_23383,N_16333,N_16737);
or U23384 (N_23384,N_16322,N_17820);
nor U23385 (N_23385,N_19669,N_18102);
and U23386 (N_23386,N_19107,N_16311);
nor U23387 (N_23387,N_16167,N_19973);
and U23388 (N_23388,N_18213,N_16974);
nand U23389 (N_23389,N_18077,N_19594);
and U23390 (N_23390,N_17616,N_16887);
or U23391 (N_23391,N_17361,N_16082);
or U23392 (N_23392,N_15307,N_16786);
and U23393 (N_23393,N_16917,N_17280);
and U23394 (N_23394,N_15443,N_18586);
nor U23395 (N_23395,N_16739,N_17581);
nor U23396 (N_23396,N_17386,N_19080);
nor U23397 (N_23397,N_18611,N_17394);
nor U23398 (N_23398,N_18591,N_15541);
nor U23399 (N_23399,N_16061,N_17407);
nand U23400 (N_23400,N_19065,N_18006);
and U23401 (N_23401,N_19847,N_15568);
nor U23402 (N_23402,N_17533,N_19024);
nor U23403 (N_23403,N_17963,N_17818);
and U23404 (N_23404,N_18887,N_19685);
nor U23405 (N_23405,N_17875,N_15868);
nand U23406 (N_23406,N_16953,N_16331);
or U23407 (N_23407,N_16908,N_19035);
xnor U23408 (N_23408,N_17625,N_15738);
xor U23409 (N_23409,N_16284,N_15468);
and U23410 (N_23410,N_19009,N_17556);
xnor U23411 (N_23411,N_19897,N_19246);
or U23412 (N_23412,N_19578,N_19909);
xor U23413 (N_23413,N_19094,N_18954);
xnor U23414 (N_23414,N_15154,N_19885);
nand U23415 (N_23415,N_16054,N_15072);
or U23416 (N_23416,N_17506,N_18445);
and U23417 (N_23417,N_15040,N_15705);
xnor U23418 (N_23418,N_17003,N_19245);
nand U23419 (N_23419,N_19375,N_16886);
xnor U23420 (N_23420,N_16596,N_18757);
and U23421 (N_23421,N_16433,N_17847);
xnor U23422 (N_23422,N_15106,N_15489);
nand U23423 (N_23423,N_17039,N_15434);
and U23424 (N_23424,N_17659,N_19027);
xor U23425 (N_23425,N_19335,N_17785);
xnor U23426 (N_23426,N_18736,N_18342);
nor U23427 (N_23427,N_15359,N_18234);
nand U23428 (N_23428,N_17997,N_17744);
and U23429 (N_23429,N_18139,N_17561);
nor U23430 (N_23430,N_17196,N_15254);
or U23431 (N_23431,N_17609,N_18927);
and U23432 (N_23432,N_17303,N_17279);
nor U23433 (N_23433,N_15596,N_17976);
and U23434 (N_23434,N_16045,N_19708);
nor U23435 (N_23435,N_18508,N_18450);
xnor U23436 (N_23436,N_15717,N_15237);
nand U23437 (N_23437,N_19911,N_18513);
xnor U23438 (N_23438,N_19925,N_15581);
xor U23439 (N_23439,N_18036,N_15950);
nor U23440 (N_23440,N_16965,N_19900);
nor U23441 (N_23441,N_18649,N_17151);
and U23442 (N_23442,N_18523,N_19834);
nor U23443 (N_23443,N_19325,N_16780);
or U23444 (N_23444,N_18068,N_17058);
xor U23445 (N_23445,N_19564,N_17949);
or U23446 (N_23446,N_16139,N_15561);
and U23447 (N_23447,N_19067,N_15268);
and U23448 (N_23448,N_15196,N_19003);
nor U23449 (N_23449,N_17832,N_16283);
nor U23450 (N_23450,N_19980,N_19957);
or U23451 (N_23451,N_18809,N_16344);
nand U23452 (N_23452,N_15825,N_18525);
nand U23453 (N_23453,N_15673,N_15865);
or U23454 (N_23454,N_18732,N_17969);
and U23455 (N_23455,N_17564,N_18639);
xor U23456 (N_23456,N_18661,N_15952);
nor U23457 (N_23457,N_18078,N_15287);
and U23458 (N_23458,N_19491,N_19538);
nor U23459 (N_23459,N_15621,N_18630);
or U23460 (N_23460,N_16800,N_15748);
nand U23461 (N_23461,N_17459,N_16911);
and U23462 (N_23462,N_15606,N_18756);
xor U23463 (N_23463,N_15512,N_16837);
nand U23464 (N_23464,N_18168,N_15904);
nor U23465 (N_23465,N_18030,N_18572);
xnor U23466 (N_23466,N_15062,N_16760);
nand U23467 (N_23467,N_18290,N_19965);
nand U23468 (N_23468,N_15099,N_15311);
nor U23469 (N_23469,N_19667,N_18147);
nor U23470 (N_23470,N_17639,N_17093);
and U23471 (N_23471,N_17269,N_17846);
xnor U23472 (N_23472,N_17260,N_19718);
and U23473 (N_23473,N_18148,N_16683);
and U23474 (N_23474,N_16684,N_17035);
nand U23475 (N_23475,N_19064,N_17442);
nand U23476 (N_23476,N_18066,N_16300);
and U23477 (N_23477,N_19854,N_18833);
or U23478 (N_23478,N_16375,N_15830);
xnor U23479 (N_23479,N_19188,N_16671);
or U23480 (N_23480,N_17205,N_16662);
or U23481 (N_23481,N_19505,N_15004);
or U23482 (N_23482,N_17496,N_18839);
nor U23483 (N_23483,N_18460,N_19634);
nor U23484 (N_23484,N_18432,N_15944);
nor U23485 (N_23485,N_19499,N_18217);
nor U23486 (N_23486,N_15926,N_18767);
and U23487 (N_23487,N_18913,N_19697);
xnor U23488 (N_23488,N_17498,N_15817);
nand U23489 (N_23489,N_19315,N_19841);
xor U23490 (N_23490,N_19288,N_18567);
nand U23491 (N_23491,N_17004,N_17836);
and U23492 (N_23492,N_18460,N_16575);
xor U23493 (N_23493,N_19540,N_16601);
nand U23494 (N_23494,N_19981,N_19212);
nor U23495 (N_23495,N_18466,N_17962);
or U23496 (N_23496,N_16332,N_17346);
nand U23497 (N_23497,N_16051,N_19740);
and U23498 (N_23498,N_19748,N_16971);
nor U23499 (N_23499,N_18366,N_16787);
or U23500 (N_23500,N_17059,N_19822);
or U23501 (N_23501,N_19567,N_19830);
nand U23502 (N_23502,N_17963,N_15588);
or U23503 (N_23503,N_17481,N_18067);
nor U23504 (N_23504,N_18249,N_18272);
and U23505 (N_23505,N_19363,N_16757);
nor U23506 (N_23506,N_17132,N_15219);
and U23507 (N_23507,N_19502,N_19942);
nand U23508 (N_23508,N_16654,N_17640);
xor U23509 (N_23509,N_16893,N_19333);
xor U23510 (N_23510,N_15034,N_19687);
or U23511 (N_23511,N_18898,N_15490);
and U23512 (N_23512,N_16272,N_16896);
nor U23513 (N_23513,N_15789,N_15772);
xnor U23514 (N_23514,N_17361,N_18319);
or U23515 (N_23515,N_15944,N_15051);
or U23516 (N_23516,N_15959,N_16014);
nand U23517 (N_23517,N_17952,N_17527);
nor U23518 (N_23518,N_16350,N_15305);
nor U23519 (N_23519,N_18448,N_17366);
and U23520 (N_23520,N_19932,N_17031);
nor U23521 (N_23521,N_18986,N_15934);
nand U23522 (N_23522,N_17294,N_16043);
xnor U23523 (N_23523,N_16186,N_17998);
nand U23524 (N_23524,N_19146,N_16268);
or U23525 (N_23525,N_18895,N_19423);
nor U23526 (N_23526,N_17373,N_18462);
nor U23527 (N_23527,N_15743,N_19921);
and U23528 (N_23528,N_19344,N_18071);
nor U23529 (N_23529,N_18474,N_16550);
nor U23530 (N_23530,N_16983,N_16984);
nand U23531 (N_23531,N_17046,N_17174);
nor U23532 (N_23532,N_16447,N_16727);
or U23533 (N_23533,N_19219,N_19636);
and U23534 (N_23534,N_16011,N_18252);
nand U23535 (N_23535,N_15686,N_19862);
nor U23536 (N_23536,N_19524,N_17347);
nand U23537 (N_23537,N_16577,N_17079);
xor U23538 (N_23538,N_15585,N_16832);
or U23539 (N_23539,N_18019,N_15139);
nor U23540 (N_23540,N_19479,N_18716);
nor U23541 (N_23541,N_19492,N_18614);
nand U23542 (N_23542,N_15987,N_15158);
and U23543 (N_23543,N_15123,N_17951);
or U23544 (N_23544,N_16175,N_18190);
nor U23545 (N_23545,N_19953,N_15405);
and U23546 (N_23546,N_19029,N_16841);
xor U23547 (N_23547,N_18969,N_16473);
and U23548 (N_23548,N_15590,N_19430);
xnor U23549 (N_23549,N_17399,N_17969);
nor U23550 (N_23550,N_16212,N_18584);
or U23551 (N_23551,N_18573,N_18538);
nor U23552 (N_23552,N_15124,N_16593);
xor U23553 (N_23553,N_17026,N_19256);
nor U23554 (N_23554,N_16207,N_19553);
or U23555 (N_23555,N_17818,N_19550);
and U23556 (N_23556,N_17252,N_17553);
and U23557 (N_23557,N_15700,N_18321);
or U23558 (N_23558,N_19019,N_16446);
xor U23559 (N_23559,N_15298,N_17278);
and U23560 (N_23560,N_16420,N_16416);
xnor U23561 (N_23561,N_17628,N_17498);
xor U23562 (N_23562,N_15017,N_15039);
nand U23563 (N_23563,N_18693,N_18437);
or U23564 (N_23564,N_15625,N_18640);
and U23565 (N_23565,N_17726,N_19534);
or U23566 (N_23566,N_19753,N_16033);
and U23567 (N_23567,N_15890,N_17377);
nor U23568 (N_23568,N_17660,N_16016);
nand U23569 (N_23569,N_19415,N_18261);
nor U23570 (N_23570,N_17672,N_15691);
nor U23571 (N_23571,N_16119,N_18925);
nor U23572 (N_23572,N_17438,N_16791);
nand U23573 (N_23573,N_17501,N_18182);
nand U23574 (N_23574,N_16394,N_15098);
and U23575 (N_23575,N_15258,N_19728);
and U23576 (N_23576,N_16101,N_16425);
nand U23577 (N_23577,N_16118,N_15585);
nor U23578 (N_23578,N_18929,N_15032);
nand U23579 (N_23579,N_18574,N_19896);
nand U23580 (N_23580,N_16364,N_19397);
nor U23581 (N_23581,N_17187,N_19004);
nand U23582 (N_23582,N_18122,N_15166);
nand U23583 (N_23583,N_17299,N_17840);
and U23584 (N_23584,N_15807,N_16601);
xor U23585 (N_23585,N_16001,N_19203);
nor U23586 (N_23586,N_18183,N_17013);
nor U23587 (N_23587,N_15532,N_19147);
nand U23588 (N_23588,N_19122,N_18904);
and U23589 (N_23589,N_19950,N_15797);
nor U23590 (N_23590,N_15428,N_16720);
nand U23591 (N_23591,N_16777,N_17840);
and U23592 (N_23592,N_15983,N_15391);
nor U23593 (N_23593,N_15320,N_18958);
or U23594 (N_23594,N_17284,N_19601);
nor U23595 (N_23595,N_16358,N_18857);
xnor U23596 (N_23596,N_18012,N_19347);
nor U23597 (N_23597,N_19030,N_17984);
nor U23598 (N_23598,N_17733,N_17148);
nor U23599 (N_23599,N_18089,N_15135);
xor U23600 (N_23600,N_18427,N_17486);
and U23601 (N_23601,N_18537,N_17832);
xnor U23602 (N_23602,N_15584,N_17671);
nand U23603 (N_23603,N_18327,N_17837);
and U23604 (N_23604,N_16170,N_18682);
nand U23605 (N_23605,N_15068,N_17173);
and U23606 (N_23606,N_18413,N_15349);
xor U23607 (N_23607,N_18491,N_19719);
or U23608 (N_23608,N_17369,N_16767);
nand U23609 (N_23609,N_17393,N_16004);
nand U23610 (N_23610,N_17002,N_17006);
xnor U23611 (N_23611,N_16117,N_18836);
xnor U23612 (N_23612,N_16419,N_18957);
nand U23613 (N_23613,N_16989,N_15470);
or U23614 (N_23614,N_19610,N_15106);
nor U23615 (N_23615,N_19754,N_16495);
and U23616 (N_23616,N_15570,N_18896);
xor U23617 (N_23617,N_17311,N_18120);
xor U23618 (N_23618,N_15761,N_15886);
and U23619 (N_23619,N_18800,N_17232);
nand U23620 (N_23620,N_16694,N_16511);
xnor U23621 (N_23621,N_17492,N_18170);
or U23622 (N_23622,N_19930,N_18401);
or U23623 (N_23623,N_18678,N_18544);
nand U23624 (N_23624,N_17400,N_17924);
nand U23625 (N_23625,N_16861,N_17055);
and U23626 (N_23626,N_18852,N_15830);
or U23627 (N_23627,N_16720,N_17721);
or U23628 (N_23628,N_17273,N_15811);
and U23629 (N_23629,N_16906,N_16993);
nand U23630 (N_23630,N_18668,N_17332);
and U23631 (N_23631,N_16180,N_19692);
or U23632 (N_23632,N_18887,N_15377);
nand U23633 (N_23633,N_19919,N_18577);
nand U23634 (N_23634,N_16134,N_17992);
or U23635 (N_23635,N_19420,N_17733);
and U23636 (N_23636,N_16642,N_18520);
and U23637 (N_23637,N_19505,N_19726);
and U23638 (N_23638,N_18129,N_18131);
and U23639 (N_23639,N_19809,N_16741);
xnor U23640 (N_23640,N_18144,N_19899);
nand U23641 (N_23641,N_16634,N_16971);
xor U23642 (N_23642,N_18641,N_18056);
or U23643 (N_23643,N_19166,N_15678);
nand U23644 (N_23644,N_18097,N_17459);
nand U23645 (N_23645,N_19061,N_19466);
nand U23646 (N_23646,N_18404,N_18717);
or U23647 (N_23647,N_15131,N_15984);
nand U23648 (N_23648,N_17324,N_17687);
xnor U23649 (N_23649,N_15712,N_15435);
nand U23650 (N_23650,N_19605,N_15353);
nor U23651 (N_23651,N_15648,N_19399);
nand U23652 (N_23652,N_15615,N_15202);
or U23653 (N_23653,N_18961,N_18155);
nor U23654 (N_23654,N_19224,N_18748);
nand U23655 (N_23655,N_18684,N_16943);
and U23656 (N_23656,N_19764,N_18019);
and U23657 (N_23657,N_17138,N_15893);
or U23658 (N_23658,N_19770,N_15333);
nand U23659 (N_23659,N_16420,N_15889);
or U23660 (N_23660,N_17227,N_19161);
and U23661 (N_23661,N_15678,N_17961);
and U23662 (N_23662,N_18635,N_16818);
xnor U23663 (N_23663,N_18225,N_18604);
and U23664 (N_23664,N_16099,N_16412);
nor U23665 (N_23665,N_16057,N_16001);
xnor U23666 (N_23666,N_19399,N_18806);
xnor U23667 (N_23667,N_16356,N_15964);
or U23668 (N_23668,N_19259,N_18344);
and U23669 (N_23669,N_17919,N_19185);
nor U23670 (N_23670,N_18259,N_17588);
nand U23671 (N_23671,N_18491,N_16914);
or U23672 (N_23672,N_16428,N_15874);
nor U23673 (N_23673,N_15434,N_16422);
or U23674 (N_23674,N_18694,N_17445);
nand U23675 (N_23675,N_15069,N_15455);
xnor U23676 (N_23676,N_17449,N_16017);
nand U23677 (N_23677,N_19900,N_15732);
nor U23678 (N_23678,N_15733,N_17217);
nor U23679 (N_23679,N_19300,N_18062);
and U23680 (N_23680,N_19473,N_15432);
and U23681 (N_23681,N_19029,N_15704);
xor U23682 (N_23682,N_17459,N_17487);
xnor U23683 (N_23683,N_18800,N_19243);
nor U23684 (N_23684,N_15702,N_15835);
and U23685 (N_23685,N_19950,N_18057);
or U23686 (N_23686,N_19318,N_16494);
or U23687 (N_23687,N_19665,N_17395);
nand U23688 (N_23688,N_17899,N_17081);
nand U23689 (N_23689,N_16979,N_17247);
xnor U23690 (N_23690,N_17776,N_19506);
or U23691 (N_23691,N_19507,N_19830);
and U23692 (N_23692,N_18918,N_17135);
nor U23693 (N_23693,N_19525,N_19342);
or U23694 (N_23694,N_15315,N_16757);
nor U23695 (N_23695,N_19019,N_17724);
nor U23696 (N_23696,N_17228,N_15788);
xor U23697 (N_23697,N_19044,N_15996);
and U23698 (N_23698,N_15483,N_16873);
xnor U23699 (N_23699,N_16956,N_16439);
nor U23700 (N_23700,N_15122,N_18277);
xor U23701 (N_23701,N_17595,N_16925);
nand U23702 (N_23702,N_15407,N_18987);
nor U23703 (N_23703,N_17030,N_16295);
xnor U23704 (N_23704,N_19187,N_15157);
and U23705 (N_23705,N_17067,N_18790);
xor U23706 (N_23706,N_16905,N_15125);
nor U23707 (N_23707,N_17507,N_15061);
nor U23708 (N_23708,N_17704,N_16516);
xor U23709 (N_23709,N_17351,N_16605);
and U23710 (N_23710,N_15315,N_19992);
and U23711 (N_23711,N_18975,N_19094);
nor U23712 (N_23712,N_18268,N_16116);
nand U23713 (N_23713,N_16552,N_18412);
xnor U23714 (N_23714,N_15946,N_15869);
or U23715 (N_23715,N_16525,N_15331);
and U23716 (N_23716,N_19502,N_17940);
and U23717 (N_23717,N_17419,N_19941);
and U23718 (N_23718,N_19118,N_19493);
and U23719 (N_23719,N_18190,N_18551);
nand U23720 (N_23720,N_15456,N_17835);
nand U23721 (N_23721,N_17505,N_19714);
and U23722 (N_23722,N_16444,N_16192);
or U23723 (N_23723,N_15745,N_19151);
xor U23724 (N_23724,N_18041,N_16872);
or U23725 (N_23725,N_18497,N_18293);
xnor U23726 (N_23726,N_18471,N_16713);
nand U23727 (N_23727,N_17019,N_18184);
nand U23728 (N_23728,N_15464,N_16467);
xor U23729 (N_23729,N_19386,N_16152);
nand U23730 (N_23730,N_18528,N_16215);
nand U23731 (N_23731,N_15452,N_16645);
xor U23732 (N_23732,N_17041,N_18105);
nor U23733 (N_23733,N_19286,N_15019);
and U23734 (N_23734,N_19188,N_17834);
and U23735 (N_23735,N_19799,N_15639);
nand U23736 (N_23736,N_15040,N_15689);
and U23737 (N_23737,N_15256,N_17517);
nand U23738 (N_23738,N_19077,N_18183);
or U23739 (N_23739,N_15421,N_17350);
and U23740 (N_23740,N_17068,N_16557);
nand U23741 (N_23741,N_17682,N_19597);
or U23742 (N_23742,N_15712,N_19898);
nand U23743 (N_23743,N_18839,N_18149);
and U23744 (N_23744,N_16791,N_16673);
and U23745 (N_23745,N_17719,N_18771);
xor U23746 (N_23746,N_15894,N_17194);
nor U23747 (N_23747,N_19177,N_18495);
nor U23748 (N_23748,N_17917,N_19797);
nand U23749 (N_23749,N_16210,N_16171);
xnor U23750 (N_23750,N_17887,N_17668);
nor U23751 (N_23751,N_18395,N_18744);
xor U23752 (N_23752,N_16159,N_17254);
nand U23753 (N_23753,N_19214,N_16524);
xnor U23754 (N_23754,N_19445,N_15407);
nor U23755 (N_23755,N_15298,N_16059);
and U23756 (N_23756,N_17117,N_18310);
nand U23757 (N_23757,N_15607,N_18975);
and U23758 (N_23758,N_19948,N_16365);
nand U23759 (N_23759,N_19773,N_15656);
xnor U23760 (N_23760,N_18121,N_18384);
or U23761 (N_23761,N_18665,N_18623);
nor U23762 (N_23762,N_18474,N_15532);
and U23763 (N_23763,N_18653,N_19433);
nor U23764 (N_23764,N_19441,N_19792);
and U23765 (N_23765,N_15369,N_17456);
or U23766 (N_23766,N_17811,N_15387);
nor U23767 (N_23767,N_18251,N_19964);
nand U23768 (N_23768,N_17392,N_19411);
or U23769 (N_23769,N_15313,N_16671);
or U23770 (N_23770,N_17816,N_16832);
and U23771 (N_23771,N_16054,N_16700);
nor U23772 (N_23772,N_17300,N_18851);
nand U23773 (N_23773,N_16461,N_18579);
nand U23774 (N_23774,N_15437,N_16167);
xnor U23775 (N_23775,N_17754,N_19148);
xnor U23776 (N_23776,N_18224,N_15475);
and U23777 (N_23777,N_17238,N_19878);
nand U23778 (N_23778,N_17903,N_16428);
xnor U23779 (N_23779,N_15684,N_19608);
nor U23780 (N_23780,N_18039,N_18313);
or U23781 (N_23781,N_17279,N_19800);
or U23782 (N_23782,N_15813,N_16604);
xor U23783 (N_23783,N_19029,N_16305);
xnor U23784 (N_23784,N_17535,N_18155);
xor U23785 (N_23785,N_19682,N_15968);
nand U23786 (N_23786,N_16030,N_18072);
xnor U23787 (N_23787,N_19297,N_19280);
or U23788 (N_23788,N_16086,N_16323);
nor U23789 (N_23789,N_17315,N_18293);
or U23790 (N_23790,N_18090,N_19619);
nor U23791 (N_23791,N_19968,N_19034);
nor U23792 (N_23792,N_15945,N_16263);
nand U23793 (N_23793,N_18476,N_17685);
nand U23794 (N_23794,N_16037,N_17534);
nor U23795 (N_23795,N_16414,N_17374);
nor U23796 (N_23796,N_17274,N_18186);
nor U23797 (N_23797,N_15343,N_16113);
nand U23798 (N_23798,N_16419,N_17634);
or U23799 (N_23799,N_17205,N_15651);
nand U23800 (N_23800,N_17457,N_15502);
nand U23801 (N_23801,N_19635,N_15549);
or U23802 (N_23802,N_18847,N_19707);
nor U23803 (N_23803,N_15651,N_17593);
xnor U23804 (N_23804,N_16192,N_19060);
and U23805 (N_23805,N_16241,N_15799);
or U23806 (N_23806,N_19364,N_15209);
and U23807 (N_23807,N_18939,N_17242);
and U23808 (N_23808,N_17316,N_15706);
and U23809 (N_23809,N_16313,N_17813);
nand U23810 (N_23810,N_17375,N_18099);
nand U23811 (N_23811,N_16404,N_17070);
xor U23812 (N_23812,N_15844,N_18539);
and U23813 (N_23813,N_19355,N_16696);
nand U23814 (N_23814,N_19188,N_17728);
xor U23815 (N_23815,N_15308,N_17777);
or U23816 (N_23816,N_17079,N_18413);
xor U23817 (N_23817,N_17511,N_15946);
and U23818 (N_23818,N_15328,N_16744);
and U23819 (N_23819,N_16452,N_15855);
nor U23820 (N_23820,N_16704,N_17631);
and U23821 (N_23821,N_19545,N_18082);
nand U23822 (N_23822,N_19394,N_15424);
and U23823 (N_23823,N_19411,N_17876);
nor U23824 (N_23824,N_17177,N_19893);
nor U23825 (N_23825,N_15811,N_17022);
nand U23826 (N_23826,N_15487,N_16242);
or U23827 (N_23827,N_15432,N_18988);
xnor U23828 (N_23828,N_19359,N_16917);
nor U23829 (N_23829,N_19714,N_17179);
nor U23830 (N_23830,N_17015,N_19664);
or U23831 (N_23831,N_17209,N_17955);
or U23832 (N_23832,N_16525,N_16792);
and U23833 (N_23833,N_19433,N_17375);
or U23834 (N_23834,N_16986,N_18667);
nor U23835 (N_23835,N_15926,N_19758);
or U23836 (N_23836,N_15837,N_19080);
nand U23837 (N_23837,N_18949,N_16529);
and U23838 (N_23838,N_18496,N_18606);
nand U23839 (N_23839,N_19692,N_17655);
and U23840 (N_23840,N_17106,N_17436);
xor U23841 (N_23841,N_18897,N_17020);
nand U23842 (N_23842,N_18025,N_17935);
xnor U23843 (N_23843,N_16646,N_15986);
nand U23844 (N_23844,N_15597,N_15975);
xnor U23845 (N_23845,N_16787,N_18431);
or U23846 (N_23846,N_17140,N_18473);
and U23847 (N_23847,N_18611,N_19485);
or U23848 (N_23848,N_18564,N_18919);
nor U23849 (N_23849,N_15725,N_19995);
nand U23850 (N_23850,N_18998,N_16876);
and U23851 (N_23851,N_15349,N_16464);
nand U23852 (N_23852,N_16297,N_17045);
and U23853 (N_23853,N_18115,N_16028);
nor U23854 (N_23854,N_18987,N_19298);
xor U23855 (N_23855,N_16701,N_15837);
nand U23856 (N_23856,N_18952,N_15132);
nand U23857 (N_23857,N_15999,N_19249);
nor U23858 (N_23858,N_15367,N_18334);
nor U23859 (N_23859,N_17060,N_17258);
and U23860 (N_23860,N_19212,N_18556);
xnor U23861 (N_23861,N_17420,N_16248);
nand U23862 (N_23862,N_18800,N_17279);
xor U23863 (N_23863,N_15419,N_19673);
nor U23864 (N_23864,N_19918,N_16863);
or U23865 (N_23865,N_17011,N_19445);
or U23866 (N_23866,N_19357,N_16912);
nor U23867 (N_23867,N_19872,N_16216);
nor U23868 (N_23868,N_16924,N_19960);
and U23869 (N_23869,N_15684,N_15915);
and U23870 (N_23870,N_17925,N_15647);
nor U23871 (N_23871,N_18767,N_15134);
or U23872 (N_23872,N_15684,N_17101);
xnor U23873 (N_23873,N_19823,N_18649);
nand U23874 (N_23874,N_16822,N_18903);
nor U23875 (N_23875,N_15909,N_19773);
nand U23876 (N_23876,N_18777,N_18848);
nor U23877 (N_23877,N_16562,N_15326);
nor U23878 (N_23878,N_17543,N_19298);
nand U23879 (N_23879,N_18001,N_15112);
nor U23880 (N_23880,N_15905,N_17995);
nor U23881 (N_23881,N_15163,N_19387);
nor U23882 (N_23882,N_17886,N_16962);
xor U23883 (N_23883,N_18328,N_19145);
nand U23884 (N_23884,N_16518,N_15600);
or U23885 (N_23885,N_16281,N_19373);
and U23886 (N_23886,N_19813,N_15287);
or U23887 (N_23887,N_15613,N_19250);
nand U23888 (N_23888,N_17681,N_16065);
and U23889 (N_23889,N_17108,N_19871);
xnor U23890 (N_23890,N_17575,N_19625);
nand U23891 (N_23891,N_18409,N_17881);
and U23892 (N_23892,N_17162,N_17187);
nand U23893 (N_23893,N_17578,N_19948);
and U23894 (N_23894,N_17066,N_17092);
nand U23895 (N_23895,N_15541,N_16040);
xnor U23896 (N_23896,N_16900,N_19162);
nand U23897 (N_23897,N_15225,N_17024);
nand U23898 (N_23898,N_18453,N_18070);
xor U23899 (N_23899,N_16921,N_19709);
xnor U23900 (N_23900,N_16875,N_15872);
xor U23901 (N_23901,N_19582,N_16289);
xor U23902 (N_23902,N_15231,N_17059);
or U23903 (N_23903,N_16889,N_17723);
nor U23904 (N_23904,N_18970,N_15453);
or U23905 (N_23905,N_19237,N_19900);
nor U23906 (N_23906,N_16711,N_16659);
nor U23907 (N_23907,N_17902,N_18176);
xnor U23908 (N_23908,N_19225,N_15346);
or U23909 (N_23909,N_19608,N_15596);
nand U23910 (N_23910,N_15455,N_16150);
and U23911 (N_23911,N_18124,N_17827);
nor U23912 (N_23912,N_17594,N_17266);
nand U23913 (N_23913,N_18050,N_19003);
xor U23914 (N_23914,N_18293,N_18076);
nor U23915 (N_23915,N_19173,N_19535);
nand U23916 (N_23916,N_17478,N_15001);
and U23917 (N_23917,N_16877,N_16434);
nor U23918 (N_23918,N_18044,N_15937);
and U23919 (N_23919,N_15568,N_19671);
and U23920 (N_23920,N_17640,N_19777);
nor U23921 (N_23921,N_17099,N_17672);
and U23922 (N_23922,N_17907,N_16738);
nand U23923 (N_23923,N_16638,N_16661);
or U23924 (N_23924,N_17277,N_15658);
or U23925 (N_23925,N_15942,N_17356);
or U23926 (N_23926,N_17297,N_17840);
or U23927 (N_23927,N_17425,N_18286);
nor U23928 (N_23928,N_18556,N_16712);
nand U23929 (N_23929,N_17612,N_18919);
or U23930 (N_23930,N_17510,N_17573);
xnor U23931 (N_23931,N_17763,N_18675);
and U23932 (N_23932,N_17368,N_15999);
nor U23933 (N_23933,N_15069,N_17332);
or U23934 (N_23934,N_16801,N_17538);
xnor U23935 (N_23935,N_16334,N_17146);
xor U23936 (N_23936,N_19703,N_16794);
or U23937 (N_23937,N_16524,N_18140);
and U23938 (N_23938,N_15061,N_17485);
xor U23939 (N_23939,N_17751,N_18878);
nor U23940 (N_23940,N_16859,N_16414);
nor U23941 (N_23941,N_18576,N_16703);
nor U23942 (N_23942,N_19110,N_17359);
xnor U23943 (N_23943,N_15453,N_18931);
or U23944 (N_23944,N_15984,N_16374);
and U23945 (N_23945,N_18699,N_16856);
and U23946 (N_23946,N_18977,N_15639);
or U23947 (N_23947,N_18846,N_18565);
and U23948 (N_23948,N_18470,N_17895);
or U23949 (N_23949,N_15936,N_18139);
and U23950 (N_23950,N_17015,N_17855);
or U23951 (N_23951,N_18396,N_18701);
xor U23952 (N_23952,N_19650,N_19022);
xor U23953 (N_23953,N_19158,N_19168);
and U23954 (N_23954,N_17083,N_17769);
nor U23955 (N_23955,N_16394,N_17922);
nor U23956 (N_23956,N_15564,N_17329);
xnor U23957 (N_23957,N_16034,N_17025);
and U23958 (N_23958,N_18283,N_19184);
nor U23959 (N_23959,N_19270,N_17984);
and U23960 (N_23960,N_15606,N_19364);
nor U23961 (N_23961,N_17401,N_18755);
or U23962 (N_23962,N_19869,N_19432);
nor U23963 (N_23963,N_17381,N_17130);
nor U23964 (N_23964,N_15791,N_18855);
nand U23965 (N_23965,N_19322,N_19787);
and U23966 (N_23966,N_16896,N_16265);
or U23967 (N_23967,N_16555,N_19371);
or U23968 (N_23968,N_17970,N_19604);
xnor U23969 (N_23969,N_15362,N_19400);
nor U23970 (N_23970,N_19547,N_17380);
nand U23971 (N_23971,N_16718,N_16564);
nor U23972 (N_23972,N_15500,N_15659);
xnor U23973 (N_23973,N_19187,N_15808);
or U23974 (N_23974,N_17013,N_17721);
nand U23975 (N_23975,N_18051,N_15568);
nor U23976 (N_23976,N_16431,N_17120);
nand U23977 (N_23977,N_19616,N_18229);
or U23978 (N_23978,N_17452,N_19220);
xor U23979 (N_23979,N_15325,N_19790);
nor U23980 (N_23980,N_19762,N_17423);
and U23981 (N_23981,N_17506,N_17752);
xor U23982 (N_23982,N_18880,N_19393);
and U23983 (N_23983,N_15984,N_18417);
or U23984 (N_23984,N_16113,N_16124);
nor U23985 (N_23985,N_19226,N_18271);
nand U23986 (N_23986,N_17968,N_17175);
or U23987 (N_23987,N_18305,N_16328);
and U23988 (N_23988,N_16714,N_16814);
nor U23989 (N_23989,N_17720,N_16886);
and U23990 (N_23990,N_16684,N_15633);
nand U23991 (N_23991,N_15711,N_19407);
nand U23992 (N_23992,N_19357,N_15587);
xor U23993 (N_23993,N_17127,N_16516);
or U23994 (N_23994,N_19386,N_19605);
nand U23995 (N_23995,N_18897,N_16147);
xor U23996 (N_23996,N_19318,N_15642);
nand U23997 (N_23997,N_18317,N_15342);
xor U23998 (N_23998,N_19671,N_16809);
or U23999 (N_23999,N_19634,N_17231);
xor U24000 (N_24000,N_16428,N_16759);
nand U24001 (N_24001,N_15461,N_17498);
xnor U24002 (N_24002,N_17201,N_16583);
or U24003 (N_24003,N_16904,N_18351);
xor U24004 (N_24004,N_15687,N_18006);
xor U24005 (N_24005,N_15814,N_17788);
or U24006 (N_24006,N_15695,N_16333);
xnor U24007 (N_24007,N_17810,N_16144);
nor U24008 (N_24008,N_15902,N_17295);
nor U24009 (N_24009,N_19551,N_15110);
nand U24010 (N_24010,N_19776,N_19052);
and U24011 (N_24011,N_16791,N_16490);
and U24012 (N_24012,N_18060,N_15414);
and U24013 (N_24013,N_15729,N_17464);
or U24014 (N_24014,N_17288,N_16649);
and U24015 (N_24015,N_19020,N_17234);
xnor U24016 (N_24016,N_16702,N_19085);
and U24017 (N_24017,N_18539,N_18649);
xor U24018 (N_24018,N_17316,N_16107);
xnor U24019 (N_24019,N_18593,N_15951);
xor U24020 (N_24020,N_19858,N_15480);
nor U24021 (N_24021,N_16401,N_16115);
and U24022 (N_24022,N_19362,N_15262);
nor U24023 (N_24023,N_19216,N_18194);
nand U24024 (N_24024,N_16674,N_17527);
nor U24025 (N_24025,N_17189,N_16561);
and U24026 (N_24026,N_15324,N_19533);
or U24027 (N_24027,N_17171,N_15414);
xor U24028 (N_24028,N_15338,N_15236);
xor U24029 (N_24029,N_15443,N_18296);
or U24030 (N_24030,N_16893,N_19121);
nand U24031 (N_24031,N_18466,N_18333);
nor U24032 (N_24032,N_17647,N_19852);
nand U24033 (N_24033,N_17408,N_15521);
nand U24034 (N_24034,N_15635,N_16975);
nor U24035 (N_24035,N_17470,N_16151);
and U24036 (N_24036,N_16778,N_15814);
and U24037 (N_24037,N_17585,N_19475);
nand U24038 (N_24038,N_19368,N_17294);
or U24039 (N_24039,N_19984,N_19469);
nor U24040 (N_24040,N_19591,N_19728);
xnor U24041 (N_24041,N_19487,N_17667);
nor U24042 (N_24042,N_19011,N_19914);
nor U24043 (N_24043,N_16153,N_18544);
nand U24044 (N_24044,N_17927,N_18196);
xnor U24045 (N_24045,N_17869,N_15129);
and U24046 (N_24046,N_19339,N_19448);
and U24047 (N_24047,N_16149,N_18314);
nor U24048 (N_24048,N_15888,N_18561);
or U24049 (N_24049,N_16298,N_18701);
nor U24050 (N_24050,N_19538,N_18711);
or U24051 (N_24051,N_18941,N_18441);
nor U24052 (N_24052,N_17695,N_15187);
and U24053 (N_24053,N_15346,N_17183);
xnor U24054 (N_24054,N_16067,N_19533);
nor U24055 (N_24055,N_16040,N_15271);
nor U24056 (N_24056,N_18302,N_18321);
and U24057 (N_24057,N_15075,N_17749);
xor U24058 (N_24058,N_18699,N_15901);
nor U24059 (N_24059,N_17118,N_19573);
xnor U24060 (N_24060,N_18021,N_19326);
nand U24061 (N_24061,N_17959,N_16783);
xnor U24062 (N_24062,N_18979,N_16436);
nand U24063 (N_24063,N_17190,N_17670);
nand U24064 (N_24064,N_17406,N_19844);
and U24065 (N_24065,N_19564,N_19272);
and U24066 (N_24066,N_16316,N_16970);
xnor U24067 (N_24067,N_15953,N_18516);
nor U24068 (N_24068,N_18524,N_19211);
nor U24069 (N_24069,N_19243,N_18036);
xor U24070 (N_24070,N_18223,N_15666);
nor U24071 (N_24071,N_19884,N_18844);
xnor U24072 (N_24072,N_15735,N_17320);
nor U24073 (N_24073,N_19328,N_15110);
nand U24074 (N_24074,N_17987,N_16669);
nor U24075 (N_24075,N_17331,N_15742);
xnor U24076 (N_24076,N_16289,N_17310);
or U24077 (N_24077,N_15537,N_18347);
nand U24078 (N_24078,N_19591,N_17334);
nand U24079 (N_24079,N_18158,N_15294);
and U24080 (N_24080,N_17953,N_19610);
xor U24081 (N_24081,N_19824,N_19904);
xnor U24082 (N_24082,N_16295,N_18708);
nor U24083 (N_24083,N_17645,N_16083);
or U24084 (N_24084,N_15677,N_17488);
nand U24085 (N_24085,N_15374,N_16321);
nand U24086 (N_24086,N_15731,N_19197);
xnor U24087 (N_24087,N_16693,N_15452);
or U24088 (N_24088,N_19262,N_19673);
nand U24089 (N_24089,N_15006,N_19462);
or U24090 (N_24090,N_15434,N_16096);
xnor U24091 (N_24091,N_18469,N_17011);
xnor U24092 (N_24092,N_18921,N_18914);
xnor U24093 (N_24093,N_17405,N_18940);
or U24094 (N_24094,N_19039,N_19968);
nor U24095 (N_24095,N_15535,N_18237);
xor U24096 (N_24096,N_18442,N_15956);
and U24097 (N_24097,N_15853,N_19865);
nand U24098 (N_24098,N_18417,N_15227);
or U24099 (N_24099,N_19801,N_15003);
and U24100 (N_24100,N_15879,N_19755);
nor U24101 (N_24101,N_16096,N_17837);
and U24102 (N_24102,N_17097,N_16004);
nor U24103 (N_24103,N_17139,N_19399);
nand U24104 (N_24104,N_17251,N_16331);
and U24105 (N_24105,N_17316,N_16615);
and U24106 (N_24106,N_17106,N_17993);
xnor U24107 (N_24107,N_15649,N_19354);
nor U24108 (N_24108,N_16813,N_17243);
xnor U24109 (N_24109,N_15708,N_19121);
xnor U24110 (N_24110,N_15042,N_17335);
xnor U24111 (N_24111,N_18446,N_16440);
or U24112 (N_24112,N_18033,N_19059);
nand U24113 (N_24113,N_17693,N_18558);
or U24114 (N_24114,N_15252,N_19498);
and U24115 (N_24115,N_19478,N_19891);
nand U24116 (N_24116,N_19297,N_19566);
nand U24117 (N_24117,N_16405,N_15855);
nand U24118 (N_24118,N_15362,N_16040);
nand U24119 (N_24119,N_18079,N_15166);
nand U24120 (N_24120,N_18219,N_18191);
nor U24121 (N_24121,N_17130,N_18645);
xor U24122 (N_24122,N_18469,N_18280);
nor U24123 (N_24123,N_17013,N_17350);
nor U24124 (N_24124,N_18342,N_19390);
or U24125 (N_24125,N_19484,N_16935);
or U24126 (N_24126,N_19442,N_15191);
nand U24127 (N_24127,N_16538,N_17621);
or U24128 (N_24128,N_18223,N_16242);
or U24129 (N_24129,N_19920,N_16280);
xor U24130 (N_24130,N_15017,N_18325);
or U24131 (N_24131,N_16359,N_18357);
nor U24132 (N_24132,N_16442,N_18388);
nor U24133 (N_24133,N_19101,N_17500);
nand U24134 (N_24134,N_16550,N_17560);
xnor U24135 (N_24135,N_19632,N_16634);
or U24136 (N_24136,N_18563,N_18887);
and U24137 (N_24137,N_16514,N_18605);
nand U24138 (N_24138,N_17417,N_18142);
nor U24139 (N_24139,N_19090,N_16399);
nand U24140 (N_24140,N_16626,N_18270);
nand U24141 (N_24141,N_18899,N_18760);
and U24142 (N_24142,N_17055,N_16239);
xnor U24143 (N_24143,N_19060,N_19264);
and U24144 (N_24144,N_18717,N_15800);
nor U24145 (N_24145,N_16466,N_16606);
xor U24146 (N_24146,N_16063,N_16633);
nor U24147 (N_24147,N_18827,N_15639);
nor U24148 (N_24148,N_19877,N_19929);
nand U24149 (N_24149,N_15968,N_17865);
and U24150 (N_24150,N_18868,N_17274);
and U24151 (N_24151,N_19591,N_19640);
and U24152 (N_24152,N_15713,N_16561);
or U24153 (N_24153,N_19470,N_16363);
nand U24154 (N_24154,N_16940,N_19337);
and U24155 (N_24155,N_17132,N_19831);
nand U24156 (N_24156,N_17274,N_16535);
nor U24157 (N_24157,N_19230,N_18383);
nand U24158 (N_24158,N_18907,N_15189);
nand U24159 (N_24159,N_18579,N_18631);
and U24160 (N_24160,N_18330,N_19157);
nand U24161 (N_24161,N_16320,N_15621);
or U24162 (N_24162,N_17381,N_16519);
xnor U24163 (N_24163,N_19659,N_15260);
xor U24164 (N_24164,N_16493,N_15874);
and U24165 (N_24165,N_17733,N_15508);
nor U24166 (N_24166,N_17092,N_16580);
nor U24167 (N_24167,N_17575,N_19618);
xnor U24168 (N_24168,N_16295,N_19556);
nand U24169 (N_24169,N_17879,N_19627);
nor U24170 (N_24170,N_16818,N_18452);
or U24171 (N_24171,N_17505,N_15830);
xnor U24172 (N_24172,N_18417,N_18825);
xnor U24173 (N_24173,N_18872,N_18373);
nand U24174 (N_24174,N_18673,N_17258);
xor U24175 (N_24175,N_18977,N_16396);
nor U24176 (N_24176,N_16453,N_18325);
xnor U24177 (N_24177,N_18748,N_19505);
xnor U24178 (N_24178,N_19407,N_16468);
nor U24179 (N_24179,N_18181,N_15190);
nor U24180 (N_24180,N_15710,N_16183);
nand U24181 (N_24181,N_19619,N_18623);
nand U24182 (N_24182,N_18849,N_18143);
nor U24183 (N_24183,N_15662,N_16620);
and U24184 (N_24184,N_15990,N_19002);
and U24185 (N_24185,N_18072,N_17917);
and U24186 (N_24186,N_17276,N_19905);
xor U24187 (N_24187,N_15761,N_15695);
xnor U24188 (N_24188,N_15931,N_16521);
nand U24189 (N_24189,N_17907,N_18395);
xnor U24190 (N_24190,N_18102,N_18940);
nor U24191 (N_24191,N_17732,N_17671);
nor U24192 (N_24192,N_15223,N_17899);
and U24193 (N_24193,N_18977,N_17728);
xor U24194 (N_24194,N_16834,N_17678);
xor U24195 (N_24195,N_15224,N_19649);
xor U24196 (N_24196,N_17509,N_19925);
xnor U24197 (N_24197,N_18638,N_19352);
nor U24198 (N_24198,N_18468,N_17285);
and U24199 (N_24199,N_16565,N_19348);
and U24200 (N_24200,N_19528,N_16439);
nand U24201 (N_24201,N_19011,N_18361);
and U24202 (N_24202,N_19069,N_17857);
or U24203 (N_24203,N_18994,N_17175);
and U24204 (N_24204,N_18668,N_15297);
xnor U24205 (N_24205,N_18119,N_19639);
or U24206 (N_24206,N_19272,N_16238);
nand U24207 (N_24207,N_17461,N_19798);
or U24208 (N_24208,N_18952,N_17001);
nor U24209 (N_24209,N_17061,N_15626);
nand U24210 (N_24210,N_15990,N_19029);
and U24211 (N_24211,N_16845,N_17478);
and U24212 (N_24212,N_18368,N_18481);
nand U24213 (N_24213,N_18979,N_17020);
xor U24214 (N_24214,N_17658,N_18211);
and U24215 (N_24215,N_19200,N_19230);
or U24216 (N_24216,N_18742,N_15737);
xor U24217 (N_24217,N_17215,N_17942);
nand U24218 (N_24218,N_18869,N_15727);
and U24219 (N_24219,N_17450,N_15459);
nand U24220 (N_24220,N_16539,N_18524);
nand U24221 (N_24221,N_18772,N_18889);
and U24222 (N_24222,N_19199,N_18894);
xnor U24223 (N_24223,N_15073,N_19690);
nor U24224 (N_24224,N_15509,N_16528);
or U24225 (N_24225,N_18747,N_19901);
nor U24226 (N_24226,N_19286,N_18049);
and U24227 (N_24227,N_15437,N_16559);
xor U24228 (N_24228,N_17877,N_16840);
and U24229 (N_24229,N_15052,N_19675);
xnor U24230 (N_24230,N_17000,N_18943);
or U24231 (N_24231,N_18493,N_19425);
xor U24232 (N_24232,N_18027,N_15738);
nor U24233 (N_24233,N_15196,N_15011);
nor U24234 (N_24234,N_16982,N_18497);
and U24235 (N_24235,N_19620,N_17264);
nor U24236 (N_24236,N_16781,N_19439);
xor U24237 (N_24237,N_16952,N_18416);
nor U24238 (N_24238,N_18582,N_17578);
xnor U24239 (N_24239,N_15230,N_16028);
xnor U24240 (N_24240,N_17331,N_18688);
xor U24241 (N_24241,N_17727,N_16374);
nand U24242 (N_24242,N_17915,N_15196);
or U24243 (N_24243,N_16732,N_19711);
nor U24244 (N_24244,N_18636,N_17107);
nand U24245 (N_24245,N_15919,N_15294);
xnor U24246 (N_24246,N_16331,N_18219);
and U24247 (N_24247,N_19678,N_15505);
or U24248 (N_24248,N_17051,N_19247);
or U24249 (N_24249,N_19012,N_19561);
nand U24250 (N_24250,N_17417,N_19113);
or U24251 (N_24251,N_16857,N_17953);
or U24252 (N_24252,N_19496,N_16543);
and U24253 (N_24253,N_19834,N_16645);
nor U24254 (N_24254,N_18904,N_19007);
or U24255 (N_24255,N_17244,N_19316);
and U24256 (N_24256,N_17978,N_16990);
or U24257 (N_24257,N_16154,N_16730);
nand U24258 (N_24258,N_16015,N_19746);
or U24259 (N_24259,N_19758,N_18070);
or U24260 (N_24260,N_17531,N_19672);
nand U24261 (N_24261,N_18762,N_18165);
nor U24262 (N_24262,N_18712,N_18595);
and U24263 (N_24263,N_16117,N_18153);
xor U24264 (N_24264,N_15233,N_16807);
or U24265 (N_24265,N_16856,N_16191);
nor U24266 (N_24266,N_15965,N_17411);
nor U24267 (N_24267,N_16479,N_15859);
and U24268 (N_24268,N_19154,N_18382);
xor U24269 (N_24269,N_16806,N_15003);
and U24270 (N_24270,N_15421,N_18918);
nand U24271 (N_24271,N_18773,N_18519);
nor U24272 (N_24272,N_19633,N_16434);
nand U24273 (N_24273,N_15737,N_18596);
nand U24274 (N_24274,N_15312,N_16419);
nor U24275 (N_24275,N_18793,N_16281);
nor U24276 (N_24276,N_19967,N_15983);
and U24277 (N_24277,N_17398,N_15628);
and U24278 (N_24278,N_15276,N_18467);
nor U24279 (N_24279,N_16451,N_15218);
nand U24280 (N_24280,N_18180,N_16771);
xnor U24281 (N_24281,N_16876,N_15942);
nor U24282 (N_24282,N_16641,N_16886);
and U24283 (N_24283,N_16491,N_18772);
and U24284 (N_24284,N_17180,N_18919);
nor U24285 (N_24285,N_16624,N_18081);
and U24286 (N_24286,N_19558,N_18734);
xnor U24287 (N_24287,N_15246,N_18816);
and U24288 (N_24288,N_17931,N_19841);
and U24289 (N_24289,N_16390,N_18317);
and U24290 (N_24290,N_16163,N_16221);
or U24291 (N_24291,N_18056,N_19546);
nand U24292 (N_24292,N_18040,N_17285);
nor U24293 (N_24293,N_18668,N_17459);
nor U24294 (N_24294,N_16118,N_18770);
and U24295 (N_24295,N_18803,N_18829);
or U24296 (N_24296,N_19315,N_18816);
xnor U24297 (N_24297,N_16757,N_16738);
nor U24298 (N_24298,N_16830,N_16150);
xnor U24299 (N_24299,N_18112,N_16527);
nand U24300 (N_24300,N_16184,N_16455);
nand U24301 (N_24301,N_17778,N_17567);
nand U24302 (N_24302,N_16781,N_17788);
xor U24303 (N_24303,N_17739,N_19194);
or U24304 (N_24304,N_16370,N_17142);
xor U24305 (N_24305,N_15588,N_19181);
xnor U24306 (N_24306,N_17317,N_19117);
nand U24307 (N_24307,N_19894,N_17009);
and U24308 (N_24308,N_16680,N_19052);
nand U24309 (N_24309,N_15764,N_18925);
nor U24310 (N_24310,N_15314,N_19260);
or U24311 (N_24311,N_16071,N_16846);
and U24312 (N_24312,N_17886,N_17889);
nand U24313 (N_24313,N_16709,N_16679);
or U24314 (N_24314,N_17743,N_19380);
nand U24315 (N_24315,N_16395,N_18670);
and U24316 (N_24316,N_16198,N_19017);
or U24317 (N_24317,N_17385,N_16778);
or U24318 (N_24318,N_19877,N_16471);
xor U24319 (N_24319,N_15729,N_16783);
nand U24320 (N_24320,N_16661,N_15747);
or U24321 (N_24321,N_18996,N_17546);
or U24322 (N_24322,N_19340,N_18960);
nand U24323 (N_24323,N_17282,N_19164);
nand U24324 (N_24324,N_15008,N_16614);
nand U24325 (N_24325,N_17065,N_16273);
nor U24326 (N_24326,N_19717,N_16674);
and U24327 (N_24327,N_17254,N_17755);
or U24328 (N_24328,N_16689,N_16615);
nand U24329 (N_24329,N_15343,N_18689);
nor U24330 (N_24330,N_17505,N_17029);
and U24331 (N_24331,N_18027,N_17800);
and U24332 (N_24332,N_19135,N_16645);
nand U24333 (N_24333,N_16310,N_19050);
xor U24334 (N_24334,N_16606,N_15814);
or U24335 (N_24335,N_16431,N_15030);
nand U24336 (N_24336,N_16149,N_17808);
xnor U24337 (N_24337,N_19790,N_18862);
and U24338 (N_24338,N_18387,N_17710);
or U24339 (N_24339,N_15400,N_16059);
nor U24340 (N_24340,N_16632,N_17409);
nand U24341 (N_24341,N_19816,N_15115);
nor U24342 (N_24342,N_15802,N_15552);
and U24343 (N_24343,N_19367,N_15513);
or U24344 (N_24344,N_15600,N_19597);
nand U24345 (N_24345,N_17587,N_19719);
xnor U24346 (N_24346,N_18456,N_15112);
nor U24347 (N_24347,N_19997,N_19643);
nand U24348 (N_24348,N_16546,N_17946);
or U24349 (N_24349,N_19500,N_16252);
nor U24350 (N_24350,N_19103,N_15580);
or U24351 (N_24351,N_16496,N_19878);
and U24352 (N_24352,N_16915,N_16560);
nor U24353 (N_24353,N_16340,N_16036);
nor U24354 (N_24354,N_17036,N_15827);
nor U24355 (N_24355,N_19973,N_19984);
nor U24356 (N_24356,N_18745,N_18813);
xnor U24357 (N_24357,N_19694,N_16259);
or U24358 (N_24358,N_19366,N_15414);
or U24359 (N_24359,N_17338,N_18086);
nand U24360 (N_24360,N_19975,N_16596);
nor U24361 (N_24361,N_17629,N_17017);
xor U24362 (N_24362,N_19186,N_17327);
nand U24363 (N_24363,N_17202,N_18553);
nor U24364 (N_24364,N_15724,N_19087);
or U24365 (N_24365,N_19987,N_16042);
nor U24366 (N_24366,N_19676,N_15922);
nor U24367 (N_24367,N_18577,N_15343);
nand U24368 (N_24368,N_16666,N_19310);
or U24369 (N_24369,N_17770,N_18301);
or U24370 (N_24370,N_17611,N_15417);
and U24371 (N_24371,N_16546,N_18862);
and U24372 (N_24372,N_17494,N_17222);
xnor U24373 (N_24373,N_19361,N_18692);
or U24374 (N_24374,N_15346,N_15894);
nand U24375 (N_24375,N_19660,N_17100);
nor U24376 (N_24376,N_16603,N_17003);
or U24377 (N_24377,N_17601,N_15715);
or U24378 (N_24378,N_16879,N_16849);
and U24379 (N_24379,N_16280,N_17173);
xnor U24380 (N_24380,N_15163,N_16653);
xnor U24381 (N_24381,N_19093,N_16811);
nor U24382 (N_24382,N_17180,N_16167);
nor U24383 (N_24383,N_18447,N_18160);
xnor U24384 (N_24384,N_17710,N_18440);
nor U24385 (N_24385,N_16405,N_19035);
xnor U24386 (N_24386,N_16413,N_16822);
nor U24387 (N_24387,N_16395,N_18816);
and U24388 (N_24388,N_15446,N_15033);
xor U24389 (N_24389,N_19131,N_17891);
nor U24390 (N_24390,N_15594,N_15868);
and U24391 (N_24391,N_15224,N_18995);
nor U24392 (N_24392,N_19718,N_17652);
nor U24393 (N_24393,N_19273,N_19930);
or U24394 (N_24394,N_17791,N_17005);
nand U24395 (N_24395,N_19935,N_16795);
nor U24396 (N_24396,N_15991,N_18511);
and U24397 (N_24397,N_19533,N_19212);
xnor U24398 (N_24398,N_15601,N_16722);
nand U24399 (N_24399,N_18527,N_17333);
xor U24400 (N_24400,N_16780,N_15826);
and U24401 (N_24401,N_19358,N_17429);
and U24402 (N_24402,N_17266,N_17280);
nand U24403 (N_24403,N_15158,N_16000);
nand U24404 (N_24404,N_19080,N_19344);
xnor U24405 (N_24405,N_17555,N_19967);
and U24406 (N_24406,N_17526,N_15133);
or U24407 (N_24407,N_19613,N_17687);
nor U24408 (N_24408,N_19925,N_19253);
nand U24409 (N_24409,N_18115,N_15645);
or U24410 (N_24410,N_19640,N_18505);
xor U24411 (N_24411,N_17076,N_17314);
and U24412 (N_24412,N_15199,N_16216);
or U24413 (N_24413,N_18962,N_19575);
or U24414 (N_24414,N_16871,N_16513);
and U24415 (N_24415,N_16107,N_15220);
nor U24416 (N_24416,N_16167,N_19085);
nor U24417 (N_24417,N_16062,N_15425);
nor U24418 (N_24418,N_15814,N_16079);
nor U24419 (N_24419,N_19310,N_17010);
nand U24420 (N_24420,N_18735,N_17267);
xor U24421 (N_24421,N_15769,N_19610);
nor U24422 (N_24422,N_18484,N_18224);
and U24423 (N_24423,N_17923,N_18653);
xnor U24424 (N_24424,N_15086,N_16054);
or U24425 (N_24425,N_17954,N_17772);
nand U24426 (N_24426,N_19646,N_16121);
and U24427 (N_24427,N_17147,N_17166);
and U24428 (N_24428,N_15833,N_17299);
xnor U24429 (N_24429,N_17338,N_17765);
and U24430 (N_24430,N_17684,N_17599);
nand U24431 (N_24431,N_15781,N_17447);
xor U24432 (N_24432,N_18650,N_15575);
nor U24433 (N_24433,N_18164,N_17648);
nor U24434 (N_24434,N_16167,N_18913);
or U24435 (N_24435,N_15033,N_18664);
nand U24436 (N_24436,N_19116,N_15764);
nor U24437 (N_24437,N_19485,N_15227);
nor U24438 (N_24438,N_19579,N_19283);
nor U24439 (N_24439,N_15069,N_16094);
or U24440 (N_24440,N_18253,N_18349);
or U24441 (N_24441,N_19195,N_16763);
and U24442 (N_24442,N_19797,N_17798);
nand U24443 (N_24443,N_18346,N_17098);
and U24444 (N_24444,N_17648,N_16811);
xnor U24445 (N_24445,N_19000,N_18201);
nor U24446 (N_24446,N_16183,N_16779);
or U24447 (N_24447,N_16094,N_15666);
and U24448 (N_24448,N_18584,N_17666);
and U24449 (N_24449,N_16482,N_18726);
xor U24450 (N_24450,N_18484,N_17724);
and U24451 (N_24451,N_17355,N_17773);
nor U24452 (N_24452,N_17286,N_16246);
nand U24453 (N_24453,N_19987,N_17881);
nor U24454 (N_24454,N_17800,N_15333);
or U24455 (N_24455,N_16089,N_15471);
and U24456 (N_24456,N_16412,N_16331);
xor U24457 (N_24457,N_18022,N_18929);
and U24458 (N_24458,N_19024,N_16438);
nand U24459 (N_24459,N_17432,N_15560);
or U24460 (N_24460,N_19205,N_15421);
and U24461 (N_24461,N_16095,N_19585);
or U24462 (N_24462,N_17923,N_16657);
or U24463 (N_24463,N_18498,N_17980);
nor U24464 (N_24464,N_18170,N_17290);
nor U24465 (N_24465,N_15579,N_15505);
xnor U24466 (N_24466,N_18895,N_15748);
or U24467 (N_24467,N_16193,N_15797);
xor U24468 (N_24468,N_15572,N_15634);
or U24469 (N_24469,N_19204,N_15312);
nand U24470 (N_24470,N_18744,N_17900);
and U24471 (N_24471,N_18642,N_17061);
or U24472 (N_24472,N_15206,N_18117);
and U24473 (N_24473,N_15026,N_15281);
xnor U24474 (N_24474,N_15606,N_18596);
or U24475 (N_24475,N_18220,N_16863);
nor U24476 (N_24476,N_17887,N_15144);
nand U24477 (N_24477,N_19544,N_17331);
nand U24478 (N_24478,N_18331,N_19117);
or U24479 (N_24479,N_15992,N_16563);
nor U24480 (N_24480,N_16786,N_15071);
xnor U24481 (N_24481,N_17563,N_19053);
and U24482 (N_24482,N_17297,N_18144);
and U24483 (N_24483,N_15832,N_19604);
nand U24484 (N_24484,N_18145,N_17043);
nand U24485 (N_24485,N_15417,N_17921);
or U24486 (N_24486,N_18451,N_17610);
nand U24487 (N_24487,N_15023,N_18724);
nand U24488 (N_24488,N_18434,N_16675);
nand U24489 (N_24489,N_19062,N_19463);
xnor U24490 (N_24490,N_18780,N_18985);
nand U24491 (N_24491,N_16583,N_15994);
xnor U24492 (N_24492,N_16374,N_16548);
and U24493 (N_24493,N_17239,N_19822);
xor U24494 (N_24494,N_16691,N_17978);
and U24495 (N_24495,N_17612,N_16795);
nand U24496 (N_24496,N_15893,N_15327);
xnor U24497 (N_24497,N_19269,N_15604);
and U24498 (N_24498,N_15644,N_16845);
nand U24499 (N_24499,N_19160,N_15655);
and U24500 (N_24500,N_16340,N_19130);
xor U24501 (N_24501,N_18138,N_19838);
nor U24502 (N_24502,N_15705,N_18093);
xor U24503 (N_24503,N_17920,N_16021);
and U24504 (N_24504,N_16859,N_19735);
nand U24505 (N_24505,N_15225,N_15865);
and U24506 (N_24506,N_16723,N_18439);
xor U24507 (N_24507,N_17331,N_17855);
xnor U24508 (N_24508,N_15514,N_17990);
or U24509 (N_24509,N_15971,N_15252);
nand U24510 (N_24510,N_16159,N_15480);
nor U24511 (N_24511,N_17048,N_15816);
nand U24512 (N_24512,N_16399,N_15026);
or U24513 (N_24513,N_15844,N_19164);
xnor U24514 (N_24514,N_16939,N_19831);
nand U24515 (N_24515,N_18961,N_18033);
nand U24516 (N_24516,N_18140,N_18832);
and U24517 (N_24517,N_19092,N_19826);
and U24518 (N_24518,N_18286,N_15902);
or U24519 (N_24519,N_16252,N_16815);
nor U24520 (N_24520,N_15413,N_15246);
xnor U24521 (N_24521,N_18684,N_18595);
or U24522 (N_24522,N_19041,N_18819);
nand U24523 (N_24523,N_15846,N_18044);
and U24524 (N_24524,N_19075,N_17279);
xnor U24525 (N_24525,N_19106,N_18276);
nand U24526 (N_24526,N_19974,N_19548);
nor U24527 (N_24527,N_15306,N_17604);
nand U24528 (N_24528,N_18848,N_16889);
or U24529 (N_24529,N_16736,N_15501);
or U24530 (N_24530,N_15346,N_19316);
nand U24531 (N_24531,N_18320,N_15000);
xnor U24532 (N_24532,N_19166,N_19311);
nor U24533 (N_24533,N_18319,N_15534);
xnor U24534 (N_24534,N_15060,N_18574);
or U24535 (N_24535,N_18534,N_16110);
xor U24536 (N_24536,N_19993,N_16751);
and U24537 (N_24537,N_18504,N_18060);
or U24538 (N_24538,N_16008,N_16132);
xnor U24539 (N_24539,N_15876,N_17664);
or U24540 (N_24540,N_17711,N_19344);
and U24541 (N_24541,N_18551,N_16018);
and U24542 (N_24542,N_17171,N_17752);
nand U24543 (N_24543,N_19831,N_18955);
and U24544 (N_24544,N_18614,N_16778);
and U24545 (N_24545,N_18906,N_15507);
and U24546 (N_24546,N_18298,N_16858);
xor U24547 (N_24547,N_16415,N_18474);
or U24548 (N_24548,N_15166,N_17047);
and U24549 (N_24549,N_17683,N_18881);
nor U24550 (N_24550,N_15154,N_16209);
or U24551 (N_24551,N_16505,N_17407);
xor U24552 (N_24552,N_15314,N_15787);
xor U24553 (N_24553,N_18483,N_17668);
or U24554 (N_24554,N_19725,N_16660);
and U24555 (N_24555,N_19934,N_16659);
xnor U24556 (N_24556,N_18836,N_16528);
xor U24557 (N_24557,N_15611,N_16656);
or U24558 (N_24558,N_15238,N_17104);
nand U24559 (N_24559,N_18634,N_16710);
nor U24560 (N_24560,N_19626,N_18289);
or U24561 (N_24561,N_19046,N_16756);
nor U24562 (N_24562,N_19461,N_16965);
xor U24563 (N_24563,N_19558,N_15099);
and U24564 (N_24564,N_16716,N_17669);
nor U24565 (N_24565,N_18288,N_19305);
nand U24566 (N_24566,N_17326,N_16300);
and U24567 (N_24567,N_17438,N_19093);
nand U24568 (N_24568,N_15432,N_16099);
or U24569 (N_24569,N_17671,N_18769);
or U24570 (N_24570,N_17656,N_16561);
and U24571 (N_24571,N_16578,N_19107);
or U24572 (N_24572,N_16915,N_16743);
nand U24573 (N_24573,N_19003,N_17026);
and U24574 (N_24574,N_19104,N_19890);
xnor U24575 (N_24575,N_18211,N_15953);
or U24576 (N_24576,N_16187,N_17390);
and U24577 (N_24577,N_16273,N_15884);
and U24578 (N_24578,N_19231,N_15102);
and U24579 (N_24579,N_17713,N_17342);
and U24580 (N_24580,N_15521,N_15245);
xnor U24581 (N_24581,N_18164,N_18279);
or U24582 (N_24582,N_17255,N_18298);
or U24583 (N_24583,N_17550,N_19292);
xor U24584 (N_24584,N_16729,N_19940);
nor U24585 (N_24585,N_15477,N_15323);
or U24586 (N_24586,N_18790,N_18655);
or U24587 (N_24587,N_18726,N_19653);
xnor U24588 (N_24588,N_19648,N_18091);
or U24589 (N_24589,N_15071,N_15179);
nor U24590 (N_24590,N_19349,N_16901);
or U24591 (N_24591,N_15184,N_16058);
nor U24592 (N_24592,N_18467,N_18417);
nand U24593 (N_24593,N_19004,N_18453);
nor U24594 (N_24594,N_16872,N_19355);
xnor U24595 (N_24595,N_18532,N_18749);
nor U24596 (N_24596,N_18617,N_16422);
nor U24597 (N_24597,N_15095,N_15710);
nor U24598 (N_24598,N_15686,N_17285);
nor U24599 (N_24599,N_15465,N_16934);
xor U24600 (N_24600,N_17466,N_19321);
or U24601 (N_24601,N_19108,N_16381);
nand U24602 (N_24602,N_16429,N_18063);
nor U24603 (N_24603,N_18842,N_17722);
xnor U24604 (N_24604,N_17148,N_16143);
and U24605 (N_24605,N_19068,N_16888);
xnor U24606 (N_24606,N_19409,N_16138);
and U24607 (N_24607,N_16565,N_18153);
xnor U24608 (N_24608,N_17713,N_18137);
nand U24609 (N_24609,N_17293,N_16283);
nand U24610 (N_24610,N_15224,N_19371);
nand U24611 (N_24611,N_18230,N_16082);
xor U24612 (N_24612,N_18671,N_18089);
nand U24613 (N_24613,N_15388,N_16886);
nor U24614 (N_24614,N_16814,N_16472);
nand U24615 (N_24615,N_15554,N_16142);
xnor U24616 (N_24616,N_18396,N_18329);
nor U24617 (N_24617,N_15728,N_17442);
or U24618 (N_24618,N_15508,N_16060);
xor U24619 (N_24619,N_15952,N_18595);
or U24620 (N_24620,N_16987,N_16015);
nand U24621 (N_24621,N_17498,N_17864);
nor U24622 (N_24622,N_18470,N_16282);
or U24623 (N_24623,N_18817,N_16104);
nor U24624 (N_24624,N_16507,N_16185);
nor U24625 (N_24625,N_19430,N_19894);
nor U24626 (N_24626,N_19155,N_15674);
and U24627 (N_24627,N_19136,N_18943);
nand U24628 (N_24628,N_17601,N_16073);
nor U24629 (N_24629,N_16242,N_19938);
or U24630 (N_24630,N_19826,N_15995);
and U24631 (N_24631,N_18684,N_17060);
and U24632 (N_24632,N_18928,N_18333);
xor U24633 (N_24633,N_16016,N_17475);
and U24634 (N_24634,N_19981,N_19732);
nor U24635 (N_24635,N_19923,N_17884);
nand U24636 (N_24636,N_19663,N_19409);
and U24637 (N_24637,N_15418,N_18689);
nand U24638 (N_24638,N_19924,N_18544);
or U24639 (N_24639,N_19478,N_16592);
or U24640 (N_24640,N_18595,N_18341);
nand U24641 (N_24641,N_15516,N_17986);
or U24642 (N_24642,N_17962,N_18578);
nor U24643 (N_24643,N_19477,N_15172);
or U24644 (N_24644,N_15292,N_18635);
nand U24645 (N_24645,N_17748,N_16674);
xnor U24646 (N_24646,N_15577,N_18169);
or U24647 (N_24647,N_15855,N_19100);
nand U24648 (N_24648,N_18720,N_18552);
or U24649 (N_24649,N_17500,N_18698);
xor U24650 (N_24650,N_15446,N_19888);
or U24651 (N_24651,N_17076,N_15131);
and U24652 (N_24652,N_18876,N_19161);
and U24653 (N_24653,N_16881,N_16645);
or U24654 (N_24654,N_18561,N_18463);
xor U24655 (N_24655,N_17332,N_18158);
nor U24656 (N_24656,N_16507,N_17591);
and U24657 (N_24657,N_19424,N_15133);
nand U24658 (N_24658,N_17700,N_16479);
nand U24659 (N_24659,N_18874,N_18596);
and U24660 (N_24660,N_19835,N_15956);
nand U24661 (N_24661,N_15997,N_17063);
or U24662 (N_24662,N_16953,N_17437);
nor U24663 (N_24663,N_15544,N_19998);
nor U24664 (N_24664,N_19432,N_15682);
and U24665 (N_24665,N_15106,N_17021);
and U24666 (N_24666,N_17403,N_16701);
or U24667 (N_24667,N_19070,N_19165);
and U24668 (N_24668,N_15752,N_17927);
or U24669 (N_24669,N_15682,N_18230);
or U24670 (N_24670,N_15601,N_19231);
nor U24671 (N_24671,N_15288,N_19226);
nand U24672 (N_24672,N_19480,N_15042);
nor U24673 (N_24673,N_15998,N_19355);
xnor U24674 (N_24674,N_15687,N_18806);
nor U24675 (N_24675,N_15307,N_17135);
or U24676 (N_24676,N_15237,N_16982);
or U24677 (N_24677,N_19565,N_16423);
xor U24678 (N_24678,N_15032,N_15274);
and U24679 (N_24679,N_18178,N_19555);
xor U24680 (N_24680,N_18220,N_15418);
xnor U24681 (N_24681,N_18794,N_18592);
xnor U24682 (N_24682,N_19351,N_19174);
nand U24683 (N_24683,N_17173,N_17819);
xor U24684 (N_24684,N_15720,N_16821);
or U24685 (N_24685,N_15802,N_16072);
or U24686 (N_24686,N_18976,N_19266);
xor U24687 (N_24687,N_15840,N_18293);
nor U24688 (N_24688,N_15296,N_16363);
xnor U24689 (N_24689,N_16620,N_17778);
nand U24690 (N_24690,N_15499,N_16508);
xor U24691 (N_24691,N_16429,N_16054);
nor U24692 (N_24692,N_16508,N_17621);
nand U24693 (N_24693,N_15884,N_16081);
or U24694 (N_24694,N_16450,N_16853);
nor U24695 (N_24695,N_17784,N_15050);
nand U24696 (N_24696,N_16515,N_18463);
or U24697 (N_24697,N_16490,N_19963);
xnor U24698 (N_24698,N_19119,N_16257);
xor U24699 (N_24699,N_18939,N_19735);
or U24700 (N_24700,N_16209,N_15081);
and U24701 (N_24701,N_19118,N_19449);
xnor U24702 (N_24702,N_17523,N_16714);
xnor U24703 (N_24703,N_16076,N_15915);
and U24704 (N_24704,N_19118,N_17987);
xor U24705 (N_24705,N_19887,N_15915);
nor U24706 (N_24706,N_15988,N_15073);
xnor U24707 (N_24707,N_17965,N_16319);
nand U24708 (N_24708,N_15840,N_19400);
nand U24709 (N_24709,N_15258,N_19960);
and U24710 (N_24710,N_16419,N_15379);
nor U24711 (N_24711,N_19452,N_18238);
nor U24712 (N_24712,N_18992,N_18924);
nand U24713 (N_24713,N_19569,N_19785);
nand U24714 (N_24714,N_16422,N_15026);
nand U24715 (N_24715,N_19915,N_17048);
nor U24716 (N_24716,N_16464,N_16495);
and U24717 (N_24717,N_15300,N_16111);
xnor U24718 (N_24718,N_16430,N_18980);
or U24719 (N_24719,N_15775,N_16137);
nor U24720 (N_24720,N_19277,N_17014);
xnor U24721 (N_24721,N_15723,N_18094);
nor U24722 (N_24722,N_16391,N_17284);
xor U24723 (N_24723,N_17709,N_19548);
nand U24724 (N_24724,N_19267,N_17429);
xor U24725 (N_24725,N_15798,N_19547);
nand U24726 (N_24726,N_15629,N_16281);
nor U24727 (N_24727,N_15193,N_18627);
or U24728 (N_24728,N_16762,N_19404);
and U24729 (N_24729,N_19183,N_18250);
and U24730 (N_24730,N_17922,N_15194);
and U24731 (N_24731,N_18044,N_16237);
and U24732 (N_24732,N_19361,N_16718);
and U24733 (N_24733,N_16411,N_17294);
or U24734 (N_24734,N_16119,N_19740);
nor U24735 (N_24735,N_15380,N_19355);
or U24736 (N_24736,N_16831,N_18601);
or U24737 (N_24737,N_19454,N_19612);
or U24738 (N_24738,N_15201,N_15701);
nand U24739 (N_24739,N_19370,N_15559);
nand U24740 (N_24740,N_18844,N_19770);
and U24741 (N_24741,N_16167,N_17567);
nor U24742 (N_24742,N_17046,N_16727);
nor U24743 (N_24743,N_19298,N_16234);
or U24744 (N_24744,N_18480,N_19642);
nand U24745 (N_24745,N_16945,N_17731);
nor U24746 (N_24746,N_15152,N_19253);
xor U24747 (N_24747,N_18994,N_18902);
or U24748 (N_24748,N_19304,N_17643);
nand U24749 (N_24749,N_18839,N_18954);
and U24750 (N_24750,N_16393,N_17386);
and U24751 (N_24751,N_19974,N_18962);
nand U24752 (N_24752,N_16144,N_18385);
and U24753 (N_24753,N_19845,N_17958);
xor U24754 (N_24754,N_19180,N_16185);
nor U24755 (N_24755,N_19962,N_16725);
or U24756 (N_24756,N_17883,N_19113);
nor U24757 (N_24757,N_15132,N_19289);
xnor U24758 (N_24758,N_17411,N_16953);
nand U24759 (N_24759,N_16941,N_19704);
nand U24760 (N_24760,N_18980,N_18518);
nand U24761 (N_24761,N_17764,N_19680);
nor U24762 (N_24762,N_15248,N_18756);
nand U24763 (N_24763,N_19284,N_16280);
xnor U24764 (N_24764,N_17444,N_17067);
nand U24765 (N_24765,N_16251,N_19747);
or U24766 (N_24766,N_18990,N_19013);
nor U24767 (N_24767,N_19277,N_19782);
xor U24768 (N_24768,N_17420,N_15379);
or U24769 (N_24769,N_16962,N_15979);
or U24770 (N_24770,N_18905,N_17972);
nand U24771 (N_24771,N_18519,N_15389);
or U24772 (N_24772,N_18186,N_15106);
xnor U24773 (N_24773,N_15597,N_16400);
xor U24774 (N_24774,N_15621,N_18309);
xnor U24775 (N_24775,N_19937,N_18265);
xnor U24776 (N_24776,N_16617,N_15425);
or U24777 (N_24777,N_19543,N_17215);
or U24778 (N_24778,N_19110,N_19913);
nor U24779 (N_24779,N_19944,N_18494);
nor U24780 (N_24780,N_15973,N_16887);
nand U24781 (N_24781,N_18169,N_17988);
or U24782 (N_24782,N_17414,N_18661);
xnor U24783 (N_24783,N_18605,N_18286);
and U24784 (N_24784,N_15689,N_17623);
and U24785 (N_24785,N_18972,N_16951);
xor U24786 (N_24786,N_17722,N_17015);
nand U24787 (N_24787,N_19687,N_16226);
or U24788 (N_24788,N_18279,N_16521);
nand U24789 (N_24789,N_15923,N_18696);
xnor U24790 (N_24790,N_19412,N_19053);
nand U24791 (N_24791,N_16329,N_17774);
xnor U24792 (N_24792,N_16569,N_15807);
nor U24793 (N_24793,N_15040,N_19705);
nand U24794 (N_24794,N_16681,N_19370);
and U24795 (N_24795,N_16528,N_16431);
nor U24796 (N_24796,N_17479,N_18287);
or U24797 (N_24797,N_16786,N_18766);
nand U24798 (N_24798,N_15481,N_17204);
nor U24799 (N_24799,N_18320,N_18918);
nand U24800 (N_24800,N_19845,N_18946);
nand U24801 (N_24801,N_18912,N_16268);
and U24802 (N_24802,N_18129,N_15675);
or U24803 (N_24803,N_15121,N_15458);
nand U24804 (N_24804,N_18798,N_17931);
nand U24805 (N_24805,N_17662,N_18023);
nand U24806 (N_24806,N_17655,N_18088);
nand U24807 (N_24807,N_17727,N_15836);
xnor U24808 (N_24808,N_18418,N_16789);
nand U24809 (N_24809,N_19878,N_17567);
xor U24810 (N_24810,N_15579,N_18721);
or U24811 (N_24811,N_16981,N_18250);
and U24812 (N_24812,N_17231,N_18622);
and U24813 (N_24813,N_17531,N_16483);
or U24814 (N_24814,N_19299,N_15814);
nand U24815 (N_24815,N_18721,N_18373);
and U24816 (N_24816,N_16581,N_15784);
xnor U24817 (N_24817,N_18055,N_16266);
and U24818 (N_24818,N_18439,N_17596);
xnor U24819 (N_24819,N_18254,N_19571);
xor U24820 (N_24820,N_18964,N_16052);
nor U24821 (N_24821,N_19741,N_16075);
nor U24822 (N_24822,N_18514,N_15406);
xor U24823 (N_24823,N_17066,N_18193);
or U24824 (N_24824,N_19229,N_17799);
nor U24825 (N_24825,N_18009,N_19916);
or U24826 (N_24826,N_19540,N_15621);
nand U24827 (N_24827,N_16422,N_18227);
xor U24828 (N_24828,N_19561,N_15793);
or U24829 (N_24829,N_17322,N_16381);
or U24830 (N_24830,N_16117,N_15088);
and U24831 (N_24831,N_17400,N_18867);
nand U24832 (N_24832,N_19958,N_16892);
xnor U24833 (N_24833,N_16356,N_17433);
nor U24834 (N_24834,N_18188,N_15050);
or U24835 (N_24835,N_19530,N_18663);
or U24836 (N_24836,N_19389,N_16346);
and U24837 (N_24837,N_19906,N_17973);
or U24838 (N_24838,N_18731,N_19211);
nand U24839 (N_24839,N_17066,N_15357);
and U24840 (N_24840,N_19475,N_19210);
or U24841 (N_24841,N_17365,N_17734);
and U24842 (N_24842,N_16869,N_15560);
nor U24843 (N_24843,N_18344,N_16383);
and U24844 (N_24844,N_18256,N_18761);
and U24845 (N_24845,N_18004,N_17819);
xnor U24846 (N_24846,N_15836,N_16573);
nor U24847 (N_24847,N_18389,N_18260);
and U24848 (N_24848,N_19142,N_16999);
and U24849 (N_24849,N_16624,N_15647);
xor U24850 (N_24850,N_19638,N_17939);
nand U24851 (N_24851,N_17090,N_19304);
nand U24852 (N_24852,N_19975,N_18019);
and U24853 (N_24853,N_19829,N_17256);
nand U24854 (N_24854,N_19585,N_17192);
or U24855 (N_24855,N_19699,N_19643);
or U24856 (N_24856,N_15283,N_16299);
xor U24857 (N_24857,N_19623,N_19312);
and U24858 (N_24858,N_16424,N_19770);
xor U24859 (N_24859,N_16238,N_19931);
nor U24860 (N_24860,N_19586,N_17749);
xor U24861 (N_24861,N_19299,N_17655);
nand U24862 (N_24862,N_18174,N_18895);
nor U24863 (N_24863,N_15200,N_15458);
xnor U24864 (N_24864,N_15585,N_16644);
and U24865 (N_24865,N_17918,N_16044);
and U24866 (N_24866,N_17490,N_17028);
or U24867 (N_24867,N_15973,N_15895);
nand U24868 (N_24868,N_17075,N_16874);
or U24869 (N_24869,N_15890,N_18490);
nor U24870 (N_24870,N_16197,N_17668);
nor U24871 (N_24871,N_18828,N_18393);
or U24872 (N_24872,N_16399,N_18266);
or U24873 (N_24873,N_18921,N_19631);
xor U24874 (N_24874,N_19391,N_17662);
nand U24875 (N_24875,N_15555,N_15045);
and U24876 (N_24876,N_19411,N_17083);
xnor U24877 (N_24877,N_16816,N_15475);
and U24878 (N_24878,N_16801,N_17428);
nand U24879 (N_24879,N_18248,N_15175);
nand U24880 (N_24880,N_15578,N_17174);
xnor U24881 (N_24881,N_18059,N_19151);
and U24882 (N_24882,N_16114,N_16785);
xor U24883 (N_24883,N_19576,N_15014);
xnor U24884 (N_24884,N_17153,N_17814);
and U24885 (N_24885,N_19761,N_15698);
xor U24886 (N_24886,N_18188,N_17124);
nand U24887 (N_24887,N_17482,N_16418);
nand U24888 (N_24888,N_18857,N_15151);
nand U24889 (N_24889,N_18218,N_15505);
nor U24890 (N_24890,N_18324,N_19287);
or U24891 (N_24891,N_18431,N_16213);
and U24892 (N_24892,N_19799,N_16488);
or U24893 (N_24893,N_17502,N_16626);
nand U24894 (N_24894,N_15346,N_18550);
and U24895 (N_24895,N_19304,N_19965);
and U24896 (N_24896,N_18970,N_16538);
nand U24897 (N_24897,N_17746,N_18490);
or U24898 (N_24898,N_18012,N_17839);
or U24899 (N_24899,N_15623,N_15534);
nand U24900 (N_24900,N_16487,N_16662);
or U24901 (N_24901,N_18210,N_17363);
and U24902 (N_24902,N_15386,N_15043);
or U24903 (N_24903,N_17240,N_15138);
or U24904 (N_24904,N_17544,N_19484);
and U24905 (N_24905,N_18238,N_15953);
nand U24906 (N_24906,N_16980,N_16303);
nor U24907 (N_24907,N_18266,N_19616);
and U24908 (N_24908,N_15138,N_18188);
nand U24909 (N_24909,N_19919,N_16416);
or U24910 (N_24910,N_16525,N_17007);
or U24911 (N_24911,N_15373,N_17949);
xnor U24912 (N_24912,N_15289,N_16172);
nand U24913 (N_24913,N_19575,N_17032);
or U24914 (N_24914,N_17003,N_15283);
nand U24915 (N_24915,N_15553,N_17900);
xnor U24916 (N_24916,N_18828,N_18640);
xnor U24917 (N_24917,N_16446,N_15645);
or U24918 (N_24918,N_17234,N_16855);
nor U24919 (N_24919,N_16973,N_17543);
and U24920 (N_24920,N_18137,N_16156);
or U24921 (N_24921,N_19576,N_18451);
xor U24922 (N_24922,N_19101,N_15295);
or U24923 (N_24923,N_16158,N_19170);
or U24924 (N_24924,N_16998,N_18168);
nor U24925 (N_24925,N_16137,N_18442);
nand U24926 (N_24926,N_15459,N_16198);
xor U24927 (N_24927,N_16198,N_15642);
xnor U24928 (N_24928,N_19123,N_18618);
and U24929 (N_24929,N_19501,N_17939);
and U24930 (N_24930,N_15848,N_15185);
nor U24931 (N_24931,N_16562,N_15888);
nand U24932 (N_24932,N_18154,N_18802);
and U24933 (N_24933,N_17681,N_16490);
nor U24934 (N_24934,N_16981,N_15826);
and U24935 (N_24935,N_16738,N_16523);
xor U24936 (N_24936,N_18739,N_19705);
xor U24937 (N_24937,N_16024,N_17712);
nor U24938 (N_24938,N_16971,N_15378);
nor U24939 (N_24939,N_15635,N_19456);
xnor U24940 (N_24940,N_17490,N_16807);
or U24941 (N_24941,N_15864,N_19311);
or U24942 (N_24942,N_15247,N_16787);
and U24943 (N_24943,N_18622,N_16919);
nand U24944 (N_24944,N_17885,N_16340);
and U24945 (N_24945,N_15815,N_15070);
nor U24946 (N_24946,N_19088,N_15575);
xor U24947 (N_24947,N_15867,N_18175);
nand U24948 (N_24948,N_16284,N_17028);
xnor U24949 (N_24949,N_16274,N_17022);
and U24950 (N_24950,N_16036,N_16256);
xnor U24951 (N_24951,N_16341,N_15369);
xor U24952 (N_24952,N_17436,N_15609);
nor U24953 (N_24953,N_17734,N_16287);
or U24954 (N_24954,N_19613,N_19095);
and U24955 (N_24955,N_17559,N_19347);
and U24956 (N_24956,N_18527,N_16818);
and U24957 (N_24957,N_16349,N_16948);
and U24958 (N_24958,N_17249,N_18367);
xor U24959 (N_24959,N_19329,N_19568);
and U24960 (N_24960,N_17183,N_15677);
xor U24961 (N_24961,N_16612,N_19348);
and U24962 (N_24962,N_18650,N_18100);
nor U24963 (N_24963,N_17348,N_16872);
and U24964 (N_24964,N_15083,N_15366);
or U24965 (N_24965,N_15981,N_19823);
or U24966 (N_24966,N_17686,N_17432);
nand U24967 (N_24967,N_18207,N_16690);
and U24968 (N_24968,N_16304,N_18864);
and U24969 (N_24969,N_17532,N_17280);
or U24970 (N_24970,N_16316,N_17045);
nor U24971 (N_24971,N_17230,N_18182);
nor U24972 (N_24972,N_16621,N_16055);
and U24973 (N_24973,N_19623,N_18398);
or U24974 (N_24974,N_15878,N_15603);
and U24975 (N_24975,N_19642,N_16197);
nor U24976 (N_24976,N_15960,N_16649);
nor U24977 (N_24977,N_16471,N_15293);
nand U24978 (N_24978,N_17717,N_17467);
and U24979 (N_24979,N_17862,N_17594);
nor U24980 (N_24980,N_18165,N_19436);
or U24981 (N_24981,N_19371,N_19028);
xnor U24982 (N_24982,N_15015,N_16047);
or U24983 (N_24983,N_15259,N_15665);
nand U24984 (N_24984,N_19506,N_15075);
xor U24985 (N_24985,N_19937,N_16758);
xnor U24986 (N_24986,N_16660,N_18310);
or U24987 (N_24987,N_19850,N_17855);
xor U24988 (N_24988,N_15632,N_18765);
nor U24989 (N_24989,N_19638,N_19851);
and U24990 (N_24990,N_15614,N_19150);
xor U24991 (N_24991,N_19421,N_17656);
xor U24992 (N_24992,N_18164,N_17435);
and U24993 (N_24993,N_17220,N_18585);
and U24994 (N_24994,N_15557,N_16988);
or U24995 (N_24995,N_15323,N_17707);
and U24996 (N_24996,N_17579,N_16947);
xnor U24997 (N_24997,N_15139,N_19885);
nand U24998 (N_24998,N_15404,N_16836);
or U24999 (N_24999,N_19648,N_15098);
nor U25000 (N_25000,N_24278,N_23906);
and U25001 (N_25001,N_23137,N_20894);
xor U25002 (N_25002,N_24657,N_21501);
nand U25003 (N_25003,N_20772,N_20814);
and U25004 (N_25004,N_21106,N_20959);
nand U25005 (N_25005,N_24312,N_22596);
nand U25006 (N_25006,N_23878,N_21203);
nor U25007 (N_25007,N_24854,N_21337);
or U25008 (N_25008,N_23218,N_20861);
and U25009 (N_25009,N_22115,N_24148);
or U25010 (N_25010,N_22559,N_23469);
nand U25011 (N_25011,N_23445,N_23520);
and U25012 (N_25012,N_21594,N_22166);
and U25013 (N_25013,N_23889,N_23779);
nor U25014 (N_25014,N_22240,N_20131);
or U25015 (N_25015,N_24228,N_22825);
nand U25016 (N_25016,N_24077,N_22198);
nand U25017 (N_25017,N_23385,N_20052);
nor U25018 (N_25018,N_20543,N_21842);
nand U25019 (N_25019,N_24808,N_24646);
xnor U25020 (N_25020,N_21676,N_20442);
and U25021 (N_25021,N_22474,N_23991);
nor U25022 (N_25022,N_23701,N_21772);
and U25023 (N_25023,N_20172,N_22645);
xnor U25024 (N_25024,N_20651,N_23910);
nand U25025 (N_25025,N_20527,N_23332);
nand U25026 (N_25026,N_24789,N_23432);
nor U25027 (N_25027,N_21146,N_22827);
xnor U25028 (N_25028,N_23002,N_21429);
or U25029 (N_25029,N_21157,N_24366);
nand U25030 (N_25030,N_20314,N_23909);
or U25031 (N_25031,N_21502,N_23744);
xor U25032 (N_25032,N_22059,N_24391);
nand U25033 (N_25033,N_23656,N_22872);
or U25034 (N_25034,N_22582,N_22100);
or U25035 (N_25035,N_20072,N_21006);
nor U25036 (N_25036,N_23290,N_24403);
nor U25037 (N_25037,N_24971,N_24661);
nand U25038 (N_25038,N_20636,N_23425);
and U25039 (N_25039,N_21549,N_20080);
nand U25040 (N_25040,N_20617,N_21237);
nand U25041 (N_25041,N_22310,N_20634);
nand U25042 (N_25042,N_21172,N_23157);
nand U25043 (N_25043,N_23920,N_24119);
nand U25044 (N_25044,N_23552,N_22667);
and U25045 (N_25045,N_20471,N_20969);
nor U25046 (N_25046,N_24844,N_24212);
xnor U25047 (N_25047,N_20414,N_21878);
nand U25048 (N_25048,N_22085,N_21789);
and U25049 (N_25049,N_21829,N_22615);
nand U25050 (N_25050,N_21022,N_22533);
xor U25051 (N_25051,N_21833,N_22965);
nand U25052 (N_25052,N_23117,N_23621);
or U25053 (N_25053,N_20307,N_21513);
nor U25054 (N_25054,N_21343,N_23562);
and U25055 (N_25055,N_23073,N_24383);
and U25056 (N_25056,N_23093,N_23817);
or U25057 (N_25057,N_20707,N_22684);
nand U25058 (N_25058,N_20335,N_20087);
xnor U25059 (N_25059,N_21793,N_24457);
nand U25060 (N_25060,N_24286,N_20368);
and U25061 (N_25061,N_21330,N_21184);
and U25062 (N_25062,N_22573,N_23215);
nor U25063 (N_25063,N_21084,N_22584);
nand U25064 (N_25064,N_23083,N_20841);
nor U25065 (N_25065,N_24542,N_21820);
xor U25066 (N_25066,N_24563,N_21065);
nor U25067 (N_25067,N_24802,N_22586);
nand U25068 (N_25068,N_20542,N_23072);
nand U25069 (N_25069,N_22818,N_23649);
xnor U25070 (N_25070,N_21450,N_20317);
and U25071 (N_25071,N_21127,N_20924);
xor U25072 (N_25072,N_23370,N_23677);
or U25073 (N_25073,N_20141,N_23455);
or U25074 (N_25074,N_24258,N_22091);
nand U25075 (N_25075,N_22366,N_22799);
nor U25076 (N_25076,N_21749,N_20182);
xnor U25077 (N_25077,N_21865,N_21807);
and U25078 (N_25078,N_24583,N_22689);
or U25079 (N_25079,N_22478,N_20193);
nand U25080 (N_25080,N_23726,N_22096);
or U25081 (N_25081,N_23317,N_22755);
nor U25082 (N_25082,N_21327,N_24071);
or U25083 (N_25083,N_22155,N_22647);
xnor U25084 (N_25084,N_20743,N_24160);
or U25085 (N_25085,N_20833,N_20316);
nand U25086 (N_25086,N_23278,N_21167);
nand U25087 (N_25087,N_24045,N_20941);
nand U25088 (N_25088,N_22433,N_22677);
nor U25089 (N_25089,N_20461,N_23930);
xnor U25090 (N_25090,N_22668,N_22144);
nand U25091 (N_25091,N_21632,N_24894);
nor U25092 (N_25092,N_21916,N_23129);
or U25093 (N_25093,N_21870,N_20809);
or U25094 (N_25094,N_21151,N_24845);
or U25095 (N_25095,N_20697,N_24096);
and U25096 (N_25096,N_20069,N_24779);
nand U25097 (N_25097,N_24699,N_24612);
and U25098 (N_25098,N_23020,N_24952);
nor U25099 (N_25099,N_24197,N_23985);
xnor U25100 (N_25100,N_20706,N_20904);
and U25101 (N_25101,N_20535,N_21741);
nor U25102 (N_25102,N_20822,N_24310);
or U25103 (N_25103,N_20658,N_24414);
xor U25104 (N_25104,N_21178,N_20585);
nand U25105 (N_25105,N_22900,N_22698);
xor U25106 (N_25106,N_24996,N_21664);
and U25107 (N_25107,N_24118,N_20023);
nor U25108 (N_25108,N_24560,N_21618);
nand U25109 (N_25109,N_20176,N_21097);
xor U25110 (N_25110,N_23448,N_23706);
nor U25111 (N_25111,N_24085,N_21525);
xnor U25112 (N_25112,N_24384,N_21771);
nand U25113 (N_25113,N_21375,N_21145);
xor U25114 (N_25114,N_23619,N_24595);
and U25115 (N_25115,N_20887,N_20754);
xor U25116 (N_25116,N_24574,N_22968);
or U25117 (N_25117,N_24040,N_23565);
or U25118 (N_25118,N_20662,N_24203);
xnor U25119 (N_25119,N_24929,N_23516);
nor U25120 (N_25120,N_23021,N_24579);
xnor U25121 (N_25121,N_20359,N_20392);
or U25122 (N_25122,N_21076,N_20510);
or U25123 (N_25123,N_21536,N_21510);
xnor U25124 (N_25124,N_23859,N_23025);
nand U25125 (N_25125,N_21709,N_21242);
xor U25126 (N_25126,N_20839,N_23932);
nand U25127 (N_25127,N_20831,N_20294);
xnor U25128 (N_25128,N_21869,N_20277);
xor U25129 (N_25129,N_22682,N_21174);
or U25130 (N_25130,N_21667,N_20411);
or U25131 (N_25131,N_24861,N_24857);
and U25132 (N_25132,N_22761,N_22153);
nor U25133 (N_25133,N_24164,N_23412);
or U25134 (N_25134,N_23915,N_23119);
and U25135 (N_25135,N_20209,N_24065);
nor U25136 (N_25136,N_24712,N_21049);
and U25137 (N_25137,N_23104,N_22276);
xor U25138 (N_25138,N_21665,N_22403);
nand U25139 (N_25139,N_23741,N_24448);
xor U25140 (N_25140,N_22214,N_21039);
nand U25141 (N_25141,N_22179,N_22369);
nand U25142 (N_25142,N_24274,N_21574);
or U25143 (N_25143,N_24733,N_20747);
xnor U25144 (N_25144,N_21126,N_24121);
nor U25145 (N_25145,N_23224,N_24573);
xor U25146 (N_25146,N_23230,N_22196);
nor U25147 (N_25147,N_24482,N_20818);
or U25148 (N_25148,N_23606,N_24248);
nor U25149 (N_25149,N_23330,N_21272);
xor U25150 (N_25150,N_24109,N_22109);
nor U25151 (N_25151,N_24257,N_21917);
or U25152 (N_25152,N_24876,N_23843);
and U25153 (N_25153,N_23705,N_20186);
or U25154 (N_25154,N_24667,N_21359);
nand U25155 (N_25155,N_22191,N_22726);
nand U25156 (N_25156,N_20273,N_22411);
and U25157 (N_25157,N_23981,N_22350);
nand U25158 (N_25158,N_20721,N_21317);
xor U25159 (N_25159,N_23989,N_24156);
and U25160 (N_25160,N_23257,N_24872);
and U25161 (N_25161,N_23814,N_21433);
xnor U25162 (N_25162,N_23854,N_23764);
nand U25163 (N_25163,N_23326,N_24389);
or U25164 (N_25164,N_20401,N_23426);
and U25165 (N_25165,N_23596,N_20106);
nor U25166 (N_25166,N_24903,N_22627);
xor U25167 (N_25167,N_20889,N_21773);
nor U25168 (N_25168,N_20219,N_23622);
or U25169 (N_25169,N_22526,N_22101);
nor U25170 (N_25170,N_23666,N_24027);
xor U25171 (N_25171,N_21743,N_22508);
and U25172 (N_25172,N_22847,N_24877);
or U25173 (N_25173,N_20019,N_20547);
xor U25174 (N_25174,N_24791,N_20583);
xor U25175 (N_25175,N_21406,N_22859);
nand U25176 (N_25176,N_23247,N_21357);
xor U25177 (N_25177,N_21465,N_20315);
xnor U25178 (N_25178,N_22282,N_20337);
nand U25179 (N_25179,N_23819,N_24581);
nor U25180 (N_25180,N_22235,N_22332);
or U25181 (N_25181,N_23947,N_22980);
or U25182 (N_25182,N_22485,N_24649);
xnor U25183 (N_25183,N_21716,N_21971);
nor U25184 (N_25184,N_21673,N_20105);
nand U25185 (N_25185,N_21363,N_21016);
xor U25186 (N_25186,N_23631,N_21800);
and U25187 (N_25187,N_24538,N_21404);
xnor U25188 (N_25188,N_22247,N_20781);
and U25189 (N_25189,N_22140,N_22700);
or U25190 (N_25190,N_23153,N_21976);
and U25191 (N_25191,N_21094,N_20823);
xor U25192 (N_25192,N_23777,N_24038);
or U25193 (N_25193,N_24343,N_20271);
nand U25194 (N_25194,N_22225,N_21722);
nor U25195 (N_25195,N_23686,N_23300);
and U25196 (N_25196,N_24735,N_22760);
nor U25197 (N_25197,N_20815,N_20264);
xnor U25198 (N_25198,N_22339,N_22583);
xor U25199 (N_25199,N_20526,N_23273);
and U25200 (N_25200,N_22525,N_23527);
and U25201 (N_25201,N_20464,N_24099);
nor U25202 (N_25202,N_24515,N_24994);
nand U25203 (N_25203,N_21496,N_24427);
and U25204 (N_25204,N_20241,N_23306);
xor U25205 (N_25205,N_23966,N_22763);
or U25206 (N_25206,N_22224,N_23390);
nor U25207 (N_25207,N_20654,N_22608);
and U25208 (N_25208,N_22076,N_22986);
nand U25209 (N_25209,N_20588,N_24732);
xor U25210 (N_25210,N_23776,N_20378);
nand U25211 (N_25211,N_21586,N_21364);
nor U25212 (N_25212,N_23479,N_24768);
and U25213 (N_25213,N_23751,N_22561);
nor U25214 (N_25214,N_21617,N_23407);
nor U25215 (N_25215,N_24607,N_24835);
xor U25216 (N_25216,N_20983,N_21639);
or U25217 (N_25217,N_20483,N_22896);
and U25218 (N_25218,N_24042,N_21810);
nand U25219 (N_25219,N_24587,N_24480);
or U25220 (N_25220,N_23387,N_20060);
xor U25221 (N_25221,N_23142,N_23891);
xnor U25222 (N_25222,N_23754,N_23853);
nor U25223 (N_25223,N_20263,N_22742);
xnor U25224 (N_25224,N_21652,N_22994);
nand U25225 (N_25225,N_20312,N_20986);
xnor U25226 (N_25226,N_24643,N_24433);
nand U25227 (N_25227,N_22190,N_24183);
nand U25228 (N_25228,N_20481,N_20003);
or U25229 (N_25229,N_24133,N_22547);
or U25230 (N_25230,N_22720,N_24984);
xnor U25231 (N_25231,N_23652,N_20285);
and U25232 (N_25232,N_21417,N_21284);
nor U25233 (N_25233,N_23654,N_24093);
xor U25234 (N_25234,N_22243,N_21514);
and U25235 (N_25235,N_20376,N_23048);
nor U25236 (N_25236,N_20750,N_23939);
or U25237 (N_25237,N_24311,N_22802);
nor U25238 (N_25238,N_22492,N_22165);
or U25239 (N_25239,N_22543,N_20643);
nand U25240 (N_25240,N_23762,N_21727);
or U25241 (N_25241,N_21655,N_23372);
and U25242 (N_25242,N_22598,N_22949);
nand U25243 (N_25243,N_23778,N_24316);
xor U25244 (N_25244,N_22992,N_21085);
or U25245 (N_25245,N_21958,N_21186);
and U25246 (N_25246,N_23862,N_23902);
or U25247 (N_25247,N_22323,N_22842);
nor U25248 (N_25248,N_20123,N_20239);
nand U25249 (N_25249,N_20455,N_24168);
nand U25250 (N_25250,N_23857,N_23155);
xor U25251 (N_25251,N_22920,N_23060);
nand U25252 (N_25252,N_21333,N_22538);
or U25253 (N_25253,N_22017,N_21908);
nor U25254 (N_25254,N_20421,N_22057);
or U25255 (N_25255,N_22367,N_24818);
nand U25256 (N_25256,N_23248,N_22452);
nand U25257 (N_25257,N_20567,N_20107);
and U25258 (N_25258,N_23279,N_22154);
nand U25259 (N_25259,N_22861,N_23844);
nand U25260 (N_25260,N_20898,N_22132);
xor U25261 (N_25261,N_24687,N_23265);
and U25262 (N_25262,N_24623,N_21608);
xnor U25263 (N_25263,N_22482,N_23995);
nand U25264 (N_25264,N_23447,N_21032);
or U25265 (N_25265,N_20674,N_20960);
nor U25266 (N_25266,N_21449,N_24362);
nand U25267 (N_25267,N_22618,N_21582);
and U25268 (N_25268,N_21424,N_20694);
xnor U25269 (N_25269,N_23397,N_22940);
nor U25270 (N_25270,N_22336,N_23028);
nor U25271 (N_25271,N_20053,N_20681);
nand U25272 (N_25272,N_20125,N_22897);
or U25273 (N_25273,N_24819,N_21471);
nor U25274 (N_25274,N_21805,N_24051);
and U25275 (N_25275,N_22047,N_21391);
and U25276 (N_25276,N_22396,N_22164);
nand U25277 (N_25277,N_24486,N_24641);
nor U25278 (N_25278,N_24327,N_22107);
xnor U25279 (N_25279,N_21314,N_24006);
nor U25280 (N_25280,N_23590,N_24204);
nor U25281 (N_25281,N_21968,N_22296);
and U25282 (N_25282,N_20065,N_21374);
or U25283 (N_25283,N_20099,N_21721);
nor U25284 (N_25284,N_21552,N_20088);
or U25285 (N_25285,N_24559,N_24941);
xnor U25286 (N_25286,N_21794,N_23244);
or U25287 (N_25287,N_20218,N_24737);
or U25288 (N_25288,N_21993,N_24678);
xnor U25289 (N_25289,N_23281,N_21483);
and U25290 (N_25290,N_24244,N_21516);
or U25291 (N_25291,N_20143,N_23496);
or U25292 (N_25292,N_22200,N_23990);
xor U25293 (N_25293,N_24376,N_20633);
nand U25294 (N_25294,N_21216,N_20614);
nor U25295 (N_25295,N_20187,N_22322);
and U25296 (N_25296,N_21179,N_22748);
xor U25297 (N_25297,N_22938,N_21936);
nand U25298 (N_25298,N_22162,N_22168);
or U25299 (N_25299,N_23979,N_22182);
and U25300 (N_25300,N_22899,N_22718);
and U25301 (N_25301,N_21836,N_20428);
nand U25302 (N_25302,N_20945,N_23888);
nor U25303 (N_25303,N_23994,N_20215);
nand U25304 (N_25304,N_22630,N_23418);
and U25305 (N_25305,N_21757,N_23312);
and U25306 (N_25306,N_24585,N_21013);
and U25307 (N_25307,N_22701,N_21418);
or U25308 (N_25308,N_22528,N_24090);
or U25309 (N_25309,N_24303,N_23406);
nand U25310 (N_25310,N_24625,N_21675);
nor U25311 (N_25311,N_24976,N_24261);
nand U25312 (N_25312,N_22564,N_23136);
xnor U25313 (N_25313,N_22395,N_24750);
xor U25314 (N_25314,N_22364,N_24163);
or U25315 (N_25315,N_20503,N_20095);
nor U25316 (N_25316,N_24477,N_20600);
nand U25317 (N_25317,N_21957,N_24755);
or U25318 (N_25318,N_22098,N_20931);
nand U25319 (N_25319,N_22130,N_24349);
nand U25320 (N_25320,N_24423,N_24606);
xnor U25321 (N_25321,N_23197,N_24548);
nand U25322 (N_25322,N_21044,N_21207);
nand U25323 (N_25323,N_22597,N_22099);
xnor U25324 (N_25324,N_20975,N_23680);
nand U25325 (N_25325,N_23113,N_20745);
nand U25326 (N_25326,N_20908,N_23258);
and U25327 (N_25327,N_24057,N_21456);
xor U25328 (N_25328,N_21199,N_22549);
xor U25329 (N_25329,N_24236,N_20801);
or U25330 (N_25330,N_20480,N_20500);
and U25331 (N_25331,N_21080,N_21297);
or U25332 (N_25332,N_24191,N_20635);
nor U25333 (N_25333,N_23052,N_21062);
nor U25334 (N_25334,N_23586,N_24114);
nand U25335 (N_25335,N_24852,N_23647);
or U25336 (N_25336,N_20696,N_20992);
nand U25337 (N_25337,N_21497,N_20557);
nand U25338 (N_25338,N_24010,N_22800);
and U25339 (N_25339,N_22127,N_21548);
and U25340 (N_25340,N_24790,N_20655);
nor U25341 (N_25341,N_24619,N_22613);
or U25342 (N_25342,N_22551,N_20160);
or U25343 (N_25343,N_20115,N_23524);
xnor U25344 (N_25344,N_22320,N_21858);
nand U25345 (N_25345,N_20332,N_22023);
xor U25346 (N_25346,N_22838,N_20008);
and U25347 (N_25347,N_23661,N_24088);
nand U25348 (N_25348,N_20789,N_23000);
nor U25349 (N_25349,N_23761,N_24751);
nor U25350 (N_25350,N_23641,N_21578);
nand U25351 (N_25351,N_20073,N_20615);
nor U25352 (N_25352,N_22446,N_23302);
nand U25353 (N_25353,N_24753,N_22913);
or U25354 (N_25354,N_24688,N_22223);
nor U25355 (N_25355,N_24353,N_21416);
nand U25356 (N_25356,N_24438,N_23949);
nor U25357 (N_25357,N_20108,N_20799);
xor U25358 (N_25358,N_23738,N_20274);
xnor U25359 (N_25359,N_23414,N_22739);
or U25360 (N_25360,N_20257,N_22066);
or U25361 (N_25361,N_23805,N_22215);
nand U25362 (N_25362,N_22562,N_24464);
nand U25363 (N_25363,N_20949,N_23353);
or U25364 (N_25364,N_20830,N_20198);
xor U25365 (N_25365,N_22619,N_23481);
or U25366 (N_25366,N_23860,N_20075);
xnor U25367 (N_25367,N_23616,N_23438);
nand U25368 (N_25368,N_20211,N_24009);
or U25369 (N_25369,N_20872,N_23168);
or U25370 (N_25370,N_21942,N_20416);
nand U25371 (N_25371,N_21295,N_21638);
and U25372 (N_25372,N_20995,N_24198);
nand U25373 (N_25373,N_21596,N_22219);
and U25374 (N_25374,N_20156,N_22628);
nand U25375 (N_25375,N_24254,N_24780);
and U25376 (N_25376,N_21346,N_24798);
nor U25377 (N_25377,N_21439,N_20756);
and U25378 (N_25378,N_20490,N_22852);
xnor U25379 (N_25379,N_23232,N_21754);
xnor U25380 (N_25380,N_23081,N_24858);
nor U25381 (N_25381,N_21806,N_21353);
xnor U25382 (N_25382,N_23732,N_23827);
or U25383 (N_25383,N_23362,N_23066);
xor U25384 (N_25384,N_24534,N_22374);
xnor U25385 (N_25385,N_20292,N_23400);
and U25386 (N_25386,N_20509,N_20403);
or U25387 (N_25387,N_22280,N_22439);
nand U25388 (N_25388,N_21656,N_23167);
nand U25389 (N_25389,N_20032,N_22775);
and U25390 (N_25390,N_20751,N_22357);
nand U25391 (N_25391,N_22242,N_22532);
and U25392 (N_25392,N_20545,N_24345);
xor U25393 (N_25393,N_23796,N_21154);
nor U25394 (N_25394,N_21141,N_24864);
nor U25395 (N_25395,N_20935,N_23340);
nand U25396 (N_25396,N_24495,N_23487);
xnor U25397 (N_25397,N_22173,N_20692);
nand U25398 (N_25398,N_21212,N_20802);
and U25399 (N_25399,N_23585,N_20339);
nor U25400 (N_25400,N_21434,N_21798);
nor U25401 (N_25401,N_21782,N_23018);
or U25402 (N_25402,N_24379,N_21234);
xor U25403 (N_25403,N_24517,N_22729);
or U25404 (N_25404,N_20163,N_23916);
xnor U25405 (N_25405,N_24672,N_24321);
xnor U25406 (N_25406,N_21073,N_21070);
or U25407 (N_25407,N_24985,N_23634);
and U25408 (N_25408,N_24137,N_24660);
nor U25409 (N_25409,N_20981,N_20015);
or U25410 (N_25410,N_21864,N_23513);
nand U25411 (N_25411,N_23404,N_24828);
and U25412 (N_25412,N_21290,N_21563);
and U25413 (N_25413,N_24966,N_24810);
or U25414 (N_25414,N_24061,N_24954);
nand U25415 (N_25415,N_20702,N_20045);
nor U25416 (N_25416,N_22033,N_24120);
and U25417 (N_25417,N_20805,N_24410);
or U25418 (N_25418,N_24425,N_21003);
nand U25419 (N_25419,N_21831,N_23746);
nor U25420 (N_25420,N_22041,N_24080);
xnor U25421 (N_25421,N_24107,N_20259);
nand U25422 (N_25422,N_20495,N_23076);
nor U25423 (N_25423,N_20854,N_21011);
and U25424 (N_25424,N_23812,N_23055);
nor U25425 (N_25425,N_21059,N_24822);
and U25426 (N_25426,N_21444,N_21408);
and U25427 (N_25427,N_22405,N_21838);
and U25428 (N_25428,N_24092,N_24350);
or U25429 (N_25429,N_20389,N_21760);
or U25430 (N_25430,N_21325,N_22150);
or U25431 (N_25431,N_20318,N_22125);
nand U25432 (N_25432,N_24617,N_21534);
or U25433 (N_25433,N_24492,N_20020);
or U25434 (N_25434,N_22398,N_23366);
xor U25435 (N_25435,N_21301,N_23533);
nor U25436 (N_25436,N_23007,N_23442);
and U25437 (N_25437,N_24825,N_24633);
and U25438 (N_25438,N_21849,N_20589);
nor U25439 (N_25439,N_24832,N_20474);
nor U25440 (N_25440,N_22693,N_21394);
xnor U25441 (N_25441,N_21572,N_23220);
xor U25442 (N_25442,N_22014,N_23420);
nor U25443 (N_25443,N_24885,N_23164);
xnor U25444 (N_25444,N_23683,N_20230);
nand U25445 (N_25445,N_24478,N_22914);
or U25446 (N_25446,N_24229,N_24547);
nor U25447 (N_25447,N_23650,N_22451);
nand U25448 (N_25448,N_23444,N_21025);
nor U25449 (N_25449,N_24184,N_20456);
xnor U25450 (N_25450,N_21998,N_20528);
or U25451 (N_25451,N_23690,N_21913);
nand U25452 (N_25452,N_24143,N_23032);
nand U25453 (N_25453,N_22520,N_24173);
and U25454 (N_25454,N_22524,N_21556);
xnor U25455 (N_25455,N_20682,N_22341);
xor U25456 (N_25456,N_20129,N_24449);
and U25457 (N_25457,N_24253,N_20086);
nand U25458 (N_25458,N_21986,N_22288);
nor U25459 (N_25459,N_20200,N_21963);
or U25460 (N_25460,N_20289,N_22746);
nor U25461 (N_25461,N_23515,N_23598);
xnor U25462 (N_25462,N_24367,N_20989);
and U25463 (N_25463,N_21294,N_20372);
and U25464 (N_25464,N_23327,N_23942);
or U25465 (N_25465,N_23096,N_23097);
nand U25466 (N_25466,N_24246,N_24497);
xor U25467 (N_25467,N_24243,N_22080);
and U25468 (N_25468,N_21054,N_21678);
nor U25469 (N_25469,N_22476,N_24030);
nor U25470 (N_25470,N_21200,N_20029);
nor U25471 (N_25471,N_20653,N_20990);
xor U25472 (N_25472,N_20321,N_23070);
or U25473 (N_25473,N_24490,N_24746);
or U25474 (N_25474,N_20406,N_23831);
nor U25475 (N_25475,N_24487,N_24050);
and U25476 (N_25476,N_20144,N_24935);
xnor U25477 (N_25477,N_20127,N_22067);
nor U25478 (N_25478,N_22928,N_24821);
or U25479 (N_25479,N_24709,N_24648);
nor U25480 (N_25480,N_21246,N_22292);
xor U25481 (N_25481,N_21012,N_24491);
nand U25482 (N_25482,N_21360,N_23031);
xnor U25483 (N_25483,N_20836,N_21226);
nor U25484 (N_25484,N_23820,N_21479);
and U25485 (N_25485,N_24473,N_22514);
nand U25486 (N_25486,N_24589,N_23088);
xnor U25487 (N_25487,N_21508,N_20699);
or U25488 (N_25488,N_22530,N_20806);
nor U25489 (N_25489,N_21862,N_20101);
xnor U25490 (N_25490,N_20356,N_22342);
nor U25491 (N_25491,N_23718,N_21669);
or U25492 (N_25492,N_23792,N_21897);
nor U25493 (N_25493,N_23768,N_20720);
nor U25494 (N_25494,N_23733,N_23504);
xnor U25495 (N_25495,N_20575,N_22629);
and U25496 (N_25496,N_24230,N_20934);
xor U25497 (N_25497,N_20443,N_22774);
nor U25498 (N_25498,N_24304,N_20735);
and U25499 (N_25499,N_21029,N_24631);
and U25500 (N_25500,N_21681,N_23806);
and U25501 (N_25501,N_23742,N_23307);
nand U25502 (N_25502,N_20306,N_23040);
nand U25503 (N_25503,N_23297,N_22021);
or U25504 (N_25504,N_20987,N_20791);
nand U25505 (N_25505,N_21352,N_22116);
and U25506 (N_25506,N_21110,N_23384);
or U25507 (N_25507,N_21075,N_23108);
xor U25508 (N_25508,N_22544,N_21001);
nor U25509 (N_25509,N_24567,N_21774);
nand U25510 (N_25510,N_24466,N_24505);
xor U25511 (N_25511,N_21755,N_21108);
and U25512 (N_25512,N_21538,N_21612);
and U25513 (N_25513,N_20656,N_21426);
nor U25514 (N_25514,N_24252,N_21589);
and U25515 (N_25515,N_22959,N_22790);
or U25516 (N_25516,N_22529,N_23027);
nand U25517 (N_25517,N_21987,N_20236);
and U25518 (N_25518,N_20905,N_22239);
nor U25519 (N_25519,N_23328,N_22979);
xnor U25520 (N_25520,N_21544,N_22848);
xnor U25521 (N_25521,N_22019,N_20649);
xnor U25522 (N_25522,N_22335,N_23983);
xor U25523 (N_25523,N_24900,N_21311);
and U25524 (N_25524,N_20524,N_23471);
nor U25525 (N_25525,N_23127,N_22244);
or U25526 (N_25526,N_24731,N_21240);
nor U25527 (N_25527,N_20859,N_23435);
xor U25528 (N_25528,N_24501,N_24296);
and U25529 (N_25529,N_20291,N_22220);
nand U25530 (N_25530,N_22347,N_20873);
xor U25531 (N_25531,N_22272,N_21153);
nand U25532 (N_25532,N_24005,N_21827);
or U25533 (N_25533,N_21308,N_20680);
or U25534 (N_25534,N_24738,N_20666);
xor U25535 (N_25535,N_23852,N_23440);
or U25536 (N_25536,N_22851,N_23632);
nand U25537 (N_25537,N_24012,N_21511);
and U25538 (N_25538,N_20952,N_21414);
and U25539 (N_25539,N_23053,N_20749);
or U25540 (N_25540,N_24078,N_24599);
nor U25541 (N_25541,N_24453,N_21017);
or U25542 (N_25542,N_24294,N_20753);
or U25543 (N_25543,N_24455,N_21350);
nand U25544 (N_25544,N_24338,N_24784);
nand U25545 (N_25545,N_22796,N_23130);
xnor U25546 (N_25546,N_22491,N_20227);
and U25547 (N_25547,N_20569,N_22961);
xnor U25548 (N_25548,N_22218,N_22875);
nor U25549 (N_25549,N_22068,N_24218);
nor U25550 (N_25550,N_20625,N_24662);
and U25551 (N_25551,N_22226,N_20328);
or U25552 (N_25552,N_22795,N_23180);
xnor U25553 (N_25553,N_21397,N_21061);
xor U25554 (N_25554,N_23213,N_21526);
nor U25555 (N_25555,N_24814,N_23646);
nand U25556 (N_25556,N_20973,N_23578);
nor U25557 (N_25557,N_22962,N_22146);
xor U25558 (N_25558,N_24195,N_24710);
nand U25559 (N_25559,N_21030,N_22557);
or U25560 (N_25560,N_21597,N_23422);
nand U25561 (N_25561,N_24552,N_20940);
nand U25562 (N_25562,N_20732,N_22927);
and U25563 (N_25563,N_22042,N_23041);
nor U25564 (N_25564,N_24874,N_24826);
xor U25565 (N_25565,N_20867,N_21887);
and U25566 (N_25566,N_21964,N_23763);
and U25567 (N_25567,N_22936,N_23266);
nor U25568 (N_25568,N_22606,N_20946);
nand U25569 (N_25569,N_24677,N_22075);
and U25570 (N_25570,N_22866,N_23467);
nor U25571 (N_25571,N_22004,N_21576);
or U25572 (N_25572,N_21546,N_21610);
or U25573 (N_25573,N_21109,N_21533);
or U25574 (N_25574,N_22589,N_23275);
xor U25575 (N_25575,N_22565,N_22723);
or U25576 (N_25576,N_20903,N_22752);
nor U25577 (N_25577,N_21615,N_20007);
or U25578 (N_25578,N_23341,N_21627);
nand U25579 (N_25579,N_24967,N_22279);
or U25580 (N_25580,N_22370,N_20433);
nor U25581 (N_25581,N_21351,N_23237);
nand U25582 (N_25582,N_24106,N_20576);
and U25583 (N_25583,N_20798,N_20149);
nor U25584 (N_25584,N_23446,N_21130);
xnor U25585 (N_25585,N_22863,N_24508);
and U25586 (N_25586,N_23645,N_23240);
xor U25587 (N_25587,N_22588,N_21103);
nand U25588 (N_25588,N_23896,N_24910);
or U25589 (N_25589,N_21818,N_24072);
nor U25590 (N_25590,N_22522,N_23263);
xnor U25591 (N_25591,N_23588,N_21005);
nor U25592 (N_25592,N_22463,N_23617);
or U25593 (N_25593,N_20438,N_20972);
nand U25594 (N_25594,N_20035,N_23739);
or U25595 (N_25595,N_23417,N_22028);
nor U25596 (N_25596,N_23901,N_22652);
nand U25597 (N_25597,N_20532,N_20084);
or U25598 (N_25598,N_24256,N_21489);
and U25599 (N_25599,N_24792,N_24771);
nand U25600 (N_25600,N_23625,N_24320);
xor U25601 (N_25601,N_23717,N_22368);
xor U25602 (N_25602,N_21366,N_22762);
nor U25603 (N_25603,N_21657,N_20254);
or U25604 (N_25604,N_23832,N_23978);
nand U25605 (N_25605,N_22660,N_22511);
xor U25606 (N_25606,N_21883,N_20892);
nand U25607 (N_25607,N_21795,N_20612);
xor U25608 (N_25608,N_21541,N_22999);
nand U25609 (N_25609,N_21796,N_23499);
nor U25610 (N_25610,N_22414,N_24866);
nand U25611 (N_25611,N_24377,N_21265);
xnor U25612 (N_25612,N_23840,N_23074);
nor U25613 (N_25613,N_20620,N_23841);
or U25614 (N_25614,N_24986,N_24014);
nand U25615 (N_25615,N_23115,N_20918);
nor U25616 (N_25616,N_21604,N_20790);
nand U25617 (N_25617,N_24445,N_24211);
nor U25618 (N_25618,N_20175,N_20712);
and U25619 (N_25619,N_23170,N_22073);
nor U25620 (N_25620,N_22889,N_24217);
nor U25621 (N_25621,N_22431,N_24293);
or U25622 (N_25622,N_22976,N_23001);
nor U25623 (N_25623,N_23503,N_23316);
xnor U25624 (N_25624,N_24479,N_22907);
or U25625 (N_25625,N_24469,N_22184);
nand U25626 (N_25626,N_23799,N_24806);
and U25627 (N_25627,N_24430,N_23664);
nand U25628 (N_25628,N_24194,N_21558);
xor U25629 (N_25629,N_21867,N_22382);
nand U25630 (N_25630,N_21322,N_20937);
or U25631 (N_25631,N_23039,N_24216);
nand U25632 (N_25632,N_22794,N_23162);
xnor U25633 (N_25633,N_24594,N_20808);
xnor U25634 (N_25634,N_20130,N_21879);
xnor U25635 (N_25635,N_21688,N_23461);
xnor U25636 (N_25636,N_22815,N_20708);
or U25637 (N_25637,N_22203,N_20173);
or U25638 (N_25638,N_20240,N_22303);
nor U25639 (N_25639,N_23769,N_23904);
nor U25640 (N_25640,N_24932,N_23251);
nor U25641 (N_25641,N_21031,N_23009);
or U25642 (N_25642,N_21250,N_23615);
or U25643 (N_25643,N_20251,N_20909);
and U25644 (N_25644,N_24701,N_20445);
nor U25645 (N_25645,N_24428,N_24992);
xor U25646 (N_25646,N_24521,N_24322);
and U25647 (N_25647,N_24708,N_23842);
or U25648 (N_25648,N_24982,N_22945);
nor U25649 (N_25649,N_22950,N_24189);
or U25650 (N_25650,N_23553,N_24730);
nand U25651 (N_25651,N_22952,N_24393);
nand U25652 (N_25652,N_24978,N_21211);
xnor U25653 (N_25653,N_23061,N_24666);
nor U25654 (N_25654,N_23694,N_23546);
xnor U25655 (N_25655,N_23721,N_21370);
nor U25656 (N_25656,N_24025,N_21717);
nor U25657 (N_25657,N_23268,N_21724);
xnor U25658 (N_25658,N_22951,N_23740);
nand U25659 (N_25659,N_24209,N_22252);
nand U25660 (N_25660,N_20938,N_20267);
xor U25661 (N_25661,N_21187,N_24609);
nor U25662 (N_25662,N_20922,N_23766);
xnor U25663 (N_25663,N_23687,N_20391);
nand U25664 (N_25664,N_23505,N_22400);
or U25665 (N_25665,N_24528,N_24671);
nor U25666 (N_25666,N_20838,N_23029);
nand U25667 (N_25667,N_22160,N_22269);
and U25668 (N_25668,N_20993,N_22941);
nor U25669 (N_25669,N_23368,N_21980);
xnor U25670 (N_25670,N_22380,N_24754);
nor U25671 (N_25671,N_23421,N_20730);
and U25672 (N_25672,N_24550,N_20630);
nor U25673 (N_25673,N_23811,N_23092);
or U25674 (N_25674,N_24152,N_20158);
xnor U25675 (N_25675,N_24945,N_23752);
nor U25676 (N_25676,N_23190,N_23325);
and U25677 (N_25677,N_24676,N_22770);
nor U25678 (N_25678,N_20661,N_24968);
xnor U25679 (N_25679,N_22764,N_23239);
nor U25680 (N_25680,N_20288,N_24933);
or U25681 (N_25681,N_23046,N_21107);
xnor U25682 (N_25682,N_22459,N_21067);
and U25683 (N_25683,N_23600,N_21950);
nand U25684 (N_25684,N_21555,N_20462);
or U25685 (N_25685,N_22783,N_22311);
xor U25686 (N_25686,N_20104,N_21072);
nand U25687 (N_25687,N_20022,N_23571);
and U25688 (N_25688,N_23727,N_22181);
nor U25689 (N_25689,N_20748,N_20499);
xor U25690 (N_25690,N_20734,N_23110);
and U25691 (N_25691,N_22114,N_22444);
xor U25692 (N_25692,N_23427,N_22108);
nand U25693 (N_25693,N_22328,N_24956);
and U25694 (N_25694,N_23620,N_24908);
or U25695 (N_25695,N_20025,N_23309);
nor U25696 (N_25696,N_23866,N_24392);
or U25697 (N_25697,N_23356,N_22186);
nand U25698 (N_25698,N_23855,N_22898);
and U25699 (N_25699,N_24245,N_23914);
or U25700 (N_25700,N_20224,N_20917);
nand U25701 (N_25701,N_24314,N_21565);
xor U25702 (N_25702,N_24155,N_22049);
xnor U25703 (N_25703,N_24186,N_21522);
xnor U25704 (N_25704,N_21874,N_22170);
and U25705 (N_25705,N_24632,N_24974);
nor U25706 (N_25706,N_22853,N_20647);
xnor U25707 (N_25707,N_24846,N_22654);
or U25708 (N_25708,N_21160,N_23688);
nand U25709 (N_25709,N_21047,N_24752);
and U25710 (N_25710,N_20048,N_21684);
and U25711 (N_25711,N_23393,N_21892);
nor U25712 (N_25712,N_24569,N_23657);
or U25713 (N_25713,N_22634,N_21045);
xor U25714 (N_25714,N_24139,N_23019);
and U25715 (N_25715,N_24953,N_21643);
or U25716 (N_25716,N_24259,N_23824);
nor U25717 (N_25717,N_20737,N_21307);
nor U25718 (N_25718,N_22227,N_23541);
and U25719 (N_25719,N_24474,N_24668);
xor U25720 (N_25720,N_20235,N_24979);
and U25721 (N_25721,N_23743,N_23201);
and U25722 (N_25722,N_21310,N_24786);
nor U25723 (N_25723,N_22471,N_23969);
xor U25724 (N_25724,N_20269,N_22205);
nor U25725 (N_25725,N_24450,N_23477);
nand U25726 (N_25726,N_23095,N_21495);
or U25727 (N_25727,N_20252,N_22707);
and U25728 (N_25728,N_22636,N_22493);
nor U25729 (N_25729,N_20465,N_23780);
nand U25730 (N_25730,N_24459,N_23269);
nand U25731 (N_25731,N_21734,N_22309);
xor U25732 (N_25732,N_23454,N_21654);
nor U25733 (N_25733,N_22176,N_21911);
xor U25734 (N_25734,N_21111,N_23638);
or U25735 (N_25735,N_24812,N_21921);
nand U25736 (N_25736,N_23975,N_23488);
nor U25737 (N_25737,N_24356,N_21959);
nand U25738 (N_25738,N_21997,N_20494);
or U25739 (N_25739,N_20701,N_23548);
xnor U25740 (N_25740,N_20824,N_23593);
nor U25741 (N_25741,N_20497,N_22990);
and U25742 (N_25742,N_22657,N_22809);
nor U25743 (N_25743,N_20212,N_24694);
xnor U25744 (N_25744,N_22572,N_22010);
and U25745 (N_25745,N_20742,N_21402);
or U25746 (N_25746,N_20595,N_24297);
xor U25747 (N_25747,N_21362,N_24718);
nand U25748 (N_25748,N_22683,N_21140);
nand U25749 (N_25749,N_23893,N_23289);
nand U25750 (N_25750,N_21881,N_23428);
and U25751 (N_25751,N_22029,N_22351);
and U25752 (N_25752,N_21163,N_21752);
xnor U25753 (N_25753,N_22418,N_22975);
nor U25754 (N_25754,N_23217,N_24456);
or U25755 (N_25755,N_21592,N_22877);
or U25756 (N_25756,N_23253,N_23903);
nor U25757 (N_25757,N_22541,N_22330);
xnor U25758 (N_25758,N_22273,N_20261);
nand U25759 (N_25759,N_20276,N_23456);
and U25760 (N_25760,N_20740,N_20713);
and U25761 (N_25761,N_22786,N_24315);
xnor U25762 (N_25762,N_20688,N_21761);
and U25763 (N_25763,N_21616,N_23791);
or U25764 (N_25764,N_24611,N_23944);
xnor U25765 (N_25765,N_24948,N_23998);
and U25766 (N_25766,N_21443,N_23556);
nand U25767 (N_25767,N_22542,N_24965);
or U25768 (N_25768,N_21812,N_20283);
nor U25769 (N_25769,N_24031,N_21316);
nand U25770 (N_25770,N_21217,N_23807);
or U25771 (N_25771,N_24796,N_24561);
and U25772 (N_25772,N_22012,N_22973);
and U25773 (N_25773,N_21991,N_22697);
nand U25774 (N_25774,N_21377,N_20984);
nand U25775 (N_25775,N_22502,N_23773);
and U25776 (N_25776,N_22401,N_24630);
and U25777 (N_25777,N_24726,N_24568);
nand U25778 (N_25778,N_21117,N_22934);
xor U25779 (N_25779,N_20210,N_24138);
or U25780 (N_25780,N_21633,N_22953);
and U25781 (N_25781,N_21068,N_20794);
nor U25782 (N_25782,N_23580,N_24650);
nor U25783 (N_25783,N_20691,N_22429);
nor U25784 (N_25784,N_21467,N_24439);
and U25785 (N_25785,N_22399,N_20362);
nor U25786 (N_25786,N_21847,N_24816);
xor U25787 (N_25787,N_21848,N_23892);
nor U25788 (N_25788,N_20479,N_24013);
and U25789 (N_25789,N_21457,N_24837);
or U25790 (N_25790,N_21898,N_21136);
and U25791 (N_25791,N_21791,N_21148);
and U25792 (N_25792,N_22050,N_22434);
nor U25793 (N_25793,N_24860,N_24295);
or U25794 (N_25794,N_21540,N_23517);
or U25795 (N_25795,N_21766,N_21122);
xor U25796 (N_25796,N_20857,N_20120);
xnor U25797 (N_25797,N_21732,N_24060);
xor U25798 (N_25798,N_20602,N_21579);
or U25799 (N_25799,N_24054,N_24889);
and U25800 (N_25800,N_22002,N_20832);
or U25801 (N_25801,N_22798,N_22747);
nor U25802 (N_25802,N_21204,N_21871);
nor U25803 (N_25803,N_24422,N_22131);
and U25804 (N_25804,N_23476,N_21464);
nand U25805 (N_25805,N_24178,N_20059);
xnor U25806 (N_25806,N_20958,N_23071);
nand U25807 (N_25807,N_24896,N_22733);
and U25808 (N_25808,N_23260,N_24993);
and U25809 (N_25809,N_22120,N_21388);
nor U25810 (N_25810,N_21719,N_22110);
xor U25811 (N_25811,N_24570,N_22171);
or U25812 (N_25812,N_22674,N_24546);
or U25813 (N_25813,N_23150,N_20517);
nand U25814 (N_25814,N_24716,N_22728);
nand U25815 (N_25815,N_21803,N_22193);
nand U25816 (N_25816,N_23484,N_21744);
nor U25817 (N_25817,N_20953,N_23051);
xor U25818 (N_25818,N_22317,N_23775);
or U25819 (N_25819,N_23584,N_23333);
nand U25820 (N_25820,N_22993,N_21334);
nand U25821 (N_25821,N_21532,N_22621);
nand U25822 (N_25822,N_21241,N_21168);
nand U25823 (N_25823,N_22699,N_21876);
and U25824 (N_25824,N_23087,N_21707);
nor U25825 (N_25825,N_24272,N_20641);
xnor U25826 (N_25826,N_20484,N_23283);
xnor U25827 (N_25827,N_21326,N_21629);
nor U25828 (N_25828,N_20453,N_24440);
nor U25829 (N_25829,N_20178,N_21662);
nand U25830 (N_25830,N_22937,N_22916);
or U25831 (N_25831,N_23555,N_20349);
nand U25832 (N_25832,N_23433,N_22655);
xor U25833 (N_25833,N_23753,N_20906);
nand U25834 (N_25834,N_23466,N_24647);
nand U25835 (N_25835,N_24043,N_21819);
nand U25836 (N_25836,N_20468,N_20420);
or U25837 (N_25837,N_23587,N_20353);
nor U25838 (N_25838,N_24605,N_20768);
and U25839 (N_25839,N_22704,N_20788);
xnor U25840 (N_25840,N_23146,N_20616);
nand U25841 (N_25841,N_22037,N_20205);
nand U25842 (N_25842,N_21961,N_20082);
xor U25843 (N_25843,N_20247,N_21910);
xnor U25844 (N_25844,N_20331,N_23659);
nand U25845 (N_25845,N_23250,N_20385);
or U25846 (N_25846,N_24799,N_21981);
and U25847 (N_25847,N_24856,N_24918);
or U25848 (N_25848,N_24618,N_20746);
or U25849 (N_25849,N_21008,N_21573);
or U25850 (N_25850,N_21587,N_21469);
xor U25851 (N_25851,N_24717,N_22307);
or U25852 (N_25852,N_20599,N_21133);
xor U25853 (N_25853,N_24575,N_21975);
nand U25854 (N_25854,N_21312,N_23378);
or U25855 (N_25855,N_23202,N_23707);
nor U25856 (N_25856,N_22388,N_21281);
nand U25857 (N_25857,N_22440,N_23651);
and U25858 (N_25858,N_23720,N_20054);
nor U25859 (N_25859,N_21296,N_23196);
and U25860 (N_25860,N_21677,N_23434);
xnor U25861 (N_25861,N_20508,N_20111);
or U25862 (N_25862,N_20793,N_21787);
and U25863 (N_25863,N_22972,N_23141);
xor U25864 (N_25864,N_20695,N_21948);
xnor U25865 (N_25865,N_23883,N_22126);
xor U25866 (N_25866,N_24598,N_24227);
nand U25867 (N_25867,N_21660,N_23633);
xor U25868 (N_25868,N_21303,N_21355);
or U25869 (N_25869,N_22540,N_24159);
and U25870 (N_25870,N_23062,N_22873);
or U25871 (N_25871,N_23043,N_20145);
nand U25872 (N_25872,N_22751,N_22624);
and U25873 (N_25873,N_24026,N_21530);
and U25874 (N_25874,N_24463,N_23212);
or U25875 (N_25875,N_20436,N_20238);
nand U25876 (N_25876,N_22460,N_21494);
nand U25877 (N_25877,N_23767,N_20529);
or U25878 (N_25878,N_22112,N_20967);
nand U25879 (N_25879,N_21057,N_24772);
nor U25880 (N_25880,N_22732,N_22886);
xor U25881 (N_25881,N_21266,N_23623);
or U25882 (N_25882,N_22692,N_24135);
nor U25883 (N_25883,N_23781,N_23951);
nor U25884 (N_25884,N_24757,N_20764);
and U25885 (N_25885,N_23176,N_20094);
nand U25886 (N_25886,N_21028,N_23693);
or U25887 (N_25887,N_23826,N_22837);
nor U25888 (N_25888,N_22882,N_23570);
or U25889 (N_25889,N_20919,N_21480);
nand U25890 (N_25890,N_21041,N_20566);
nand U25891 (N_25891,N_24628,N_24728);
or U25892 (N_25892,N_23107,N_22537);
or U25893 (N_25893,N_24781,N_23547);
nor U25894 (N_25894,N_21988,N_21230);
xor U25895 (N_25895,N_24721,N_20606);
nand U25896 (N_25896,N_20844,N_22915);
xor U25897 (N_25897,N_20693,N_22711);
or U25898 (N_25898,N_22604,N_21493);
xor U25899 (N_25899,N_21321,N_23945);
nor U25900 (N_25900,N_24592,N_23177);
xnor U25901 (N_25901,N_21535,N_20270);
xor U25902 (N_25902,N_23719,N_23509);
nor U25903 (N_25903,N_23785,N_22772);
nor U25904 (N_25904,N_23277,N_23211);
nor U25905 (N_25905,N_21120,N_24048);
nand U25906 (N_25906,N_23411,N_20133);
or U25907 (N_25907,N_21809,N_20856);
nor U25908 (N_25908,N_20074,N_23292);
nor U25909 (N_25909,N_20369,N_21915);
nand U25910 (N_25910,N_20667,N_23195);
or U25911 (N_25911,N_24800,N_22416);
xnor U25912 (N_25912,N_22921,N_21227);
nand U25913 (N_25913,N_20155,N_24842);
or U25914 (N_25914,N_23249,N_24762);
or U25915 (N_25915,N_21720,N_24680);
and U25916 (N_25916,N_24084,N_20923);
xor U25917 (N_25917,N_23574,N_20869);
or U25918 (N_25918,N_22138,N_21422);
nor U25919 (N_25919,N_23507,N_20229);
and U25920 (N_25920,N_21247,N_22981);
xnor U25921 (N_25921,N_21252,N_23198);
xor U25922 (N_25922,N_21248,N_24600);
nand U25923 (N_25923,N_20049,N_20570);
and U25924 (N_25924,N_23126,N_20979);
nor U25925 (N_25925,N_20319,N_21463);
and U25926 (N_25926,N_22237,N_24333);
nor U25927 (N_25927,N_24242,N_22024);
or U25928 (N_25928,N_24262,N_24939);
xor U25929 (N_25929,N_22834,N_20016);
or U25930 (N_25930,N_20466,N_24251);
or U25931 (N_25931,N_23489,N_23012);
nand U25932 (N_25932,N_20638,N_20329);
xor U25933 (N_25933,N_21021,N_23301);
and U25934 (N_25934,N_23676,N_21839);
or U25935 (N_25935,N_21725,N_21613);
and U25936 (N_25936,N_21093,N_21801);
and U25937 (N_25937,N_22879,N_23798);
nand U25938 (N_25938,N_23858,N_22721);
or U25939 (N_25939,N_22991,N_23879);
and U25940 (N_25940,N_20928,N_24529);
nand U25941 (N_25941,N_22688,N_22383);
and U25942 (N_25942,N_24880,N_22513);
xnor U25943 (N_25943,N_22820,N_21659);
nor U25944 (N_25944,N_21764,N_24745);
nor U25945 (N_25945,N_22142,N_20226);
xnor U25946 (N_25946,N_21515,N_22649);
and U25947 (N_25947,N_22466,N_21636);
or U25948 (N_25948,N_23145,N_23997);
nor U25949 (N_25949,N_23098,N_22813);
nand U25950 (N_25950,N_21663,N_20439);
nor U25951 (N_25951,N_21846,N_24336);
xor U25952 (N_25952,N_24836,N_24950);
nand U25953 (N_25953,N_20816,N_20624);
nor U25954 (N_25954,N_20716,N_22187);
nand U25955 (N_25955,N_24446,N_20469);
xnor U25956 (N_25956,N_24670,N_21441);
and U25957 (N_25957,N_21802,N_23669);
nand U25958 (N_25958,N_24622,N_23345);
xor U25959 (N_25959,N_20220,N_20883);
nor U25960 (N_25960,N_22935,N_24162);
nand U25961 (N_25961,N_23613,N_21710);
or U25962 (N_25962,N_24179,N_24140);
nand U25963 (N_25963,N_22982,N_22705);
and U25964 (N_25964,N_24201,N_21445);
nand U25965 (N_25965,N_23988,N_21648);
and U25966 (N_25966,N_23643,N_24123);
nand U25967 (N_25967,N_21896,N_20762);
and U25968 (N_25968,N_20519,N_24372);
and U25969 (N_25969,N_24934,N_21239);
or U25970 (N_25970,N_23464,N_20305);
xor U25971 (N_25971,N_22483,N_24615);
and U25972 (N_25972,N_24210,N_24307);
nor U25973 (N_25973,N_22512,N_20309);
or U25974 (N_25974,N_23782,N_24614);
xnor U25975 (N_25975,N_21191,N_24037);
or U25976 (N_25976,N_24240,N_24947);
nand U25977 (N_25977,N_22056,N_20840);
xnor U25978 (N_25978,N_23100,N_22251);
nor U25979 (N_25979,N_24185,N_23216);
xnor U25980 (N_25980,N_22811,N_21451);
and U25981 (N_25981,N_20902,N_22575);
or U25982 (N_25982,N_21115,N_24074);
xor U25983 (N_25983,N_20214,N_21484);
or U25984 (N_25984,N_24557,N_22609);
or U25985 (N_25985,N_20248,N_24224);
or U25986 (N_25986,N_22128,N_20607);
nor U25987 (N_25987,N_21953,N_20755);
nor U25988 (N_25988,N_20412,N_23538);
xor U25989 (N_25989,N_22826,N_24167);
xor U25990 (N_25990,N_22180,N_24095);
nand U25991 (N_25991,N_22261,N_23965);
and U25992 (N_25992,N_24951,N_20631);
nor U25993 (N_25993,N_20231,N_22420);
and U25994 (N_25994,N_21861,N_21996);
nand U25995 (N_25995,N_24878,N_20136);
nor U25996 (N_25996,N_23534,N_24997);
or U25997 (N_25997,N_20431,N_23304);
xor U25998 (N_25998,N_24895,N_22327);
or U25999 (N_25999,N_22777,N_23394);
nand U26000 (N_26000,N_22878,N_22792);
nor U26001 (N_26001,N_20165,N_24983);
nor U26002 (N_26002,N_22858,N_22498);
or U26003 (N_26003,N_20689,N_20287);
or U26004 (N_26004,N_22409,N_20835);
nor U26005 (N_26005,N_22246,N_23640);
nand U26006 (N_26006,N_24499,N_22521);
or U26007 (N_26007,N_24973,N_22298);
nor U26008 (N_26008,N_20584,N_23188);
or U26009 (N_26009,N_24586,N_20042);
nor U26010 (N_26010,N_23219,N_22964);
xor U26011 (N_26011,N_20450,N_21349);
nand U26012 (N_26012,N_24540,N_24341);
and U26013 (N_26013,N_24972,N_24269);
and U26014 (N_26014,N_21621,N_23940);
or U26015 (N_26015,N_21336,N_24034);
nand U26016 (N_26016,N_23478,N_23848);
nor U26017 (N_26017,N_24988,N_22441);
and U26018 (N_26018,N_22422,N_21192);
or U26019 (N_26019,N_24995,N_20930);
nor U26020 (N_26020,N_24990,N_22806);
or U26021 (N_26021,N_21421,N_20921);
and U26022 (N_26022,N_21689,N_20915);
nand U26023 (N_26023,N_23044,N_20581);
xor U26024 (N_26024,N_23474,N_22197);
nand U26025 (N_26025,N_24231,N_24335);
nand U26026 (N_26026,N_20410,N_20322);
nor U26027 (N_26027,N_24719,N_22750);
xor U26028 (N_26028,N_23453,N_22048);
or U26029 (N_26029,N_21275,N_23875);
and U26030 (N_26030,N_23528,N_24378);
or U26031 (N_26031,N_22217,N_22230);
nor U26032 (N_26032,N_21169,N_23984);
nand U26033 (N_26033,N_24213,N_21427);
nand U26034 (N_26034,N_21929,N_21091);
and U26035 (N_26035,N_21475,N_24729);
nand U26036 (N_26036,N_21219,N_24181);
or U26037 (N_26037,N_20551,N_24018);
nor U26038 (N_26038,N_22316,N_20070);
nand U26039 (N_26039,N_22359,N_21817);
xnor U26040 (N_26040,N_22829,N_24805);
or U26041 (N_26041,N_21195,N_24593);
nor U26042 (N_26042,N_21285,N_20683);
nor U26043 (N_26043,N_21300,N_22034);
nand U26044 (N_26044,N_22923,N_22695);
nand U26045 (N_26045,N_23639,N_24279);
and U26046 (N_26046,N_24725,N_22472);
nand U26047 (N_26047,N_22759,N_20715);
and U26048 (N_26048,N_24916,N_21264);
xnor U26049 (N_26049,N_22871,N_22717);
or U26050 (N_26050,N_20482,N_23022);
xnor U26051 (N_26051,N_23861,N_24020);
and U26052 (N_26052,N_22862,N_20081);
nand U26053 (N_26053,N_23731,N_23728);
and U26054 (N_26054,N_21591,N_23120);
nand U26055 (N_26055,N_21837,N_23987);
and U26056 (N_26056,N_22287,N_21347);
and U26057 (N_26057,N_20448,N_23329);
nor U26058 (N_26058,N_22648,N_24145);
nand U26059 (N_26059,N_22488,N_22553);
or U26060 (N_26060,N_24112,N_22231);
nand U26061 (N_26061,N_22967,N_23243);
xor U26062 (N_26062,N_20345,N_22306);
nor U26063 (N_26063,N_20463,N_24404);
or U26064 (N_26064,N_20541,N_23498);
nor U26065 (N_26065,N_21381,N_20021);
nor U26066 (N_26066,N_22841,N_24961);
or U26067 (N_26067,N_24288,N_21504);
and U26068 (N_26068,N_21271,N_23788);
xnor U26069 (N_26069,N_22458,N_24371);
or U26070 (N_26070,N_23724,N_21699);
xnor U26071 (N_26071,N_23786,N_23475);
and U26072 (N_26072,N_22000,N_21972);
nor U26073 (N_26073,N_24292,N_22464);
or U26074 (N_26074,N_22070,N_21951);
nand U26075 (N_26075,N_20034,N_23736);
xor U26076 (N_26076,N_20895,N_22534);
nor U26077 (N_26077,N_22054,N_23342);
and U26078 (N_26078,N_24704,N_20409);
or U26079 (N_26079,N_23252,N_23315);
nand U26080 (N_26080,N_23321,N_22278);
nand U26081 (N_26081,N_21777,N_20167);
and U26082 (N_26082,N_20507,N_23054);
xnor U26083 (N_26083,N_21748,N_20344);
and U26084 (N_26084,N_20171,N_20604);
or U26085 (N_26085,N_20787,N_23236);
or U26086 (N_26086,N_21243,N_24840);
nand U26087 (N_26087,N_24070,N_20534);
or U26088 (N_26088,N_24028,N_21505);
nand U26089 (N_26089,N_22901,N_23770);
xor U26090 (N_26090,N_20148,N_21545);
or U26091 (N_26091,N_24693,N_24309);
or U26092 (N_26092,N_20323,N_23270);
xnor U26093 (N_26093,N_22009,N_22266);
or U26094 (N_26094,N_20676,N_21703);
nor U26095 (N_26095,N_23809,N_24323);
nand U26096 (N_26096,N_23229,N_24019);
and U26097 (N_26097,N_23572,N_21413);
xnor U26098 (N_26098,N_24921,N_20677);
and U26099 (N_26099,N_23460,N_22397);
or U26100 (N_26100,N_20812,N_22808);
and U26101 (N_26101,N_21392,N_21679);
or U26102 (N_26102,N_22633,N_22424);
and U26103 (N_26103,N_24829,N_20897);
xor U26104 (N_26104,N_24642,N_21607);
or U26105 (N_26105,N_22202,N_22555);
or U26106 (N_26106,N_20626,N_24405);
nor U26107 (N_26107,N_23838,N_23847);
nand U26108 (N_26108,N_22373,N_23016);
nor U26109 (N_26109,N_20804,N_24354);
xor U26110 (N_26110,N_21834,N_24969);
or U26111 (N_26111,N_21020,N_23545);
or U26112 (N_26112,N_24749,N_22605);
nor U26113 (N_26113,N_20738,N_20068);
nor U26114 (N_26114,N_23605,N_21279);
nand U26115 (N_26115,N_21517,N_23759);
and U26116 (N_26116,N_21693,N_22281);
or U26117 (N_26117,N_22722,N_24306);
xor U26118 (N_26118,N_23116,N_24087);
xnor U26119 (N_26119,N_24283,N_24412);
nand U26120 (N_26120,N_23856,N_21932);
nand U26121 (N_26121,N_24461,N_24536);
or U26122 (N_26122,N_21649,N_21423);
nand U26123 (N_26123,N_23629,N_20157);
nand U26124 (N_26124,N_23377,N_21197);
and U26125 (N_26125,N_21539,N_24504);
nand U26126 (N_26126,N_24029,N_24919);
or U26127 (N_26127,N_21973,N_20669);
or U26128 (N_26128,N_21568,N_24226);
nand U26129 (N_26129,N_22500,N_20803);
or U26130 (N_26130,N_22869,N_21822);
nor U26131 (N_26131,N_24419,N_20382);
nor U26132 (N_26132,N_20262,N_20404);
nor U26133 (N_26133,N_23200,N_23050);
xnor U26134 (N_26134,N_24284,N_24901);
nand U26135 (N_26135,N_22855,N_22159);
and U26136 (N_26136,N_20121,N_22381);
and U26137 (N_26137,N_23678,N_21338);
xnor U26138 (N_26138,N_24624,N_23873);
nor U26139 (N_26139,N_23355,N_23182);
nand U26140 (N_26140,N_21024,N_23109);
nor U26141 (N_26141,N_21694,N_20326);
nand U26142 (N_26142,N_20761,N_23194);
nor U26143 (N_26143,N_23187,N_21967);
or U26144 (N_26144,N_24416,N_23462);
nand U26145 (N_26145,N_20538,N_23501);
nor U26146 (N_26146,N_23402,N_20177);
xnor U26147 (N_26147,N_22426,N_24520);
nor U26148 (N_26148,N_21899,N_23159);
and U26149 (N_26149,N_24475,N_23458);
or U26150 (N_26150,N_21431,N_24937);
and U26151 (N_26151,N_22743,N_22145);
and U26152 (N_26152,N_20554,N_22669);
xnor U26153 (N_26153,N_24300,N_24912);
nor U26154 (N_26154,N_20286,N_23014);
nor U26155 (N_26155,N_20487,N_24268);
xor U26156 (N_26156,N_23204,N_24957);
nor U26157 (N_26157,N_21023,N_23758);
nor U26158 (N_26158,N_24221,N_21697);
xor U26159 (N_26159,N_21984,N_23452);
nor U26160 (N_26160,N_24365,N_20330);
and U26161 (N_26161,N_23549,N_20169);
nor U26162 (N_26162,N_20726,N_23133);
and U26163 (N_26163,N_22207,N_22484);
or U26164 (N_26164,N_20038,N_20057);
nand U26165 (N_26165,N_24131,N_23712);
nor U26166 (N_26166,N_21570,N_21466);
xnor U26167 (N_26167,N_21875,N_21358);
or U26168 (N_26168,N_20013,N_21448);
nor U26169 (N_26169,N_24266,N_20228);
xor U26170 (N_26170,N_22527,N_23047);
nor U26171 (N_26171,N_20357,N_22253);
xor U26172 (N_26172,N_24734,N_22523);
nand U26173 (N_26173,N_23024,N_24496);
nor U26174 (N_26174,N_24571,N_21156);
nand U26175 (N_26175,N_20033,N_23181);
and U26176 (N_26176,N_21634,N_23711);
nor U26177 (N_26177,N_24576,N_20272);
nor U26178 (N_26178,N_22504,N_21118);
and U26179 (N_26179,N_24702,N_23535);
xnor U26180 (N_26180,N_22662,N_22773);
and U26181 (N_26181,N_22229,N_21704);
xnor U26182 (N_26182,N_21090,N_24398);
and U26183 (N_26183,N_22590,N_20342);
nand U26184 (N_26184,N_23974,N_21873);
nor U26185 (N_26185,N_22731,N_24241);
nand U26186 (N_26186,N_22233,N_21753);
and U26187 (N_26187,N_23057,N_24193);
xor U26188 (N_26188,N_20100,N_20377);
xor U26189 (N_26189,N_20293,N_20152);
xnor U26190 (N_26190,N_23674,N_21924);
xor U26191 (N_26191,N_22005,N_24219);
xor U26192 (N_26192,N_23286,N_21123);
xnor U26193 (N_26193,N_24281,N_24691);
nand U26194 (N_26194,N_23178,N_20018);
nor U26195 (N_26195,N_22078,N_21600);
nand U26196 (N_26196,N_24920,N_24363);
nor U26197 (N_26197,N_23439,N_21158);
nor U26198 (N_26198,N_22515,N_20939);
and U26199 (N_26199,N_24483,N_23124);
xnor U26200 (N_26200,N_20381,N_23063);
and U26201 (N_26201,N_22228,N_22206);
or U26202 (N_26202,N_24513,N_23564);
and U26203 (N_26203,N_23948,N_20168);
xor U26204 (N_26204,N_21651,N_24017);
and U26205 (N_26205,N_24059,N_24905);
nor U26206 (N_26206,N_23502,N_22581);
nand U26207 (N_26207,N_21173,N_22580);
and U26208 (N_26208,N_22064,N_24841);
and U26209 (N_26209,N_21528,N_23210);
nand U26210 (N_26210,N_20673,N_21776);
nor U26211 (N_26211,N_24498,N_22912);
and U26212 (N_26212,N_24938,N_24553);
and U26213 (N_26213,N_21293,N_23231);
xnor U26214 (N_26214,N_21941,N_22831);
and U26215 (N_26215,N_24192,N_23702);
and U26216 (N_26216,N_24773,N_22641);
or U26217 (N_26217,N_23310,N_24509);
nand U26218 (N_26218,N_20134,N_21785);
and U26219 (N_26219,N_24675,N_21344);
and U26220 (N_26220,N_20496,N_22823);
nand U26221 (N_26221,N_20562,N_21982);
nor U26222 (N_26222,N_21965,N_21905);
nor U26223 (N_26223,N_20629,N_20046);
or U26224 (N_26224,N_22734,N_21149);
xor U26225 (N_26225,N_21486,N_23403);
xor U26226 (N_26226,N_22353,N_24604);
nand U26227 (N_26227,N_23950,N_22030);
nand U26228 (N_26228,N_23280,N_24748);
or U26229 (N_26229,N_23784,N_20550);
nor U26230 (N_26230,N_22665,N_23876);
or U26231 (N_26231,N_22337,N_21577);
xnor U26232 (N_26232,N_21387,N_24989);
nor U26233 (N_26233,N_23846,N_24387);
xnor U26234 (N_26234,N_23143,N_24358);
and U26235 (N_26235,N_20885,N_24696);
or U26236 (N_26236,N_20191,N_24330);
xor U26237 (N_26237,N_20829,N_21010);
nand U26238 (N_26238,N_21702,N_22832);
nor U26239 (N_26239,N_23491,N_23675);
or U26240 (N_26240,N_21903,N_21139);
or U26241 (N_26241,N_20525,N_23673);
or U26242 (N_26242,N_24724,N_20437);
and U26243 (N_26243,N_24124,N_23299);
or U26244 (N_26244,N_23392,N_21931);
or U26245 (N_26245,N_24831,N_22039);
or U26246 (N_26246,N_21599,N_20780);
xor U26247 (N_26247,N_22082,N_23272);
nand U26248 (N_26248,N_24402,N_23049);
and U26249 (N_26249,N_23630,N_23305);
or U26250 (N_26250,N_23577,N_21575);
and U26251 (N_26251,N_24564,N_21625);
and U26252 (N_26252,N_23871,N_24868);
and U26253 (N_26253,N_23689,N_21095);
xor U26254 (N_26254,N_22865,N_23470);
xnor U26255 (N_26255,N_22494,N_21714);
and U26256 (N_26256,N_22673,N_22753);
xnor U26257 (N_26257,N_22468,N_24859);
nand U26258 (N_26258,N_22467,N_20010);
or U26259 (N_26259,N_23492,N_23870);
xor U26260 (N_26260,N_20548,N_20670);
and U26261 (N_26261,N_20204,N_21543);
nand U26262 (N_26262,N_23575,N_22725);
xor U26263 (N_26263,N_24663,N_20565);
nand U26264 (N_26264,N_21257,N_21531);
or U26265 (N_26265,N_24264,N_20206);
or U26266 (N_26266,N_20668,N_21482);
nor U26267 (N_26267,N_21430,N_24827);
xor U26268 (N_26268,N_23015,N_21036);
and U26269 (N_26269,N_20821,N_24823);
nor U26270 (N_26270,N_22780,N_22248);
and U26271 (N_26271,N_24603,N_24665);
nand U26272 (N_26272,N_24465,N_21974);
nand U26273 (N_26273,N_22081,N_22801);
xnor U26274 (N_26274,N_21745,N_20961);
xnor U26275 (N_26275,N_20454,N_23075);
or U26276 (N_26276,N_22413,N_22546);
nand U26277 (N_26277,N_24601,N_22430);
nor U26278 (N_26278,N_22204,N_20278);
xnor U26279 (N_26279,N_22939,N_23226);
or U26280 (N_26280,N_22404,N_20183);
and U26281 (N_26281,N_20978,N_22324);
xnor U26282 (N_26282,N_22386,N_21396);
nand U26283 (N_26283,N_23156,N_22824);
xor U26284 (N_26284,N_24187,N_22867);
nor U26285 (N_26285,N_24205,N_23810);
xor U26286 (N_26286,N_24838,N_24200);
and U26287 (N_26287,N_24267,N_24562);
and U26288 (N_26288,N_22881,N_20752);
or U26289 (N_26289,N_21189,N_21949);
xor U26290 (N_26290,N_23056,N_20489);
xnor U26291 (N_26291,N_21206,N_20395);
nor U26292 (N_26292,N_23599,N_22211);
and U26293 (N_26293,N_20776,N_24620);
nand U26294 (N_26294,N_24134,N_23006);
nor U26295 (N_26295,N_20350,N_21190);
nand U26296 (N_26296,N_22393,N_21046);
or U26297 (N_26297,N_22062,N_20295);
xnor U26298 (N_26298,N_24299,N_23134);
or U26299 (N_26299,N_20446,N_24094);
nand U26300 (N_26300,N_24282,N_23845);
nor U26301 (N_26301,N_24756,N_23174);
nor U26302 (N_26302,N_20203,N_21114);
or U26303 (N_26303,N_22325,N_24022);
xnor U26304 (N_26304,N_21823,N_24098);
nor U26305 (N_26305,N_23911,N_20580);
and U26306 (N_26306,N_23926,N_21278);
xnor U26307 (N_26307,N_22462,N_20140);
or U26308 (N_26308,N_23597,N_21792);
or U26309 (N_26309,N_24637,N_21198);
and U26310 (N_26310,N_22566,N_23285);
or U26311 (N_26311,N_20520,N_20671);
and U26312 (N_26312,N_24108,N_22850);
or U26313 (N_26313,N_23525,N_23246);
nand U26314 (N_26314,N_23589,N_24907);
and U26315 (N_26315,N_24769,N_21790);
nor U26316 (N_26316,N_24869,N_24149);
and U26317 (N_26317,N_20051,N_24411);
and U26318 (N_26318,N_21306,N_24640);
and U26319 (N_26319,N_20717,N_21225);
nor U26320 (N_26320,N_20998,N_24233);
xor U26321 (N_26321,N_24122,N_22210);
xor U26322 (N_26322,N_21922,N_23973);
xnor U26323 (N_26323,N_20333,N_21176);
and U26324 (N_26324,N_21373,N_22135);
xnor U26325 (N_26325,N_24714,N_24452);
and U26326 (N_26326,N_22807,N_22570);
nor U26327 (N_26327,N_20334,N_20996);
nand U26328 (N_26328,N_24765,N_23144);
and U26329 (N_26329,N_23042,N_22258);
nand U26330 (N_26330,N_22857,N_24126);
nand U26331 (N_26331,N_23010,N_23036);
xor U26332 (N_26332,N_23551,N_23078);
and U26333 (N_26333,N_21081,N_20700);
or U26334 (N_26334,N_20572,N_24766);
nor U26335 (N_26335,N_23003,N_24083);
nor U26336 (N_26336,N_21485,N_24011);
nor U26337 (N_26337,N_22607,N_21332);
nand U26338 (N_26338,N_24651,N_22563);
or U26339 (N_26339,N_24537,N_24468);
xor U26340 (N_26340,N_21261,N_20907);
and U26341 (N_26341,N_23106,N_23813);
xor U26342 (N_26342,N_20275,N_24639);
nand U26343 (N_26343,N_23199,N_23334);
or U26344 (N_26344,N_23209,N_24298);
nand U26345 (N_26345,N_21581,N_24285);
xor U26346 (N_26346,N_21825,N_22284);
xnor U26347 (N_26347,N_22730,N_22263);
nand U26348 (N_26348,N_20846,N_22143);
and U26349 (N_26349,N_21989,N_20942);
xnor U26350 (N_26350,N_20447,N_23090);
nand U26351 (N_26351,N_23713,N_20097);
and U26352 (N_26352,N_22232,N_21927);
nand U26353 (N_26353,N_22929,N_23214);
nor U26354 (N_26354,N_22727,N_23225);
nand U26355 (N_26355,N_21920,N_23749);
xnor U26356 (N_26356,N_22283,N_21935);
nor U26357 (N_26357,N_21309,N_23628);
nand U26358 (N_26358,N_21378,N_21040);
nor U26359 (N_26359,N_21769,N_22158);
xnor U26360 (N_26360,N_22340,N_24317);
nor U26361 (N_26361,N_23183,N_23008);
xnor U26362 (N_26362,N_23877,N_23351);
and U26363 (N_26363,N_24578,N_20138);
and U26364 (N_26364,N_24692,N_24471);
nand U26365 (N_26365,N_23821,N_23352);
nand U26366 (N_26366,N_24435,N_24136);
or U26367 (N_26367,N_23919,N_24429);
nand U26368 (N_26368,N_24417,N_23933);
nand U26369 (N_26369,N_20375,N_21680);
nand U26370 (N_26370,N_21318,N_24141);
and U26371 (N_26371,N_20083,N_23725);
xnor U26372 (N_26372,N_24626,N_23699);
nand U26373 (N_26373,N_21009,N_21393);
xnor U26374 (N_26374,N_23882,N_23867);
and U26375 (N_26375,N_21407,N_24922);
nand U26376 (N_26376,N_21458,N_22797);
or U26377 (N_26377,N_20870,N_22828);
nor U26378 (N_26378,N_22989,N_22771);
nand U26379 (N_26379,N_20540,N_24925);
or U26380 (N_26380,N_22816,N_20063);
or U26381 (N_26381,N_24153,N_23354);
nand U26382 (N_26382,N_23405,N_20522);
nor U26383 (N_26383,N_23256,N_20610);
nor U26384 (N_26384,N_20733,N_22904);
and U26385 (N_26385,N_24462,N_21509);
and U26386 (N_26386,N_24382,N_21726);
nand U26387 (N_26387,N_23993,N_21124);
nor U26388 (N_26388,N_24234,N_22086);
and U26389 (N_26389,N_22599,N_20076);
nand U26390 (N_26390,N_23864,N_24793);
xnor U26391 (N_26391,N_24390,N_22305);
nor U26392 (N_26392,N_24001,N_21491);
nand U26393 (N_26393,N_22769,N_21171);
nand U26394 (N_26394,N_23222,N_21473);
nand U26395 (N_26395,N_23802,N_21650);
xor U26396 (N_26396,N_21894,N_24451);
nand U26397 (N_26397,N_21386,N_22175);
nand U26398 (N_26398,N_23522,N_22577);
nand U26399 (N_26399,N_20770,N_22497);
or U26400 (N_26400,N_24871,N_22372);
xnor U26401 (N_26401,N_21853,N_22666);
and U26402 (N_26402,N_24987,N_20645);
nand U26403 (N_26403,N_20810,N_21708);
nand U26404 (N_26404,N_22151,N_21079);
or U26405 (N_26405,N_20971,N_21432);
nor U26406 (N_26406,N_24785,N_23276);
nor U26407 (N_26407,N_22479,N_21500);
xor U26408 (N_26408,N_23668,N_23158);
or U26409 (N_26409,N_23094,N_24125);
nor U26410 (N_26410,N_21788,N_24523);
nand U26411 (N_26411,N_23887,N_20586);
nand U26412 (N_26412,N_20184,N_20555);
nand U26413 (N_26413,N_20237,N_22892);
nand U26414 (N_26414,N_23550,N_21658);
nand U26415 (N_26415,N_22192,N_20400);
and U26416 (N_26416,N_21074,N_23086);
or U26417 (N_26417,N_23540,N_22058);
nand U26418 (N_26418,N_24220,N_21728);
and U26419 (N_26419,N_23348,N_21371);
xnor U26420 (N_26420,N_21183,N_21069);
or U26421 (N_26421,N_24346,N_20858);
nor U26422 (N_26422,N_24068,N_20408);
xnor U26423 (N_26423,N_24669,N_24161);
xor U26424 (N_26424,N_24770,N_23320);
or U26425 (N_26425,N_22854,N_23207);
nor U26426 (N_26426,N_23139,N_21685);
xnor U26427 (N_26427,N_23667,N_22026);
nor U26428 (N_26428,N_22740,N_24436);
or U26429 (N_26429,N_21159,N_21101);
or U26430 (N_26430,N_21231,N_21182);
or U26431 (N_26431,N_24421,N_23065);
or U26432 (N_26432,N_21550,N_24686);
nand U26433 (N_26433,N_22680,N_20820);
xor U26434 (N_26434,N_24235,N_23601);
or U26435 (N_26435,N_22392,N_22840);
and U26436 (N_26436,N_24543,N_23271);
and U26437 (N_26437,N_21273,N_22295);
nand U26438 (N_26438,N_23992,N_21653);
xnor U26439 (N_26439,N_24722,N_24271);
and U26440 (N_26440,N_21104,N_24290);
or U26441 (N_26441,N_20888,N_23644);
xnor U26442 (N_26442,N_24531,N_20800);
xor U26443 (N_26443,N_24890,N_23519);
xor U26444 (N_26444,N_21524,N_20473);
or U26445 (N_26445,N_22435,N_20116);
xnor U26446 (N_26446,N_22507,N_20911);
xnor U26447 (N_26447,N_20343,N_21238);
xnor U26448 (N_26448,N_22174,N_24558);
and U26449 (N_26449,N_23242,N_24368);
and U26450 (N_26450,N_24113,N_22712);
xor U26451 (N_26451,N_21914,N_20796);
xnor U26452 (N_26452,N_20927,N_24924);
nor U26453 (N_26453,N_22696,N_23193);
nor U26454 (N_26454,N_20159,N_21814);
nand U26455 (N_26455,N_24776,N_22410);
or U26456 (N_26456,N_23529,N_23319);
nand U26457 (N_26457,N_23148,N_24590);
or U26458 (N_26458,N_24064,N_21690);
nor U26459 (N_26459,N_22574,N_23968);
nor U26460 (N_26460,N_20659,N_21389);
xnor U26461 (N_26461,N_20475,N_20423);
xor U26462 (N_26462,N_20258,N_24214);
nor U26463 (N_26463,N_24172,N_24132);
xor U26464 (N_26464,N_24046,N_21635);
or U26465 (N_26465,N_20771,N_21966);
nor U26466 (N_26466,N_21808,N_22954);
xor U26467 (N_26467,N_20310,N_20591);
and U26468 (N_26468,N_22356,N_21490);
nor U26469 (N_26469,N_24069,N_24887);
xnor U26470 (N_26470,N_23582,N_20594);
xnor U26471 (N_26471,N_21882,N_20213);
nand U26472 (N_26472,N_22027,N_24848);
or U26473 (N_26473,N_20744,N_20536);
nor U26474 (N_26474,N_24326,N_23935);
xor U26475 (N_26475,N_23642,N_24104);
nand U26476 (N_26476,N_23897,N_20741);
nand U26477 (N_26477,N_20398,N_20492);
xnor U26478 (N_26478,N_21630,N_22610);
and U26479 (N_26479,N_22334,N_20884);
nor U26480 (N_26480,N_23037,N_21770);
xor U26481 (N_26481,N_21224,N_20040);
and U26482 (N_26482,N_20518,N_22123);
nor U26483 (N_26483,N_23696,N_23059);
nor U26484 (N_26484,N_22804,N_20962);
and U26485 (N_26485,N_22022,N_20485);
nor U26486 (N_26486,N_20964,N_23531);
or U26487 (N_26487,N_21038,N_24963);
nor U26488 (N_26488,N_22299,N_23101);
nand U26489 (N_26489,N_20675,N_24596);
nand U26490 (N_26490,N_21453,N_21706);
nor U26491 (N_26491,N_21215,N_20011);
xor U26492 (N_26492,N_23609,N_23336);
or U26493 (N_26493,N_22671,N_20587);
or U26494 (N_26494,N_24926,N_22319);
and U26495 (N_26495,N_21672,N_20850);
or U26496 (N_26496,N_23829,N_24016);
nor U26497 (N_26497,N_24850,N_20910);
nor U26498 (N_26498,N_22631,N_24331);
or U26499 (N_26499,N_23709,N_21886);
nand U26500 (N_26500,N_23103,N_22554);
or U26501 (N_26501,N_21228,N_21739);
nor U26502 (N_26502,N_22506,N_21315);
nand U26503 (N_26503,N_22365,N_20166);
xnor U26504 (N_26504,N_20621,N_20628);
xnor U26505 (N_26505,N_21222,N_20758);
xnor U26506 (N_26506,N_21188,N_20901);
or U26507 (N_26507,N_24086,N_21398);
nand U26508 (N_26508,N_23371,N_20096);
nand U26509 (N_26509,N_20974,N_20619);
or U26510 (N_26510,N_20030,N_23671);
nor U26511 (N_26511,N_20298,N_21521);
and U26512 (N_26512,N_20513,N_24041);
nor U26513 (N_26513,N_20221,N_20553);
and U26514 (N_26514,N_22361,N_23423);
nor U26515 (N_26515,N_23886,N_23410);
nand U26516 (N_26516,N_24289,N_22784);
xnor U26517 (N_26517,N_20727,N_24645);
nand U26518 (N_26518,N_20092,N_24076);
and U26519 (N_26519,N_20002,N_22911);
xnor U26520 (N_26520,N_20932,N_21116);
xor U26521 (N_26521,N_24400,N_23636);
and U26522 (N_26522,N_20093,N_22344);
nand U26523 (N_26523,N_21715,N_24565);
and U26524 (N_26524,N_21687,N_23077);
and U26525 (N_26525,N_23344,N_24862);
nand U26526 (N_26526,N_20605,N_20613);
nand U26527 (N_26527,N_22122,N_24627);
or U26528 (N_26528,N_21900,N_22265);
or U26529 (N_26529,N_24280,N_20601);
nor U26530 (N_26530,N_24655,N_23512);
or U26531 (N_26531,N_22314,N_20056);
or U26532 (N_26532,N_21768,N_23128);
xor U26533 (N_26533,N_24342,N_24171);
nor U26534 (N_26534,N_21078,N_21804);
or U26535 (N_26535,N_20544,N_24847);
nand U26536 (N_26536,N_22738,N_22601);
nand U26537 (N_26537,N_23568,N_22354);
and U26538 (N_26538,N_22065,N_23970);
nor U26539 (N_26539,N_20703,N_20460);
nor U26540 (N_26540,N_20797,N_23343);
nor U26541 (N_26541,N_23704,N_21860);
nand U26542 (N_26542,N_24588,N_22833);
nand U26543 (N_26543,N_21233,N_23982);
and U26544 (N_26544,N_23324,N_20364);
nor U26545 (N_26545,N_23804,N_20865);
nand U26546 (N_26546,N_21255,N_23373);
or U26547 (N_26547,N_20622,N_22097);
xor U26548 (N_26548,N_21695,N_21995);
xnor U26549 (N_26549,N_21569,N_23118);
nand U26550 (N_26550,N_21175,N_22432);
xor U26551 (N_26551,N_24881,N_23756);
nor U26552 (N_26552,N_22256,N_21129);
xor U26553 (N_26553,N_20250,N_22960);
or U26554 (N_26554,N_24049,N_21288);
nor U26555 (N_26555,N_20564,N_23815);
xor U26556 (N_26556,N_20311,N_23241);
xnor U26557 (N_26557,N_24443,N_24082);
and U26558 (N_26558,N_23708,N_20146);
or U26559 (N_26559,N_20955,N_21696);
nor U26560 (N_26560,N_23734,N_20879);
and U26561 (N_26561,N_21738,N_24541);
or U26562 (N_26562,N_22117,N_20684);
nor U26563 (N_26563,N_24554,N_21590);
xnor U26564 (N_26564,N_23913,N_20122);
xor U26565 (N_26565,N_24959,N_22517);
or U26566 (N_26566,N_22201,N_22406);
nor U26567 (N_26567,N_24067,N_22141);
xor U26568 (N_26568,N_23493,N_24319);
and U26569 (N_26569,N_21134,N_22917);
xnor U26570 (N_26570,N_20281,N_22933);
nor U26571 (N_26571,N_22481,N_21713);
nand U26572 (N_26572,N_23233,N_21947);
nand U26573 (N_26573,N_24727,N_22821);
and U26574 (N_26574,N_23132,N_24767);
and U26575 (N_26575,N_24813,N_20242);
and U26576 (N_26576,N_23147,N_21880);
nor U26577 (N_26577,N_21083,N_21855);
and U26578 (N_26578,N_20813,N_21244);
or U26579 (N_26579,N_20608,N_22644);
xnor U26580 (N_26580,N_21066,N_20325);
or U26581 (N_26581,N_22714,N_21474);
xnor U26582 (N_26582,N_21050,N_20817);
xor U26583 (N_26583,N_22716,N_23607);
xor U26584 (N_26584,N_21863,N_23977);
nand U26585 (N_26585,N_20067,N_22267);
nor U26586 (N_26586,N_23808,N_21854);
xnor U26587 (N_26587,N_24169,N_20351);
nor U26588 (N_26588,N_21007,N_20009);
nor U26589 (N_26589,N_22375,N_21756);
nand U26590 (N_26590,N_23463,N_21859);
or U26591 (N_26591,N_22450,N_21821);
nor U26592 (N_26592,N_21937,N_24273);
nor U26593 (N_26593,N_24597,N_24943);
and U26594 (N_26594,N_23173,N_24361);
xor U26595 (N_26595,N_20449,N_23030);
nand U26596 (N_26596,N_24237,N_20050);
nand U26597 (N_26597,N_20201,N_20855);
and U26598 (N_26598,N_21166,N_21185);
xnor U26599 (N_26599,N_23311,N_24824);
nor U26600 (N_26600,N_22791,N_24518);
xnor U26601 (N_26601,N_24958,N_20153);
and U26602 (N_26602,N_23960,N_24980);
xnor U26603 (N_26603,N_22995,N_21701);
xnor U26604 (N_26604,N_24875,N_22617);
and U26605 (N_26605,N_20690,N_22032);
xnor U26606 (N_26606,N_22735,N_24355);
xnor U26607 (N_26607,N_24652,N_21666);
or U26608 (N_26608,N_20725,N_20249);
nor U26609 (N_26609,N_24506,N_21841);
or U26610 (N_26610,N_23648,N_21970);
or U26611 (N_26611,N_22626,N_20365);
or U26612 (N_26612,N_22868,N_20384);
and U26613 (N_26613,N_22001,N_24883);
and U26614 (N_26614,N_21622,N_20413);
nor U26615 (N_26615,N_23473,N_20970);
and U26616 (N_26616,N_21299,N_23710);
xor U26617 (N_26617,N_24764,N_21368);
or U26618 (N_26618,N_21561,N_24021);
xor U26619 (N_26619,N_22394,N_20162);
xnor U26620 (N_26620,N_23112,N_21828);
nand U26621 (N_26621,N_23560,N_21866);
and U26622 (N_26622,N_20091,N_22709);
and U26623 (N_26623,N_24898,N_24879);
nand U26624 (N_26624,N_23794,N_21645);
and U26625 (N_26625,N_22503,N_20402);
xor U26626 (N_26626,N_20501,N_23360);
nor U26627 (N_26627,N_21584,N_23282);
nand U26628 (N_26628,N_21305,N_24664);
nand U26629 (N_26629,N_20642,N_24936);
and U26630 (N_26630,N_21938,N_22052);
or U26631 (N_26631,N_23542,N_21405);
or U26632 (N_26632,N_24369,N_22156);
or U26633 (N_26633,N_20556,N_23539);
or U26634 (N_26634,N_22118,N_23735);
xnor U26635 (N_26635,N_20077,N_21323);
or U26636 (N_26636,N_20929,N_20000);
xor U26637 (N_26637,N_24777,N_23924);
and U26638 (N_26638,N_23895,N_23228);
xnor U26639 (N_26639,N_21778,N_24533);
nor U26640 (N_26640,N_23363,N_20066);
nor U26641 (N_26641,N_20302,N_22756);
nor U26642 (N_26642,N_21885,N_24102);
and U26643 (N_26643,N_24886,N_20458);
xnor U26644 (N_26644,N_22776,N_23670);
nand U26645 (N_26645,N_23608,N_20968);
nand U26646 (N_26646,N_22576,N_22035);
or U26647 (N_26647,N_23554,N_21400);
and U26648 (N_26648,N_23931,N_23510);
xnor U26649 (N_26649,N_23868,N_23663);
or U26650 (N_26650,N_23884,N_22051);
xor U26651 (N_26651,N_21585,N_20361);
nor U26652 (N_26652,N_20358,N_21092);
nor U26653 (N_26653,N_21365,N_20304);
or U26654 (N_26654,N_22736,N_20977);
nor U26655 (N_26655,N_20985,N_21641);
nand U26656 (N_26656,N_22385,N_21588);
and U26657 (N_26657,N_23672,N_22670);
nor U26658 (N_26658,N_22043,N_23085);
nor U26659 (N_26659,N_22031,N_24865);
and U26660 (N_26660,N_20426,N_21002);
xnor U26661 (N_26661,N_24634,N_20346);
nand U26662 (N_26662,N_20336,N_21043);
xor U26663 (N_26663,N_22661,N_22106);
nand U26664 (N_26664,N_24373,N_21893);
or U26665 (N_26665,N_20827,N_21593);
nand U26666 (N_26666,N_21602,N_21815);
xnor U26667 (N_26667,N_20988,N_21447);
or U26668 (N_26668,N_23308,N_21283);
nor U26669 (N_26669,N_21952,N_24103);
nand U26670 (N_26670,N_20244,N_24357);
xnor U26671 (N_26671,N_23105,N_24441);
or U26672 (N_26672,N_20957,N_21201);
or U26673 (N_26673,N_22465,N_20516);
nor U26674 (N_26674,N_22167,N_22436);
xnor U26675 (N_26675,N_21138,N_21425);
xor U26676 (N_26676,N_21291,N_24129);
and U26677 (N_26677,N_23165,N_20603);
nor U26678 (N_26678,N_20976,N_24397);
xor U26679 (N_26679,N_22213,N_20347);
nor U26680 (N_26680,N_20852,N_23765);
nor U26681 (N_26681,N_22103,N_20514);
nor U26682 (N_26682,N_23558,N_21004);
xor U26683 (N_26683,N_21888,N_24328);
nand U26684 (N_26684,N_21620,N_24270);
and U26685 (N_26685,N_22346,N_22587);
nand U26686 (N_26686,N_22274,N_20190);
and U26687 (N_26687,N_23523,N_22955);
or U26688 (N_26688,N_22163,N_21797);
nor U26689 (N_26689,N_23123,N_22069);
nand U26690 (N_26690,N_20452,N_24795);
or U26691 (N_26691,N_21498,N_22971);
and U26692 (N_26692,N_22469,N_23468);
nand U26693 (N_26693,N_21411,N_20113);
or U26694 (N_26694,N_23184,N_21609);
and U26695 (N_26695,N_21926,N_20828);
or U26696 (N_26696,N_23267,N_23760);
or U26697 (N_26697,N_21452,N_21254);
or U26698 (N_26698,N_21767,N_23254);
or U26699 (N_26699,N_23494,N_22741);
nor U26700 (N_26700,N_21399,N_21436);
or U26701 (N_26701,N_21890,N_24580);
xnor U26702 (N_26702,N_24105,N_24176);
or U26703 (N_26703,N_23450,N_21060);
nor U26704 (N_26704,N_21918,N_22656);
and U26705 (N_26705,N_23976,N_24741);
nor U26706 (N_26706,N_22766,N_22194);
nand U26707 (N_26707,N_20759,N_21144);
or U26708 (N_26708,N_21518,N_24150);
nand U26709 (N_26709,N_23102,N_22663);
and U26710 (N_26710,N_23635,N_23380);
nand U26711 (N_26711,N_22338,N_22676);
and U26712 (N_26712,N_22053,N_22417);
xor U26713 (N_26713,N_20005,N_20568);
or U26714 (N_26714,N_21208,N_21372);
or U26715 (N_26715,N_20533,N_24467);
or U26716 (N_26716,N_24434,N_23303);
nand U26717 (N_26717,N_20864,N_21232);
nor U26718 (N_26718,N_24843,N_23863);
and U26719 (N_26719,N_24519,N_21557);
and U26720 (N_26720,N_21048,N_23298);
nand U26721 (N_26721,N_23849,N_24930);
or U26722 (N_26722,N_20896,N_24399);
xnor U26723 (N_26723,N_24891,N_22216);
or U26724 (N_26724,N_20842,N_24502);
or U26725 (N_26725,N_24413,N_24142);
or U26726 (N_26726,N_20880,N_20719);
nand U26727 (N_26727,N_24301,N_22997);
or U26728 (N_26728,N_22754,N_23684);
xnor U26729 (N_26729,N_21087,N_21292);
nor U26730 (N_26730,N_21711,N_20422);
xor U26731 (N_26731,N_22454,N_20893);
nand U26732 (N_26732,N_21909,N_21401);
nor U26733 (N_26733,N_21161,N_24927);
or U26734 (N_26734,N_24458,N_22102);
nand U26735 (N_26735,N_22477,N_20933);
xor U26736 (N_26736,N_23881,N_23959);
nor U26737 (N_26737,N_24923,N_20900);
xnor U26738 (N_26738,N_22706,N_23941);
nand U26739 (N_26739,N_20394,N_20174);
xnor U26740 (N_26740,N_22016,N_22658);
or U26741 (N_26741,N_24196,N_20775);
xor U26742 (N_26742,N_21758,N_22910);
and U26743 (N_26743,N_23500,N_22819);
nand U26744 (N_26744,N_24147,N_20055);
nand U26745 (N_26745,N_20425,N_24052);
nor U26746 (N_26746,N_22442,N_23898);
and U26747 (N_26747,N_24834,N_20300);
or U26748 (N_26748,N_24659,N_24556);
or U26749 (N_26749,N_20825,N_23179);
xor U26750 (N_26750,N_22379,N_22105);
or U26751 (N_26751,N_21221,N_24089);
xor U26752 (N_26752,N_20194,N_23872);
xor U26753 (N_26753,N_22445,N_20757);
nor U26754 (N_26754,N_24008,N_24291);
nand U26755 (N_26755,N_21994,N_21736);
and U26756 (N_26756,N_23874,N_22830);
nand U26757 (N_26757,N_23971,N_21403);
nand U26758 (N_26758,N_20705,N_20161);
and U26759 (N_26759,N_23602,N_21014);
nand U26760 (N_26760,N_20578,N_23322);
xor U26761 (N_26761,N_21956,N_22304);
nor U26762 (N_26762,N_20845,N_21253);
nor U26763 (N_26763,N_20644,N_22789);
nand U26764 (N_26764,N_22558,N_23692);
and U26765 (N_26765,N_21249,N_22810);
nand U26766 (N_26766,N_24917,N_21686);
xnor U26767 (N_26767,N_23506,N_22302);
or U26768 (N_26768,N_24673,N_22480);
nand U26769 (N_26769,N_20014,N_20920);
or U26770 (N_26770,N_24158,N_23388);
nand U26771 (N_26771,N_20388,N_24783);
nor U26772 (N_26772,N_22856,N_21674);
xnor U26773 (N_26773,N_23401,N_22996);
nand U26774 (N_26774,N_20407,N_24494);
or U26775 (N_26775,N_24340,N_24329);
nand U26776 (N_26776,N_22315,N_24739);
nand U26777 (N_26777,N_24444,N_20925);
or U26778 (N_26778,N_24870,N_24999);
nor U26779 (N_26779,N_20678,N_23624);
nand U26780 (N_26780,N_20354,N_21933);
or U26781 (N_26781,N_23465,N_24629);
or U26782 (N_26782,N_21180,N_21580);
or U26783 (N_26783,N_22902,N_20223);
nand U26784 (N_26784,N_24432,N_22475);
and U26785 (N_26785,N_24803,N_22183);
and U26786 (N_26786,N_20650,N_23737);
or U26787 (N_26787,N_24807,N_21042);
xnor U26788 (N_26788,N_23172,N_20405);
nor U26789 (N_26789,N_20012,N_23339);
xor U26790 (N_26790,N_21143,N_21313);
and U26791 (N_26791,N_22708,N_24527);
nand U26792 (N_26792,N_21382,N_22172);
nor U26793 (N_26793,N_23223,N_24062);
or U26794 (N_26794,N_23561,N_23803);
or U26795 (N_26795,N_22518,N_23530);
nor U26796 (N_26796,N_22614,N_23980);
nand U26797 (N_26797,N_20611,N_20117);
xnor U26798 (N_26798,N_23703,N_20192);
or U26799 (N_26799,N_22767,N_21419);
or U26800 (N_26800,N_23033,N_20429);
nor U26801 (N_26801,N_24638,N_21142);
or U26802 (N_26802,N_21902,N_23185);
or U26803 (N_26803,N_22969,N_21623);
xor U26804 (N_26804,N_22072,N_21165);
or U26805 (N_26805,N_24706,N_20393);
xor U26806 (N_26806,N_21527,N_22188);
and U26807 (N_26807,N_20760,N_24260);
or U26808 (N_26808,N_22664,N_22040);
nand U26809 (N_26809,N_23399,N_23449);
nor U26810 (N_26810,N_20916,N_23787);
or U26811 (N_26811,N_24584,N_20124);
nor U26812 (N_26812,N_23004,N_20763);
or U26813 (N_26813,N_24127,N_24811);
or U26814 (N_26814,N_24206,N_24644);
nor U26815 (N_26815,N_22254,N_20039);
xnor U26816 (N_26816,N_20994,N_24058);
nor U26817 (N_26817,N_23457,N_22421);
nor U26818 (N_26818,N_21137,N_23038);
nand U26819 (N_26819,N_24899,N_20089);
or U26820 (N_26820,N_24955,N_20137);
nor U26821 (N_26821,N_20477,N_24902);
or U26822 (N_26822,N_24003,N_22473);
xnor U26823 (N_26823,N_22060,N_24809);
nor U26824 (N_26824,N_24374,N_24616);
and U26825 (N_26825,N_23023,N_21470);
xnor U26826 (N_26826,N_20253,N_23262);
nand U26827 (N_26827,N_24636,N_22602);
xor U26828 (N_26828,N_22702,N_20573);
xor U26829 (N_26829,N_22679,N_20478);
xor U26830 (N_26830,N_24116,N_22591);
nor U26831 (N_26831,N_24977,N_24863);
xnor U26832 (N_26832,N_22329,N_23905);
or U26833 (N_26833,N_20114,N_22352);
nand U26834 (N_26834,N_20860,N_21646);
and U26835 (N_26835,N_20189,N_21595);
nor U26836 (N_26836,N_20546,N_20188);
xor U26837 (N_26837,N_20926,N_24532);
xor U26838 (N_26838,N_23259,N_21954);
nand U26839 (N_26839,N_24683,N_24740);
xor U26840 (N_26840,N_21476,N_21194);
or U26841 (N_26841,N_23833,N_20303);
and U26842 (N_26842,N_21096,N_22620);
or U26843 (N_26843,N_23604,N_21598);
nor U26844 (N_26844,N_21551,N_22870);
nand U26845 (N_26845,N_21235,N_24855);
and U26846 (N_26846,N_24447,N_23208);
or U26847 (N_26847,N_22486,N_20847);
nor U26848 (N_26848,N_20950,N_21410);
and U26849 (N_26849,N_24359,N_20767);
or U26850 (N_26850,N_20028,N_24111);
and U26851 (N_26851,N_24962,N_23581);
and U26852 (N_26852,N_22758,N_20627);
nand U26853 (N_26853,N_22286,N_21229);
or U26854 (N_26854,N_22768,N_20997);
and U26855 (N_26855,N_20216,N_23865);
nor U26856 (N_26856,N_20470,N_20685);
nand U26857 (N_26857,N_22277,N_22157);
xor U26858 (N_26858,N_22509,N_24942);
nand U26859 (N_26859,N_22139,N_24981);
nor U26860 (N_26860,N_21298,N_21872);
and U26861 (N_26861,N_23443,N_22212);
xor U26862 (N_26862,N_22489,N_21251);
xnor U26863 (N_26863,N_20663,N_21125);
nand U26864 (N_26864,N_20360,N_21459);
xor U26865 (N_26865,N_24489,N_21428);
xor U26866 (N_26866,N_20418,N_23612);
xor U26867 (N_26867,N_23681,N_24685);
nand U26868 (N_26868,N_20954,N_20320);
nor U26869 (N_26869,N_20891,N_20723);
nand U26870 (N_26870,N_23869,N_21274);
xor U26871 (N_26871,N_21631,N_22594);
nand U26872 (N_26872,N_24906,N_20936);
and U26873 (N_26873,N_20255,N_20881);
xnor U26874 (N_26874,N_21058,N_20434);
nand U26875 (N_26875,N_22249,N_24222);
and U26876 (N_26876,N_23583,N_20951);
or U26877 (N_26877,N_23835,N_20778);
and U26878 (N_26878,N_21383,N_20430);
or U26879 (N_26879,N_23318,N_23691);
or U26880 (N_26880,N_24151,N_23313);
xor U26881 (N_26881,N_23511,N_24313);
nor U26882 (N_26882,N_20777,N_23451);
nand U26883 (N_26883,N_23485,N_23890);
and U26884 (N_26884,N_23836,N_20593);
and U26885 (N_26885,N_23381,N_23594);
nand U26886 (N_26886,N_24555,N_24190);
xor U26887 (N_26887,N_20539,N_23934);
xnor U26888 (N_26888,N_21671,N_24073);
and U26889 (N_26889,N_20637,N_20383);
and U26890 (N_26890,N_21390,N_22616);
xor U26891 (N_26891,N_23626,N_22501);
nor U26892 (N_26892,N_22496,N_23946);
nand U26893 (N_26893,N_23161,N_24232);
nand U26894 (N_26894,N_20786,N_24395);
nor U26895 (N_26895,N_24884,N_23907);
and U26896 (N_26896,N_21765,N_21614);
xnor U26897 (N_26897,N_23967,N_22297);
and U26898 (N_26898,N_20440,N_22611);
nor U26899 (N_26899,N_24830,N_24146);
nand U26900 (N_26900,N_24715,N_20001);
nand U26901 (N_26901,N_21733,N_23482);
or U26902 (N_26902,N_22428,N_22593);
and U26903 (N_26903,N_23961,N_21033);
and U26904 (N_26904,N_23894,N_22888);
nand U26905 (N_26905,N_22389,N_22612);
and U26906 (N_26906,N_20698,N_24275);
and U26907 (N_26907,N_21529,N_20180);
and U26908 (N_26908,N_23483,N_23745);
or U26909 (N_26909,N_24408,N_23367);
nand U26910 (N_26910,N_23850,N_22922);
and U26911 (N_26911,N_22094,N_23480);
and U26912 (N_26912,N_22321,N_23437);
or U26913 (N_26913,N_20085,N_22710);
or U26914 (N_26914,N_23151,N_23912);
nor U26915 (N_26915,N_20736,N_22985);
and U26916 (N_26916,N_20773,N_20504);
nand U26917 (N_26917,N_20196,N_22448);
or U26918 (N_26918,N_24723,N_23261);
nand U26919 (N_26919,N_20948,N_23537);
xnor U26920 (N_26920,N_22678,N_22595);
and U26921 (N_26921,N_23953,N_24250);
nor U26922 (N_26922,N_20505,N_22074);
or U26923 (N_26923,N_20582,N_24004);
or U26924 (N_26924,N_20006,N_20139);
and U26925 (N_26925,N_21718,N_24998);
or U26926 (N_26926,N_23518,N_21560);
nor U26927 (N_26927,N_20472,N_24476);
nand U26928 (N_26928,N_24545,N_23900);
nor U26929 (N_26929,N_20202,N_22550);
or U26930 (N_26930,N_24778,N_24385);
xnor U26931 (N_26931,N_24375,N_23383);
or U26932 (N_26932,N_21919,N_23698);
xnor U26933 (N_26933,N_20324,N_24949);
nand U26934 (N_26934,N_20782,N_23954);
nand U26935 (N_26935,N_23823,N_23521);
and U26936 (N_26936,N_23797,N_23929);
and U26937 (N_26937,N_23486,N_24225);
or U26938 (N_26938,N_21735,N_22765);
nor U26939 (N_26939,N_22779,N_24839);
or U26940 (N_26940,N_24002,N_21112);
nand U26941 (N_26941,N_21415,N_21960);
and U26942 (N_26942,N_22308,N_22944);
xnor U26943 (N_26943,N_22077,N_22849);
nand U26944 (N_26944,N_21089,N_24177);
xnor U26945 (N_26945,N_20863,N_23166);
xor U26946 (N_26946,N_24055,N_22839);
nor U26947 (N_26947,N_22640,N_22343);
or U26948 (N_26948,N_24503,N_24166);
xnor U26949 (N_26949,N_24873,N_20299);
nand U26950 (N_26950,N_20367,N_22536);
nor U26951 (N_26951,N_21105,N_22585);
nand U26952 (N_26952,N_21884,N_22942);
nor U26953 (N_26953,N_24380,N_22622);
nor U26954 (N_26954,N_23293,N_22088);
and U26955 (N_26955,N_23679,N_23175);
nand U26956 (N_26956,N_23169,N_23365);
or U26957 (N_26957,N_20563,N_21811);
nand U26958 (N_26958,N_22625,N_22691);
and U26959 (N_26959,N_20531,N_20982);
nor U26960 (N_26960,N_24539,N_24208);
xnor U26961 (N_26961,N_21267,N_22638);
nor U26962 (N_26962,N_22044,N_22987);
and U26963 (N_26963,N_21737,N_21868);
or U26964 (N_26964,N_23714,N_20886);
xor U26965 (N_26965,N_24705,N_20966);
nand U26966 (N_26966,N_21478,N_22245);
nand U26967 (N_26967,N_24713,N_22427);
nor U26968 (N_26968,N_24157,N_20232);
xor U26969 (N_26969,N_22453,N_20807);
xnor U26970 (N_26970,N_20207,N_24101);
nor U26971 (N_26971,N_21889,N_20195);
or U26972 (N_26972,N_22495,N_20370);
or U26973 (N_26973,N_21979,N_22402);
xnor U26974 (N_26974,N_23825,N_23357);
and U26975 (N_26975,N_21740,N_21435);
nand U26976 (N_26976,N_20459,N_22687);
or U26977 (N_26977,N_22983,N_23497);
or U26978 (N_26978,N_24247,N_22089);
nand U26979 (N_26979,N_20871,N_20024);
or U26980 (N_26980,N_23369,N_24188);
nor U26981 (N_26981,N_22894,N_24348);
nor U26982 (N_26982,N_22045,N_21566);
nand U26983 (N_26983,N_21925,N_22924);
or U26984 (N_26984,N_24544,N_20965);
and U26985 (N_26985,N_21367,N_20710);
or U26986 (N_26986,N_21747,N_23957);
xnor U26987 (N_26987,N_24512,N_21128);
or U26988 (N_26988,N_22510,N_24407);
nand U26989 (N_26989,N_21019,N_22918);
and U26990 (N_26990,N_22681,N_23295);
nand U26991 (N_26991,N_21071,N_21218);
and U26992 (N_26992,N_22378,N_23035);
nand U26993 (N_26993,N_23291,N_21845);
or U26994 (N_26994,N_20639,N_23618);
nand U26995 (N_26995,N_22134,N_21780);
and U26996 (N_26996,N_21642,N_22222);
xnor U26997 (N_26997,N_23114,N_24867);
nand U26998 (N_26998,N_21830,N_24454);
xnor U26999 (N_26999,N_24684,N_21983);
nor U27000 (N_27000,N_24658,N_24360);
nor U27001 (N_27001,N_20664,N_24394);
nand U27002 (N_27002,N_20722,N_20623);
or U27003 (N_27003,N_24897,N_22822);
and U27004 (N_27004,N_23801,N_20245);
nand U27005 (N_27005,N_21385,N_22300);
and U27006 (N_27006,N_21121,N_22943);
and U27007 (N_27007,N_23655,N_21270);
nor U27008 (N_27008,N_21990,N_20062);
xnor U27009 (N_27009,N_21784,N_21824);
xnor U27010 (N_27010,N_21619,N_23899);
nor U27011 (N_27011,N_21152,N_23192);
and U27012 (N_27012,N_22947,N_24931);
or U27013 (N_27013,N_21940,N_21468);
and U27014 (N_27014,N_22457,N_22749);
or U27015 (N_27015,N_22623,N_22262);
xor U27016 (N_27016,N_20340,N_23972);
nand U27017 (N_27017,N_24115,N_22013);
or U27018 (N_27018,N_20784,N_22963);
and U27019 (N_27019,N_22071,N_20837);
and U27020 (N_27020,N_23408,N_21260);
nand U27021 (N_27021,N_24928,N_24063);
and U27022 (N_27022,N_22817,N_21519);
nand U27023 (N_27023,N_21354,N_21460);
nor U27024 (N_27024,N_20112,N_24566);
nor U27025 (N_27025,N_21000,N_24207);
or U27026 (N_27026,N_24621,N_22782);
or U27027 (N_27027,N_22241,N_24763);
or U27028 (N_27028,N_20352,N_24656);
nor U27029 (N_27029,N_21542,N_24602);
xor U27030 (N_27030,N_20266,N_22449);
or U27031 (N_27031,N_23963,N_20561);
or U27032 (N_27032,N_23089,N_20297);
and U27033 (N_27033,N_23755,N_23559);
and U27034 (N_27034,N_20427,N_24305);
and U27035 (N_27035,N_24577,N_23885);
nand U27036 (N_27036,N_23816,N_22946);
nor U27037 (N_27037,N_20308,N_20296);
nor U27038 (N_27038,N_22719,N_22578);
xnor U27039 (N_27039,N_22516,N_23595);
nor U27040 (N_27040,N_20142,N_20646);
nor U27041 (N_27041,N_21637,N_23938);
and U27042 (N_27042,N_22447,N_24797);
xor U27043 (N_27043,N_23543,N_22650);
or U27044 (N_27044,N_20225,N_23774);
nor U27045 (N_27045,N_22535,N_21562);
nand U27046 (N_27046,N_21302,N_22025);
nand U27047 (N_27047,N_22036,N_21329);
xor U27048 (N_27048,N_20819,N_20765);
nand U27049 (N_27049,N_21099,N_22084);
xnor U27050 (N_27050,N_23922,N_20728);
nand U27051 (N_27051,N_22423,N_22737);
and U27052 (N_27052,N_22694,N_23221);
nor U27053 (N_27053,N_22147,N_21205);
or U27054 (N_27054,N_21852,N_23986);
nor U27055 (N_27055,N_22757,N_23068);
nor U27056 (N_27056,N_20571,N_20373);
nand U27057 (N_27057,N_23928,N_20371);
nand U27058 (N_27058,N_21670,N_24485);
or U27059 (N_27059,N_23034,N_21746);
xnor U27060 (N_27060,N_22632,N_23296);
or U27061 (N_27061,N_21835,N_21035);
nor U27062 (N_27062,N_22169,N_24743);
and U27063 (N_27063,N_24287,N_23364);
or U27064 (N_27064,N_23069,N_22846);
nand U27065 (N_27065,N_23430,N_22345);
nand U27066 (N_27066,N_22055,N_20774);
or U27067 (N_27067,N_21698,N_23818);
and U27068 (N_27068,N_23771,N_24091);
and U27069 (N_27069,N_23921,N_20596);
xnor U27070 (N_27070,N_23274,N_24325);
or U27071 (N_27071,N_22438,N_23508);
and U27072 (N_27072,N_23234,N_21462);
xor U27073 (N_27073,N_23441,N_23722);
xnor U27074 (N_27074,N_22289,N_23099);
and U27075 (N_27075,N_24170,N_24760);
xor U27076 (N_27076,N_23611,N_21945);
nand U27077 (N_27077,N_24888,N_24472);
nand U27078 (N_27078,N_21442,N_22531);
nand U27079 (N_27079,N_23490,N_22639);
or U27080 (N_27080,N_21554,N_23660);
nor U27081 (N_27081,N_21077,N_22312);
xnor U27082 (N_27082,N_23603,N_22845);
nand U27083 (N_27083,N_22384,N_20882);
nand U27084 (N_27084,N_22083,N_20444);
nand U27085 (N_27085,N_21339,N_23685);
and U27086 (N_27086,N_24033,N_21813);
nor U27087 (N_27087,N_24804,N_21132);
and U27088 (N_27088,N_24075,N_23171);
and U27089 (N_27089,N_21268,N_21901);
xor U27090 (N_27090,N_22234,N_24352);
and U27091 (N_27091,N_23189,N_20432);
nand U27092 (N_27092,N_23419,N_24653);
and U27093 (N_27093,N_20109,N_24524);
and U27094 (N_27094,N_23653,N_20256);
or U27095 (N_27095,N_21826,N_21904);
nor U27096 (N_27096,N_24700,N_23658);
nand U27097 (N_27097,N_22291,N_22061);
or U27098 (N_27098,N_20874,N_23697);
nor U27099 (N_27099,N_24787,N_23962);
nand U27100 (N_27100,N_21786,N_22006);
nand U27101 (N_27101,N_22568,N_20853);
nor U27102 (N_27102,N_22864,N_20498);
and U27103 (N_27103,N_20386,N_23386);
and U27104 (N_27104,N_24035,N_22812);
and U27105 (N_27105,N_24238,N_20185);
nand U27106 (N_27106,N_20387,N_23287);
and U27107 (N_27107,N_20890,N_21603);
xnor U27108 (N_27108,N_20665,N_20679);
and U27109 (N_27109,N_21213,N_21034);
xor U27110 (N_27110,N_21723,N_24535);
nand U27111 (N_27111,N_22545,N_22285);
and U27112 (N_27112,N_23338,N_21341);
xor U27113 (N_27113,N_22552,N_22793);
and U27114 (N_27114,N_20004,N_24406);
nor U27115 (N_27115,N_24882,N_22984);
or U27116 (N_27116,N_22651,N_22236);
or U27117 (N_27117,N_21499,N_20150);
nand U27118 (N_27118,N_22208,N_24514);
and U27119 (N_27119,N_21606,N_20766);
nor U27120 (N_27120,N_21340,N_23927);
and U27121 (N_27121,N_21731,N_21282);
nor U27122 (N_27122,N_21269,N_20785);
nand U27123 (N_27123,N_23431,N_22805);
nand U27124 (N_27124,N_20590,N_21583);
or U27125 (N_27125,N_23772,N_24817);
xnor U27126 (N_27126,N_22930,N_21856);
xnor U27127 (N_27127,N_23079,N_24424);
nand U27128 (N_27128,N_20424,N_22932);
nor U27129 (N_27129,N_23579,N_24175);
xnor U27130 (N_27130,N_22642,N_21605);
nand U27131 (N_27131,N_24351,N_22333);
and U27132 (N_27132,N_21799,N_23067);
and U27133 (N_27133,N_23140,N_21775);
xnor U27134 (N_27134,N_20355,N_21280);
or U27135 (N_27135,N_24470,N_24610);
and U27136 (N_27136,N_23964,N_20574);
nor U27137 (N_27137,N_21683,N_21944);
and U27138 (N_27138,N_23937,N_21891);
or U27139 (N_27139,N_24202,N_20037);
and U27140 (N_27140,N_22124,N_22958);
nand U27141 (N_27141,N_20476,N_21763);
nand U27142 (N_27142,N_22884,N_23235);
xnor U27143 (N_27143,N_20036,N_20652);
nor U27144 (N_27144,N_20729,N_21601);
and U27145 (N_27145,N_21162,N_22020);
and U27146 (N_27146,N_22978,N_24853);
or U27147 (N_27147,N_22703,N_22178);
xnor U27148 (N_27148,N_23409,N_24344);
xnor U27149 (N_27149,N_23789,N_24904);
nor U27150 (N_27150,N_22948,N_22556);
xor U27151 (N_27151,N_23923,N_23080);
xor U27152 (N_27152,N_23716,N_23436);
and U27153 (N_27153,N_22271,N_22390);
xor U27154 (N_27154,N_23790,N_20058);
xor U27155 (N_27155,N_24097,N_23839);
or U27156 (N_27156,N_21236,N_20079);
and U27157 (N_27157,N_23337,N_23424);
nand U27158 (N_27158,N_20779,N_24337);
and U27159 (N_27159,N_23154,N_24117);
or U27160 (N_27160,N_21955,N_21906);
nor U27161 (N_27161,N_20549,N_20486);
nand U27162 (N_27162,N_23314,N_22744);
nor U27163 (N_27163,N_22113,N_24991);
or U27164 (N_27164,N_23747,N_20284);
xnor U27165 (N_27165,N_24488,N_20374);
and U27166 (N_27166,N_24302,N_24510);
or U27167 (N_27167,N_22185,N_21564);
nand U27168 (N_27168,N_24324,N_24758);
nor U27169 (N_27169,N_22876,N_23576);
nor U27170 (N_27170,N_22499,N_24549);
xor U27171 (N_27171,N_20217,N_20327);
xor U27172 (N_27172,N_24420,N_24007);
or U27173 (N_27173,N_21155,N_20041);
xnor U27174 (N_27174,N_20944,N_21626);
and U27175 (N_27175,N_20843,N_24370);
or U27176 (N_27176,N_21193,N_20243);
or U27177 (N_27177,N_20552,N_21640);
or U27178 (N_27178,N_22363,N_23614);
and U27179 (N_27179,N_20963,N_20640);
xnor U27180 (N_27180,N_21053,N_21611);
and U27181 (N_27181,N_21361,N_24066);
nor U27182 (N_27182,N_22885,N_20980);
xor U27183 (N_27183,N_24525,N_24024);
or U27184 (N_27184,N_20338,N_21304);
xnor U27185 (N_27185,N_22257,N_21277);
nor U27186 (N_27186,N_21923,N_24401);
xnor U27187 (N_27187,N_23084,N_23495);
nor U27188 (N_27188,N_24174,N_23429);
and U27189 (N_27189,N_21356,N_24110);
and U27190 (N_27190,N_22675,N_24332);
and U27191 (N_27191,N_20396,N_24484);
or U27192 (N_27192,N_23918,N_23943);
nor U27193 (N_27193,N_21287,N_21342);
and U27194 (N_27194,N_22290,N_22377);
nand U27195 (N_27195,N_23627,N_23288);
nand U27196 (N_27196,N_20811,N_24154);
nor U27197 (N_27197,N_24481,N_24911);
or U27198 (N_27198,N_20943,N_24500);
nand U27199 (N_27199,N_24318,N_22893);
and U27200 (N_27200,N_22007,N_22313);
or U27201 (N_27201,N_22860,N_22136);
nand U27202 (N_27202,N_22974,N_21210);
xnor U27203 (N_27203,N_21985,N_22011);
nor U27204 (N_27204,N_22903,N_24199);
nand U27205 (N_27205,N_20313,N_23335);
nand U27206 (N_27206,N_23349,N_23880);
xor U27207 (N_27207,N_21170,N_22487);
and U27208 (N_27208,N_22560,N_21454);
or U27209 (N_27209,N_22880,N_20415);
or U27210 (N_27210,N_22891,N_21730);
nor U27211 (N_27211,N_24276,N_23715);
xor U27212 (N_27212,N_24426,N_20301);
nand U27213 (N_27213,N_23557,N_22152);
and U27214 (N_27214,N_20512,N_23396);
nor U27215 (N_27215,N_21220,N_21289);
or U27216 (N_27216,N_20632,N_22505);
nand U27217 (N_27217,N_20222,N_24308);
xor U27218 (N_27218,N_21164,N_22293);
nor U27219 (N_27219,N_21895,N_24334);
and U27220 (N_27220,N_20914,N_23064);
xor U27221 (N_27221,N_23996,N_22221);
and U27222 (N_27222,N_20711,N_24530);
xnor U27223 (N_27223,N_20848,N_24975);
and U27224 (N_27224,N_22685,N_20348);
nor U27225 (N_27225,N_23459,N_21331);
or U27226 (N_27226,N_21086,N_21052);
or U27227 (N_27227,N_22015,N_22919);
and U27228 (N_27228,N_23152,N_24697);
and U27229 (N_27229,N_22603,N_24849);
nor U27230 (N_27230,N_22908,N_22844);
nand U27231 (N_27231,N_20577,N_22874);
nand U27232 (N_27232,N_21446,N_20417);
nor U27233 (N_27233,N_23205,N_21328);
or U27234 (N_27234,N_22419,N_24703);
nand U27235 (N_27235,N_24893,N_20119);
nand U27236 (N_27236,N_21027,N_23026);
xnor U27237 (N_27237,N_23415,N_22724);
and U27238 (N_27238,N_20132,N_20090);
or U27239 (N_27239,N_23592,N_20687);
nor U27240 (N_27240,N_20103,N_23757);
and U27241 (N_27241,N_22490,N_24396);
nand U27242 (N_27242,N_21256,N_24381);
nor U27243 (N_27243,N_23149,N_21345);
xnor U27244 (N_27244,N_20877,N_23382);
nand U27245 (N_27245,N_21844,N_20078);
or U27246 (N_27246,N_21437,N_24079);
xor U27247 (N_27247,N_21700,N_20530);
or U27248 (N_27248,N_21729,N_24782);
or U27249 (N_27249,N_24000,N_24761);
nor U27250 (N_27250,N_22571,N_24613);
xnor U27251 (N_27251,N_21571,N_24689);
or U27252 (N_27252,N_23358,N_20718);
and U27253 (N_27253,N_22137,N_23186);
xor U27254 (N_27254,N_20672,N_24036);
and U27255 (N_27255,N_22966,N_22148);
xor U27256 (N_27256,N_24128,N_22259);
xnor U27257 (N_27257,N_20282,N_22836);
or U27258 (N_27258,N_24815,N_21056);
and U27259 (N_27259,N_23682,N_24720);
and U27260 (N_27260,N_20071,N_22133);
nor U27261 (N_27261,N_21202,N_20506);
and U27262 (N_27262,N_22569,N_21978);
and U27263 (N_27263,N_24970,N_22111);
or U27264 (N_27264,N_22659,N_21781);
and U27265 (N_27265,N_20826,N_22209);
or U27266 (N_27266,N_24940,N_23536);
xor U27267 (N_27267,N_20102,N_24654);
nor U27268 (N_27268,N_23005,N_21258);
xnor U27269 (N_27269,N_23138,N_23375);
or U27270 (N_27270,N_23416,N_20061);
nor U27271 (N_27271,N_20515,N_23111);
nand U27272 (N_27272,N_24635,N_21547);
or U27273 (N_27273,N_21520,N_23793);
nand U27274 (N_27274,N_20868,N_20027);
or U27275 (N_27275,N_22905,N_21369);
nand U27276 (N_27276,N_24526,N_24892);
or U27277 (N_27277,N_20875,N_22713);
nor U27278 (N_27278,N_23135,N_24180);
or U27279 (N_27279,N_21647,N_23526);
and U27280 (N_27280,N_24023,N_20118);
or U27281 (N_27281,N_24788,N_21850);
or U27282 (N_27282,N_23908,N_24681);
nand U27283 (N_27283,N_21668,N_20126);
and U27284 (N_27284,N_24053,N_21380);
nor U27285 (N_27285,N_21705,N_20849);
nor U27286 (N_27286,N_22883,N_21102);
nor U27287 (N_27287,N_24551,N_20135);
nor U27288 (N_27288,N_21276,N_23379);
or U27289 (N_27289,N_21209,N_21051);
nor U27290 (N_27290,N_23999,N_21851);
xnor U27291 (N_27291,N_22199,N_23532);
and U27292 (N_27292,N_23122,N_21832);
nor U27293 (N_27293,N_22926,N_20457);
xor U27294 (N_27294,N_20795,N_24833);
nand U27295 (N_27295,N_21559,N_24265);
nand U27296 (N_27296,N_20265,N_20154);
and U27297 (N_27297,N_22643,N_20660);
nand U27298 (N_27298,N_24015,N_20511);
and U27299 (N_27299,N_24182,N_23795);
xnor U27300 (N_27300,N_24736,N_21098);
and U27301 (N_27301,N_22690,N_21245);
nand U27302 (N_27302,N_23837,N_22592);
xor U27303 (N_27303,N_21440,N_24774);
and U27304 (N_27304,N_22046,N_24759);
xor U27305 (N_27305,N_21523,N_21135);
nor U27306 (N_27306,N_21661,N_21691);
nor U27307 (N_27307,N_20704,N_21181);
or U27308 (N_27308,N_21214,N_23567);
nand U27309 (N_27309,N_21384,N_24364);
xnor U27310 (N_27310,N_20714,N_20724);
or U27311 (N_27311,N_24044,N_22260);
xor U27312 (N_27312,N_22294,N_20657);
and U27313 (N_27313,N_23227,N_20026);
nor U27314 (N_27314,N_21943,N_22270);
and U27315 (N_27315,N_20031,N_21461);
xor U27316 (N_27316,N_21503,N_21783);
or U27317 (N_27317,N_24913,N_22090);
nand U27318 (N_27318,N_22456,N_22977);
nor U27319 (N_27319,N_24960,N_21286);
nor U27320 (N_27320,N_20558,N_21177);
or U27321 (N_27321,N_23082,N_20290);
and U27322 (N_27322,N_20435,N_21259);
or U27323 (N_27323,N_20792,N_24695);
and U27324 (N_27324,N_20441,N_20047);
and U27325 (N_27325,N_20991,N_22250);
or U27326 (N_27326,N_22455,N_22415);
nand U27327 (N_27327,N_23331,N_20709);
nand U27328 (N_27328,N_21100,N_21481);
or U27329 (N_27329,N_23255,N_21912);
or U27330 (N_27330,N_23665,N_21438);
nor U27331 (N_27331,N_22391,N_20419);
nand U27332 (N_27332,N_21420,N_22539);
nor U27333 (N_27333,N_22785,N_21324);
xnor U27334 (N_27334,N_23955,N_23591);
nand U27335 (N_27335,N_23830,N_23573);
and U27336 (N_27336,N_20609,N_22781);
nor U27337 (N_27337,N_20128,N_23395);
nor U27338 (N_27338,N_22063,N_20380);
and U27339 (N_27339,N_20912,N_23822);
or U27340 (N_27340,N_20560,N_23925);
xnor U27341 (N_27341,N_22331,N_21376);
nor U27342 (N_27342,N_22238,N_21335);
nor U27343 (N_27343,N_22161,N_23936);
and U27344 (N_27344,N_24608,N_22301);
nand U27345 (N_27345,N_22275,N_22408);
xor U27346 (N_27346,N_20502,N_24493);
or U27347 (N_27347,N_21877,N_21977);
or U27348 (N_27348,N_24047,N_21379);
and U27349 (N_27349,N_22360,N_22788);
xor U27350 (N_27350,N_20731,N_20451);
and U27351 (N_27351,N_20739,N_22348);
xnor U27352 (N_27352,N_23203,N_23013);
and U27353 (N_27353,N_24056,N_21113);
and U27354 (N_27354,N_21150,N_23563);
and U27355 (N_27355,N_20467,N_20147);
xnor U27356 (N_27356,N_23346,N_20862);
nor U27357 (N_27357,N_23389,N_21946);
and U27358 (N_27358,N_23730,N_23017);
nor U27359 (N_27359,N_23851,N_24442);
or U27360 (N_27360,N_20618,N_24032);
and U27361 (N_27361,N_21348,N_21223);
nand U27362 (N_27362,N_22255,N_23723);
xor U27363 (N_27363,N_22189,N_22003);
nor U27364 (N_27364,N_21477,N_22326);
nand U27365 (N_27365,N_24909,N_22988);
nor U27366 (N_27366,N_24915,N_23610);
nor U27367 (N_27367,N_22412,N_24742);
nor U27368 (N_27368,N_20234,N_24263);
xnor U27369 (N_27369,N_22318,N_24255);
and U27370 (N_27370,N_20279,N_20260);
or U27371 (N_27371,N_20999,N_22358);
nor U27372 (N_27372,N_20110,N_23750);
nor U27373 (N_27373,N_22931,N_22895);
or U27374 (N_27374,N_22095,N_20390);
and U27375 (N_27375,N_20493,N_21262);
xnor U27376 (N_27376,N_21196,N_21320);
or U27377 (N_27377,N_23391,N_20164);
or U27378 (N_27378,N_24851,N_24507);
and U27379 (N_27379,N_24682,N_23472);
or U27380 (N_27380,N_20592,N_20523);
and U27381 (N_27381,N_22672,N_23011);
and U27382 (N_27382,N_23163,N_22149);
nor U27383 (N_27383,N_20233,N_20363);
or U27384 (N_27384,N_20783,N_22637);
nor U27385 (N_27385,N_22092,N_21962);
or U27386 (N_27386,N_21537,N_21026);
or U27387 (N_27387,N_21055,N_22843);
xor U27388 (N_27388,N_21712,N_20851);
nand U27389 (N_27389,N_23729,N_23828);
xnor U27390 (N_27390,N_23347,N_22579);
nand U27391 (N_27391,N_24801,N_24946);
and U27392 (N_27392,N_20181,N_22745);
or U27393 (N_27393,N_22909,N_24039);
or U27394 (N_27394,N_21857,N_20648);
nand U27395 (N_27395,N_21395,N_24388);
nor U27396 (N_27396,N_21487,N_22177);
xnor U27397 (N_27397,N_24431,N_22519);
and U27398 (N_27398,N_23058,N_23125);
and U27399 (N_27399,N_20044,N_21131);
or U27400 (N_27400,N_23361,N_24130);
nand U27401 (N_27401,N_24165,N_20280);
or U27402 (N_27402,N_23569,N_20537);
xnor U27403 (N_27403,N_23191,N_21816);
nor U27404 (N_27404,N_20876,N_23398);
xor U27405 (N_27405,N_20686,N_20098);
nor U27406 (N_27406,N_24522,N_22548);
or U27407 (N_27407,N_23284,N_24415);
nand U27408 (N_27408,N_22129,N_23131);
or U27409 (N_27409,N_21969,N_23917);
and U27410 (N_27410,N_20017,N_20064);
and U27411 (N_27411,N_21063,N_24775);
or U27412 (N_27412,N_21064,N_21037);
nor U27413 (N_27413,N_23800,N_23374);
xnor U27414 (N_27414,N_20379,N_23662);
nand U27415 (N_27415,N_22778,N_23359);
nand U27416 (N_27416,N_21742,N_24747);
nor U27417 (N_27417,N_21759,N_20043);
and U27418 (N_27418,N_21319,N_20246);
nand U27419 (N_27419,N_22119,N_23376);
and U27420 (N_27420,N_24144,N_20913);
or U27421 (N_27421,N_22646,N_21412);
and U27422 (N_27422,N_24711,N_23294);
and U27423 (N_27423,N_21682,N_21082);
nand U27424 (N_27424,N_21624,N_20597);
or U27425 (N_27425,N_22890,N_21840);
and U27426 (N_27426,N_20208,N_20598);
nand U27427 (N_27427,N_24339,N_22093);
xnor U27428 (N_27428,N_22376,N_20341);
or U27429 (N_27429,N_21492,N_24511);
xor U27430 (N_27430,N_22038,N_21992);
and U27431 (N_27431,N_22970,N_23264);
and U27432 (N_27432,N_23637,N_22715);
nor U27433 (N_27433,N_20366,N_24591);
nor U27434 (N_27434,N_21088,N_23695);
and U27435 (N_27435,N_22079,N_20151);
and U27436 (N_27436,N_20956,N_24794);
xnor U27437 (N_27437,N_23514,N_22121);
or U27438 (N_27438,N_21455,N_21934);
or U27439 (N_27439,N_22461,N_22803);
nand U27440 (N_27440,N_22998,N_22087);
and U27441 (N_27441,N_21779,N_20491);
or U27442 (N_27442,N_24239,N_23956);
nor U27443 (N_27443,N_21928,N_23958);
nand U27444 (N_27444,N_22600,N_21488);
nand U27445 (N_27445,N_22018,N_23091);
and U27446 (N_27446,N_20399,N_23160);
nor U27447 (N_27447,N_21567,N_24944);
and U27448 (N_27448,N_21119,N_21553);
and U27449 (N_27449,N_22355,N_21018);
and U27450 (N_27450,N_24674,N_22686);
and U27451 (N_27451,N_23323,N_24277);
and U27452 (N_27452,N_22814,N_23952);
xnor U27453 (N_27453,N_20866,N_24820);
xnor U27454 (N_27454,N_20878,N_23748);
and U27455 (N_27455,N_22349,N_21015);
nor U27456 (N_27456,N_24744,N_23413);
xnor U27457 (N_27457,N_20899,N_21999);
nand U27458 (N_27458,N_21507,N_23834);
nor U27459 (N_27459,N_24249,N_20199);
nand U27460 (N_27460,N_24572,N_21628);
xor U27461 (N_27461,N_24409,N_22567);
or U27462 (N_27462,N_23544,N_21751);
nand U27463 (N_27463,N_23045,N_24386);
nor U27464 (N_27464,N_22407,N_22787);
nor U27465 (N_27465,N_24516,N_24582);
nand U27466 (N_27466,N_24081,N_20397);
or U27467 (N_27467,N_21843,N_22362);
xnor U27468 (N_27468,N_20521,N_21147);
nand U27469 (N_27469,N_24690,N_20579);
or U27470 (N_27470,N_21762,N_21692);
or U27471 (N_27471,N_24437,N_23206);
nor U27472 (N_27472,N_23566,N_20488);
nand U27473 (N_27473,N_24418,N_22008);
or U27474 (N_27474,N_22925,N_22653);
xnor U27475 (N_27475,N_23700,N_23245);
nor U27476 (N_27476,N_20179,N_22437);
nor U27477 (N_27477,N_20170,N_21512);
xor U27478 (N_27478,N_22887,N_22387);
and U27479 (N_27479,N_20559,N_24223);
nand U27480 (N_27480,N_21409,N_21263);
nand U27481 (N_27481,N_22443,N_21506);
nor U27482 (N_27482,N_22268,N_22104);
and U27483 (N_27483,N_22635,N_22835);
or U27484 (N_27484,N_23238,N_23783);
or U27485 (N_27485,N_20834,N_22264);
xnor U27486 (N_27486,N_22956,N_20197);
nand U27487 (N_27487,N_20947,N_22957);
or U27488 (N_27488,N_22906,N_21907);
nand U27489 (N_27489,N_20769,N_21930);
nor U27490 (N_27490,N_24964,N_20268);
nor U27491 (N_27491,N_21939,N_21750);
and U27492 (N_27492,N_22425,N_22470);
nand U27493 (N_27493,N_24460,N_22371);
xor U27494 (N_27494,N_23121,N_24679);
and U27495 (N_27495,N_24100,N_22195);
xnor U27496 (N_27496,N_24698,N_24707);
nor U27497 (N_27497,N_21644,N_24914);
xnor U27498 (N_27498,N_24215,N_24347);
xnor U27499 (N_27499,N_21472,N_23350);
nor U27500 (N_27500,N_20163,N_23569);
xnor U27501 (N_27501,N_21819,N_22744);
xnor U27502 (N_27502,N_21342,N_23688);
xor U27503 (N_27503,N_22457,N_23380);
xnor U27504 (N_27504,N_24673,N_23280);
or U27505 (N_27505,N_21547,N_24538);
nor U27506 (N_27506,N_21129,N_24571);
or U27507 (N_27507,N_21864,N_22773);
xor U27508 (N_27508,N_23262,N_24839);
xnor U27509 (N_27509,N_23057,N_21820);
nor U27510 (N_27510,N_24497,N_23260);
nand U27511 (N_27511,N_20916,N_24533);
nor U27512 (N_27512,N_23116,N_20040);
xor U27513 (N_27513,N_24103,N_24741);
nor U27514 (N_27514,N_24285,N_20783);
xnor U27515 (N_27515,N_24178,N_21782);
nor U27516 (N_27516,N_24805,N_20666);
xor U27517 (N_27517,N_20775,N_21519);
nor U27518 (N_27518,N_22125,N_24882);
or U27519 (N_27519,N_20650,N_24362);
xnor U27520 (N_27520,N_20208,N_24671);
nor U27521 (N_27521,N_21125,N_22281);
xor U27522 (N_27522,N_24664,N_20607);
nor U27523 (N_27523,N_23336,N_24287);
nor U27524 (N_27524,N_22945,N_23721);
xnor U27525 (N_27525,N_21895,N_21362);
or U27526 (N_27526,N_20550,N_23684);
or U27527 (N_27527,N_20843,N_21418);
nor U27528 (N_27528,N_22350,N_24816);
xnor U27529 (N_27529,N_24443,N_23883);
and U27530 (N_27530,N_21186,N_22015);
nor U27531 (N_27531,N_22335,N_23387);
nor U27532 (N_27532,N_20672,N_22722);
or U27533 (N_27533,N_24401,N_20856);
xnor U27534 (N_27534,N_22051,N_24479);
and U27535 (N_27535,N_21129,N_22005);
or U27536 (N_27536,N_21260,N_22845);
or U27537 (N_27537,N_20188,N_21727);
nor U27538 (N_27538,N_22120,N_20675);
nand U27539 (N_27539,N_21715,N_24206);
or U27540 (N_27540,N_22043,N_21642);
and U27541 (N_27541,N_22621,N_21420);
nor U27542 (N_27542,N_20713,N_23213);
or U27543 (N_27543,N_23547,N_22291);
nand U27544 (N_27544,N_22025,N_21513);
or U27545 (N_27545,N_24940,N_23032);
or U27546 (N_27546,N_21100,N_21796);
nand U27547 (N_27547,N_24732,N_23073);
or U27548 (N_27548,N_22091,N_21187);
and U27549 (N_27549,N_20134,N_23026);
nor U27550 (N_27550,N_24113,N_24036);
nand U27551 (N_27551,N_24967,N_23580);
xnor U27552 (N_27552,N_20446,N_21204);
nand U27553 (N_27553,N_22577,N_23333);
and U27554 (N_27554,N_23660,N_20750);
and U27555 (N_27555,N_21733,N_24470);
and U27556 (N_27556,N_21997,N_20624);
xnor U27557 (N_27557,N_21441,N_20955);
xor U27558 (N_27558,N_24396,N_22745);
xor U27559 (N_27559,N_24253,N_22921);
xnor U27560 (N_27560,N_23868,N_20418);
or U27561 (N_27561,N_20451,N_20557);
xor U27562 (N_27562,N_20774,N_21097);
xnor U27563 (N_27563,N_20827,N_20395);
xor U27564 (N_27564,N_21133,N_22219);
or U27565 (N_27565,N_20555,N_23548);
xnor U27566 (N_27566,N_22858,N_23477);
or U27567 (N_27567,N_20379,N_23456);
nor U27568 (N_27568,N_23770,N_24191);
nand U27569 (N_27569,N_21036,N_24607);
and U27570 (N_27570,N_22435,N_20210);
nand U27571 (N_27571,N_20636,N_22648);
nor U27572 (N_27572,N_22541,N_20773);
and U27573 (N_27573,N_22279,N_20809);
xor U27574 (N_27574,N_24120,N_24714);
and U27575 (N_27575,N_22656,N_20296);
or U27576 (N_27576,N_24045,N_20602);
or U27577 (N_27577,N_23387,N_24536);
or U27578 (N_27578,N_20886,N_24787);
and U27579 (N_27579,N_20711,N_20029);
nor U27580 (N_27580,N_20241,N_20141);
nand U27581 (N_27581,N_22167,N_24380);
nor U27582 (N_27582,N_22585,N_24923);
xnor U27583 (N_27583,N_21811,N_21720);
nand U27584 (N_27584,N_23028,N_23352);
and U27585 (N_27585,N_20327,N_22150);
or U27586 (N_27586,N_21264,N_20542);
xnor U27587 (N_27587,N_22431,N_20156);
xor U27588 (N_27588,N_24152,N_24694);
and U27589 (N_27589,N_24187,N_23095);
nand U27590 (N_27590,N_24696,N_21200);
xnor U27591 (N_27591,N_20534,N_22642);
nand U27592 (N_27592,N_24265,N_21500);
xor U27593 (N_27593,N_22895,N_21221);
and U27594 (N_27594,N_22364,N_22737);
and U27595 (N_27595,N_21464,N_24127);
or U27596 (N_27596,N_20928,N_20286);
nand U27597 (N_27597,N_23477,N_20461);
or U27598 (N_27598,N_21657,N_24395);
nor U27599 (N_27599,N_22313,N_23249);
or U27600 (N_27600,N_23214,N_24658);
nand U27601 (N_27601,N_23346,N_24811);
or U27602 (N_27602,N_23796,N_20130);
nor U27603 (N_27603,N_23687,N_22565);
xor U27604 (N_27604,N_20428,N_20184);
and U27605 (N_27605,N_21767,N_24801);
xnor U27606 (N_27606,N_24446,N_23512);
nand U27607 (N_27607,N_23185,N_22240);
xnor U27608 (N_27608,N_22928,N_22395);
nand U27609 (N_27609,N_22127,N_20961);
xor U27610 (N_27610,N_20394,N_22059);
or U27611 (N_27611,N_22960,N_23815);
and U27612 (N_27612,N_20022,N_22671);
or U27613 (N_27613,N_24672,N_23051);
nor U27614 (N_27614,N_22102,N_24838);
xor U27615 (N_27615,N_21831,N_23488);
nor U27616 (N_27616,N_20999,N_23235);
xnor U27617 (N_27617,N_22268,N_23866);
nand U27618 (N_27618,N_22267,N_23080);
or U27619 (N_27619,N_23349,N_23216);
nand U27620 (N_27620,N_20088,N_23004);
or U27621 (N_27621,N_23918,N_22793);
xnor U27622 (N_27622,N_23566,N_24788);
xnor U27623 (N_27623,N_23602,N_21082);
nor U27624 (N_27624,N_22071,N_24314);
or U27625 (N_27625,N_22163,N_23415);
xnor U27626 (N_27626,N_24408,N_21873);
or U27627 (N_27627,N_21273,N_20744);
xnor U27628 (N_27628,N_23783,N_22753);
nor U27629 (N_27629,N_20574,N_22093);
or U27630 (N_27630,N_24932,N_22057);
nand U27631 (N_27631,N_23893,N_22770);
nor U27632 (N_27632,N_24999,N_22720);
nand U27633 (N_27633,N_22270,N_21443);
nand U27634 (N_27634,N_24755,N_20298);
xor U27635 (N_27635,N_24129,N_21618);
or U27636 (N_27636,N_21631,N_21763);
nor U27637 (N_27637,N_21595,N_22526);
nand U27638 (N_27638,N_23493,N_24886);
nor U27639 (N_27639,N_23190,N_22891);
xor U27640 (N_27640,N_23615,N_21757);
and U27641 (N_27641,N_22083,N_24804);
nor U27642 (N_27642,N_23490,N_21471);
nand U27643 (N_27643,N_22891,N_21605);
xor U27644 (N_27644,N_21132,N_23132);
and U27645 (N_27645,N_24209,N_20903);
and U27646 (N_27646,N_23451,N_20518);
nor U27647 (N_27647,N_22485,N_20901);
nand U27648 (N_27648,N_21080,N_24033);
or U27649 (N_27649,N_24471,N_22267);
and U27650 (N_27650,N_23443,N_24964);
nand U27651 (N_27651,N_23157,N_23694);
nand U27652 (N_27652,N_24066,N_22936);
nand U27653 (N_27653,N_23782,N_20648);
and U27654 (N_27654,N_23751,N_20904);
nand U27655 (N_27655,N_22465,N_20210);
nor U27656 (N_27656,N_24628,N_23910);
and U27657 (N_27657,N_22347,N_21708);
xor U27658 (N_27658,N_24635,N_20493);
and U27659 (N_27659,N_20807,N_21585);
or U27660 (N_27660,N_21164,N_24857);
and U27661 (N_27661,N_22115,N_22228);
nand U27662 (N_27662,N_22521,N_23352);
nor U27663 (N_27663,N_23244,N_22861);
and U27664 (N_27664,N_23494,N_22356);
xor U27665 (N_27665,N_22471,N_23281);
nor U27666 (N_27666,N_22714,N_23293);
nand U27667 (N_27667,N_22878,N_20093);
and U27668 (N_27668,N_24730,N_21444);
nand U27669 (N_27669,N_24031,N_20683);
xor U27670 (N_27670,N_24835,N_24291);
and U27671 (N_27671,N_20405,N_23589);
or U27672 (N_27672,N_20864,N_22383);
nand U27673 (N_27673,N_22031,N_20806);
nor U27674 (N_27674,N_21825,N_20915);
nor U27675 (N_27675,N_21518,N_20853);
or U27676 (N_27676,N_21898,N_21611);
nand U27677 (N_27677,N_20541,N_20858);
or U27678 (N_27678,N_24394,N_24895);
nor U27679 (N_27679,N_21859,N_21888);
xor U27680 (N_27680,N_24671,N_22210);
and U27681 (N_27681,N_21405,N_21178);
or U27682 (N_27682,N_20284,N_24122);
and U27683 (N_27683,N_20141,N_21456);
nand U27684 (N_27684,N_21429,N_22061);
xor U27685 (N_27685,N_24088,N_23481);
xnor U27686 (N_27686,N_21570,N_22535);
or U27687 (N_27687,N_23677,N_22786);
xnor U27688 (N_27688,N_24459,N_22409);
and U27689 (N_27689,N_22311,N_23046);
and U27690 (N_27690,N_23386,N_23098);
nand U27691 (N_27691,N_24088,N_24457);
xor U27692 (N_27692,N_20956,N_21004);
nor U27693 (N_27693,N_23834,N_21275);
nand U27694 (N_27694,N_22916,N_22144);
and U27695 (N_27695,N_21635,N_21870);
or U27696 (N_27696,N_22803,N_23489);
nand U27697 (N_27697,N_24359,N_24772);
nand U27698 (N_27698,N_22011,N_21962);
and U27699 (N_27699,N_22471,N_23956);
nand U27700 (N_27700,N_24101,N_22694);
nor U27701 (N_27701,N_23211,N_23903);
or U27702 (N_27702,N_20399,N_24300);
nor U27703 (N_27703,N_20363,N_23218);
and U27704 (N_27704,N_20478,N_20812);
xnor U27705 (N_27705,N_20213,N_23514);
and U27706 (N_27706,N_22022,N_22933);
xnor U27707 (N_27707,N_24630,N_23405);
and U27708 (N_27708,N_23828,N_23249);
and U27709 (N_27709,N_22069,N_22092);
and U27710 (N_27710,N_22049,N_23217);
and U27711 (N_27711,N_22805,N_24493);
or U27712 (N_27712,N_21114,N_21621);
nand U27713 (N_27713,N_24878,N_23973);
or U27714 (N_27714,N_24339,N_23868);
and U27715 (N_27715,N_20093,N_22635);
nor U27716 (N_27716,N_23405,N_23505);
nand U27717 (N_27717,N_23890,N_23707);
nor U27718 (N_27718,N_21195,N_21336);
nand U27719 (N_27719,N_22670,N_23217);
nand U27720 (N_27720,N_23757,N_20760);
nand U27721 (N_27721,N_21033,N_22614);
nand U27722 (N_27722,N_20170,N_22463);
nor U27723 (N_27723,N_24179,N_22262);
xnor U27724 (N_27724,N_21830,N_20397);
nor U27725 (N_27725,N_20831,N_21071);
and U27726 (N_27726,N_21746,N_23598);
xor U27727 (N_27727,N_24980,N_22381);
nand U27728 (N_27728,N_22978,N_21796);
nand U27729 (N_27729,N_22801,N_21730);
nand U27730 (N_27730,N_20404,N_23833);
and U27731 (N_27731,N_20508,N_24453);
nor U27732 (N_27732,N_22373,N_24119);
or U27733 (N_27733,N_21917,N_24296);
and U27734 (N_27734,N_24927,N_23294);
xor U27735 (N_27735,N_21328,N_24681);
nand U27736 (N_27736,N_20202,N_23714);
and U27737 (N_27737,N_21699,N_23231);
or U27738 (N_27738,N_22044,N_23947);
nand U27739 (N_27739,N_21471,N_22730);
and U27740 (N_27740,N_21372,N_21011);
nor U27741 (N_27741,N_20355,N_20498);
nand U27742 (N_27742,N_20239,N_22407);
nor U27743 (N_27743,N_23119,N_24551);
or U27744 (N_27744,N_22237,N_22592);
nor U27745 (N_27745,N_21449,N_20635);
and U27746 (N_27746,N_21493,N_20362);
or U27747 (N_27747,N_21935,N_23945);
nand U27748 (N_27748,N_21594,N_20027);
and U27749 (N_27749,N_20167,N_24731);
or U27750 (N_27750,N_21770,N_24370);
nor U27751 (N_27751,N_24894,N_24082);
nor U27752 (N_27752,N_20460,N_20215);
and U27753 (N_27753,N_22498,N_22118);
nor U27754 (N_27754,N_21029,N_22908);
xnor U27755 (N_27755,N_21826,N_23125);
nor U27756 (N_27756,N_20051,N_23580);
nor U27757 (N_27757,N_24052,N_21701);
nor U27758 (N_27758,N_23413,N_20473);
or U27759 (N_27759,N_24300,N_22669);
and U27760 (N_27760,N_20570,N_23282);
and U27761 (N_27761,N_24773,N_21945);
or U27762 (N_27762,N_21317,N_21893);
nor U27763 (N_27763,N_20478,N_22834);
xnor U27764 (N_27764,N_20264,N_22197);
nor U27765 (N_27765,N_21949,N_24065);
or U27766 (N_27766,N_20586,N_22855);
nand U27767 (N_27767,N_21102,N_22705);
or U27768 (N_27768,N_22674,N_21136);
and U27769 (N_27769,N_20863,N_20522);
or U27770 (N_27770,N_24195,N_24296);
or U27771 (N_27771,N_23528,N_20050);
or U27772 (N_27772,N_23972,N_24788);
and U27773 (N_27773,N_21109,N_22396);
xor U27774 (N_27774,N_21580,N_22158);
nand U27775 (N_27775,N_21773,N_21265);
nand U27776 (N_27776,N_20438,N_22775);
or U27777 (N_27777,N_23214,N_21549);
nand U27778 (N_27778,N_22520,N_22972);
xor U27779 (N_27779,N_23499,N_23052);
and U27780 (N_27780,N_20914,N_20457);
xor U27781 (N_27781,N_20874,N_21966);
nor U27782 (N_27782,N_21975,N_23853);
or U27783 (N_27783,N_24655,N_23135);
and U27784 (N_27784,N_23954,N_20522);
and U27785 (N_27785,N_22904,N_24402);
or U27786 (N_27786,N_23255,N_22135);
and U27787 (N_27787,N_20288,N_24330);
nand U27788 (N_27788,N_24853,N_23296);
xnor U27789 (N_27789,N_24149,N_20171);
or U27790 (N_27790,N_21541,N_20286);
nor U27791 (N_27791,N_20208,N_22190);
and U27792 (N_27792,N_20920,N_23368);
nor U27793 (N_27793,N_21368,N_21869);
nand U27794 (N_27794,N_23393,N_24350);
or U27795 (N_27795,N_24882,N_21274);
nand U27796 (N_27796,N_21840,N_20736);
or U27797 (N_27797,N_23926,N_24054);
nor U27798 (N_27798,N_20005,N_22202);
and U27799 (N_27799,N_20393,N_21446);
and U27800 (N_27800,N_24104,N_24017);
or U27801 (N_27801,N_22859,N_22138);
and U27802 (N_27802,N_21186,N_22622);
or U27803 (N_27803,N_23528,N_21202);
nor U27804 (N_27804,N_22180,N_20673);
nor U27805 (N_27805,N_23922,N_23748);
and U27806 (N_27806,N_23942,N_24946);
nor U27807 (N_27807,N_20634,N_24293);
nor U27808 (N_27808,N_22524,N_20740);
and U27809 (N_27809,N_24334,N_24837);
and U27810 (N_27810,N_21764,N_24671);
nand U27811 (N_27811,N_24448,N_24886);
or U27812 (N_27812,N_21239,N_20053);
and U27813 (N_27813,N_21459,N_21992);
and U27814 (N_27814,N_24733,N_24545);
or U27815 (N_27815,N_20250,N_24515);
nor U27816 (N_27816,N_22392,N_24270);
or U27817 (N_27817,N_22633,N_24909);
and U27818 (N_27818,N_24127,N_23924);
nand U27819 (N_27819,N_22031,N_23584);
xnor U27820 (N_27820,N_21923,N_23030);
or U27821 (N_27821,N_23709,N_24100);
nand U27822 (N_27822,N_23612,N_20186);
nor U27823 (N_27823,N_23950,N_24358);
nor U27824 (N_27824,N_24193,N_21416);
or U27825 (N_27825,N_22510,N_21887);
nor U27826 (N_27826,N_24511,N_24346);
or U27827 (N_27827,N_22160,N_20877);
nand U27828 (N_27828,N_20225,N_21443);
or U27829 (N_27829,N_22297,N_21354);
xor U27830 (N_27830,N_23068,N_21675);
and U27831 (N_27831,N_21420,N_24034);
xor U27832 (N_27832,N_20668,N_22754);
nand U27833 (N_27833,N_21096,N_21909);
nand U27834 (N_27834,N_24085,N_21967);
and U27835 (N_27835,N_20363,N_24283);
nand U27836 (N_27836,N_21429,N_22270);
nor U27837 (N_27837,N_21641,N_24303);
nand U27838 (N_27838,N_20577,N_24722);
nor U27839 (N_27839,N_21726,N_22229);
or U27840 (N_27840,N_22066,N_22095);
xnor U27841 (N_27841,N_20240,N_22895);
xnor U27842 (N_27842,N_22363,N_23112);
and U27843 (N_27843,N_23380,N_24065);
and U27844 (N_27844,N_21653,N_22949);
and U27845 (N_27845,N_20198,N_24556);
xor U27846 (N_27846,N_22810,N_20149);
xnor U27847 (N_27847,N_24410,N_23987);
nor U27848 (N_27848,N_20783,N_21821);
xor U27849 (N_27849,N_23609,N_22142);
and U27850 (N_27850,N_23142,N_23774);
xnor U27851 (N_27851,N_22521,N_23914);
nand U27852 (N_27852,N_24669,N_23715);
nor U27853 (N_27853,N_21683,N_21060);
xor U27854 (N_27854,N_22648,N_20838);
nor U27855 (N_27855,N_24034,N_23577);
or U27856 (N_27856,N_22206,N_21841);
nand U27857 (N_27857,N_24176,N_20368);
nor U27858 (N_27858,N_24881,N_24931);
or U27859 (N_27859,N_24185,N_20930);
nor U27860 (N_27860,N_24107,N_20067);
xnor U27861 (N_27861,N_21421,N_20227);
and U27862 (N_27862,N_23459,N_24486);
nor U27863 (N_27863,N_21595,N_24750);
nor U27864 (N_27864,N_22332,N_20577);
xnor U27865 (N_27865,N_22763,N_23838);
xor U27866 (N_27866,N_23996,N_23924);
and U27867 (N_27867,N_22105,N_23488);
nor U27868 (N_27868,N_24850,N_24580);
nand U27869 (N_27869,N_20092,N_23555);
xnor U27870 (N_27870,N_21017,N_20004);
nand U27871 (N_27871,N_22552,N_23529);
and U27872 (N_27872,N_23137,N_22666);
xor U27873 (N_27873,N_20626,N_21589);
nor U27874 (N_27874,N_24535,N_23551);
nor U27875 (N_27875,N_23436,N_20012);
and U27876 (N_27876,N_22010,N_23095);
nand U27877 (N_27877,N_21783,N_24354);
and U27878 (N_27878,N_23664,N_24880);
xor U27879 (N_27879,N_21441,N_23827);
xor U27880 (N_27880,N_20471,N_21789);
and U27881 (N_27881,N_20786,N_20928);
and U27882 (N_27882,N_21007,N_20749);
nor U27883 (N_27883,N_20013,N_23569);
xnor U27884 (N_27884,N_21406,N_22988);
nand U27885 (N_27885,N_20049,N_20384);
and U27886 (N_27886,N_22568,N_23606);
and U27887 (N_27887,N_20586,N_22966);
or U27888 (N_27888,N_20928,N_22855);
and U27889 (N_27889,N_23084,N_22637);
xnor U27890 (N_27890,N_20919,N_22347);
xnor U27891 (N_27891,N_24509,N_24999);
or U27892 (N_27892,N_23747,N_20021);
and U27893 (N_27893,N_22130,N_20292);
xor U27894 (N_27894,N_21487,N_20074);
nand U27895 (N_27895,N_22246,N_21003);
xnor U27896 (N_27896,N_23775,N_21675);
xnor U27897 (N_27897,N_23837,N_23527);
xor U27898 (N_27898,N_23987,N_21296);
xor U27899 (N_27899,N_23458,N_23415);
xnor U27900 (N_27900,N_20269,N_23350);
or U27901 (N_27901,N_23014,N_22648);
and U27902 (N_27902,N_21643,N_24633);
nand U27903 (N_27903,N_20626,N_23361);
or U27904 (N_27904,N_20326,N_22547);
xor U27905 (N_27905,N_22340,N_22889);
or U27906 (N_27906,N_22730,N_21190);
nor U27907 (N_27907,N_22905,N_24279);
nor U27908 (N_27908,N_22399,N_23256);
and U27909 (N_27909,N_23995,N_24197);
and U27910 (N_27910,N_24854,N_24603);
or U27911 (N_27911,N_22279,N_24360);
and U27912 (N_27912,N_24434,N_20346);
nand U27913 (N_27913,N_22040,N_23695);
nor U27914 (N_27914,N_22996,N_21772);
nand U27915 (N_27915,N_22857,N_20997);
nand U27916 (N_27916,N_20633,N_24085);
xnor U27917 (N_27917,N_22484,N_23919);
xor U27918 (N_27918,N_24803,N_23609);
nor U27919 (N_27919,N_22377,N_22440);
xnor U27920 (N_27920,N_20213,N_24166);
nor U27921 (N_27921,N_23488,N_24868);
or U27922 (N_27922,N_20343,N_24587);
and U27923 (N_27923,N_21565,N_20088);
nand U27924 (N_27924,N_24375,N_21037);
nor U27925 (N_27925,N_20329,N_23931);
or U27926 (N_27926,N_21801,N_23530);
xnor U27927 (N_27927,N_21450,N_23523);
or U27928 (N_27928,N_21729,N_21288);
nor U27929 (N_27929,N_20255,N_22924);
or U27930 (N_27930,N_24229,N_23664);
xnor U27931 (N_27931,N_20996,N_22672);
nor U27932 (N_27932,N_22976,N_21094);
or U27933 (N_27933,N_24099,N_20002);
nor U27934 (N_27934,N_23210,N_22810);
xnor U27935 (N_27935,N_21833,N_24939);
xor U27936 (N_27936,N_24976,N_22014);
or U27937 (N_27937,N_20595,N_22871);
xnor U27938 (N_27938,N_24206,N_23139);
or U27939 (N_27939,N_23102,N_22173);
xor U27940 (N_27940,N_21691,N_20450);
and U27941 (N_27941,N_20437,N_20208);
xor U27942 (N_27942,N_23579,N_20720);
xnor U27943 (N_27943,N_24875,N_23466);
nand U27944 (N_27944,N_22137,N_21225);
or U27945 (N_27945,N_20034,N_22438);
or U27946 (N_27946,N_21070,N_20821);
nand U27947 (N_27947,N_20579,N_22510);
or U27948 (N_27948,N_23598,N_20467);
nor U27949 (N_27949,N_22827,N_20857);
xnor U27950 (N_27950,N_24091,N_24279);
xor U27951 (N_27951,N_21900,N_20741);
or U27952 (N_27952,N_21980,N_23530);
nand U27953 (N_27953,N_22616,N_21971);
or U27954 (N_27954,N_22456,N_22967);
and U27955 (N_27955,N_21063,N_21104);
nand U27956 (N_27956,N_20986,N_24831);
xor U27957 (N_27957,N_22541,N_23384);
nand U27958 (N_27958,N_23758,N_20917);
xor U27959 (N_27959,N_21606,N_22882);
xnor U27960 (N_27960,N_23930,N_20567);
nand U27961 (N_27961,N_21513,N_24817);
xor U27962 (N_27962,N_20350,N_23766);
or U27963 (N_27963,N_21619,N_24118);
xor U27964 (N_27964,N_24724,N_24559);
or U27965 (N_27965,N_22065,N_20849);
nor U27966 (N_27966,N_20515,N_23125);
nor U27967 (N_27967,N_24167,N_21755);
nor U27968 (N_27968,N_24584,N_24868);
xnor U27969 (N_27969,N_24074,N_22992);
nor U27970 (N_27970,N_20050,N_22162);
or U27971 (N_27971,N_24140,N_20097);
or U27972 (N_27972,N_22072,N_23483);
nor U27973 (N_27973,N_24514,N_21717);
nand U27974 (N_27974,N_20757,N_21173);
nand U27975 (N_27975,N_22875,N_23537);
xor U27976 (N_27976,N_20624,N_22023);
xnor U27977 (N_27977,N_20456,N_23526);
or U27978 (N_27978,N_21254,N_23684);
or U27979 (N_27979,N_21328,N_23616);
nor U27980 (N_27980,N_23177,N_22589);
nand U27981 (N_27981,N_22214,N_22831);
nor U27982 (N_27982,N_21976,N_22181);
nor U27983 (N_27983,N_20551,N_22884);
nand U27984 (N_27984,N_20083,N_22415);
nor U27985 (N_27985,N_20807,N_22091);
nand U27986 (N_27986,N_23892,N_24998);
or U27987 (N_27987,N_23685,N_20446);
xor U27988 (N_27988,N_20424,N_24779);
and U27989 (N_27989,N_22444,N_20135);
or U27990 (N_27990,N_22691,N_20330);
xor U27991 (N_27991,N_22104,N_23565);
nor U27992 (N_27992,N_20547,N_21039);
nand U27993 (N_27993,N_21422,N_20613);
xnor U27994 (N_27994,N_20712,N_22730);
and U27995 (N_27995,N_20738,N_23978);
or U27996 (N_27996,N_20182,N_24301);
nor U27997 (N_27997,N_22188,N_21610);
and U27998 (N_27998,N_21286,N_22567);
xnor U27999 (N_27999,N_21856,N_21633);
and U28000 (N_28000,N_24050,N_22499);
xnor U28001 (N_28001,N_22198,N_20817);
nor U28002 (N_28002,N_21815,N_22120);
nand U28003 (N_28003,N_23074,N_23123);
nand U28004 (N_28004,N_22800,N_23431);
xor U28005 (N_28005,N_24669,N_22997);
nand U28006 (N_28006,N_22362,N_24398);
nand U28007 (N_28007,N_24295,N_24151);
nor U28008 (N_28008,N_21912,N_24913);
nand U28009 (N_28009,N_21068,N_23161);
nand U28010 (N_28010,N_23182,N_23218);
xor U28011 (N_28011,N_22727,N_21749);
or U28012 (N_28012,N_20272,N_23815);
and U28013 (N_28013,N_24689,N_21315);
or U28014 (N_28014,N_20719,N_21568);
nor U28015 (N_28015,N_24945,N_22716);
xnor U28016 (N_28016,N_24200,N_20641);
or U28017 (N_28017,N_20047,N_24424);
or U28018 (N_28018,N_21746,N_22322);
and U28019 (N_28019,N_22251,N_24964);
xnor U28020 (N_28020,N_21680,N_22006);
nand U28021 (N_28021,N_20451,N_24018);
nand U28022 (N_28022,N_24490,N_20878);
and U28023 (N_28023,N_24326,N_20112);
and U28024 (N_28024,N_22925,N_24237);
or U28025 (N_28025,N_24180,N_21768);
and U28026 (N_28026,N_24836,N_22519);
or U28027 (N_28027,N_21585,N_21015);
nand U28028 (N_28028,N_21777,N_21298);
or U28029 (N_28029,N_22837,N_21920);
nand U28030 (N_28030,N_22699,N_20273);
nor U28031 (N_28031,N_23423,N_21198);
nand U28032 (N_28032,N_23724,N_21717);
xor U28033 (N_28033,N_21888,N_23128);
nand U28034 (N_28034,N_24368,N_22294);
nor U28035 (N_28035,N_24841,N_23909);
and U28036 (N_28036,N_21146,N_24622);
nand U28037 (N_28037,N_24784,N_22789);
nor U28038 (N_28038,N_23885,N_21654);
nand U28039 (N_28039,N_20611,N_21464);
and U28040 (N_28040,N_22227,N_21681);
or U28041 (N_28041,N_20676,N_24876);
and U28042 (N_28042,N_22117,N_22797);
and U28043 (N_28043,N_22657,N_24834);
xor U28044 (N_28044,N_23264,N_21778);
or U28045 (N_28045,N_20013,N_21699);
and U28046 (N_28046,N_20994,N_23683);
and U28047 (N_28047,N_21981,N_23574);
and U28048 (N_28048,N_23061,N_23910);
nand U28049 (N_28049,N_22230,N_20954);
or U28050 (N_28050,N_20660,N_24376);
and U28051 (N_28051,N_20829,N_24433);
xor U28052 (N_28052,N_21551,N_22551);
nor U28053 (N_28053,N_22601,N_24095);
xor U28054 (N_28054,N_24323,N_21379);
or U28055 (N_28055,N_20539,N_22380);
xnor U28056 (N_28056,N_20966,N_24847);
nand U28057 (N_28057,N_24029,N_24817);
nor U28058 (N_28058,N_21204,N_23692);
and U28059 (N_28059,N_22962,N_21729);
or U28060 (N_28060,N_22756,N_20096);
nor U28061 (N_28061,N_20705,N_24004);
and U28062 (N_28062,N_21770,N_21383);
nand U28063 (N_28063,N_22235,N_23573);
and U28064 (N_28064,N_24522,N_20583);
and U28065 (N_28065,N_20134,N_22032);
or U28066 (N_28066,N_21866,N_22950);
nor U28067 (N_28067,N_24293,N_22221);
or U28068 (N_28068,N_24583,N_24383);
nand U28069 (N_28069,N_24288,N_20626);
and U28070 (N_28070,N_24634,N_20087);
or U28071 (N_28071,N_21029,N_22315);
and U28072 (N_28072,N_23519,N_20831);
or U28073 (N_28073,N_22408,N_23283);
nand U28074 (N_28074,N_24149,N_22631);
xnor U28075 (N_28075,N_20619,N_22973);
xor U28076 (N_28076,N_22166,N_20206);
xor U28077 (N_28077,N_21931,N_21727);
xnor U28078 (N_28078,N_22593,N_22924);
xnor U28079 (N_28079,N_24165,N_23229);
nand U28080 (N_28080,N_21032,N_24930);
or U28081 (N_28081,N_20841,N_23535);
or U28082 (N_28082,N_24351,N_22102);
nor U28083 (N_28083,N_24143,N_23895);
nor U28084 (N_28084,N_22609,N_20504);
nand U28085 (N_28085,N_21719,N_23469);
xnor U28086 (N_28086,N_20892,N_24116);
xnor U28087 (N_28087,N_24834,N_23225);
nor U28088 (N_28088,N_24936,N_22679);
nor U28089 (N_28089,N_21836,N_22804);
nand U28090 (N_28090,N_21574,N_20360);
nand U28091 (N_28091,N_21859,N_23506);
nand U28092 (N_28092,N_22685,N_22511);
or U28093 (N_28093,N_23269,N_21350);
or U28094 (N_28094,N_24023,N_20049);
or U28095 (N_28095,N_24362,N_23299);
nor U28096 (N_28096,N_21632,N_24669);
xor U28097 (N_28097,N_20234,N_21484);
nand U28098 (N_28098,N_22412,N_22954);
and U28099 (N_28099,N_23635,N_23742);
nand U28100 (N_28100,N_23961,N_24660);
or U28101 (N_28101,N_22053,N_23129);
nor U28102 (N_28102,N_23401,N_24302);
nand U28103 (N_28103,N_22084,N_24092);
nor U28104 (N_28104,N_22018,N_24926);
nor U28105 (N_28105,N_20754,N_20212);
and U28106 (N_28106,N_24639,N_23296);
nand U28107 (N_28107,N_21734,N_22189);
nor U28108 (N_28108,N_23057,N_23493);
xnor U28109 (N_28109,N_22280,N_21018);
nand U28110 (N_28110,N_20920,N_24100);
and U28111 (N_28111,N_20356,N_24907);
or U28112 (N_28112,N_24871,N_24074);
and U28113 (N_28113,N_20045,N_23956);
nand U28114 (N_28114,N_20877,N_20649);
or U28115 (N_28115,N_21642,N_20419);
nor U28116 (N_28116,N_20226,N_22483);
and U28117 (N_28117,N_21836,N_22684);
and U28118 (N_28118,N_23426,N_23482);
or U28119 (N_28119,N_24643,N_22913);
nor U28120 (N_28120,N_20444,N_24207);
and U28121 (N_28121,N_21650,N_22935);
nor U28122 (N_28122,N_22211,N_20522);
nand U28123 (N_28123,N_23053,N_24044);
xnor U28124 (N_28124,N_22091,N_22712);
nor U28125 (N_28125,N_20678,N_23957);
or U28126 (N_28126,N_20573,N_23266);
and U28127 (N_28127,N_23988,N_23889);
and U28128 (N_28128,N_24860,N_22428);
xor U28129 (N_28129,N_22243,N_24394);
nand U28130 (N_28130,N_24969,N_21990);
nand U28131 (N_28131,N_22715,N_24417);
xor U28132 (N_28132,N_21311,N_21320);
and U28133 (N_28133,N_23809,N_24762);
and U28134 (N_28134,N_24452,N_20336);
nor U28135 (N_28135,N_22899,N_22789);
and U28136 (N_28136,N_24688,N_22531);
and U28137 (N_28137,N_21079,N_21772);
or U28138 (N_28138,N_24571,N_24507);
and U28139 (N_28139,N_22833,N_22371);
nor U28140 (N_28140,N_22193,N_23677);
xor U28141 (N_28141,N_21474,N_20258);
nor U28142 (N_28142,N_22042,N_21067);
nand U28143 (N_28143,N_21912,N_21932);
and U28144 (N_28144,N_24754,N_21650);
nand U28145 (N_28145,N_21972,N_21558);
nand U28146 (N_28146,N_21149,N_24918);
or U28147 (N_28147,N_23685,N_22363);
nand U28148 (N_28148,N_22951,N_21719);
nand U28149 (N_28149,N_24162,N_24228);
or U28150 (N_28150,N_21592,N_24297);
nor U28151 (N_28151,N_23094,N_22275);
xor U28152 (N_28152,N_20654,N_23295);
and U28153 (N_28153,N_23826,N_23568);
nand U28154 (N_28154,N_22265,N_24144);
nor U28155 (N_28155,N_22048,N_24108);
nor U28156 (N_28156,N_22440,N_22131);
or U28157 (N_28157,N_20011,N_21983);
or U28158 (N_28158,N_21695,N_22520);
or U28159 (N_28159,N_24672,N_20362);
and U28160 (N_28160,N_24687,N_23632);
nor U28161 (N_28161,N_22819,N_21719);
and U28162 (N_28162,N_21842,N_23516);
xor U28163 (N_28163,N_22452,N_20845);
and U28164 (N_28164,N_20803,N_21820);
or U28165 (N_28165,N_21980,N_20294);
or U28166 (N_28166,N_23411,N_22602);
xor U28167 (N_28167,N_24360,N_24142);
or U28168 (N_28168,N_23574,N_22609);
and U28169 (N_28169,N_21792,N_21842);
and U28170 (N_28170,N_21885,N_20706);
nand U28171 (N_28171,N_20143,N_22083);
xnor U28172 (N_28172,N_23038,N_23828);
or U28173 (N_28173,N_21315,N_23745);
nor U28174 (N_28174,N_22100,N_24728);
nand U28175 (N_28175,N_20088,N_24867);
xor U28176 (N_28176,N_24231,N_20140);
xnor U28177 (N_28177,N_23094,N_24482);
xnor U28178 (N_28178,N_22989,N_21889);
or U28179 (N_28179,N_24055,N_20367);
nand U28180 (N_28180,N_20769,N_23565);
or U28181 (N_28181,N_21401,N_20116);
and U28182 (N_28182,N_21545,N_21200);
xor U28183 (N_28183,N_22494,N_23354);
nand U28184 (N_28184,N_24896,N_24216);
xor U28185 (N_28185,N_20435,N_20824);
nand U28186 (N_28186,N_20410,N_23331);
xor U28187 (N_28187,N_20602,N_21013);
nand U28188 (N_28188,N_22721,N_20044);
and U28189 (N_28189,N_21000,N_24033);
nand U28190 (N_28190,N_21048,N_20187);
and U28191 (N_28191,N_24419,N_20875);
nor U28192 (N_28192,N_23110,N_22958);
or U28193 (N_28193,N_22082,N_23004);
or U28194 (N_28194,N_24372,N_20989);
and U28195 (N_28195,N_23948,N_21202);
xor U28196 (N_28196,N_22065,N_22072);
nor U28197 (N_28197,N_24534,N_23231);
xnor U28198 (N_28198,N_20579,N_24107);
xor U28199 (N_28199,N_22053,N_22065);
and U28200 (N_28200,N_24439,N_23997);
nor U28201 (N_28201,N_21425,N_21315);
xnor U28202 (N_28202,N_24691,N_20777);
nor U28203 (N_28203,N_22674,N_22060);
nor U28204 (N_28204,N_21409,N_24372);
xor U28205 (N_28205,N_21806,N_24162);
and U28206 (N_28206,N_23890,N_21553);
nand U28207 (N_28207,N_22361,N_22127);
nand U28208 (N_28208,N_22350,N_20167);
and U28209 (N_28209,N_20536,N_20685);
or U28210 (N_28210,N_23707,N_23967);
nand U28211 (N_28211,N_22032,N_22673);
xor U28212 (N_28212,N_20193,N_22573);
nor U28213 (N_28213,N_21041,N_22125);
nor U28214 (N_28214,N_21487,N_20760);
and U28215 (N_28215,N_23848,N_24981);
nor U28216 (N_28216,N_24923,N_24740);
and U28217 (N_28217,N_20101,N_21327);
and U28218 (N_28218,N_24813,N_20187);
xnor U28219 (N_28219,N_20238,N_22345);
nor U28220 (N_28220,N_20263,N_24481);
and U28221 (N_28221,N_20131,N_20921);
and U28222 (N_28222,N_20191,N_23408);
and U28223 (N_28223,N_21779,N_22664);
xor U28224 (N_28224,N_22313,N_23934);
nand U28225 (N_28225,N_20640,N_21111);
or U28226 (N_28226,N_24968,N_20453);
and U28227 (N_28227,N_20676,N_23721);
xnor U28228 (N_28228,N_24406,N_24310);
nand U28229 (N_28229,N_20375,N_23052);
and U28230 (N_28230,N_21209,N_20158);
xor U28231 (N_28231,N_22861,N_24174);
nor U28232 (N_28232,N_24322,N_20758);
and U28233 (N_28233,N_24754,N_24304);
and U28234 (N_28234,N_22221,N_22359);
and U28235 (N_28235,N_21350,N_22224);
and U28236 (N_28236,N_24515,N_23932);
nor U28237 (N_28237,N_23324,N_20575);
nand U28238 (N_28238,N_22688,N_21357);
xnor U28239 (N_28239,N_23727,N_22038);
nor U28240 (N_28240,N_21905,N_23819);
xnor U28241 (N_28241,N_24281,N_20134);
and U28242 (N_28242,N_21920,N_22857);
and U28243 (N_28243,N_24453,N_21511);
xnor U28244 (N_28244,N_22064,N_24905);
xor U28245 (N_28245,N_23805,N_24014);
or U28246 (N_28246,N_21455,N_21747);
or U28247 (N_28247,N_21899,N_22915);
nand U28248 (N_28248,N_22992,N_23982);
nor U28249 (N_28249,N_21461,N_20943);
nand U28250 (N_28250,N_22903,N_22600);
xnor U28251 (N_28251,N_24550,N_21947);
and U28252 (N_28252,N_20130,N_23119);
nor U28253 (N_28253,N_21046,N_23609);
nor U28254 (N_28254,N_20551,N_22552);
nor U28255 (N_28255,N_21025,N_21856);
nor U28256 (N_28256,N_24074,N_24697);
xnor U28257 (N_28257,N_22740,N_24590);
or U28258 (N_28258,N_24560,N_24389);
and U28259 (N_28259,N_20226,N_20901);
and U28260 (N_28260,N_23087,N_20437);
nor U28261 (N_28261,N_21619,N_20718);
nor U28262 (N_28262,N_24265,N_24448);
and U28263 (N_28263,N_23354,N_21753);
nand U28264 (N_28264,N_24962,N_22617);
and U28265 (N_28265,N_20571,N_24206);
xor U28266 (N_28266,N_22667,N_24863);
nor U28267 (N_28267,N_22098,N_20742);
nand U28268 (N_28268,N_20367,N_21102);
xnor U28269 (N_28269,N_22901,N_24490);
or U28270 (N_28270,N_20428,N_24966);
nand U28271 (N_28271,N_24797,N_22121);
or U28272 (N_28272,N_20182,N_23988);
and U28273 (N_28273,N_22634,N_21110);
or U28274 (N_28274,N_21100,N_23788);
nand U28275 (N_28275,N_21479,N_23177);
and U28276 (N_28276,N_21201,N_24224);
nor U28277 (N_28277,N_20349,N_20273);
or U28278 (N_28278,N_20311,N_20412);
xor U28279 (N_28279,N_23253,N_20376);
or U28280 (N_28280,N_22684,N_23704);
nor U28281 (N_28281,N_22757,N_23831);
and U28282 (N_28282,N_23641,N_24260);
nor U28283 (N_28283,N_20376,N_22373);
or U28284 (N_28284,N_21448,N_23331);
or U28285 (N_28285,N_22847,N_23949);
and U28286 (N_28286,N_24765,N_23616);
xor U28287 (N_28287,N_20325,N_20735);
and U28288 (N_28288,N_24894,N_21926);
nand U28289 (N_28289,N_20150,N_23667);
nor U28290 (N_28290,N_20873,N_24363);
and U28291 (N_28291,N_21051,N_23772);
nand U28292 (N_28292,N_22643,N_23968);
nor U28293 (N_28293,N_23519,N_23786);
or U28294 (N_28294,N_21994,N_23354);
or U28295 (N_28295,N_22397,N_24564);
nor U28296 (N_28296,N_23674,N_22004);
nand U28297 (N_28297,N_22063,N_23456);
or U28298 (N_28298,N_23972,N_20123);
and U28299 (N_28299,N_20284,N_22106);
and U28300 (N_28300,N_21000,N_20700);
nor U28301 (N_28301,N_21710,N_21321);
or U28302 (N_28302,N_21295,N_22787);
nor U28303 (N_28303,N_20233,N_24352);
and U28304 (N_28304,N_20860,N_22799);
and U28305 (N_28305,N_20461,N_23814);
nor U28306 (N_28306,N_23244,N_21898);
xor U28307 (N_28307,N_23631,N_24509);
nor U28308 (N_28308,N_22568,N_20289);
and U28309 (N_28309,N_20675,N_24534);
nor U28310 (N_28310,N_24433,N_23684);
or U28311 (N_28311,N_21581,N_23788);
xnor U28312 (N_28312,N_24509,N_22513);
or U28313 (N_28313,N_22425,N_22797);
or U28314 (N_28314,N_22395,N_23341);
nor U28315 (N_28315,N_22597,N_24450);
nor U28316 (N_28316,N_20545,N_23741);
nor U28317 (N_28317,N_21854,N_22384);
nor U28318 (N_28318,N_20760,N_23279);
and U28319 (N_28319,N_24482,N_20868);
nor U28320 (N_28320,N_21912,N_23589);
nor U28321 (N_28321,N_22408,N_20823);
nand U28322 (N_28322,N_22291,N_24143);
or U28323 (N_28323,N_20518,N_20131);
and U28324 (N_28324,N_22489,N_22803);
or U28325 (N_28325,N_21127,N_24867);
nor U28326 (N_28326,N_22937,N_24625);
and U28327 (N_28327,N_20737,N_23350);
or U28328 (N_28328,N_22993,N_23004);
xor U28329 (N_28329,N_20030,N_24178);
and U28330 (N_28330,N_21852,N_21834);
or U28331 (N_28331,N_23331,N_21228);
xnor U28332 (N_28332,N_24299,N_20819);
xnor U28333 (N_28333,N_21255,N_23394);
xnor U28334 (N_28334,N_22481,N_20023);
xnor U28335 (N_28335,N_21912,N_21778);
nor U28336 (N_28336,N_21472,N_21422);
and U28337 (N_28337,N_23667,N_24582);
and U28338 (N_28338,N_22288,N_21021);
nand U28339 (N_28339,N_23528,N_24835);
nand U28340 (N_28340,N_24314,N_22286);
nor U28341 (N_28341,N_21353,N_20404);
or U28342 (N_28342,N_20473,N_22684);
or U28343 (N_28343,N_20452,N_21201);
nor U28344 (N_28344,N_20265,N_23745);
xor U28345 (N_28345,N_22825,N_22347);
nor U28346 (N_28346,N_23265,N_23279);
and U28347 (N_28347,N_24725,N_22062);
nor U28348 (N_28348,N_23481,N_23769);
nand U28349 (N_28349,N_22326,N_21605);
xnor U28350 (N_28350,N_24933,N_24160);
nand U28351 (N_28351,N_22827,N_22994);
and U28352 (N_28352,N_20654,N_24243);
xnor U28353 (N_28353,N_24098,N_21532);
xor U28354 (N_28354,N_23058,N_23488);
nand U28355 (N_28355,N_23522,N_20332);
and U28356 (N_28356,N_20228,N_23975);
or U28357 (N_28357,N_20542,N_22859);
and U28358 (N_28358,N_22760,N_20069);
or U28359 (N_28359,N_20445,N_21082);
xor U28360 (N_28360,N_24344,N_22847);
xnor U28361 (N_28361,N_23458,N_24719);
or U28362 (N_28362,N_22767,N_23987);
nand U28363 (N_28363,N_23689,N_24850);
nand U28364 (N_28364,N_20962,N_20545);
and U28365 (N_28365,N_20993,N_23712);
and U28366 (N_28366,N_20162,N_22727);
nand U28367 (N_28367,N_24576,N_24599);
nor U28368 (N_28368,N_24362,N_24784);
nor U28369 (N_28369,N_23683,N_23085);
nand U28370 (N_28370,N_24412,N_22302);
and U28371 (N_28371,N_20444,N_22078);
nor U28372 (N_28372,N_24058,N_23371);
and U28373 (N_28373,N_20881,N_21837);
nor U28374 (N_28374,N_24670,N_23082);
xor U28375 (N_28375,N_21491,N_22374);
and U28376 (N_28376,N_21869,N_22387);
or U28377 (N_28377,N_22811,N_20187);
nor U28378 (N_28378,N_22442,N_21518);
or U28379 (N_28379,N_22496,N_23475);
nor U28380 (N_28380,N_20385,N_21408);
and U28381 (N_28381,N_20002,N_20722);
and U28382 (N_28382,N_21240,N_24208);
nand U28383 (N_28383,N_21974,N_23529);
nand U28384 (N_28384,N_24222,N_20346);
xnor U28385 (N_28385,N_20275,N_21527);
and U28386 (N_28386,N_22784,N_21160);
nand U28387 (N_28387,N_24812,N_21952);
or U28388 (N_28388,N_24522,N_24814);
or U28389 (N_28389,N_22132,N_20195);
or U28390 (N_28390,N_22712,N_22276);
and U28391 (N_28391,N_23458,N_21178);
xnor U28392 (N_28392,N_20410,N_23962);
nor U28393 (N_28393,N_20030,N_23964);
nand U28394 (N_28394,N_24343,N_22873);
or U28395 (N_28395,N_23269,N_21452);
or U28396 (N_28396,N_21896,N_23122);
and U28397 (N_28397,N_24245,N_22519);
nor U28398 (N_28398,N_22896,N_22757);
or U28399 (N_28399,N_20751,N_22709);
and U28400 (N_28400,N_22173,N_24296);
xor U28401 (N_28401,N_20017,N_23354);
xor U28402 (N_28402,N_24240,N_23731);
or U28403 (N_28403,N_20846,N_24199);
nor U28404 (N_28404,N_20392,N_22059);
nor U28405 (N_28405,N_23031,N_20793);
and U28406 (N_28406,N_20395,N_23389);
nand U28407 (N_28407,N_20435,N_23289);
nand U28408 (N_28408,N_24384,N_24639);
nor U28409 (N_28409,N_20398,N_20858);
nor U28410 (N_28410,N_21258,N_22303);
or U28411 (N_28411,N_20112,N_21436);
and U28412 (N_28412,N_21045,N_20867);
nor U28413 (N_28413,N_22066,N_23053);
xor U28414 (N_28414,N_22090,N_20358);
and U28415 (N_28415,N_23513,N_23596);
nor U28416 (N_28416,N_20300,N_24682);
or U28417 (N_28417,N_21117,N_20767);
xor U28418 (N_28418,N_21174,N_23414);
and U28419 (N_28419,N_22149,N_20535);
and U28420 (N_28420,N_23889,N_20820);
xor U28421 (N_28421,N_24088,N_23197);
and U28422 (N_28422,N_21554,N_20702);
or U28423 (N_28423,N_20278,N_24031);
and U28424 (N_28424,N_22434,N_22314);
or U28425 (N_28425,N_24098,N_24216);
nand U28426 (N_28426,N_22929,N_21554);
and U28427 (N_28427,N_20949,N_23296);
and U28428 (N_28428,N_20084,N_23686);
xor U28429 (N_28429,N_22454,N_20355);
xnor U28430 (N_28430,N_23830,N_24292);
xnor U28431 (N_28431,N_20593,N_22849);
xnor U28432 (N_28432,N_24557,N_21516);
xor U28433 (N_28433,N_20071,N_22269);
and U28434 (N_28434,N_24726,N_24455);
xor U28435 (N_28435,N_21579,N_22913);
and U28436 (N_28436,N_22349,N_20179);
xor U28437 (N_28437,N_20070,N_22322);
or U28438 (N_28438,N_20268,N_21330);
and U28439 (N_28439,N_23356,N_21463);
nand U28440 (N_28440,N_24886,N_24417);
and U28441 (N_28441,N_23078,N_23510);
nand U28442 (N_28442,N_22395,N_21060);
nand U28443 (N_28443,N_22874,N_23012);
or U28444 (N_28444,N_23188,N_22844);
nor U28445 (N_28445,N_20463,N_23513);
nor U28446 (N_28446,N_22374,N_23629);
nor U28447 (N_28447,N_22553,N_22422);
xnor U28448 (N_28448,N_24956,N_21728);
xnor U28449 (N_28449,N_20342,N_24778);
nor U28450 (N_28450,N_21551,N_24753);
or U28451 (N_28451,N_23522,N_21409);
nor U28452 (N_28452,N_22656,N_20715);
and U28453 (N_28453,N_24189,N_24261);
nor U28454 (N_28454,N_24597,N_20661);
xnor U28455 (N_28455,N_21899,N_23083);
nor U28456 (N_28456,N_23902,N_21930);
and U28457 (N_28457,N_21826,N_22599);
or U28458 (N_28458,N_23458,N_23444);
and U28459 (N_28459,N_24937,N_23004);
nor U28460 (N_28460,N_23584,N_22604);
and U28461 (N_28461,N_21357,N_20145);
or U28462 (N_28462,N_24602,N_23196);
nor U28463 (N_28463,N_23843,N_22230);
or U28464 (N_28464,N_22668,N_24325);
xnor U28465 (N_28465,N_22906,N_24076);
xor U28466 (N_28466,N_21423,N_21412);
nor U28467 (N_28467,N_20334,N_22105);
nand U28468 (N_28468,N_20692,N_20171);
xnor U28469 (N_28469,N_21855,N_24635);
nor U28470 (N_28470,N_22339,N_23334);
xor U28471 (N_28471,N_24223,N_24210);
or U28472 (N_28472,N_21770,N_24591);
and U28473 (N_28473,N_24656,N_20742);
nand U28474 (N_28474,N_20834,N_21018);
xnor U28475 (N_28475,N_22982,N_22755);
xor U28476 (N_28476,N_21659,N_23039);
nand U28477 (N_28477,N_22497,N_23682);
or U28478 (N_28478,N_21070,N_21880);
and U28479 (N_28479,N_22297,N_23435);
nor U28480 (N_28480,N_23292,N_24162);
nand U28481 (N_28481,N_20931,N_20170);
and U28482 (N_28482,N_22983,N_21466);
nand U28483 (N_28483,N_20247,N_24049);
and U28484 (N_28484,N_24190,N_24100);
nand U28485 (N_28485,N_22910,N_21648);
and U28486 (N_28486,N_23511,N_24489);
nand U28487 (N_28487,N_23287,N_24576);
nand U28488 (N_28488,N_22846,N_20254);
and U28489 (N_28489,N_21116,N_21003);
nor U28490 (N_28490,N_24476,N_20248);
and U28491 (N_28491,N_21272,N_20765);
xnor U28492 (N_28492,N_24730,N_24591);
and U28493 (N_28493,N_23158,N_21864);
xor U28494 (N_28494,N_24061,N_24381);
and U28495 (N_28495,N_21038,N_21291);
and U28496 (N_28496,N_24869,N_20068);
nand U28497 (N_28497,N_23683,N_22123);
and U28498 (N_28498,N_22327,N_23046);
and U28499 (N_28499,N_24801,N_20144);
xnor U28500 (N_28500,N_24700,N_22398);
and U28501 (N_28501,N_22664,N_22029);
nand U28502 (N_28502,N_23109,N_23024);
nand U28503 (N_28503,N_20158,N_22732);
or U28504 (N_28504,N_24613,N_24244);
nand U28505 (N_28505,N_21563,N_20321);
xor U28506 (N_28506,N_21876,N_23609);
nand U28507 (N_28507,N_24548,N_21523);
xnor U28508 (N_28508,N_23117,N_22578);
xor U28509 (N_28509,N_24612,N_20401);
or U28510 (N_28510,N_20492,N_21773);
or U28511 (N_28511,N_21315,N_22464);
and U28512 (N_28512,N_23095,N_20936);
xor U28513 (N_28513,N_23469,N_24225);
nand U28514 (N_28514,N_24312,N_22879);
nor U28515 (N_28515,N_20145,N_23479);
and U28516 (N_28516,N_22311,N_24337);
nor U28517 (N_28517,N_21250,N_20904);
xnor U28518 (N_28518,N_23954,N_22940);
nor U28519 (N_28519,N_20551,N_20528);
nor U28520 (N_28520,N_21667,N_23072);
xor U28521 (N_28521,N_23995,N_22106);
nand U28522 (N_28522,N_20741,N_22347);
nand U28523 (N_28523,N_20652,N_22060);
and U28524 (N_28524,N_23860,N_21400);
xor U28525 (N_28525,N_22635,N_20548);
nor U28526 (N_28526,N_20979,N_21848);
nand U28527 (N_28527,N_23756,N_20693);
xnor U28528 (N_28528,N_20364,N_22443);
xor U28529 (N_28529,N_24975,N_20745);
or U28530 (N_28530,N_24868,N_23346);
nand U28531 (N_28531,N_22405,N_23592);
nor U28532 (N_28532,N_21303,N_21293);
nor U28533 (N_28533,N_20994,N_24560);
xor U28534 (N_28534,N_20927,N_21357);
or U28535 (N_28535,N_20432,N_22686);
xor U28536 (N_28536,N_20617,N_24835);
xor U28537 (N_28537,N_20224,N_23065);
nor U28538 (N_28538,N_22129,N_23949);
or U28539 (N_28539,N_24552,N_23994);
xor U28540 (N_28540,N_21067,N_24347);
nand U28541 (N_28541,N_21325,N_21178);
or U28542 (N_28542,N_22847,N_21480);
or U28543 (N_28543,N_22762,N_22318);
or U28544 (N_28544,N_20179,N_24934);
and U28545 (N_28545,N_23114,N_21199);
xnor U28546 (N_28546,N_24015,N_24800);
nor U28547 (N_28547,N_22424,N_20886);
nor U28548 (N_28548,N_22852,N_22258);
and U28549 (N_28549,N_24688,N_22247);
and U28550 (N_28550,N_22980,N_24865);
xnor U28551 (N_28551,N_22374,N_23281);
or U28552 (N_28552,N_21484,N_20135);
xnor U28553 (N_28553,N_23020,N_20229);
nor U28554 (N_28554,N_22856,N_23149);
nand U28555 (N_28555,N_21795,N_23755);
and U28556 (N_28556,N_23350,N_21850);
xor U28557 (N_28557,N_23232,N_20971);
nand U28558 (N_28558,N_23591,N_23575);
nand U28559 (N_28559,N_23479,N_23109);
or U28560 (N_28560,N_22850,N_21770);
nor U28561 (N_28561,N_21964,N_22226);
or U28562 (N_28562,N_22714,N_20467);
and U28563 (N_28563,N_22426,N_23272);
or U28564 (N_28564,N_24103,N_23069);
nor U28565 (N_28565,N_22357,N_23464);
or U28566 (N_28566,N_22741,N_21828);
or U28567 (N_28567,N_24439,N_21988);
nor U28568 (N_28568,N_24504,N_23641);
nand U28569 (N_28569,N_24863,N_20155);
xor U28570 (N_28570,N_23615,N_23696);
xor U28571 (N_28571,N_23700,N_24082);
or U28572 (N_28572,N_20569,N_21871);
nand U28573 (N_28573,N_24283,N_21898);
nand U28574 (N_28574,N_22907,N_22139);
nand U28575 (N_28575,N_20857,N_23240);
and U28576 (N_28576,N_23712,N_23959);
and U28577 (N_28577,N_22119,N_22648);
nor U28578 (N_28578,N_22360,N_21773);
xor U28579 (N_28579,N_20137,N_21793);
and U28580 (N_28580,N_23997,N_23670);
nand U28581 (N_28581,N_23114,N_20557);
and U28582 (N_28582,N_24973,N_22657);
and U28583 (N_28583,N_23861,N_20797);
xnor U28584 (N_28584,N_22266,N_23939);
and U28585 (N_28585,N_21488,N_21709);
nand U28586 (N_28586,N_21249,N_24828);
and U28587 (N_28587,N_24653,N_21920);
xnor U28588 (N_28588,N_21735,N_23726);
nor U28589 (N_28589,N_24683,N_21870);
nor U28590 (N_28590,N_23661,N_21020);
xor U28591 (N_28591,N_23626,N_23942);
xor U28592 (N_28592,N_20869,N_20214);
and U28593 (N_28593,N_23263,N_24756);
nand U28594 (N_28594,N_22813,N_21531);
or U28595 (N_28595,N_20590,N_21498);
nand U28596 (N_28596,N_20906,N_21189);
nor U28597 (N_28597,N_21001,N_20141);
and U28598 (N_28598,N_23821,N_24472);
xor U28599 (N_28599,N_23730,N_21386);
nor U28600 (N_28600,N_24642,N_24503);
nand U28601 (N_28601,N_22831,N_23944);
xor U28602 (N_28602,N_24469,N_23968);
nor U28603 (N_28603,N_24645,N_23585);
or U28604 (N_28604,N_21280,N_21106);
and U28605 (N_28605,N_20745,N_22806);
and U28606 (N_28606,N_24582,N_20865);
and U28607 (N_28607,N_20906,N_22954);
or U28608 (N_28608,N_23391,N_20552);
or U28609 (N_28609,N_23808,N_21713);
nand U28610 (N_28610,N_24781,N_24528);
and U28611 (N_28611,N_23746,N_21584);
nand U28612 (N_28612,N_24809,N_24420);
or U28613 (N_28613,N_22613,N_23683);
nand U28614 (N_28614,N_20198,N_20346);
and U28615 (N_28615,N_21338,N_21080);
and U28616 (N_28616,N_22327,N_24771);
nand U28617 (N_28617,N_22555,N_22805);
nand U28618 (N_28618,N_22482,N_22640);
nand U28619 (N_28619,N_21506,N_22392);
nand U28620 (N_28620,N_21686,N_23729);
nor U28621 (N_28621,N_23848,N_20458);
or U28622 (N_28622,N_22275,N_20102);
or U28623 (N_28623,N_22548,N_24091);
and U28624 (N_28624,N_21955,N_22726);
nand U28625 (N_28625,N_20798,N_24881);
or U28626 (N_28626,N_20437,N_20359);
and U28627 (N_28627,N_20906,N_24692);
or U28628 (N_28628,N_21285,N_24081);
and U28629 (N_28629,N_22473,N_22639);
xor U28630 (N_28630,N_21426,N_20668);
and U28631 (N_28631,N_22755,N_24590);
xnor U28632 (N_28632,N_23348,N_21398);
nand U28633 (N_28633,N_20729,N_24550);
and U28634 (N_28634,N_21828,N_20665);
or U28635 (N_28635,N_22747,N_20890);
nor U28636 (N_28636,N_20869,N_20797);
nand U28637 (N_28637,N_23712,N_23440);
nand U28638 (N_28638,N_23560,N_22183);
nor U28639 (N_28639,N_24612,N_20666);
xor U28640 (N_28640,N_22613,N_20458);
or U28641 (N_28641,N_23376,N_24237);
or U28642 (N_28642,N_23186,N_24325);
and U28643 (N_28643,N_22257,N_24779);
or U28644 (N_28644,N_21434,N_24248);
xnor U28645 (N_28645,N_21552,N_22149);
nor U28646 (N_28646,N_24110,N_24073);
or U28647 (N_28647,N_22348,N_20895);
nand U28648 (N_28648,N_23071,N_21265);
or U28649 (N_28649,N_21394,N_21537);
nor U28650 (N_28650,N_22569,N_20702);
xnor U28651 (N_28651,N_21143,N_22257);
and U28652 (N_28652,N_20186,N_23092);
and U28653 (N_28653,N_24484,N_22650);
xnor U28654 (N_28654,N_21205,N_21346);
nor U28655 (N_28655,N_24819,N_22063);
nand U28656 (N_28656,N_23857,N_24375);
xor U28657 (N_28657,N_22474,N_22734);
nand U28658 (N_28658,N_21339,N_20486);
nand U28659 (N_28659,N_22184,N_20352);
xor U28660 (N_28660,N_23579,N_22151);
or U28661 (N_28661,N_20866,N_23044);
xor U28662 (N_28662,N_20735,N_24722);
nand U28663 (N_28663,N_24439,N_20074);
and U28664 (N_28664,N_21069,N_24898);
and U28665 (N_28665,N_21622,N_23152);
or U28666 (N_28666,N_22819,N_20134);
and U28667 (N_28667,N_24058,N_23870);
nand U28668 (N_28668,N_24248,N_24057);
xor U28669 (N_28669,N_24845,N_23463);
nor U28670 (N_28670,N_24483,N_22224);
nor U28671 (N_28671,N_24564,N_23830);
nor U28672 (N_28672,N_20384,N_20348);
nand U28673 (N_28673,N_23908,N_20347);
and U28674 (N_28674,N_20097,N_20222);
nor U28675 (N_28675,N_24424,N_20255);
nor U28676 (N_28676,N_23778,N_24705);
or U28677 (N_28677,N_21321,N_23768);
nand U28678 (N_28678,N_24377,N_22161);
xnor U28679 (N_28679,N_20637,N_24897);
nand U28680 (N_28680,N_20600,N_20931);
or U28681 (N_28681,N_23517,N_24646);
nand U28682 (N_28682,N_21121,N_20349);
or U28683 (N_28683,N_24259,N_24062);
xnor U28684 (N_28684,N_23234,N_24523);
or U28685 (N_28685,N_21917,N_24477);
or U28686 (N_28686,N_20528,N_22221);
nor U28687 (N_28687,N_21012,N_20602);
nand U28688 (N_28688,N_22143,N_23614);
and U28689 (N_28689,N_24187,N_20923);
or U28690 (N_28690,N_22983,N_24991);
nor U28691 (N_28691,N_20976,N_23332);
nand U28692 (N_28692,N_22180,N_23867);
nor U28693 (N_28693,N_24422,N_21139);
and U28694 (N_28694,N_23909,N_20397);
or U28695 (N_28695,N_21222,N_22406);
and U28696 (N_28696,N_22809,N_20481);
and U28697 (N_28697,N_21022,N_24313);
or U28698 (N_28698,N_22523,N_21000);
and U28699 (N_28699,N_21625,N_21721);
xnor U28700 (N_28700,N_24783,N_22763);
xnor U28701 (N_28701,N_20994,N_23036);
nand U28702 (N_28702,N_20067,N_22044);
nor U28703 (N_28703,N_21921,N_22217);
nor U28704 (N_28704,N_20458,N_20976);
xor U28705 (N_28705,N_21316,N_21041);
and U28706 (N_28706,N_22861,N_21702);
nand U28707 (N_28707,N_20914,N_24543);
and U28708 (N_28708,N_21564,N_22549);
nor U28709 (N_28709,N_22238,N_23914);
and U28710 (N_28710,N_23096,N_21541);
nand U28711 (N_28711,N_23950,N_24934);
nor U28712 (N_28712,N_21102,N_24348);
and U28713 (N_28713,N_23407,N_23159);
nor U28714 (N_28714,N_21990,N_24724);
xnor U28715 (N_28715,N_24140,N_22461);
or U28716 (N_28716,N_24091,N_20792);
nor U28717 (N_28717,N_23172,N_20049);
nand U28718 (N_28718,N_24862,N_20462);
or U28719 (N_28719,N_21836,N_22735);
nor U28720 (N_28720,N_21560,N_24295);
nand U28721 (N_28721,N_23599,N_20651);
xor U28722 (N_28722,N_21611,N_21005);
or U28723 (N_28723,N_20045,N_22608);
nand U28724 (N_28724,N_20780,N_20093);
and U28725 (N_28725,N_20094,N_23099);
or U28726 (N_28726,N_24927,N_22388);
and U28727 (N_28727,N_24757,N_24548);
or U28728 (N_28728,N_23901,N_20634);
nand U28729 (N_28729,N_23863,N_20495);
or U28730 (N_28730,N_21455,N_23228);
or U28731 (N_28731,N_22478,N_23366);
nor U28732 (N_28732,N_24812,N_22202);
xnor U28733 (N_28733,N_21820,N_22178);
nand U28734 (N_28734,N_24718,N_24078);
and U28735 (N_28735,N_24044,N_21448);
xnor U28736 (N_28736,N_21739,N_24219);
nor U28737 (N_28737,N_21162,N_21700);
xnor U28738 (N_28738,N_23538,N_21997);
or U28739 (N_28739,N_23373,N_24557);
nand U28740 (N_28740,N_24962,N_22809);
nand U28741 (N_28741,N_24207,N_24430);
nand U28742 (N_28742,N_24915,N_20906);
nand U28743 (N_28743,N_22236,N_22423);
xnor U28744 (N_28744,N_22976,N_20660);
nand U28745 (N_28745,N_23007,N_24093);
xor U28746 (N_28746,N_21585,N_22054);
nand U28747 (N_28747,N_20774,N_22771);
nor U28748 (N_28748,N_24601,N_23937);
and U28749 (N_28749,N_24723,N_20471);
or U28750 (N_28750,N_23384,N_24986);
nand U28751 (N_28751,N_24241,N_21076);
xor U28752 (N_28752,N_20919,N_23704);
xnor U28753 (N_28753,N_22235,N_22551);
nand U28754 (N_28754,N_23436,N_24810);
or U28755 (N_28755,N_21095,N_20150);
nor U28756 (N_28756,N_24864,N_23439);
xor U28757 (N_28757,N_24313,N_24773);
or U28758 (N_28758,N_22345,N_21045);
nor U28759 (N_28759,N_24927,N_20056);
or U28760 (N_28760,N_22781,N_21735);
nand U28761 (N_28761,N_20353,N_24496);
xor U28762 (N_28762,N_23044,N_20522);
nor U28763 (N_28763,N_24633,N_23090);
nor U28764 (N_28764,N_24257,N_23854);
xnor U28765 (N_28765,N_21048,N_21619);
nor U28766 (N_28766,N_23411,N_24688);
xnor U28767 (N_28767,N_20511,N_21050);
nor U28768 (N_28768,N_21026,N_24144);
nand U28769 (N_28769,N_23745,N_22141);
and U28770 (N_28770,N_24644,N_24488);
and U28771 (N_28771,N_22575,N_20826);
and U28772 (N_28772,N_20770,N_21040);
or U28773 (N_28773,N_22479,N_23753);
nand U28774 (N_28774,N_24460,N_23406);
nor U28775 (N_28775,N_24062,N_21749);
nor U28776 (N_28776,N_22815,N_20175);
and U28777 (N_28777,N_24327,N_20350);
nor U28778 (N_28778,N_23844,N_20564);
xor U28779 (N_28779,N_24081,N_22251);
xor U28780 (N_28780,N_21980,N_20827);
nor U28781 (N_28781,N_20329,N_24014);
or U28782 (N_28782,N_21417,N_23690);
nand U28783 (N_28783,N_22814,N_24426);
nor U28784 (N_28784,N_21128,N_23640);
nor U28785 (N_28785,N_22053,N_22326);
nor U28786 (N_28786,N_23358,N_22816);
xor U28787 (N_28787,N_24414,N_24791);
and U28788 (N_28788,N_21905,N_21797);
xnor U28789 (N_28789,N_23416,N_23675);
and U28790 (N_28790,N_20268,N_20380);
and U28791 (N_28791,N_21186,N_24812);
or U28792 (N_28792,N_24672,N_22875);
nand U28793 (N_28793,N_21345,N_21263);
and U28794 (N_28794,N_21229,N_21103);
nand U28795 (N_28795,N_24169,N_21722);
xor U28796 (N_28796,N_22972,N_21829);
and U28797 (N_28797,N_20502,N_20355);
nor U28798 (N_28798,N_21982,N_20566);
xor U28799 (N_28799,N_23967,N_24254);
nor U28800 (N_28800,N_20210,N_23307);
or U28801 (N_28801,N_22747,N_24990);
nor U28802 (N_28802,N_22853,N_21457);
xor U28803 (N_28803,N_23557,N_22485);
nor U28804 (N_28804,N_23081,N_22321);
xnor U28805 (N_28805,N_23027,N_22169);
and U28806 (N_28806,N_24142,N_21019);
nand U28807 (N_28807,N_22032,N_24164);
or U28808 (N_28808,N_24760,N_20714);
xor U28809 (N_28809,N_22928,N_23399);
or U28810 (N_28810,N_21811,N_24404);
nor U28811 (N_28811,N_22782,N_20330);
nor U28812 (N_28812,N_21874,N_24294);
xor U28813 (N_28813,N_21680,N_22082);
xor U28814 (N_28814,N_20144,N_20951);
nand U28815 (N_28815,N_21144,N_22570);
nand U28816 (N_28816,N_22374,N_23191);
and U28817 (N_28817,N_21695,N_20620);
xor U28818 (N_28818,N_20432,N_24914);
and U28819 (N_28819,N_21664,N_20182);
xor U28820 (N_28820,N_23559,N_24949);
nor U28821 (N_28821,N_23287,N_21199);
nand U28822 (N_28822,N_23608,N_20963);
or U28823 (N_28823,N_23717,N_21113);
nor U28824 (N_28824,N_22337,N_22932);
and U28825 (N_28825,N_24244,N_23818);
nand U28826 (N_28826,N_22277,N_23925);
xnor U28827 (N_28827,N_23873,N_21094);
or U28828 (N_28828,N_23302,N_20221);
and U28829 (N_28829,N_23554,N_24019);
or U28830 (N_28830,N_24192,N_20183);
xor U28831 (N_28831,N_20049,N_23993);
xnor U28832 (N_28832,N_22827,N_23003);
xor U28833 (N_28833,N_24445,N_20642);
xor U28834 (N_28834,N_20364,N_22083);
or U28835 (N_28835,N_21690,N_22985);
and U28836 (N_28836,N_24329,N_23857);
and U28837 (N_28837,N_24948,N_20167);
nand U28838 (N_28838,N_21444,N_23120);
nand U28839 (N_28839,N_20983,N_20522);
or U28840 (N_28840,N_24003,N_24904);
nand U28841 (N_28841,N_24594,N_20157);
nand U28842 (N_28842,N_24857,N_20722);
nand U28843 (N_28843,N_24547,N_22798);
nor U28844 (N_28844,N_22121,N_24852);
xor U28845 (N_28845,N_20935,N_22301);
nand U28846 (N_28846,N_21749,N_24463);
xnor U28847 (N_28847,N_21794,N_23694);
and U28848 (N_28848,N_24690,N_20586);
or U28849 (N_28849,N_22448,N_24663);
or U28850 (N_28850,N_24367,N_23587);
xnor U28851 (N_28851,N_21528,N_20249);
or U28852 (N_28852,N_22809,N_22474);
nor U28853 (N_28853,N_24710,N_24655);
and U28854 (N_28854,N_22401,N_20719);
and U28855 (N_28855,N_24713,N_23778);
nand U28856 (N_28856,N_24050,N_20836);
xor U28857 (N_28857,N_20303,N_22526);
and U28858 (N_28858,N_22152,N_22914);
and U28859 (N_28859,N_20383,N_20703);
nand U28860 (N_28860,N_24335,N_21490);
or U28861 (N_28861,N_24114,N_20782);
and U28862 (N_28862,N_20700,N_21181);
xnor U28863 (N_28863,N_24834,N_24995);
xor U28864 (N_28864,N_20801,N_24604);
nand U28865 (N_28865,N_22493,N_20320);
nor U28866 (N_28866,N_24999,N_22451);
and U28867 (N_28867,N_23387,N_21593);
nand U28868 (N_28868,N_20679,N_20680);
xor U28869 (N_28869,N_23455,N_22955);
nand U28870 (N_28870,N_24102,N_22033);
and U28871 (N_28871,N_22542,N_22288);
and U28872 (N_28872,N_21001,N_22016);
xnor U28873 (N_28873,N_22526,N_23093);
and U28874 (N_28874,N_22709,N_22784);
nand U28875 (N_28875,N_23683,N_22814);
nand U28876 (N_28876,N_21916,N_21541);
nand U28877 (N_28877,N_23231,N_22854);
nand U28878 (N_28878,N_22490,N_23343);
nand U28879 (N_28879,N_24345,N_21912);
xnor U28880 (N_28880,N_20778,N_23435);
and U28881 (N_28881,N_21572,N_20339);
nor U28882 (N_28882,N_21302,N_24688);
xor U28883 (N_28883,N_20476,N_20726);
nor U28884 (N_28884,N_24506,N_23275);
or U28885 (N_28885,N_22813,N_24268);
or U28886 (N_28886,N_20843,N_22174);
or U28887 (N_28887,N_22492,N_20661);
xnor U28888 (N_28888,N_21019,N_24324);
xor U28889 (N_28889,N_22243,N_24278);
nand U28890 (N_28890,N_21498,N_23281);
or U28891 (N_28891,N_23860,N_23975);
xor U28892 (N_28892,N_21885,N_24779);
nor U28893 (N_28893,N_20575,N_22073);
and U28894 (N_28894,N_20306,N_21847);
xor U28895 (N_28895,N_21044,N_22822);
nor U28896 (N_28896,N_20785,N_20756);
or U28897 (N_28897,N_22227,N_21871);
nor U28898 (N_28898,N_24778,N_23499);
or U28899 (N_28899,N_20852,N_23527);
nor U28900 (N_28900,N_22608,N_24528);
and U28901 (N_28901,N_20508,N_23669);
nor U28902 (N_28902,N_23614,N_22760);
and U28903 (N_28903,N_22128,N_22282);
xor U28904 (N_28904,N_21489,N_24603);
nand U28905 (N_28905,N_23636,N_24036);
nand U28906 (N_28906,N_21037,N_20459);
or U28907 (N_28907,N_22813,N_23915);
and U28908 (N_28908,N_24349,N_22164);
nand U28909 (N_28909,N_21226,N_20994);
nand U28910 (N_28910,N_20259,N_22119);
xnor U28911 (N_28911,N_23067,N_22789);
nor U28912 (N_28912,N_23917,N_20104);
and U28913 (N_28913,N_20086,N_24255);
nor U28914 (N_28914,N_21408,N_20442);
or U28915 (N_28915,N_21163,N_21027);
or U28916 (N_28916,N_20631,N_23256);
and U28917 (N_28917,N_22855,N_24078);
xnor U28918 (N_28918,N_22842,N_21549);
nor U28919 (N_28919,N_23373,N_22009);
nor U28920 (N_28920,N_23626,N_22310);
xnor U28921 (N_28921,N_21590,N_22447);
or U28922 (N_28922,N_23285,N_23095);
and U28923 (N_28923,N_21482,N_23267);
nand U28924 (N_28924,N_21065,N_24240);
or U28925 (N_28925,N_21078,N_20211);
nand U28926 (N_28926,N_21119,N_21716);
nand U28927 (N_28927,N_24886,N_21618);
and U28928 (N_28928,N_23605,N_21507);
nor U28929 (N_28929,N_22858,N_24338);
and U28930 (N_28930,N_22342,N_22800);
xor U28931 (N_28931,N_22534,N_22711);
nor U28932 (N_28932,N_21360,N_20159);
or U28933 (N_28933,N_24795,N_20229);
nand U28934 (N_28934,N_21846,N_21157);
nor U28935 (N_28935,N_20016,N_23170);
nand U28936 (N_28936,N_20039,N_22513);
nand U28937 (N_28937,N_20979,N_23119);
xnor U28938 (N_28938,N_21936,N_21547);
xor U28939 (N_28939,N_20978,N_20859);
xor U28940 (N_28940,N_24913,N_24835);
and U28941 (N_28941,N_20753,N_21855);
xor U28942 (N_28942,N_24581,N_23308);
and U28943 (N_28943,N_24039,N_20768);
or U28944 (N_28944,N_22217,N_23738);
and U28945 (N_28945,N_24663,N_20873);
or U28946 (N_28946,N_24475,N_20935);
and U28947 (N_28947,N_22147,N_22405);
nor U28948 (N_28948,N_20883,N_24673);
nor U28949 (N_28949,N_23133,N_24824);
nor U28950 (N_28950,N_22837,N_21232);
nor U28951 (N_28951,N_22701,N_23227);
nor U28952 (N_28952,N_22557,N_24637);
and U28953 (N_28953,N_21261,N_24859);
and U28954 (N_28954,N_20461,N_20813);
xnor U28955 (N_28955,N_23173,N_24027);
xor U28956 (N_28956,N_22041,N_24211);
nor U28957 (N_28957,N_22813,N_24720);
nor U28958 (N_28958,N_20284,N_20192);
nor U28959 (N_28959,N_24529,N_23878);
and U28960 (N_28960,N_24069,N_21952);
nor U28961 (N_28961,N_21374,N_21372);
and U28962 (N_28962,N_21916,N_20449);
and U28963 (N_28963,N_22740,N_21131);
nor U28964 (N_28964,N_22157,N_22310);
and U28965 (N_28965,N_24735,N_21046);
and U28966 (N_28966,N_22605,N_23574);
or U28967 (N_28967,N_21452,N_22360);
or U28968 (N_28968,N_24497,N_22919);
xor U28969 (N_28969,N_21433,N_20444);
nor U28970 (N_28970,N_23232,N_24625);
and U28971 (N_28971,N_21243,N_23107);
xnor U28972 (N_28972,N_24943,N_23369);
nor U28973 (N_28973,N_20885,N_23623);
or U28974 (N_28974,N_23814,N_20363);
xnor U28975 (N_28975,N_20637,N_22854);
xor U28976 (N_28976,N_24927,N_20359);
xnor U28977 (N_28977,N_21704,N_21843);
xnor U28978 (N_28978,N_24712,N_22833);
or U28979 (N_28979,N_20364,N_23266);
and U28980 (N_28980,N_20443,N_24899);
xnor U28981 (N_28981,N_22741,N_21807);
or U28982 (N_28982,N_24362,N_22044);
or U28983 (N_28983,N_20411,N_23746);
nor U28984 (N_28984,N_20918,N_23269);
xor U28985 (N_28985,N_22295,N_22033);
xnor U28986 (N_28986,N_22627,N_24344);
nand U28987 (N_28987,N_20326,N_20971);
nor U28988 (N_28988,N_20345,N_21801);
nand U28989 (N_28989,N_22240,N_20965);
or U28990 (N_28990,N_22811,N_22177);
nand U28991 (N_28991,N_20278,N_24132);
or U28992 (N_28992,N_21302,N_21781);
nand U28993 (N_28993,N_23362,N_24970);
nor U28994 (N_28994,N_23313,N_24674);
and U28995 (N_28995,N_22664,N_21704);
nand U28996 (N_28996,N_20234,N_23698);
nor U28997 (N_28997,N_22930,N_22659);
nand U28998 (N_28998,N_23710,N_23788);
nand U28999 (N_28999,N_23428,N_22962);
xnor U29000 (N_29000,N_21313,N_22515);
and U29001 (N_29001,N_24279,N_21550);
xor U29002 (N_29002,N_23457,N_24319);
nor U29003 (N_29003,N_24020,N_20323);
nand U29004 (N_29004,N_23364,N_21228);
xnor U29005 (N_29005,N_20844,N_23947);
nand U29006 (N_29006,N_21061,N_24866);
xnor U29007 (N_29007,N_22345,N_22371);
or U29008 (N_29008,N_21856,N_21742);
nor U29009 (N_29009,N_21402,N_20612);
or U29010 (N_29010,N_24882,N_20437);
nand U29011 (N_29011,N_20366,N_24162);
nor U29012 (N_29012,N_20100,N_23218);
or U29013 (N_29013,N_24252,N_23687);
or U29014 (N_29014,N_23853,N_20868);
or U29015 (N_29015,N_21961,N_22756);
xnor U29016 (N_29016,N_24978,N_23870);
nand U29017 (N_29017,N_21048,N_23401);
nor U29018 (N_29018,N_20025,N_22550);
or U29019 (N_29019,N_20962,N_22078);
nand U29020 (N_29020,N_21142,N_24686);
and U29021 (N_29021,N_20000,N_20196);
or U29022 (N_29022,N_20623,N_22553);
xnor U29023 (N_29023,N_24423,N_24916);
xor U29024 (N_29024,N_23344,N_24095);
xor U29025 (N_29025,N_21546,N_24372);
xor U29026 (N_29026,N_20277,N_23269);
nor U29027 (N_29027,N_23548,N_21629);
nor U29028 (N_29028,N_23532,N_22810);
xor U29029 (N_29029,N_20385,N_21486);
nand U29030 (N_29030,N_24094,N_23536);
nor U29031 (N_29031,N_20319,N_21783);
nand U29032 (N_29032,N_21411,N_21712);
and U29033 (N_29033,N_24711,N_24823);
nand U29034 (N_29034,N_20994,N_24261);
xor U29035 (N_29035,N_23314,N_23111);
xor U29036 (N_29036,N_24638,N_23768);
nor U29037 (N_29037,N_21857,N_24720);
or U29038 (N_29038,N_23745,N_24145);
nor U29039 (N_29039,N_21423,N_22437);
nand U29040 (N_29040,N_23867,N_20097);
nand U29041 (N_29041,N_21024,N_22339);
xnor U29042 (N_29042,N_20219,N_21384);
nand U29043 (N_29043,N_21609,N_21703);
nor U29044 (N_29044,N_24221,N_20159);
nor U29045 (N_29045,N_23701,N_20956);
nor U29046 (N_29046,N_21364,N_22879);
nor U29047 (N_29047,N_24002,N_21363);
nand U29048 (N_29048,N_22560,N_24350);
or U29049 (N_29049,N_23116,N_24002);
xnor U29050 (N_29050,N_21661,N_23947);
nor U29051 (N_29051,N_24420,N_23101);
and U29052 (N_29052,N_21441,N_22949);
or U29053 (N_29053,N_23461,N_20065);
nand U29054 (N_29054,N_20080,N_23469);
nand U29055 (N_29055,N_22564,N_20096);
nor U29056 (N_29056,N_23372,N_24907);
and U29057 (N_29057,N_20314,N_21837);
xnor U29058 (N_29058,N_20904,N_24061);
and U29059 (N_29059,N_21668,N_20733);
or U29060 (N_29060,N_20235,N_22135);
xor U29061 (N_29061,N_20176,N_21640);
nor U29062 (N_29062,N_22443,N_24164);
xnor U29063 (N_29063,N_24292,N_22314);
nand U29064 (N_29064,N_24399,N_24812);
xor U29065 (N_29065,N_21890,N_22381);
nand U29066 (N_29066,N_22623,N_22817);
or U29067 (N_29067,N_23293,N_20260);
and U29068 (N_29068,N_21095,N_23417);
and U29069 (N_29069,N_20569,N_21227);
nand U29070 (N_29070,N_21230,N_22756);
nand U29071 (N_29071,N_21840,N_23920);
xor U29072 (N_29072,N_24847,N_24010);
xor U29073 (N_29073,N_23638,N_22551);
nor U29074 (N_29074,N_21965,N_20000);
or U29075 (N_29075,N_21655,N_21828);
nand U29076 (N_29076,N_24001,N_22722);
and U29077 (N_29077,N_21254,N_24321);
and U29078 (N_29078,N_23096,N_23032);
xor U29079 (N_29079,N_21616,N_23044);
nand U29080 (N_29080,N_20704,N_22240);
and U29081 (N_29081,N_20547,N_20798);
and U29082 (N_29082,N_20063,N_24808);
or U29083 (N_29083,N_23103,N_23111);
and U29084 (N_29084,N_23131,N_22961);
nand U29085 (N_29085,N_24601,N_22686);
and U29086 (N_29086,N_24285,N_23595);
nand U29087 (N_29087,N_24201,N_23380);
and U29088 (N_29088,N_20866,N_23553);
or U29089 (N_29089,N_20534,N_22325);
nor U29090 (N_29090,N_23843,N_23983);
and U29091 (N_29091,N_22237,N_24811);
nor U29092 (N_29092,N_23867,N_24303);
and U29093 (N_29093,N_24713,N_22525);
xor U29094 (N_29094,N_23124,N_21076);
nand U29095 (N_29095,N_21690,N_22446);
and U29096 (N_29096,N_21131,N_23549);
or U29097 (N_29097,N_22671,N_22782);
xor U29098 (N_29098,N_20437,N_21888);
nand U29099 (N_29099,N_21209,N_23078);
nand U29100 (N_29100,N_20590,N_24497);
nor U29101 (N_29101,N_20636,N_22729);
or U29102 (N_29102,N_21350,N_22254);
xor U29103 (N_29103,N_20035,N_20441);
and U29104 (N_29104,N_22523,N_21698);
or U29105 (N_29105,N_20235,N_22940);
nand U29106 (N_29106,N_24885,N_24905);
nor U29107 (N_29107,N_20907,N_20997);
or U29108 (N_29108,N_20044,N_20484);
nor U29109 (N_29109,N_22611,N_24182);
or U29110 (N_29110,N_24643,N_20492);
xor U29111 (N_29111,N_23994,N_21415);
or U29112 (N_29112,N_22719,N_20782);
nor U29113 (N_29113,N_24224,N_24263);
xnor U29114 (N_29114,N_21286,N_24060);
nor U29115 (N_29115,N_21562,N_23657);
nand U29116 (N_29116,N_22181,N_21953);
nor U29117 (N_29117,N_22263,N_24605);
and U29118 (N_29118,N_20686,N_20966);
xnor U29119 (N_29119,N_20489,N_21317);
or U29120 (N_29120,N_22852,N_24572);
xor U29121 (N_29121,N_24823,N_21669);
and U29122 (N_29122,N_20237,N_20258);
nor U29123 (N_29123,N_20657,N_24239);
nand U29124 (N_29124,N_22871,N_23176);
xnor U29125 (N_29125,N_20822,N_23043);
xnor U29126 (N_29126,N_24394,N_21541);
and U29127 (N_29127,N_20067,N_24425);
nor U29128 (N_29128,N_21298,N_22509);
nand U29129 (N_29129,N_22967,N_24255);
xnor U29130 (N_29130,N_20072,N_22690);
or U29131 (N_29131,N_20687,N_21461);
and U29132 (N_29132,N_23854,N_22189);
and U29133 (N_29133,N_22231,N_24208);
and U29134 (N_29134,N_20538,N_22023);
nor U29135 (N_29135,N_24748,N_23594);
xor U29136 (N_29136,N_21462,N_23551);
xor U29137 (N_29137,N_23610,N_24089);
nand U29138 (N_29138,N_20602,N_23036);
nor U29139 (N_29139,N_23272,N_24270);
nand U29140 (N_29140,N_20864,N_22477);
and U29141 (N_29141,N_20661,N_20690);
nand U29142 (N_29142,N_23240,N_24133);
and U29143 (N_29143,N_23460,N_22038);
or U29144 (N_29144,N_22778,N_20341);
xor U29145 (N_29145,N_22061,N_23122);
nand U29146 (N_29146,N_21389,N_20378);
or U29147 (N_29147,N_24861,N_24791);
xnor U29148 (N_29148,N_23756,N_21829);
nand U29149 (N_29149,N_23941,N_22101);
or U29150 (N_29150,N_21873,N_24265);
or U29151 (N_29151,N_21243,N_23512);
or U29152 (N_29152,N_20694,N_21185);
xnor U29153 (N_29153,N_22398,N_24480);
nand U29154 (N_29154,N_23722,N_24628);
and U29155 (N_29155,N_21555,N_24643);
and U29156 (N_29156,N_23203,N_21323);
xnor U29157 (N_29157,N_24591,N_23403);
xor U29158 (N_29158,N_24468,N_22757);
and U29159 (N_29159,N_24507,N_24665);
xnor U29160 (N_29160,N_21534,N_23802);
xnor U29161 (N_29161,N_24519,N_24660);
and U29162 (N_29162,N_21591,N_22914);
and U29163 (N_29163,N_23793,N_22380);
xor U29164 (N_29164,N_24879,N_23060);
and U29165 (N_29165,N_21564,N_20305);
and U29166 (N_29166,N_21361,N_20333);
nor U29167 (N_29167,N_24846,N_24309);
or U29168 (N_29168,N_21189,N_24963);
nand U29169 (N_29169,N_22962,N_21927);
or U29170 (N_29170,N_20285,N_21886);
and U29171 (N_29171,N_22774,N_23242);
or U29172 (N_29172,N_21899,N_23860);
nor U29173 (N_29173,N_20204,N_24911);
or U29174 (N_29174,N_20286,N_22302);
or U29175 (N_29175,N_20471,N_20143);
xnor U29176 (N_29176,N_24497,N_23627);
nor U29177 (N_29177,N_21347,N_22788);
and U29178 (N_29178,N_21903,N_21073);
xor U29179 (N_29179,N_21692,N_22345);
xor U29180 (N_29180,N_22996,N_20892);
or U29181 (N_29181,N_20587,N_21249);
xor U29182 (N_29182,N_22230,N_23059);
and U29183 (N_29183,N_23576,N_24475);
and U29184 (N_29184,N_22716,N_21813);
nand U29185 (N_29185,N_20710,N_20307);
nor U29186 (N_29186,N_23988,N_23860);
nand U29187 (N_29187,N_22685,N_23877);
nand U29188 (N_29188,N_22818,N_21116);
nand U29189 (N_29189,N_21902,N_24617);
xor U29190 (N_29190,N_22928,N_22742);
or U29191 (N_29191,N_24209,N_24808);
xnor U29192 (N_29192,N_20120,N_22307);
and U29193 (N_29193,N_21022,N_21784);
or U29194 (N_29194,N_20627,N_23672);
or U29195 (N_29195,N_20447,N_20522);
or U29196 (N_29196,N_22380,N_20059);
nor U29197 (N_29197,N_20506,N_20519);
xor U29198 (N_29198,N_22821,N_24931);
nand U29199 (N_29199,N_23942,N_22051);
nand U29200 (N_29200,N_23154,N_20344);
or U29201 (N_29201,N_24143,N_23655);
nor U29202 (N_29202,N_21468,N_21289);
xnor U29203 (N_29203,N_21194,N_20469);
nor U29204 (N_29204,N_24270,N_22337);
and U29205 (N_29205,N_24062,N_23617);
nand U29206 (N_29206,N_21311,N_21172);
nor U29207 (N_29207,N_20670,N_24844);
and U29208 (N_29208,N_21468,N_21502);
or U29209 (N_29209,N_20324,N_21371);
nor U29210 (N_29210,N_20765,N_22993);
xor U29211 (N_29211,N_22691,N_20282);
nor U29212 (N_29212,N_23651,N_20627);
and U29213 (N_29213,N_22539,N_20344);
nor U29214 (N_29214,N_23295,N_23868);
or U29215 (N_29215,N_23351,N_24836);
or U29216 (N_29216,N_22713,N_22374);
xnor U29217 (N_29217,N_22356,N_24123);
or U29218 (N_29218,N_24668,N_22829);
xnor U29219 (N_29219,N_24451,N_20743);
or U29220 (N_29220,N_23471,N_21494);
nand U29221 (N_29221,N_23835,N_24839);
or U29222 (N_29222,N_20883,N_22218);
and U29223 (N_29223,N_24070,N_22293);
nand U29224 (N_29224,N_21989,N_23409);
or U29225 (N_29225,N_24379,N_22640);
and U29226 (N_29226,N_22255,N_20413);
xnor U29227 (N_29227,N_23683,N_23255);
nand U29228 (N_29228,N_24502,N_20283);
or U29229 (N_29229,N_23272,N_22281);
nor U29230 (N_29230,N_21239,N_21578);
or U29231 (N_29231,N_23112,N_24530);
nor U29232 (N_29232,N_23282,N_23542);
nor U29233 (N_29233,N_23670,N_24310);
nand U29234 (N_29234,N_21112,N_21264);
nor U29235 (N_29235,N_24956,N_22465);
nor U29236 (N_29236,N_23361,N_22001);
xnor U29237 (N_29237,N_23845,N_20099);
nor U29238 (N_29238,N_22591,N_21910);
nor U29239 (N_29239,N_21525,N_22782);
xor U29240 (N_29240,N_22829,N_24328);
or U29241 (N_29241,N_20770,N_23227);
xor U29242 (N_29242,N_23823,N_22251);
nand U29243 (N_29243,N_23178,N_24021);
xor U29244 (N_29244,N_21015,N_24207);
and U29245 (N_29245,N_24235,N_24189);
nand U29246 (N_29246,N_24785,N_24221);
and U29247 (N_29247,N_23385,N_20348);
xor U29248 (N_29248,N_24634,N_22312);
xnor U29249 (N_29249,N_22572,N_24418);
and U29250 (N_29250,N_20884,N_23408);
and U29251 (N_29251,N_21209,N_21961);
xor U29252 (N_29252,N_20981,N_20328);
nor U29253 (N_29253,N_20009,N_22744);
or U29254 (N_29254,N_22810,N_23868);
xnor U29255 (N_29255,N_21353,N_21147);
or U29256 (N_29256,N_20147,N_23491);
nor U29257 (N_29257,N_23494,N_23070);
nor U29258 (N_29258,N_20933,N_20420);
and U29259 (N_29259,N_23662,N_23931);
or U29260 (N_29260,N_24774,N_24921);
or U29261 (N_29261,N_21754,N_24546);
nand U29262 (N_29262,N_21840,N_22402);
and U29263 (N_29263,N_24944,N_24437);
xor U29264 (N_29264,N_23691,N_21236);
nand U29265 (N_29265,N_20118,N_22952);
and U29266 (N_29266,N_24917,N_23753);
and U29267 (N_29267,N_20129,N_21942);
xor U29268 (N_29268,N_24437,N_20007);
nand U29269 (N_29269,N_22904,N_20861);
nor U29270 (N_29270,N_23000,N_20901);
and U29271 (N_29271,N_22213,N_22529);
nor U29272 (N_29272,N_22111,N_22321);
or U29273 (N_29273,N_23043,N_23211);
nor U29274 (N_29274,N_22165,N_21820);
xor U29275 (N_29275,N_24712,N_24419);
nor U29276 (N_29276,N_23484,N_22830);
or U29277 (N_29277,N_21186,N_23747);
xnor U29278 (N_29278,N_23810,N_22820);
xor U29279 (N_29279,N_22274,N_23024);
or U29280 (N_29280,N_20737,N_21863);
nand U29281 (N_29281,N_24038,N_24077);
and U29282 (N_29282,N_24591,N_23474);
and U29283 (N_29283,N_20627,N_24150);
xnor U29284 (N_29284,N_21267,N_22162);
nand U29285 (N_29285,N_24336,N_23833);
nor U29286 (N_29286,N_22990,N_22808);
xor U29287 (N_29287,N_22876,N_24695);
or U29288 (N_29288,N_21816,N_21189);
or U29289 (N_29289,N_20091,N_24014);
and U29290 (N_29290,N_22005,N_23210);
xor U29291 (N_29291,N_22035,N_24238);
xor U29292 (N_29292,N_23797,N_21582);
nand U29293 (N_29293,N_20095,N_22577);
or U29294 (N_29294,N_23805,N_20375);
or U29295 (N_29295,N_23013,N_20108);
nor U29296 (N_29296,N_20475,N_21580);
xnor U29297 (N_29297,N_20178,N_21897);
nor U29298 (N_29298,N_20526,N_22119);
nor U29299 (N_29299,N_20004,N_21019);
or U29300 (N_29300,N_24943,N_20117);
or U29301 (N_29301,N_22090,N_20920);
xnor U29302 (N_29302,N_21575,N_22109);
nand U29303 (N_29303,N_23446,N_23424);
nand U29304 (N_29304,N_21789,N_21615);
or U29305 (N_29305,N_24036,N_21036);
or U29306 (N_29306,N_20252,N_23542);
and U29307 (N_29307,N_20883,N_21372);
and U29308 (N_29308,N_24933,N_21434);
and U29309 (N_29309,N_21381,N_21327);
nor U29310 (N_29310,N_20307,N_24807);
nor U29311 (N_29311,N_20785,N_24046);
xor U29312 (N_29312,N_23074,N_23130);
xor U29313 (N_29313,N_21102,N_23576);
xnor U29314 (N_29314,N_24972,N_24153);
nor U29315 (N_29315,N_22441,N_21808);
nand U29316 (N_29316,N_22979,N_20755);
nand U29317 (N_29317,N_22311,N_20713);
or U29318 (N_29318,N_24174,N_24411);
or U29319 (N_29319,N_20648,N_24111);
or U29320 (N_29320,N_20166,N_24949);
and U29321 (N_29321,N_21634,N_21367);
and U29322 (N_29322,N_24951,N_24698);
or U29323 (N_29323,N_23015,N_21718);
nor U29324 (N_29324,N_23054,N_23502);
xnor U29325 (N_29325,N_21856,N_22689);
nand U29326 (N_29326,N_23695,N_20537);
and U29327 (N_29327,N_21755,N_24287);
nor U29328 (N_29328,N_20570,N_23020);
nand U29329 (N_29329,N_20054,N_20515);
and U29330 (N_29330,N_23262,N_22942);
and U29331 (N_29331,N_21687,N_21685);
or U29332 (N_29332,N_24597,N_23897);
or U29333 (N_29333,N_22459,N_24228);
and U29334 (N_29334,N_20131,N_22819);
nor U29335 (N_29335,N_24019,N_21859);
and U29336 (N_29336,N_23614,N_22888);
or U29337 (N_29337,N_21476,N_23240);
nand U29338 (N_29338,N_24276,N_24842);
or U29339 (N_29339,N_20063,N_22401);
xor U29340 (N_29340,N_22220,N_20701);
nor U29341 (N_29341,N_21458,N_21459);
nor U29342 (N_29342,N_24593,N_22315);
or U29343 (N_29343,N_23133,N_20027);
nand U29344 (N_29344,N_24520,N_24031);
or U29345 (N_29345,N_20936,N_23578);
and U29346 (N_29346,N_24020,N_22455);
nor U29347 (N_29347,N_23878,N_23916);
nor U29348 (N_29348,N_23236,N_23376);
or U29349 (N_29349,N_20203,N_20809);
or U29350 (N_29350,N_22054,N_20051);
or U29351 (N_29351,N_22970,N_20322);
xor U29352 (N_29352,N_23122,N_22922);
and U29353 (N_29353,N_24434,N_24134);
and U29354 (N_29354,N_23213,N_23414);
and U29355 (N_29355,N_24460,N_21949);
nor U29356 (N_29356,N_22221,N_20563);
nand U29357 (N_29357,N_22024,N_22430);
nand U29358 (N_29358,N_22888,N_21993);
xor U29359 (N_29359,N_24203,N_20420);
xnor U29360 (N_29360,N_22060,N_23838);
nand U29361 (N_29361,N_22325,N_21088);
nand U29362 (N_29362,N_23595,N_23550);
nand U29363 (N_29363,N_21284,N_24508);
nor U29364 (N_29364,N_22795,N_22500);
or U29365 (N_29365,N_23359,N_23374);
or U29366 (N_29366,N_23731,N_24297);
nand U29367 (N_29367,N_20596,N_24333);
nor U29368 (N_29368,N_24231,N_20844);
and U29369 (N_29369,N_22019,N_22553);
xnor U29370 (N_29370,N_24052,N_24965);
or U29371 (N_29371,N_22688,N_20337);
nor U29372 (N_29372,N_21984,N_20280);
nand U29373 (N_29373,N_20028,N_20225);
and U29374 (N_29374,N_20257,N_22162);
xor U29375 (N_29375,N_23714,N_24585);
and U29376 (N_29376,N_24136,N_22539);
or U29377 (N_29377,N_23366,N_21129);
and U29378 (N_29378,N_22805,N_22417);
xnor U29379 (N_29379,N_23246,N_24582);
nand U29380 (N_29380,N_23320,N_21318);
or U29381 (N_29381,N_20701,N_21531);
nor U29382 (N_29382,N_23885,N_20390);
or U29383 (N_29383,N_21212,N_23152);
or U29384 (N_29384,N_20566,N_24421);
nor U29385 (N_29385,N_20519,N_20780);
nand U29386 (N_29386,N_20909,N_21532);
xor U29387 (N_29387,N_24699,N_22409);
nand U29388 (N_29388,N_20002,N_23438);
and U29389 (N_29389,N_22290,N_20800);
nand U29390 (N_29390,N_21872,N_20143);
and U29391 (N_29391,N_22224,N_22574);
xnor U29392 (N_29392,N_24527,N_24315);
nor U29393 (N_29393,N_20630,N_21979);
or U29394 (N_29394,N_21089,N_20825);
nor U29395 (N_29395,N_20459,N_22888);
xnor U29396 (N_29396,N_21486,N_21056);
xor U29397 (N_29397,N_22661,N_20647);
nand U29398 (N_29398,N_24842,N_20574);
and U29399 (N_29399,N_20616,N_24282);
or U29400 (N_29400,N_23201,N_20222);
or U29401 (N_29401,N_23531,N_20789);
nand U29402 (N_29402,N_22080,N_20614);
and U29403 (N_29403,N_20239,N_22382);
nor U29404 (N_29404,N_20837,N_22759);
nand U29405 (N_29405,N_21229,N_21939);
xor U29406 (N_29406,N_24403,N_23378);
or U29407 (N_29407,N_21105,N_21656);
nand U29408 (N_29408,N_24121,N_21900);
nand U29409 (N_29409,N_24433,N_20720);
xor U29410 (N_29410,N_24169,N_22752);
xnor U29411 (N_29411,N_20869,N_23794);
nor U29412 (N_29412,N_23146,N_21112);
nand U29413 (N_29413,N_22460,N_21242);
nor U29414 (N_29414,N_22757,N_24873);
nor U29415 (N_29415,N_23213,N_20439);
nor U29416 (N_29416,N_20856,N_21174);
or U29417 (N_29417,N_21665,N_21623);
xnor U29418 (N_29418,N_24225,N_22768);
and U29419 (N_29419,N_22467,N_22984);
and U29420 (N_29420,N_24974,N_21771);
nand U29421 (N_29421,N_20861,N_20436);
nor U29422 (N_29422,N_23595,N_23018);
nand U29423 (N_29423,N_23599,N_24031);
xnor U29424 (N_29424,N_22950,N_24751);
nand U29425 (N_29425,N_21718,N_21044);
or U29426 (N_29426,N_24023,N_24488);
nand U29427 (N_29427,N_23368,N_21367);
nand U29428 (N_29428,N_24171,N_22835);
nand U29429 (N_29429,N_20998,N_21026);
or U29430 (N_29430,N_23648,N_22265);
nand U29431 (N_29431,N_20069,N_23226);
or U29432 (N_29432,N_24724,N_23366);
or U29433 (N_29433,N_22612,N_23694);
or U29434 (N_29434,N_24351,N_22371);
and U29435 (N_29435,N_24714,N_22724);
or U29436 (N_29436,N_21737,N_24623);
or U29437 (N_29437,N_24986,N_21313);
nor U29438 (N_29438,N_20316,N_20743);
nor U29439 (N_29439,N_22475,N_22278);
xor U29440 (N_29440,N_21884,N_22402);
xnor U29441 (N_29441,N_21369,N_20988);
nand U29442 (N_29442,N_23273,N_22374);
and U29443 (N_29443,N_20656,N_24354);
nor U29444 (N_29444,N_20610,N_21075);
nor U29445 (N_29445,N_22108,N_20223);
nor U29446 (N_29446,N_24275,N_21752);
nor U29447 (N_29447,N_23166,N_24256);
xnor U29448 (N_29448,N_20851,N_20371);
nor U29449 (N_29449,N_24706,N_21061);
nor U29450 (N_29450,N_24524,N_22402);
nor U29451 (N_29451,N_23457,N_23483);
nor U29452 (N_29452,N_23482,N_20129);
or U29453 (N_29453,N_22502,N_22781);
or U29454 (N_29454,N_24237,N_21227);
xnor U29455 (N_29455,N_20848,N_22080);
or U29456 (N_29456,N_24732,N_20030);
nand U29457 (N_29457,N_22689,N_22272);
xnor U29458 (N_29458,N_24656,N_23752);
nor U29459 (N_29459,N_23400,N_20740);
or U29460 (N_29460,N_20834,N_20766);
or U29461 (N_29461,N_21434,N_23805);
nand U29462 (N_29462,N_21719,N_20875);
xnor U29463 (N_29463,N_23223,N_20575);
and U29464 (N_29464,N_23672,N_24127);
nand U29465 (N_29465,N_23451,N_23824);
nor U29466 (N_29466,N_22167,N_23791);
and U29467 (N_29467,N_23272,N_22636);
xnor U29468 (N_29468,N_23253,N_20317);
and U29469 (N_29469,N_24170,N_24797);
nor U29470 (N_29470,N_22212,N_23510);
nor U29471 (N_29471,N_22153,N_23518);
or U29472 (N_29472,N_24810,N_20482);
nor U29473 (N_29473,N_23068,N_24141);
xor U29474 (N_29474,N_20076,N_23985);
nand U29475 (N_29475,N_21609,N_23696);
or U29476 (N_29476,N_24899,N_20246);
and U29477 (N_29477,N_24321,N_24278);
or U29478 (N_29478,N_22523,N_23469);
xnor U29479 (N_29479,N_22976,N_20479);
and U29480 (N_29480,N_20703,N_21601);
and U29481 (N_29481,N_20688,N_20617);
and U29482 (N_29482,N_21381,N_23359);
xnor U29483 (N_29483,N_20364,N_21582);
xnor U29484 (N_29484,N_21356,N_24116);
nand U29485 (N_29485,N_23425,N_24821);
xor U29486 (N_29486,N_20878,N_23837);
xnor U29487 (N_29487,N_23020,N_22599);
nand U29488 (N_29488,N_24677,N_23341);
nor U29489 (N_29489,N_20778,N_22870);
and U29490 (N_29490,N_22437,N_22746);
nor U29491 (N_29491,N_24002,N_22282);
nor U29492 (N_29492,N_24070,N_20603);
and U29493 (N_29493,N_21248,N_24220);
nand U29494 (N_29494,N_24352,N_22366);
nor U29495 (N_29495,N_20859,N_22074);
or U29496 (N_29496,N_22928,N_24784);
or U29497 (N_29497,N_22380,N_24987);
nor U29498 (N_29498,N_22945,N_24695);
or U29499 (N_29499,N_22693,N_20373);
nand U29500 (N_29500,N_21583,N_24005);
nand U29501 (N_29501,N_24021,N_21834);
nand U29502 (N_29502,N_22869,N_24839);
nor U29503 (N_29503,N_20295,N_21854);
or U29504 (N_29504,N_20489,N_22521);
or U29505 (N_29505,N_20556,N_22002);
nor U29506 (N_29506,N_22136,N_20783);
xnor U29507 (N_29507,N_21671,N_22048);
and U29508 (N_29508,N_23809,N_21215);
nor U29509 (N_29509,N_24083,N_21273);
xnor U29510 (N_29510,N_21282,N_24142);
and U29511 (N_29511,N_20722,N_23479);
and U29512 (N_29512,N_21428,N_24631);
nand U29513 (N_29513,N_24669,N_24254);
nand U29514 (N_29514,N_20786,N_20422);
and U29515 (N_29515,N_24395,N_24052);
xor U29516 (N_29516,N_20158,N_21658);
nand U29517 (N_29517,N_23585,N_22971);
and U29518 (N_29518,N_23755,N_20154);
xor U29519 (N_29519,N_20384,N_20486);
xnor U29520 (N_29520,N_22312,N_21122);
and U29521 (N_29521,N_21800,N_20992);
and U29522 (N_29522,N_24670,N_24842);
nand U29523 (N_29523,N_21987,N_23397);
xnor U29524 (N_29524,N_24174,N_20261);
xnor U29525 (N_29525,N_20905,N_22033);
nand U29526 (N_29526,N_22159,N_20353);
xor U29527 (N_29527,N_23714,N_24817);
or U29528 (N_29528,N_24264,N_23061);
nand U29529 (N_29529,N_20632,N_20436);
xor U29530 (N_29530,N_24391,N_21683);
or U29531 (N_29531,N_24828,N_24646);
nand U29532 (N_29532,N_21973,N_23319);
nor U29533 (N_29533,N_23128,N_23359);
and U29534 (N_29534,N_24338,N_21237);
nor U29535 (N_29535,N_21297,N_24561);
nand U29536 (N_29536,N_23424,N_21946);
nor U29537 (N_29537,N_23347,N_24489);
and U29538 (N_29538,N_21589,N_23424);
nand U29539 (N_29539,N_22034,N_24033);
or U29540 (N_29540,N_24452,N_23076);
nand U29541 (N_29541,N_22670,N_23287);
nor U29542 (N_29542,N_21201,N_21013);
nand U29543 (N_29543,N_22393,N_21844);
nor U29544 (N_29544,N_20289,N_23941);
and U29545 (N_29545,N_21605,N_24464);
nor U29546 (N_29546,N_21270,N_22397);
nand U29547 (N_29547,N_21798,N_22665);
and U29548 (N_29548,N_23241,N_22435);
or U29549 (N_29549,N_24161,N_23978);
or U29550 (N_29550,N_24851,N_22034);
nor U29551 (N_29551,N_23952,N_20451);
nor U29552 (N_29552,N_23977,N_21498);
xor U29553 (N_29553,N_24922,N_22698);
xor U29554 (N_29554,N_23496,N_22179);
and U29555 (N_29555,N_21549,N_22911);
nor U29556 (N_29556,N_21343,N_21162);
and U29557 (N_29557,N_24370,N_20615);
nand U29558 (N_29558,N_21245,N_24638);
nor U29559 (N_29559,N_21499,N_23767);
nand U29560 (N_29560,N_21046,N_22540);
nor U29561 (N_29561,N_23557,N_20498);
or U29562 (N_29562,N_24208,N_20332);
nand U29563 (N_29563,N_23375,N_20766);
and U29564 (N_29564,N_20124,N_20175);
or U29565 (N_29565,N_22528,N_21277);
nand U29566 (N_29566,N_22971,N_20758);
and U29567 (N_29567,N_20688,N_22696);
xnor U29568 (N_29568,N_24878,N_22384);
or U29569 (N_29569,N_20387,N_23719);
nand U29570 (N_29570,N_20078,N_23052);
nor U29571 (N_29571,N_22633,N_21653);
xor U29572 (N_29572,N_20297,N_20645);
or U29573 (N_29573,N_20561,N_24212);
xnor U29574 (N_29574,N_20617,N_20341);
and U29575 (N_29575,N_20836,N_20371);
nor U29576 (N_29576,N_22840,N_22244);
xnor U29577 (N_29577,N_20635,N_21958);
nand U29578 (N_29578,N_23636,N_20707);
nand U29579 (N_29579,N_21901,N_22519);
nand U29580 (N_29580,N_20648,N_22336);
and U29581 (N_29581,N_23570,N_23495);
nor U29582 (N_29582,N_21752,N_20928);
nand U29583 (N_29583,N_23664,N_22310);
nand U29584 (N_29584,N_21551,N_24872);
or U29585 (N_29585,N_24222,N_23551);
nor U29586 (N_29586,N_20337,N_20864);
or U29587 (N_29587,N_23539,N_22264);
or U29588 (N_29588,N_22552,N_22444);
nand U29589 (N_29589,N_21053,N_23547);
and U29590 (N_29590,N_20410,N_23394);
or U29591 (N_29591,N_24043,N_22722);
and U29592 (N_29592,N_24570,N_23648);
nand U29593 (N_29593,N_23962,N_21175);
or U29594 (N_29594,N_21110,N_24933);
xor U29595 (N_29595,N_22824,N_23461);
and U29596 (N_29596,N_23890,N_20915);
nand U29597 (N_29597,N_22772,N_23181);
and U29598 (N_29598,N_20687,N_21359);
and U29599 (N_29599,N_21559,N_23993);
and U29600 (N_29600,N_24204,N_24285);
and U29601 (N_29601,N_24866,N_22086);
and U29602 (N_29602,N_21551,N_23200);
nand U29603 (N_29603,N_21521,N_22562);
xor U29604 (N_29604,N_21057,N_22446);
nand U29605 (N_29605,N_20559,N_24114);
xor U29606 (N_29606,N_22914,N_21060);
xnor U29607 (N_29607,N_24298,N_23533);
xor U29608 (N_29608,N_23264,N_21028);
nor U29609 (N_29609,N_23728,N_22102);
xnor U29610 (N_29610,N_23816,N_22408);
nor U29611 (N_29611,N_23386,N_20613);
and U29612 (N_29612,N_24281,N_21112);
nand U29613 (N_29613,N_22351,N_24610);
or U29614 (N_29614,N_22651,N_21484);
and U29615 (N_29615,N_20727,N_20364);
nand U29616 (N_29616,N_22224,N_22562);
xor U29617 (N_29617,N_24506,N_24635);
or U29618 (N_29618,N_21921,N_20436);
and U29619 (N_29619,N_20347,N_23068);
xor U29620 (N_29620,N_22374,N_24073);
and U29621 (N_29621,N_22802,N_23689);
and U29622 (N_29622,N_24833,N_22455);
nor U29623 (N_29623,N_21860,N_24727);
and U29624 (N_29624,N_20378,N_24593);
or U29625 (N_29625,N_21332,N_21653);
nor U29626 (N_29626,N_21243,N_23669);
xor U29627 (N_29627,N_21500,N_20203);
and U29628 (N_29628,N_23730,N_22902);
nand U29629 (N_29629,N_24940,N_23392);
nand U29630 (N_29630,N_20426,N_22375);
and U29631 (N_29631,N_21996,N_21544);
nor U29632 (N_29632,N_20060,N_22698);
nor U29633 (N_29633,N_22636,N_24031);
xor U29634 (N_29634,N_20874,N_24955);
nand U29635 (N_29635,N_24278,N_20200);
and U29636 (N_29636,N_21431,N_22753);
nor U29637 (N_29637,N_20943,N_24643);
and U29638 (N_29638,N_22415,N_20868);
and U29639 (N_29639,N_24175,N_23614);
nand U29640 (N_29640,N_21252,N_23035);
nor U29641 (N_29641,N_20590,N_22245);
nor U29642 (N_29642,N_20699,N_23877);
and U29643 (N_29643,N_23470,N_20110);
nor U29644 (N_29644,N_20412,N_24079);
or U29645 (N_29645,N_22112,N_23535);
nor U29646 (N_29646,N_21924,N_21557);
nand U29647 (N_29647,N_24040,N_21934);
nand U29648 (N_29648,N_20182,N_22186);
or U29649 (N_29649,N_23307,N_23688);
nand U29650 (N_29650,N_20665,N_24282);
or U29651 (N_29651,N_24772,N_20471);
nand U29652 (N_29652,N_20593,N_24499);
xor U29653 (N_29653,N_23863,N_22212);
and U29654 (N_29654,N_22191,N_21349);
and U29655 (N_29655,N_23934,N_23298);
or U29656 (N_29656,N_23129,N_22059);
and U29657 (N_29657,N_22976,N_21260);
nor U29658 (N_29658,N_21890,N_23515);
and U29659 (N_29659,N_21877,N_23183);
or U29660 (N_29660,N_20135,N_21346);
or U29661 (N_29661,N_24513,N_21174);
nor U29662 (N_29662,N_20769,N_24006);
and U29663 (N_29663,N_22702,N_22056);
and U29664 (N_29664,N_23136,N_20695);
or U29665 (N_29665,N_20632,N_24054);
xor U29666 (N_29666,N_23970,N_23009);
or U29667 (N_29667,N_23100,N_24620);
nand U29668 (N_29668,N_20225,N_23226);
nor U29669 (N_29669,N_24144,N_20812);
nand U29670 (N_29670,N_20212,N_20472);
and U29671 (N_29671,N_21486,N_21900);
or U29672 (N_29672,N_21094,N_20638);
nor U29673 (N_29673,N_21499,N_22542);
and U29674 (N_29674,N_23683,N_23927);
nor U29675 (N_29675,N_21006,N_24418);
or U29676 (N_29676,N_22709,N_22308);
xnor U29677 (N_29677,N_22253,N_24852);
nor U29678 (N_29678,N_20619,N_21710);
or U29679 (N_29679,N_22428,N_23128);
nand U29680 (N_29680,N_20665,N_20584);
and U29681 (N_29681,N_20449,N_22137);
nand U29682 (N_29682,N_20370,N_24388);
nor U29683 (N_29683,N_20306,N_24650);
or U29684 (N_29684,N_22793,N_22008);
and U29685 (N_29685,N_23036,N_22915);
and U29686 (N_29686,N_22392,N_22634);
nor U29687 (N_29687,N_23229,N_23624);
and U29688 (N_29688,N_23076,N_22483);
nand U29689 (N_29689,N_20918,N_21829);
nor U29690 (N_29690,N_23754,N_23935);
nor U29691 (N_29691,N_24545,N_24557);
and U29692 (N_29692,N_20720,N_23540);
nor U29693 (N_29693,N_22243,N_24466);
and U29694 (N_29694,N_24901,N_23972);
and U29695 (N_29695,N_21244,N_20487);
nor U29696 (N_29696,N_23061,N_21075);
and U29697 (N_29697,N_21338,N_23643);
and U29698 (N_29698,N_23486,N_23755);
nor U29699 (N_29699,N_21668,N_22738);
and U29700 (N_29700,N_21787,N_21769);
xor U29701 (N_29701,N_22717,N_20555);
nand U29702 (N_29702,N_20191,N_24794);
nor U29703 (N_29703,N_22598,N_20828);
and U29704 (N_29704,N_23203,N_24765);
and U29705 (N_29705,N_22310,N_20429);
or U29706 (N_29706,N_22874,N_21571);
or U29707 (N_29707,N_24907,N_23206);
xor U29708 (N_29708,N_20763,N_20198);
and U29709 (N_29709,N_24692,N_20760);
and U29710 (N_29710,N_23304,N_21154);
nor U29711 (N_29711,N_24997,N_24061);
nand U29712 (N_29712,N_24329,N_22003);
or U29713 (N_29713,N_22870,N_21596);
and U29714 (N_29714,N_21376,N_22260);
nand U29715 (N_29715,N_21870,N_21701);
and U29716 (N_29716,N_21097,N_23821);
nand U29717 (N_29717,N_20097,N_21138);
nand U29718 (N_29718,N_20789,N_24220);
nand U29719 (N_29719,N_21299,N_22056);
nor U29720 (N_29720,N_23719,N_22732);
nand U29721 (N_29721,N_20365,N_24188);
and U29722 (N_29722,N_24584,N_21983);
xor U29723 (N_29723,N_20246,N_23293);
nand U29724 (N_29724,N_22058,N_23310);
or U29725 (N_29725,N_20274,N_20059);
xor U29726 (N_29726,N_20839,N_20732);
or U29727 (N_29727,N_20305,N_20408);
nor U29728 (N_29728,N_20688,N_20082);
nand U29729 (N_29729,N_24566,N_24400);
xnor U29730 (N_29730,N_23338,N_22353);
and U29731 (N_29731,N_22917,N_20245);
nor U29732 (N_29732,N_22289,N_21578);
nor U29733 (N_29733,N_22140,N_24011);
or U29734 (N_29734,N_23792,N_22527);
xnor U29735 (N_29735,N_20938,N_22673);
nand U29736 (N_29736,N_22386,N_23259);
and U29737 (N_29737,N_21942,N_24987);
xor U29738 (N_29738,N_22209,N_20327);
nor U29739 (N_29739,N_23988,N_23573);
and U29740 (N_29740,N_22407,N_24709);
and U29741 (N_29741,N_20331,N_21924);
or U29742 (N_29742,N_21887,N_21984);
or U29743 (N_29743,N_24294,N_20051);
and U29744 (N_29744,N_24715,N_21047);
nor U29745 (N_29745,N_24398,N_21558);
xnor U29746 (N_29746,N_22490,N_21249);
and U29747 (N_29747,N_20629,N_24861);
and U29748 (N_29748,N_24680,N_23557);
xnor U29749 (N_29749,N_21715,N_22645);
nor U29750 (N_29750,N_20008,N_23345);
nor U29751 (N_29751,N_20112,N_23992);
and U29752 (N_29752,N_20579,N_23671);
or U29753 (N_29753,N_20961,N_23842);
xnor U29754 (N_29754,N_22835,N_20070);
or U29755 (N_29755,N_24457,N_20661);
xor U29756 (N_29756,N_24005,N_23968);
nand U29757 (N_29757,N_21902,N_20775);
and U29758 (N_29758,N_24345,N_22792);
or U29759 (N_29759,N_21086,N_22134);
nor U29760 (N_29760,N_22500,N_22991);
nor U29761 (N_29761,N_22795,N_24486);
and U29762 (N_29762,N_22427,N_20573);
nand U29763 (N_29763,N_21315,N_23046);
nand U29764 (N_29764,N_22058,N_23897);
or U29765 (N_29765,N_22112,N_22117);
or U29766 (N_29766,N_21291,N_22287);
nor U29767 (N_29767,N_23935,N_24612);
nor U29768 (N_29768,N_21203,N_24256);
xnor U29769 (N_29769,N_22775,N_21906);
nor U29770 (N_29770,N_21200,N_21483);
nor U29771 (N_29771,N_21472,N_24021);
xor U29772 (N_29772,N_24119,N_24477);
nand U29773 (N_29773,N_24866,N_21404);
nor U29774 (N_29774,N_22342,N_21788);
xnor U29775 (N_29775,N_22896,N_24095);
nor U29776 (N_29776,N_24625,N_22840);
xor U29777 (N_29777,N_21364,N_24695);
xnor U29778 (N_29778,N_20848,N_22130);
nor U29779 (N_29779,N_20169,N_22406);
xor U29780 (N_29780,N_20711,N_23107);
and U29781 (N_29781,N_22883,N_24693);
and U29782 (N_29782,N_20270,N_22184);
and U29783 (N_29783,N_23704,N_20911);
nor U29784 (N_29784,N_20204,N_22327);
nand U29785 (N_29785,N_20841,N_20761);
xor U29786 (N_29786,N_21351,N_24775);
nand U29787 (N_29787,N_20284,N_24948);
xor U29788 (N_29788,N_24374,N_21549);
nor U29789 (N_29789,N_24995,N_22912);
or U29790 (N_29790,N_20947,N_20218);
nor U29791 (N_29791,N_22835,N_22702);
and U29792 (N_29792,N_22810,N_24191);
and U29793 (N_29793,N_22601,N_22726);
and U29794 (N_29794,N_23978,N_22074);
nand U29795 (N_29795,N_20581,N_21901);
or U29796 (N_29796,N_20551,N_23622);
or U29797 (N_29797,N_21497,N_24996);
nand U29798 (N_29798,N_21851,N_24712);
or U29799 (N_29799,N_24721,N_22341);
nor U29800 (N_29800,N_24668,N_20052);
nand U29801 (N_29801,N_21808,N_20140);
nor U29802 (N_29802,N_21483,N_22710);
or U29803 (N_29803,N_22784,N_22071);
xor U29804 (N_29804,N_24046,N_23617);
and U29805 (N_29805,N_24564,N_20603);
or U29806 (N_29806,N_24530,N_22111);
nand U29807 (N_29807,N_20745,N_23314);
xnor U29808 (N_29808,N_23742,N_24273);
nand U29809 (N_29809,N_21147,N_20549);
xnor U29810 (N_29810,N_22037,N_21628);
xor U29811 (N_29811,N_23294,N_21384);
nor U29812 (N_29812,N_22224,N_23587);
and U29813 (N_29813,N_20519,N_20709);
nand U29814 (N_29814,N_21511,N_24638);
and U29815 (N_29815,N_20077,N_21037);
or U29816 (N_29816,N_20461,N_23925);
or U29817 (N_29817,N_20440,N_22405);
nor U29818 (N_29818,N_24000,N_21544);
and U29819 (N_29819,N_22811,N_20958);
nor U29820 (N_29820,N_22708,N_23743);
nand U29821 (N_29821,N_24548,N_23508);
or U29822 (N_29822,N_22698,N_20441);
nor U29823 (N_29823,N_21090,N_22486);
or U29824 (N_29824,N_22616,N_24619);
and U29825 (N_29825,N_20430,N_21412);
nand U29826 (N_29826,N_21536,N_21159);
and U29827 (N_29827,N_22260,N_22715);
nor U29828 (N_29828,N_24310,N_23619);
nand U29829 (N_29829,N_22789,N_23209);
and U29830 (N_29830,N_24601,N_20483);
and U29831 (N_29831,N_24708,N_24052);
or U29832 (N_29832,N_21799,N_22588);
nand U29833 (N_29833,N_22072,N_21635);
nor U29834 (N_29834,N_22391,N_21043);
xor U29835 (N_29835,N_23182,N_24201);
and U29836 (N_29836,N_23213,N_23043);
nor U29837 (N_29837,N_24409,N_24726);
nand U29838 (N_29838,N_23911,N_20591);
nand U29839 (N_29839,N_22155,N_24046);
nor U29840 (N_29840,N_24584,N_24116);
and U29841 (N_29841,N_23133,N_22315);
nand U29842 (N_29842,N_20884,N_22747);
xnor U29843 (N_29843,N_23226,N_20594);
xnor U29844 (N_29844,N_24440,N_20264);
nand U29845 (N_29845,N_23450,N_23478);
nor U29846 (N_29846,N_22740,N_21662);
nand U29847 (N_29847,N_22414,N_20958);
nand U29848 (N_29848,N_21991,N_24716);
and U29849 (N_29849,N_22116,N_22946);
xor U29850 (N_29850,N_23950,N_20079);
nand U29851 (N_29851,N_22382,N_22354);
and U29852 (N_29852,N_22588,N_22033);
or U29853 (N_29853,N_22248,N_23717);
xor U29854 (N_29854,N_24148,N_24146);
and U29855 (N_29855,N_22414,N_24050);
or U29856 (N_29856,N_22064,N_22200);
nand U29857 (N_29857,N_24706,N_24442);
nand U29858 (N_29858,N_24867,N_21778);
nor U29859 (N_29859,N_22481,N_21482);
nand U29860 (N_29860,N_23682,N_21878);
or U29861 (N_29861,N_23316,N_20631);
or U29862 (N_29862,N_23654,N_20626);
nand U29863 (N_29863,N_20377,N_23233);
xor U29864 (N_29864,N_24417,N_22644);
or U29865 (N_29865,N_23903,N_20110);
and U29866 (N_29866,N_22262,N_24632);
or U29867 (N_29867,N_22035,N_20031);
xor U29868 (N_29868,N_20745,N_21019);
or U29869 (N_29869,N_22732,N_24802);
or U29870 (N_29870,N_22247,N_21378);
nor U29871 (N_29871,N_23136,N_23554);
nand U29872 (N_29872,N_24850,N_23239);
and U29873 (N_29873,N_24460,N_20693);
or U29874 (N_29874,N_23408,N_20228);
nor U29875 (N_29875,N_22801,N_24815);
or U29876 (N_29876,N_22509,N_21667);
nand U29877 (N_29877,N_20354,N_24689);
xor U29878 (N_29878,N_24254,N_21590);
nor U29879 (N_29879,N_21693,N_22608);
and U29880 (N_29880,N_22577,N_22134);
and U29881 (N_29881,N_24121,N_24137);
nor U29882 (N_29882,N_21495,N_24269);
nand U29883 (N_29883,N_22049,N_20568);
nor U29884 (N_29884,N_24661,N_20823);
nand U29885 (N_29885,N_22388,N_21730);
and U29886 (N_29886,N_21271,N_24724);
xor U29887 (N_29887,N_20864,N_24164);
nor U29888 (N_29888,N_24265,N_20058);
or U29889 (N_29889,N_21112,N_23882);
xnor U29890 (N_29890,N_23334,N_23984);
nand U29891 (N_29891,N_21515,N_22849);
xnor U29892 (N_29892,N_23916,N_23662);
or U29893 (N_29893,N_22570,N_23361);
xor U29894 (N_29894,N_22647,N_23033);
nand U29895 (N_29895,N_22592,N_22054);
xnor U29896 (N_29896,N_20736,N_22136);
or U29897 (N_29897,N_21600,N_24574);
or U29898 (N_29898,N_24285,N_22097);
xor U29899 (N_29899,N_22399,N_22838);
or U29900 (N_29900,N_20200,N_22027);
nor U29901 (N_29901,N_23459,N_21631);
nor U29902 (N_29902,N_23680,N_22447);
and U29903 (N_29903,N_20553,N_22183);
and U29904 (N_29904,N_23625,N_21854);
nand U29905 (N_29905,N_22733,N_20175);
nand U29906 (N_29906,N_23726,N_20884);
xor U29907 (N_29907,N_22250,N_21252);
nand U29908 (N_29908,N_20178,N_20875);
xnor U29909 (N_29909,N_21570,N_23657);
nand U29910 (N_29910,N_22104,N_20416);
or U29911 (N_29911,N_20621,N_23245);
xnor U29912 (N_29912,N_23235,N_21812);
nor U29913 (N_29913,N_22722,N_22810);
and U29914 (N_29914,N_22142,N_20834);
nand U29915 (N_29915,N_24332,N_23567);
xor U29916 (N_29916,N_22241,N_22160);
or U29917 (N_29917,N_22511,N_21678);
nor U29918 (N_29918,N_22839,N_20839);
nand U29919 (N_29919,N_20432,N_22079);
or U29920 (N_29920,N_24788,N_23355);
and U29921 (N_29921,N_22853,N_22687);
and U29922 (N_29922,N_23901,N_23831);
nand U29923 (N_29923,N_24000,N_21011);
xnor U29924 (N_29924,N_23258,N_22932);
nand U29925 (N_29925,N_22585,N_20672);
nor U29926 (N_29926,N_23515,N_20191);
nand U29927 (N_29927,N_24731,N_23282);
nor U29928 (N_29928,N_20656,N_22718);
xor U29929 (N_29929,N_21253,N_21539);
nand U29930 (N_29930,N_23250,N_22846);
or U29931 (N_29931,N_20712,N_23092);
xnor U29932 (N_29932,N_22800,N_22721);
nor U29933 (N_29933,N_24271,N_23084);
nand U29934 (N_29934,N_20158,N_23707);
or U29935 (N_29935,N_24732,N_23742);
and U29936 (N_29936,N_23427,N_21986);
or U29937 (N_29937,N_20440,N_20787);
and U29938 (N_29938,N_22314,N_20807);
and U29939 (N_29939,N_20101,N_20718);
xor U29940 (N_29940,N_24264,N_23889);
and U29941 (N_29941,N_23400,N_20618);
or U29942 (N_29942,N_24132,N_24555);
and U29943 (N_29943,N_21818,N_22127);
and U29944 (N_29944,N_21399,N_20245);
and U29945 (N_29945,N_23153,N_20633);
nor U29946 (N_29946,N_24791,N_23230);
or U29947 (N_29947,N_24115,N_21176);
or U29948 (N_29948,N_21067,N_23854);
or U29949 (N_29949,N_22819,N_21553);
nand U29950 (N_29950,N_21194,N_22857);
nor U29951 (N_29951,N_22976,N_24443);
xnor U29952 (N_29952,N_21111,N_23212);
and U29953 (N_29953,N_23683,N_20983);
or U29954 (N_29954,N_24911,N_20694);
and U29955 (N_29955,N_20270,N_23721);
xnor U29956 (N_29956,N_22435,N_24940);
nand U29957 (N_29957,N_23507,N_20493);
nand U29958 (N_29958,N_20932,N_23600);
nand U29959 (N_29959,N_20366,N_22812);
nor U29960 (N_29960,N_20869,N_21076);
and U29961 (N_29961,N_20684,N_23538);
nor U29962 (N_29962,N_22942,N_24633);
nand U29963 (N_29963,N_21772,N_23105);
or U29964 (N_29964,N_22752,N_23877);
nand U29965 (N_29965,N_23659,N_20921);
nand U29966 (N_29966,N_24955,N_23417);
or U29967 (N_29967,N_22253,N_23044);
and U29968 (N_29968,N_22326,N_22932);
nand U29969 (N_29969,N_21464,N_20198);
nor U29970 (N_29970,N_21569,N_22098);
or U29971 (N_29971,N_21063,N_23220);
or U29972 (N_29972,N_22466,N_24588);
or U29973 (N_29973,N_21400,N_21933);
and U29974 (N_29974,N_22072,N_22206);
xor U29975 (N_29975,N_21838,N_23764);
xnor U29976 (N_29976,N_24753,N_24473);
nand U29977 (N_29977,N_24013,N_20360);
or U29978 (N_29978,N_21865,N_23384);
nand U29979 (N_29979,N_23300,N_24260);
xor U29980 (N_29980,N_23799,N_20750);
or U29981 (N_29981,N_21872,N_24380);
and U29982 (N_29982,N_24282,N_23199);
xnor U29983 (N_29983,N_21127,N_22745);
and U29984 (N_29984,N_21979,N_21799);
or U29985 (N_29985,N_22936,N_20249);
xnor U29986 (N_29986,N_24663,N_24994);
xnor U29987 (N_29987,N_21428,N_23069);
xnor U29988 (N_29988,N_24530,N_20162);
nor U29989 (N_29989,N_20976,N_23834);
xnor U29990 (N_29990,N_20939,N_20545);
and U29991 (N_29991,N_20725,N_24411);
xnor U29992 (N_29992,N_21602,N_22398);
nand U29993 (N_29993,N_21578,N_23051);
nor U29994 (N_29994,N_21830,N_20927);
or U29995 (N_29995,N_24020,N_22566);
nor U29996 (N_29996,N_24806,N_22956);
or U29997 (N_29997,N_24040,N_22021);
nand U29998 (N_29998,N_24238,N_23125);
nand U29999 (N_29999,N_23498,N_23284);
nand UO_0 (O_0,N_27124,N_29184);
nand UO_1 (O_1,N_29976,N_26754);
nor UO_2 (O_2,N_25284,N_27985);
nor UO_3 (O_3,N_29781,N_25704);
and UO_4 (O_4,N_29622,N_28675);
nor UO_5 (O_5,N_26596,N_25805);
nand UO_6 (O_6,N_26755,N_26594);
xor UO_7 (O_7,N_28927,N_25330);
nor UO_8 (O_8,N_26468,N_27462);
nand UO_9 (O_9,N_28357,N_27548);
and UO_10 (O_10,N_29129,N_27580);
nor UO_11 (O_11,N_29078,N_26285);
xor UO_12 (O_12,N_27507,N_26688);
and UO_13 (O_13,N_26588,N_27719);
and UO_14 (O_14,N_26020,N_28176);
nor UO_15 (O_15,N_28003,N_29346);
or UO_16 (O_16,N_28402,N_26905);
nand UO_17 (O_17,N_29283,N_27598);
or UO_18 (O_18,N_29165,N_25645);
and UO_19 (O_19,N_26088,N_26400);
xnor UO_20 (O_20,N_28628,N_26912);
xor UO_21 (O_21,N_26550,N_28784);
nand UO_22 (O_22,N_27140,N_25475);
xnor UO_23 (O_23,N_28332,N_25355);
nor UO_24 (O_24,N_25473,N_29607);
xnor UO_25 (O_25,N_25509,N_27976);
nand UO_26 (O_26,N_26960,N_26707);
nand UO_27 (O_27,N_27804,N_29577);
nor UO_28 (O_28,N_26178,N_27585);
nand UO_29 (O_29,N_25906,N_25630);
nand UO_30 (O_30,N_28672,N_27289);
or UO_31 (O_31,N_27223,N_25610);
nand UO_32 (O_32,N_28345,N_28616);
nand UO_33 (O_33,N_29090,N_29025);
nor UO_34 (O_34,N_28701,N_27991);
xnor UO_35 (O_35,N_27736,N_25295);
or UO_36 (O_36,N_29169,N_25121);
nand UO_37 (O_37,N_27351,N_27744);
or UO_38 (O_38,N_29814,N_27635);
and UO_39 (O_39,N_29952,N_28949);
or UO_40 (O_40,N_29718,N_25700);
and UO_41 (O_41,N_25480,N_26577);
nand UO_42 (O_42,N_28319,N_27849);
xor UO_43 (O_43,N_29995,N_26925);
and UO_44 (O_44,N_29344,N_27317);
nand UO_45 (O_45,N_28638,N_27735);
nand UO_46 (O_46,N_26263,N_27931);
and UO_47 (O_47,N_26555,N_25343);
nand UO_48 (O_48,N_29270,N_25593);
or UO_49 (O_49,N_28414,N_28940);
nor UO_50 (O_50,N_27691,N_27499);
or UO_51 (O_51,N_28432,N_28517);
xor UO_52 (O_52,N_25799,N_27158);
nand UO_53 (O_53,N_28886,N_25926);
nand UO_54 (O_54,N_27162,N_26337);
nor UO_55 (O_55,N_27536,N_29942);
and UO_56 (O_56,N_29110,N_25611);
or UO_57 (O_57,N_28437,N_25241);
nor UO_58 (O_58,N_26028,N_28774);
and UO_59 (O_59,N_27305,N_29771);
xnor UO_60 (O_60,N_25770,N_29725);
or UO_61 (O_61,N_28843,N_25697);
nor UO_62 (O_62,N_27771,N_28876);
and UO_63 (O_63,N_27617,N_29943);
xor UO_64 (O_64,N_29980,N_27712);
xor UO_65 (O_65,N_26006,N_26981);
nand UO_66 (O_66,N_28561,N_28852);
or UO_67 (O_67,N_27412,N_25349);
or UO_68 (O_68,N_29039,N_25763);
xor UO_69 (O_69,N_26237,N_26019);
or UO_70 (O_70,N_26112,N_29961);
nor UO_71 (O_71,N_29068,N_25572);
nand UO_72 (O_72,N_25790,N_26748);
xor UO_73 (O_73,N_27438,N_27559);
nand UO_74 (O_74,N_29438,N_27323);
or UO_75 (O_75,N_25250,N_26252);
nand UO_76 (O_76,N_26916,N_29533);
and UO_77 (O_77,N_29256,N_25338);
nand UO_78 (O_78,N_29323,N_28819);
or UO_79 (O_79,N_28216,N_25052);
nand UO_80 (O_80,N_29712,N_27599);
nor UO_81 (O_81,N_25915,N_28869);
and UO_82 (O_82,N_27873,N_28566);
and UO_83 (O_83,N_27402,N_26266);
nand UO_84 (O_84,N_25108,N_26012);
xor UO_85 (O_85,N_29233,N_26447);
nor UO_86 (O_86,N_29757,N_29565);
nand UO_87 (O_87,N_27489,N_29773);
nor UO_88 (O_88,N_28148,N_29208);
nor UO_89 (O_89,N_26639,N_28063);
nor UO_90 (O_90,N_29195,N_28746);
xor UO_91 (O_91,N_27163,N_27994);
or UO_92 (O_92,N_29595,N_29625);
xnor UO_93 (O_93,N_29618,N_27298);
nor UO_94 (O_94,N_29998,N_27503);
nand UO_95 (O_95,N_25526,N_28583);
nand UO_96 (O_96,N_28861,N_29353);
xnor UO_97 (O_97,N_29471,N_29485);
or UO_98 (O_98,N_29237,N_26246);
xnor UO_99 (O_99,N_26305,N_28854);
xor UO_100 (O_100,N_29633,N_29464);
or UO_101 (O_101,N_27566,N_28917);
xor UO_102 (O_102,N_29951,N_28247);
nor UO_103 (O_103,N_26693,N_29540);
or UO_104 (O_104,N_26378,N_26842);
xor UO_105 (O_105,N_26568,N_25647);
nor UO_106 (O_106,N_27509,N_28849);
nor UO_107 (O_107,N_27715,N_25626);
nor UO_108 (O_108,N_27043,N_26223);
nor UO_109 (O_109,N_25754,N_29430);
xor UO_110 (O_110,N_26073,N_26728);
or UO_111 (O_111,N_27666,N_25225);
and UO_112 (O_112,N_28356,N_29907);
and UO_113 (O_113,N_29305,N_26827);
nand UO_114 (O_114,N_29893,N_29067);
or UO_115 (O_115,N_25598,N_26749);
or UO_116 (O_116,N_28095,N_25129);
xor UO_117 (O_117,N_25416,N_29212);
nor UO_118 (O_118,N_29659,N_25567);
xnor UO_119 (O_119,N_29704,N_27961);
xnor UO_120 (O_120,N_27600,N_26092);
or UO_121 (O_121,N_25551,N_26167);
xnor UO_122 (O_122,N_29535,N_29710);
xor UO_123 (O_123,N_26957,N_26431);
nor UO_124 (O_124,N_25076,N_26722);
and UO_125 (O_125,N_25286,N_25372);
or UO_126 (O_126,N_29468,N_29593);
and UO_127 (O_127,N_27819,N_25163);
nor UO_128 (O_128,N_25390,N_25171);
and UO_129 (O_129,N_27777,N_29437);
xor UO_130 (O_130,N_28966,N_25822);
xnor UO_131 (O_131,N_26674,N_27947);
or UO_132 (O_132,N_27946,N_28707);
and UO_133 (O_133,N_29677,N_25318);
or UO_134 (O_134,N_26949,N_25079);
or UO_135 (O_135,N_29063,N_26430);
nand UO_136 (O_136,N_28469,N_25890);
or UO_137 (O_137,N_29466,N_28403);
xor UO_138 (O_138,N_25333,N_28604);
nor UO_139 (O_139,N_27921,N_28633);
or UO_140 (O_140,N_28637,N_26318);
and UO_141 (O_141,N_26018,N_25094);
or UO_142 (O_142,N_27386,N_27549);
xor UO_143 (O_143,N_28549,N_26881);
nor UO_144 (O_144,N_28687,N_25077);
and UO_145 (O_145,N_27123,N_27663);
or UO_146 (O_146,N_28931,N_25635);
or UO_147 (O_147,N_28121,N_26498);
nand UO_148 (O_148,N_29138,N_27579);
nand UO_149 (O_149,N_27710,N_26801);
xnor UO_150 (O_150,N_28735,N_28495);
xor UO_151 (O_151,N_27825,N_26240);
nand UO_152 (O_152,N_27845,N_27775);
nor UO_153 (O_153,N_25054,N_26220);
and UO_154 (O_154,N_25975,N_26419);
xor UO_155 (O_155,N_28499,N_28941);
xor UO_156 (O_156,N_26816,N_26775);
xor UO_157 (O_157,N_27066,N_26614);
nand UO_158 (O_158,N_27679,N_29339);
nor UO_159 (O_159,N_25796,N_26093);
nor UO_160 (O_160,N_26806,N_27618);
xor UO_161 (O_161,N_25582,N_28807);
nor UO_162 (O_162,N_28490,N_27091);
or UO_163 (O_163,N_26288,N_26508);
nor UO_164 (O_164,N_25298,N_27912);
nand UO_165 (O_165,N_28202,N_25989);
and UO_166 (O_166,N_25281,N_28799);
nor UO_167 (O_167,N_25184,N_27854);
nor UO_168 (O_168,N_25707,N_27619);
nand UO_169 (O_169,N_25973,N_28359);
nand UO_170 (O_170,N_27109,N_28004);
and UO_171 (O_171,N_29366,N_28000);
xor UO_172 (O_172,N_25090,N_29307);
or UO_173 (O_173,N_28040,N_28393);
and UO_174 (O_174,N_26225,N_28162);
xor UO_175 (O_175,N_25191,N_25395);
or UO_176 (O_176,N_27723,N_29018);
nand UO_177 (O_177,N_27400,N_26098);
nor UO_178 (O_178,N_29738,N_25378);
and UO_179 (O_179,N_25933,N_27424);
nand UO_180 (O_180,N_27702,N_26231);
and UO_181 (O_181,N_26044,N_28433);
nor UO_182 (O_182,N_27522,N_26574);
or UO_183 (O_183,N_28791,N_29141);
or UO_184 (O_184,N_26527,N_26179);
nor UO_185 (O_185,N_26583,N_26280);
and UO_186 (O_186,N_29946,N_25251);
nand UO_187 (O_187,N_28986,N_29524);
xor UO_188 (O_188,N_26696,N_27369);
xor UO_189 (O_189,N_27379,N_25178);
xnor UO_190 (O_190,N_29094,N_29403);
nand UO_191 (O_191,N_28906,N_28903);
or UO_192 (O_192,N_28871,N_25049);
xor UO_193 (O_193,N_26154,N_27781);
nand UO_194 (O_194,N_25968,N_29823);
and UO_195 (O_195,N_25888,N_28089);
xor UO_196 (O_196,N_26956,N_28109);
nor UO_197 (O_197,N_25447,N_26773);
nor UO_198 (O_198,N_26163,N_28454);
or UO_199 (O_199,N_26831,N_25938);
and UO_200 (O_200,N_28624,N_27256);
and UO_201 (O_201,N_27714,N_28221);
nor UO_202 (O_202,N_27383,N_26055);
or UO_203 (O_203,N_28772,N_29003);
xor UO_204 (O_204,N_29147,N_25501);
nor UO_205 (O_205,N_28948,N_25239);
nor UO_206 (O_206,N_26175,N_28296);
nand UO_207 (O_207,N_27115,N_28766);
nand UO_208 (O_208,N_26871,N_27042);
nand UO_209 (O_209,N_26517,N_28896);
xor UO_210 (O_210,N_27512,N_28962);
nor UO_211 (O_211,N_26499,N_26269);
xnor UO_212 (O_212,N_28771,N_27620);
nand UO_213 (O_213,N_28997,N_29467);
and UO_214 (O_214,N_29229,N_28987);
xnor UO_215 (O_215,N_27765,N_28483);
nor UO_216 (O_216,N_26353,N_29744);
nor UO_217 (O_217,N_25006,N_27005);
and UO_218 (O_218,N_27944,N_27477);
nand UO_219 (O_219,N_26565,N_26504);
or UO_220 (O_220,N_28778,N_25921);
or UO_221 (O_221,N_28123,N_25379);
nand UO_222 (O_222,N_27544,N_28084);
or UO_223 (O_223,N_27230,N_26564);
xnor UO_224 (O_224,N_28032,N_29768);
or UO_225 (O_225,N_26680,N_27076);
and UO_226 (O_226,N_29192,N_29614);
nand UO_227 (O_227,N_28899,N_26065);
or UO_228 (O_228,N_28211,N_27546);
xnor UO_229 (O_229,N_29257,N_27125);
nand UO_230 (O_230,N_25951,N_29228);
or UO_231 (O_231,N_26078,N_28353);
xnor UO_232 (O_232,N_26771,N_29882);
nand UO_233 (O_233,N_28270,N_27540);
and UO_234 (O_234,N_26165,N_29691);
xnor UO_235 (O_235,N_27907,N_29042);
or UO_236 (O_236,N_26041,N_29729);
and UO_237 (O_237,N_29360,N_29956);
xnor UO_238 (O_238,N_29364,N_28417);
xor UO_239 (O_239,N_26144,N_25808);
nand UO_240 (O_240,N_26657,N_27979);
and UO_241 (O_241,N_26100,N_26438);
nand UO_242 (O_242,N_25169,N_29827);
nor UO_243 (O_243,N_25325,N_25037);
nand UO_244 (O_244,N_25026,N_25183);
or UO_245 (O_245,N_29848,N_26169);
and UO_246 (O_246,N_28447,N_26611);
nor UO_247 (O_247,N_26545,N_27959);
and UO_248 (O_248,N_26199,N_27356);
and UO_249 (O_249,N_25821,N_27682);
nor UO_250 (O_250,N_26514,N_28969);
nand UO_251 (O_251,N_25439,N_25453);
or UO_252 (O_252,N_26976,N_26810);
xnor UO_253 (O_253,N_28297,N_26477);
nand UO_254 (O_254,N_26377,N_28373);
or UO_255 (O_255,N_25740,N_27945);
nor UO_256 (O_256,N_25722,N_29988);
xor UO_257 (O_257,N_27293,N_29086);
nand UO_258 (O_258,N_27989,N_27277);
nand UO_259 (O_259,N_28477,N_28430);
and UO_260 (O_260,N_29440,N_25463);
or UO_261 (O_261,N_27127,N_29815);
or UO_262 (O_262,N_25963,N_28007);
or UO_263 (O_263,N_28146,N_25749);
and UO_264 (O_264,N_26413,N_25929);
nand UO_265 (O_265,N_29661,N_29680);
or UO_266 (O_266,N_27319,N_27044);
and UO_267 (O_267,N_25024,N_25606);
and UO_268 (O_268,N_27866,N_27964);
xnor UO_269 (O_269,N_26376,N_27496);
or UO_270 (O_270,N_28410,N_28328);
or UO_271 (O_271,N_28654,N_26540);
xor UO_272 (O_272,N_28266,N_25721);
nor UO_273 (O_273,N_25166,N_26177);
xor UO_274 (O_274,N_28634,N_27228);
xor UO_275 (O_275,N_25413,N_25323);
xor UO_276 (O_276,N_25159,N_29185);
xor UO_277 (O_277,N_29335,N_28075);
nand UO_278 (O_278,N_25471,N_29746);
xnor UO_279 (O_279,N_25916,N_29280);
nand UO_280 (O_280,N_28779,N_27645);
or UO_281 (O_281,N_25341,N_27862);
or UO_282 (O_282,N_27032,N_29845);
or UO_283 (O_283,N_27161,N_29643);
and UO_284 (O_284,N_25880,N_27108);
nor UO_285 (O_285,N_29146,N_25555);
or UO_286 (O_286,N_28456,N_26166);
and UO_287 (O_287,N_27285,N_26620);
and UO_288 (O_288,N_25699,N_26474);
xor UO_289 (O_289,N_25138,N_29584);
xnor UO_290 (O_290,N_27650,N_27478);
or UO_291 (O_291,N_29516,N_29758);
xor UO_292 (O_292,N_28998,N_26740);
or UO_293 (O_293,N_27527,N_26228);
or UO_294 (O_294,N_29557,N_27794);
nor UO_295 (O_295,N_25393,N_29298);
nand UO_296 (O_296,N_29069,N_29809);
nor UO_297 (O_297,N_28898,N_27810);
nand UO_298 (O_298,N_29373,N_29405);
nand UO_299 (O_299,N_26149,N_28996);
nand UO_300 (O_300,N_25039,N_28196);
nand UO_301 (O_301,N_27829,N_29537);
xnor UO_302 (O_302,N_25527,N_28354);
nand UO_303 (O_303,N_28814,N_29262);
nand UO_304 (O_304,N_28846,N_28048);
nor UO_305 (O_305,N_25521,N_27479);
nor UO_306 (O_306,N_28602,N_28983);
nand UO_307 (O_307,N_28912,N_28406);
nor UO_308 (O_308,N_29365,N_29077);
xnor UO_309 (O_309,N_28191,N_27800);
xnor UO_310 (O_310,N_27080,N_28439);
or UO_311 (O_311,N_29453,N_25080);
xnor UO_312 (O_312,N_25110,N_25181);
nor UO_313 (O_313,N_28632,N_26210);
nor UO_314 (O_314,N_28054,N_26987);
xor UO_315 (O_315,N_29450,N_27494);
nor UO_316 (O_316,N_27891,N_29843);
xor UO_317 (O_317,N_29561,N_27088);
xnor UO_318 (O_318,N_26042,N_28520);
xnor UO_319 (O_319,N_26450,N_27545);
xnor UO_320 (O_320,N_28474,N_27261);
nand UO_321 (O_321,N_25505,N_27466);
xnor UO_322 (O_322,N_26315,N_26965);
or UO_323 (O_323,N_25544,N_29784);
nand UO_324 (O_324,N_29321,N_26535);
xor UO_325 (O_325,N_27428,N_26996);
xnor UO_326 (O_326,N_25566,N_25846);
or UO_327 (O_327,N_25204,N_27365);
or UO_328 (O_328,N_25269,N_29984);
nor UO_329 (O_329,N_25476,N_28770);
or UO_330 (O_330,N_27476,N_29277);
and UO_331 (O_331,N_27733,N_29079);
nor UO_332 (O_332,N_26350,N_25779);
or UO_333 (O_333,N_29322,N_28630);
nand UO_334 (O_334,N_25798,N_29439);
nor UO_335 (O_335,N_29356,N_27766);
nand UO_336 (O_336,N_27890,N_27035);
and UO_337 (O_337,N_27729,N_26648);
or UO_338 (O_338,N_25857,N_28115);
or UO_339 (O_339,N_28990,N_29302);
or UO_340 (O_340,N_27166,N_28156);
or UO_341 (O_341,N_27037,N_26913);
nor UO_342 (O_342,N_27500,N_29551);
nand UO_343 (O_343,N_28358,N_27529);
nand UO_344 (O_344,N_27220,N_25106);
xor UO_345 (O_345,N_26772,N_29276);
or UO_346 (O_346,N_29272,N_27071);
nand UO_347 (O_347,N_28227,N_25685);
nor UO_348 (O_348,N_26389,N_29197);
xor UO_349 (O_349,N_27904,N_26443);
nand UO_350 (O_350,N_27493,N_28677);
nand UO_351 (O_351,N_27008,N_27593);
or UO_352 (O_352,N_26001,N_28641);
or UO_353 (O_353,N_28182,N_29045);
nor UO_354 (O_354,N_28288,N_26462);
nor UO_355 (O_355,N_27562,N_28157);
xor UO_356 (O_356,N_29311,N_27187);
or UO_357 (O_357,N_27189,N_28485);
xnor UO_358 (O_358,N_25315,N_27858);
xnor UO_359 (O_359,N_29030,N_26973);
xnor UO_360 (O_360,N_27069,N_25461);
nor UO_361 (O_361,N_25038,N_25990);
and UO_362 (O_362,N_29544,N_29662);
or UO_363 (O_363,N_29454,N_25708);
and UO_364 (O_364,N_28957,N_29244);
and UO_365 (O_365,N_28737,N_29760);
or UO_366 (O_366,N_26578,N_29451);
or UO_367 (O_367,N_28829,N_29745);
and UO_368 (O_368,N_27055,N_25876);
xnor UO_369 (O_369,N_26396,N_26512);
xnor UO_370 (O_370,N_28509,N_25474);
nor UO_371 (O_371,N_26161,N_26494);
xnor UO_372 (O_372,N_26638,N_28978);
nor UO_373 (O_373,N_27171,N_26752);
nand UO_374 (O_374,N_29029,N_25132);
nand UO_375 (O_375,N_29384,N_26254);
xor UO_376 (O_376,N_26975,N_28408);
nand UO_377 (O_377,N_26692,N_27583);
nor UO_378 (O_378,N_27421,N_25227);
or UO_379 (O_379,N_25173,N_25587);
and UO_380 (O_380,N_29979,N_28662);
xnor UO_381 (O_381,N_26039,N_28132);
and UO_382 (O_382,N_25569,N_28163);
or UO_383 (O_383,N_29100,N_29431);
and UO_384 (O_384,N_26126,N_25747);
or UO_385 (O_385,N_27611,N_29473);
and UO_386 (O_386,N_25455,N_28331);
and UO_387 (O_387,N_29955,N_26776);
xnor UO_388 (O_388,N_29116,N_28037);
nor UO_389 (O_389,N_29786,N_27322);
or UO_390 (O_390,N_27518,N_27920);
or UO_391 (O_391,N_25910,N_28181);
or UO_392 (O_392,N_27625,N_26652);
xor UO_393 (O_393,N_25119,N_29911);
or UO_394 (O_394,N_26856,N_27070);
nor UO_395 (O_395,N_29461,N_27960);
nand UO_396 (O_396,N_28045,N_26335);
or UO_397 (O_397,N_28611,N_25041);
xnor UO_398 (O_398,N_25875,N_26080);
nand UO_399 (O_399,N_27672,N_26854);
or UO_400 (O_400,N_28065,N_29967);
nand UO_401 (O_401,N_28754,N_27668);
or UO_402 (O_402,N_26851,N_26857);
or UO_403 (O_403,N_27610,N_26287);
nand UO_404 (O_404,N_28467,N_28850);
or UO_405 (O_405,N_28968,N_29620);
or UO_406 (O_406,N_26519,N_29130);
nor UO_407 (O_407,N_27254,N_25503);
nand UO_408 (O_408,N_25398,N_25945);
nor UO_409 (O_409,N_27252,N_26616);
and UO_410 (O_410,N_25422,N_27399);
or UO_411 (O_411,N_26466,N_25943);
xnor UO_412 (O_412,N_28568,N_27515);
and UO_413 (O_413,N_28133,N_27779);
and UO_414 (O_414,N_27553,N_28575);
nor UO_415 (O_415,N_27885,N_25705);
and UO_416 (O_416,N_25290,N_28744);
xor UO_417 (O_417,N_28047,N_25369);
xor UO_418 (O_418,N_27950,N_25959);
and UO_419 (O_419,N_26841,N_25688);
xnor UO_420 (O_420,N_29944,N_29177);
nor UO_421 (O_421,N_27910,N_29196);
nor UO_422 (O_422,N_27996,N_29675);
nor UO_423 (O_423,N_25291,N_28971);
nand UO_424 (O_424,N_26989,N_26689);
nand UO_425 (O_425,N_25553,N_29133);
xor UO_426 (O_426,N_28431,N_29987);
or UO_427 (O_427,N_29857,N_27456);
nor UO_428 (O_428,N_26123,N_27887);
xnor UO_429 (O_429,N_29336,N_26451);
or UO_430 (O_430,N_25053,N_29238);
nand UO_431 (O_431,N_27889,N_26129);
xor UO_432 (O_432,N_25470,N_29137);
or UO_433 (O_433,N_26467,N_25732);
nor UO_434 (O_434,N_26838,N_26265);
or UO_435 (O_435,N_25155,N_27903);
nor UO_436 (O_436,N_26272,N_29400);
or UO_437 (O_437,N_29598,N_27865);
nor UO_438 (O_438,N_28205,N_26381);
xnor UO_439 (O_439,N_27826,N_27357);
and UO_440 (O_440,N_25619,N_26829);
nor UO_441 (O_441,N_27977,N_28421);
nor UO_442 (O_442,N_29796,N_29251);
nor UO_443 (O_443,N_27231,N_27533);
nor UO_444 (O_444,N_29858,N_27701);
and UO_445 (O_445,N_28803,N_28334);
xnor UO_446 (O_446,N_27345,N_28972);
xnor UO_447 (O_447,N_29793,N_29330);
nor UO_448 (O_448,N_25842,N_28755);
and UO_449 (O_449,N_25113,N_27151);
nor UO_450 (O_450,N_26878,N_29309);
nor UO_451 (O_451,N_26085,N_28060);
and UO_452 (O_452,N_29660,N_26083);
or UO_453 (O_453,N_26507,N_27731);
and UO_454 (O_454,N_25706,N_25276);
nor UO_455 (O_455,N_27876,N_26992);
xor UO_456 (O_456,N_28072,N_26985);
or UO_457 (O_457,N_28925,N_25502);
xor UO_458 (O_458,N_26698,N_25033);
nand UO_459 (O_459,N_26770,N_27306);
and UO_460 (O_460,N_25901,N_27911);
and UO_461 (O_461,N_27801,N_27856);
xor UO_462 (O_462,N_27122,N_26792);
nor UO_463 (O_463,N_27848,N_27260);
and UO_464 (O_464,N_26029,N_27396);
or UO_465 (O_465,N_27949,N_26130);
nor UO_466 (O_466,N_25366,N_25666);
or UO_467 (O_467,N_25971,N_27646);
and UO_468 (O_468,N_27867,N_28016);
nand UO_469 (O_469,N_26475,N_26662);
or UO_470 (O_470,N_29287,N_29780);
and UO_471 (O_471,N_29520,N_27208);
and UO_472 (O_472,N_29171,N_26298);
nand UO_473 (O_473,N_28411,N_28204);
or UO_474 (O_474,N_26384,N_28481);
or UO_475 (O_475,N_27391,N_25001);
and UO_476 (O_476,N_25022,N_25232);
xor UO_477 (O_477,N_27739,N_25099);
xor UO_478 (O_478,N_28419,N_27495);
xnor UO_479 (O_479,N_28683,N_29070);
xnor UO_480 (O_480,N_26623,N_28255);
xnor UO_481 (O_481,N_25782,N_25683);
xnor UO_482 (O_482,N_28936,N_29297);
and UO_483 (O_483,N_26522,N_25440);
or UO_484 (O_484,N_29774,N_27587);
and UO_485 (O_485,N_29981,N_28543);
xnor UO_486 (O_486,N_26515,N_27393);
nor UO_487 (O_487,N_25238,N_25283);
or UO_488 (O_488,N_29688,N_26355);
nor UO_489 (O_489,N_29555,N_26945);
nor UO_490 (O_490,N_29409,N_28752);
nand UO_491 (O_491,N_28079,N_27327);
or UO_492 (O_492,N_27215,N_25564);
xor UO_493 (O_493,N_26155,N_26908);
nand UO_494 (O_494,N_28550,N_27259);
nand UO_495 (O_495,N_29011,N_25804);
or UO_496 (O_496,N_28688,N_28859);
xor UO_497 (O_497,N_25152,N_25042);
nor UO_498 (O_498,N_25142,N_28476);
nand UO_499 (O_499,N_25426,N_28183);
and UO_500 (O_500,N_26900,N_26602);
and UO_501 (O_501,N_27570,N_29676);
or UO_502 (O_502,N_28866,N_25278);
nor UO_503 (O_503,N_27068,N_26296);
or UO_504 (O_504,N_27269,N_27089);
or UO_505 (O_505,N_29698,N_26882);
nor UO_506 (O_506,N_25858,N_28389);
nand UO_507 (O_507,N_27730,N_25500);
xnor UO_508 (O_508,N_26595,N_26232);
and UO_509 (O_509,N_25151,N_26744);
nand UO_510 (O_510,N_26138,N_28923);
or UO_511 (O_511,N_29462,N_27175);
and UO_512 (O_512,N_26994,N_27309);
and UO_513 (O_513,N_27286,N_25240);
nand UO_514 (O_514,N_26730,N_27818);
nor UO_515 (O_515,N_27660,N_26991);
xnor UO_516 (O_516,N_26877,N_27508);
and UO_517 (O_517,N_25852,N_29264);
or UO_518 (O_518,N_26453,N_28789);
and UO_519 (O_519,N_29091,N_26759);
or UO_520 (O_520,N_26509,N_26262);
nand UO_521 (O_521,N_25467,N_29805);
or UO_522 (O_522,N_28979,N_29393);
and UO_523 (O_523,N_25019,N_29378);
xor UO_524 (O_524,N_29076,N_28908);
xor UO_525 (O_525,N_27366,N_27460);
nand UO_526 (O_526,N_27700,N_28346);
or UO_527 (O_527,N_27116,N_29463);
and UO_528 (O_528,N_26035,N_27382);
or UO_529 (O_529,N_28096,N_29396);
nand UO_530 (O_530,N_28284,N_26747);
nor UO_531 (O_531,N_28235,N_27967);
or UO_532 (O_532,N_28666,N_29190);
nand UO_533 (O_533,N_28203,N_26146);
nor UO_534 (O_534,N_25691,N_29588);
or UO_535 (O_535,N_28011,N_25194);
and UO_536 (O_536,N_27689,N_28840);
nor UO_537 (O_537,N_29268,N_26089);
nand UO_538 (O_538,N_27673,N_25082);
xor UO_539 (O_539,N_27419,N_26694);
nor UO_540 (O_540,N_28946,N_28815);
and UO_541 (O_541,N_27706,N_25743);
nor UO_542 (O_542,N_26673,N_25466);
nor UO_543 (O_543,N_27567,N_26308);
or UO_544 (O_544,N_29507,N_28868);
and UO_545 (O_545,N_27446,N_27420);
xor UO_546 (O_546,N_25556,N_25252);
nor UO_547 (O_547,N_29172,N_27839);
nor UO_548 (O_548,N_26449,N_26618);
and UO_549 (O_549,N_27033,N_28035);
nand UO_550 (O_550,N_26892,N_25955);
nand UO_551 (O_551,N_25522,N_25816);
or UO_552 (O_552,N_25177,N_28725);
or UO_553 (O_553,N_27838,N_26513);
xnor UO_554 (O_554,N_28186,N_28907);
or UO_555 (O_555,N_25187,N_28152);
nand UO_556 (O_556,N_26142,N_28193);
xor UO_557 (O_557,N_26518,N_29333);
or UO_558 (O_558,N_26132,N_27359);
and UO_559 (O_559,N_25615,N_29053);
nand UO_560 (O_560,N_28658,N_25891);
and UO_561 (O_561,N_28518,N_28381);
or UO_562 (O_562,N_25456,N_28159);
nor UO_563 (O_563,N_29299,N_28885);
nor UO_564 (O_564,N_29634,N_29021);
or UO_565 (O_565,N_29678,N_26329);
and UO_566 (O_566,N_27321,N_25158);
xor UO_567 (O_567,N_27782,N_26713);
or UO_568 (O_568,N_26300,N_27929);
nor UO_569 (O_569,N_29436,N_26387);
or UO_570 (O_570,N_27146,N_29166);
or UO_571 (O_571,N_27516,N_27853);
or UO_572 (O_572,N_26173,N_25718);
nor UO_573 (O_573,N_27995,N_25307);
nor UO_574 (O_574,N_25056,N_26855);
and UO_575 (O_575,N_28295,N_26847);
and UO_576 (O_576,N_25727,N_28895);
and UO_577 (O_577,N_25117,N_25812);
and UO_578 (O_578,N_29124,N_27018);
nor UO_579 (O_579,N_26802,N_28164);
or UO_580 (O_580,N_27126,N_25837);
nand UO_581 (O_581,N_26567,N_25385);
or UO_582 (O_582,N_29708,N_26576);
or UO_583 (O_583,N_27803,N_29719);
nand UO_584 (O_584,N_27506,N_27767);
xnor UO_585 (O_585,N_28073,N_27112);
nand UO_586 (O_586,N_27922,N_28781);
or UO_587 (O_587,N_27096,N_28922);
xor UO_588 (O_588,N_29150,N_28067);
nor UO_589 (O_589,N_29418,N_28083);
and UO_590 (O_590,N_26815,N_28504);
and UO_591 (O_591,N_26062,N_27000);
or UO_592 (O_592,N_25927,N_25321);
and UO_593 (O_593,N_25516,N_27007);
nor UO_594 (O_594,N_26071,N_25005);
or UO_595 (O_595,N_27784,N_28993);
or UO_596 (O_596,N_27627,N_29890);
nor UO_597 (O_597,N_27902,N_28339);
or UO_598 (O_598,N_27772,N_28349);
nor UO_599 (O_599,N_26593,N_28625);
xnor UO_600 (O_600,N_28705,N_26120);
and UO_601 (O_601,N_26922,N_28900);
and UO_602 (O_602,N_29355,N_27915);
and UO_603 (O_603,N_26731,N_28913);
nor UO_604 (O_604,N_27678,N_25625);
nor UO_605 (O_605,N_26709,N_29087);
nand UO_606 (O_606,N_28555,N_25603);
or UO_607 (O_607,N_25709,N_29271);
and UO_608 (O_608,N_29059,N_28951);
xnor UO_609 (O_609,N_29898,N_27556);
nor UO_610 (O_610,N_28617,N_25563);
nor UO_611 (O_611,N_26667,N_26984);
nand UO_612 (O_612,N_25198,N_29145);
nand UO_613 (O_613,N_29479,N_27128);
nand UO_614 (O_614,N_27555,N_29031);
nor UO_615 (O_615,N_28511,N_27290);
nor UO_616 (O_616,N_25524,N_28434);
or UO_617 (O_617,N_26763,N_25118);
and UO_618 (O_618,N_27452,N_27401);
and UO_619 (O_619,N_26880,N_29230);
or UO_620 (O_620,N_29160,N_28596);
and UO_621 (O_621,N_25964,N_26302);
xnor UO_622 (O_622,N_28386,N_28017);
nand UO_623 (O_623,N_26777,N_25230);
xnor UO_624 (O_624,N_29015,N_25414);
and UO_625 (O_625,N_26629,N_26082);
and UO_626 (O_626,N_26094,N_26095);
or UO_627 (O_627,N_26950,N_25735);
or UO_628 (O_628,N_29940,N_26313);
or UO_629 (O_629,N_25078,N_28404);
xor UO_630 (O_630,N_28606,N_27082);
xor UO_631 (O_631,N_28673,N_26721);
nor UO_632 (O_632,N_29095,N_29879);
or UO_633 (O_633,N_27750,N_29222);
and UO_634 (O_634,N_29304,N_27058);
and UO_635 (O_635,N_29685,N_26553);
and UO_636 (O_636,N_29813,N_26186);
xnor UO_637 (O_637,N_29702,N_27087);
nand UO_638 (O_638,N_25135,N_29476);
nand UO_639 (O_639,N_25612,N_25088);
or UO_640 (O_640,N_25179,N_29159);
nand UO_641 (O_641,N_28260,N_27759);
or UO_642 (O_642,N_26153,N_29155);
or UO_643 (O_643,N_26195,N_26170);
nor UO_644 (O_644,N_27693,N_25755);
nand UO_645 (O_645,N_26291,N_27155);
or UO_646 (O_646,N_28144,N_27732);
and UO_647 (O_647,N_29803,N_28765);
or UO_648 (O_648,N_28087,N_25141);
or UO_649 (O_649,N_29664,N_27144);
nand UO_650 (O_650,N_28427,N_25753);
xor UO_651 (O_651,N_29819,N_26448);
and UO_652 (O_652,N_25047,N_29647);
xor UO_653 (O_653,N_27975,N_26480);
xnor UO_654 (O_654,N_25174,N_25271);
or UO_655 (O_655,N_29687,N_26970);
nand UO_656 (O_656,N_25539,N_26294);
and UO_657 (O_657,N_26822,N_25308);
nand UO_658 (O_658,N_29876,N_26794);
nor UO_659 (O_659,N_26277,N_27734);
xnor UO_660 (O_660,N_28647,N_26097);
or UO_661 (O_661,N_25868,N_29093);
nand UO_662 (O_662,N_29118,N_28883);
nor UO_663 (O_663,N_27963,N_26157);
nor UO_664 (O_664,N_29218,N_26445);
and UO_665 (O_665,N_25419,N_28710);
xnor UO_666 (O_666,N_25698,N_29044);
or UO_667 (O_667,N_29441,N_26585);
nor UO_668 (O_668,N_25188,N_28192);
xnor UO_669 (O_669,N_25277,N_25221);
xnor UO_670 (O_670,N_26551,N_26539);
xor UO_671 (O_671,N_25654,N_28453);
nor UO_672 (O_672,N_26557,N_25180);
or UO_673 (O_673,N_25748,N_29447);
nand UO_674 (O_674,N_28076,N_26853);
or UO_675 (O_675,N_25562,N_28140);
and UO_676 (O_676,N_28692,N_28232);
nand UO_677 (O_677,N_25879,N_27751);
and UO_678 (O_678,N_25604,N_28370);
or UO_679 (O_679,N_25484,N_28873);
or UO_680 (O_680,N_29478,N_27461);
xor UO_681 (O_681,N_26889,N_29404);
nor UO_682 (O_682,N_25206,N_26279);
and UO_683 (O_683,N_25860,N_27469);
and UO_684 (O_684,N_28416,N_28118);
and UO_685 (O_685,N_29652,N_27685);
and UO_686 (O_686,N_27737,N_28052);
and UO_687 (O_687,N_28642,N_25084);
and UO_688 (O_688,N_28494,N_26766);
and UO_689 (O_689,N_26779,N_25040);
and UO_690 (O_690,N_25673,N_29085);
nor UO_691 (O_691,N_25982,N_27062);
or UO_692 (O_692,N_27884,N_25850);
nor UO_693 (O_693,N_26686,N_29669);
xor UO_694 (O_694,N_29111,N_27809);
xnor UO_695 (O_695,N_28315,N_28388);
nand UO_696 (O_696,N_29562,N_26971);
or UO_697 (O_697,N_28712,N_28418);
and UO_698 (O_698,N_25534,N_29239);
or UO_699 (O_699,N_25356,N_27755);
nand UO_700 (O_700,N_25541,N_28881);
xnor UO_701 (O_701,N_27925,N_29416);
nor UO_702 (O_702,N_27575,N_27244);
and UO_703 (O_703,N_27333,N_25789);
xnor UO_704 (O_704,N_28878,N_25375);
xnor UO_705 (O_705,N_28179,N_29549);
nand UO_706 (O_706,N_25870,N_29434);
or UO_707 (O_707,N_25272,N_29609);
or UO_708 (O_708,N_25093,N_25361);
xnor UO_709 (O_709,N_29089,N_27787);
nand UO_710 (O_710,N_26844,N_26250);
or UO_711 (O_711,N_26104,N_26658);
nand UO_712 (O_712,N_28579,N_25658);
nand UO_713 (O_713,N_25928,N_26328);
xnor UO_714 (O_714,N_29343,N_27361);
or UO_715 (O_715,N_28320,N_27811);
xor UO_716 (O_716,N_25998,N_29638);
and UO_717 (O_717,N_25249,N_28524);
nor UO_718 (O_718,N_28924,N_25021);
and UO_719 (O_719,N_27100,N_25386);
xor UO_720 (O_720,N_29554,N_27786);
and UO_721 (O_721,N_26193,N_29289);
nor UO_722 (O_722,N_25263,N_25613);
nor UO_723 (O_723,N_28828,N_29965);
nand UO_724 (O_724,N_26205,N_25777);
xnor UO_725 (O_725,N_25596,N_25364);
or UO_726 (O_726,N_25176,N_28131);
xor UO_727 (O_727,N_27565,N_29512);
xnor UO_728 (O_728,N_27117,N_27248);
and UO_729 (O_729,N_25552,N_28835);
nor UO_730 (O_730,N_28210,N_26244);
xnor UO_731 (O_731,N_25073,N_29569);
and UO_732 (O_732,N_26233,N_27659);
and UO_733 (O_733,N_26874,N_28158);
nor UO_734 (O_734,N_27951,N_26040);
nand UO_735 (O_735,N_26953,N_29923);
nand UO_736 (O_736,N_25760,N_25231);
xor UO_737 (O_737,N_26774,N_26897);
xor UO_738 (O_738,N_26860,N_26678);
or UO_739 (O_739,N_27595,N_28603);
xor UO_740 (O_740,N_29993,N_25617);
xnor UO_741 (O_741,N_25497,N_26066);
xor UO_742 (O_742,N_28587,N_26172);
xor UO_743 (O_743,N_29474,N_25646);
and UO_744 (O_744,N_25060,N_26666);
or UO_745 (O_745,N_25855,N_27820);
and UO_746 (O_746,N_27823,N_28243);
and UO_747 (O_747,N_29927,N_27749);
nor UO_748 (O_748,N_26724,N_29475);
nand UO_749 (O_749,N_27677,N_29619);
or UO_750 (O_750,N_25067,N_28920);
nand UO_751 (O_751,N_28317,N_27704);
xnor UO_752 (O_752,N_29377,N_28278);
nor UO_753 (O_753,N_27653,N_27240);
nand UO_754 (O_754,N_27339,N_26869);
nand UO_755 (O_755,N_25784,N_25624);
and UO_756 (O_756,N_26858,N_29682);
nand UO_757 (O_757,N_26995,N_26790);
xor UO_758 (O_758,N_26821,N_27030);
xor UO_759 (O_759,N_29973,N_28548);
xnor UO_760 (O_760,N_27074,N_29724);
xnor UO_761 (O_761,N_28853,N_29278);
or UO_762 (O_762,N_29253,N_28733);
xor UO_763 (O_763,N_25608,N_29072);
nor UO_764 (O_764,N_29258,N_26612);
nand UO_765 (O_765,N_27806,N_25629);
or UO_766 (O_766,N_26562,N_28013);
nor UO_767 (O_767,N_28491,N_26780);
or UO_768 (O_768,N_25840,N_29179);
xnor UO_769 (O_769,N_26898,N_26192);
and UO_770 (O_770,N_27937,N_25565);
nor UO_771 (O_771,N_28031,N_26603);
nand UO_772 (O_772,N_26799,N_25669);
nor UO_773 (O_773,N_29217,N_29349);
xnor UO_774 (O_774,N_25884,N_28874);
nor UO_775 (O_775,N_29284,N_26349);
or UO_776 (O_776,N_27436,N_27085);
or UO_777 (O_777,N_26086,N_28826);
or UO_778 (O_778,N_28992,N_25157);
xor UO_779 (O_779,N_29107,N_29938);
nand UO_780 (O_780,N_28019,N_27615);
nor UO_781 (O_781,N_25014,N_27760);
or UO_782 (O_782,N_25091,N_27019);
or UO_783 (O_783,N_29423,N_28837);
or UO_784 (O_784,N_25069,N_27013);
xnor UO_785 (O_785,N_25279,N_27232);
xor UO_786 (O_786,N_29009,N_26124);
and UO_787 (O_787,N_29917,N_25510);
and UO_788 (O_788,N_27973,N_27987);
and UO_789 (O_789,N_25599,N_26151);
nand UO_790 (O_790,N_25761,N_29064);
nor UO_791 (O_791,N_25992,N_25872);
and UO_792 (O_792,N_25792,N_27186);
nor UO_793 (O_793,N_25444,N_27006);
nor UO_794 (O_794,N_25601,N_26278);
nor UO_795 (O_795,N_27774,N_28166);
nand UO_796 (O_796,N_26164,N_25358);
nand UO_797 (O_797,N_25383,N_26339);
or UO_798 (O_798,N_25967,N_28463);
nor UO_799 (O_799,N_25211,N_28327);
or UO_800 (O_800,N_29249,N_25288);
nand UO_801 (O_801,N_28757,N_26397);
nor UO_802 (O_802,N_28461,N_25614);
or UO_803 (O_803,N_27370,N_27622);
or UO_804 (O_804,N_25340,N_28294);
xor UO_805 (O_805,N_27047,N_28351);
xor UO_806 (O_806,N_26103,N_26804);
and UO_807 (O_807,N_27348,N_28487);
nand UO_808 (O_808,N_25742,N_29637);
and UO_809 (O_809,N_26461,N_27928);
xor UO_810 (O_810,N_28413,N_25207);
nand UO_811 (O_811,N_26714,N_26032);
and UO_812 (O_812,N_26152,N_26536);
nand UO_813 (O_813,N_25514,N_28750);
nor UO_814 (O_814,N_27793,N_25570);
or UO_815 (O_815,N_29325,N_28290);
xor UO_816 (O_816,N_26746,N_26361);
nor UO_817 (O_817,N_29157,N_25882);
xnor UO_818 (O_818,N_26293,N_28120);
nor UO_819 (O_819,N_29816,N_29830);
and UO_820 (O_820,N_28092,N_27713);
nand UO_821 (O_821,N_29666,N_26702);
xor UO_822 (O_822,N_26715,N_26870);
or UO_823 (O_823,N_28559,N_29722);
xor UO_824 (O_824,N_29406,N_28030);
or UO_825 (O_825,N_27429,N_28535);
nand UO_826 (O_826,N_27897,N_25745);
and UO_827 (O_827,N_25273,N_29580);
nor UO_828 (O_828,N_29048,N_25417);
xor UO_829 (O_829,N_27221,N_28333);
or UO_830 (O_830,N_28136,N_29515);
nor UO_831 (O_831,N_25253,N_28631);
nor UO_832 (O_832,N_26716,N_28457);
nor UO_833 (O_833,N_29023,N_28578);
or UO_834 (O_834,N_27275,N_26619);
and UO_835 (O_835,N_25436,N_29672);
or UO_836 (O_836,N_27031,N_25725);
nor UO_837 (O_837,N_29567,N_25153);
nand UO_838 (O_838,N_25498,N_26485);
and UO_839 (O_839,N_27482,N_28249);
and UO_840 (O_840,N_26656,N_25744);
nor UO_841 (O_841,N_29395,N_26418);
and UO_842 (O_842,N_29285,N_26783);
or UO_843 (O_843,N_27084,N_27024);
nor UO_844 (O_844,N_27572,N_26317);
and UO_845 (O_845,N_26481,N_27745);
nor UO_846 (O_846,N_25558,N_29380);
and UO_847 (O_847,N_27184,N_29231);
xor UO_848 (O_848,N_26180,N_28607);
and UO_849 (O_849,N_27667,N_27236);
and UO_850 (O_850,N_29402,N_25543);
xor UO_851 (O_851,N_26782,N_28257);
xnor UO_852 (O_852,N_27060,N_29376);
nor UO_853 (O_853,N_27993,N_27796);
or UO_854 (O_854,N_27307,N_28887);
nor UO_855 (O_855,N_29639,N_29167);
xor UO_856 (O_856,N_29332,N_26227);
nand UO_857 (O_857,N_27778,N_25781);
and UO_858 (O_858,N_28739,N_28656);
xnor UO_859 (O_859,N_27754,N_28198);
xor UO_860 (O_860,N_29982,N_29046);
or UO_861 (O_861,N_27325,N_28502);
nor UO_862 (O_862,N_25292,N_25663);
nor UO_863 (O_863,N_29777,N_25316);
xor UO_864 (O_864,N_25621,N_29027);
nand UO_865 (O_865,N_29200,N_28190);
and UO_866 (O_866,N_29521,N_29968);
xnor UO_867 (O_867,N_28756,N_26059);
nor UO_868 (O_868,N_26076,N_29556);
nand UO_869 (O_869,N_27020,N_25387);
xor UO_870 (O_870,N_29178,N_29424);
and UO_871 (O_871,N_29849,N_28581);
nor UO_872 (O_872,N_28777,N_28595);
xnor UO_873 (O_873,N_29657,N_25653);
or UO_874 (O_874,N_27970,N_26888);
or UO_875 (O_875,N_28961,N_25776);
nand UO_876 (O_876,N_28580,N_26344);
or UO_877 (O_877,N_25210,N_27203);
nand UO_878 (O_878,N_26352,N_29340);
nor UO_879 (O_879,N_29363,N_27156);
nand UO_880 (O_880,N_27093,N_28233);
nand UO_881 (O_881,N_27978,N_28300);
nand UO_882 (O_882,N_29694,N_28714);
and UO_883 (O_883,N_28661,N_27131);
or UO_884 (O_884,N_29368,N_26592);
or UO_885 (O_885,N_25764,N_27695);
and UO_886 (O_886,N_26031,N_28811);
nand UO_887 (O_887,N_28174,N_26712);
and UO_888 (O_888,N_26408,N_25410);
and UO_889 (O_889,N_25145,N_28911);
nand UO_890 (O_890,N_25217,N_29459);
or UO_891 (O_891,N_25048,N_29493);
nand UO_892 (O_892,N_26962,N_28208);
or UO_893 (O_893,N_28696,N_27986);
or UO_894 (O_894,N_26275,N_27272);
and UO_895 (O_895,N_27416,N_26379);
and UO_896 (O_896,N_26027,N_29248);
xor UO_897 (O_897,N_26803,N_26023);
xnor UO_898 (O_898,N_27139,N_27861);
or UO_899 (O_899,N_28665,N_26546);
xnor UO_900 (O_900,N_28836,N_25354);
or UO_901 (O_901,N_25681,N_26924);
nor UO_902 (O_902,N_27304,N_25954);
nor UO_903 (O_903,N_26681,N_29869);
and UO_904 (O_904,N_25317,N_25579);
xnor UO_905 (O_905,N_26582,N_25442);
nand UO_906 (O_906,N_25991,N_26064);
nand UO_907 (O_907,N_29627,N_29600);
and UO_908 (O_908,N_28218,N_29347);
or UO_909 (O_909,N_27021,N_26903);
nand UO_910 (O_910,N_29317,N_29480);
nor UO_911 (O_911,N_29591,N_28307);
and UO_912 (O_912,N_26789,N_26520);
or UO_913 (O_913,N_28376,N_26276);
or UO_914 (O_914,N_25778,N_29175);
nand UO_915 (O_915,N_25259,N_25715);
nand UO_916 (O_916,N_29818,N_28851);
nand UO_917 (O_917,N_28646,N_25486);
nand UO_918 (O_918,N_26492,N_29726);
or UO_919 (O_919,N_28805,N_25944);
and UO_920 (O_920,N_26428,N_29700);
xor UO_921 (O_921,N_28810,N_27194);
xnor UO_922 (O_922,N_26457,N_26605);
and UO_923 (O_923,N_27414,N_26817);
or UO_924 (O_924,N_29530,N_26118);
xnor UO_925 (O_925,N_27984,N_26135);
or UO_926 (O_926,N_25939,N_25847);
or UO_927 (O_927,N_26650,N_26690);
nor UO_928 (O_928,N_27758,N_26634);
nand UO_929 (O_929,N_26909,N_27385);
nand UO_930 (O_930,N_25512,N_25650);
or UO_931 (O_931,N_28890,N_27358);
xor UO_932 (O_932,N_29088,N_27218);
and UO_933 (O_933,N_26672,N_28407);
and UO_934 (O_934,N_29350,N_27101);
nand UO_935 (O_935,N_27776,N_27472);
or UO_936 (O_936,N_25342,N_29918);
or UO_937 (O_937,N_29206,N_25574);
and UO_938 (O_938,N_28228,N_27387);
xnor UO_939 (O_939,N_25089,N_26257);
nor UO_940 (O_940,N_29259,N_27113);
nor UO_941 (O_941,N_26182,N_27608);
or UO_942 (O_942,N_26655,N_29415);
or UO_943 (O_943,N_25679,N_29586);
xor UO_944 (O_944,N_29452,N_26663);
nor UO_945 (O_945,N_29975,N_25493);
or UO_946 (O_946,N_26204,N_27094);
nor UO_947 (O_947,N_27930,N_25724);
nand UO_948 (O_948,N_28038,N_26322);
or UO_949 (O_949,N_29002,N_27210);
or UO_950 (O_950,N_27990,N_25200);
nand UO_951 (O_951,N_28619,N_26580);
nor UO_952 (O_952,N_28390,N_27504);
nand UO_953 (O_953,N_25978,N_29008);
or UO_954 (O_954,N_28348,N_26586);
xnor UO_955 (O_955,N_26274,N_28893);
nand UO_956 (O_956,N_29314,N_26340);
nor UO_957 (O_957,N_29640,N_26720);
xnor UO_958 (O_958,N_26421,N_29590);
nor UO_959 (O_959,N_29096,N_26798);
nor UO_960 (O_960,N_27647,N_29351);
xor UO_961 (O_961,N_27243,N_27039);
nand UO_962 (O_962,N_29282,N_29419);
nor UO_963 (O_963,N_26114,N_27742);
xnor UO_964 (O_964,N_28711,N_26584);
xor UO_965 (O_965,N_29313,N_27699);
xor UO_966 (O_966,N_28918,N_25362);
xor UO_967 (O_967,N_27159,N_26865);
nand UO_968 (O_968,N_25011,N_28959);
nand UO_969 (O_969,N_25686,N_28762);
nand UO_970 (O_970,N_28834,N_27012);
or UO_971 (O_971,N_27384,N_26370);
nand UO_972 (O_972,N_26613,N_27688);
and UO_973 (O_973,N_27004,N_28445);
nand UO_974 (O_974,N_27842,N_29985);
xnor UO_975 (O_975,N_27141,N_29626);
nor UO_976 (O_976,N_25578,N_26944);
nor UO_977 (O_977,N_29303,N_28171);
or UO_978 (O_978,N_29615,N_26938);
or UO_979 (O_979,N_29041,N_29749);
nand UO_980 (O_980,N_27711,N_25548);
nand UO_981 (O_981,N_29899,N_27833);
xor UO_982 (O_982,N_25002,N_28891);
and UO_983 (O_983,N_27170,N_26581);
nor UO_984 (O_984,N_29616,N_28287);
or UO_985 (O_985,N_27107,N_27756);
nor UO_986 (O_986,N_25144,N_26862);
nand UO_987 (O_987,N_29789,N_25947);
xor UO_988 (O_988,N_28175,N_26326);
and UO_989 (O_989,N_26750,N_26416);
nand UO_990 (O_990,N_27198,N_28340);
and UO_991 (O_991,N_28577,N_28049);
xor UO_992 (O_992,N_27528,N_26247);
xor UO_993 (O_993,N_26659,N_25717);
nor UO_994 (O_994,N_27028,N_29458);
xor UO_995 (O_995,N_26506,N_27335);
xor UO_996 (O_996,N_27757,N_25443);
xor UO_997 (O_997,N_28994,N_27791);
nand UO_998 (O_998,N_26946,N_27449);
nor UO_999 (O_999,N_25495,N_28817);
and UO_1000 (O_1000,N_29432,N_27877);
nand UO_1001 (O_1001,N_25492,N_26437);
xor UO_1002 (O_1002,N_26359,N_26530);
or UO_1003 (O_1003,N_26834,N_26491);
nor UO_1004 (O_1004,N_25713,N_28039);
nand UO_1005 (O_1005,N_25874,N_27918);
and UO_1006 (O_1006,N_29936,N_26476);
nand UO_1007 (O_1007,N_25644,N_28222);
nor UO_1008 (O_1008,N_29629,N_27237);
nand UO_1009 (O_1009,N_29875,N_28077);
xor UO_1010 (O_1010,N_25499,N_27388);
nor UO_1011 (O_1011,N_25346,N_25692);
and UO_1012 (O_1012,N_25786,N_27135);
and UO_1013 (O_1013,N_28678,N_29267);
xnor UO_1014 (O_1014,N_27288,N_29635);
and UO_1015 (O_1015,N_26967,N_25134);
xor UO_1016 (O_1016,N_29741,N_28074);
xnor UO_1017 (O_1017,N_28337,N_28585);
and UO_1018 (O_1018,N_28314,N_25695);
nor UO_1019 (O_1019,N_29686,N_26670);
xnor UO_1020 (O_1020,N_25245,N_26840);
nand UO_1021 (O_1021,N_26524,N_27114);
and UO_1022 (O_1022,N_25661,N_28117);
nor UO_1023 (O_1023,N_28250,N_27497);
nor UO_1024 (O_1024,N_29862,N_28719);
nand UO_1025 (O_1025,N_27652,N_25452);
xnor UO_1026 (O_1026,N_27181,N_25680);
nand UO_1027 (O_1027,N_27315,N_25432);
and UO_1028 (O_1028,N_27078,N_28472);
nand UO_1029 (O_1029,N_26446,N_27762);
nor UO_1030 (O_1030,N_29958,N_29382);
or UO_1031 (O_1031,N_27454,N_25672);
and UO_1032 (O_1032,N_26289,N_27919);
or UO_1033 (O_1033,N_29019,N_25146);
nand UO_1034 (O_1034,N_25209,N_28248);
nand UO_1035 (O_1035,N_29608,N_26735);
xnor UO_1036 (O_1036,N_25430,N_25373);
nor UO_1037 (O_1037,N_29663,N_27453);
nand UO_1038 (O_1038,N_27417,N_27072);
and UO_1039 (O_1039,N_26249,N_29026);
nand UO_1040 (O_1040,N_28768,N_28542);
nand UO_1041 (O_1041,N_27296,N_26273);
nand UO_1042 (O_1042,N_27629,N_27654);
and UO_1043 (O_1043,N_27352,N_26426);
nor UO_1044 (O_1044,N_26572,N_25137);
and UO_1045 (O_1045,N_25075,N_26049);
or UO_1046 (O_1046,N_27690,N_26926);
xnor UO_1047 (O_1047,N_28571,N_28237);
nand UO_1048 (O_1048,N_27280,N_28858);
and UO_1049 (O_1049,N_29919,N_26048);
nand UO_1050 (O_1050,N_26067,N_26999);
and UO_1051 (O_1051,N_25806,N_26105);
or UO_1052 (O_1052,N_27628,N_29763);
nor UO_1053 (O_1053,N_26500,N_29606);
nor UO_1054 (O_1054,N_25071,N_28738);
xor UO_1055 (O_1055,N_26101,N_29080);
nor UO_1056 (O_1056,N_29573,N_28363);
nor UO_1057 (O_1057,N_25219,N_26000);
or UO_1058 (O_1058,N_27095,N_26941);
nand UO_1059 (O_1059,N_25116,N_25854);
nand UO_1060 (O_1060,N_28055,N_27434);
and UO_1061 (O_1061,N_27251,N_29817);
and UO_1062 (O_1062,N_29173,N_25787);
nand UO_1063 (O_1063,N_27642,N_25542);
and UO_1064 (O_1064,N_29861,N_27560);
nor UO_1065 (O_1065,N_28856,N_28942);
xor UO_1066 (O_1066,N_28636,N_29912);
nand UO_1067 (O_1067,N_26380,N_29017);
nand UO_1068 (O_1068,N_29306,N_28824);
and UO_1069 (O_1069,N_27537,N_26920);
xor UO_1070 (O_1070,N_28668,N_26420);
nand UO_1071 (O_1071,N_29889,N_29469);
or UO_1072 (O_1072,N_26145,N_26510);
or UO_1073 (O_1073,N_29223,N_28538);
or UO_1074 (O_1074,N_28761,N_29560);
or UO_1075 (O_1075,N_29667,N_28981);
xnor UO_1076 (O_1076,N_25032,N_25063);
nand UO_1077 (O_1077,N_29742,N_28383);
nand UO_1078 (O_1078,N_25023,N_25730);
or UO_1079 (O_1079,N_25168,N_25581);
nand UO_1080 (O_1080,N_28794,N_27870);
or UO_1081 (O_1081,N_29444,N_28239);
and UO_1082 (O_1082,N_27687,N_28306);
nand UO_1083 (O_1083,N_28558,N_28302);
nand UO_1084 (O_1084,N_28135,N_26543);
xor UO_1085 (O_1085,N_28528,N_25072);
nor UO_1086 (O_1086,N_25803,N_29885);
and UO_1087 (O_1087,N_28527,N_26134);
and UO_1088 (O_1088,N_28259,N_25100);
nand UO_1089 (O_1089,N_25639,N_29470);
and UO_1090 (O_1090,N_28621,N_29681);
nor UO_1091 (O_1091,N_29545,N_26534);
xnor UO_1092 (O_1092,N_27936,N_28143);
or UO_1093 (O_1093,N_25659,N_29052);
and UO_1094 (O_1094,N_29559,N_25923);
and UO_1095 (O_1095,N_25438,N_25958);
xor UO_1096 (O_1096,N_28062,N_29139);
or UO_1097 (O_1097,N_26675,N_26560);
nor UO_1098 (O_1098,N_27191,N_26357);
nor UO_1099 (O_1099,N_25511,N_28704);
nand UO_1100 (O_1100,N_25115,N_27120);
or UO_1101 (O_1101,N_27665,N_27773);
and UO_1102 (O_1102,N_26365,N_25111);
nor UO_1103 (O_1103,N_28635,N_28088);
nor UO_1104 (O_1104,N_25182,N_28310);
xor UO_1105 (O_1105,N_28268,N_27099);
or UO_1106 (O_1106,N_25487,N_26525);
and UO_1107 (O_1107,N_29645,N_25449);
and UO_1108 (O_1108,N_28450,N_25795);
or UO_1109 (O_1109,N_25222,N_25310);
nor UO_1110 (O_1110,N_29734,N_25919);
or UO_1111 (O_1111,N_27616,N_28180);
and UO_1112 (O_1112,N_27353,N_28283);
nor UO_1113 (O_1113,N_26122,N_29716);
nor UO_1114 (O_1114,N_25734,N_26737);
xor UO_1115 (O_1115,N_27405,N_27747);
and UO_1116 (O_1116,N_26478,N_27581);
xnor UO_1117 (O_1117,N_25866,N_26119);
nand UO_1118 (O_1118,N_26398,N_28787);
nor UO_1119 (O_1119,N_28282,N_29083);
nand UO_1120 (O_1120,N_29670,N_27859);
xor UO_1121 (O_1121,N_29630,N_27397);
and UO_1122 (O_1122,N_27864,N_27312);
nor UO_1123 (O_1123,N_29456,N_26470);
nor UO_1124 (O_1124,N_27670,N_28610);
nand UO_1125 (O_1125,N_27313,N_27814);
nand UO_1126 (O_1126,N_27444,N_26861);
nand UO_1127 (O_1127,N_26587,N_26148);
and UO_1128 (O_1128,N_27780,N_26820);
nor UO_1129 (O_1129,N_27510,N_29122);
nor UO_1130 (O_1130,N_25628,N_25297);
xnor UO_1131 (O_1131,N_25594,N_26901);
and UO_1132 (O_1132,N_28355,N_28448);
xor UO_1133 (O_1133,N_29189,N_25961);
nand UO_1134 (O_1134,N_29121,N_26823);
and UO_1135 (O_1135,N_26403,N_26948);
nand UO_1136 (O_1136,N_28944,N_27658);
nor UO_1137 (O_1137,N_26819,N_29293);
or UO_1138 (O_1138,N_28574,N_25160);
nand UO_1139 (O_1139,N_28150,N_29511);
nand UO_1140 (O_1140,N_29807,N_28801);
and UO_1141 (O_1141,N_28482,N_27300);
or UO_1142 (O_1142,N_29457,N_28552);
xnor UO_1143 (O_1143,N_25112,N_25371);
and UO_1144 (O_1144,N_27487,N_27255);
nor UO_1145 (O_1145,N_26311,N_25833);
xnor UO_1146 (O_1146,N_29013,N_25549);
xor UO_1147 (O_1147,N_25791,N_28276);
nand UO_1148 (O_1148,N_26875,N_28734);
or UO_1149 (O_1149,N_28870,N_25059);
and UO_1150 (O_1150,N_28091,N_27169);
xor UO_1151 (O_1151,N_26108,N_28372);
or UO_1152 (O_1152,N_28335,N_27276);
nor UO_1153 (O_1153,N_29836,N_28894);
and UO_1154 (O_1154,N_29296,N_29460);
xnor UO_1155 (O_1155,N_25143,N_26646);
xnor UO_1156 (O_1156,N_28100,N_28875);
xnor UO_1157 (O_1157,N_27694,N_27145);
xor UO_1158 (O_1158,N_25957,N_25903);
nor UO_1159 (O_1159,N_29957,N_28783);
nor UO_1160 (O_1160,N_28400,N_27863);
xor UO_1161 (O_1161,N_27017,N_25425);
or UO_1162 (O_1162,N_27265,N_27458);
and UO_1163 (O_1163,N_25050,N_29187);
nand UO_1164 (O_1164,N_27938,N_26056);
nor UO_1165 (O_1165,N_25170,N_25757);
or UO_1166 (O_1166,N_26969,N_26531);
or UO_1167 (O_1167,N_25266,N_27485);
nor UO_1168 (O_1168,N_29903,N_25746);
nor UO_1169 (O_1169,N_27851,N_29581);
and UO_1170 (O_1170,N_25819,N_27795);
and UO_1171 (O_1171,N_29065,N_29563);
or UO_1172 (O_1172,N_29126,N_27875);
nand UO_1173 (O_1173,N_26011,N_29770);
or UO_1174 (O_1174,N_29202,N_29035);
nand UO_1175 (O_1175,N_26955,N_29410);
nand UO_1176 (O_1176,N_25433,N_28904);
or UO_1177 (O_1177,N_27881,N_26281);
nand UO_1178 (O_1178,N_26532,N_26653);
xor UO_1179 (O_1179,N_29324,N_27129);
nand UO_1180 (O_1180,N_27338,N_26342);
xnor UO_1181 (O_1181,N_28521,N_26742);
or UO_1182 (O_1182,N_28508,N_29194);
and UO_1183 (O_1183,N_25136,N_29225);
or UO_1184 (O_1184,N_25918,N_26705);
xnor UO_1185 (O_1185,N_29497,N_29611);
xor UO_1186 (O_1186,N_27923,N_28240);
nor UO_1187 (O_1187,N_29733,N_28612);
or UO_1188 (O_1188,N_28212,N_25774);
or UO_1189 (O_1189,N_25300,N_26765);
xnor UO_1190 (O_1190,N_28142,N_29054);
or UO_1191 (O_1191,N_25199,N_25977);
nand UO_1192 (O_1192,N_28795,N_26951);
and UO_1193 (O_1193,N_27568,N_26026);
or UO_1194 (O_1194,N_26751,N_27046);
nor UO_1195 (O_1195,N_29539,N_28214);
or UO_1196 (O_1196,N_28446,N_27034);
xor UO_1197 (O_1197,N_26549,N_28697);
xor UO_1198 (O_1198,N_25127,N_25256);
and UO_1199 (O_1199,N_29947,N_28716);
and UO_1200 (O_1200,N_27172,N_27188);
nor UO_1201 (O_1201,N_28594,N_28556);
xor UO_1202 (O_1202,N_26899,N_26936);
nand UO_1203 (O_1203,N_29102,N_25061);
xor UO_1204 (O_1204,N_29526,N_26685);
nand UO_1205 (O_1205,N_25682,N_25437);
or UO_1206 (O_1206,N_28820,N_27372);
nor UO_1207 (O_1207,N_29542,N_29038);
and UO_1208 (O_1208,N_29697,N_29703);
nor UO_1209 (O_1209,N_28800,N_27835);
and UO_1210 (O_1210,N_29502,N_29932);
and UO_1211 (O_1211,N_26736,N_26003);
xor UO_1212 (O_1212,N_29782,N_25737);
and UO_1213 (O_1213,N_28420,N_29245);
and UO_1214 (O_1214,N_27708,N_29644);
and UO_1215 (O_1215,N_25092,N_25793);
nor UO_1216 (O_1216,N_27278,N_29795);
or UO_1217 (O_1217,N_26701,N_26767);
nor UO_1218 (O_1218,N_27234,N_29477);
nor UO_1219 (O_1219,N_26940,N_28024);
nor UO_1220 (O_1220,N_29799,N_26188);
or UO_1221 (O_1221,N_26762,N_26221);
nor UO_1222 (O_1222,N_29583,N_29541);
or UO_1223 (O_1223,N_26805,N_26495);
or UO_1224 (O_1224,N_29822,N_28364);
and UO_1225 (O_1225,N_29057,N_29509);
nor UO_1226 (O_1226,N_25641,N_28371);
nand UO_1227 (O_1227,N_28970,N_25930);
xnor UO_1228 (O_1228,N_29835,N_27457);
xnor UO_1229 (O_1229,N_28569,N_26537);
nor UO_1230 (O_1230,N_28185,N_26626);
nand UO_1231 (O_1231,N_28028,N_25068);
nor UO_1232 (O_1232,N_25751,N_29327);
nand UO_1233 (O_1233,N_26045,N_29168);
xor UO_1234 (O_1234,N_26150,N_28336);
and UO_1235 (O_1235,N_28051,N_27380);
xnor UO_1236 (O_1236,N_26127,N_26921);
xnor UO_1237 (O_1237,N_26677,N_25900);
or UO_1238 (O_1238,N_28324,N_28230);
and UO_1239 (O_1239,N_26942,N_26271);
or UO_1240 (O_1240,N_26297,N_27514);
or UO_1241 (O_1241,N_26137,N_25415);
and UO_1242 (O_1242,N_26654,N_29061);
and UO_1243 (O_1243,N_25058,N_27422);
and UO_1244 (O_1244,N_29125,N_26022);
nand UO_1245 (O_1245,N_27430,N_28412);
xnor UO_1246 (O_1246,N_25907,N_27065);
or UO_1247 (O_1247,N_27639,N_25248);
and UO_1248 (O_1248,N_28706,N_28640);
nor UO_1249 (O_1249,N_28693,N_28350);
and UO_1250 (O_1250,N_28126,N_27054);
or UO_1251 (O_1251,N_28360,N_28498);
and UO_1252 (O_1252,N_27303,N_27847);
xor UO_1253 (O_1253,N_28515,N_29641);
nand UO_1254 (O_1254,N_27852,N_25752);
nor UO_1255 (O_1255,N_29550,N_26573);
and UO_1256 (O_1256,N_26606,N_28916);
nor UO_1257 (O_1257,N_25125,N_25327);
and UO_1258 (O_1258,N_29612,N_25268);
nor UO_1259 (O_1259,N_25665,N_29930);
or UO_1260 (O_1260,N_27988,N_27045);
xor UO_1261 (O_1261,N_29449,N_28352);
and UO_1262 (O_1262,N_28723,N_25451);
xnor UO_1263 (O_1263,N_29833,N_28790);
xor UO_1264 (O_1264,N_27717,N_29853);
nor UO_1265 (O_1265,N_25347,N_28379);
or UO_1266 (O_1266,N_27728,N_29750);
nor UO_1267 (O_1267,N_27209,N_26321);
nand UO_1268 (O_1268,N_27738,N_28676);
nand UO_1269 (O_1269,N_29098,N_26074);
or UO_1270 (O_1270,N_27441,N_28618);
nor UO_1271 (O_1271,N_26615,N_27501);
or UO_1272 (O_1272,N_28792,N_25813);
nor UO_1273 (O_1273,N_29538,N_28699);
nor UO_1274 (O_1274,N_29714,N_26201);
nand UO_1275 (O_1275,N_27769,N_27026);
nor UO_1276 (O_1276,N_27090,N_27392);
nor UO_1277 (O_1277,N_28921,N_25365);
nor UO_1278 (O_1278,N_28058,N_27199);
or UO_1279 (O_1279,N_25214,N_26493);
nand UO_1280 (O_1280,N_27971,N_29674);
xnor UO_1281 (O_1281,N_28586,N_29636);
nand UO_1282 (O_1282,N_28080,N_29723);
or UO_1283 (O_1283,N_28822,N_29162);
nand UO_1284 (O_1284,N_28405,N_25412);
xnor UO_1285 (O_1285,N_25994,N_29154);
or UO_1286 (O_1286,N_29486,N_28471);
xnor UO_1287 (O_1287,N_27214,N_29390);
nand UO_1288 (O_1288,N_25985,N_28724);
nand UO_1289 (O_1289,N_28644,N_25309);
and UO_1290 (O_1290,N_29684,N_27118);
nand UO_1291 (O_1291,N_26896,N_27607);
and UO_1292 (O_1292,N_29273,N_25065);
or UO_1293 (O_1293,N_27283,N_27105);
nand UO_1294 (O_1294,N_25710,N_27411);
or UO_1295 (O_1295,N_27843,N_28056);
nor UO_1296 (O_1296,N_29972,N_29522);
xor UO_1297 (O_1297,N_25353,N_26236);
xnor UO_1298 (O_1298,N_28932,N_25261);
nand UO_1299 (O_1299,N_27709,N_28492);
xor UO_1300 (O_1300,N_28234,N_29433);
nor UO_1301 (O_1301,N_25719,N_27443);
nand UO_1302 (O_1302,N_26632,N_28137);
or UO_1303 (O_1303,N_26885,N_27798);
and UO_1304 (O_1304,N_27692,N_28465);
or UO_1305 (O_1305,N_27442,N_26917);
nor UO_1306 (O_1306,N_25434,N_26891);
xnor UO_1307 (O_1307,N_26700,N_28217);
or UO_1308 (O_1308,N_26338,N_25797);
nand UO_1309 (O_1309,N_28241,N_25949);
xnor UO_1310 (O_1310,N_27941,N_28398);
nor UO_1311 (O_1311,N_28539,N_26373);
xor UO_1312 (O_1312,N_27192,N_25733);
nor UO_1313 (O_1313,N_28847,N_27883);
and UO_1314 (O_1314,N_26708,N_25736);
or UO_1315 (O_1315,N_27061,N_28989);
nor UO_1316 (O_1316,N_26979,N_27075);
xnor UO_1317 (O_1317,N_29354,N_26726);
xnor UO_1318 (O_1318,N_25887,N_29909);
xnor UO_1319 (O_1319,N_25738,N_25627);
and UO_1320 (O_1320,N_27648,N_29226);
nor UO_1321 (O_1321,N_29421,N_25585);
xor UO_1322 (O_1322,N_25892,N_29504);
nand UO_1323 (O_1323,N_25454,N_29735);
and UO_1324 (O_1324,N_26434,N_28888);
nand UO_1325 (O_1325,N_29274,N_29594);
nor UO_1326 (O_1326,N_29896,N_28952);
nor UO_1327 (O_1327,N_25009,N_29099);
or UO_1328 (O_1328,N_25258,N_28435);
or UO_1329 (O_1329,N_25823,N_25103);
nand UO_1330 (O_1330,N_25215,N_28500);
or UO_1331 (O_1331,N_28667,N_26621);
nand UO_1332 (O_1332,N_25012,N_25105);
and UO_1333 (O_1333,N_28748,N_27153);
nand UO_1334 (O_1334,N_26191,N_27900);
xnor UO_1335 (O_1335,N_27924,N_27609);
xnor UO_1336 (O_1336,N_29131,N_25296);
nor UO_1337 (O_1337,N_26972,N_25402);
nand UO_1338 (O_1338,N_25859,N_25828);
nor UO_1339 (O_1339,N_29892,N_25370);
and UO_1340 (O_1340,N_27415,N_25637);
or UO_1341 (O_1341,N_28600,N_25537);
or UO_1342 (O_1342,N_25427,N_29934);
or UO_1343 (O_1343,N_27542,N_28468);
and UO_1344 (O_1344,N_29367,N_28188);
nor UO_1345 (O_1345,N_28033,N_26341);
or UO_1346 (O_1346,N_28395,N_25098);
nand UO_1347 (O_1347,N_29997,N_26106);
and UO_1348 (O_1348,N_28833,N_27603);
xor UO_1349 (O_1349,N_27596,N_27326);
nor UO_1350 (O_1350,N_28867,N_25101);
and UO_1351 (O_1351,N_26372,N_27002);
nand UO_1352 (O_1352,N_27435,N_28622);
and UO_1353 (O_1353,N_25584,N_25814);
nor UO_1354 (O_1354,N_25015,N_27630);
nor UO_1355 (O_1355,N_25986,N_27968);
nor UO_1356 (O_1356,N_28590,N_25535);
xor UO_1357 (O_1357,N_29049,N_27346);
xor UO_1358 (O_1358,N_29428,N_29214);
xnor UO_1359 (O_1359,N_29518,N_26207);
or UO_1360 (O_1360,N_25247,N_25329);
nand UO_1361 (O_1361,N_29292,N_27972);
xor UO_1362 (O_1362,N_25314,N_29759);
nand UO_1363 (O_1363,N_25609,N_28455);
and UO_1364 (O_1364,N_27827,N_29328);
nor UO_1365 (O_1365,N_28484,N_27808);
and UO_1366 (O_1366,N_29007,N_28155);
nor UO_1367 (O_1367,N_26017,N_27273);
and UO_1368 (O_1368,N_25203,N_27180);
xnor UO_1369 (O_1369,N_29748,N_27589);
xor UO_1370 (O_1370,N_27894,N_25794);
or UO_1371 (O_1371,N_28444,N_26640);
nand UO_1372 (O_1372,N_25408,N_27869);
and UO_1373 (O_1373,N_26435,N_29552);
nor UO_1374 (O_1374,N_26414,N_26208);
nand UO_1375 (O_1375,N_25995,N_27174);
nand UO_1376 (O_1376,N_28042,N_25491);
xor UO_1377 (O_1377,N_28532,N_26472);
nand UO_1378 (O_1378,N_27427,N_27235);
and UO_1379 (O_1379,N_29492,N_27106);
nor UO_1380 (O_1380,N_29227,N_26284);
or UO_1381 (O_1381,N_27056,N_25783);
and UO_1382 (O_1382,N_26733,N_27634);
xor UO_1383 (O_1383,N_28884,N_27716);
nand UO_1384 (O_1384,N_28740,N_28601);
xor UO_1385 (O_1385,N_25264,N_29097);
and UO_1386 (O_1386,N_29572,N_27253);
nor UO_1387 (O_1387,N_27764,N_28391);
or UO_1388 (O_1388,N_27407,N_29963);
and UO_1389 (O_1389,N_27802,N_27433);
nand UO_1390 (O_1390,N_28564,N_27926);
nand UO_1391 (O_1391,N_26943,N_25312);
or UO_1392 (O_1392,N_27651,N_28960);
nand UO_1393 (O_1393,N_25999,N_28764);
or UO_1394 (O_1394,N_27097,N_27250);
xnor UO_1395 (O_1395,N_28975,N_25085);
nor UO_1396 (O_1396,N_25925,N_26887);
nor UO_1397 (O_1397,N_29908,N_27807);
xnor UO_1398 (O_1398,N_25192,N_27119);
or UO_1399 (O_1399,N_28809,N_25147);
or UO_1400 (O_1400,N_28006,N_25714);
or UO_1401 (O_1401,N_27328,N_26198);
and UO_1402 (O_1402,N_28215,N_27226);
nand UO_1403 (O_1403,N_28369,N_27404);
nor UO_1404 (O_1404,N_29579,N_28976);
nand UO_1405 (O_1405,N_28512,N_28199);
nor UO_1406 (O_1406,N_29650,N_28977);
xnor UO_1407 (O_1407,N_26343,N_27543);
or UO_1408 (O_1408,N_28449,N_25904);
xor UO_1409 (O_1409,N_27167,N_25739);
nand UO_1410 (O_1410,N_29924,N_29747);
or UO_1411 (O_1411,N_26497,N_27965);
or UO_1412 (O_1412,N_25213,N_25381);
or UO_1413 (O_1413,N_26412,N_25638);
nand UO_1414 (O_1414,N_25102,N_25508);
nor UO_1415 (O_1415,N_27601,N_26813);
and UO_1416 (O_1416,N_28841,N_28523);
or UO_1417 (O_1417,N_25800,N_26332);
nor UO_1418 (O_1418,N_28103,N_27892);
and UO_1419 (O_1419,N_27638,N_28362);
nand UO_1420 (O_1420,N_25756,N_25845);
nor UO_1421 (O_1421,N_26117,N_29732);
nor UO_1422 (O_1422,N_28728,N_28187);
nor UO_1423 (O_1423,N_25301,N_25482);
nand UO_1424 (O_1424,N_28929,N_28825);
xnor UO_1425 (O_1425,N_28980,N_28679);
nand UO_1426 (O_1426,N_27563,N_29543);
or UO_1427 (O_1427,N_28950,N_26423);
nor UO_1428 (O_1428,N_29016,N_28293);
xnor UO_1429 (O_1429,N_29727,N_27029);
nor UO_1430 (O_1430,N_29865,N_27003);
and UO_1431 (O_1431,N_28265,N_26826);
xnor UO_1432 (O_1432,N_29668,N_27331);
xor UO_1433 (O_1433,N_29756,N_28743);
or UO_1434 (O_1434,N_25878,N_28134);
nand UO_1435 (O_1435,N_27133,N_27373);
xor UO_1436 (O_1436,N_26382,N_27577);
nand UO_1437 (O_1437,N_26563,N_25409);
xor UO_1438 (O_1438,N_29235,N_26471);
nor UO_1439 (O_1439,N_27830,N_26243);
xnor UO_1440 (O_1440,N_28012,N_27908);
nor UO_1441 (O_1441,N_27086,N_26627);
nand UO_1442 (O_1442,N_26795,N_26526);
nand UO_1443 (O_1443,N_28008,N_29775);
nor UO_1444 (O_1444,N_29844,N_27059);
nor UO_1445 (O_1445,N_29109,N_27073);
nor UO_1446 (O_1446,N_28609,N_29989);
xor UO_1447 (O_1447,N_29870,N_26719);
and UO_1448 (O_1448,N_26947,N_26558);
or UO_1449 (O_1449,N_25942,N_29886);
or UO_1450 (O_1450,N_29375,N_26402);
xor UO_1451 (O_1451,N_25407,N_25148);
or UO_1452 (O_1452,N_27792,N_29443);
and UO_1453 (O_1453,N_26710,N_25848);
nor UO_1454 (O_1454,N_29568,N_27149);
nand UO_1455 (O_1455,N_26630,N_25459);
xor UO_1456 (O_1456,N_29232,N_25550);
and UO_1457 (O_1457,N_28715,N_29914);
nand UO_1458 (O_1458,N_26635,N_26839);
xor UO_1459 (O_1459,N_26218,N_27942);
xnor UO_1460 (O_1460,N_25531,N_26440);
and UO_1461 (O_1461,N_28525,N_26631);
and UO_1462 (O_1462,N_29236,N_25720);
nor UO_1463 (O_1463,N_27178,N_26286);
and UO_1464 (O_1464,N_29501,N_29730);
nand UO_1465 (O_1465,N_29037,N_28629);
or UO_1466 (O_1466,N_29812,N_26679);
or UO_1467 (O_1467,N_29383,N_26484);
xor UO_1468 (O_1468,N_25836,N_25605);
xor UO_1469 (O_1469,N_26859,N_29164);
nor UO_1470 (O_1470,N_28110,N_28113);
or UO_1471 (O_1471,N_25948,N_28785);
or UO_1472 (O_1472,N_25392,N_26156);
or UO_1473 (O_1473,N_29536,N_27267);
or UO_1474 (O_1474,N_27813,N_29894);
xnor UO_1475 (O_1475,N_25937,N_26439);
nand UO_1476 (O_1476,N_26256,N_25299);
nor UO_1477 (O_1477,N_27724,N_25824);
nand UO_1478 (O_1478,N_29603,N_26283);
xnor UO_1479 (O_1479,N_27898,N_26660);
nand UO_1480 (O_1480,N_27274,N_29990);
xor UO_1481 (O_1481,N_27205,N_26399);
nand UO_1482 (O_1482,N_27297,N_28367);
or UO_1483 (O_1483,N_25843,N_25851);
nor UO_1484 (O_1484,N_25462,N_27530);
or UO_1485 (O_1485,N_28101,N_29092);
nand UO_1486 (O_1486,N_28541,N_29915);
and UO_1487 (O_1487,N_29602,N_26292);
and UO_1488 (O_1488,N_25162,N_28169);
and UO_1489 (O_1489,N_29216,N_27671);
xor UO_1490 (O_1490,N_28544,N_26911);
and UO_1491 (O_1491,N_27797,N_25877);
nand UO_1492 (O_1492,N_29242,N_27282);
xor UO_1493 (O_1493,N_29488,N_28231);
xor UO_1494 (O_1494,N_28053,N_26609);
and UO_1495 (O_1495,N_29051,N_25423);
xor UO_1496 (O_1496,N_27176,N_25883);
and UO_1497 (O_1497,N_28050,N_28671);
xnor UO_1498 (O_1498,N_29193,N_25424);
nor UO_1499 (O_1499,N_29877,N_29499);
nor UO_1500 (O_1500,N_28380,N_28488);
or UO_1501 (O_1501,N_25917,N_26482);
xor UO_1502 (O_1502,N_25831,N_28674);
xnor UO_1503 (O_1503,N_25826,N_29254);
nand UO_1504 (O_1504,N_27281,N_25632);
xor UO_1505 (O_1505,N_29804,N_27999);
and UO_1506 (O_1506,N_27664,N_28592);
xnor UO_1507 (O_1507,N_26797,N_27656);
nand UO_1508 (O_1508,N_27294,N_29884);
nand UO_1509 (O_1509,N_27641,N_29005);
or UO_1510 (O_1510,N_29855,N_27917);
or UO_1511 (O_1511,N_25515,N_27268);
or UO_1512 (O_1512,N_26523,N_25897);
nand UO_1513 (O_1513,N_26047,N_26441);
xnor UO_1514 (O_1514,N_28973,N_29649);
or UO_1515 (O_1515,N_26295,N_25345);
nand UO_1516 (O_1516,N_25380,N_26964);
nor UO_1517 (O_1517,N_25150,N_29628);
or UO_1518 (O_1518,N_26718,N_26354);
nand UO_1519 (O_1519,N_26503,N_29103);
nand UO_1520 (O_1520,N_29856,N_25712);
xnor UO_1521 (O_1521,N_26015,N_26599);
nand UO_1522 (O_1522,N_28813,N_25952);
nor UO_1523 (O_1523,N_25003,N_27413);
xor UO_1524 (O_1524,N_29623,N_29891);
nor UO_1525 (O_1525,N_25898,N_29762);
or UO_1526 (O_1526,N_26601,N_25908);
nand UO_1527 (O_1527,N_27841,N_28401);
xnor UO_1528 (O_1528,N_28167,N_26009);
or UO_1529 (O_1529,N_26697,N_29797);
nand UO_1530 (O_1530,N_25285,N_28741);
or UO_1531 (O_1531,N_27136,N_25577);
xnor UO_1532 (O_1532,N_25303,N_27879);
nor UO_1533 (O_1533,N_29241,N_25825);
and UO_1534 (O_1534,N_26054,N_28910);
nor UO_1535 (O_1535,N_27850,N_26211);
nand UO_1536 (O_1536,N_26258,N_28207);
nand UO_1537 (O_1537,N_29337,N_29135);
nand UO_1538 (O_1538,N_25768,N_27410);
and UO_1539 (O_1539,N_26216,N_28105);
nor UO_1540 (O_1540,N_25305,N_26259);
and UO_1541 (O_1541,N_27377,N_25018);
xor UO_1542 (O_1542,N_28147,N_27355);
nor UO_1543 (O_1543,N_28591,N_27914);
nor UO_1544 (O_1544,N_28442,N_28639);
or UO_1545 (O_1545,N_26033,N_29935);
nand UO_1546 (O_1546,N_27450,N_29489);
nor UO_1547 (O_1547,N_25590,N_25895);
xnor UO_1548 (O_1548,N_29913,N_27637);
nand UO_1549 (O_1549,N_28576,N_29933);
or UO_1550 (O_1550,N_25260,N_27640);
nand UO_1551 (O_1551,N_28470,N_29888);
or UO_1552 (O_1552,N_27535,N_29883);
and UO_1553 (O_1553,N_29901,N_26824);
xor UO_1554 (O_1554,N_28763,N_28366);
nand UO_1555 (O_1555,N_27130,N_26090);
nand UO_1556 (O_1556,N_28026,N_26465);
and UO_1557 (O_1557,N_27871,N_28396);
or UO_1558 (O_1558,N_28323,N_25131);
and UO_1559 (O_1559,N_26253,N_27201);
nor UO_1560 (O_1560,N_25311,N_29191);
nor UO_1561 (O_1561,N_25913,N_27681);
nor UO_1562 (O_1562,N_26533,N_29158);
nor UO_1563 (O_1563,N_26929,N_25668);
xnor UO_1564 (O_1564,N_28149,N_29709);
nand UO_1565 (O_1565,N_27064,N_29381);
nand UO_1566 (O_1566,N_29731,N_25233);
nor UO_1567 (O_1567,N_26057,N_26025);
and UO_1568 (O_1568,N_29873,N_26811);
or UO_1569 (O_1569,N_27722,N_28459);
and UO_1570 (O_1570,N_26183,N_25690);
and UO_1571 (O_1571,N_26141,N_27079);
xor UO_1572 (O_1572,N_25817,N_26046);
and UO_1573 (O_1573,N_27011,N_28620);
nor UO_1574 (O_1574,N_25465,N_25656);
nor UO_1575 (O_1575,N_25064,N_29066);
nand UO_1576 (O_1576,N_26388,N_26369);
nor UO_1577 (O_1577,N_27368,N_26251);
nand UO_1578 (O_1578,N_26429,N_29939);
xor UO_1579 (O_1579,N_29207,N_26939);
and UO_1580 (O_1580,N_25017,N_27783);
nand UO_1581 (O_1581,N_26699,N_26669);
and UO_1582 (O_1582,N_25306,N_27901);
nor UO_1583 (O_1583,N_25767,N_28311);
nor UO_1584 (O_1584,N_26643,N_29490);
or UO_1585 (O_1585,N_28857,N_27815);
nor UO_1586 (O_1586,N_28572,N_27104);
and UO_1587 (O_1587,N_25571,N_29587);
and UO_1588 (O_1588,N_25861,N_29646);
xnor UO_1589 (O_1589,N_25280,N_25765);
nand UO_1590 (O_1590,N_25889,N_25458);
nand UO_1591 (O_1591,N_27241,N_28584);
nor UO_1592 (O_1592,N_27233,N_28424);
nor UO_1593 (O_1593,N_26628,N_29247);
or UO_1594 (O_1594,N_28014,N_29401);
nor UO_1595 (O_1595,N_29152,N_27707);
and UO_1596 (O_1596,N_27425,N_29692);
nor UO_1597 (O_1597,N_26863,N_25205);
nor UO_1598 (O_1598,N_27344,N_28289);
nor UO_1599 (O_1599,N_28727,N_28797);
nor UO_1600 (O_1600,N_26084,N_26902);
and UO_1601 (O_1601,N_28533,N_27217);
xnor UO_1602 (O_1602,N_29864,N_28044);
xnor UO_1603 (O_1603,N_27896,N_28547);
nand UO_1604 (O_1604,N_28177,N_29082);
or UO_1605 (O_1605,N_26140,N_29132);
nand UO_1606 (O_1606,N_25468,N_28440);
or UO_1607 (O_1607,N_25337,N_29372);
xor UO_1608 (O_1608,N_26391,N_25560);
nor UO_1609 (O_1609,N_29106,N_25262);
nand UO_1610 (O_1610,N_27703,N_28415);
xor UO_1611 (O_1611,N_26125,N_25616);
or UO_1612 (O_1612,N_25809,N_29397);
nand UO_1613 (O_1613,N_26189,N_27245);
nand UO_1614 (O_1614,N_29566,N_28901);
or UO_1615 (O_1615,N_29900,N_26706);
xor UO_1616 (O_1616,N_28582,N_26998);
nand UO_1617 (O_1617,N_25377,N_26505);
xnor UO_1618 (O_1618,N_25124,N_29345);
nand UO_1619 (O_1619,N_28312,N_27470);
and UO_1620 (O_1620,N_28281,N_29028);
xor UO_1621 (O_1621,N_29720,N_27718);
nor UO_1622 (O_1622,N_25400,N_28130);
or UO_1623 (O_1623,N_25664,N_29874);
nand UO_1624 (O_1624,N_27997,N_27207);
xor UO_1625 (O_1625,N_29281,N_25490);
nand UO_1626 (O_1626,N_26486,N_25934);
nand UO_1627 (O_1627,N_26238,N_27336);
nand UO_1628 (O_1628,N_28685,N_29866);
nand UO_1629 (O_1629,N_25518,N_27432);
and UO_1630 (O_1630,N_27445,N_29205);
or UO_1631 (O_1631,N_28107,N_27371);
and UO_1632 (O_1632,N_26894,N_27375);
xnor UO_1633 (O_1633,N_25046,N_25479);
and UO_1634 (O_1634,N_27498,N_29180);
xnor UO_1635 (O_1635,N_26346,N_25856);
nand UO_1636 (O_1636,N_27675,N_26778);
or UO_1637 (O_1637,N_26415,N_26395);
or UO_1638 (O_1638,N_29334,N_28093);
or UO_1639 (O_1639,N_29361,N_28930);
and UO_1640 (O_1640,N_29713,N_25087);
xnor UO_1641 (O_1641,N_28780,N_26608);
nor UO_1642 (O_1642,N_26310,N_27103);
xor UO_1643 (O_1643,N_28838,N_26312);
xor UO_1644 (O_1644,N_25528,N_25723);
and UO_1645 (O_1645,N_28557,N_27177);
or UO_1646 (O_1646,N_27491,N_25095);
or UO_1647 (O_1647,N_28709,N_25081);
nor UO_1648 (O_1648,N_27040,N_29359);
nor UO_1649 (O_1649,N_27448,N_29413);
nand UO_1650 (O_1650,N_26711,N_29435);
nand UO_1651 (O_1651,N_26162,N_27574);
xnor UO_1652 (O_1652,N_29523,N_29269);
xor UO_1653 (O_1653,N_28209,N_26968);
xnor UO_1654 (O_1654,N_27893,N_25128);
nor UO_1655 (O_1655,N_27455,N_26835);
and UO_1656 (O_1656,N_27812,N_28493);
or UO_1657 (O_1657,N_27258,N_29331);
xnor UO_1658 (O_1658,N_26363,N_29058);
xnor UO_1659 (O_1659,N_27538,N_26547);
xnor UO_1660 (O_1660,N_28721,N_26561);
nor UO_1661 (O_1661,N_28034,N_26502);
xor UO_1662 (O_1662,N_25525,N_26575);
xor UO_1663 (O_1663,N_26833,N_28375);
xor UO_1664 (O_1664,N_29769,N_29201);
or UO_1665 (O_1665,N_28119,N_25031);
and UO_1666 (O_1666,N_29971,N_29802);
and UO_1667 (O_1667,N_28695,N_27958);
nand UO_1668 (O_1668,N_29887,N_27483);
and UO_1669 (O_1669,N_27206,N_27212);
nor UO_1670 (O_1670,N_25600,N_29842);
or UO_1671 (O_1671,N_25228,N_28786);
nand UO_1672 (O_1672,N_27481,N_27557);
xor UO_1673 (O_1673,N_25139,N_26769);
and UO_1674 (O_1674,N_25922,N_29319);
or UO_1675 (O_1675,N_27966,N_26362);
and UO_1676 (O_1676,N_28736,N_29487);
nor UO_1677 (O_1677,N_25236,N_27643);
or UO_1678 (O_1678,N_28816,N_26212);
nand UO_1679 (O_1679,N_26171,N_26454);
xnor UO_1680 (O_1680,N_29182,N_28473);
xor UO_1681 (O_1681,N_28522,N_26872);
nor UO_1682 (O_1682,N_25388,N_26394);
nor UO_1683 (O_1683,N_29905,N_26808);
xnor UO_1684 (O_1684,N_25838,N_28220);
nor UO_1685 (O_1685,N_26756,N_29904);
nor UO_1686 (O_1686,N_27023,N_29210);
xnor UO_1687 (O_1687,N_27164,N_26600);
nor UO_1688 (O_1688,N_27302,N_28964);
nand UO_1689 (O_1689,N_28643,N_27418);
nor UO_1690 (O_1690,N_26636,N_26850);
nor UO_1691 (O_1691,N_25580,N_28070);
nand UO_1692 (O_1692,N_27271,N_27279);
nor UO_1693 (O_1693,N_28253,N_28285);
nand UO_1694 (O_1694,N_26219,N_26215);
or UO_1695 (O_1695,N_27789,N_27395);
and UO_1696 (O_1696,N_26738,N_25631);
xnor UO_1697 (O_1697,N_29791,N_25701);
nor UO_1698 (O_1698,N_27347,N_25368);
or UO_1699 (O_1699,N_25313,N_27511);
or UO_1700 (O_1700,N_25960,N_25161);
nor UO_1701 (O_1701,N_26907,N_26665);
nand UO_1702 (O_1702,N_27821,N_27053);
and UO_1703 (O_1703,N_28689,N_28889);
xnor UO_1704 (O_1704,N_29941,N_29128);
nand UO_1705 (O_1705,N_29778,N_29753);
nand UO_1706 (O_1706,N_26556,N_26793);
or UO_1707 (O_1707,N_27655,N_26390);
and UO_1708 (O_1708,N_26919,N_29392);
nand UO_1709 (O_1709,N_26591,N_28104);
and UO_1710 (O_1710,N_26786,N_26617);
and UO_1711 (O_1711,N_26604,N_27398);
and UO_1712 (O_1712,N_29945,N_27519);
nor UO_1713 (O_1713,N_26158,N_26345);
nor UO_1714 (O_1714,N_29617,N_26016);
nor UO_1715 (O_1715,N_25633,N_29371);
and UO_1716 (O_1716,N_27242,N_25477);
nand UO_1717 (O_1717,N_26309,N_25448);
nor UO_1718 (O_1718,N_29084,N_28343);
xnor UO_1719 (O_1719,N_28953,N_25726);
nand UO_1720 (O_1720,N_29656,N_28645);
nand UO_1721 (O_1721,N_28127,N_25830);
xnor UO_1722 (O_1722,N_28905,N_28292);
xor UO_1723 (O_1723,N_28703,N_28974);
nand UO_1724 (O_1724,N_26405,N_25689);
nor UO_1725 (O_1725,N_27447,N_27050);
xor UO_1726 (O_1726,N_28361,N_29370);
and UO_1727 (O_1727,N_27592,N_26334);
nor UO_1728 (O_1728,N_27913,N_26460);
nor UO_1729 (O_1729,N_27933,N_29527);
and UO_1730 (O_1730,N_27727,N_29950);
nand UO_1731 (O_1731,N_26645,N_25962);
xor UO_1732 (O_1732,N_29108,N_25083);
nor UO_1733 (O_1733,N_25363,N_29387);
nand UO_1734 (O_1734,N_25953,N_26764);
and UO_1735 (O_1735,N_27740,N_28273);
nor UO_1736 (O_1736,N_29751,N_28021);
nor UO_1737 (O_1737,N_27001,N_25841);
or UO_1738 (O_1738,N_28338,N_27423);
or UO_1739 (O_1739,N_27525,N_29114);
or UO_1740 (O_1740,N_29151,N_27110);
or UO_1741 (O_1741,N_26570,N_27337);
xor UO_1742 (O_1742,N_29916,N_25618);
nor UO_1743 (O_1743,N_29728,N_25728);
nor UO_1744 (O_1744,N_28291,N_25507);
nor UO_1745 (O_1745,N_25013,N_26021);
and UO_1746 (O_1746,N_27354,N_26432);
or UO_1747 (O_1747,N_29648,N_29846);
nor UO_1748 (O_1748,N_29810,N_26222);
or UO_1749 (O_1749,N_28018,N_26371);
nand UO_1750 (O_1750,N_25242,N_26270);
and UO_1751 (O_1751,N_26061,N_25519);
xor UO_1752 (O_1752,N_26516,N_25185);
nand UO_1753 (O_1753,N_27266,N_28934);
and UO_1754 (O_1754,N_25788,N_28099);
nand UO_1755 (O_1755,N_26425,N_27569);
nor UO_1756 (O_1756,N_29571,N_29821);
and UO_1757 (O_1757,N_26351,N_26473);
xnor UO_1758 (O_1758,N_26923,N_29300);
nor UO_1759 (O_1759,N_25920,N_26030);
nand UO_1760 (O_1760,N_26190,N_28982);
or UO_1761 (O_1761,N_25863,N_28452);
xnor UO_1762 (O_1762,N_28939,N_26217);
or UO_1763 (O_1763,N_28475,N_25156);
nor UO_1764 (O_1764,N_26375,N_27523);
and UO_1765 (O_1765,N_29558,N_26717);
and UO_1766 (O_1766,N_29388,N_26883);
and UO_1767 (O_1767,N_27550,N_29613);
nand UO_1768 (O_1768,N_26214,N_27263);
nand UO_1769 (O_1769,N_26739,N_29320);
nand UO_1770 (O_1770,N_28462,N_27154);
or UO_1771 (O_1771,N_27878,N_25623);
or UO_1772 (O_1772,N_26876,N_27363);
nand UO_1773 (O_1773,N_27360,N_28682);
or UO_1774 (O_1774,N_28236,N_27644);
nor UO_1775 (O_1775,N_28036,N_27247);
xor UO_1776 (O_1776,N_25405,N_25976);
xnor UO_1777 (O_1777,N_29902,N_29417);
xor UO_1778 (O_1778,N_28947,N_29369);
nor UO_1779 (O_1779,N_28141,N_28726);
and UO_1780 (O_1780,N_26456,N_29183);
xnor UO_1781 (O_1781,N_27451,N_28002);
nand UO_1782 (O_1782,N_29570,N_29004);
nor UO_1783 (O_1783,N_27957,N_26729);
nor UO_1784 (O_1784,N_29294,N_28059);
xnor UO_1785 (O_1785,N_26255,N_29829);
or UO_1786 (O_1786,N_28108,N_28842);
and UO_1787 (O_1787,N_26323,N_26809);
nand UO_1788 (O_1788,N_28392,N_28758);
or UO_1789 (O_1789,N_27081,N_28020);
nor UO_1790 (O_1790,N_26818,N_27524);
nand UO_1791 (O_1791,N_29308,N_28935);
and UO_1792 (O_1792,N_26607,N_29806);
and UO_1793 (O_1793,N_28985,N_28698);
xnor UO_1794 (O_1794,N_26058,N_26464);
nor UO_1795 (O_1795,N_29575,N_25956);
and UO_1796 (O_1796,N_26038,N_27534);
nand UO_1797 (O_1797,N_28537,N_25504);
nor UO_1798 (O_1798,N_28195,N_29117);
xnor UO_1799 (O_1799,N_26393,N_28496);
or UO_1800 (O_1800,N_27475,N_25896);
and UO_1801 (O_1801,N_25293,N_29149);
or UO_1802 (O_1802,N_26407,N_27195);
and UO_1803 (O_1803,N_26143,N_26934);
and UO_1804 (O_1804,N_29034,N_26890);
and UO_1805 (O_1805,N_28464,N_29689);
nor UO_1806 (O_1806,N_29519,N_27662);
nand UO_1807 (O_1807,N_25762,N_27222);
nor UO_1808 (O_1808,N_29604,N_26417);
nand UO_1809 (O_1809,N_27872,N_29592);
and UO_1810 (O_1810,N_29868,N_25302);
nor UO_1811 (O_1811,N_25359,N_27190);
and UO_1812 (O_1812,N_26571,N_25970);
nand UO_1813 (O_1813,N_28428,N_26559);
nor UO_1814 (O_1814,N_27486,N_27905);
and UO_1815 (O_1815,N_25536,N_29056);
or UO_1816 (O_1816,N_29219,N_29794);
xor UO_1817 (O_1817,N_28102,N_25421);
and UO_1818 (O_1818,N_29531,N_29445);
nand UO_1819 (O_1819,N_27157,N_25651);
xnor UO_1820 (O_1820,N_28933,N_27471);
nand UO_1821 (O_1821,N_25983,N_26642);
and UO_1822 (O_1822,N_29695,N_29906);
or UO_1823 (O_1823,N_28570,N_29970);
or UO_1824 (O_1824,N_25530,N_29012);
and UO_1825 (O_1825,N_26895,N_27308);
and UO_1826 (O_1826,N_27063,N_27349);
or UO_1827 (O_1827,N_26927,N_27582);
xnor UO_1828 (O_1828,N_25172,N_25517);
and UO_1829 (O_1829,N_28226,N_25020);
nand UO_1830 (O_1830,N_26213,N_28479);
xor UO_1831 (O_1831,N_28184,N_27246);
or UO_1832 (O_1832,N_27173,N_26196);
xor UO_1833 (O_1833,N_27394,N_25045);
nor UO_1834 (O_1834,N_26483,N_26661);
or UO_1835 (O_1835,N_26846,N_27661);
nand UO_1836 (O_1836,N_28271,N_29136);
xor UO_1837 (O_1837,N_28122,N_28860);
and UO_1838 (O_1838,N_28399,N_29534);
nand UO_1839 (O_1839,N_27770,N_27632);
nand UO_1840 (O_1840,N_29740,N_27025);
nand UO_1841 (O_1841,N_25344,N_27341);
nor UO_1842 (O_1842,N_27374,N_27576);
and UO_1843 (O_1843,N_29642,N_29978);
nor UO_1844 (O_1844,N_25469,N_25445);
nand UO_1845 (O_1845,N_26051,N_25034);
or UO_1846 (O_1846,N_29513,N_26704);
or UO_1847 (O_1847,N_26229,N_27350);
or UO_1848 (O_1848,N_26521,N_29316);
nand UO_1849 (O_1849,N_29001,N_27137);
or UO_1850 (O_1850,N_28425,N_26121);
xor UO_1851 (O_1851,N_27992,N_29715);
nor UO_1852 (O_1852,N_28608,N_29506);
or UO_1853 (O_1853,N_27152,N_27561);
or UO_1854 (O_1854,N_26852,N_26664);
xor UO_1855 (O_1855,N_27052,N_29928);
nand UO_1856 (O_1856,N_28139,N_27597);
nor UO_1857 (O_1857,N_29465,N_25660);
or UO_1858 (O_1858,N_29755,N_28670);
xnor UO_1859 (O_1859,N_27262,N_28009);
xnor UO_1860 (O_1860,N_28823,N_28534);
nor UO_1861 (O_1861,N_27874,N_25399);
and UO_1862 (O_1862,N_27935,N_25592);
or UO_1863 (O_1863,N_29389,N_25687);
xnor UO_1864 (O_1864,N_29240,N_28251);
nor UO_1865 (O_1865,N_27822,N_28298);
xor UO_1866 (O_1866,N_26668,N_28154);
and UO_1867 (O_1867,N_28560,N_26590);
or UO_1868 (O_1868,N_26745,N_26884);
and UO_1869 (O_1869,N_25684,N_25936);
and UO_1870 (O_1870,N_25750,N_28098);
nand UO_1871 (O_1871,N_25027,N_29491);
or UO_1872 (O_1872,N_29318,N_26202);
and UO_1873 (O_1873,N_26974,N_29508);
or UO_1874 (O_1874,N_25675,N_29188);
xnor UO_1875 (O_1875,N_28663,N_29425);
or UO_1876 (O_1876,N_27868,N_29033);
or UO_1877 (O_1877,N_27403,N_27551);
nor UO_1878 (O_1878,N_25004,N_29412);
xor UO_1879 (O_1879,N_27022,N_26264);
or UO_1880 (O_1880,N_26682,N_28686);
nor UO_1881 (O_1881,N_25559,N_28845);
xnor UO_1882 (O_1882,N_25335,N_27340);
nand UO_1883 (O_1883,N_29983,N_29224);
xor UO_1884 (O_1884,N_27459,N_29140);
or UO_1885 (O_1885,N_28599,N_28802);
or UO_1886 (O_1886,N_27239,N_25140);
nand UO_1887 (O_1887,N_29500,N_25979);
nor UO_1888 (O_1888,N_26203,N_27594);
and UO_1889 (O_1889,N_27517,N_25428);
or UO_1890 (O_1890,N_29156,N_28540);
xor UO_1891 (O_1891,N_29772,N_29104);
xnor UO_1892 (O_1892,N_28330,N_28793);
nor UO_1893 (O_1893,N_27953,N_28882);
and UO_1894 (O_1894,N_27390,N_29484);
nand UO_1895 (O_1895,N_28717,N_25122);
or UO_1896 (O_1896,N_25867,N_26935);
or UO_1897 (O_1897,N_26676,N_27142);
or UO_1898 (O_1898,N_28426,N_26490);
nand UO_1899 (O_1899,N_28242,N_28066);
or UO_1900 (O_1900,N_28821,N_28984);
nor UO_1901 (O_1901,N_27591,N_29494);
xor UO_1902 (O_1902,N_29181,N_25450);
xor UO_1903 (O_1903,N_25670,N_27389);
or UO_1904 (O_1904,N_27974,N_29948);
nor UO_1905 (O_1905,N_28200,N_28168);
nand UO_1906 (O_1906,N_25197,N_25010);
or UO_1907 (O_1907,N_29785,N_29326);
or UO_1908 (O_1908,N_25941,N_28316);
nor UO_1909 (O_1909,N_29422,N_27257);
xor UO_1910 (O_1910,N_29960,N_29839);
nor UO_1911 (O_1911,N_28865,N_26268);
nor UO_1912 (O_1912,N_26647,N_26316);
nor UO_1913 (O_1913,N_26107,N_25935);
nand UO_1914 (O_1914,N_29265,N_29651);
nor UO_1915 (O_1915,N_27520,N_28775);
xor UO_1916 (O_1916,N_28138,N_28589);
xor UO_1917 (O_1917,N_28125,N_27983);
xnor UO_1918 (O_1918,N_29653,N_26695);
or UO_1919 (O_1919,N_26541,N_26455);
nand UO_1920 (O_1920,N_25834,N_29455);
nor UO_1921 (O_1921,N_25576,N_25676);
nor UO_1922 (O_1922,N_28827,N_28279);
xnor UO_1923 (O_1923,N_28573,N_26544);
or UO_1924 (O_1924,N_25328,N_28015);
and UO_1925 (O_1925,N_26542,N_26364);
nand UO_1926 (O_1926,N_28321,N_26548);
xor UO_1927 (O_1927,N_28598,N_28507);
nand UO_1928 (O_1928,N_27998,N_28409);
nor UO_1929 (O_1929,N_26304,N_25643);
nand UO_1930 (O_1930,N_27613,N_27229);
and UO_1931 (O_1931,N_28536,N_25331);
or UO_1932 (O_1932,N_25591,N_27721);
and UO_1933 (O_1933,N_25981,N_27541);
xor UO_1934 (O_1934,N_28382,N_29937);
and UO_1935 (O_1935,N_28713,N_26002);
nand UO_1936 (O_1936,N_25807,N_27010);
nand UO_1937 (O_1937,N_28963,N_25648);
or UO_1938 (O_1938,N_29841,N_29482);
xor UO_1939 (O_1939,N_27531,N_29101);
and UO_1940 (O_1940,N_28832,N_28262);
nand UO_1941 (O_1941,N_29209,N_26368);
nor UO_1942 (O_1942,N_26226,N_29498);
nor UO_1943 (O_1943,N_28129,N_28954);
nand UO_1944 (O_1944,N_29481,N_28374);
nand UO_1945 (O_1945,N_27720,N_28530);
and UO_1946 (O_1946,N_28909,N_27753);
and UO_1947 (O_1947,N_29631,N_25716);
and UO_1948 (O_1948,N_26299,N_29532);
xnor UO_1949 (O_1949,N_25886,N_26982);
or UO_1950 (O_1950,N_26828,N_29824);
nand UO_1951 (O_1951,N_29831,N_26761);
and UO_1952 (O_1952,N_26864,N_29546);
xnor UO_1953 (O_1953,N_25674,N_26004);
and UO_1954 (O_1954,N_29852,N_27249);
or UO_1955 (O_1955,N_29472,N_27940);
or UO_1956 (O_1956,N_26597,N_25899);
xor UO_1957 (O_1957,N_27147,N_28531);
and UO_1958 (O_1958,N_26197,N_25693);
nand UO_1959 (O_1959,N_29047,N_29071);
xnor UO_1960 (O_1960,N_28614,N_25729);
nand UO_1961 (O_1961,N_26187,N_29929);
or UO_1962 (O_1962,N_26977,N_27906);
xnor UO_1963 (O_1963,N_25324,N_29203);
or UO_1964 (O_1964,N_28064,N_29338);
or UO_1965 (O_1965,N_26386,N_29352);
or UO_1966 (O_1966,N_26469,N_26622);
nand UO_1967 (O_1967,N_28804,N_25540);
and UO_1968 (O_1968,N_26906,N_28830);
xor UO_1969 (O_1969,N_25832,N_26206);
and UO_1970 (O_1970,N_27343,N_26651);
and UO_1971 (O_1971,N_26401,N_25950);
nand UO_1972 (O_1972,N_28855,N_25980);
nor UO_1973 (O_1973,N_29161,N_26096);
xor UO_1974 (O_1974,N_29142,N_25811);
nor UO_1975 (O_1975,N_29032,N_25573);
and UO_1976 (O_1976,N_25201,N_26324);
nand UO_1977 (O_1977,N_28669,N_25193);
xnor UO_1978 (O_1978,N_29342,N_25016);
nand UO_1979 (O_1979,N_27179,N_26825);
nand UO_1980 (O_1980,N_26358,N_25109);
nand UO_1981 (O_1981,N_27934,N_28272);
nor UO_1982 (O_1982,N_26444,N_29851);
or UO_1983 (O_1983,N_29420,N_29711);
or UO_1984 (O_1984,N_26184,N_27439);
nor UO_1985 (O_1985,N_25677,N_26116);
xor UO_1986 (O_1986,N_28844,N_28153);
nand UO_1987 (O_1987,N_25226,N_28818);
nor UO_1988 (O_1988,N_25270,N_29992);
nor UO_1989 (O_1989,N_29153,N_25696);
nand UO_1990 (O_1990,N_28731,N_26330);
nand UO_1991 (O_1991,N_26176,N_26131);
nand UO_1992 (O_1992,N_25583,N_29621);
and UO_1993 (O_1993,N_27954,N_27292);
nand UO_1994 (O_1994,N_28161,N_29081);
nand UO_1995 (O_1995,N_26757,N_25350);
and UO_1996 (O_1996,N_27196,N_29765);
nand UO_1997 (O_1997,N_28246,N_25326);
or UO_1998 (O_1998,N_25441,N_27009);
nor UO_1999 (O_1999,N_28478,N_29808);
nor UO_2000 (O_2000,N_25360,N_29683);
xor UO_2001 (O_2001,N_29341,N_27364);
nor UO_2002 (O_2002,N_25575,N_28956);
or UO_2003 (O_2003,N_25382,N_27431);
xnor UO_2004 (O_2004,N_29910,N_28588);
xnor UO_2005 (O_2005,N_28877,N_26014);
nor UO_2006 (O_2006,N_29446,N_29199);
or UO_2007 (O_2007,N_25030,N_26052);
nor UO_2008 (O_2008,N_27211,N_28041);
nor UO_2009 (O_2009,N_27943,N_25212);
and UO_2010 (O_2010,N_25104,N_25588);
or UO_2011 (O_2011,N_25202,N_29250);
nand UO_2012 (O_2012,N_29348,N_28057);
nand UO_2013 (O_2013,N_26367,N_25397);
nand UO_2014 (O_2014,N_28660,N_25678);
nand UO_2015 (O_2015,N_25844,N_26133);
and UO_2016 (O_2016,N_26788,N_28274);
xor UO_2017 (O_2017,N_28938,N_25218);
nor UO_2018 (O_2018,N_25244,N_29926);
and UO_2019 (O_2019,N_25294,N_27038);
or UO_2020 (O_2020,N_27160,N_28806);
or UO_2021 (O_2021,N_29252,N_25216);
nand UO_2022 (O_2022,N_26314,N_25932);
nand UO_2023 (O_2023,N_25394,N_25902);
and UO_2024 (O_2024,N_29574,N_28256);
and UO_2025 (O_2025,N_29291,N_26374);
nor UO_2026 (O_2026,N_25446,N_29878);
nand UO_2027 (O_2027,N_26918,N_25771);
nand UO_2028 (O_2028,N_28078,N_28301);
nand UO_2029 (O_2029,N_27318,N_29693);
nor UO_2030 (O_2030,N_26868,N_26366);
and UO_2031 (O_2031,N_25208,N_28368);
nand UO_2032 (O_2032,N_26319,N_25993);
or UO_2033 (O_2033,N_25391,N_29585);
nor UO_2034 (O_2034,N_29394,N_26034);
or UO_2035 (O_2035,N_28238,N_28085);
xor UO_2036 (O_2036,N_27697,N_29632);
and UO_2037 (O_2037,N_25988,N_26978);
or UO_2038 (O_2038,N_27490,N_25246);
nor UO_2039 (O_2039,N_27492,N_25051);
or UO_2040 (O_2040,N_26037,N_29783);
nand UO_2041 (O_2041,N_26832,N_26734);
nor UO_2042 (O_2042,N_28269,N_27909);
xnor UO_2043 (O_2043,N_29279,N_29779);
xor UO_2044 (O_2044,N_25404,N_28694);
xnor UO_2045 (O_2045,N_29547,N_25254);
xor UO_2046 (O_2046,N_28776,N_25234);
xnor UO_2047 (O_2047,N_28151,N_26109);
xor UO_2048 (O_2048,N_26301,N_27138);
nand UO_2049 (O_2049,N_26442,N_26966);
nor UO_2050 (O_2050,N_25513,N_25431);
and UO_2051 (O_2051,N_25662,N_27182);
nor UO_2052 (O_2052,N_25255,N_26036);
xnor UO_2053 (O_2053,N_28341,N_29266);
xnor UO_2054 (O_2054,N_28513,N_27048);
and UO_2055 (O_2055,N_27049,N_26959);
and UO_2056 (O_2056,N_25289,N_27752);
xnor UO_2057 (O_2057,N_25485,N_25914);
xnor UO_2058 (O_2058,N_28286,N_28623);
nor UO_2059 (O_2059,N_26904,N_29014);
nor UO_2060 (O_2060,N_25130,N_26013);
xnor UO_2061 (O_2061,N_27831,N_27185);
xor UO_2062 (O_2062,N_28094,N_25533);
xnor UO_2063 (O_2063,N_28114,N_28022);
nor UO_2064 (O_2064,N_25772,N_28796);
nor UO_2065 (O_2065,N_29176,N_26684);
or UO_2066 (O_2066,N_29215,N_28010);
or UO_2067 (O_2067,N_25460,N_27224);
nand UO_2068 (O_2068,N_27408,N_27790);
and UO_2069 (O_2069,N_26008,N_27480);
nor UO_2070 (O_2070,N_29717,N_25597);
xnor UO_2071 (O_2071,N_28651,N_27463);
and UO_2072 (O_2072,N_27502,N_28839);
or UO_2073 (O_2073,N_27310,N_29213);
nor UO_2074 (O_2074,N_26010,N_26930);
and UO_2075 (O_2075,N_25420,N_25389);
and UO_2076 (O_2076,N_26110,N_28563);
and UO_2077 (O_2077,N_25984,N_28189);
or UO_2078 (O_2078,N_29386,N_27684);
xor UO_2079 (O_2079,N_27982,N_26230);
nand UO_2080 (O_2080,N_29221,N_28429);
and UO_2081 (O_2081,N_26886,N_27376);
and UO_2082 (O_2082,N_27513,N_25758);
nor UO_2083 (O_2083,N_28510,N_27342);
and UO_2084 (O_2084,N_29315,N_29260);
or UO_2085 (O_2085,N_29043,N_28503);
and UO_2086 (O_2086,N_26993,N_28325);
nor UO_2087 (O_2087,N_26997,N_28681);
nor UO_2088 (O_2088,N_28378,N_28915);
nand UO_2089 (O_2089,N_28937,N_28313);
nor UO_2090 (O_2090,N_29696,N_27440);
xnor UO_2091 (O_2091,N_25496,N_26807);
and UO_2092 (O_2092,N_25520,N_28489);
xnor UO_2093 (O_2093,N_27334,N_26986);
xnor UO_2094 (O_2094,N_28261,N_27204);
nand UO_2095 (O_2095,N_26641,N_25384);
nand UO_2096 (O_2096,N_25237,N_26479);
and UO_2097 (O_2097,N_26235,N_25731);
xor UO_2098 (O_2098,N_28732,N_25523);
and UO_2099 (O_2099,N_29075,N_26356);
xnor UO_2100 (O_2100,N_29391,N_26625);
or UO_2101 (O_2101,N_28864,N_26160);
or UO_2102 (O_2102,N_25561,N_26768);
nand UO_2103 (O_2103,N_27612,N_26072);
or UO_2104 (O_2104,N_28342,N_29977);
xor UO_2105 (O_2105,N_26102,N_26063);
nor UO_2106 (O_2106,N_26260,N_25322);
and UO_2107 (O_2107,N_27299,N_25097);
or UO_2108 (O_2108,N_28742,N_25853);
nand UO_2109 (O_2109,N_26489,N_27962);
or UO_2110 (O_2110,N_28788,N_27623);
xor UO_2111 (O_2111,N_29739,N_29610);
nor UO_2112 (O_2112,N_25996,N_26168);
nand UO_2113 (O_2113,N_28275,N_28749);
or UO_2114 (O_2114,N_26758,N_29954);
and UO_2115 (O_2115,N_28194,N_29847);
nand UO_2116 (O_2116,N_26070,N_27484);
nor UO_2117 (O_2117,N_29174,N_27027);
nor UO_2118 (O_2118,N_26732,N_27828);
and UO_2119 (O_2119,N_29665,N_25759);
xnor UO_2120 (O_2120,N_29050,N_29243);
and UO_2121 (O_2121,N_26569,N_26914);
xor UO_2122 (O_2122,N_28229,N_27381);
or UO_2123 (O_2123,N_26404,N_29860);
xor UO_2124 (O_2124,N_25554,N_27586);
and UO_2125 (O_2125,N_27532,N_29589);
xor UO_2126 (O_2126,N_26385,N_29790);
or UO_2127 (O_2127,N_29496,N_29144);
nor UO_2128 (O_2128,N_28263,N_27324);
or UO_2129 (O_2129,N_25403,N_27860);
and UO_2130 (O_2130,N_25107,N_27788);
nand UO_2131 (O_2131,N_26867,N_28988);
or UO_2132 (O_2132,N_28880,N_25997);
nor UO_2133 (O_2133,N_28773,N_29798);
or UO_2134 (O_2134,N_25881,N_29120);
or UO_2135 (O_2135,N_26424,N_27539);
nand UO_2136 (O_2136,N_28422,N_26360);
xnor UO_2137 (O_2137,N_25494,N_26784);
nand UO_2138 (O_2138,N_27183,N_25243);
nor UO_2139 (O_2139,N_28655,N_26422);
nand UO_2140 (O_2140,N_25401,N_25940);
nor UO_2141 (O_2141,N_28244,N_25547);
nand UO_2142 (O_2142,N_27467,N_27981);
and UO_2143 (O_2143,N_26791,N_28627);
xor UO_2144 (O_2144,N_29825,N_25275);
nor UO_2145 (O_2145,N_25657,N_27473);
xor UO_2146 (O_2146,N_29204,N_25538);
nor UO_2147 (O_2147,N_29655,N_26459);
nand UO_2148 (O_2148,N_29949,N_29198);
and UO_2149 (O_2149,N_25694,N_28529);
xnor UO_2150 (O_2150,N_29062,N_25348);
and UO_2151 (O_2151,N_27741,N_28505);
and UO_2152 (O_2152,N_28691,N_25873);
nand UO_2153 (O_2153,N_27521,N_25924);
xor UO_2154 (O_2154,N_29966,N_26245);
nand UO_2155 (O_2155,N_29707,N_25457);
and UO_2156 (O_2156,N_25586,N_29701);
and UO_2157 (O_2157,N_25818,N_26837);
and UO_2158 (O_2158,N_26053,N_25703);
xor UO_2159 (O_2159,N_29510,N_26091);
xnor UO_2160 (O_2160,N_27969,N_27227);
and UO_2161 (O_2161,N_27332,N_27785);
nor UO_2162 (O_2162,N_25711,N_29000);
and UO_2163 (O_2163,N_25532,N_29792);
xor UO_2164 (O_2164,N_29310,N_26113);
and UO_2165 (O_2165,N_28605,N_28224);
or UO_2166 (O_2166,N_29576,N_28326);
nand UO_2167 (O_2167,N_28213,N_26005);
nor UO_2168 (O_2168,N_25972,N_28926);
or UO_2169 (O_2169,N_27213,N_29863);
xor UO_2170 (O_2170,N_25869,N_29514);
xnor UO_2171 (O_2171,N_29959,N_29787);
nand UO_2172 (O_2172,N_25351,N_26307);
nand UO_2173 (O_2173,N_25780,N_27939);
nor UO_2174 (O_2174,N_26933,N_27036);
and UO_2175 (O_2175,N_26043,N_29290);
or UO_2176 (O_2176,N_28862,N_29505);
nand UO_2177 (O_2177,N_29671,N_26320);
nand UO_2178 (O_2178,N_29261,N_25164);
nor UO_2179 (O_2179,N_27464,N_25931);
xor UO_2180 (O_2180,N_25352,N_28025);
nor UO_2181 (O_2181,N_26683,N_29953);
or UO_2182 (O_2182,N_29699,N_25224);
nor UO_2183 (O_2183,N_29024,N_27588);
and UO_2184 (O_2184,N_27014,N_28225);
and UO_2185 (O_2185,N_27148,N_25589);
or UO_2186 (O_2186,N_28111,N_26589);
and UO_2187 (O_2187,N_26501,N_26843);
nor UO_2188 (O_2188,N_29119,N_25862);
xnor UO_2189 (O_2189,N_28769,N_29986);
and UO_2190 (O_2190,N_25154,N_29255);
xnor UO_2191 (O_2191,N_27763,N_25367);
and UO_2192 (O_2192,N_29820,N_27165);
or UO_2193 (O_2193,N_25257,N_25189);
nor UO_2194 (O_2194,N_25406,N_25652);
nand UO_2195 (O_2195,N_25396,N_27698);
xor UO_2196 (O_2196,N_28551,N_29127);
and UO_2197 (O_2197,N_25304,N_29374);
nand UO_2198 (O_2198,N_25865,N_28178);
and UO_2199 (O_2199,N_26649,N_26303);
or UO_2200 (O_2200,N_29826,N_27614);
nand UO_2201 (O_2201,N_29010,N_29596);
nor UO_2202 (O_2202,N_25149,N_27726);
nand UO_2203 (O_2203,N_25220,N_25062);
nor UO_2204 (O_2204,N_28514,N_26963);
nor UO_2205 (O_2205,N_29503,N_27578);
nor UO_2206 (O_2206,N_28280,N_25472);
nor UO_2207 (O_2207,N_29105,N_26743);
and UO_2208 (O_2208,N_25074,N_27132);
nand UO_2209 (O_2209,N_28201,N_29113);
and UO_2210 (O_2210,N_28097,N_29362);
nor UO_2211 (O_2211,N_29288,N_28322);
xor UO_2212 (O_2212,N_29991,N_28747);
nand UO_2213 (O_2213,N_25007,N_26348);
and UO_2214 (O_2214,N_25043,N_26159);
nor UO_2215 (O_2215,N_25035,N_26069);
or UO_2216 (O_2216,N_26932,N_28197);
nand UO_2217 (O_2217,N_29624,N_29408);
xor UO_2218 (O_2218,N_28782,N_25196);
nand UO_2219 (O_2219,N_26727,N_25357);
and UO_2220 (O_2220,N_26598,N_27150);
or UO_2221 (O_2221,N_25120,N_25481);
nand UO_2222 (O_2222,N_26781,N_29597);
or UO_2223 (O_2223,N_29832,N_27602);
nand UO_2224 (O_2224,N_29705,N_29654);
or UO_2225 (O_2225,N_26306,N_28438);
or UO_2226 (O_2226,N_28497,N_25622);
xnor UO_2227 (O_2227,N_25086,N_29996);
or UO_2228 (O_2228,N_26224,N_26079);
nand UO_2229 (O_2229,N_28466,N_26099);
nand UO_2230 (O_2230,N_25815,N_27554);
nor UO_2231 (O_2231,N_28460,N_25000);
and UO_2232 (O_2232,N_26336,N_26610);
and UO_2233 (O_2233,N_26409,N_25066);
and UO_2234 (O_2234,N_28173,N_27676);
or UO_2235 (O_2235,N_27857,N_25607);
nand UO_2236 (O_2236,N_28546,N_25974);
nand UO_2237 (O_2237,N_26411,N_25114);
or UO_2238 (O_2238,N_28160,N_25229);
and UO_2239 (O_2239,N_29134,N_28219);
and UO_2240 (O_2240,N_28751,N_27291);
nand UO_2241 (O_2241,N_26139,N_28106);
nor UO_2242 (O_2242,N_28848,N_27526);
or UO_2243 (O_2243,N_28145,N_28501);
xnor UO_2244 (O_2244,N_27980,N_27505);
xor UO_2245 (O_2245,N_26812,N_29880);
nor UO_2246 (O_2246,N_26406,N_28112);
xnor UO_2247 (O_2247,N_25810,N_28967);
and UO_2248 (O_2248,N_26814,N_26458);
xor UO_2249 (O_2249,N_29564,N_29036);
or UO_2250 (O_2250,N_28344,N_25008);
and UO_2251 (O_2251,N_25702,N_25912);
or UO_2252 (O_2252,N_29867,N_28863);
nor UO_2253 (O_2253,N_27882,N_28626);
nor UO_2254 (O_2254,N_26990,N_28165);
nand UO_2255 (O_2255,N_29528,N_29517);
xnor UO_2256 (O_2256,N_28650,N_26879);
nor UO_2257 (O_2257,N_28252,N_29529);
xor UO_2258 (O_2258,N_29234,N_27636);
nor UO_2259 (O_2259,N_25096,N_29123);
nand UO_2260 (O_2260,N_29055,N_25829);
and UO_2261 (O_2261,N_25773,N_25282);
and UO_2262 (O_2262,N_27558,N_28023);
xor UO_2263 (O_2263,N_25655,N_25766);
nor UO_2264 (O_2264,N_26529,N_29895);
and UO_2265 (O_2265,N_28519,N_28458);
or UO_2266 (O_2266,N_25339,N_26282);
or UO_2267 (O_2267,N_28005,N_28116);
nor UO_2268 (O_2268,N_25649,N_28172);
or UO_2269 (O_2269,N_27406,N_28308);
xor UO_2270 (O_2270,N_26081,N_29969);
nand UO_2271 (O_2271,N_28545,N_28090);
and UO_2272 (O_2272,N_25133,N_29143);
xor UO_2273 (O_2273,N_27041,N_25057);
nand UO_2274 (O_2274,N_28480,N_25640);
xor UO_2275 (O_2275,N_25905,N_27844);
xor UO_2276 (O_2276,N_26111,N_28318);
or UO_2277 (O_2277,N_26687,N_29358);
xor UO_2278 (O_2278,N_27956,N_25839);
nand UO_2279 (O_2279,N_27888,N_27200);
nand UO_2280 (O_2280,N_29398,N_27193);
nand UO_2281 (O_2281,N_27316,N_25336);
nand UO_2282 (O_2282,N_29658,N_27899);
or UO_2283 (O_2283,N_27552,N_28914);
and UO_2284 (O_2284,N_27886,N_27952);
nor UO_2285 (O_2285,N_27696,N_27746);
nand UO_2286 (O_2286,N_26463,N_27051);
xor UO_2287 (O_2287,N_27817,N_27102);
nor UO_2288 (O_2288,N_25871,N_27468);
or UO_2289 (O_2289,N_28593,N_29553);
and UO_2290 (O_2290,N_29220,N_29838);
and UO_2291 (O_2291,N_27571,N_29483);
nand UO_2292 (O_2292,N_27409,N_25332);
xnor UO_2293 (O_2293,N_29379,N_29964);
nor UO_2294 (O_2294,N_29962,N_28436);
or UO_2295 (O_2295,N_25969,N_29871);
and UO_2296 (O_2296,N_28526,N_26937);
and UO_2297 (O_2297,N_26487,N_29931);
and UO_2298 (O_2298,N_26836,N_28648);
nand UO_2299 (O_2299,N_28958,N_27805);
nor UO_2300 (O_2300,N_25029,N_29442);
xor UO_2301 (O_2301,N_29186,N_28124);
xor UO_2302 (O_2302,N_28029,N_26830);
nor UO_2303 (O_2303,N_27083,N_29275);
nor UO_2304 (O_2304,N_27674,N_27621);
xnor UO_2305 (O_2305,N_26579,N_27799);
nor UO_2306 (O_2306,N_29764,N_25602);
and UO_2307 (O_2307,N_25636,N_26760);
xor UO_2308 (O_2308,N_29112,N_26703);
xnor UO_2309 (O_2309,N_26075,N_26893);
nand UO_2310 (O_2310,N_26242,N_28567);
xnor UO_2311 (O_2311,N_27649,N_29999);
nor UO_2312 (O_2312,N_28562,N_26691);
or UO_2313 (O_2313,N_29357,N_26928);
and UO_2314 (O_2314,N_27705,N_27573);
nand UO_2315 (O_2315,N_27015,N_27168);
or UO_2316 (O_2316,N_28516,N_27631);
nand UO_2317 (O_2317,N_25801,N_26200);
xnor UO_2318 (O_2318,N_25820,N_27426);
and UO_2319 (O_2319,N_28303,N_25911);
nand UO_2320 (O_2320,N_29385,N_27092);
and UO_2321 (O_2321,N_27834,N_28872);
nor UO_2322 (O_2322,N_25267,N_25287);
nor UO_2323 (O_2323,N_29495,N_28720);
or UO_2324 (O_2324,N_29974,N_28730);
or UO_2325 (O_2325,N_27840,N_25642);
xor UO_2326 (O_2326,N_28615,N_27761);
xor UO_2327 (O_2327,N_29737,N_28759);
nand UO_2328 (O_2328,N_25987,N_25190);
and UO_2329 (O_2329,N_27330,N_26961);
and UO_2330 (O_2330,N_26174,N_25165);
and UO_2331 (O_2331,N_25235,N_25055);
nand UO_2332 (O_2332,N_25223,N_25827);
and UO_2333 (O_2333,N_29801,N_26954);
xor UO_2334 (O_2334,N_26552,N_27626);
and UO_2335 (O_2335,N_29925,N_27016);
xor UO_2336 (O_2336,N_28299,N_25265);
nor UO_2337 (O_2337,N_29837,N_28001);
xor UO_2338 (O_2338,N_25741,N_27932);
or UO_2339 (O_2339,N_28071,N_25568);
nand UO_2340 (O_2340,N_27547,N_28086);
and UO_2341 (O_2341,N_25802,N_28928);
or UO_2342 (O_2342,N_29834,N_25849);
nand UO_2343 (O_2343,N_26566,N_26050);
nor UO_2344 (O_2344,N_27329,N_26181);
xor UO_2345 (O_2345,N_25946,N_29736);
nand UO_2346 (O_2346,N_25025,N_28943);
xnor UO_2347 (O_2347,N_27067,N_28377);
nand UO_2348 (O_2348,N_27238,N_29163);
xnor UO_2349 (O_2349,N_27437,N_27725);
nor UO_2350 (O_2350,N_26915,N_25965);
nand UO_2351 (O_2351,N_29407,N_28892);
nor UO_2352 (O_2352,N_25595,N_29690);
nor UO_2353 (O_2353,N_25435,N_28081);
and UO_2354 (O_2354,N_26800,N_25671);
xor UO_2355 (O_2355,N_25175,N_27768);
and UO_2356 (O_2356,N_27488,N_26866);
or UO_2357 (O_2357,N_28659,N_26261);
nor UO_2358 (O_2358,N_27134,N_25411);
nor UO_2359 (O_2359,N_25028,N_28223);
or UO_2360 (O_2360,N_29881,N_27098);
nand UO_2361 (O_2361,N_29776,N_29872);
and UO_2362 (O_2362,N_28760,N_29399);
or UO_2363 (O_2363,N_26983,N_28879);
nand UO_2364 (O_2364,N_27216,N_26267);
and UO_2365 (O_2365,N_29850,N_29605);
xnor UO_2366 (O_2366,N_25529,N_27633);
and UO_2367 (O_2367,N_29263,N_29411);
and UO_2368 (O_2368,N_25126,N_26528);
or UO_2369 (O_2369,N_29074,N_28027);
nor UO_2370 (O_2370,N_27824,N_27121);
nor UO_2371 (O_2371,N_28553,N_26290);
nor UO_2372 (O_2372,N_27270,N_25044);
and UO_2373 (O_2373,N_25885,N_28767);
and UO_2374 (O_2374,N_25966,N_26194);
or UO_2375 (O_2375,N_29582,N_27846);
nor UO_2376 (O_2376,N_26644,N_27225);
nor UO_2377 (O_2377,N_27057,N_26723);
and UO_2378 (O_2378,N_29673,N_25374);
nor UO_2379 (O_2379,N_25769,N_25186);
or UO_2380 (O_2380,N_29922,N_27077);
and UO_2381 (O_2381,N_28451,N_28919);
xor UO_2382 (O_2382,N_28991,N_29800);
or UO_2383 (O_2383,N_26848,N_28329);
or UO_2384 (O_2384,N_28264,N_26496);
nor UO_2385 (O_2385,N_26753,N_28309);
xnor UO_2386 (O_2386,N_29286,N_25620);
nand UO_2387 (O_2387,N_27743,N_26637);
or UO_2388 (O_2388,N_28729,N_27657);
xor UO_2389 (O_2389,N_29828,N_29761);
or UO_2390 (O_2390,N_27605,N_28128);
or UO_2391 (O_2391,N_26241,N_25894);
nor UO_2392 (O_2392,N_26327,N_28897);
xor UO_2393 (O_2393,N_27683,N_28441);
nand UO_2394 (O_2394,N_26538,N_28554);
nand UO_2395 (O_2395,N_25545,N_28384);
and UO_2396 (O_2396,N_27295,N_27320);
or UO_2397 (O_2397,N_27680,N_29721);
nand UO_2398 (O_2398,N_26007,N_28245);
xnor UO_2399 (O_2399,N_26234,N_25835);
and UO_2400 (O_2400,N_28657,N_28423);
nor UO_2401 (O_2401,N_26725,N_28387);
xnor UO_2402 (O_2402,N_26931,N_26554);
nand UO_2403 (O_2403,N_28613,N_26511);
or UO_2404 (O_2404,N_27832,N_27197);
and UO_2405 (O_2405,N_27837,N_28718);
or UO_2406 (O_2406,N_26383,N_28267);
nor UO_2407 (O_2407,N_28684,N_29788);
or UO_2408 (O_2408,N_28304,N_25418);
xnor UO_2409 (O_2409,N_29525,N_25667);
xor UO_2410 (O_2410,N_27311,N_25634);
and UO_2411 (O_2411,N_29897,N_26068);
nand UO_2412 (O_2412,N_29752,N_26910);
and UO_2413 (O_2413,N_27287,N_28753);
or UO_2414 (O_2414,N_29329,N_28565);
and UO_2415 (O_2415,N_26849,N_29548);
and UO_2416 (O_2416,N_26410,N_29073);
or UO_2417 (O_2417,N_26952,N_25775);
nor UO_2418 (O_2418,N_27624,N_29414);
or UO_2419 (O_2419,N_26873,N_27855);
and UO_2420 (O_2420,N_25893,N_26427);
nor UO_2421 (O_2421,N_26347,N_26785);
xnor UO_2422 (O_2422,N_28831,N_25070);
or UO_2423 (O_2423,N_25909,N_26147);
or UO_2424 (O_2424,N_27564,N_26060);
nand UO_2425 (O_2425,N_25195,N_26787);
nor UO_2426 (O_2426,N_28486,N_28061);
or UO_2427 (O_2427,N_29766,N_27264);
xnor UO_2428 (O_2428,N_26436,N_27836);
or UO_2429 (O_2429,N_29920,N_28745);
or UO_2430 (O_2430,N_27219,N_29448);
nor UO_2431 (O_2431,N_27284,N_27465);
nor UO_2432 (O_2432,N_25489,N_28254);
or UO_2433 (O_2433,N_27895,N_28690);
xor UO_2434 (O_2434,N_29006,N_27584);
nand UO_2435 (O_2435,N_28902,N_26845);
and UO_2436 (O_2436,N_27362,N_29170);
nand UO_2437 (O_2437,N_27474,N_27111);
nor UO_2438 (O_2438,N_28170,N_29246);
nand UO_2439 (O_2439,N_27202,N_28955);
nand UO_2440 (O_2440,N_26452,N_29020);
xor UO_2441 (O_2441,N_25274,N_27948);
and UO_2442 (O_2442,N_28385,N_29578);
nand UO_2443 (O_2443,N_28652,N_29811);
xnor UO_2444 (O_2444,N_29859,N_28995);
and UO_2445 (O_2445,N_27367,N_28812);
xnor UO_2446 (O_2446,N_28597,N_26433);
xnor UO_2447 (O_2447,N_28443,N_29706);
xor UO_2448 (O_2448,N_28702,N_28397);
xnor UO_2449 (O_2449,N_25319,N_28506);
and UO_2450 (O_2450,N_26128,N_26392);
xor UO_2451 (O_2451,N_28649,N_29312);
or UO_2452 (O_2452,N_26087,N_29022);
xor UO_2453 (O_2453,N_28046,N_26333);
nor UO_2454 (O_2454,N_28999,N_28945);
nor UO_2455 (O_2455,N_26136,N_27378);
or UO_2456 (O_2456,N_28277,N_28798);
nor UO_2457 (O_2457,N_28206,N_26741);
and UO_2458 (O_2458,N_29148,N_25464);
xnor UO_2459 (O_2459,N_26980,N_28722);
xnor UO_2460 (O_2460,N_29427,N_25123);
and UO_2461 (O_2461,N_26331,N_29060);
and UO_2462 (O_2462,N_29599,N_26077);
and UO_2463 (O_2463,N_27143,N_26796);
nand UO_2464 (O_2464,N_28305,N_29211);
nand UO_2465 (O_2465,N_29295,N_25546);
or UO_2466 (O_2466,N_25478,N_27916);
nand UO_2467 (O_2467,N_29840,N_27880);
xnor UO_2468 (O_2468,N_27669,N_29115);
xor UO_2469 (O_2469,N_29921,N_27686);
nand UO_2470 (O_2470,N_26248,N_25429);
xor UO_2471 (O_2471,N_25864,N_28664);
and UO_2472 (O_2472,N_26624,N_26115);
nand UO_2473 (O_2473,N_29601,N_26633);
or UO_2474 (O_2474,N_27816,N_29429);
xnor UO_2475 (O_2475,N_28708,N_26185);
xor UO_2476 (O_2476,N_29767,N_27314);
and UO_2477 (O_2477,N_28680,N_25785);
nor UO_2478 (O_2478,N_29040,N_28347);
or UO_2479 (O_2479,N_29679,N_25483);
nand UO_2480 (O_2480,N_25506,N_25376);
nand UO_2481 (O_2481,N_28700,N_29301);
xnor UO_2482 (O_2482,N_28808,N_26325);
nand UO_2483 (O_2483,N_25334,N_27606);
xor UO_2484 (O_2484,N_26488,N_29994);
nand UO_2485 (O_2485,N_27927,N_27604);
nor UO_2486 (O_2486,N_26958,N_26239);
or UO_2487 (O_2487,N_29426,N_29743);
nor UO_2488 (O_2488,N_28653,N_25320);
nor UO_2489 (O_2489,N_29854,N_28394);
or UO_2490 (O_2490,N_28069,N_26671);
nor UO_2491 (O_2491,N_25036,N_28258);
and UO_2492 (O_2492,N_28365,N_27301);
or UO_2493 (O_2493,N_26988,N_27748);
xnor UO_2494 (O_2494,N_28068,N_25488);
xnor UO_2495 (O_2495,N_26024,N_26209);
and UO_2496 (O_2496,N_28965,N_28082);
and UO_2497 (O_2497,N_25167,N_27955);
nor UO_2498 (O_2498,N_28043,N_25557);
or UO_2499 (O_2499,N_29754,N_27590);
or UO_2500 (O_2500,N_25983,N_25214);
nand UO_2501 (O_2501,N_25548,N_25033);
nand UO_2502 (O_2502,N_26258,N_29018);
and UO_2503 (O_2503,N_25933,N_25047);
and UO_2504 (O_2504,N_25444,N_29866);
nand UO_2505 (O_2505,N_28341,N_28930);
or UO_2506 (O_2506,N_29260,N_25204);
and UO_2507 (O_2507,N_29374,N_28630);
and UO_2508 (O_2508,N_26012,N_29606);
nand UO_2509 (O_2509,N_27495,N_27208);
and UO_2510 (O_2510,N_26194,N_28658);
nand UO_2511 (O_2511,N_27017,N_29883);
and UO_2512 (O_2512,N_26707,N_27420);
or UO_2513 (O_2513,N_27955,N_27927);
xnor UO_2514 (O_2514,N_27445,N_25858);
and UO_2515 (O_2515,N_26632,N_29351);
and UO_2516 (O_2516,N_25072,N_27644);
nand UO_2517 (O_2517,N_25903,N_25962);
or UO_2518 (O_2518,N_28312,N_29815);
xnor UO_2519 (O_2519,N_28804,N_28376);
nand UO_2520 (O_2520,N_25755,N_26840);
nand UO_2521 (O_2521,N_28540,N_27872);
or UO_2522 (O_2522,N_28663,N_25412);
xnor UO_2523 (O_2523,N_25739,N_27568);
or UO_2524 (O_2524,N_29562,N_29714);
or UO_2525 (O_2525,N_26626,N_25577);
nor UO_2526 (O_2526,N_25339,N_27782);
xnor UO_2527 (O_2527,N_29316,N_29582);
xor UO_2528 (O_2528,N_25826,N_25973);
nand UO_2529 (O_2529,N_29184,N_26927);
or UO_2530 (O_2530,N_29049,N_29933);
nor UO_2531 (O_2531,N_26207,N_27313);
or UO_2532 (O_2532,N_27547,N_29829);
or UO_2533 (O_2533,N_25015,N_28927);
and UO_2534 (O_2534,N_29688,N_25291);
and UO_2535 (O_2535,N_26090,N_29652);
and UO_2536 (O_2536,N_27426,N_28405);
nor UO_2537 (O_2537,N_29852,N_26249);
nor UO_2538 (O_2538,N_25033,N_28790);
and UO_2539 (O_2539,N_26939,N_28250);
nor UO_2540 (O_2540,N_29919,N_28468);
or UO_2541 (O_2541,N_29083,N_25820);
and UO_2542 (O_2542,N_26216,N_27428);
nand UO_2543 (O_2543,N_29951,N_28350);
or UO_2544 (O_2544,N_28015,N_27052);
nand UO_2545 (O_2545,N_29666,N_26929);
or UO_2546 (O_2546,N_26416,N_26332);
xnor UO_2547 (O_2547,N_26334,N_25526);
nand UO_2548 (O_2548,N_28304,N_29754);
nor UO_2549 (O_2549,N_26629,N_25912);
and UO_2550 (O_2550,N_26527,N_25871);
nor UO_2551 (O_2551,N_29641,N_25603);
xnor UO_2552 (O_2552,N_26490,N_28801);
and UO_2553 (O_2553,N_25691,N_25142);
nand UO_2554 (O_2554,N_28453,N_27815);
or UO_2555 (O_2555,N_29058,N_27433);
nor UO_2556 (O_2556,N_28521,N_29775);
xor UO_2557 (O_2557,N_28828,N_28812);
nand UO_2558 (O_2558,N_27587,N_26906);
nand UO_2559 (O_2559,N_28935,N_28264);
xor UO_2560 (O_2560,N_25961,N_29278);
nor UO_2561 (O_2561,N_25385,N_28242);
xnor UO_2562 (O_2562,N_29144,N_25064);
nand UO_2563 (O_2563,N_28535,N_29275);
nor UO_2564 (O_2564,N_29034,N_28409);
or UO_2565 (O_2565,N_28275,N_26100);
and UO_2566 (O_2566,N_27189,N_26618);
nand UO_2567 (O_2567,N_28878,N_26042);
nor UO_2568 (O_2568,N_29823,N_29275);
xor UO_2569 (O_2569,N_25901,N_28658);
or UO_2570 (O_2570,N_28947,N_29735);
nand UO_2571 (O_2571,N_25618,N_28157);
nand UO_2572 (O_2572,N_29910,N_25373);
xor UO_2573 (O_2573,N_28453,N_28285);
or UO_2574 (O_2574,N_27775,N_25025);
or UO_2575 (O_2575,N_29440,N_25689);
or UO_2576 (O_2576,N_26472,N_29657);
nand UO_2577 (O_2577,N_27754,N_26409);
and UO_2578 (O_2578,N_28273,N_27396);
nor UO_2579 (O_2579,N_25611,N_29366);
or UO_2580 (O_2580,N_29979,N_29436);
and UO_2581 (O_2581,N_28616,N_27428);
and UO_2582 (O_2582,N_26210,N_26647);
and UO_2583 (O_2583,N_29862,N_27972);
and UO_2584 (O_2584,N_25693,N_28855);
or UO_2585 (O_2585,N_25763,N_26876);
or UO_2586 (O_2586,N_28943,N_29163);
nor UO_2587 (O_2587,N_25706,N_26323);
or UO_2588 (O_2588,N_25581,N_29130);
nand UO_2589 (O_2589,N_27555,N_26061);
xor UO_2590 (O_2590,N_29919,N_29986);
nand UO_2591 (O_2591,N_29715,N_26190);
nand UO_2592 (O_2592,N_25105,N_28072);
nand UO_2593 (O_2593,N_28979,N_26021);
and UO_2594 (O_2594,N_28822,N_28121);
xor UO_2595 (O_2595,N_25020,N_29169);
xor UO_2596 (O_2596,N_25727,N_29738);
or UO_2597 (O_2597,N_29090,N_28272);
nor UO_2598 (O_2598,N_29858,N_26303);
or UO_2599 (O_2599,N_26970,N_28341);
or UO_2600 (O_2600,N_29857,N_29960);
nand UO_2601 (O_2601,N_26061,N_26699);
nor UO_2602 (O_2602,N_26091,N_26888);
nor UO_2603 (O_2603,N_28732,N_25011);
nor UO_2604 (O_2604,N_25338,N_26552);
nor UO_2605 (O_2605,N_27133,N_28422);
nand UO_2606 (O_2606,N_29423,N_28242);
nor UO_2607 (O_2607,N_25220,N_25279);
nand UO_2608 (O_2608,N_27598,N_29107);
or UO_2609 (O_2609,N_25781,N_27097);
xnor UO_2610 (O_2610,N_25094,N_28418);
xor UO_2611 (O_2611,N_29042,N_26713);
nand UO_2612 (O_2612,N_29960,N_26829);
and UO_2613 (O_2613,N_28256,N_26322);
or UO_2614 (O_2614,N_26496,N_26869);
nor UO_2615 (O_2615,N_28255,N_29783);
xor UO_2616 (O_2616,N_27992,N_29554);
xor UO_2617 (O_2617,N_26305,N_25647);
nand UO_2618 (O_2618,N_25566,N_27172);
and UO_2619 (O_2619,N_25633,N_26242);
nand UO_2620 (O_2620,N_26761,N_28525);
and UO_2621 (O_2621,N_28769,N_27981);
nor UO_2622 (O_2622,N_26696,N_26837);
and UO_2623 (O_2623,N_28448,N_25936);
and UO_2624 (O_2624,N_29826,N_25405);
nor UO_2625 (O_2625,N_28721,N_27393);
xor UO_2626 (O_2626,N_26712,N_28125);
or UO_2627 (O_2627,N_29639,N_28336);
xor UO_2628 (O_2628,N_27024,N_29380);
xor UO_2629 (O_2629,N_29763,N_26046);
nor UO_2630 (O_2630,N_27456,N_25950);
or UO_2631 (O_2631,N_28711,N_29546);
or UO_2632 (O_2632,N_25075,N_27034);
and UO_2633 (O_2633,N_26421,N_28354);
and UO_2634 (O_2634,N_26917,N_27219);
or UO_2635 (O_2635,N_26732,N_29714);
or UO_2636 (O_2636,N_27620,N_28728);
nor UO_2637 (O_2637,N_25840,N_28765);
and UO_2638 (O_2638,N_29793,N_26126);
and UO_2639 (O_2639,N_29878,N_29096);
or UO_2640 (O_2640,N_26681,N_25250);
xnor UO_2641 (O_2641,N_27108,N_29579);
xor UO_2642 (O_2642,N_27448,N_27061);
xor UO_2643 (O_2643,N_27662,N_28517);
and UO_2644 (O_2644,N_26986,N_29264);
or UO_2645 (O_2645,N_27034,N_25384);
nor UO_2646 (O_2646,N_28116,N_26754);
xnor UO_2647 (O_2647,N_25148,N_25518);
or UO_2648 (O_2648,N_28560,N_27653);
nand UO_2649 (O_2649,N_28256,N_25550);
or UO_2650 (O_2650,N_25196,N_29060);
nand UO_2651 (O_2651,N_27991,N_26119);
or UO_2652 (O_2652,N_28284,N_26932);
and UO_2653 (O_2653,N_28709,N_28563);
or UO_2654 (O_2654,N_28075,N_29099);
or UO_2655 (O_2655,N_26905,N_25185);
nor UO_2656 (O_2656,N_25295,N_26488);
nand UO_2657 (O_2657,N_25898,N_29856);
nor UO_2658 (O_2658,N_25800,N_25783);
nor UO_2659 (O_2659,N_25425,N_25847);
nand UO_2660 (O_2660,N_25853,N_25949);
xor UO_2661 (O_2661,N_28662,N_28424);
xnor UO_2662 (O_2662,N_28321,N_28524);
or UO_2663 (O_2663,N_26829,N_26143);
nor UO_2664 (O_2664,N_26044,N_27213);
nand UO_2665 (O_2665,N_27732,N_29443);
or UO_2666 (O_2666,N_27584,N_29539);
or UO_2667 (O_2667,N_26426,N_28135);
xor UO_2668 (O_2668,N_25769,N_28299);
or UO_2669 (O_2669,N_26486,N_26540);
xor UO_2670 (O_2670,N_29576,N_27603);
xnor UO_2671 (O_2671,N_26919,N_25648);
and UO_2672 (O_2672,N_29206,N_25885);
and UO_2673 (O_2673,N_28123,N_27680);
nor UO_2674 (O_2674,N_29250,N_27042);
nor UO_2675 (O_2675,N_25621,N_29706);
nor UO_2676 (O_2676,N_25299,N_28747);
xnor UO_2677 (O_2677,N_25054,N_25688);
and UO_2678 (O_2678,N_28402,N_26392);
and UO_2679 (O_2679,N_28751,N_28708);
xor UO_2680 (O_2680,N_29163,N_28289);
xnor UO_2681 (O_2681,N_27513,N_28490);
nand UO_2682 (O_2682,N_27764,N_29115);
nand UO_2683 (O_2683,N_25423,N_26570);
nor UO_2684 (O_2684,N_27510,N_26644);
nand UO_2685 (O_2685,N_28005,N_27611);
or UO_2686 (O_2686,N_28824,N_29390);
xnor UO_2687 (O_2687,N_27106,N_28892);
nor UO_2688 (O_2688,N_29478,N_25037);
xnor UO_2689 (O_2689,N_28180,N_27176);
or UO_2690 (O_2690,N_26243,N_26652);
or UO_2691 (O_2691,N_28836,N_26282);
nor UO_2692 (O_2692,N_26930,N_28421);
nand UO_2693 (O_2693,N_27930,N_27354);
and UO_2694 (O_2694,N_27307,N_28972);
or UO_2695 (O_2695,N_26077,N_29086);
xnor UO_2696 (O_2696,N_27567,N_26210);
or UO_2697 (O_2697,N_29530,N_29104);
and UO_2698 (O_2698,N_27216,N_25227);
and UO_2699 (O_2699,N_28767,N_27004);
xor UO_2700 (O_2700,N_29672,N_28797);
and UO_2701 (O_2701,N_25153,N_27100);
or UO_2702 (O_2702,N_25011,N_28357);
or UO_2703 (O_2703,N_25363,N_29919);
or UO_2704 (O_2704,N_26660,N_25112);
nor UO_2705 (O_2705,N_27916,N_25013);
nand UO_2706 (O_2706,N_29402,N_29843);
nor UO_2707 (O_2707,N_29365,N_29560);
or UO_2708 (O_2708,N_28279,N_28689);
xnor UO_2709 (O_2709,N_27897,N_26191);
nor UO_2710 (O_2710,N_25160,N_29536);
nand UO_2711 (O_2711,N_28500,N_27082);
or UO_2712 (O_2712,N_25171,N_25160);
nand UO_2713 (O_2713,N_29563,N_26590);
or UO_2714 (O_2714,N_28765,N_29219);
xor UO_2715 (O_2715,N_25614,N_28283);
xor UO_2716 (O_2716,N_27694,N_28996);
nand UO_2717 (O_2717,N_29149,N_26097);
xnor UO_2718 (O_2718,N_26666,N_25224);
or UO_2719 (O_2719,N_26177,N_27069);
nand UO_2720 (O_2720,N_28102,N_25476);
nand UO_2721 (O_2721,N_27718,N_27979);
xnor UO_2722 (O_2722,N_27449,N_26234);
and UO_2723 (O_2723,N_29641,N_29235);
and UO_2724 (O_2724,N_26936,N_25550);
xor UO_2725 (O_2725,N_28609,N_27276);
or UO_2726 (O_2726,N_25020,N_25561);
nand UO_2727 (O_2727,N_26503,N_28356);
nor UO_2728 (O_2728,N_28500,N_29081);
and UO_2729 (O_2729,N_25284,N_29489);
xor UO_2730 (O_2730,N_29659,N_26766);
nand UO_2731 (O_2731,N_25007,N_25383);
nor UO_2732 (O_2732,N_26257,N_29661);
or UO_2733 (O_2733,N_26464,N_28527);
or UO_2734 (O_2734,N_25176,N_26437);
xnor UO_2735 (O_2735,N_27820,N_27035);
and UO_2736 (O_2736,N_26105,N_29060);
and UO_2737 (O_2737,N_26435,N_29251);
nor UO_2738 (O_2738,N_26013,N_25365);
nor UO_2739 (O_2739,N_26342,N_29644);
xnor UO_2740 (O_2740,N_27625,N_25442);
nor UO_2741 (O_2741,N_25030,N_25843);
and UO_2742 (O_2742,N_29656,N_26471);
and UO_2743 (O_2743,N_25121,N_26519);
xor UO_2744 (O_2744,N_28505,N_25952);
xnor UO_2745 (O_2745,N_29484,N_29669);
and UO_2746 (O_2746,N_26946,N_28786);
and UO_2747 (O_2747,N_27383,N_28650);
nand UO_2748 (O_2748,N_27016,N_26630);
and UO_2749 (O_2749,N_26682,N_27947);
and UO_2750 (O_2750,N_26992,N_27065);
nor UO_2751 (O_2751,N_26201,N_25478);
xor UO_2752 (O_2752,N_28321,N_26421);
nor UO_2753 (O_2753,N_25859,N_28132);
or UO_2754 (O_2754,N_25448,N_27036);
xor UO_2755 (O_2755,N_28575,N_27708);
and UO_2756 (O_2756,N_28976,N_25020);
nand UO_2757 (O_2757,N_25736,N_27234);
xnor UO_2758 (O_2758,N_27127,N_28362);
nand UO_2759 (O_2759,N_27651,N_25488);
nor UO_2760 (O_2760,N_28240,N_26766);
nor UO_2761 (O_2761,N_27243,N_26961);
or UO_2762 (O_2762,N_27363,N_29781);
or UO_2763 (O_2763,N_27991,N_26943);
and UO_2764 (O_2764,N_26098,N_26863);
nand UO_2765 (O_2765,N_28221,N_29709);
nor UO_2766 (O_2766,N_28609,N_29975);
and UO_2767 (O_2767,N_26845,N_28362);
and UO_2768 (O_2768,N_27956,N_29459);
and UO_2769 (O_2769,N_27814,N_28756);
nor UO_2770 (O_2770,N_27192,N_26814);
and UO_2771 (O_2771,N_27806,N_28380);
or UO_2772 (O_2772,N_26069,N_25639);
and UO_2773 (O_2773,N_27782,N_28127);
nand UO_2774 (O_2774,N_29908,N_28494);
nand UO_2775 (O_2775,N_29426,N_26227);
xnor UO_2776 (O_2776,N_28528,N_27806);
nor UO_2777 (O_2777,N_26875,N_28993);
nand UO_2778 (O_2778,N_29352,N_28507);
nor UO_2779 (O_2779,N_28340,N_26092);
nor UO_2780 (O_2780,N_28882,N_29012);
and UO_2781 (O_2781,N_25577,N_28375);
nand UO_2782 (O_2782,N_28005,N_29597);
nand UO_2783 (O_2783,N_28608,N_25696);
xnor UO_2784 (O_2784,N_28033,N_27179);
nand UO_2785 (O_2785,N_28161,N_28935);
nor UO_2786 (O_2786,N_27193,N_25810);
nand UO_2787 (O_2787,N_27715,N_29657);
nor UO_2788 (O_2788,N_27398,N_28972);
xnor UO_2789 (O_2789,N_26099,N_26179);
or UO_2790 (O_2790,N_28939,N_26968);
nand UO_2791 (O_2791,N_27256,N_29003);
nand UO_2792 (O_2792,N_25536,N_26669);
and UO_2793 (O_2793,N_29843,N_27519);
and UO_2794 (O_2794,N_28787,N_27345);
nand UO_2795 (O_2795,N_25921,N_29184);
nand UO_2796 (O_2796,N_29988,N_26403);
or UO_2797 (O_2797,N_25630,N_29125);
and UO_2798 (O_2798,N_26600,N_28522);
nand UO_2799 (O_2799,N_29370,N_28618);
xnor UO_2800 (O_2800,N_28989,N_26109);
nand UO_2801 (O_2801,N_25013,N_27492);
nor UO_2802 (O_2802,N_27890,N_28090);
xnor UO_2803 (O_2803,N_26264,N_25008);
and UO_2804 (O_2804,N_25544,N_28920);
and UO_2805 (O_2805,N_29818,N_27559);
or UO_2806 (O_2806,N_29622,N_26477);
or UO_2807 (O_2807,N_27619,N_26829);
nand UO_2808 (O_2808,N_29920,N_29068);
nand UO_2809 (O_2809,N_29983,N_25178);
nor UO_2810 (O_2810,N_25608,N_25666);
or UO_2811 (O_2811,N_29902,N_28421);
or UO_2812 (O_2812,N_25751,N_26549);
and UO_2813 (O_2813,N_28229,N_25728);
xnor UO_2814 (O_2814,N_29594,N_26646);
and UO_2815 (O_2815,N_25491,N_29728);
and UO_2816 (O_2816,N_27285,N_27588);
nor UO_2817 (O_2817,N_26536,N_29052);
or UO_2818 (O_2818,N_27446,N_25314);
or UO_2819 (O_2819,N_26722,N_28694);
or UO_2820 (O_2820,N_25519,N_25222);
and UO_2821 (O_2821,N_26953,N_29465);
and UO_2822 (O_2822,N_26035,N_29512);
nor UO_2823 (O_2823,N_25745,N_29547);
or UO_2824 (O_2824,N_26570,N_29014);
nand UO_2825 (O_2825,N_28799,N_25942);
nand UO_2826 (O_2826,N_26039,N_29694);
nand UO_2827 (O_2827,N_27165,N_29238);
xnor UO_2828 (O_2828,N_28040,N_26850);
nor UO_2829 (O_2829,N_27468,N_29885);
nand UO_2830 (O_2830,N_29626,N_25229);
nor UO_2831 (O_2831,N_26708,N_29112);
or UO_2832 (O_2832,N_26037,N_26459);
and UO_2833 (O_2833,N_26867,N_26334);
or UO_2834 (O_2834,N_27767,N_28228);
nor UO_2835 (O_2835,N_27076,N_28257);
xor UO_2836 (O_2836,N_25796,N_25547);
xor UO_2837 (O_2837,N_25315,N_27827);
nand UO_2838 (O_2838,N_26475,N_28377);
and UO_2839 (O_2839,N_26520,N_29934);
and UO_2840 (O_2840,N_28957,N_29946);
or UO_2841 (O_2841,N_25639,N_28701);
xnor UO_2842 (O_2842,N_29771,N_28400);
and UO_2843 (O_2843,N_28528,N_26914);
xnor UO_2844 (O_2844,N_28364,N_28756);
nor UO_2845 (O_2845,N_26924,N_28897);
and UO_2846 (O_2846,N_25233,N_28145);
xnor UO_2847 (O_2847,N_26234,N_28304);
and UO_2848 (O_2848,N_29988,N_29019);
xor UO_2849 (O_2849,N_28136,N_27598);
or UO_2850 (O_2850,N_25388,N_29208);
xnor UO_2851 (O_2851,N_28422,N_28960);
nor UO_2852 (O_2852,N_26599,N_29136);
nor UO_2853 (O_2853,N_26703,N_27744);
xnor UO_2854 (O_2854,N_29048,N_25837);
nor UO_2855 (O_2855,N_26441,N_25102);
xor UO_2856 (O_2856,N_28066,N_25653);
and UO_2857 (O_2857,N_25212,N_26143);
xnor UO_2858 (O_2858,N_29696,N_27441);
xor UO_2859 (O_2859,N_25821,N_27356);
nor UO_2860 (O_2860,N_25248,N_28349);
xnor UO_2861 (O_2861,N_26050,N_27959);
or UO_2862 (O_2862,N_26636,N_27364);
nand UO_2863 (O_2863,N_27267,N_27694);
and UO_2864 (O_2864,N_27656,N_29391);
or UO_2865 (O_2865,N_26361,N_27179);
nand UO_2866 (O_2866,N_28652,N_26227);
xnor UO_2867 (O_2867,N_29698,N_27422);
or UO_2868 (O_2868,N_27511,N_26658);
and UO_2869 (O_2869,N_26683,N_25840);
nor UO_2870 (O_2870,N_27434,N_26487);
or UO_2871 (O_2871,N_27648,N_27174);
or UO_2872 (O_2872,N_29134,N_27389);
nor UO_2873 (O_2873,N_28354,N_26801);
xor UO_2874 (O_2874,N_28014,N_28725);
nor UO_2875 (O_2875,N_25949,N_25470);
nor UO_2876 (O_2876,N_25051,N_28008);
or UO_2877 (O_2877,N_27231,N_27120);
nor UO_2878 (O_2878,N_28706,N_28433);
or UO_2879 (O_2879,N_25071,N_27388);
nand UO_2880 (O_2880,N_28912,N_25349);
and UO_2881 (O_2881,N_27295,N_26348);
nand UO_2882 (O_2882,N_27627,N_29903);
xor UO_2883 (O_2883,N_25586,N_27188);
nand UO_2884 (O_2884,N_27284,N_25915);
and UO_2885 (O_2885,N_29468,N_27909);
and UO_2886 (O_2886,N_28721,N_29204);
or UO_2887 (O_2887,N_28397,N_28013);
or UO_2888 (O_2888,N_26166,N_27180);
and UO_2889 (O_2889,N_27706,N_29070);
nor UO_2890 (O_2890,N_25645,N_25486);
or UO_2891 (O_2891,N_29005,N_25211);
nand UO_2892 (O_2892,N_27804,N_29610);
nor UO_2893 (O_2893,N_26381,N_26546);
nand UO_2894 (O_2894,N_29727,N_27636);
nor UO_2895 (O_2895,N_28502,N_28109);
and UO_2896 (O_2896,N_27215,N_26451);
xnor UO_2897 (O_2897,N_29906,N_25446);
or UO_2898 (O_2898,N_29973,N_28613);
or UO_2899 (O_2899,N_28406,N_29510);
xor UO_2900 (O_2900,N_28707,N_26699);
xnor UO_2901 (O_2901,N_29032,N_29751);
nor UO_2902 (O_2902,N_26235,N_28331);
nand UO_2903 (O_2903,N_27394,N_27159);
or UO_2904 (O_2904,N_29223,N_27212);
and UO_2905 (O_2905,N_29401,N_29644);
nor UO_2906 (O_2906,N_29014,N_27490);
nor UO_2907 (O_2907,N_28263,N_28193);
xor UO_2908 (O_2908,N_25415,N_26602);
and UO_2909 (O_2909,N_29018,N_28193);
or UO_2910 (O_2910,N_29962,N_25004);
or UO_2911 (O_2911,N_25010,N_25630);
nand UO_2912 (O_2912,N_29799,N_25696);
and UO_2913 (O_2913,N_25485,N_26570);
or UO_2914 (O_2914,N_29566,N_25538);
or UO_2915 (O_2915,N_28099,N_28324);
nor UO_2916 (O_2916,N_28230,N_27552);
and UO_2917 (O_2917,N_27110,N_29430);
or UO_2918 (O_2918,N_26242,N_29209);
nor UO_2919 (O_2919,N_25370,N_27051);
or UO_2920 (O_2920,N_26185,N_25615);
nand UO_2921 (O_2921,N_25969,N_27206);
nand UO_2922 (O_2922,N_25237,N_26874);
nor UO_2923 (O_2923,N_26641,N_25275);
nor UO_2924 (O_2924,N_26856,N_28386);
and UO_2925 (O_2925,N_27802,N_26158);
and UO_2926 (O_2926,N_27885,N_28817);
nor UO_2927 (O_2927,N_27984,N_26789);
and UO_2928 (O_2928,N_28115,N_28216);
and UO_2929 (O_2929,N_27439,N_26605);
xnor UO_2930 (O_2930,N_28405,N_27836);
nor UO_2931 (O_2931,N_26057,N_28699);
xor UO_2932 (O_2932,N_26211,N_28653);
or UO_2933 (O_2933,N_26736,N_29428);
nor UO_2934 (O_2934,N_28560,N_26889);
and UO_2935 (O_2935,N_27455,N_25270);
xor UO_2936 (O_2936,N_27744,N_29700);
nand UO_2937 (O_2937,N_29402,N_26839);
nand UO_2938 (O_2938,N_28426,N_27551);
xnor UO_2939 (O_2939,N_25066,N_29724);
or UO_2940 (O_2940,N_27383,N_26414);
or UO_2941 (O_2941,N_25238,N_29778);
and UO_2942 (O_2942,N_28740,N_25316);
xnor UO_2943 (O_2943,N_28125,N_28585);
xnor UO_2944 (O_2944,N_29315,N_26870);
xor UO_2945 (O_2945,N_28108,N_26345);
and UO_2946 (O_2946,N_26709,N_25463);
nand UO_2947 (O_2947,N_25030,N_29424);
or UO_2948 (O_2948,N_28124,N_26732);
nor UO_2949 (O_2949,N_26060,N_27358);
and UO_2950 (O_2950,N_27486,N_26571);
and UO_2951 (O_2951,N_28410,N_27368);
xor UO_2952 (O_2952,N_28305,N_28948);
xor UO_2953 (O_2953,N_29282,N_28244);
and UO_2954 (O_2954,N_29527,N_27921);
nor UO_2955 (O_2955,N_28563,N_26850);
and UO_2956 (O_2956,N_28218,N_29341);
nor UO_2957 (O_2957,N_29270,N_29744);
or UO_2958 (O_2958,N_25523,N_29132);
nand UO_2959 (O_2959,N_27021,N_27141);
nor UO_2960 (O_2960,N_27239,N_27597);
and UO_2961 (O_2961,N_28153,N_26753);
xnor UO_2962 (O_2962,N_27449,N_29500);
xor UO_2963 (O_2963,N_25058,N_26203);
or UO_2964 (O_2964,N_26849,N_25674);
or UO_2965 (O_2965,N_25796,N_28212);
nand UO_2966 (O_2966,N_25686,N_28081);
xnor UO_2967 (O_2967,N_26977,N_29129);
or UO_2968 (O_2968,N_27194,N_26725);
and UO_2969 (O_2969,N_26894,N_27014);
or UO_2970 (O_2970,N_26867,N_29617);
nand UO_2971 (O_2971,N_26551,N_28964);
and UO_2972 (O_2972,N_28952,N_25147);
nand UO_2973 (O_2973,N_27937,N_29640);
or UO_2974 (O_2974,N_27439,N_29762);
xor UO_2975 (O_2975,N_27948,N_26602);
nand UO_2976 (O_2976,N_25168,N_29013);
xor UO_2977 (O_2977,N_26245,N_28333);
or UO_2978 (O_2978,N_26966,N_28295);
xnor UO_2979 (O_2979,N_25537,N_26630);
and UO_2980 (O_2980,N_29207,N_29174);
and UO_2981 (O_2981,N_26984,N_28181);
nor UO_2982 (O_2982,N_27963,N_26462);
xnor UO_2983 (O_2983,N_25948,N_25178);
xnor UO_2984 (O_2984,N_28875,N_26119);
nor UO_2985 (O_2985,N_29968,N_29089);
or UO_2986 (O_2986,N_29026,N_27145);
nor UO_2987 (O_2987,N_25939,N_29249);
nand UO_2988 (O_2988,N_27331,N_28469);
or UO_2989 (O_2989,N_28395,N_25343);
nand UO_2990 (O_2990,N_29819,N_26438);
xor UO_2991 (O_2991,N_28656,N_26736);
nor UO_2992 (O_2992,N_29705,N_28300);
and UO_2993 (O_2993,N_28590,N_25940);
or UO_2994 (O_2994,N_29485,N_25987);
nor UO_2995 (O_2995,N_25106,N_26281);
or UO_2996 (O_2996,N_26638,N_28857);
xnor UO_2997 (O_2997,N_29302,N_25633);
xnor UO_2998 (O_2998,N_29246,N_26796);
nor UO_2999 (O_2999,N_27296,N_27596);
xnor UO_3000 (O_3000,N_29803,N_25419);
or UO_3001 (O_3001,N_26787,N_28137);
nor UO_3002 (O_3002,N_28349,N_26755);
nor UO_3003 (O_3003,N_28101,N_25478);
xnor UO_3004 (O_3004,N_25248,N_27022);
or UO_3005 (O_3005,N_28404,N_26313);
or UO_3006 (O_3006,N_27826,N_25705);
nor UO_3007 (O_3007,N_26820,N_27154);
nand UO_3008 (O_3008,N_29538,N_26892);
nor UO_3009 (O_3009,N_29144,N_29360);
or UO_3010 (O_3010,N_28323,N_26182);
and UO_3011 (O_3011,N_28982,N_27211);
xor UO_3012 (O_3012,N_26314,N_27437);
and UO_3013 (O_3013,N_29707,N_28108);
or UO_3014 (O_3014,N_27845,N_25621);
nor UO_3015 (O_3015,N_25294,N_29177);
xor UO_3016 (O_3016,N_25637,N_28236);
xor UO_3017 (O_3017,N_27779,N_28596);
nand UO_3018 (O_3018,N_27703,N_29366);
nand UO_3019 (O_3019,N_28998,N_28458);
xor UO_3020 (O_3020,N_26231,N_27927);
xor UO_3021 (O_3021,N_28255,N_28409);
nand UO_3022 (O_3022,N_29828,N_28027);
nand UO_3023 (O_3023,N_25313,N_26000);
and UO_3024 (O_3024,N_27789,N_29928);
nand UO_3025 (O_3025,N_25091,N_26477);
and UO_3026 (O_3026,N_25111,N_28253);
nor UO_3027 (O_3027,N_26511,N_28751);
and UO_3028 (O_3028,N_29763,N_26621);
nand UO_3029 (O_3029,N_26173,N_25855);
xnor UO_3030 (O_3030,N_27429,N_28386);
xor UO_3031 (O_3031,N_29942,N_26425);
nor UO_3032 (O_3032,N_26885,N_26072);
or UO_3033 (O_3033,N_27021,N_27366);
nor UO_3034 (O_3034,N_28869,N_28135);
nand UO_3035 (O_3035,N_26588,N_29987);
nand UO_3036 (O_3036,N_27807,N_29823);
nor UO_3037 (O_3037,N_27951,N_28859);
nand UO_3038 (O_3038,N_26282,N_25527);
and UO_3039 (O_3039,N_27133,N_27798);
and UO_3040 (O_3040,N_27915,N_25000);
xor UO_3041 (O_3041,N_25857,N_29215);
and UO_3042 (O_3042,N_27510,N_29866);
or UO_3043 (O_3043,N_28690,N_29553);
nand UO_3044 (O_3044,N_26394,N_25427);
xnor UO_3045 (O_3045,N_25326,N_26115);
xnor UO_3046 (O_3046,N_29403,N_29205);
and UO_3047 (O_3047,N_27526,N_28749);
xnor UO_3048 (O_3048,N_28827,N_27638);
xor UO_3049 (O_3049,N_26675,N_28529);
nand UO_3050 (O_3050,N_29011,N_25029);
and UO_3051 (O_3051,N_25471,N_28680);
and UO_3052 (O_3052,N_29826,N_29115);
xnor UO_3053 (O_3053,N_28920,N_28873);
nor UO_3054 (O_3054,N_25800,N_26034);
or UO_3055 (O_3055,N_28519,N_27960);
nand UO_3056 (O_3056,N_27103,N_28655);
nor UO_3057 (O_3057,N_26226,N_26288);
or UO_3058 (O_3058,N_28639,N_27059);
nand UO_3059 (O_3059,N_28833,N_27777);
and UO_3060 (O_3060,N_25293,N_26299);
or UO_3061 (O_3061,N_29031,N_27415);
nand UO_3062 (O_3062,N_25236,N_28291);
nor UO_3063 (O_3063,N_25869,N_29971);
and UO_3064 (O_3064,N_28613,N_29846);
or UO_3065 (O_3065,N_28518,N_25872);
nor UO_3066 (O_3066,N_29307,N_28504);
nor UO_3067 (O_3067,N_25964,N_27080);
and UO_3068 (O_3068,N_28714,N_25947);
nand UO_3069 (O_3069,N_26050,N_26301);
nand UO_3070 (O_3070,N_26291,N_28912);
nand UO_3071 (O_3071,N_27851,N_29056);
or UO_3072 (O_3072,N_26449,N_26102);
nor UO_3073 (O_3073,N_26729,N_28486);
or UO_3074 (O_3074,N_28971,N_28579);
nand UO_3075 (O_3075,N_28875,N_28247);
nand UO_3076 (O_3076,N_28980,N_26999);
or UO_3077 (O_3077,N_27642,N_26018);
or UO_3078 (O_3078,N_26065,N_26942);
and UO_3079 (O_3079,N_27290,N_25882);
and UO_3080 (O_3080,N_28284,N_26794);
or UO_3081 (O_3081,N_25312,N_26684);
or UO_3082 (O_3082,N_28449,N_29771);
nand UO_3083 (O_3083,N_25796,N_27217);
xor UO_3084 (O_3084,N_28290,N_26551);
nor UO_3085 (O_3085,N_28588,N_27085);
xor UO_3086 (O_3086,N_29473,N_28919);
or UO_3087 (O_3087,N_29141,N_29812);
nor UO_3088 (O_3088,N_26678,N_27493);
nor UO_3089 (O_3089,N_28273,N_28647);
nor UO_3090 (O_3090,N_27828,N_27201);
nand UO_3091 (O_3091,N_26402,N_29377);
nor UO_3092 (O_3092,N_29602,N_25522);
nand UO_3093 (O_3093,N_27334,N_27723);
or UO_3094 (O_3094,N_29080,N_28708);
xor UO_3095 (O_3095,N_28610,N_27541);
nand UO_3096 (O_3096,N_29975,N_25266);
nor UO_3097 (O_3097,N_26888,N_27555);
xor UO_3098 (O_3098,N_28351,N_29535);
or UO_3099 (O_3099,N_26837,N_29788);
and UO_3100 (O_3100,N_25755,N_25473);
xnor UO_3101 (O_3101,N_26623,N_26810);
nor UO_3102 (O_3102,N_28707,N_27157);
nor UO_3103 (O_3103,N_26337,N_27478);
nand UO_3104 (O_3104,N_27131,N_25864);
and UO_3105 (O_3105,N_29482,N_29226);
nor UO_3106 (O_3106,N_27772,N_27753);
and UO_3107 (O_3107,N_27756,N_29701);
and UO_3108 (O_3108,N_25875,N_26708);
nand UO_3109 (O_3109,N_28025,N_29683);
nor UO_3110 (O_3110,N_27111,N_28267);
nand UO_3111 (O_3111,N_27512,N_29479);
xor UO_3112 (O_3112,N_28058,N_28916);
nand UO_3113 (O_3113,N_28653,N_28649);
xnor UO_3114 (O_3114,N_28798,N_29546);
xnor UO_3115 (O_3115,N_27397,N_25323);
or UO_3116 (O_3116,N_25307,N_27665);
and UO_3117 (O_3117,N_28927,N_25567);
or UO_3118 (O_3118,N_27914,N_29573);
nand UO_3119 (O_3119,N_28689,N_28240);
or UO_3120 (O_3120,N_28625,N_25305);
or UO_3121 (O_3121,N_29784,N_25267);
nand UO_3122 (O_3122,N_28638,N_28691);
or UO_3123 (O_3123,N_29605,N_29892);
nand UO_3124 (O_3124,N_26257,N_27277);
xnor UO_3125 (O_3125,N_29103,N_25349);
xor UO_3126 (O_3126,N_25302,N_28023);
or UO_3127 (O_3127,N_25109,N_28283);
xor UO_3128 (O_3128,N_28797,N_29924);
xor UO_3129 (O_3129,N_27441,N_29788);
nor UO_3130 (O_3130,N_28646,N_28563);
nor UO_3131 (O_3131,N_28730,N_27458);
or UO_3132 (O_3132,N_27616,N_29643);
nor UO_3133 (O_3133,N_28548,N_28185);
xnor UO_3134 (O_3134,N_29267,N_27845);
or UO_3135 (O_3135,N_26906,N_29236);
xnor UO_3136 (O_3136,N_29662,N_25415);
nand UO_3137 (O_3137,N_25999,N_25259);
nor UO_3138 (O_3138,N_25622,N_26225);
or UO_3139 (O_3139,N_28874,N_29824);
nor UO_3140 (O_3140,N_27042,N_25959);
and UO_3141 (O_3141,N_26625,N_25008);
xnor UO_3142 (O_3142,N_28688,N_29312);
or UO_3143 (O_3143,N_27397,N_26727);
nand UO_3144 (O_3144,N_26058,N_28098);
xnor UO_3145 (O_3145,N_25591,N_28207);
and UO_3146 (O_3146,N_29299,N_29086);
xor UO_3147 (O_3147,N_27330,N_28706);
xor UO_3148 (O_3148,N_28431,N_27122);
and UO_3149 (O_3149,N_27483,N_29002);
and UO_3150 (O_3150,N_28123,N_26427);
nand UO_3151 (O_3151,N_25524,N_26458);
nand UO_3152 (O_3152,N_26798,N_29791);
or UO_3153 (O_3153,N_27539,N_25448);
nand UO_3154 (O_3154,N_28570,N_29056);
nand UO_3155 (O_3155,N_27907,N_26251);
nor UO_3156 (O_3156,N_28825,N_25256);
xnor UO_3157 (O_3157,N_28319,N_29447);
nor UO_3158 (O_3158,N_26695,N_26061);
or UO_3159 (O_3159,N_27298,N_28201);
nor UO_3160 (O_3160,N_28121,N_28514);
nand UO_3161 (O_3161,N_29134,N_26386);
xor UO_3162 (O_3162,N_29440,N_28418);
and UO_3163 (O_3163,N_27875,N_26302);
nor UO_3164 (O_3164,N_26154,N_25072);
nor UO_3165 (O_3165,N_29006,N_29617);
nor UO_3166 (O_3166,N_25182,N_28789);
or UO_3167 (O_3167,N_28783,N_27591);
xor UO_3168 (O_3168,N_29984,N_25586);
nand UO_3169 (O_3169,N_25784,N_25210);
nand UO_3170 (O_3170,N_27542,N_29727);
nor UO_3171 (O_3171,N_29216,N_25324);
nor UO_3172 (O_3172,N_25094,N_27551);
or UO_3173 (O_3173,N_26079,N_29477);
xor UO_3174 (O_3174,N_28459,N_26006);
or UO_3175 (O_3175,N_28453,N_28302);
xor UO_3176 (O_3176,N_27402,N_27253);
nor UO_3177 (O_3177,N_29962,N_27048);
nand UO_3178 (O_3178,N_28339,N_27715);
nor UO_3179 (O_3179,N_28394,N_27097);
xnor UO_3180 (O_3180,N_28406,N_27780);
or UO_3181 (O_3181,N_27908,N_29566);
xor UO_3182 (O_3182,N_28275,N_27566);
xor UO_3183 (O_3183,N_26208,N_25207);
xor UO_3184 (O_3184,N_27613,N_25157);
and UO_3185 (O_3185,N_29063,N_27576);
xnor UO_3186 (O_3186,N_27417,N_26735);
nand UO_3187 (O_3187,N_28004,N_29077);
xnor UO_3188 (O_3188,N_29522,N_28868);
or UO_3189 (O_3189,N_27061,N_28023);
nand UO_3190 (O_3190,N_26901,N_29638);
xor UO_3191 (O_3191,N_26306,N_29881);
and UO_3192 (O_3192,N_26814,N_25840);
nand UO_3193 (O_3193,N_26326,N_27599);
or UO_3194 (O_3194,N_26819,N_27682);
nand UO_3195 (O_3195,N_26379,N_26501);
nand UO_3196 (O_3196,N_27240,N_29360);
and UO_3197 (O_3197,N_28971,N_26479);
nor UO_3198 (O_3198,N_26406,N_27657);
or UO_3199 (O_3199,N_28856,N_26650);
nand UO_3200 (O_3200,N_27665,N_28112);
nand UO_3201 (O_3201,N_25024,N_27765);
nor UO_3202 (O_3202,N_27988,N_25748);
nor UO_3203 (O_3203,N_27464,N_29345);
xnor UO_3204 (O_3204,N_29778,N_27717);
nor UO_3205 (O_3205,N_26644,N_26562);
and UO_3206 (O_3206,N_29539,N_29074);
nand UO_3207 (O_3207,N_25109,N_29506);
and UO_3208 (O_3208,N_28616,N_25032);
or UO_3209 (O_3209,N_29589,N_29470);
xnor UO_3210 (O_3210,N_27595,N_27710);
or UO_3211 (O_3211,N_27591,N_25176);
or UO_3212 (O_3212,N_25555,N_28082);
or UO_3213 (O_3213,N_25096,N_28907);
nand UO_3214 (O_3214,N_28979,N_28081);
xnor UO_3215 (O_3215,N_26624,N_26318);
xnor UO_3216 (O_3216,N_27814,N_29800);
and UO_3217 (O_3217,N_25902,N_26623);
nor UO_3218 (O_3218,N_27575,N_29531);
nor UO_3219 (O_3219,N_29306,N_25617);
nor UO_3220 (O_3220,N_29313,N_27823);
nor UO_3221 (O_3221,N_25066,N_28352);
or UO_3222 (O_3222,N_26848,N_26900);
nor UO_3223 (O_3223,N_26737,N_25218);
and UO_3224 (O_3224,N_28944,N_25671);
or UO_3225 (O_3225,N_29156,N_25316);
xnor UO_3226 (O_3226,N_29064,N_29008);
and UO_3227 (O_3227,N_26159,N_29034);
xor UO_3228 (O_3228,N_27395,N_27085);
nor UO_3229 (O_3229,N_26810,N_27899);
or UO_3230 (O_3230,N_28590,N_26894);
nor UO_3231 (O_3231,N_26765,N_28083);
xor UO_3232 (O_3232,N_26138,N_29969);
nor UO_3233 (O_3233,N_25414,N_27658);
and UO_3234 (O_3234,N_29814,N_26458);
nor UO_3235 (O_3235,N_27379,N_25707);
or UO_3236 (O_3236,N_28356,N_28379);
or UO_3237 (O_3237,N_26679,N_26156);
nor UO_3238 (O_3238,N_28171,N_25727);
or UO_3239 (O_3239,N_26674,N_26951);
nor UO_3240 (O_3240,N_27554,N_29128);
nand UO_3241 (O_3241,N_28569,N_28214);
xnor UO_3242 (O_3242,N_28790,N_26514);
nor UO_3243 (O_3243,N_28914,N_26719);
nand UO_3244 (O_3244,N_29244,N_27371);
or UO_3245 (O_3245,N_26335,N_28220);
or UO_3246 (O_3246,N_25854,N_28742);
or UO_3247 (O_3247,N_28337,N_28425);
nor UO_3248 (O_3248,N_25869,N_25248);
or UO_3249 (O_3249,N_26967,N_26988);
nand UO_3250 (O_3250,N_27365,N_25263);
nand UO_3251 (O_3251,N_29946,N_26962);
nand UO_3252 (O_3252,N_28899,N_29622);
or UO_3253 (O_3253,N_25355,N_29092);
or UO_3254 (O_3254,N_27319,N_27907);
nand UO_3255 (O_3255,N_26743,N_28840);
nand UO_3256 (O_3256,N_29489,N_29208);
nor UO_3257 (O_3257,N_28884,N_28298);
nor UO_3258 (O_3258,N_27655,N_29496);
or UO_3259 (O_3259,N_25103,N_29912);
and UO_3260 (O_3260,N_26380,N_26454);
nand UO_3261 (O_3261,N_26520,N_26073);
and UO_3262 (O_3262,N_25006,N_29467);
xnor UO_3263 (O_3263,N_27706,N_26426);
nand UO_3264 (O_3264,N_26880,N_28996);
and UO_3265 (O_3265,N_29697,N_29354);
nand UO_3266 (O_3266,N_26266,N_26259);
or UO_3267 (O_3267,N_27119,N_27049);
or UO_3268 (O_3268,N_28315,N_28954);
or UO_3269 (O_3269,N_25008,N_28175);
and UO_3270 (O_3270,N_27611,N_26782);
nor UO_3271 (O_3271,N_25570,N_26822);
or UO_3272 (O_3272,N_27366,N_29930);
nor UO_3273 (O_3273,N_26769,N_25783);
nor UO_3274 (O_3274,N_28232,N_29156);
nor UO_3275 (O_3275,N_29997,N_28335);
nand UO_3276 (O_3276,N_28912,N_27212);
xnor UO_3277 (O_3277,N_25519,N_27943);
xnor UO_3278 (O_3278,N_28291,N_26929);
xor UO_3279 (O_3279,N_28640,N_25471);
nand UO_3280 (O_3280,N_27007,N_25056);
nand UO_3281 (O_3281,N_27611,N_26687);
or UO_3282 (O_3282,N_26739,N_26478);
and UO_3283 (O_3283,N_26369,N_26250);
and UO_3284 (O_3284,N_26060,N_25892);
nor UO_3285 (O_3285,N_25382,N_25728);
nor UO_3286 (O_3286,N_26864,N_29378);
or UO_3287 (O_3287,N_25240,N_29250);
and UO_3288 (O_3288,N_25146,N_26390);
or UO_3289 (O_3289,N_28636,N_26610);
or UO_3290 (O_3290,N_27283,N_25410);
nor UO_3291 (O_3291,N_27393,N_25246);
nor UO_3292 (O_3292,N_26182,N_29656);
xnor UO_3293 (O_3293,N_29382,N_26640);
nand UO_3294 (O_3294,N_26336,N_26126);
xnor UO_3295 (O_3295,N_26125,N_29357);
or UO_3296 (O_3296,N_26401,N_25856);
or UO_3297 (O_3297,N_28272,N_29983);
and UO_3298 (O_3298,N_28666,N_25833);
xor UO_3299 (O_3299,N_25929,N_28574);
nand UO_3300 (O_3300,N_26385,N_26238);
and UO_3301 (O_3301,N_28339,N_29975);
or UO_3302 (O_3302,N_26956,N_26425);
nor UO_3303 (O_3303,N_25163,N_26432);
or UO_3304 (O_3304,N_27383,N_27147);
xor UO_3305 (O_3305,N_25177,N_28836);
or UO_3306 (O_3306,N_27637,N_28656);
nor UO_3307 (O_3307,N_27985,N_29723);
nand UO_3308 (O_3308,N_26966,N_28468);
nand UO_3309 (O_3309,N_26517,N_28375);
and UO_3310 (O_3310,N_28194,N_27725);
or UO_3311 (O_3311,N_27303,N_28077);
nor UO_3312 (O_3312,N_29851,N_29043);
nand UO_3313 (O_3313,N_26750,N_27958);
nor UO_3314 (O_3314,N_27985,N_26768);
and UO_3315 (O_3315,N_29092,N_27304);
xor UO_3316 (O_3316,N_27546,N_25232);
xnor UO_3317 (O_3317,N_26645,N_27896);
or UO_3318 (O_3318,N_29565,N_26430);
nor UO_3319 (O_3319,N_29413,N_29736);
nand UO_3320 (O_3320,N_25664,N_25385);
nand UO_3321 (O_3321,N_26606,N_26852);
or UO_3322 (O_3322,N_27268,N_27019);
or UO_3323 (O_3323,N_28190,N_27341);
xnor UO_3324 (O_3324,N_26115,N_25948);
nand UO_3325 (O_3325,N_29140,N_28371);
nand UO_3326 (O_3326,N_26282,N_29317);
xnor UO_3327 (O_3327,N_29298,N_27146);
or UO_3328 (O_3328,N_29270,N_26227);
or UO_3329 (O_3329,N_27953,N_27565);
nand UO_3330 (O_3330,N_27682,N_27857);
and UO_3331 (O_3331,N_25255,N_26192);
or UO_3332 (O_3332,N_28311,N_26516);
or UO_3333 (O_3333,N_26989,N_28256);
xor UO_3334 (O_3334,N_29632,N_25779);
nand UO_3335 (O_3335,N_25440,N_28566);
or UO_3336 (O_3336,N_25359,N_25139);
nor UO_3337 (O_3337,N_26005,N_29182);
xnor UO_3338 (O_3338,N_29569,N_27670);
and UO_3339 (O_3339,N_29866,N_25219);
or UO_3340 (O_3340,N_29989,N_29392);
nor UO_3341 (O_3341,N_25988,N_26580);
and UO_3342 (O_3342,N_28166,N_27244);
xnor UO_3343 (O_3343,N_27454,N_25677);
nand UO_3344 (O_3344,N_26927,N_28973);
xnor UO_3345 (O_3345,N_28483,N_26218);
nor UO_3346 (O_3346,N_26640,N_29636);
and UO_3347 (O_3347,N_26523,N_27980);
nor UO_3348 (O_3348,N_26380,N_25368);
xnor UO_3349 (O_3349,N_26622,N_28186);
and UO_3350 (O_3350,N_26056,N_28038);
or UO_3351 (O_3351,N_27234,N_27977);
xnor UO_3352 (O_3352,N_25690,N_27745);
nor UO_3353 (O_3353,N_26227,N_26139);
nand UO_3354 (O_3354,N_26588,N_26945);
nand UO_3355 (O_3355,N_25531,N_26010);
xnor UO_3356 (O_3356,N_28136,N_28497);
or UO_3357 (O_3357,N_25197,N_29975);
or UO_3358 (O_3358,N_29243,N_28857);
and UO_3359 (O_3359,N_25949,N_28988);
and UO_3360 (O_3360,N_27119,N_26187);
nand UO_3361 (O_3361,N_29873,N_28357);
xor UO_3362 (O_3362,N_25323,N_25273);
and UO_3363 (O_3363,N_27137,N_26514);
nand UO_3364 (O_3364,N_28516,N_25619);
nor UO_3365 (O_3365,N_27578,N_25259);
or UO_3366 (O_3366,N_28600,N_28627);
nor UO_3367 (O_3367,N_26923,N_26675);
nand UO_3368 (O_3368,N_27965,N_26377);
or UO_3369 (O_3369,N_28509,N_25175);
or UO_3370 (O_3370,N_28213,N_26109);
nor UO_3371 (O_3371,N_27698,N_29905);
nor UO_3372 (O_3372,N_28248,N_28346);
and UO_3373 (O_3373,N_27502,N_25262);
or UO_3374 (O_3374,N_25079,N_26361);
xor UO_3375 (O_3375,N_28929,N_29347);
or UO_3376 (O_3376,N_28214,N_27270);
nand UO_3377 (O_3377,N_26520,N_28174);
nand UO_3378 (O_3378,N_28763,N_28435);
nor UO_3379 (O_3379,N_29109,N_25205);
nor UO_3380 (O_3380,N_27639,N_29625);
and UO_3381 (O_3381,N_25439,N_27852);
nand UO_3382 (O_3382,N_26793,N_26651);
xor UO_3383 (O_3383,N_26926,N_28581);
nor UO_3384 (O_3384,N_27632,N_29697);
nand UO_3385 (O_3385,N_29260,N_27796);
or UO_3386 (O_3386,N_27956,N_26008);
nor UO_3387 (O_3387,N_27162,N_25716);
nor UO_3388 (O_3388,N_25576,N_25000);
and UO_3389 (O_3389,N_29303,N_29537);
nor UO_3390 (O_3390,N_26799,N_25414);
and UO_3391 (O_3391,N_25967,N_28663);
nor UO_3392 (O_3392,N_29150,N_26206);
and UO_3393 (O_3393,N_25692,N_25862);
and UO_3394 (O_3394,N_26029,N_28537);
nand UO_3395 (O_3395,N_29467,N_29231);
nor UO_3396 (O_3396,N_25180,N_29812);
nor UO_3397 (O_3397,N_29566,N_25918);
xnor UO_3398 (O_3398,N_28577,N_28315);
xnor UO_3399 (O_3399,N_25579,N_29522);
xnor UO_3400 (O_3400,N_27495,N_25163);
nor UO_3401 (O_3401,N_25090,N_26168);
xnor UO_3402 (O_3402,N_26805,N_25843);
nor UO_3403 (O_3403,N_28760,N_26753);
or UO_3404 (O_3404,N_26772,N_29583);
nand UO_3405 (O_3405,N_27167,N_25694);
nand UO_3406 (O_3406,N_26759,N_28566);
xnor UO_3407 (O_3407,N_27836,N_28285);
nor UO_3408 (O_3408,N_28847,N_27827);
xnor UO_3409 (O_3409,N_25207,N_29107);
and UO_3410 (O_3410,N_26978,N_27109);
nand UO_3411 (O_3411,N_26142,N_28253);
or UO_3412 (O_3412,N_27117,N_28762);
and UO_3413 (O_3413,N_29857,N_27119);
and UO_3414 (O_3414,N_29657,N_25721);
nor UO_3415 (O_3415,N_27595,N_28037);
and UO_3416 (O_3416,N_27774,N_27006);
or UO_3417 (O_3417,N_25709,N_26254);
and UO_3418 (O_3418,N_26628,N_25691);
xor UO_3419 (O_3419,N_27484,N_27641);
xor UO_3420 (O_3420,N_29989,N_28972);
xnor UO_3421 (O_3421,N_25093,N_27851);
and UO_3422 (O_3422,N_29485,N_26482);
nand UO_3423 (O_3423,N_25277,N_28311);
and UO_3424 (O_3424,N_28891,N_29725);
nor UO_3425 (O_3425,N_28190,N_25957);
nand UO_3426 (O_3426,N_29973,N_28601);
and UO_3427 (O_3427,N_28694,N_27419);
or UO_3428 (O_3428,N_27849,N_28520);
nor UO_3429 (O_3429,N_29546,N_26520);
nand UO_3430 (O_3430,N_26394,N_25981);
and UO_3431 (O_3431,N_25952,N_27633);
nand UO_3432 (O_3432,N_25625,N_25473);
nor UO_3433 (O_3433,N_26437,N_25477);
nand UO_3434 (O_3434,N_25233,N_26222);
nor UO_3435 (O_3435,N_26042,N_29053);
nand UO_3436 (O_3436,N_25958,N_29071);
nand UO_3437 (O_3437,N_29281,N_27945);
and UO_3438 (O_3438,N_25986,N_29251);
or UO_3439 (O_3439,N_29343,N_25667);
and UO_3440 (O_3440,N_26866,N_26223);
or UO_3441 (O_3441,N_27789,N_26190);
nor UO_3442 (O_3442,N_29144,N_26365);
nand UO_3443 (O_3443,N_25416,N_26086);
or UO_3444 (O_3444,N_29947,N_26462);
nand UO_3445 (O_3445,N_25957,N_27291);
nor UO_3446 (O_3446,N_27984,N_25181);
xor UO_3447 (O_3447,N_29637,N_29229);
and UO_3448 (O_3448,N_25101,N_27815);
and UO_3449 (O_3449,N_28256,N_26785);
or UO_3450 (O_3450,N_26735,N_26376);
nand UO_3451 (O_3451,N_29427,N_28795);
nor UO_3452 (O_3452,N_26972,N_27783);
nor UO_3453 (O_3453,N_29673,N_28809);
or UO_3454 (O_3454,N_25711,N_27371);
nand UO_3455 (O_3455,N_28932,N_28192);
nor UO_3456 (O_3456,N_27111,N_26988);
nand UO_3457 (O_3457,N_25533,N_27162);
nand UO_3458 (O_3458,N_25320,N_29768);
and UO_3459 (O_3459,N_25482,N_29580);
nand UO_3460 (O_3460,N_27825,N_28400);
xor UO_3461 (O_3461,N_25984,N_28294);
xor UO_3462 (O_3462,N_29310,N_25859);
nand UO_3463 (O_3463,N_25724,N_26476);
or UO_3464 (O_3464,N_26992,N_28294);
nand UO_3465 (O_3465,N_28972,N_29699);
nor UO_3466 (O_3466,N_28128,N_29833);
or UO_3467 (O_3467,N_27528,N_28282);
nand UO_3468 (O_3468,N_26582,N_27637);
nor UO_3469 (O_3469,N_28735,N_25070);
nor UO_3470 (O_3470,N_29065,N_28243);
nand UO_3471 (O_3471,N_27583,N_26402);
nor UO_3472 (O_3472,N_27162,N_27660);
and UO_3473 (O_3473,N_25883,N_29521);
or UO_3474 (O_3474,N_28030,N_26710);
nand UO_3475 (O_3475,N_25576,N_26415);
xnor UO_3476 (O_3476,N_29621,N_26390);
and UO_3477 (O_3477,N_28349,N_27626);
or UO_3478 (O_3478,N_29093,N_27909);
nand UO_3479 (O_3479,N_29179,N_26236);
nand UO_3480 (O_3480,N_27937,N_27960);
or UO_3481 (O_3481,N_28936,N_29664);
or UO_3482 (O_3482,N_29054,N_26656);
xor UO_3483 (O_3483,N_28398,N_26454);
xor UO_3484 (O_3484,N_25595,N_25526);
and UO_3485 (O_3485,N_26850,N_29496);
nand UO_3486 (O_3486,N_29361,N_26759);
nor UO_3487 (O_3487,N_29022,N_26470);
and UO_3488 (O_3488,N_28786,N_29347);
nor UO_3489 (O_3489,N_26102,N_28475);
and UO_3490 (O_3490,N_29033,N_29249);
or UO_3491 (O_3491,N_25266,N_28443);
nand UO_3492 (O_3492,N_29899,N_25922);
or UO_3493 (O_3493,N_28908,N_25638);
and UO_3494 (O_3494,N_27809,N_25686);
nand UO_3495 (O_3495,N_25117,N_27223);
or UO_3496 (O_3496,N_27083,N_26320);
nand UO_3497 (O_3497,N_28368,N_28956);
or UO_3498 (O_3498,N_28703,N_28750);
or UO_3499 (O_3499,N_25948,N_27376);
endmodule