module basic_2500_25000_3000_8_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_894,In_1033);
and U1 (N_1,In_718,In_965);
nor U2 (N_2,In_873,In_1218);
or U3 (N_3,In_809,In_1562);
nor U4 (N_4,In_1829,In_790);
nor U5 (N_5,In_1843,In_1666);
or U6 (N_6,In_282,In_1793);
and U7 (N_7,In_1437,In_814);
and U8 (N_8,In_2271,In_1587);
xnor U9 (N_9,In_1897,In_1947);
nand U10 (N_10,In_594,In_767);
nand U11 (N_11,In_2317,In_1154);
or U12 (N_12,In_373,In_748);
xor U13 (N_13,In_128,In_1151);
xor U14 (N_14,In_380,In_1962);
nand U15 (N_15,In_1588,In_242);
nor U16 (N_16,In_2399,In_1935);
and U17 (N_17,In_1410,In_1697);
nand U18 (N_18,In_110,In_835);
or U19 (N_19,In_354,In_688);
or U20 (N_20,In_1084,In_243);
or U21 (N_21,In_1135,In_1176);
xor U22 (N_22,In_685,In_2262);
xor U23 (N_23,In_761,In_1488);
and U24 (N_24,In_1535,In_1003);
nor U25 (N_25,In_609,In_94);
and U26 (N_26,In_165,In_1435);
xnor U27 (N_27,In_1441,In_105);
nand U28 (N_28,In_41,In_1508);
nor U29 (N_29,In_2015,In_1881);
xor U30 (N_30,In_987,In_1018);
and U31 (N_31,In_285,In_1740);
or U32 (N_32,In_513,In_1335);
nor U33 (N_33,In_1326,In_113);
and U34 (N_34,In_2246,In_1858);
nand U35 (N_35,In_910,In_645);
nand U36 (N_36,In_531,In_2441);
xor U37 (N_37,In_1366,In_1266);
xor U38 (N_38,In_430,In_786);
nand U39 (N_39,In_2190,In_481);
or U40 (N_40,In_367,In_615);
and U41 (N_41,In_565,In_2429);
and U42 (N_42,In_2493,In_184);
and U43 (N_43,In_997,In_1049);
and U44 (N_44,In_2151,In_1857);
xnor U45 (N_45,In_358,In_439);
xnor U46 (N_46,In_1316,In_706);
nand U47 (N_47,In_1701,In_1452);
nand U48 (N_48,In_1870,In_981);
xnor U49 (N_49,In_507,In_2153);
nor U50 (N_50,In_2230,In_6);
and U51 (N_51,In_630,In_2118);
xnor U52 (N_52,In_1998,In_344);
xnor U53 (N_53,In_172,In_2411);
or U54 (N_54,In_1337,In_231);
nor U55 (N_55,In_823,In_723);
nor U56 (N_56,In_67,In_1856);
and U57 (N_57,In_2165,In_2098);
or U58 (N_58,In_1372,In_2415);
nand U59 (N_59,In_224,In_148);
or U60 (N_60,In_1346,In_1997);
xor U61 (N_61,In_500,In_551);
nor U62 (N_62,In_625,In_549);
or U63 (N_63,In_730,In_1627);
xnor U64 (N_64,In_1411,In_1388);
nand U65 (N_65,In_784,In_1582);
xnor U66 (N_66,In_2345,In_222);
and U67 (N_67,In_2244,In_794);
xor U68 (N_68,In_2397,In_752);
and U69 (N_69,In_1097,In_2203);
and U70 (N_70,In_80,In_2075);
or U71 (N_71,In_785,In_1663);
xor U72 (N_72,In_1568,In_2319);
or U73 (N_73,In_2475,In_632);
nor U74 (N_74,In_2217,In_432);
nand U75 (N_75,In_872,In_484);
xor U76 (N_76,In_1132,In_1912);
xor U77 (N_77,In_808,In_1470);
or U78 (N_78,In_1491,In_1436);
nor U79 (N_79,In_735,In_475);
xor U80 (N_80,In_174,In_1404);
nand U81 (N_81,In_1817,In_250);
nor U82 (N_82,In_1550,In_750);
xor U83 (N_83,In_1516,In_1930);
or U84 (N_84,In_686,In_1636);
xor U85 (N_85,In_877,In_1290);
nor U86 (N_86,In_1024,In_2160);
nand U87 (N_87,In_1548,In_1527);
or U88 (N_88,In_406,In_300);
or U89 (N_89,In_1333,In_419);
or U90 (N_90,In_1917,In_661);
or U91 (N_91,In_1838,In_364);
nor U92 (N_92,In_1732,In_2081);
or U93 (N_93,In_1791,In_47);
nand U94 (N_94,In_332,In_1685);
or U95 (N_95,In_1541,In_1932);
xnor U96 (N_96,In_137,In_399);
or U97 (N_97,In_2329,In_2456);
nor U98 (N_98,In_1728,In_2152);
xor U99 (N_99,In_1986,In_2284);
and U100 (N_100,In_431,In_2472);
nor U101 (N_101,In_1731,In_1776);
and U102 (N_102,In_1832,In_130);
and U103 (N_103,In_1131,In_2068);
xor U104 (N_104,In_852,In_653);
nand U105 (N_105,In_51,In_534);
xor U106 (N_106,In_1754,In_55);
and U107 (N_107,In_1345,In_745);
and U108 (N_108,In_308,In_792);
or U109 (N_109,In_186,In_1785);
nand U110 (N_110,In_1678,In_162);
nor U111 (N_111,In_1051,In_1072);
or U112 (N_112,In_1798,In_783);
and U113 (N_113,In_1540,In_969);
nor U114 (N_114,In_1647,In_962);
nor U115 (N_115,In_1958,In_2448);
xnor U116 (N_116,In_1652,In_271);
nand U117 (N_117,In_2099,In_279);
nor U118 (N_118,In_712,In_1193);
nor U119 (N_119,In_1042,In_1542);
nor U120 (N_120,In_2418,In_1030);
xnor U121 (N_121,In_1751,In_401);
nor U122 (N_122,In_921,In_1323);
xor U123 (N_123,In_2181,In_2471);
nor U124 (N_124,In_870,In_1208);
nand U125 (N_125,In_988,In_2186);
nand U126 (N_126,In_9,In_1122);
nand U127 (N_127,In_1510,In_1683);
nand U128 (N_128,In_485,In_1309);
xor U129 (N_129,In_311,In_2221);
or U130 (N_130,In_2466,In_2102);
and U131 (N_131,In_1005,In_132);
nor U132 (N_132,In_1268,In_1862);
xnor U133 (N_133,In_2458,In_116);
xnor U134 (N_134,In_1118,In_1270);
xnor U135 (N_135,In_2247,In_1430);
or U136 (N_136,In_1524,In_896);
nor U137 (N_137,In_683,In_1492);
nand U138 (N_138,In_230,In_1416);
nand U139 (N_139,In_1708,In_1318);
and U140 (N_140,In_106,In_844);
and U141 (N_141,In_952,In_2120);
nand U142 (N_142,In_1669,In_540);
nand U143 (N_143,In_1913,In_700);
or U144 (N_144,In_2467,In_23);
nor U145 (N_145,In_1235,In_360);
and U146 (N_146,In_2114,In_621);
xor U147 (N_147,In_1996,In_1014);
nand U148 (N_148,In_978,In_490);
or U149 (N_149,In_1210,In_2242);
and U150 (N_150,In_2282,In_212);
xnor U151 (N_151,In_1393,In_1970);
xnor U152 (N_152,In_1584,In_1168);
xor U153 (N_153,In_2142,In_1760);
or U154 (N_154,In_307,In_1400);
and U155 (N_155,In_2009,In_562);
nand U156 (N_156,In_984,In_1690);
and U157 (N_157,In_1674,In_990);
nor U158 (N_158,In_1528,In_888);
nand U159 (N_159,In_780,In_1717);
xor U160 (N_160,In_8,In_355);
xor U161 (N_161,In_428,In_1392);
xnor U162 (N_162,In_881,In_273);
nor U163 (N_163,In_2440,In_1257);
nor U164 (N_164,In_711,In_1745);
and U165 (N_165,In_438,In_1088);
or U166 (N_166,In_710,In_2260);
nand U167 (N_167,In_1981,In_1872);
or U168 (N_168,In_2220,In_839);
nand U169 (N_169,In_33,In_1579);
xnor U170 (N_170,In_693,In_2128);
nand U171 (N_171,In_810,In_54);
or U172 (N_172,In_681,In_1432);
nor U173 (N_173,In_1306,In_1352);
nor U174 (N_174,In_474,In_538);
and U175 (N_175,In_1753,In_335);
xnor U176 (N_176,In_297,In_2078);
nor U177 (N_177,In_58,In_2460);
nor U178 (N_178,In_2163,In_851);
xnor U179 (N_179,In_833,In_1212);
xor U180 (N_180,In_1505,In_555);
or U181 (N_181,In_1001,In_1580);
xor U182 (N_182,In_383,In_442);
or U183 (N_183,In_180,In_679);
and U184 (N_184,In_49,In_83);
and U185 (N_185,In_2453,In_1818);
and U186 (N_186,In_150,In_1296);
or U187 (N_187,In_568,In_328);
nand U188 (N_188,In_1223,In_2047);
nor U189 (N_189,In_1476,In_1121);
or U190 (N_190,In_2245,In_691);
or U191 (N_191,In_1882,In_415);
xor U192 (N_192,In_665,In_86);
nor U193 (N_193,In_214,In_2174);
and U194 (N_194,In_429,In_1291);
and U195 (N_195,In_1120,In_575);
and U196 (N_196,In_1729,In_228);
and U197 (N_197,In_149,In_2499);
or U198 (N_198,In_1028,In_22);
xnor U199 (N_199,In_295,In_496);
and U200 (N_200,In_2111,In_1171);
xnor U201 (N_201,In_1609,In_1529);
or U202 (N_202,In_570,In_1720);
nand U203 (N_203,In_1639,In_2264);
or U204 (N_204,In_1147,In_445);
nand U205 (N_205,In_1280,In_1321);
and U206 (N_206,In_392,In_518);
nand U207 (N_207,In_2044,In_734);
or U208 (N_208,In_1234,In_1515);
nor U209 (N_209,In_1890,In_2090);
xnor U210 (N_210,In_202,In_862);
nor U211 (N_211,In_1427,In_283);
or U212 (N_212,In_1189,In_1407);
and U213 (N_213,In_650,In_1401);
xnor U214 (N_214,In_1297,In_1463);
nand U215 (N_215,In_1381,In_618);
nor U216 (N_216,In_1809,In_2088);
xor U217 (N_217,In_2011,In_427);
xnor U218 (N_218,In_372,In_741);
or U219 (N_219,In_329,In_1282);
or U220 (N_220,In_2483,In_1842);
nand U221 (N_221,In_1111,In_1713);
nor U222 (N_222,In_613,In_1702);
nand U223 (N_223,In_13,In_1828);
nand U224 (N_224,In_1968,In_371);
and U225 (N_225,In_304,In_1148);
xor U226 (N_226,In_529,In_504);
xnor U227 (N_227,In_40,In_1556);
nor U228 (N_228,In_902,In_325);
or U229 (N_229,In_1971,In_539);
or U230 (N_230,In_1197,In_1465);
xnor U231 (N_231,In_2119,In_2211);
or U232 (N_232,In_1156,In_664);
nor U233 (N_233,In_409,In_127);
nand U234 (N_234,In_1815,In_2234);
nor U235 (N_235,In_692,In_853);
nor U236 (N_236,In_2263,In_2383);
nor U237 (N_237,In_842,In_2177);
nor U238 (N_238,In_1705,In_1383);
xor U239 (N_239,In_2268,In_2107);
nand U240 (N_240,In_938,In_2269);
and U241 (N_241,In_1806,In_1403);
and U242 (N_242,In_2393,In_1274);
nand U243 (N_243,In_973,In_1987);
and U244 (N_244,In_1625,In_2310);
nand U245 (N_245,In_1139,In_722);
nand U246 (N_246,In_2478,In_2084);
or U247 (N_247,In_2249,In_2183);
and U248 (N_248,In_1692,In_829);
nor U249 (N_249,In_516,In_2089);
or U250 (N_250,In_1009,In_802);
and U251 (N_251,In_778,In_1460);
nand U252 (N_252,In_2117,In_804);
or U253 (N_253,In_1490,In_70);
xor U254 (N_254,In_1547,In_714);
and U255 (N_255,In_694,In_405);
and U256 (N_256,In_1106,In_2086);
nor U257 (N_257,In_1765,In_617);
nor U258 (N_258,In_2199,In_1953);
or U259 (N_259,In_2178,In_1482);
xnor U260 (N_260,In_155,In_1721);
and U261 (N_261,In_912,In_2083);
nor U262 (N_262,In_1672,In_227);
nor U263 (N_263,In_2469,In_577);
nor U264 (N_264,In_846,In_942);
nand U265 (N_265,In_2306,In_2402);
and U266 (N_266,In_2058,In_254);
nor U267 (N_267,In_2379,In_1076);
xnor U268 (N_268,In_2134,In_1596);
and U269 (N_269,In_397,In_179);
nand U270 (N_270,In_1397,In_261);
nor U271 (N_271,In_1389,In_1841);
and U272 (N_272,In_1831,In_1474);
or U273 (N_273,In_2170,In_606);
and U274 (N_274,In_1469,In_478);
nand U275 (N_275,In_1205,In_889);
xnor U276 (N_276,In_766,In_1440);
or U277 (N_277,In_582,In_1906);
and U278 (N_278,In_2455,In_1331);
nand U279 (N_279,In_2233,In_472);
nand U280 (N_280,In_751,In_1904);
and U281 (N_281,In_2433,In_1426);
and U282 (N_282,In_2039,In_1999);
xnor U283 (N_283,In_991,In_933);
nand U284 (N_284,In_1819,In_1050);
nand U285 (N_285,In_1812,In_1613);
nor U286 (N_286,In_567,In_211);
nor U287 (N_287,In_1353,In_1065);
or U288 (N_288,In_471,In_1376);
nand U289 (N_289,In_2474,In_977);
or U290 (N_290,In_1356,In_199);
nand U291 (N_291,In_1628,In_920);
nor U292 (N_292,In_1735,In_1633);
xnor U293 (N_293,In_158,In_1421);
xnor U294 (N_294,In_402,In_2238);
nor U295 (N_295,In_52,In_1433);
nor U296 (N_296,In_1926,In_119);
xnor U297 (N_297,In_1518,In_1115);
and U298 (N_298,In_90,In_1875);
and U299 (N_299,In_779,In_937);
nor U300 (N_300,In_334,In_499);
or U301 (N_301,In_2095,In_733);
nor U302 (N_302,In_233,In_1211);
and U303 (N_303,In_259,In_2452);
nor U304 (N_304,In_1676,In_1365);
nand U305 (N_305,In_2108,In_458);
nor U306 (N_306,In_299,In_2126);
xnor U307 (N_307,In_200,In_1902);
or U308 (N_308,In_1727,In_972);
or U309 (N_309,In_2293,In_1017);
nor U310 (N_310,In_1873,In_2320);
nand U311 (N_311,In_1934,In_886);
and U312 (N_312,In_337,In_943);
and U313 (N_313,In_2158,In_2156);
nor U314 (N_314,In_1044,In_219);
xor U315 (N_315,In_1431,In_1138);
and U316 (N_316,In_1157,In_684);
xor U317 (N_317,In_1308,In_528);
xnor U318 (N_318,In_1185,In_1093);
nand U319 (N_319,In_2387,In_201);
nor U320 (N_320,In_1718,In_1418);
xor U321 (N_321,In_1839,In_296);
or U322 (N_322,In_1425,In_2106);
xnor U323 (N_323,In_350,In_1772);
xnor U324 (N_324,In_689,In_1334);
nor U325 (N_325,In_2129,In_2045);
and U326 (N_326,In_362,In_89);
xnor U327 (N_327,In_1845,In_1561);
xor U328 (N_328,In_1680,In_1083);
and U329 (N_329,In_604,In_2321);
or U330 (N_330,In_607,In_1313);
or U331 (N_331,In_1612,In_448);
nor U332 (N_332,In_623,In_1480);
nor U333 (N_333,In_1060,In_1712);
and U334 (N_334,In_1204,In_1077);
nor U335 (N_335,In_1219,In_1513);
and U336 (N_336,In_1670,In_1378);
nor U337 (N_337,In_2332,In_619);
and U338 (N_338,In_584,In_2025);
xnor U339 (N_339,In_1834,In_263);
xor U340 (N_340,In_1850,In_1814);
nor U341 (N_341,In_930,In_1177);
nor U342 (N_342,In_1444,In_1927);
or U343 (N_343,In_1501,In_272);
or U344 (N_344,In_561,In_167);
and U345 (N_345,In_1933,In_860);
or U346 (N_346,In_897,In_1799);
or U347 (N_347,In_1153,In_444);
nand U348 (N_348,In_166,In_2139);
nand U349 (N_349,In_1586,In_1022);
nand U350 (N_350,In_1206,In_2037);
xor U351 (N_351,In_111,In_17);
or U352 (N_352,In_1395,In_1302);
nor U353 (N_353,In_426,In_236);
xnor U354 (N_354,In_620,In_563);
and U355 (N_355,In_2240,In_289);
nand U356 (N_356,In_390,In_2333);
or U357 (N_357,In_2331,In_1011);
nor U358 (N_358,In_1645,In_2278);
xnor U359 (N_359,In_787,In_2363);
xnor U360 (N_360,In_649,In_375);
or U361 (N_361,In_806,In_892);
nor U362 (N_362,In_1959,In_1107);
and U363 (N_363,In_477,In_2307);
and U364 (N_364,In_893,In_2372);
or U365 (N_365,In_460,In_1013);
or U366 (N_366,In_365,In_320);
or U367 (N_367,In_1922,In_363);
xnor U368 (N_368,In_1537,In_103);
or U369 (N_369,In_2096,In_736);
and U370 (N_370,In_1632,In_2354);
nand U371 (N_371,In_1459,In_2141);
xnor U372 (N_372,In_2228,In_2390);
and U373 (N_373,In_1551,In_2131);
xor U374 (N_374,In_2193,In_2135);
nor U375 (N_375,In_294,In_2255);
or U376 (N_376,In_194,In_2032);
nand U377 (N_377,In_151,In_672);
or U378 (N_378,In_868,In_1067);
nand U379 (N_379,In_1844,In_2154);
nor U380 (N_380,In_2484,In_879);
xor U381 (N_381,In_1938,In_321);
nor U382 (N_382,In_2150,In_797);
and U383 (N_383,In_935,In_1598);
xnor U384 (N_384,In_2005,In_455);
and U385 (N_385,In_1668,In_2373);
or U386 (N_386,In_2382,In_1174);
xor U387 (N_387,In_2326,In_2185);
nand U388 (N_388,In_264,In_817);
xnor U389 (N_389,In_945,In_1878);
nor U390 (N_390,In_265,In_1553);
and U391 (N_391,In_2130,In_1454);
nand U392 (N_392,In_2194,In_1545);
and U393 (N_393,In_709,In_660);
nand U394 (N_394,In_2406,In_2189);
and U395 (N_395,In_1945,In_655);
xor U396 (N_396,In_932,In_2376);
and U397 (N_397,In_403,In_1203);
and U398 (N_398,In_773,In_596);
nand U399 (N_399,In_1124,In_916);
nand U400 (N_400,In_639,In_1662);
nor U401 (N_401,In_2007,In_1347);
or U402 (N_402,In_2029,In_1591);
xnor U403 (N_403,In_1687,In_284);
nor U404 (N_404,In_953,In_85);
or U405 (N_405,In_1142,In_2212);
nor U406 (N_406,In_848,In_2392);
xor U407 (N_407,In_1349,In_196);
nor U408 (N_408,In_1034,In_1526);
nor U409 (N_409,In_1716,In_1993);
xnor U410 (N_410,In_520,In_443);
and U411 (N_411,In_1737,In_280);
or U412 (N_412,In_1752,In_1936);
nand U413 (N_413,In_732,In_2143);
nand U414 (N_414,In_828,In_985);
nor U415 (N_415,In_2124,In_2368);
and U416 (N_416,In_1258,In_274);
or U417 (N_417,In_922,In_1254);
or U418 (N_418,In_2358,In_1758);
nand U419 (N_419,In_715,In_322);
nand U420 (N_420,In_2366,In_1242);
xnor U421 (N_421,In_216,In_1538);
xnor U422 (N_422,In_2175,In_1523);
and U423 (N_423,In_407,In_2054);
xnor U424 (N_424,In_2496,In_1181);
nor U425 (N_425,In_2049,In_2051);
nor U426 (N_426,In_675,In_290);
xnor U427 (N_427,In_217,In_338);
and U428 (N_428,In_1464,In_1689);
nand U429 (N_429,In_2295,In_1849);
xnor U430 (N_430,In_2481,In_2276);
nor U431 (N_431,In_1769,In_386);
nor U432 (N_432,In_118,In_1653);
xnor U433 (N_433,In_69,In_244);
nand U434 (N_434,In_1,In_1607);
nand U435 (N_435,In_341,In_855);
xnor U436 (N_436,In_1114,In_117);
xor U437 (N_437,In_349,In_2146);
nor U438 (N_438,In_913,In_178);
or U439 (N_439,In_612,In_2482);
or U440 (N_440,In_854,In_676);
or U441 (N_441,In_359,In_1054);
nand U442 (N_442,In_421,In_998);
or U443 (N_443,In_1169,In_2407);
and U444 (N_444,In_1047,In_1946);
or U445 (N_445,In_1826,In_2087);
xor U446 (N_446,In_2223,In_2115);
nor U447 (N_447,In_915,In_1100);
nand U448 (N_448,In_1424,In_12);
xnor U449 (N_449,In_2201,In_64);
and U450 (N_450,In_0,In_286);
nand U451 (N_451,In_1412,In_759);
nor U452 (N_452,In_1246,In_849);
nand U453 (N_453,In_2436,In_648);
nor U454 (N_454,In_1789,In_2251);
nor U455 (N_455,In_742,In_19);
or U456 (N_456,In_1601,In_1081);
or U457 (N_457,In_2435,In_1599);
nor U458 (N_458,In_1822,In_62);
and U459 (N_459,In_1301,In_586);
or U460 (N_460,In_1236,In_1429);
or U461 (N_461,In_453,In_221);
nand U462 (N_462,In_2125,In_1907);
xnor U463 (N_463,In_1278,In_642);
xnor U464 (N_464,In_46,In_215);
nor U465 (N_465,In_1565,In_968);
or U466 (N_466,In_1281,In_2027);
and U467 (N_467,In_724,In_356);
and U468 (N_468,In_97,In_2327);
xnor U469 (N_469,In_588,In_2442);
nand U470 (N_470,In_267,In_883);
and U471 (N_471,In_1434,In_1207);
xor U472 (N_472,In_2001,In_827);
or U473 (N_473,In_1190,In_501);
xor U474 (N_474,In_2477,In_368);
nand U475 (N_475,In_28,In_1534);
nor U476 (N_476,In_1863,In_63);
nand U477 (N_477,In_975,In_547);
and U478 (N_478,In_807,In_1295);
nor U479 (N_479,In_4,In_2405);
xnor U480 (N_480,In_1357,In_345);
xor U481 (N_481,In_1507,In_417);
xor U482 (N_482,In_2064,In_2316);
and U483 (N_483,In_2267,In_1359);
xor U484 (N_484,In_826,In_1891);
nor U485 (N_485,In_2046,In_1626);
nand U486 (N_486,In_1773,In_581);
nor U487 (N_487,In_1191,In_1445);
and U488 (N_488,In_133,In_2384);
and U489 (N_489,In_1200,In_353);
nor U490 (N_490,In_1784,In_856);
xor U491 (N_491,In_319,In_1780);
nand U492 (N_492,In_2497,In_396);
xor U493 (N_493,In_2318,In_824);
nor U494 (N_494,In_566,In_776);
and U495 (N_495,In_2014,In_695);
and U496 (N_496,In_656,In_20);
nand U497 (N_497,In_2476,In_946);
nand U498 (N_498,In_2022,In_1555);
nor U499 (N_499,In_91,In_393);
xor U500 (N_500,In_1846,In_1575);
xnor U501 (N_501,In_2439,In_1649);
xnor U502 (N_502,In_1140,In_1982);
and U503 (N_503,In_1835,In_101);
nor U504 (N_504,In_1770,In_843);
nor U505 (N_505,In_1499,In_1063);
or U506 (N_506,In_772,In_2296);
xor U507 (N_507,In_11,In_936);
xnor U508 (N_508,In_1883,In_1387);
or U509 (N_509,In_1696,In_1559);
or U510 (N_510,In_763,In_1125);
nand U511 (N_511,In_1602,In_1825);
xnor U512 (N_512,In_963,In_96);
or U513 (N_513,In_815,In_775);
or U514 (N_514,In_2023,In_2216);
nor U515 (N_515,In_1859,In_674);
nor U516 (N_516,In_1643,In_2285);
xnor U517 (N_517,In_2343,In_2494);
and U518 (N_518,In_1008,In_2042);
nor U519 (N_519,In_2008,In_1025);
and U520 (N_520,In_731,In_292);
or U521 (N_521,In_887,In_951);
or U522 (N_522,In_234,In_1238);
or U523 (N_523,In_527,In_2202);
nor U524 (N_524,In_603,In_1150);
nor U525 (N_525,In_521,In_905);
or U526 (N_526,In_125,In_1711);
xnor U527 (N_527,In_554,In_2237);
nand U528 (N_528,In_605,In_1778);
or U529 (N_529,In_717,In_408);
or U530 (N_530,In_39,In_1929);
xor U531 (N_531,In_239,In_2155);
nor U532 (N_532,In_95,In_611);
nand U533 (N_533,In_2434,In_447);
and U534 (N_534,In_995,In_754);
xnor U535 (N_535,In_812,In_1126);
or U536 (N_536,In_1078,In_670);
nor U537 (N_537,In_1664,In_313);
or U538 (N_538,In_1213,In_1657);
and U539 (N_539,In_2398,In_1759);
or U540 (N_540,In_1983,In_1228);
nor U541 (N_541,In_2004,In_904);
or U542 (N_542,In_1225,In_2450);
xor U543 (N_543,In_1802,In_1417);
xnor U544 (N_544,In_1794,In_1133);
and U545 (N_545,In_316,In_366);
or U546 (N_546,In_771,In_2348);
nor U547 (N_547,In_2300,In_2182);
xnor U548 (N_548,In_558,In_713);
nand U549 (N_549,In_1438,In_268);
and U550 (N_550,In_108,In_958);
and U551 (N_551,In_542,In_845);
and U552 (N_552,In_791,In_1289);
nor U553 (N_553,In_1823,In_1976);
or U554 (N_554,In_1605,In_2301);
nor U555 (N_555,In_589,In_1055);
nor U556 (N_556,In_2180,In_1975);
xor U557 (N_557,In_1833,In_744);
nand U558 (N_558,In_2243,In_1312);
nor U559 (N_559,In_1450,In_1723);
xnor U560 (N_560,In_587,In_960);
xor U561 (N_561,In_394,In_2495);
or U562 (N_562,In_1233,In_1648);
xor U563 (N_563,In_1851,In_914);
xor U564 (N_564,In_1382,In_25);
and U565 (N_565,In_126,In_1340);
and U566 (N_566,In_1145,In_508);
nor U567 (N_567,In_470,In_2171);
and U568 (N_568,In_2097,In_1898);
and U569 (N_569,In_1116,In_1455);
and U570 (N_570,In_1532,In_30);
xor U571 (N_571,In_1837,In_1284);
nand U572 (N_572,In_1925,In_43);
or U573 (N_573,In_1762,In_781);
xnor U574 (N_574,In_1059,In_452);
and U575 (N_575,In_1944,In_1298);
nor U576 (N_576,In_2020,In_2371);
nor U577 (N_577,In_1056,In_2449);
or U578 (N_578,In_2082,In_1057);
or U579 (N_579,In_2077,In_1221);
or U580 (N_580,In_1667,In_1187);
or U581 (N_581,In_147,In_1245);
nor U582 (N_582,In_2352,In_2281);
xnor U583 (N_583,In_885,In_598);
nand U584 (N_584,In_2294,In_831);
or U585 (N_585,In_424,In_2258);
nor U586 (N_586,In_35,In_2377);
xor U587 (N_587,In_87,In_1869);
xor U588 (N_588,In_1373,In_2322);
nand U589 (N_589,In_107,In_629);
or U590 (N_590,In_2364,In_1475);
nand U591 (N_591,In_2279,In_595);
nand U592 (N_592,In_1506,In_1606);
or U593 (N_593,In_1194,In_2034);
nor U594 (N_594,In_1631,In_1006);
or U595 (N_595,In_1592,In_479);
nand U596 (N_596,In_777,In_1594);
xnor U597 (N_597,In_1774,In_2259);
and U598 (N_598,In_2445,In_2437);
or U599 (N_599,In_34,In_1827);
xnor U600 (N_600,In_663,In_600);
nor U601 (N_601,In_2145,In_1724);
or U602 (N_602,In_1682,In_213);
xnor U603 (N_603,In_1744,In_1027);
and U604 (N_604,In_466,In_1800);
xor U605 (N_605,In_1546,In_2166);
nand U606 (N_606,In_2314,In_1002);
nand U607 (N_607,In_1805,In_1761);
or U608 (N_608,In_1487,In_73);
nand U609 (N_609,In_138,In_1237);
xor U610 (N_610,In_161,In_1918);
nor U611 (N_611,In_530,In_1196);
and U612 (N_612,In_1250,In_1495);
nor U613 (N_613,In_1144,In_1368);
xor U614 (N_614,In_1162,In_1865);
and U615 (N_615,In_841,In_2250);
xnor U616 (N_616,In_884,In_303);
or U617 (N_617,In_287,In_369);
xnor U618 (N_618,In_2487,In_1739);
nor U619 (N_619,In_29,In_99);
nor U620 (N_620,In_1276,In_1484);
and U621 (N_621,In_514,In_805);
xor U622 (N_622,In_2167,In_2133);
nor U623 (N_623,In_467,In_871);
nand U624 (N_624,In_919,In_768);
xor U625 (N_625,In_1654,In_1288);
and U626 (N_626,In_2400,In_728);
or U627 (N_627,In_1707,In_2218);
nor U628 (N_628,In_1175,In_1031);
xor U629 (N_629,In_758,In_1231);
and U630 (N_630,In_602,In_976);
or U631 (N_631,In_1328,In_1889);
nand U632 (N_632,In_796,In_398);
or U633 (N_633,In_1449,In_610);
or U634 (N_634,In_677,In_2328);
xor U635 (N_635,In_1700,In_387);
and U636 (N_636,In_2413,In_309);
and U637 (N_637,In_659,In_1714);
xnor U638 (N_638,In_970,In_2370);
nor U639 (N_639,In_908,In_425);
or U640 (N_640,In_1600,In_310);
or U641 (N_641,In_720,In_226);
nand U642 (N_642,In_974,In_446);
nor U643 (N_643,In_240,In_2313);
nor U644 (N_644,In_1748,In_2432);
nand U645 (N_645,In_861,In_1956);
or U646 (N_646,In_160,In_374);
xor U647 (N_647,In_737,In_2138);
nor U648 (N_648,In_1887,In_1380);
nor U649 (N_649,In_865,In_1581);
nor U650 (N_650,In_293,In_1262);
and U651 (N_651,In_464,In_2116);
or U652 (N_652,In_580,In_255);
or U653 (N_653,In_1267,In_1964);
nand U654 (N_654,In_1094,In_1655);
nor U655 (N_655,In_971,In_1152);
or U656 (N_656,In_1766,In_2395);
and U657 (N_657,In_498,In_191);
or U658 (N_658,In_1489,In_223);
and U659 (N_659,In_2280,In_1572);
nand U660 (N_660,In_1422,In_1277);
nor U661 (N_661,In_2021,In_330);
nand U662 (N_662,In_2464,In_2465);
xnor U663 (N_663,In_757,In_15);
nor U664 (N_664,In_765,In_1779);
nor U665 (N_665,In_2289,In_2344);
xor U666 (N_666,In_901,In_1589);
and U667 (N_667,In_2113,In_1146);
or U668 (N_668,In_2149,In_2498);
or U669 (N_669,In_449,In_2374);
and U670 (N_670,In_1409,In_1217);
or U671 (N_671,In_1951,In_959);
nand U672 (N_672,In_298,In_66);
and U673 (N_673,In_1597,In_2380);
and U674 (N_674,In_1180,In_1261);
and U675 (N_675,In_1804,In_1738);
xnor U676 (N_676,In_1629,In_1016);
nor U677 (N_677,In_800,In_899);
nand U678 (N_678,In_1375,In_112);
or U679 (N_679,In_858,In_834);
and U680 (N_680,In_1021,In_545);
nor U681 (N_681,In_2016,In_237);
or U682 (N_682,In_1896,In_579);
and U683 (N_683,In_1260,In_666);
nor U684 (N_684,In_926,In_654);
or U685 (N_685,In_1004,In_1746);
xnor U686 (N_686,In_2428,In_2225);
and U687 (N_687,In_2347,In_1036);
xnor U688 (N_688,In_140,In_635);
and U689 (N_689,In_2311,In_1497);
nor U690 (N_690,In_1069,In_404);
nor U691 (N_691,In_1466,In_1188);
and U692 (N_692,In_726,In_2067);
nor U693 (N_693,In_1567,In_640);
nand U694 (N_694,In_188,In_2219);
xor U695 (N_695,In_535,In_177);
or U696 (N_696,In_818,In_75);
and U697 (N_697,In_1179,In_989);
or U698 (N_698,In_60,In_2360);
xor U699 (N_699,In_2071,In_2248);
nor U700 (N_700,In_515,In_348);
nand U701 (N_701,In_1243,In_1184);
nand U702 (N_702,In_1183,In_585);
xor U703 (N_703,In_2454,In_413);
and U704 (N_704,In_14,In_2222);
nor U705 (N_705,In_1350,In_537);
or U706 (N_706,In_591,In_799);
nor U707 (N_707,In_2463,In_44);
and U708 (N_708,In_190,In_157);
and U709 (N_709,In_257,In_1136);
xnor U710 (N_710,In_1972,In_2198);
nand U711 (N_711,In_400,In_2443);
and U712 (N_712,In_774,In_192);
or U713 (N_713,In_2479,In_154);
nor U714 (N_714,In_1610,In_1319);
nor U715 (N_715,In_1471,In_1920);
or U716 (N_716,In_135,In_2018);
and U717 (N_717,In_462,In_376);
xnor U718 (N_718,In_176,In_512);
and U719 (N_719,In_1719,In_2069);
xor U720 (N_720,In_1075,In_927);
xnor U721 (N_721,In_1062,In_1195);
nor U722 (N_722,In_100,In_788);
xor U723 (N_723,In_473,In_519);
nand U724 (N_724,In_2486,In_61);
or U725 (N_725,In_2195,In_1332);
or U726 (N_726,In_2420,In_533);
nor U727 (N_727,In_2061,In_1038);
and U728 (N_728,In_532,In_71);
or U729 (N_729,In_696,In_2210);
or U730 (N_730,In_2335,In_2036);
nand U731 (N_731,In_253,In_2419);
xnor U732 (N_732,In_7,In_1498);
nor U733 (N_733,In_2388,In_262);
or U734 (N_734,In_2169,In_2191);
xnor U735 (N_735,In_2299,In_420);
nand U736 (N_736,In_948,In_1155);
nor U737 (N_737,In_1836,In_2341);
nand U738 (N_738,In_77,In_816);
xnor U739 (N_739,In_144,In_1453);
nand U740 (N_740,In_1980,In_708);
nor U741 (N_741,In_1186,In_869);
nand U742 (N_742,In_1390,In_1994);
xor U743 (N_743,In_251,In_2346);
nand U744 (N_744,In_246,In_204);
or U745 (N_745,In_830,In_275);
or U746 (N_746,In_1103,In_2339);
nor U747 (N_747,In_2309,In_1477);
and U748 (N_748,In_26,In_1595);
and U749 (N_749,In_2275,In_1656);
or U750 (N_750,In_2200,In_57);
and U751 (N_751,In_647,In_10);
xor U752 (N_752,In_2144,In_301);
nor U753 (N_753,In_1514,In_1533);
or U754 (N_754,In_1519,In_1767);
nand U755 (N_755,In_822,In_56);
or U756 (N_756,In_1989,In_336);
or U757 (N_757,In_1677,In_2030);
xor U758 (N_758,In_2215,In_182);
nor U759 (N_759,In_510,In_638);
xnor U760 (N_760,In_1026,In_27);
nor U761 (N_761,In_2303,In_1377);
nor U762 (N_762,In_1473,In_185);
xnor U763 (N_763,In_941,In_964);
or U764 (N_764,In_1315,In_900);
or U765 (N_765,In_572,In_1128);
and U766 (N_766,In_2002,In_258);
or U767 (N_767,In_2459,In_2013);
and U768 (N_768,In_1660,In_1880);
or U769 (N_769,In_1096,In_2072);
nor U770 (N_770,In_2076,In_1924);
and U771 (N_771,In_705,In_2101);
nand U772 (N_772,In_152,In_459);
nor U773 (N_773,In_2489,In_318);
nand U774 (N_774,In_1420,In_955);
and U775 (N_775,In_1374,In_1706);
and U776 (N_776,In_1747,In_2257);
nand U777 (N_777,In_1867,In_622);
nand U778 (N_778,In_967,In_1364);
and U779 (N_779,In_662,In_1684);
or U780 (N_780,In_1895,In_1264);
or U781 (N_781,In_2031,In_1984);
nor U782 (N_782,In_680,In_1265);
nor U783 (N_783,In_379,In_1307);
or U784 (N_784,In_2362,In_323);
nand U785 (N_785,In_170,In_1446);
and U786 (N_786,In_1292,In_1415);
nand U787 (N_787,In_1909,In_1066);
or U788 (N_788,In_1901,In_1327);
xor U789 (N_789,In_198,In_357);
nand U790 (N_790,In_2168,In_1624);
nand U791 (N_791,In_898,In_382);
nor U792 (N_792,In_1325,In_1462);
xnor U793 (N_793,In_1406,In_1079);
nor U794 (N_794,In_2367,In_923);
and U795 (N_795,In_1950,In_143);
nand U796 (N_796,In_1113,In_1709);
nand U797 (N_797,In_564,In_450);
or U798 (N_798,In_1019,In_1486);
xor U799 (N_799,In_544,In_247);
or U800 (N_800,In_702,In_996);
xor U801 (N_801,In_574,In_1080);
and U802 (N_802,In_482,In_42);
and U803 (N_803,In_895,In_276);
or U804 (N_804,In_131,In_489);
nand U805 (N_805,In_782,In_631);
and U806 (N_806,In_747,In_821);
nor U807 (N_807,In_1886,In_187);
xnor U808 (N_808,In_753,In_1240);
or U809 (N_809,In_994,In_525);
and U810 (N_810,In_1099,In_1801);
or U811 (N_811,In_719,In_523);
nand U812 (N_812,In_314,In_1900);
or U813 (N_813,In_2369,In_1394);
nor U814 (N_814,In_1868,In_2056);
nor U815 (N_815,In_1082,In_92);
nor U816 (N_816,In_2298,In_2359);
nor U817 (N_817,In_249,In_1511);
xor U818 (N_818,In_1222,In_1803);
or U819 (N_819,In_361,In_1230);
or U820 (N_820,In_2425,In_1611);
or U821 (N_821,In_1644,In_281);
and U822 (N_822,In_2239,In_813);
nand U823 (N_823,In_1137,In_2355);
nand U824 (N_824,In_16,In_1554);
and U825 (N_825,In_2122,In_2035);
or U826 (N_826,In_793,In_385);
nand U827 (N_827,In_626,In_164);
xor U828 (N_828,In_1071,In_1379);
and U829 (N_829,In_1630,In_911);
nor U830 (N_830,In_2147,In_1447);
nor U831 (N_831,In_1675,In_480);
nand U832 (N_832,In_2232,In_1992);
and U833 (N_833,In_939,In_1336);
nand U834 (N_834,In_1879,In_1304);
or U835 (N_835,In_391,In_1178);
or U836 (N_836,In_1339,In_1130);
and U837 (N_837,In_434,In_1894);
nor U838 (N_838,In_2470,In_457);
nor U839 (N_839,In_526,In_124);
and U840 (N_840,In_351,In_2006);
or U841 (N_841,In_1960,In_1522);
nand U842 (N_842,In_2334,In_838);
nand U843 (N_843,In_1402,In_1160);
nand U844 (N_844,In_1092,In_2140);
or U845 (N_845,In_488,In_120);
and U846 (N_846,In_673,In_2438);
xnor U847 (N_847,In_2396,In_193);
or U848 (N_848,In_1967,In_1248);
nor U849 (N_849,In_252,In_1949);
nor U850 (N_850,In_1941,In_949);
xnor U851 (N_851,In_950,In_1860);
and U852 (N_852,In_451,In_1439);
or U853 (N_853,In_608,In_465);
nand U854 (N_854,In_1286,In_440);
and U855 (N_855,In_1253,In_1173);
xor U856 (N_856,In_1348,In_907);
xor U857 (N_857,In_1214,In_68);
nor U858 (N_858,In_505,In_836);
nor U859 (N_859,In_1903,In_218);
and U860 (N_860,In_59,In_1688);
nand U861 (N_861,In_1661,In_614);
nand U862 (N_862,In_377,In_1671);
nor U863 (N_863,In_168,In_2254);
nand U864 (N_864,In_1423,In_1303);
nor U865 (N_865,In_1216,In_1876);
nor U866 (N_866,In_669,In_5);
nor U867 (N_867,In_739,In_1635);
or U868 (N_868,In_1811,In_1517);
nor U869 (N_869,In_1256,In_241);
or U870 (N_870,In_1244,In_1608);
and U871 (N_871,In_560,In_1419);
nor U872 (N_872,In_21,In_1979);
or U873 (N_873,In_2209,In_389);
and U874 (N_874,In_1961,In_1010);
nor U875 (N_875,In_1029,In_667);
xor U876 (N_876,In_2017,In_1468);
nor U877 (N_877,In_552,In_2485);
or U878 (N_878,In_2110,In_1543);
nor U879 (N_879,In_1892,In_2184);
or U880 (N_880,In_463,In_550);
or U881 (N_881,In_2003,In_1743);
nor U882 (N_882,In_1158,In_1525);
or U883 (N_883,In_1782,In_2253);
nand U884 (N_884,In_2043,In_2094);
or U885 (N_885,In_1615,In_2266);
or U886 (N_886,In_2426,In_536);
xor U887 (N_887,In_1369,In_1557);
and U888 (N_888,In_1921,In_2375);
or U889 (N_889,In_1263,In_1847);
nor U890 (N_890,In_1048,In_2337);
nor U891 (N_891,In_468,In_789);
nand U892 (N_892,In_671,In_1202);
nand U893 (N_893,In_743,In_1991);
and U894 (N_894,In_2336,In_208);
or U895 (N_895,In_1558,In_1691);
and U896 (N_896,In_1255,In_2208);
nand U897 (N_897,In_378,In_1621);
nand U898 (N_898,In_553,In_487);
xor U899 (N_899,In_1252,In_436);
nor U900 (N_900,In_1919,In_1413);
xnor U901 (N_901,In_1651,In_764);
nand U902 (N_902,In_1940,In_1681);
nor U903 (N_903,In_1590,In_1808);
nand U904 (N_904,In_74,In_104);
and U905 (N_905,In_2461,In_1923);
nand U906 (N_906,In_1064,In_495);
xnor U907 (N_907,In_2059,In_1172);
nand U908 (N_908,In_1990,In_2048);
and U909 (N_909,In_1300,In_98);
xnor U910 (N_910,In_414,In_1816);
or U911 (N_911,In_1703,In_1247);
or U912 (N_912,In_2315,In_1456);
nand U913 (N_913,In_2132,In_2403);
xor U914 (N_914,In_769,In_1905);
or U915 (N_915,In_2123,In_1616);
and U916 (N_916,In_1650,In_3);
and U917 (N_917,In_1091,In_1915);
or U918 (N_918,In_1694,In_866);
xnor U919 (N_919,In_343,In_1848);
or U920 (N_920,In_2421,In_388);
xnor U921 (N_921,In_601,In_1916);
xnor U922 (N_922,In_1215,In_109);
nand U923 (N_923,In_1777,In_2028);
and U924 (N_924,In_992,In_229);
or U925 (N_925,In_1496,In_770);
or U926 (N_926,In_2277,In_628);
or U927 (N_927,In_760,In_1698);
xnor U928 (N_928,In_153,In_1583);
xor U929 (N_929,In_646,In_1560);
and U930 (N_930,In_1884,In_1324);
xor U931 (N_931,In_2353,In_1166);
or U932 (N_932,In_2350,In_2308);
xnor U933 (N_933,In_1974,In_524);
xor U934 (N_934,In_122,In_1965);
and U935 (N_935,In_2424,In_1398);
or U936 (N_936,In_1201,In_925);
nor U937 (N_937,In_2229,In_2091);
xor U938 (N_938,In_1220,In_1399);
and U939 (N_939,In_592,In_986);
or U940 (N_940,In_1509,In_1618);
nand U941 (N_941,In_716,In_1763);
nand U942 (N_942,In_2214,In_1229);
or U943 (N_943,In_2324,In_2);
nor U944 (N_944,In_1396,In_1502);
or U945 (N_945,In_93,In_175);
xnor U946 (N_946,In_979,In_347);
nor U947 (N_947,In_333,In_1614);
or U948 (N_948,In_1161,In_1914);
nor U949 (N_949,In_78,In_1129);
and U950 (N_950,In_1820,In_556);
nand U951 (N_951,In_79,In_721);
nand U952 (N_952,In_1531,In_183);
xor U953 (N_953,In_2224,In_1512);
nand U954 (N_954,In_1552,In_701);
nor U955 (N_955,In_352,In_260);
nand U956 (N_956,In_1102,In_1855);
xnor U957 (N_957,In_2062,In_2148);
nor U958 (N_958,In_476,In_1311);
nor U959 (N_959,In_756,In_2074);
and U960 (N_960,In_2287,In_1043);
nor U961 (N_961,In_738,In_1854);
xnor U962 (N_962,In_2112,In_1127);
and U963 (N_963,In_1741,In_1749);
nor U964 (N_964,In_210,In_1757);
nor U965 (N_965,In_245,In_599);
or U966 (N_966,In_32,In_1090);
nor U967 (N_967,In_1141,In_2231);
and U968 (N_968,In_929,In_1622);
nor U969 (N_969,In_1977,In_1893);
or U970 (N_970,In_411,In_2446);
or U971 (N_971,In_980,In_1032);
and U972 (N_972,In_1659,In_1479);
nor U973 (N_973,In_880,In_2480);
xor U974 (N_974,In_2391,In_37);
nand U975 (N_975,In_102,In_2207);
xnor U976 (N_976,In_418,In_2070);
or U977 (N_977,In_1226,In_454);
or U978 (N_978,In_410,In_2386);
xor U979 (N_979,In_53,In_966);
xor U980 (N_980,In_2427,In_129);
nand U981 (N_981,In_1578,In_206);
nor U982 (N_982,In_370,In_2261);
and U983 (N_983,In_2236,In_637);
nor U984 (N_984,In_1358,In_982);
xnor U985 (N_985,In_145,In_1771);
and U986 (N_986,In_1037,In_502);
nor U987 (N_987,In_2291,In_84);
nand U988 (N_988,In_2026,In_1973);
xor U989 (N_989,In_1370,In_340);
or U990 (N_990,In_209,In_1361);
xor U991 (N_991,In_578,In_2100);
nor U992 (N_992,In_331,In_658);
xor U993 (N_993,In_859,In_2491);
nor U994 (N_994,In_2162,In_136);
nor U995 (N_995,In_837,In_1408);
xnor U996 (N_996,In_571,In_1098);
xor U997 (N_997,In_2137,In_291);
nor U998 (N_998,In_1840,In_2197);
xnor U999 (N_999,In_494,In_456);
nand U1000 (N_1000,In_755,In_1391);
nor U1001 (N_1001,In_1734,In_1658);
and U1002 (N_1002,In_1722,In_1199);
nand U1003 (N_1003,In_493,In_1619);
xnor U1004 (N_1004,In_342,In_1764);
nor U1005 (N_1005,In_2092,In_1061);
xor U1006 (N_1006,In_1317,In_1259);
xor U1007 (N_1007,In_2447,In_1360);
and U1008 (N_1008,In_1733,In_1481);
and U1009 (N_1009,In_2389,In_189);
or U1010 (N_1010,In_339,In_1045);
nand U1011 (N_1011,In_2410,In_2265);
nand U1012 (N_1012,In_2416,In_1007);
and U1013 (N_1013,In_1937,In_668);
nand U1014 (N_1014,In_1686,In_517);
xnor U1015 (N_1015,In_2109,In_1750);
nand U1016 (N_1016,In_678,In_2179);
and U1017 (N_1017,In_1952,In_1058);
or U1018 (N_1018,In_1405,In_433);
xor U1019 (N_1019,In_1149,In_1467);
and U1020 (N_1020,In_1693,In_906);
xor U1021 (N_1021,In_1363,In_593);
or U1022 (N_1022,In_957,In_875);
nor U1023 (N_1023,In_548,In_840);
nor U1024 (N_1024,In_511,In_801);
or U1025 (N_1025,In_643,In_1143);
and U1026 (N_1026,In_441,In_509);
xor U1027 (N_1027,In_2401,In_2357);
xnor U1028 (N_1028,In_2127,In_1123);
xor U1029 (N_1029,In_931,In_1603);
or U1030 (N_1030,In_2270,In_123);
and U1031 (N_1031,In_1813,In_1955);
xnor U1032 (N_1032,In_1638,In_248);
nor U1033 (N_1033,In_469,In_1275);
or U1034 (N_1034,In_2422,In_2351);
and U1035 (N_1035,In_1314,In_1617);
xnor U1036 (N_1036,In_644,In_1119);
and U1037 (N_1037,In_2256,In_2252);
and U1038 (N_1038,In_2121,In_2206);
or U1039 (N_1039,In_423,In_346);
xnor U1040 (N_1040,In_381,In_627);
xnor U1041 (N_1041,In_121,In_2338);
nand U1042 (N_1042,In_1530,In_878);
and U1043 (N_1043,In_1574,In_1797);
nand U1044 (N_1044,In_1783,In_690);
nor U1045 (N_1045,In_847,In_2297);
or U1046 (N_1046,In_497,In_2161);
xor U1047 (N_1047,In_1775,In_2409);
or U1048 (N_1048,In_2423,In_1414);
xor U1049 (N_1049,In_2414,In_1888);
nand U1050 (N_1050,In_1117,In_1338);
and U1051 (N_1051,In_1112,In_1232);
xor U1052 (N_1052,In_173,In_1279);
xor U1053 (N_1053,In_2093,In_1159);
nor U1054 (N_1054,In_867,In_2381);
and U1055 (N_1055,In_864,In_81);
and U1056 (N_1056,In_1566,In_1461);
or U1057 (N_1057,In_2235,In_633);
and U1058 (N_1058,In_1493,In_1699);
and U1059 (N_1059,In_541,In_163);
and U1060 (N_1060,In_727,In_1355);
nor U1061 (N_1061,In_1871,In_1041);
xor U1062 (N_1062,In_2000,In_1320);
and U1063 (N_1063,In_2024,In_65);
and U1064 (N_1064,In_2431,In_909);
and U1065 (N_1065,In_954,In_2394);
and U1066 (N_1066,In_1351,In_863);
xnor U1067 (N_1067,In_50,In_2290);
or U1068 (N_1068,In_1877,In_197);
nor U1069 (N_1069,In_278,In_1874);
or U1070 (N_1070,In_220,In_2019);
and U1071 (N_1071,In_850,In_1985);
or U1072 (N_1072,In_416,In_1908);
nand U1073 (N_1073,In_2408,In_195);
nor U1074 (N_1074,In_288,In_687);
or U1075 (N_1075,In_546,In_2473);
and U1076 (N_1076,In_1167,In_82);
or U1077 (N_1077,In_2103,In_636);
xnor U1078 (N_1078,In_395,In_1478);
xor U1079 (N_1079,In_1053,In_890);
nand U1080 (N_1080,In_1085,In_857);
and U1081 (N_1081,In_1969,In_384);
and U1082 (N_1082,In_2272,In_1371);
xor U1083 (N_1083,In_1928,In_1679);
xnor U1084 (N_1084,In_1164,In_1073);
nand U1085 (N_1085,In_1269,In_437);
nor U1086 (N_1086,In_651,In_876);
or U1087 (N_1087,In_506,In_704);
and U1088 (N_1088,In_762,In_1571);
nand U1089 (N_1089,In_1249,In_1807);
xor U1090 (N_1090,In_1521,In_2055);
nor U1091 (N_1091,In_306,In_1105);
and U1092 (N_1092,In_2274,In_917);
nor U1093 (N_1093,In_1577,In_703);
or U1094 (N_1094,In_1227,In_1885);
xnor U1095 (N_1095,In_1251,In_1852);
and U1096 (N_1096,In_1343,In_2085);
nor U1097 (N_1097,In_1443,In_2157);
or U1098 (N_1098,In_305,In_2105);
or U1099 (N_1099,In_1585,In_2033);
or U1100 (N_1100,In_142,In_819);
and U1101 (N_1101,In_2468,In_2187);
nand U1102 (N_1102,In_1241,In_2213);
nor U1103 (N_1103,In_412,In_983);
nor U1104 (N_1104,In_232,In_1911);
xor U1105 (N_1105,In_317,In_1451);
nand U1106 (N_1106,In_492,In_159);
nand U1107 (N_1107,In_2292,In_2457);
or U1108 (N_1108,In_1576,In_1500);
and U1109 (N_1109,In_2378,In_1790);
xnor U1110 (N_1110,In_1954,In_31);
nand U1111 (N_1111,In_1942,In_1285);
nand U1112 (N_1112,In_1310,In_1442);
xnor U1113 (N_1113,In_1549,In_1725);
nand U1114 (N_1114,In_1978,In_2412);
or U1115 (N_1115,In_171,In_461);
nor U1116 (N_1116,In_2451,In_422);
or U1117 (N_1117,In_2038,In_891);
and U1118 (N_1118,In_1293,In_1386);
or U1119 (N_1119,In_1861,In_1287);
nand U1120 (N_1120,In_597,In_1074);
nand U1121 (N_1121,In_256,In_557);
xnor U1122 (N_1122,In_114,In_181);
nor U1123 (N_1123,In_1988,In_1095);
nor U1124 (N_1124,In_2057,In_1544);
and U1125 (N_1125,In_1640,In_1012);
nand U1126 (N_1126,In_486,In_1756);
nand U1127 (N_1127,In_2226,In_2196);
or U1128 (N_1128,In_503,In_940);
nor U1129 (N_1129,In_326,In_2349);
nor U1130 (N_1130,In_1198,In_115);
nor U1131 (N_1131,In_2188,In_697);
and U1132 (N_1132,In_1385,In_1035);
nor U1133 (N_1133,In_1642,In_2340);
nor U1134 (N_1134,In_1726,In_1821);
and U1135 (N_1135,In_1623,In_2041);
and U1136 (N_1136,In_573,In_146);
nor U1137 (N_1137,In_1939,In_45);
nand U1138 (N_1138,In_1272,In_2159);
or U1139 (N_1139,In_2192,In_203);
xor U1140 (N_1140,In_1646,In_874);
and U1141 (N_1141,In_2356,In_2063);
or U1142 (N_1142,In_1344,In_2492);
nor U1143 (N_1143,In_740,In_1485);
or U1144 (N_1144,In_795,In_1995);
or U1145 (N_1145,In_1367,In_798);
and U1146 (N_1146,In_1736,In_2164);
and U1147 (N_1147,In_269,In_2052);
or U1148 (N_1148,In_1015,In_207);
and U1149 (N_1149,In_657,In_2104);
xnor U1150 (N_1150,In_2330,In_1020);
nand U1151 (N_1151,In_1787,In_2227);
nand U1152 (N_1152,In_1910,In_1299);
and U1153 (N_1153,In_956,In_1824);
nor U1154 (N_1154,In_1182,In_1192);
nor U1155 (N_1155,In_616,In_48);
or U1156 (N_1156,In_1330,In_1294);
and U1157 (N_1157,In_1362,In_1087);
nor U1158 (N_1158,In_1704,In_2065);
nor U1159 (N_1159,In_2073,In_1341);
nand U1160 (N_1160,In_2172,In_1209);
and U1161 (N_1161,In_1569,In_2490);
and U1162 (N_1162,In_1931,In_1239);
xor U1163 (N_1163,In_1070,In_729);
or U1164 (N_1164,In_1641,In_1110);
nor U1165 (N_1165,In_624,In_1170);
nand U1166 (N_1166,In_803,In_559);
and U1167 (N_1167,In_924,In_1108);
nor U1168 (N_1168,In_1966,In_1039);
nand U1169 (N_1169,In_315,In_435);
nor U1170 (N_1170,In_1354,In_1957);
xnor U1171 (N_1171,In_1963,In_1810);
or U1172 (N_1172,In_1273,In_1472);
nand U1173 (N_1173,In_2342,In_1564);
nand U1174 (N_1174,In_134,In_72);
nand U1175 (N_1175,In_1864,In_169);
nor U1176 (N_1176,In_2273,In_2241);
xor U1177 (N_1177,In_2080,In_918);
and U1178 (N_1178,In_1795,In_1504);
nor U1179 (N_1179,In_1742,In_1695);
nand U1180 (N_1180,In_139,In_1305);
nand U1181 (N_1181,In_999,In_1101);
xor U1182 (N_1182,In_1089,In_1023);
xor U1183 (N_1183,In_2079,In_76);
nor U1184 (N_1184,In_1948,In_1715);
nor U1185 (N_1185,In_1109,In_1342);
nand U1186 (N_1186,In_944,In_1483);
and U1187 (N_1187,In_491,In_24);
nand U1188 (N_1188,In_725,In_576);
or U1189 (N_1189,In_1329,In_2060);
or U1190 (N_1190,In_1604,In_1673);
and U1191 (N_1191,In_993,In_2012);
nand U1192 (N_1192,In_1796,In_2312);
or U1193 (N_1193,In_1428,In_1384);
or U1194 (N_1194,In_522,In_2283);
or U1195 (N_1195,In_1520,In_88);
and U1196 (N_1196,In_682,In_2053);
xnor U1197 (N_1197,In_2173,In_882);
or U1198 (N_1198,In_1458,In_1755);
or U1199 (N_1199,In_1539,In_2385);
xor U1200 (N_1200,In_1853,In_634);
xnor U1201 (N_1201,In_1866,In_2040);
nor U1202 (N_1202,In_947,In_1781);
and U1203 (N_1203,In_1104,In_2404);
nor U1204 (N_1204,In_36,In_1536);
or U1205 (N_1205,In_1224,In_1046);
and U1206 (N_1206,In_1788,In_1768);
nor U1207 (N_1207,In_2066,In_1134);
nor U1208 (N_1208,In_205,In_1730);
or U1209 (N_1209,In_1494,In_749);
xor U1210 (N_1210,In_1830,In_324);
nor U1211 (N_1211,In_652,In_1665);
or U1212 (N_1212,In_590,In_238);
nand U1213 (N_1213,In_1786,In_832);
xnor U1214 (N_1214,In_2323,In_2361);
nor U1215 (N_1215,In_934,In_38);
xnor U1216 (N_1216,In_1052,In_698);
and U1217 (N_1217,In_811,In_2462);
nor U1218 (N_1218,In_1899,In_327);
nor U1219 (N_1219,In_1593,In_707);
xor U1220 (N_1220,In_1163,In_1792);
and U1221 (N_1221,In_18,In_277);
nor U1222 (N_1222,In_1710,In_2325);
and U1223 (N_1223,In_2176,In_1271);
and U1224 (N_1224,In_483,In_1448);
xor U1225 (N_1225,In_2417,In_2365);
nand U1226 (N_1226,In_2288,In_2050);
and U1227 (N_1227,In_699,In_1068);
nand U1228 (N_1228,In_1634,In_543);
and U1229 (N_1229,In_2488,In_825);
and U1230 (N_1230,In_1283,In_2444);
nor U1231 (N_1231,In_141,In_270);
or U1232 (N_1232,In_1165,In_1620);
nor U1233 (N_1233,In_1000,In_583);
nand U1234 (N_1234,In_266,In_1563);
and U1235 (N_1235,In_903,In_2136);
xnor U1236 (N_1236,In_2204,In_1086);
nor U1237 (N_1237,In_1943,In_820);
or U1238 (N_1238,In_225,In_156);
or U1239 (N_1239,In_641,In_2010);
or U1240 (N_1240,In_235,In_1040);
xor U1241 (N_1241,In_2286,In_2305);
and U1242 (N_1242,In_961,In_1573);
nand U1243 (N_1243,In_2205,In_1637);
nor U1244 (N_1244,In_302,In_1457);
and U1245 (N_1245,In_1503,In_1322);
nand U1246 (N_1246,In_2430,In_928);
or U1247 (N_1247,In_2302,In_569);
xor U1248 (N_1248,In_746,In_1570);
or U1249 (N_1249,In_312,In_2304);
xnor U1250 (N_1250,In_1344,In_465);
nor U1251 (N_1251,In_2208,In_913);
and U1252 (N_1252,In_2248,In_959);
nand U1253 (N_1253,In_1410,In_1357);
and U1254 (N_1254,In_1366,In_404);
nor U1255 (N_1255,In_1314,In_1174);
nand U1256 (N_1256,In_1966,In_104);
nor U1257 (N_1257,In_1140,In_90);
and U1258 (N_1258,In_1508,In_2446);
or U1259 (N_1259,In_729,In_1407);
nor U1260 (N_1260,In_855,In_2255);
and U1261 (N_1261,In_618,In_655);
or U1262 (N_1262,In_649,In_2201);
nor U1263 (N_1263,In_616,In_2025);
xnor U1264 (N_1264,In_155,In_15);
xnor U1265 (N_1265,In_835,In_731);
or U1266 (N_1266,In_80,In_2343);
or U1267 (N_1267,In_1285,In_106);
nand U1268 (N_1268,In_1541,In_1416);
nor U1269 (N_1269,In_1095,In_599);
and U1270 (N_1270,In_1532,In_767);
or U1271 (N_1271,In_424,In_2049);
nor U1272 (N_1272,In_2166,In_370);
nand U1273 (N_1273,In_190,In_892);
nand U1274 (N_1274,In_510,In_2158);
and U1275 (N_1275,In_2011,In_844);
or U1276 (N_1276,In_1807,In_232);
or U1277 (N_1277,In_75,In_1561);
and U1278 (N_1278,In_1842,In_2129);
nor U1279 (N_1279,In_2136,In_1137);
xnor U1280 (N_1280,In_913,In_2368);
nand U1281 (N_1281,In_1261,In_2071);
and U1282 (N_1282,In_2172,In_1068);
nor U1283 (N_1283,In_429,In_1268);
nor U1284 (N_1284,In_47,In_1446);
nand U1285 (N_1285,In_637,In_1154);
xor U1286 (N_1286,In_1289,In_725);
nand U1287 (N_1287,In_1697,In_1047);
xnor U1288 (N_1288,In_2042,In_181);
or U1289 (N_1289,In_2486,In_2366);
nand U1290 (N_1290,In_1665,In_2307);
nor U1291 (N_1291,In_1537,In_917);
nand U1292 (N_1292,In_782,In_336);
and U1293 (N_1293,In_577,In_2309);
xor U1294 (N_1294,In_475,In_1145);
and U1295 (N_1295,In_1991,In_2214);
or U1296 (N_1296,In_1347,In_933);
and U1297 (N_1297,In_1688,In_2063);
or U1298 (N_1298,In_2142,In_1433);
nand U1299 (N_1299,In_1686,In_1312);
nand U1300 (N_1300,In_264,In_1389);
nor U1301 (N_1301,In_2143,In_1041);
and U1302 (N_1302,In_1725,In_2022);
and U1303 (N_1303,In_2083,In_2037);
nor U1304 (N_1304,In_1294,In_1581);
nor U1305 (N_1305,In_243,In_2479);
nand U1306 (N_1306,In_1578,In_1082);
nand U1307 (N_1307,In_1957,In_221);
xor U1308 (N_1308,In_183,In_733);
nand U1309 (N_1309,In_129,In_551);
nor U1310 (N_1310,In_2171,In_1989);
or U1311 (N_1311,In_1627,In_175);
or U1312 (N_1312,In_2254,In_1555);
nand U1313 (N_1313,In_2328,In_1416);
and U1314 (N_1314,In_846,In_563);
or U1315 (N_1315,In_427,In_2056);
nand U1316 (N_1316,In_1507,In_692);
or U1317 (N_1317,In_1789,In_1214);
nor U1318 (N_1318,In_1370,In_1160);
and U1319 (N_1319,In_589,In_900);
or U1320 (N_1320,In_1101,In_818);
and U1321 (N_1321,In_1066,In_1970);
and U1322 (N_1322,In_2141,In_2365);
xnor U1323 (N_1323,In_937,In_140);
xor U1324 (N_1324,In_1339,In_1729);
or U1325 (N_1325,In_871,In_305);
xnor U1326 (N_1326,In_135,In_1473);
nor U1327 (N_1327,In_408,In_1829);
or U1328 (N_1328,In_1695,In_1558);
nand U1329 (N_1329,In_804,In_1135);
and U1330 (N_1330,In_1288,In_93);
nand U1331 (N_1331,In_510,In_847);
nor U1332 (N_1332,In_1947,In_1100);
nor U1333 (N_1333,In_172,In_2209);
nand U1334 (N_1334,In_1654,In_2151);
nand U1335 (N_1335,In_267,In_1999);
xnor U1336 (N_1336,In_203,In_2306);
xnor U1337 (N_1337,In_234,In_1883);
nor U1338 (N_1338,In_52,In_2428);
and U1339 (N_1339,In_1784,In_401);
nand U1340 (N_1340,In_819,In_1985);
nand U1341 (N_1341,In_1824,In_335);
nand U1342 (N_1342,In_2166,In_1399);
xnor U1343 (N_1343,In_1901,In_1476);
or U1344 (N_1344,In_2256,In_1141);
or U1345 (N_1345,In_414,In_480);
or U1346 (N_1346,In_674,In_775);
nand U1347 (N_1347,In_578,In_2250);
or U1348 (N_1348,In_334,In_1989);
nor U1349 (N_1349,In_2233,In_827);
nand U1350 (N_1350,In_1708,In_1455);
and U1351 (N_1351,In_975,In_1000);
or U1352 (N_1352,In_343,In_736);
xnor U1353 (N_1353,In_1256,In_1094);
nor U1354 (N_1354,In_1339,In_27);
xnor U1355 (N_1355,In_2255,In_1561);
nor U1356 (N_1356,In_3,In_1444);
and U1357 (N_1357,In_1936,In_2161);
nor U1358 (N_1358,In_1386,In_805);
nor U1359 (N_1359,In_115,In_2093);
and U1360 (N_1360,In_1096,In_2034);
and U1361 (N_1361,In_2407,In_2498);
xnor U1362 (N_1362,In_855,In_2211);
nor U1363 (N_1363,In_207,In_651);
nor U1364 (N_1364,In_1109,In_1322);
xor U1365 (N_1365,In_2107,In_1687);
and U1366 (N_1366,In_1262,In_1823);
xnor U1367 (N_1367,In_2496,In_2303);
and U1368 (N_1368,In_1199,In_16);
or U1369 (N_1369,In_1511,In_780);
xor U1370 (N_1370,In_650,In_67);
or U1371 (N_1371,In_171,In_938);
nor U1372 (N_1372,In_26,In_253);
or U1373 (N_1373,In_2438,In_1193);
xnor U1374 (N_1374,In_2320,In_2430);
or U1375 (N_1375,In_845,In_2424);
or U1376 (N_1376,In_1253,In_1093);
and U1377 (N_1377,In_2110,In_959);
nand U1378 (N_1378,In_835,In_2210);
nor U1379 (N_1379,In_57,In_244);
nand U1380 (N_1380,In_1617,In_1847);
nor U1381 (N_1381,In_401,In_741);
xor U1382 (N_1382,In_592,In_1831);
or U1383 (N_1383,In_769,In_336);
and U1384 (N_1384,In_636,In_788);
and U1385 (N_1385,In_98,In_1521);
nand U1386 (N_1386,In_482,In_1239);
and U1387 (N_1387,In_1572,In_1021);
xor U1388 (N_1388,In_212,In_720);
nand U1389 (N_1389,In_2143,In_680);
xor U1390 (N_1390,In_1010,In_1657);
xor U1391 (N_1391,In_1756,In_1214);
and U1392 (N_1392,In_1787,In_87);
nor U1393 (N_1393,In_956,In_111);
nor U1394 (N_1394,In_1590,In_1542);
or U1395 (N_1395,In_1884,In_1917);
nand U1396 (N_1396,In_2001,In_2085);
nand U1397 (N_1397,In_2086,In_706);
or U1398 (N_1398,In_833,In_1336);
and U1399 (N_1399,In_1793,In_32);
nor U1400 (N_1400,In_486,In_2226);
and U1401 (N_1401,In_1051,In_1605);
nand U1402 (N_1402,In_1727,In_1335);
nor U1403 (N_1403,In_775,In_1520);
xor U1404 (N_1404,In_2384,In_1674);
or U1405 (N_1405,In_2135,In_1397);
or U1406 (N_1406,In_1453,In_822);
and U1407 (N_1407,In_272,In_2189);
or U1408 (N_1408,In_1101,In_1091);
and U1409 (N_1409,In_66,In_1619);
xor U1410 (N_1410,In_2251,In_417);
nand U1411 (N_1411,In_216,In_112);
and U1412 (N_1412,In_931,In_2105);
and U1413 (N_1413,In_2340,In_2475);
and U1414 (N_1414,In_1756,In_2276);
and U1415 (N_1415,In_1195,In_443);
or U1416 (N_1416,In_445,In_832);
nor U1417 (N_1417,In_1667,In_1220);
nor U1418 (N_1418,In_681,In_501);
nand U1419 (N_1419,In_1724,In_2049);
and U1420 (N_1420,In_941,In_1028);
nand U1421 (N_1421,In_504,In_954);
and U1422 (N_1422,In_83,In_2085);
and U1423 (N_1423,In_2392,In_1978);
or U1424 (N_1424,In_1466,In_1598);
nor U1425 (N_1425,In_97,In_440);
xor U1426 (N_1426,In_1181,In_2043);
nor U1427 (N_1427,In_731,In_1602);
nor U1428 (N_1428,In_1948,In_2286);
nand U1429 (N_1429,In_1380,In_1370);
or U1430 (N_1430,In_763,In_1091);
nor U1431 (N_1431,In_2196,In_2278);
or U1432 (N_1432,In_2274,In_1431);
nand U1433 (N_1433,In_487,In_560);
nand U1434 (N_1434,In_1362,In_1465);
nand U1435 (N_1435,In_2098,In_362);
nor U1436 (N_1436,In_1413,In_1552);
nor U1437 (N_1437,In_1246,In_141);
xnor U1438 (N_1438,In_12,In_289);
nand U1439 (N_1439,In_1113,In_343);
and U1440 (N_1440,In_306,In_492);
xnor U1441 (N_1441,In_1206,In_1510);
nor U1442 (N_1442,In_1629,In_1787);
nor U1443 (N_1443,In_619,In_1073);
nor U1444 (N_1444,In_200,In_705);
nor U1445 (N_1445,In_1345,In_140);
or U1446 (N_1446,In_353,In_925);
and U1447 (N_1447,In_1497,In_300);
nor U1448 (N_1448,In_1672,In_15);
or U1449 (N_1449,In_2249,In_2161);
or U1450 (N_1450,In_934,In_2242);
nor U1451 (N_1451,In_1422,In_1409);
and U1452 (N_1452,In_793,In_13);
nand U1453 (N_1453,In_244,In_313);
and U1454 (N_1454,In_1636,In_563);
nand U1455 (N_1455,In_1836,In_806);
xnor U1456 (N_1456,In_1385,In_678);
nand U1457 (N_1457,In_742,In_2352);
nand U1458 (N_1458,In_1889,In_1336);
nor U1459 (N_1459,In_749,In_1554);
and U1460 (N_1460,In_1046,In_2495);
and U1461 (N_1461,In_1676,In_1736);
or U1462 (N_1462,In_979,In_1561);
and U1463 (N_1463,In_1826,In_1271);
nand U1464 (N_1464,In_332,In_921);
nor U1465 (N_1465,In_1583,In_587);
nor U1466 (N_1466,In_1476,In_1435);
or U1467 (N_1467,In_101,In_1179);
nand U1468 (N_1468,In_48,In_720);
xnor U1469 (N_1469,In_1974,In_2169);
xor U1470 (N_1470,In_1918,In_1162);
or U1471 (N_1471,In_1478,In_2113);
and U1472 (N_1472,In_840,In_755);
or U1473 (N_1473,In_763,In_789);
and U1474 (N_1474,In_2446,In_908);
or U1475 (N_1475,In_923,In_1716);
nor U1476 (N_1476,In_976,In_841);
nor U1477 (N_1477,In_467,In_1940);
and U1478 (N_1478,In_1325,In_2272);
nand U1479 (N_1479,In_1666,In_1684);
or U1480 (N_1480,In_1705,In_1129);
or U1481 (N_1481,In_2392,In_2438);
and U1482 (N_1482,In_1191,In_1859);
xnor U1483 (N_1483,In_1353,In_1624);
nand U1484 (N_1484,In_1905,In_1110);
xor U1485 (N_1485,In_1504,In_1907);
and U1486 (N_1486,In_422,In_2491);
and U1487 (N_1487,In_1356,In_2056);
or U1488 (N_1488,In_1447,In_139);
or U1489 (N_1489,In_1220,In_133);
and U1490 (N_1490,In_636,In_1750);
and U1491 (N_1491,In_1909,In_2048);
and U1492 (N_1492,In_1811,In_19);
or U1493 (N_1493,In_434,In_1830);
xor U1494 (N_1494,In_668,In_392);
nor U1495 (N_1495,In_2377,In_2040);
xnor U1496 (N_1496,In_20,In_255);
nor U1497 (N_1497,In_1972,In_907);
nor U1498 (N_1498,In_15,In_255);
nor U1499 (N_1499,In_2218,In_156);
nor U1500 (N_1500,In_235,In_912);
nand U1501 (N_1501,In_1015,In_67);
xnor U1502 (N_1502,In_2445,In_711);
nand U1503 (N_1503,In_206,In_829);
nand U1504 (N_1504,In_2493,In_1926);
or U1505 (N_1505,In_744,In_1579);
and U1506 (N_1506,In_2284,In_2329);
xnor U1507 (N_1507,In_1935,In_1286);
xor U1508 (N_1508,In_620,In_948);
nor U1509 (N_1509,In_1486,In_2003);
xnor U1510 (N_1510,In_1845,In_247);
and U1511 (N_1511,In_2013,In_2177);
nand U1512 (N_1512,In_1361,In_1524);
nor U1513 (N_1513,In_316,In_581);
nand U1514 (N_1514,In_2496,In_1084);
nand U1515 (N_1515,In_626,In_769);
and U1516 (N_1516,In_2428,In_583);
or U1517 (N_1517,In_1129,In_825);
xor U1518 (N_1518,In_874,In_1248);
or U1519 (N_1519,In_1540,In_1633);
nor U1520 (N_1520,In_2011,In_347);
xor U1521 (N_1521,In_1201,In_2379);
xnor U1522 (N_1522,In_311,In_1847);
or U1523 (N_1523,In_742,In_657);
or U1524 (N_1524,In_181,In_1555);
or U1525 (N_1525,In_1459,In_1225);
nand U1526 (N_1526,In_1261,In_2078);
nand U1527 (N_1527,In_2225,In_1108);
and U1528 (N_1528,In_2170,In_1823);
nor U1529 (N_1529,In_89,In_1991);
and U1530 (N_1530,In_1192,In_1920);
xnor U1531 (N_1531,In_129,In_1034);
xor U1532 (N_1532,In_973,In_1076);
and U1533 (N_1533,In_1634,In_2203);
xnor U1534 (N_1534,In_791,In_1810);
and U1535 (N_1535,In_1009,In_1662);
nor U1536 (N_1536,In_683,In_2104);
or U1537 (N_1537,In_604,In_1540);
or U1538 (N_1538,In_1450,In_1258);
and U1539 (N_1539,In_2484,In_2416);
nand U1540 (N_1540,In_2023,In_1970);
xor U1541 (N_1541,In_1418,In_2254);
and U1542 (N_1542,In_696,In_1277);
or U1543 (N_1543,In_36,In_1388);
and U1544 (N_1544,In_380,In_2259);
xor U1545 (N_1545,In_1753,In_1886);
nand U1546 (N_1546,In_1013,In_948);
and U1547 (N_1547,In_1423,In_331);
nand U1548 (N_1548,In_515,In_642);
or U1549 (N_1549,In_2272,In_1792);
nor U1550 (N_1550,In_36,In_1234);
nand U1551 (N_1551,In_914,In_583);
and U1552 (N_1552,In_356,In_1052);
nor U1553 (N_1553,In_966,In_1775);
nor U1554 (N_1554,In_156,In_2069);
nor U1555 (N_1555,In_1349,In_1449);
xnor U1556 (N_1556,In_122,In_43);
nor U1557 (N_1557,In_525,In_2322);
xor U1558 (N_1558,In_612,In_1409);
nand U1559 (N_1559,In_1130,In_1420);
and U1560 (N_1560,In_1255,In_1923);
or U1561 (N_1561,In_879,In_2261);
nand U1562 (N_1562,In_246,In_1845);
nand U1563 (N_1563,In_910,In_1993);
nand U1564 (N_1564,In_1468,In_2110);
nor U1565 (N_1565,In_627,In_773);
or U1566 (N_1566,In_960,In_1680);
nor U1567 (N_1567,In_674,In_339);
nor U1568 (N_1568,In_1764,In_2190);
nand U1569 (N_1569,In_359,In_46);
and U1570 (N_1570,In_827,In_1207);
or U1571 (N_1571,In_1450,In_317);
nand U1572 (N_1572,In_1833,In_1331);
nor U1573 (N_1573,In_1324,In_1042);
nor U1574 (N_1574,In_1037,In_959);
or U1575 (N_1575,In_524,In_1395);
and U1576 (N_1576,In_630,In_2148);
xor U1577 (N_1577,In_1825,In_2060);
or U1578 (N_1578,In_1374,In_1480);
nor U1579 (N_1579,In_1236,In_1133);
xor U1580 (N_1580,In_1025,In_1091);
nand U1581 (N_1581,In_766,In_1979);
xor U1582 (N_1582,In_1516,In_761);
and U1583 (N_1583,In_216,In_1777);
nor U1584 (N_1584,In_46,In_744);
xnor U1585 (N_1585,In_790,In_2096);
or U1586 (N_1586,In_969,In_1044);
or U1587 (N_1587,In_742,In_1742);
nand U1588 (N_1588,In_2042,In_986);
nor U1589 (N_1589,In_2457,In_83);
nand U1590 (N_1590,In_2339,In_1439);
nor U1591 (N_1591,In_2412,In_1657);
nor U1592 (N_1592,In_1368,In_1334);
xnor U1593 (N_1593,In_1373,In_3);
nand U1594 (N_1594,In_674,In_925);
or U1595 (N_1595,In_117,In_249);
or U1596 (N_1596,In_24,In_1712);
nor U1597 (N_1597,In_52,In_1417);
xnor U1598 (N_1598,In_2097,In_1793);
and U1599 (N_1599,In_2274,In_1108);
xnor U1600 (N_1600,In_419,In_2236);
nand U1601 (N_1601,In_1892,In_9);
and U1602 (N_1602,In_378,In_2234);
and U1603 (N_1603,In_439,In_743);
nor U1604 (N_1604,In_77,In_101);
nand U1605 (N_1605,In_1811,In_1911);
nor U1606 (N_1606,In_2211,In_2499);
xor U1607 (N_1607,In_2316,In_581);
nor U1608 (N_1608,In_1481,In_1677);
and U1609 (N_1609,In_1548,In_2037);
and U1610 (N_1610,In_1000,In_1619);
or U1611 (N_1611,In_344,In_2163);
xnor U1612 (N_1612,In_1198,In_1178);
nor U1613 (N_1613,In_2133,In_286);
nor U1614 (N_1614,In_3,In_975);
nor U1615 (N_1615,In_717,In_2170);
or U1616 (N_1616,In_2261,In_2157);
xnor U1617 (N_1617,In_1826,In_498);
or U1618 (N_1618,In_1327,In_1416);
nor U1619 (N_1619,In_1552,In_117);
and U1620 (N_1620,In_862,In_1761);
nand U1621 (N_1621,In_1126,In_1320);
or U1622 (N_1622,In_252,In_2386);
xor U1623 (N_1623,In_685,In_634);
and U1624 (N_1624,In_715,In_1630);
xor U1625 (N_1625,In_1710,In_937);
or U1626 (N_1626,In_1384,In_2107);
or U1627 (N_1627,In_1383,In_499);
nand U1628 (N_1628,In_2003,In_2363);
nor U1629 (N_1629,In_1379,In_393);
nor U1630 (N_1630,In_2435,In_668);
or U1631 (N_1631,In_84,In_1419);
or U1632 (N_1632,In_2002,In_515);
xnor U1633 (N_1633,In_810,In_2369);
nand U1634 (N_1634,In_2386,In_1485);
xor U1635 (N_1635,In_1903,In_399);
xnor U1636 (N_1636,In_1495,In_402);
and U1637 (N_1637,In_1058,In_170);
and U1638 (N_1638,In_280,In_1635);
xor U1639 (N_1639,In_758,In_642);
and U1640 (N_1640,In_1224,In_778);
and U1641 (N_1641,In_943,In_226);
xor U1642 (N_1642,In_1941,In_2221);
or U1643 (N_1643,In_112,In_538);
or U1644 (N_1644,In_1193,In_860);
nand U1645 (N_1645,In_2028,In_1691);
nand U1646 (N_1646,In_1569,In_1327);
and U1647 (N_1647,In_149,In_1004);
xnor U1648 (N_1648,In_2483,In_1537);
nand U1649 (N_1649,In_1671,In_870);
or U1650 (N_1650,In_1806,In_2225);
nand U1651 (N_1651,In_546,In_1300);
and U1652 (N_1652,In_1444,In_737);
and U1653 (N_1653,In_291,In_1274);
nand U1654 (N_1654,In_1155,In_1585);
or U1655 (N_1655,In_92,In_1876);
xnor U1656 (N_1656,In_1487,In_573);
xnor U1657 (N_1657,In_231,In_233);
nand U1658 (N_1658,In_946,In_245);
xnor U1659 (N_1659,In_1963,In_2322);
or U1660 (N_1660,In_1022,In_2371);
or U1661 (N_1661,In_1608,In_463);
nand U1662 (N_1662,In_260,In_2071);
and U1663 (N_1663,In_1967,In_2291);
or U1664 (N_1664,In_192,In_1167);
or U1665 (N_1665,In_2031,In_1526);
or U1666 (N_1666,In_868,In_2232);
nand U1667 (N_1667,In_1650,In_2220);
nand U1668 (N_1668,In_2017,In_226);
and U1669 (N_1669,In_512,In_1730);
and U1670 (N_1670,In_76,In_1931);
or U1671 (N_1671,In_2375,In_269);
xnor U1672 (N_1672,In_57,In_1732);
or U1673 (N_1673,In_2443,In_1697);
xor U1674 (N_1674,In_1383,In_454);
nor U1675 (N_1675,In_1032,In_1951);
xor U1676 (N_1676,In_1117,In_840);
xnor U1677 (N_1677,In_2028,In_1960);
nand U1678 (N_1678,In_1238,In_1627);
or U1679 (N_1679,In_2491,In_685);
or U1680 (N_1680,In_2090,In_927);
and U1681 (N_1681,In_1641,In_1325);
xor U1682 (N_1682,In_1600,In_444);
nor U1683 (N_1683,In_1242,In_1305);
nand U1684 (N_1684,In_965,In_2127);
xnor U1685 (N_1685,In_2128,In_999);
or U1686 (N_1686,In_1806,In_2329);
nand U1687 (N_1687,In_1082,In_538);
and U1688 (N_1688,In_2175,In_903);
and U1689 (N_1689,In_360,In_1434);
nor U1690 (N_1690,In_165,In_375);
or U1691 (N_1691,In_756,In_2387);
nand U1692 (N_1692,In_1091,In_1667);
nand U1693 (N_1693,In_2399,In_1977);
nand U1694 (N_1694,In_2299,In_834);
or U1695 (N_1695,In_1729,In_819);
xnor U1696 (N_1696,In_365,In_98);
nand U1697 (N_1697,In_1457,In_554);
and U1698 (N_1698,In_2103,In_1885);
and U1699 (N_1699,In_1920,In_1898);
xnor U1700 (N_1700,In_1332,In_127);
xor U1701 (N_1701,In_2392,In_2149);
or U1702 (N_1702,In_542,In_2067);
and U1703 (N_1703,In_1634,In_515);
and U1704 (N_1704,In_2137,In_1969);
nand U1705 (N_1705,In_1023,In_226);
and U1706 (N_1706,In_576,In_437);
nor U1707 (N_1707,In_2332,In_2461);
nor U1708 (N_1708,In_1268,In_2389);
nor U1709 (N_1709,In_2140,In_1804);
xor U1710 (N_1710,In_1996,In_1696);
or U1711 (N_1711,In_647,In_1815);
nor U1712 (N_1712,In_1259,In_2282);
or U1713 (N_1713,In_609,In_2141);
and U1714 (N_1714,In_1673,In_1206);
or U1715 (N_1715,In_2491,In_238);
nand U1716 (N_1716,In_1846,In_541);
nand U1717 (N_1717,In_1232,In_295);
nand U1718 (N_1718,In_502,In_2317);
nand U1719 (N_1719,In_2023,In_1844);
xor U1720 (N_1720,In_1781,In_788);
xor U1721 (N_1721,In_35,In_2049);
and U1722 (N_1722,In_327,In_8);
nor U1723 (N_1723,In_2139,In_767);
xor U1724 (N_1724,In_1671,In_1791);
and U1725 (N_1725,In_1728,In_1173);
or U1726 (N_1726,In_74,In_490);
nand U1727 (N_1727,In_835,In_1476);
or U1728 (N_1728,In_1061,In_1889);
and U1729 (N_1729,In_1990,In_1672);
or U1730 (N_1730,In_1965,In_676);
nor U1731 (N_1731,In_529,In_2189);
nand U1732 (N_1732,In_2496,In_2049);
and U1733 (N_1733,In_1289,In_560);
xor U1734 (N_1734,In_1125,In_1777);
nand U1735 (N_1735,In_1652,In_686);
xor U1736 (N_1736,In_290,In_909);
or U1737 (N_1737,In_1912,In_2138);
nor U1738 (N_1738,In_1066,In_2229);
or U1739 (N_1739,In_1809,In_1041);
nor U1740 (N_1740,In_566,In_334);
xnor U1741 (N_1741,In_2411,In_329);
nor U1742 (N_1742,In_1283,In_988);
xor U1743 (N_1743,In_1234,In_1443);
nand U1744 (N_1744,In_489,In_2015);
nor U1745 (N_1745,In_1946,In_758);
nand U1746 (N_1746,In_2333,In_1069);
and U1747 (N_1747,In_1007,In_860);
or U1748 (N_1748,In_523,In_80);
nor U1749 (N_1749,In_430,In_1267);
xnor U1750 (N_1750,In_1926,In_1735);
nor U1751 (N_1751,In_1843,In_2055);
or U1752 (N_1752,In_111,In_1854);
nor U1753 (N_1753,In_981,In_386);
nand U1754 (N_1754,In_2022,In_774);
nand U1755 (N_1755,In_1092,In_2147);
and U1756 (N_1756,In_1087,In_2385);
or U1757 (N_1757,In_1895,In_617);
and U1758 (N_1758,In_222,In_15);
nor U1759 (N_1759,In_1070,In_832);
and U1760 (N_1760,In_1469,In_1485);
nand U1761 (N_1761,In_431,In_573);
nand U1762 (N_1762,In_700,In_2402);
nor U1763 (N_1763,In_633,In_1572);
and U1764 (N_1764,In_1660,In_1959);
nor U1765 (N_1765,In_859,In_2129);
or U1766 (N_1766,In_206,In_823);
xor U1767 (N_1767,In_2458,In_2304);
nor U1768 (N_1768,In_2089,In_2414);
and U1769 (N_1769,In_2422,In_149);
nor U1770 (N_1770,In_1491,In_1851);
or U1771 (N_1771,In_22,In_1682);
or U1772 (N_1772,In_362,In_1022);
or U1773 (N_1773,In_1395,In_24);
nor U1774 (N_1774,In_2170,In_753);
xor U1775 (N_1775,In_952,In_1696);
and U1776 (N_1776,In_2133,In_2124);
and U1777 (N_1777,In_156,In_1960);
nand U1778 (N_1778,In_2489,In_38);
or U1779 (N_1779,In_1528,In_1445);
or U1780 (N_1780,In_192,In_2339);
nor U1781 (N_1781,In_734,In_350);
xor U1782 (N_1782,In_939,In_2466);
nand U1783 (N_1783,In_275,In_2464);
nor U1784 (N_1784,In_2260,In_2286);
nor U1785 (N_1785,In_329,In_1281);
xnor U1786 (N_1786,In_470,In_39);
and U1787 (N_1787,In_274,In_2187);
or U1788 (N_1788,In_1692,In_629);
and U1789 (N_1789,In_887,In_2308);
xor U1790 (N_1790,In_2125,In_935);
or U1791 (N_1791,In_1452,In_2302);
nor U1792 (N_1792,In_538,In_692);
and U1793 (N_1793,In_2431,In_1719);
xnor U1794 (N_1794,In_784,In_1589);
or U1795 (N_1795,In_2135,In_1785);
nand U1796 (N_1796,In_1473,In_1358);
or U1797 (N_1797,In_909,In_109);
xnor U1798 (N_1798,In_1709,In_1890);
nand U1799 (N_1799,In_851,In_2238);
or U1800 (N_1800,In_2074,In_713);
or U1801 (N_1801,In_805,In_104);
nand U1802 (N_1802,In_461,In_115);
nand U1803 (N_1803,In_480,In_1000);
xor U1804 (N_1804,In_54,In_207);
or U1805 (N_1805,In_1296,In_1624);
and U1806 (N_1806,In_217,In_1594);
xnor U1807 (N_1807,In_1181,In_1429);
nand U1808 (N_1808,In_577,In_1107);
or U1809 (N_1809,In_893,In_1526);
nand U1810 (N_1810,In_1915,In_1029);
nand U1811 (N_1811,In_18,In_2234);
or U1812 (N_1812,In_2209,In_1024);
nand U1813 (N_1813,In_2029,In_2424);
or U1814 (N_1814,In_1958,In_2414);
and U1815 (N_1815,In_2468,In_1425);
nor U1816 (N_1816,In_1006,In_1322);
and U1817 (N_1817,In_1890,In_2370);
or U1818 (N_1818,In_1785,In_1662);
nand U1819 (N_1819,In_1939,In_273);
and U1820 (N_1820,In_2429,In_1703);
xor U1821 (N_1821,In_2126,In_274);
nand U1822 (N_1822,In_1448,In_71);
nand U1823 (N_1823,In_1316,In_1025);
nor U1824 (N_1824,In_1946,In_1052);
nor U1825 (N_1825,In_713,In_1586);
nand U1826 (N_1826,In_152,In_563);
nor U1827 (N_1827,In_1745,In_891);
nor U1828 (N_1828,In_524,In_410);
nand U1829 (N_1829,In_2201,In_1598);
nand U1830 (N_1830,In_1476,In_2085);
nor U1831 (N_1831,In_1621,In_397);
xor U1832 (N_1832,In_2262,In_2028);
nor U1833 (N_1833,In_341,In_1391);
or U1834 (N_1834,In_1998,In_1182);
and U1835 (N_1835,In_170,In_247);
or U1836 (N_1836,In_1233,In_2027);
nor U1837 (N_1837,In_512,In_1713);
nand U1838 (N_1838,In_1570,In_2242);
or U1839 (N_1839,In_868,In_1789);
nand U1840 (N_1840,In_1610,In_843);
xor U1841 (N_1841,In_1058,In_1697);
xnor U1842 (N_1842,In_624,In_1555);
nor U1843 (N_1843,In_2280,In_1573);
nor U1844 (N_1844,In_160,In_2318);
or U1845 (N_1845,In_525,In_1660);
and U1846 (N_1846,In_258,In_205);
nor U1847 (N_1847,In_702,In_1524);
or U1848 (N_1848,In_154,In_1339);
xnor U1849 (N_1849,In_1296,In_1203);
and U1850 (N_1850,In_473,In_1688);
xor U1851 (N_1851,In_1496,In_614);
and U1852 (N_1852,In_1231,In_347);
or U1853 (N_1853,In_249,In_2427);
nand U1854 (N_1854,In_1964,In_829);
xor U1855 (N_1855,In_111,In_211);
xor U1856 (N_1856,In_1198,In_2251);
nor U1857 (N_1857,In_952,In_2463);
xor U1858 (N_1858,In_812,In_2156);
xnor U1859 (N_1859,In_2433,In_1053);
and U1860 (N_1860,In_2463,In_1951);
and U1861 (N_1861,In_181,In_1068);
and U1862 (N_1862,In_1620,In_2200);
nand U1863 (N_1863,In_2023,In_2486);
xor U1864 (N_1864,In_947,In_1376);
xnor U1865 (N_1865,In_941,In_1620);
nand U1866 (N_1866,In_1650,In_2021);
or U1867 (N_1867,In_1191,In_2422);
and U1868 (N_1868,In_1044,In_544);
xnor U1869 (N_1869,In_905,In_2099);
nand U1870 (N_1870,In_1224,In_376);
or U1871 (N_1871,In_229,In_632);
xor U1872 (N_1872,In_330,In_609);
xor U1873 (N_1873,In_108,In_809);
nand U1874 (N_1874,In_616,In_737);
and U1875 (N_1875,In_806,In_2347);
xnor U1876 (N_1876,In_332,In_405);
nand U1877 (N_1877,In_678,In_609);
and U1878 (N_1878,In_1049,In_499);
xnor U1879 (N_1879,In_2038,In_947);
xor U1880 (N_1880,In_1123,In_968);
or U1881 (N_1881,In_1439,In_1229);
nand U1882 (N_1882,In_1707,In_1198);
or U1883 (N_1883,In_192,In_1510);
xnor U1884 (N_1884,In_1652,In_1159);
xor U1885 (N_1885,In_1111,In_1038);
nand U1886 (N_1886,In_249,In_257);
and U1887 (N_1887,In_118,In_928);
nor U1888 (N_1888,In_2211,In_1835);
nand U1889 (N_1889,In_717,In_1059);
and U1890 (N_1890,In_172,In_550);
nand U1891 (N_1891,In_2442,In_281);
nor U1892 (N_1892,In_2384,In_2155);
nor U1893 (N_1893,In_1262,In_279);
xnor U1894 (N_1894,In_235,In_1774);
nand U1895 (N_1895,In_239,In_2041);
nand U1896 (N_1896,In_1941,In_1572);
nand U1897 (N_1897,In_2424,In_1344);
xnor U1898 (N_1898,In_1303,In_2360);
xnor U1899 (N_1899,In_2429,In_1209);
or U1900 (N_1900,In_768,In_2051);
xnor U1901 (N_1901,In_1289,In_409);
and U1902 (N_1902,In_857,In_727);
and U1903 (N_1903,In_2178,In_2257);
xnor U1904 (N_1904,In_1386,In_1753);
and U1905 (N_1905,In_1531,In_174);
and U1906 (N_1906,In_1580,In_1742);
xor U1907 (N_1907,In_1150,In_1912);
and U1908 (N_1908,In_359,In_740);
and U1909 (N_1909,In_1524,In_1597);
or U1910 (N_1910,In_1894,In_37);
or U1911 (N_1911,In_1816,In_1330);
and U1912 (N_1912,In_888,In_1894);
xor U1913 (N_1913,In_2147,In_936);
and U1914 (N_1914,In_856,In_1445);
nand U1915 (N_1915,In_1126,In_1124);
or U1916 (N_1916,In_2039,In_1697);
or U1917 (N_1917,In_1345,In_644);
or U1918 (N_1918,In_720,In_2092);
and U1919 (N_1919,In_1761,In_2245);
nand U1920 (N_1920,In_38,In_1795);
nor U1921 (N_1921,In_2122,In_1175);
nor U1922 (N_1922,In_629,In_1886);
xor U1923 (N_1923,In_502,In_358);
xnor U1924 (N_1924,In_2044,In_1503);
and U1925 (N_1925,In_1529,In_2167);
nand U1926 (N_1926,In_90,In_449);
or U1927 (N_1927,In_1644,In_0);
nand U1928 (N_1928,In_1184,In_1562);
and U1929 (N_1929,In_328,In_472);
nor U1930 (N_1930,In_2362,In_2036);
xor U1931 (N_1931,In_680,In_360);
and U1932 (N_1932,In_1676,In_816);
and U1933 (N_1933,In_2144,In_2409);
nand U1934 (N_1934,In_2370,In_1853);
nand U1935 (N_1935,In_273,In_1465);
xor U1936 (N_1936,In_1242,In_1080);
or U1937 (N_1937,In_1333,In_824);
or U1938 (N_1938,In_638,In_2395);
nand U1939 (N_1939,In_1397,In_1720);
nand U1940 (N_1940,In_1763,In_2134);
nor U1941 (N_1941,In_744,In_725);
nand U1942 (N_1942,In_1273,In_1888);
and U1943 (N_1943,In_1081,In_2191);
xor U1944 (N_1944,In_248,In_433);
nand U1945 (N_1945,In_1277,In_1571);
and U1946 (N_1946,In_2090,In_202);
or U1947 (N_1947,In_661,In_432);
nand U1948 (N_1948,In_906,In_346);
xor U1949 (N_1949,In_2286,In_768);
and U1950 (N_1950,In_1521,In_9);
or U1951 (N_1951,In_2466,In_1849);
xnor U1952 (N_1952,In_2496,In_2050);
or U1953 (N_1953,In_805,In_1948);
xnor U1954 (N_1954,In_1801,In_439);
and U1955 (N_1955,In_557,In_2318);
nor U1956 (N_1956,In_2413,In_1239);
nor U1957 (N_1957,In_701,In_1348);
and U1958 (N_1958,In_1665,In_2091);
nand U1959 (N_1959,In_816,In_1389);
and U1960 (N_1960,In_239,In_633);
xor U1961 (N_1961,In_616,In_812);
nand U1962 (N_1962,In_1448,In_1796);
nand U1963 (N_1963,In_1530,In_535);
or U1964 (N_1964,In_369,In_1182);
xnor U1965 (N_1965,In_335,In_2038);
and U1966 (N_1966,In_548,In_1829);
and U1967 (N_1967,In_2253,In_1796);
nand U1968 (N_1968,In_1750,In_961);
or U1969 (N_1969,In_2091,In_804);
xor U1970 (N_1970,In_2200,In_763);
and U1971 (N_1971,In_570,In_2418);
and U1972 (N_1972,In_1710,In_1995);
nor U1973 (N_1973,In_916,In_781);
or U1974 (N_1974,In_95,In_1178);
nor U1975 (N_1975,In_1819,In_1753);
xor U1976 (N_1976,In_1891,In_1060);
xor U1977 (N_1977,In_1699,In_1212);
nor U1978 (N_1978,In_1497,In_2227);
or U1979 (N_1979,In_1945,In_1343);
nand U1980 (N_1980,In_466,In_2155);
nor U1981 (N_1981,In_2324,In_274);
nand U1982 (N_1982,In_136,In_1559);
nand U1983 (N_1983,In_1836,In_1588);
or U1984 (N_1984,In_2096,In_480);
xor U1985 (N_1985,In_1776,In_642);
and U1986 (N_1986,In_2330,In_869);
or U1987 (N_1987,In_1722,In_2195);
nand U1988 (N_1988,In_918,In_713);
nor U1989 (N_1989,In_2310,In_1159);
and U1990 (N_1990,In_1645,In_1182);
or U1991 (N_1991,In_880,In_1912);
xor U1992 (N_1992,In_1042,In_142);
and U1993 (N_1993,In_375,In_2277);
xor U1994 (N_1994,In_482,In_440);
and U1995 (N_1995,In_2041,In_1118);
or U1996 (N_1996,In_137,In_1552);
nor U1997 (N_1997,In_168,In_2472);
and U1998 (N_1998,In_587,In_1109);
nand U1999 (N_1999,In_45,In_881);
xnor U2000 (N_2000,In_169,In_987);
nor U2001 (N_2001,In_1271,In_1725);
xnor U2002 (N_2002,In_579,In_1778);
and U2003 (N_2003,In_515,In_1081);
nand U2004 (N_2004,In_854,In_397);
nor U2005 (N_2005,In_2463,In_2266);
xor U2006 (N_2006,In_529,In_2368);
or U2007 (N_2007,In_1819,In_2034);
nand U2008 (N_2008,In_1007,In_2269);
nor U2009 (N_2009,In_479,In_1646);
or U2010 (N_2010,In_701,In_1251);
nor U2011 (N_2011,In_632,In_445);
nand U2012 (N_2012,In_599,In_2473);
or U2013 (N_2013,In_1904,In_2229);
nand U2014 (N_2014,In_1493,In_2081);
nor U2015 (N_2015,In_11,In_1114);
xor U2016 (N_2016,In_383,In_2026);
nor U2017 (N_2017,In_2020,In_438);
and U2018 (N_2018,In_1998,In_2430);
nand U2019 (N_2019,In_568,In_2243);
nand U2020 (N_2020,In_2359,In_477);
nor U2021 (N_2021,In_1515,In_20);
nand U2022 (N_2022,In_410,In_489);
or U2023 (N_2023,In_1897,In_339);
nand U2024 (N_2024,In_469,In_1773);
xor U2025 (N_2025,In_160,In_2135);
or U2026 (N_2026,In_1805,In_2357);
xor U2027 (N_2027,In_1898,In_2311);
xnor U2028 (N_2028,In_828,In_2359);
nor U2029 (N_2029,In_620,In_2326);
or U2030 (N_2030,In_2196,In_490);
or U2031 (N_2031,In_1069,In_1357);
nand U2032 (N_2032,In_2114,In_2270);
nand U2033 (N_2033,In_16,In_1735);
nand U2034 (N_2034,In_2007,In_1091);
nor U2035 (N_2035,In_1268,In_503);
and U2036 (N_2036,In_198,In_2071);
nand U2037 (N_2037,In_1903,In_1361);
or U2038 (N_2038,In_798,In_2136);
xor U2039 (N_2039,In_1347,In_2162);
nand U2040 (N_2040,In_1697,In_1556);
or U2041 (N_2041,In_1462,In_898);
and U2042 (N_2042,In_389,In_2153);
nand U2043 (N_2043,In_1633,In_1389);
xor U2044 (N_2044,In_1827,In_2063);
xor U2045 (N_2045,In_2316,In_1982);
nand U2046 (N_2046,In_1291,In_1163);
and U2047 (N_2047,In_2272,In_1777);
xnor U2048 (N_2048,In_498,In_766);
or U2049 (N_2049,In_2248,In_2047);
xnor U2050 (N_2050,In_1095,In_1607);
and U2051 (N_2051,In_1129,In_2436);
nand U2052 (N_2052,In_1443,In_88);
xor U2053 (N_2053,In_985,In_1558);
xor U2054 (N_2054,In_2118,In_1636);
or U2055 (N_2055,In_1320,In_1068);
nand U2056 (N_2056,In_401,In_1753);
and U2057 (N_2057,In_1103,In_1809);
nand U2058 (N_2058,In_1396,In_1733);
nand U2059 (N_2059,In_677,In_1795);
and U2060 (N_2060,In_2365,In_1854);
xnor U2061 (N_2061,In_228,In_2470);
nand U2062 (N_2062,In_89,In_1976);
and U2063 (N_2063,In_1227,In_1721);
xor U2064 (N_2064,In_2392,In_298);
nand U2065 (N_2065,In_555,In_316);
or U2066 (N_2066,In_557,In_1563);
nor U2067 (N_2067,In_2057,In_1955);
xnor U2068 (N_2068,In_550,In_1581);
or U2069 (N_2069,In_1880,In_2494);
and U2070 (N_2070,In_1237,In_622);
and U2071 (N_2071,In_2223,In_1304);
and U2072 (N_2072,In_1492,In_650);
nand U2073 (N_2073,In_910,In_1318);
xnor U2074 (N_2074,In_1378,In_1369);
nand U2075 (N_2075,In_1682,In_31);
or U2076 (N_2076,In_541,In_1042);
or U2077 (N_2077,In_403,In_1151);
nand U2078 (N_2078,In_1844,In_1455);
and U2079 (N_2079,In_1983,In_269);
or U2080 (N_2080,In_587,In_1455);
and U2081 (N_2081,In_50,In_2032);
or U2082 (N_2082,In_1780,In_334);
or U2083 (N_2083,In_505,In_2481);
nand U2084 (N_2084,In_927,In_2208);
nor U2085 (N_2085,In_111,In_1980);
nor U2086 (N_2086,In_1203,In_60);
xor U2087 (N_2087,In_1004,In_1275);
or U2088 (N_2088,In_879,In_595);
xnor U2089 (N_2089,In_566,In_1475);
or U2090 (N_2090,In_1490,In_1164);
nand U2091 (N_2091,In_2165,In_776);
nor U2092 (N_2092,In_1058,In_146);
and U2093 (N_2093,In_990,In_82);
nand U2094 (N_2094,In_1221,In_2249);
nand U2095 (N_2095,In_672,In_1710);
nor U2096 (N_2096,In_1363,In_1478);
nor U2097 (N_2097,In_2366,In_614);
nor U2098 (N_2098,In_2326,In_1499);
xor U2099 (N_2099,In_628,In_2312);
or U2100 (N_2100,In_1549,In_1532);
xnor U2101 (N_2101,In_1228,In_511);
or U2102 (N_2102,In_2301,In_349);
nor U2103 (N_2103,In_72,In_227);
nand U2104 (N_2104,In_1124,In_855);
and U2105 (N_2105,In_1453,In_2433);
and U2106 (N_2106,In_1947,In_2234);
or U2107 (N_2107,In_709,In_456);
or U2108 (N_2108,In_87,In_1709);
nand U2109 (N_2109,In_2124,In_2173);
xnor U2110 (N_2110,In_2323,In_1744);
nand U2111 (N_2111,In_832,In_56);
or U2112 (N_2112,In_1274,In_1302);
nand U2113 (N_2113,In_2413,In_1230);
or U2114 (N_2114,In_269,In_579);
or U2115 (N_2115,In_1215,In_282);
nand U2116 (N_2116,In_2130,In_1500);
xnor U2117 (N_2117,In_244,In_1502);
nand U2118 (N_2118,In_755,In_137);
nand U2119 (N_2119,In_503,In_1357);
nand U2120 (N_2120,In_169,In_36);
or U2121 (N_2121,In_247,In_782);
and U2122 (N_2122,In_1188,In_1202);
or U2123 (N_2123,In_945,In_578);
or U2124 (N_2124,In_231,In_1607);
and U2125 (N_2125,In_2191,In_1135);
nor U2126 (N_2126,In_2012,In_395);
or U2127 (N_2127,In_65,In_2431);
and U2128 (N_2128,In_14,In_355);
nand U2129 (N_2129,In_1474,In_493);
xnor U2130 (N_2130,In_728,In_1928);
xnor U2131 (N_2131,In_2307,In_2280);
nand U2132 (N_2132,In_365,In_1986);
nor U2133 (N_2133,In_1047,In_666);
or U2134 (N_2134,In_973,In_53);
nor U2135 (N_2135,In_409,In_550);
xor U2136 (N_2136,In_1334,In_581);
nand U2137 (N_2137,In_1904,In_1102);
or U2138 (N_2138,In_1145,In_1703);
nand U2139 (N_2139,In_2134,In_1917);
nor U2140 (N_2140,In_1255,In_304);
and U2141 (N_2141,In_723,In_1570);
nor U2142 (N_2142,In_1067,In_1845);
or U2143 (N_2143,In_1806,In_165);
xnor U2144 (N_2144,In_549,In_470);
xor U2145 (N_2145,In_626,In_2415);
nand U2146 (N_2146,In_1234,In_22);
nor U2147 (N_2147,In_2268,In_1611);
nor U2148 (N_2148,In_1670,In_2233);
nor U2149 (N_2149,In_839,In_1469);
and U2150 (N_2150,In_891,In_2448);
and U2151 (N_2151,In_1765,In_2396);
xnor U2152 (N_2152,In_60,In_140);
nand U2153 (N_2153,In_2259,In_489);
nand U2154 (N_2154,In_1788,In_547);
xor U2155 (N_2155,In_1555,In_1270);
nor U2156 (N_2156,In_1897,In_428);
and U2157 (N_2157,In_1556,In_22);
nand U2158 (N_2158,In_843,In_414);
or U2159 (N_2159,In_1066,In_1981);
xor U2160 (N_2160,In_237,In_2045);
and U2161 (N_2161,In_1298,In_1368);
xor U2162 (N_2162,In_56,In_2230);
and U2163 (N_2163,In_2030,In_45);
or U2164 (N_2164,In_2048,In_329);
nor U2165 (N_2165,In_795,In_1678);
nor U2166 (N_2166,In_1449,In_1765);
nand U2167 (N_2167,In_1661,In_692);
nand U2168 (N_2168,In_1469,In_1394);
nand U2169 (N_2169,In_1872,In_1024);
nor U2170 (N_2170,In_554,In_732);
nor U2171 (N_2171,In_2380,In_645);
nand U2172 (N_2172,In_1363,In_1725);
and U2173 (N_2173,In_1429,In_1889);
xor U2174 (N_2174,In_1696,In_284);
or U2175 (N_2175,In_2395,In_2165);
or U2176 (N_2176,In_582,In_712);
nand U2177 (N_2177,In_271,In_2259);
and U2178 (N_2178,In_2347,In_423);
and U2179 (N_2179,In_1898,In_1096);
nor U2180 (N_2180,In_1553,In_883);
nor U2181 (N_2181,In_227,In_582);
nand U2182 (N_2182,In_26,In_207);
nand U2183 (N_2183,In_1511,In_1313);
nor U2184 (N_2184,In_1946,In_807);
nor U2185 (N_2185,In_2300,In_1606);
nor U2186 (N_2186,In_1433,In_1964);
or U2187 (N_2187,In_1566,In_335);
nor U2188 (N_2188,In_237,In_988);
nor U2189 (N_2189,In_1598,In_76);
or U2190 (N_2190,In_1425,In_1613);
nor U2191 (N_2191,In_1684,In_1327);
and U2192 (N_2192,In_1621,In_1245);
nor U2193 (N_2193,In_1884,In_1569);
and U2194 (N_2194,In_413,In_1809);
nor U2195 (N_2195,In_1333,In_2096);
and U2196 (N_2196,In_2134,In_1840);
nor U2197 (N_2197,In_1954,In_433);
nor U2198 (N_2198,In_1049,In_709);
nand U2199 (N_2199,In_1338,In_2001);
or U2200 (N_2200,In_181,In_914);
and U2201 (N_2201,In_1898,In_1070);
xnor U2202 (N_2202,In_1678,In_1033);
nand U2203 (N_2203,In_683,In_2436);
nor U2204 (N_2204,In_252,In_1820);
nand U2205 (N_2205,In_2216,In_1905);
or U2206 (N_2206,In_2154,In_1000);
and U2207 (N_2207,In_566,In_835);
or U2208 (N_2208,In_2177,In_2350);
nand U2209 (N_2209,In_972,In_2015);
nand U2210 (N_2210,In_1780,In_595);
and U2211 (N_2211,In_409,In_1729);
or U2212 (N_2212,In_278,In_1383);
nor U2213 (N_2213,In_2118,In_1225);
xor U2214 (N_2214,In_783,In_1465);
nor U2215 (N_2215,In_2238,In_1806);
xnor U2216 (N_2216,In_61,In_1143);
nand U2217 (N_2217,In_1608,In_2382);
or U2218 (N_2218,In_1344,In_2095);
nor U2219 (N_2219,In_979,In_984);
nor U2220 (N_2220,In_2222,In_1837);
xor U2221 (N_2221,In_1421,In_2052);
nand U2222 (N_2222,In_1005,In_1867);
nand U2223 (N_2223,In_1818,In_1579);
nand U2224 (N_2224,In_1689,In_2110);
nor U2225 (N_2225,In_2287,In_2200);
or U2226 (N_2226,In_993,In_1280);
or U2227 (N_2227,In_101,In_1045);
nor U2228 (N_2228,In_1337,In_2362);
nand U2229 (N_2229,In_1691,In_335);
or U2230 (N_2230,In_1583,In_2387);
and U2231 (N_2231,In_237,In_406);
xnor U2232 (N_2232,In_2265,In_49);
xor U2233 (N_2233,In_1141,In_1789);
or U2234 (N_2234,In_605,In_792);
and U2235 (N_2235,In_640,In_1680);
nand U2236 (N_2236,In_790,In_1129);
and U2237 (N_2237,In_2108,In_1796);
nand U2238 (N_2238,In_1162,In_2390);
and U2239 (N_2239,In_2338,In_4);
and U2240 (N_2240,In_68,In_1345);
nand U2241 (N_2241,In_155,In_558);
xor U2242 (N_2242,In_653,In_1047);
nor U2243 (N_2243,In_2417,In_729);
nor U2244 (N_2244,In_1385,In_72);
nor U2245 (N_2245,In_268,In_1436);
xnor U2246 (N_2246,In_239,In_1361);
nor U2247 (N_2247,In_876,In_1011);
nand U2248 (N_2248,In_2358,In_2450);
xnor U2249 (N_2249,In_1132,In_523);
or U2250 (N_2250,In_1246,In_664);
or U2251 (N_2251,In_157,In_1004);
or U2252 (N_2252,In_1815,In_2405);
or U2253 (N_2253,In_2275,In_1703);
and U2254 (N_2254,In_2139,In_1859);
nor U2255 (N_2255,In_65,In_1160);
or U2256 (N_2256,In_2291,In_1762);
nor U2257 (N_2257,In_2162,In_2292);
xnor U2258 (N_2258,In_1021,In_1288);
nor U2259 (N_2259,In_2198,In_1510);
xnor U2260 (N_2260,In_144,In_1294);
nand U2261 (N_2261,In_128,In_2435);
or U2262 (N_2262,In_1696,In_102);
xnor U2263 (N_2263,In_1431,In_1188);
and U2264 (N_2264,In_1100,In_1669);
and U2265 (N_2265,In_1256,In_247);
xnor U2266 (N_2266,In_1445,In_1799);
and U2267 (N_2267,In_1371,In_157);
or U2268 (N_2268,In_295,In_659);
nand U2269 (N_2269,In_1561,In_1275);
nor U2270 (N_2270,In_979,In_1881);
nor U2271 (N_2271,In_512,In_1193);
and U2272 (N_2272,In_314,In_1370);
nand U2273 (N_2273,In_1338,In_2303);
or U2274 (N_2274,In_1980,In_840);
or U2275 (N_2275,In_1801,In_2060);
and U2276 (N_2276,In_1475,In_76);
or U2277 (N_2277,In_2116,In_1602);
nand U2278 (N_2278,In_58,In_2427);
nand U2279 (N_2279,In_402,In_245);
xnor U2280 (N_2280,In_2399,In_493);
xnor U2281 (N_2281,In_187,In_2107);
nor U2282 (N_2282,In_198,In_1122);
or U2283 (N_2283,In_151,In_1568);
nand U2284 (N_2284,In_2224,In_51);
nand U2285 (N_2285,In_954,In_2432);
or U2286 (N_2286,In_227,In_1885);
nand U2287 (N_2287,In_387,In_212);
nor U2288 (N_2288,In_1836,In_1932);
and U2289 (N_2289,In_1510,In_1825);
or U2290 (N_2290,In_2481,In_2333);
and U2291 (N_2291,In_1865,In_1925);
nand U2292 (N_2292,In_2425,In_918);
and U2293 (N_2293,In_2163,In_1167);
nor U2294 (N_2294,In_1467,In_1104);
and U2295 (N_2295,In_2041,In_1396);
or U2296 (N_2296,In_833,In_1920);
nand U2297 (N_2297,In_2429,In_1596);
xor U2298 (N_2298,In_2438,In_913);
and U2299 (N_2299,In_1249,In_2069);
xor U2300 (N_2300,In_2098,In_473);
nand U2301 (N_2301,In_474,In_302);
and U2302 (N_2302,In_1956,In_2420);
nand U2303 (N_2303,In_2180,In_1303);
or U2304 (N_2304,In_1258,In_76);
nor U2305 (N_2305,In_1177,In_1803);
nand U2306 (N_2306,In_133,In_2397);
xor U2307 (N_2307,In_826,In_2053);
or U2308 (N_2308,In_884,In_25);
and U2309 (N_2309,In_2121,In_2013);
nor U2310 (N_2310,In_1199,In_303);
or U2311 (N_2311,In_2478,In_1791);
and U2312 (N_2312,In_405,In_2138);
nand U2313 (N_2313,In_958,In_1527);
xnor U2314 (N_2314,In_652,In_1896);
xnor U2315 (N_2315,In_1750,In_1051);
xnor U2316 (N_2316,In_150,In_906);
xnor U2317 (N_2317,In_2246,In_1229);
or U2318 (N_2318,In_876,In_1001);
nor U2319 (N_2319,In_1915,In_1580);
xor U2320 (N_2320,In_1184,In_2367);
or U2321 (N_2321,In_1217,In_2316);
xnor U2322 (N_2322,In_527,In_2032);
nor U2323 (N_2323,In_1590,In_166);
and U2324 (N_2324,In_994,In_921);
nor U2325 (N_2325,In_834,In_2395);
xor U2326 (N_2326,In_1642,In_568);
xor U2327 (N_2327,In_1221,In_2071);
nor U2328 (N_2328,In_1097,In_376);
nor U2329 (N_2329,In_2365,In_2375);
xor U2330 (N_2330,In_936,In_1478);
nand U2331 (N_2331,In_666,In_390);
and U2332 (N_2332,In_869,In_1461);
xor U2333 (N_2333,In_2443,In_1558);
and U2334 (N_2334,In_1062,In_142);
or U2335 (N_2335,In_1203,In_2071);
xnor U2336 (N_2336,In_1104,In_160);
nor U2337 (N_2337,In_2174,In_2052);
or U2338 (N_2338,In_1981,In_106);
xor U2339 (N_2339,In_205,In_1272);
and U2340 (N_2340,In_735,In_2454);
xor U2341 (N_2341,In_2090,In_392);
xnor U2342 (N_2342,In_40,In_1619);
or U2343 (N_2343,In_618,In_775);
and U2344 (N_2344,In_1118,In_60);
or U2345 (N_2345,In_1928,In_1153);
or U2346 (N_2346,In_2451,In_2383);
xor U2347 (N_2347,In_1196,In_893);
nor U2348 (N_2348,In_2180,In_411);
nand U2349 (N_2349,In_2346,In_1610);
or U2350 (N_2350,In_2008,In_982);
or U2351 (N_2351,In_1232,In_1162);
or U2352 (N_2352,In_1917,In_195);
xnor U2353 (N_2353,In_892,In_2358);
and U2354 (N_2354,In_803,In_775);
nand U2355 (N_2355,In_2223,In_2477);
and U2356 (N_2356,In_1795,In_358);
and U2357 (N_2357,In_780,In_1743);
and U2358 (N_2358,In_359,In_540);
or U2359 (N_2359,In_323,In_1484);
and U2360 (N_2360,In_1080,In_341);
nand U2361 (N_2361,In_683,In_1061);
nand U2362 (N_2362,In_1222,In_532);
xor U2363 (N_2363,In_2141,In_1093);
nand U2364 (N_2364,In_644,In_482);
nand U2365 (N_2365,In_1712,In_276);
nand U2366 (N_2366,In_1360,In_911);
nor U2367 (N_2367,In_891,In_1507);
nand U2368 (N_2368,In_1781,In_1864);
or U2369 (N_2369,In_2450,In_1282);
or U2370 (N_2370,In_387,In_2287);
nor U2371 (N_2371,In_1670,In_891);
or U2372 (N_2372,In_180,In_278);
and U2373 (N_2373,In_1947,In_909);
and U2374 (N_2374,In_886,In_2353);
nand U2375 (N_2375,In_716,In_129);
and U2376 (N_2376,In_2372,In_971);
xnor U2377 (N_2377,In_746,In_1204);
or U2378 (N_2378,In_2009,In_1674);
or U2379 (N_2379,In_779,In_101);
nor U2380 (N_2380,In_1902,In_245);
and U2381 (N_2381,In_1350,In_1108);
and U2382 (N_2382,In_2265,In_510);
nand U2383 (N_2383,In_2023,In_2094);
xnor U2384 (N_2384,In_2243,In_1048);
xnor U2385 (N_2385,In_1517,In_860);
nand U2386 (N_2386,In_1242,In_1267);
nor U2387 (N_2387,In_2464,In_1308);
nor U2388 (N_2388,In_719,In_563);
xnor U2389 (N_2389,In_712,In_588);
nor U2390 (N_2390,In_1883,In_997);
nor U2391 (N_2391,In_1526,In_212);
xnor U2392 (N_2392,In_286,In_2140);
and U2393 (N_2393,In_1037,In_1688);
and U2394 (N_2394,In_1216,In_1584);
nor U2395 (N_2395,In_1983,In_2320);
nand U2396 (N_2396,In_2288,In_690);
or U2397 (N_2397,In_1981,In_2341);
nor U2398 (N_2398,In_649,In_2270);
or U2399 (N_2399,In_115,In_986);
nand U2400 (N_2400,In_2308,In_1696);
or U2401 (N_2401,In_750,In_733);
and U2402 (N_2402,In_1265,In_1726);
xor U2403 (N_2403,In_1590,In_870);
nor U2404 (N_2404,In_2080,In_1592);
and U2405 (N_2405,In_1935,In_1823);
nor U2406 (N_2406,In_45,In_879);
nand U2407 (N_2407,In_537,In_224);
and U2408 (N_2408,In_326,In_2198);
nand U2409 (N_2409,In_1308,In_197);
nor U2410 (N_2410,In_1549,In_1529);
xnor U2411 (N_2411,In_1983,In_1389);
and U2412 (N_2412,In_1784,In_961);
nor U2413 (N_2413,In_1123,In_1283);
and U2414 (N_2414,In_1183,In_1352);
xor U2415 (N_2415,In_2226,In_1538);
and U2416 (N_2416,In_718,In_694);
nor U2417 (N_2417,In_2467,In_2442);
and U2418 (N_2418,In_1503,In_733);
xnor U2419 (N_2419,In_1818,In_1088);
nand U2420 (N_2420,In_185,In_827);
and U2421 (N_2421,In_1324,In_1759);
and U2422 (N_2422,In_1350,In_241);
nor U2423 (N_2423,In_1086,In_2268);
nor U2424 (N_2424,In_45,In_616);
or U2425 (N_2425,In_477,In_1902);
and U2426 (N_2426,In_1982,In_1931);
and U2427 (N_2427,In_2163,In_876);
and U2428 (N_2428,In_1384,In_361);
xor U2429 (N_2429,In_2458,In_555);
xnor U2430 (N_2430,In_2192,In_2191);
nor U2431 (N_2431,In_1423,In_1769);
and U2432 (N_2432,In_2451,In_2419);
nor U2433 (N_2433,In_1657,In_920);
or U2434 (N_2434,In_2178,In_2464);
nand U2435 (N_2435,In_1831,In_1909);
and U2436 (N_2436,In_1923,In_79);
nand U2437 (N_2437,In_1591,In_1276);
xor U2438 (N_2438,In_805,In_1500);
and U2439 (N_2439,In_302,In_1537);
xor U2440 (N_2440,In_1958,In_758);
or U2441 (N_2441,In_177,In_953);
and U2442 (N_2442,In_335,In_1764);
nand U2443 (N_2443,In_2480,In_557);
nand U2444 (N_2444,In_1901,In_1214);
and U2445 (N_2445,In_2426,In_881);
nor U2446 (N_2446,In_976,In_2213);
and U2447 (N_2447,In_1007,In_938);
or U2448 (N_2448,In_311,In_1277);
and U2449 (N_2449,In_938,In_727);
or U2450 (N_2450,In_1510,In_1800);
or U2451 (N_2451,In_214,In_1109);
nor U2452 (N_2452,In_1657,In_190);
xnor U2453 (N_2453,In_1650,In_2247);
or U2454 (N_2454,In_1319,In_1218);
and U2455 (N_2455,In_1435,In_285);
nor U2456 (N_2456,In_534,In_1893);
nand U2457 (N_2457,In_2396,In_1045);
nor U2458 (N_2458,In_1472,In_735);
and U2459 (N_2459,In_965,In_2183);
xnor U2460 (N_2460,In_1117,In_2277);
nor U2461 (N_2461,In_2133,In_2222);
or U2462 (N_2462,In_1263,In_1225);
nand U2463 (N_2463,In_2341,In_1898);
and U2464 (N_2464,In_2357,In_1622);
and U2465 (N_2465,In_1170,In_1408);
and U2466 (N_2466,In_300,In_1664);
and U2467 (N_2467,In_778,In_359);
xor U2468 (N_2468,In_1233,In_304);
and U2469 (N_2469,In_2135,In_2078);
nand U2470 (N_2470,In_1423,In_899);
xor U2471 (N_2471,In_1132,In_2089);
or U2472 (N_2472,In_135,In_332);
nand U2473 (N_2473,In_48,In_1738);
xor U2474 (N_2474,In_1017,In_380);
nand U2475 (N_2475,In_1211,In_1310);
or U2476 (N_2476,In_1613,In_1683);
nor U2477 (N_2477,In_1774,In_1063);
or U2478 (N_2478,In_2043,In_2142);
xor U2479 (N_2479,In_1520,In_1103);
nor U2480 (N_2480,In_758,In_2456);
or U2481 (N_2481,In_633,In_38);
or U2482 (N_2482,In_802,In_590);
or U2483 (N_2483,In_1692,In_1993);
nand U2484 (N_2484,In_1998,In_347);
nand U2485 (N_2485,In_79,In_1030);
nand U2486 (N_2486,In_2249,In_1232);
and U2487 (N_2487,In_1792,In_1497);
nor U2488 (N_2488,In_2093,In_2198);
nor U2489 (N_2489,In_1489,In_1445);
or U2490 (N_2490,In_459,In_1120);
nand U2491 (N_2491,In_2091,In_1100);
xnor U2492 (N_2492,In_1653,In_1989);
nor U2493 (N_2493,In_418,In_98);
or U2494 (N_2494,In_1647,In_1437);
or U2495 (N_2495,In_943,In_1014);
and U2496 (N_2496,In_1161,In_1446);
or U2497 (N_2497,In_11,In_1259);
and U2498 (N_2498,In_838,In_1590);
xnor U2499 (N_2499,In_1420,In_1873);
nor U2500 (N_2500,In_356,In_1134);
nor U2501 (N_2501,In_1058,In_1322);
or U2502 (N_2502,In_1148,In_1225);
nor U2503 (N_2503,In_2066,In_1425);
or U2504 (N_2504,In_1666,In_2496);
nand U2505 (N_2505,In_1207,In_45);
nand U2506 (N_2506,In_2197,In_216);
nand U2507 (N_2507,In_1014,In_623);
and U2508 (N_2508,In_2465,In_1036);
or U2509 (N_2509,In_533,In_174);
or U2510 (N_2510,In_2242,In_1832);
or U2511 (N_2511,In_1378,In_1049);
xnor U2512 (N_2512,In_718,In_1509);
or U2513 (N_2513,In_1811,In_1271);
and U2514 (N_2514,In_677,In_1988);
nor U2515 (N_2515,In_632,In_1871);
xnor U2516 (N_2516,In_348,In_463);
and U2517 (N_2517,In_1766,In_1223);
xor U2518 (N_2518,In_1913,In_2310);
nand U2519 (N_2519,In_825,In_397);
nand U2520 (N_2520,In_641,In_1337);
xnor U2521 (N_2521,In_1758,In_948);
xnor U2522 (N_2522,In_15,In_392);
xor U2523 (N_2523,In_1266,In_616);
or U2524 (N_2524,In_2173,In_12);
xnor U2525 (N_2525,In_2406,In_1571);
and U2526 (N_2526,In_2016,In_2453);
nor U2527 (N_2527,In_847,In_129);
or U2528 (N_2528,In_1644,In_1680);
nor U2529 (N_2529,In_1047,In_1264);
nor U2530 (N_2530,In_601,In_532);
or U2531 (N_2531,In_1672,In_1476);
or U2532 (N_2532,In_1091,In_1674);
or U2533 (N_2533,In_1281,In_2322);
nor U2534 (N_2534,In_555,In_2147);
or U2535 (N_2535,In_743,In_1197);
nand U2536 (N_2536,In_491,In_877);
xnor U2537 (N_2537,In_1700,In_2226);
nand U2538 (N_2538,In_40,In_1298);
xor U2539 (N_2539,In_2433,In_1943);
xnor U2540 (N_2540,In_1037,In_1392);
and U2541 (N_2541,In_607,In_2211);
xnor U2542 (N_2542,In_564,In_1322);
or U2543 (N_2543,In_752,In_735);
nor U2544 (N_2544,In_1627,In_231);
or U2545 (N_2545,In_2053,In_1013);
and U2546 (N_2546,In_641,In_2474);
or U2547 (N_2547,In_1899,In_1664);
and U2548 (N_2548,In_1177,In_1978);
xor U2549 (N_2549,In_1895,In_2070);
nor U2550 (N_2550,In_2114,In_822);
or U2551 (N_2551,In_1840,In_427);
nor U2552 (N_2552,In_1263,In_1451);
and U2553 (N_2553,In_1129,In_276);
nand U2554 (N_2554,In_1734,In_1793);
nor U2555 (N_2555,In_2236,In_1694);
and U2556 (N_2556,In_2232,In_1974);
or U2557 (N_2557,In_340,In_1352);
or U2558 (N_2558,In_1170,In_1192);
nor U2559 (N_2559,In_1432,In_298);
and U2560 (N_2560,In_1830,In_526);
nand U2561 (N_2561,In_1225,In_405);
and U2562 (N_2562,In_1509,In_2346);
xor U2563 (N_2563,In_959,In_883);
or U2564 (N_2564,In_1985,In_85);
nor U2565 (N_2565,In_2309,In_1170);
nand U2566 (N_2566,In_352,In_1065);
or U2567 (N_2567,In_2489,In_84);
nor U2568 (N_2568,In_1934,In_756);
xnor U2569 (N_2569,In_310,In_137);
and U2570 (N_2570,In_210,In_2145);
nand U2571 (N_2571,In_1429,In_1066);
nor U2572 (N_2572,In_674,In_1471);
or U2573 (N_2573,In_1303,In_1851);
nand U2574 (N_2574,In_806,In_1621);
nand U2575 (N_2575,In_756,In_625);
or U2576 (N_2576,In_668,In_864);
nor U2577 (N_2577,In_435,In_2343);
nand U2578 (N_2578,In_2454,In_1622);
or U2579 (N_2579,In_377,In_1664);
xor U2580 (N_2580,In_380,In_113);
nand U2581 (N_2581,In_1708,In_1019);
xnor U2582 (N_2582,In_1603,In_1682);
xor U2583 (N_2583,In_1432,In_617);
nor U2584 (N_2584,In_2330,In_1039);
and U2585 (N_2585,In_1507,In_2308);
nor U2586 (N_2586,In_1957,In_401);
xor U2587 (N_2587,In_871,In_514);
nand U2588 (N_2588,In_256,In_967);
xnor U2589 (N_2589,In_1951,In_1708);
nor U2590 (N_2590,In_1258,In_2374);
or U2591 (N_2591,In_836,In_203);
xnor U2592 (N_2592,In_1383,In_1189);
and U2593 (N_2593,In_233,In_2449);
nand U2594 (N_2594,In_1346,In_321);
or U2595 (N_2595,In_1330,In_1325);
nor U2596 (N_2596,In_1311,In_570);
and U2597 (N_2597,In_1680,In_1119);
xnor U2598 (N_2598,In_1814,In_1924);
and U2599 (N_2599,In_2066,In_888);
nand U2600 (N_2600,In_1828,In_1935);
and U2601 (N_2601,In_2180,In_489);
xnor U2602 (N_2602,In_718,In_1455);
or U2603 (N_2603,In_25,In_441);
nor U2604 (N_2604,In_875,In_406);
nand U2605 (N_2605,In_1913,In_345);
xnor U2606 (N_2606,In_406,In_355);
xor U2607 (N_2607,In_2431,In_307);
nand U2608 (N_2608,In_1923,In_34);
xnor U2609 (N_2609,In_1732,In_253);
or U2610 (N_2610,In_1409,In_800);
or U2611 (N_2611,In_2199,In_427);
nand U2612 (N_2612,In_640,In_2052);
nand U2613 (N_2613,In_2220,In_2006);
xor U2614 (N_2614,In_575,In_2133);
or U2615 (N_2615,In_1544,In_1627);
and U2616 (N_2616,In_2484,In_153);
nor U2617 (N_2617,In_2091,In_2092);
and U2618 (N_2618,In_239,In_824);
xnor U2619 (N_2619,In_1799,In_259);
nor U2620 (N_2620,In_1875,In_391);
and U2621 (N_2621,In_852,In_1189);
nor U2622 (N_2622,In_1398,In_1731);
xor U2623 (N_2623,In_2210,In_1227);
or U2624 (N_2624,In_2085,In_1341);
nor U2625 (N_2625,In_215,In_2089);
xnor U2626 (N_2626,In_2420,In_218);
or U2627 (N_2627,In_1270,In_2354);
nor U2628 (N_2628,In_189,In_1861);
or U2629 (N_2629,In_1803,In_2141);
nor U2630 (N_2630,In_1758,In_2177);
xor U2631 (N_2631,In_1212,In_1386);
and U2632 (N_2632,In_840,In_1875);
or U2633 (N_2633,In_55,In_1791);
xor U2634 (N_2634,In_2114,In_902);
or U2635 (N_2635,In_2163,In_1166);
xnor U2636 (N_2636,In_1883,In_1761);
and U2637 (N_2637,In_1472,In_2156);
xnor U2638 (N_2638,In_2246,In_673);
or U2639 (N_2639,In_2105,In_1457);
nor U2640 (N_2640,In_47,In_15);
nand U2641 (N_2641,In_53,In_1860);
xor U2642 (N_2642,In_2095,In_788);
nor U2643 (N_2643,In_137,In_1443);
nand U2644 (N_2644,In_1589,In_2462);
nand U2645 (N_2645,In_1731,In_2197);
or U2646 (N_2646,In_1012,In_1306);
or U2647 (N_2647,In_966,In_1745);
nor U2648 (N_2648,In_2298,In_95);
nor U2649 (N_2649,In_2048,In_880);
xor U2650 (N_2650,In_1651,In_526);
nor U2651 (N_2651,In_1942,In_1625);
or U2652 (N_2652,In_2182,In_1721);
and U2653 (N_2653,In_945,In_1700);
nor U2654 (N_2654,In_1888,In_1486);
nor U2655 (N_2655,In_106,In_2091);
or U2656 (N_2656,In_2153,In_2326);
xnor U2657 (N_2657,In_288,In_847);
nand U2658 (N_2658,In_2405,In_2002);
nand U2659 (N_2659,In_658,In_2396);
nor U2660 (N_2660,In_654,In_100);
or U2661 (N_2661,In_1487,In_738);
or U2662 (N_2662,In_2272,In_1981);
nor U2663 (N_2663,In_984,In_2145);
or U2664 (N_2664,In_766,In_1132);
nor U2665 (N_2665,In_223,In_2394);
xnor U2666 (N_2666,In_1354,In_1920);
nand U2667 (N_2667,In_2153,In_1182);
or U2668 (N_2668,In_571,In_1288);
nor U2669 (N_2669,In_894,In_642);
nand U2670 (N_2670,In_2271,In_2243);
and U2671 (N_2671,In_1232,In_23);
nand U2672 (N_2672,In_2176,In_1093);
and U2673 (N_2673,In_1721,In_2141);
nand U2674 (N_2674,In_2233,In_2020);
and U2675 (N_2675,In_1343,In_1126);
xor U2676 (N_2676,In_1032,In_1232);
nor U2677 (N_2677,In_11,In_2011);
nand U2678 (N_2678,In_541,In_932);
xor U2679 (N_2679,In_1301,In_1692);
and U2680 (N_2680,In_2166,In_836);
and U2681 (N_2681,In_675,In_1946);
xor U2682 (N_2682,In_2281,In_1352);
or U2683 (N_2683,In_1392,In_553);
xor U2684 (N_2684,In_1502,In_1256);
nor U2685 (N_2685,In_1239,In_1109);
xor U2686 (N_2686,In_887,In_2166);
or U2687 (N_2687,In_992,In_2320);
nand U2688 (N_2688,In_2178,In_1706);
xnor U2689 (N_2689,In_561,In_204);
or U2690 (N_2690,In_2011,In_24);
xnor U2691 (N_2691,In_581,In_1979);
nand U2692 (N_2692,In_73,In_2119);
or U2693 (N_2693,In_1603,In_351);
nand U2694 (N_2694,In_1787,In_1258);
xor U2695 (N_2695,In_453,In_1127);
nand U2696 (N_2696,In_2127,In_160);
or U2697 (N_2697,In_502,In_908);
or U2698 (N_2698,In_591,In_2109);
or U2699 (N_2699,In_1511,In_1260);
or U2700 (N_2700,In_711,In_225);
and U2701 (N_2701,In_2356,In_1291);
or U2702 (N_2702,In_2262,In_1974);
nor U2703 (N_2703,In_263,In_2001);
and U2704 (N_2704,In_1110,In_2063);
nand U2705 (N_2705,In_1,In_2052);
nand U2706 (N_2706,In_1664,In_2489);
nand U2707 (N_2707,In_732,In_1831);
xnor U2708 (N_2708,In_692,In_1366);
nand U2709 (N_2709,In_1916,In_2226);
xnor U2710 (N_2710,In_1246,In_804);
nor U2711 (N_2711,In_726,In_326);
or U2712 (N_2712,In_1014,In_2038);
or U2713 (N_2713,In_1927,In_1762);
xor U2714 (N_2714,In_1584,In_796);
and U2715 (N_2715,In_1690,In_1457);
nor U2716 (N_2716,In_2438,In_1842);
and U2717 (N_2717,In_1747,In_1416);
or U2718 (N_2718,In_2199,In_2020);
nor U2719 (N_2719,In_2212,In_1946);
and U2720 (N_2720,In_2499,In_1811);
nand U2721 (N_2721,In_51,In_417);
xnor U2722 (N_2722,In_575,In_18);
or U2723 (N_2723,In_2262,In_733);
and U2724 (N_2724,In_617,In_890);
nand U2725 (N_2725,In_2091,In_1729);
and U2726 (N_2726,In_1381,In_2340);
or U2727 (N_2727,In_1891,In_618);
nor U2728 (N_2728,In_1744,In_2384);
xnor U2729 (N_2729,In_738,In_839);
nand U2730 (N_2730,In_104,In_1693);
nor U2731 (N_2731,In_1594,In_2471);
or U2732 (N_2732,In_2083,In_936);
nand U2733 (N_2733,In_1473,In_697);
or U2734 (N_2734,In_892,In_1447);
nor U2735 (N_2735,In_1599,In_1687);
xnor U2736 (N_2736,In_1643,In_606);
nand U2737 (N_2737,In_1060,In_937);
xor U2738 (N_2738,In_1905,In_862);
nand U2739 (N_2739,In_1424,In_125);
nor U2740 (N_2740,In_1073,In_1652);
and U2741 (N_2741,In_1191,In_1328);
nand U2742 (N_2742,In_294,In_169);
xor U2743 (N_2743,In_17,In_2068);
or U2744 (N_2744,In_1203,In_610);
or U2745 (N_2745,In_546,In_1455);
xnor U2746 (N_2746,In_1320,In_1174);
xnor U2747 (N_2747,In_834,In_1084);
nor U2748 (N_2748,In_403,In_1841);
xor U2749 (N_2749,In_162,In_751);
nand U2750 (N_2750,In_1081,In_1135);
xor U2751 (N_2751,In_1554,In_1685);
or U2752 (N_2752,In_144,In_1935);
nand U2753 (N_2753,In_696,In_489);
and U2754 (N_2754,In_1316,In_21);
or U2755 (N_2755,In_725,In_1368);
nor U2756 (N_2756,In_1522,In_1744);
xor U2757 (N_2757,In_394,In_1305);
nand U2758 (N_2758,In_1519,In_896);
nor U2759 (N_2759,In_2226,In_272);
nor U2760 (N_2760,In_247,In_558);
xnor U2761 (N_2761,In_1357,In_2196);
xor U2762 (N_2762,In_717,In_5);
nand U2763 (N_2763,In_206,In_1209);
and U2764 (N_2764,In_2077,In_1721);
nor U2765 (N_2765,In_472,In_1216);
and U2766 (N_2766,In_305,In_1136);
xor U2767 (N_2767,In_687,In_131);
nand U2768 (N_2768,In_947,In_1446);
nand U2769 (N_2769,In_153,In_1445);
nand U2770 (N_2770,In_2377,In_1986);
and U2771 (N_2771,In_2416,In_851);
or U2772 (N_2772,In_653,In_1081);
xor U2773 (N_2773,In_2356,In_801);
nand U2774 (N_2774,In_2143,In_2345);
nor U2775 (N_2775,In_1083,In_1206);
nor U2776 (N_2776,In_1712,In_342);
nor U2777 (N_2777,In_2080,In_1054);
xnor U2778 (N_2778,In_23,In_1052);
xnor U2779 (N_2779,In_933,In_1367);
nor U2780 (N_2780,In_628,In_618);
and U2781 (N_2781,In_830,In_1049);
nor U2782 (N_2782,In_1489,In_1343);
or U2783 (N_2783,In_1528,In_1824);
nand U2784 (N_2784,In_1193,In_867);
nand U2785 (N_2785,In_2312,In_205);
nand U2786 (N_2786,In_1837,In_1665);
and U2787 (N_2787,In_1208,In_2244);
or U2788 (N_2788,In_124,In_190);
and U2789 (N_2789,In_1929,In_178);
xor U2790 (N_2790,In_551,In_1341);
and U2791 (N_2791,In_2110,In_1917);
and U2792 (N_2792,In_883,In_430);
nor U2793 (N_2793,In_1768,In_2249);
and U2794 (N_2794,In_1256,In_503);
nand U2795 (N_2795,In_2190,In_1617);
nor U2796 (N_2796,In_1851,In_1809);
and U2797 (N_2797,In_1832,In_2180);
nor U2798 (N_2798,In_369,In_2155);
xor U2799 (N_2799,In_308,In_2112);
xor U2800 (N_2800,In_385,In_1128);
nand U2801 (N_2801,In_307,In_1862);
nor U2802 (N_2802,In_971,In_830);
and U2803 (N_2803,In_1282,In_56);
nand U2804 (N_2804,In_83,In_465);
xnor U2805 (N_2805,In_1331,In_3);
and U2806 (N_2806,In_1240,In_527);
xor U2807 (N_2807,In_2374,In_322);
nor U2808 (N_2808,In_202,In_63);
or U2809 (N_2809,In_722,In_1555);
nor U2810 (N_2810,In_430,In_2461);
nand U2811 (N_2811,In_485,In_768);
xor U2812 (N_2812,In_2111,In_1091);
and U2813 (N_2813,In_509,In_1582);
nand U2814 (N_2814,In_522,In_2036);
xor U2815 (N_2815,In_605,In_133);
xor U2816 (N_2816,In_667,In_927);
or U2817 (N_2817,In_1637,In_2398);
or U2818 (N_2818,In_1910,In_1265);
xnor U2819 (N_2819,In_720,In_2461);
xor U2820 (N_2820,In_1112,In_1670);
and U2821 (N_2821,In_1278,In_678);
nand U2822 (N_2822,In_1428,In_2051);
nor U2823 (N_2823,In_89,In_2373);
or U2824 (N_2824,In_532,In_2497);
nand U2825 (N_2825,In_102,In_484);
and U2826 (N_2826,In_1439,In_96);
nand U2827 (N_2827,In_1127,In_543);
nor U2828 (N_2828,In_1435,In_1978);
nor U2829 (N_2829,In_811,In_35);
nand U2830 (N_2830,In_549,In_524);
xnor U2831 (N_2831,In_2106,In_905);
and U2832 (N_2832,In_79,In_483);
or U2833 (N_2833,In_676,In_1643);
and U2834 (N_2834,In_2226,In_2015);
and U2835 (N_2835,In_678,In_2176);
xor U2836 (N_2836,In_728,In_800);
or U2837 (N_2837,In_1922,In_1346);
nand U2838 (N_2838,In_1995,In_1182);
nor U2839 (N_2839,In_1403,In_71);
and U2840 (N_2840,In_68,In_2300);
or U2841 (N_2841,In_1546,In_1188);
xnor U2842 (N_2842,In_2277,In_530);
or U2843 (N_2843,In_2286,In_2481);
nor U2844 (N_2844,In_2000,In_2034);
or U2845 (N_2845,In_1629,In_1776);
nor U2846 (N_2846,In_1836,In_1945);
or U2847 (N_2847,In_298,In_481);
or U2848 (N_2848,In_490,In_2421);
or U2849 (N_2849,In_2417,In_2380);
xnor U2850 (N_2850,In_1708,In_1536);
and U2851 (N_2851,In_1089,In_491);
xor U2852 (N_2852,In_615,In_2090);
or U2853 (N_2853,In_1155,In_2280);
and U2854 (N_2854,In_858,In_500);
nor U2855 (N_2855,In_607,In_370);
nand U2856 (N_2856,In_1934,In_802);
xor U2857 (N_2857,In_1329,In_846);
nor U2858 (N_2858,In_108,In_775);
and U2859 (N_2859,In_2037,In_447);
xnor U2860 (N_2860,In_412,In_1646);
nand U2861 (N_2861,In_1401,In_1340);
or U2862 (N_2862,In_1318,In_681);
and U2863 (N_2863,In_1054,In_1928);
or U2864 (N_2864,In_1482,In_1751);
or U2865 (N_2865,In_1805,In_880);
xnor U2866 (N_2866,In_963,In_2112);
or U2867 (N_2867,In_2211,In_319);
and U2868 (N_2868,In_2303,In_1385);
nor U2869 (N_2869,In_179,In_2152);
xor U2870 (N_2870,In_1205,In_1991);
nand U2871 (N_2871,In_1172,In_3);
nand U2872 (N_2872,In_336,In_548);
xor U2873 (N_2873,In_2203,In_322);
xor U2874 (N_2874,In_792,In_1042);
nand U2875 (N_2875,In_1391,In_901);
xnor U2876 (N_2876,In_1951,In_58);
or U2877 (N_2877,In_530,In_2157);
and U2878 (N_2878,In_607,In_1535);
nor U2879 (N_2879,In_5,In_1041);
or U2880 (N_2880,In_571,In_910);
and U2881 (N_2881,In_1820,In_808);
xnor U2882 (N_2882,In_1012,In_1137);
xnor U2883 (N_2883,In_83,In_377);
or U2884 (N_2884,In_434,In_1574);
nand U2885 (N_2885,In_238,In_1829);
and U2886 (N_2886,In_189,In_2062);
xnor U2887 (N_2887,In_1685,In_1838);
nor U2888 (N_2888,In_1803,In_1063);
nand U2889 (N_2889,In_503,In_1651);
and U2890 (N_2890,In_2430,In_2429);
and U2891 (N_2891,In_359,In_2413);
nand U2892 (N_2892,In_835,In_1313);
nand U2893 (N_2893,In_656,In_179);
or U2894 (N_2894,In_2326,In_1274);
nand U2895 (N_2895,In_1892,In_240);
xor U2896 (N_2896,In_1788,In_388);
and U2897 (N_2897,In_1645,In_435);
nor U2898 (N_2898,In_551,In_558);
xnor U2899 (N_2899,In_1748,In_1371);
and U2900 (N_2900,In_1385,In_1794);
or U2901 (N_2901,In_1702,In_2146);
xor U2902 (N_2902,In_607,In_2047);
and U2903 (N_2903,In_642,In_1718);
nand U2904 (N_2904,In_437,In_2148);
and U2905 (N_2905,In_2221,In_1067);
and U2906 (N_2906,In_1292,In_523);
or U2907 (N_2907,In_86,In_1622);
nor U2908 (N_2908,In_433,In_2404);
nor U2909 (N_2909,In_1787,In_867);
and U2910 (N_2910,In_1979,In_957);
nor U2911 (N_2911,In_1203,In_362);
xnor U2912 (N_2912,In_867,In_668);
xnor U2913 (N_2913,In_1698,In_1627);
nand U2914 (N_2914,In_2364,In_563);
nor U2915 (N_2915,In_2172,In_520);
xor U2916 (N_2916,In_1372,In_363);
or U2917 (N_2917,In_2330,In_164);
and U2918 (N_2918,In_1306,In_382);
nor U2919 (N_2919,In_2075,In_912);
and U2920 (N_2920,In_2003,In_1386);
and U2921 (N_2921,In_916,In_1188);
nor U2922 (N_2922,In_2386,In_22);
nor U2923 (N_2923,In_34,In_563);
xnor U2924 (N_2924,In_1549,In_1399);
nor U2925 (N_2925,In_1562,In_844);
and U2926 (N_2926,In_1214,In_301);
and U2927 (N_2927,In_1050,In_1376);
nor U2928 (N_2928,In_682,In_1335);
and U2929 (N_2929,In_170,In_1288);
nor U2930 (N_2930,In_56,In_264);
nand U2931 (N_2931,In_689,In_1587);
xnor U2932 (N_2932,In_258,In_871);
nor U2933 (N_2933,In_2117,In_1999);
or U2934 (N_2934,In_530,In_2132);
or U2935 (N_2935,In_257,In_2459);
nor U2936 (N_2936,In_1999,In_50);
or U2937 (N_2937,In_2150,In_839);
or U2938 (N_2938,In_2083,In_42);
and U2939 (N_2939,In_765,In_1155);
nor U2940 (N_2940,In_999,In_2323);
xor U2941 (N_2941,In_1028,In_152);
nor U2942 (N_2942,In_2251,In_2317);
or U2943 (N_2943,In_1540,In_889);
or U2944 (N_2944,In_1984,In_1588);
or U2945 (N_2945,In_2077,In_2222);
nand U2946 (N_2946,In_1575,In_460);
xnor U2947 (N_2947,In_25,In_848);
nor U2948 (N_2948,In_1543,In_68);
nand U2949 (N_2949,In_2119,In_373);
or U2950 (N_2950,In_190,In_2180);
nor U2951 (N_2951,In_2428,In_2063);
nor U2952 (N_2952,In_1838,In_898);
xnor U2953 (N_2953,In_829,In_1449);
nor U2954 (N_2954,In_1763,In_1753);
or U2955 (N_2955,In_1738,In_2066);
xor U2956 (N_2956,In_650,In_1010);
nor U2957 (N_2957,In_1086,In_668);
xnor U2958 (N_2958,In_1430,In_2122);
nand U2959 (N_2959,In_2453,In_445);
or U2960 (N_2960,In_1290,In_1635);
nand U2961 (N_2961,In_2025,In_661);
nand U2962 (N_2962,In_1374,In_2321);
and U2963 (N_2963,In_1450,In_1192);
nor U2964 (N_2964,In_2052,In_2487);
nand U2965 (N_2965,In_390,In_640);
xor U2966 (N_2966,In_278,In_1960);
nand U2967 (N_2967,In_902,In_1240);
or U2968 (N_2968,In_2131,In_485);
nor U2969 (N_2969,In_952,In_1728);
nand U2970 (N_2970,In_2424,In_969);
nor U2971 (N_2971,In_1898,In_501);
or U2972 (N_2972,In_1166,In_553);
nor U2973 (N_2973,In_219,In_280);
and U2974 (N_2974,In_1476,In_1609);
nor U2975 (N_2975,In_667,In_788);
nor U2976 (N_2976,In_75,In_170);
nor U2977 (N_2977,In_704,In_965);
nor U2978 (N_2978,In_1185,In_1651);
and U2979 (N_2979,In_453,In_2286);
and U2980 (N_2980,In_135,In_1307);
xor U2981 (N_2981,In_1432,In_2023);
nor U2982 (N_2982,In_1823,In_52);
nand U2983 (N_2983,In_2103,In_793);
nor U2984 (N_2984,In_1909,In_437);
xnor U2985 (N_2985,In_2303,In_1251);
nand U2986 (N_2986,In_382,In_1912);
and U2987 (N_2987,In_1076,In_1226);
nor U2988 (N_2988,In_291,In_1361);
nand U2989 (N_2989,In_2084,In_1123);
and U2990 (N_2990,In_782,In_88);
xnor U2991 (N_2991,In_127,In_2378);
or U2992 (N_2992,In_168,In_1857);
nand U2993 (N_2993,In_1224,In_2083);
nor U2994 (N_2994,In_825,In_1241);
nor U2995 (N_2995,In_2338,In_2084);
xnor U2996 (N_2996,In_265,In_213);
and U2997 (N_2997,In_118,In_2153);
xnor U2998 (N_2998,In_1825,In_2197);
and U2999 (N_2999,In_1331,In_2472);
and U3000 (N_3000,In_1975,In_2008);
and U3001 (N_3001,In_2307,In_367);
nand U3002 (N_3002,In_396,In_1699);
and U3003 (N_3003,In_1858,In_261);
xnor U3004 (N_3004,In_459,In_2025);
nor U3005 (N_3005,In_1776,In_2359);
nand U3006 (N_3006,In_1890,In_767);
or U3007 (N_3007,In_348,In_361);
or U3008 (N_3008,In_1825,In_2430);
nand U3009 (N_3009,In_1210,In_2425);
nor U3010 (N_3010,In_1744,In_581);
or U3011 (N_3011,In_613,In_1580);
and U3012 (N_3012,In_157,In_673);
xnor U3013 (N_3013,In_2054,In_48);
or U3014 (N_3014,In_2021,In_1038);
nor U3015 (N_3015,In_189,In_1091);
or U3016 (N_3016,In_2224,In_391);
and U3017 (N_3017,In_1954,In_25);
nand U3018 (N_3018,In_1769,In_613);
nor U3019 (N_3019,In_525,In_169);
nor U3020 (N_3020,In_2192,In_1129);
nor U3021 (N_3021,In_1649,In_1021);
and U3022 (N_3022,In_1006,In_1372);
xnor U3023 (N_3023,In_2373,In_1298);
or U3024 (N_3024,In_1398,In_1059);
nor U3025 (N_3025,In_331,In_2393);
nor U3026 (N_3026,In_1136,In_1101);
nand U3027 (N_3027,In_520,In_1553);
nor U3028 (N_3028,In_2499,In_4);
nand U3029 (N_3029,In_1224,In_2436);
nand U3030 (N_3030,In_1304,In_2472);
nand U3031 (N_3031,In_1578,In_2093);
xnor U3032 (N_3032,In_2018,In_347);
and U3033 (N_3033,In_2450,In_748);
xnor U3034 (N_3034,In_9,In_887);
or U3035 (N_3035,In_1702,In_1307);
nor U3036 (N_3036,In_1310,In_1686);
and U3037 (N_3037,In_577,In_2174);
nor U3038 (N_3038,In_270,In_2410);
and U3039 (N_3039,In_61,In_490);
and U3040 (N_3040,In_129,In_1289);
xor U3041 (N_3041,In_415,In_704);
nand U3042 (N_3042,In_1654,In_2294);
or U3043 (N_3043,In_150,In_1955);
nand U3044 (N_3044,In_1883,In_856);
nand U3045 (N_3045,In_502,In_1493);
xnor U3046 (N_3046,In_794,In_1545);
xor U3047 (N_3047,In_239,In_1301);
nor U3048 (N_3048,In_2390,In_357);
or U3049 (N_3049,In_269,In_1768);
xnor U3050 (N_3050,In_1543,In_1297);
nand U3051 (N_3051,In_1795,In_1380);
and U3052 (N_3052,In_1877,In_2125);
xor U3053 (N_3053,In_1062,In_408);
or U3054 (N_3054,In_724,In_666);
nand U3055 (N_3055,In_1618,In_1616);
and U3056 (N_3056,In_292,In_2411);
nor U3057 (N_3057,In_560,In_1325);
nand U3058 (N_3058,In_2337,In_49);
or U3059 (N_3059,In_1927,In_1462);
nor U3060 (N_3060,In_2496,In_1380);
xor U3061 (N_3061,In_580,In_551);
xor U3062 (N_3062,In_1495,In_2107);
xnor U3063 (N_3063,In_606,In_703);
nor U3064 (N_3064,In_1203,In_494);
xnor U3065 (N_3065,In_215,In_2246);
nor U3066 (N_3066,In_1042,In_882);
and U3067 (N_3067,In_2000,In_2351);
nand U3068 (N_3068,In_555,In_2455);
nor U3069 (N_3069,In_1082,In_1812);
or U3070 (N_3070,In_550,In_849);
nand U3071 (N_3071,In_1969,In_1605);
nand U3072 (N_3072,In_838,In_42);
and U3073 (N_3073,In_290,In_1200);
nand U3074 (N_3074,In_1547,In_1282);
or U3075 (N_3075,In_1320,In_920);
and U3076 (N_3076,In_1073,In_146);
xor U3077 (N_3077,In_869,In_75);
or U3078 (N_3078,In_411,In_1095);
nand U3079 (N_3079,In_1120,In_821);
xor U3080 (N_3080,In_652,In_26);
xor U3081 (N_3081,In_2451,In_1493);
nor U3082 (N_3082,In_1102,In_1593);
or U3083 (N_3083,In_2493,In_594);
and U3084 (N_3084,In_1008,In_1625);
xor U3085 (N_3085,In_867,In_1720);
xor U3086 (N_3086,In_820,In_1283);
xor U3087 (N_3087,In_1910,In_294);
nand U3088 (N_3088,In_967,In_368);
nand U3089 (N_3089,In_1054,In_1577);
nor U3090 (N_3090,In_1311,In_841);
nor U3091 (N_3091,In_2176,In_2336);
or U3092 (N_3092,In_597,In_2341);
or U3093 (N_3093,In_1154,In_1698);
nand U3094 (N_3094,In_2416,In_563);
nand U3095 (N_3095,In_2175,In_2228);
or U3096 (N_3096,In_2226,In_504);
xor U3097 (N_3097,In_559,In_414);
and U3098 (N_3098,In_1093,In_742);
nor U3099 (N_3099,In_2260,In_358);
nand U3100 (N_3100,In_1671,In_20);
nand U3101 (N_3101,In_68,In_1999);
nor U3102 (N_3102,In_1493,In_1611);
xor U3103 (N_3103,In_835,In_1298);
nor U3104 (N_3104,In_2478,In_2268);
nand U3105 (N_3105,In_1449,In_460);
and U3106 (N_3106,In_490,In_1470);
and U3107 (N_3107,In_1529,In_2423);
and U3108 (N_3108,In_2131,In_2030);
nor U3109 (N_3109,In_516,In_1691);
and U3110 (N_3110,In_425,In_2054);
nor U3111 (N_3111,In_250,In_2126);
and U3112 (N_3112,In_924,In_1666);
or U3113 (N_3113,In_1843,In_774);
and U3114 (N_3114,In_1054,In_1570);
nor U3115 (N_3115,In_12,In_1538);
nand U3116 (N_3116,In_2198,In_333);
and U3117 (N_3117,In_733,In_1080);
and U3118 (N_3118,In_1743,In_314);
xor U3119 (N_3119,In_2218,In_911);
nand U3120 (N_3120,In_1308,In_1136);
nand U3121 (N_3121,In_2091,In_166);
nand U3122 (N_3122,In_2208,In_503);
or U3123 (N_3123,In_539,In_182);
nand U3124 (N_3124,In_1402,In_1144);
xnor U3125 (N_3125,N_1347,N_1031);
nand U3126 (N_3126,N_3073,N_368);
nor U3127 (N_3127,N_1682,N_1806);
xor U3128 (N_3128,N_290,N_2487);
xor U3129 (N_3129,N_1913,N_1043);
nor U3130 (N_3130,N_2801,N_1679);
and U3131 (N_3131,N_935,N_1281);
nand U3132 (N_3132,N_2970,N_1760);
xnor U3133 (N_3133,N_2850,N_1571);
xnor U3134 (N_3134,N_576,N_2459);
nand U3135 (N_3135,N_396,N_690);
and U3136 (N_3136,N_2825,N_666);
nor U3137 (N_3137,N_1385,N_1631);
nand U3138 (N_3138,N_2642,N_2686);
nand U3139 (N_3139,N_670,N_2753);
or U3140 (N_3140,N_2506,N_990);
and U3141 (N_3141,N_411,N_2289);
or U3142 (N_3142,N_2169,N_1113);
nand U3143 (N_3143,N_2925,N_1795);
nor U3144 (N_3144,N_2582,N_162);
nor U3145 (N_3145,N_2629,N_916);
nand U3146 (N_3146,N_1002,N_2119);
xor U3147 (N_3147,N_209,N_2494);
nand U3148 (N_3148,N_2144,N_112);
or U3149 (N_3149,N_1250,N_37);
nand U3150 (N_3150,N_1363,N_1577);
nand U3151 (N_3151,N_1625,N_2823);
nand U3152 (N_3152,N_1070,N_2946);
nor U3153 (N_3153,N_1857,N_2658);
nand U3154 (N_3154,N_2124,N_1223);
or U3155 (N_3155,N_2226,N_2343);
or U3156 (N_3156,N_3042,N_2670);
xnor U3157 (N_3157,N_2295,N_1602);
nor U3158 (N_3158,N_2796,N_1620);
nor U3159 (N_3159,N_1697,N_383);
nor U3160 (N_3160,N_2117,N_249);
and U3161 (N_3161,N_1032,N_2942);
nor U3162 (N_3162,N_2348,N_1457);
xnor U3163 (N_3163,N_1337,N_2442);
and U3164 (N_3164,N_2517,N_951);
nor U3165 (N_3165,N_1816,N_1300);
nand U3166 (N_3166,N_2976,N_969);
xor U3167 (N_3167,N_2574,N_2473);
nand U3168 (N_3168,N_1506,N_1555);
or U3169 (N_3169,N_1288,N_3047);
nor U3170 (N_3170,N_2937,N_1196);
nor U3171 (N_3171,N_696,N_1238);
nand U3172 (N_3172,N_3003,N_1025);
or U3173 (N_3173,N_1659,N_315);
nand U3174 (N_3174,N_1447,N_2607);
nor U3175 (N_3175,N_2860,N_2725);
nand U3176 (N_3176,N_3059,N_321);
nor U3177 (N_3177,N_2519,N_848);
and U3178 (N_3178,N_2004,N_2088);
xnor U3179 (N_3179,N_2047,N_755);
nand U3180 (N_3180,N_634,N_2974);
or U3181 (N_3181,N_2278,N_1314);
nor U3182 (N_3182,N_3070,N_1943);
xnor U3183 (N_3183,N_159,N_2125);
nand U3184 (N_3184,N_344,N_508);
xor U3185 (N_3185,N_355,N_29);
and U3186 (N_3186,N_2560,N_809);
nor U3187 (N_3187,N_78,N_2965);
nand U3188 (N_3188,N_2094,N_2692);
and U3189 (N_3189,N_1080,N_2966);
and U3190 (N_3190,N_597,N_1428);
xor U3191 (N_3191,N_122,N_550);
or U3192 (N_3192,N_1882,N_635);
nor U3193 (N_3193,N_1282,N_563);
xnor U3194 (N_3194,N_347,N_950);
or U3195 (N_3195,N_2889,N_2528);
and U3196 (N_3196,N_1029,N_2208);
nor U3197 (N_3197,N_2844,N_1563);
or U3198 (N_3198,N_1218,N_1399);
and U3199 (N_3199,N_999,N_1634);
nor U3200 (N_3200,N_2997,N_844);
xnor U3201 (N_3201,N_2501,N_2312);
nand U3202 (N_3202,N_2795,N_1619);
or U3203 (N_3203,N_2783,N_1586);
xnor U3204 (N_3204,N_1729,N_1813);
and U3205 (N_3205,N_2379,N_907);
nand U3206 (N_3206,N_1064,N_2014);
nor U3207 (N_3207,N_762,N_1662);
xnor U3208 (N_3208,N_1011,N_1312);
nand U3209 (N_3209,N_2475,N_1996);
nor U3210 (N_3210,N_2490,N_3055);
xor U3211 (N_3211,N_998,N_2839);
nand U3212 (N_3212,N_1910,N_806);
nand U3213 (N_3213,N_136,N_240);
nand U3214 (N_3214,N_1158,N_747);
or U3215 (N_3215,N_2690,N_335);
or U3216 (N_3216,N_220,N_1712);
nor U3217 (N_3217,N_1986,N_2341);
nand U3218 (N_3218,N_19,N_2051);
or U3219 (N_3219,N_2485,N_2621);
and U3220 (N_3220,N_1397,N_2881);
or U3221 (N_3221,N_577,N_1187);
and U3222 (N_3222,N_2918,N_1511);
or U3223 (N_3223,N_2645,N_2986);
nor U3224 (N_3224,N_202,N_3037);
nand U3225 (N_3225,N_2427,N_1713);
nor U3226 (N_3226,N_46,N_1832);
nand U3227 (N_3227,N_1524,N_1854);
and U3228 (N_3228,N_312,N_2573);
or U3229 (N_3229,N_1472,N_1872);
or U3230 (N_3230,N_1933,N_2806);
and U3231 (N_3231,N_233,N_408);
nor U3232 (N_3232,N_3061,N_660);
nor U3233 (N_3233,N_764,N_2838);
or U3234 (N_3234,N_573,N_1042);
nand U3235 (N_3235,N_1408,N_2064);
or U3236 (N_3236,N_58,N_1800);
nor U3237 (N_3237,N_2050,N_1351);
and U3238 (N_3238,N_1975,N_307);
xor U3239 (N_3239,N_2428,N_614);
nand U3240 (N_3240,N_526,N_1426);
or U3241 (N_3241,N_1174,N_2044);
xor U3242 (N_3242,N_2352,N_783);
or U3243 (N_3243,N_2462,N_1019);
or U3244 (N_3244,N_2488,N_2274);
or U3245 (N_3245,N_1834,N_2276);
and U3246 (N_3246,N_2127,N_878);
or U3247 (N_3247,N_1100,N_2131);
or U3248 (N_3248,N_3013,N_9);
xnor U3249 (N_3249,N_2010,N_2548);
xor U3250 (N_3250,N_1690,N_1862);
nor U3251 (N_3251,N_1074,N_2283);
xnor U3252 (N_3252,N_946,N_1455);
or U3253 (N_3253,N_2882,N_1664);
nand U3254 (N_3254,N_1983,N_535);
xnor U3255 (N_3255,N_2852,N_2675);
and U3256 (N_3256,N_1692,N_2681);
nand U3257 (N_3257,N_1463,N_322);
and U3258 (N_3258,N_425,N_324);
xnor U3259 (N_3259,N_1893,N_1876);
xor U3260 (N_3260,N_3072,N_2515);
nand U3261 (N_3261,N_2189,N_919);
and U3262 (N_3262,N_113,N_2359);
nor U3263 (N_3263,N_164,N_285);
or U3264 (N_3264,N_1583,N_1299);
xor U3265 (N_3265,N_981,N_2677);
and U3266 (N_3266,N_2406,N_5);
xnor U3267 (N_3267,N_475,N_2721);
nor U3268 (N_3268,N_673,N_2985);
nor U3269 (N_3269,N_2614,N_2322);
and U3270 (N_3270,N_1459,N_241);
nand U3271 (N_3271,N_1992,N_207);
and U3272 (N_3272,N_832,N_1473);
nand U3273 (N_3273,N_2931,N_1791);
nand U3274 (N_3274,N_449,N_2719);
xnor U3275 (N_3275,N_774,N_874);
xor U3276 (N_3276,N_1564,N_849);
nand U3277 (N_3277,N_403,N_936);
nand U3278 (N_3278,N_967,N_1);
and U3279 (N_3279,N_609,N_2708);
nand U3280 (N_3280,N_1181,N_1120);
and U3281 (N_3281,N_704,N_2258);
nor U3282 (N_3282,N_2296,N_3038);
xor U3283 (N_3283,N_2268,N_2203);
xor U3284 (N_3284,N_984,N_323);
nand U3285 (N_3285,N_43,N_2045);
nand U3286 (N_3286,N_638,N_2869);
xnor U3287 (N_3287,N_1771,N_617);
nor U3288 (N_3288,N_1444,N_549);
nor U3289 (N_3289,N_1931,N_474);
xnor U3290 (N_3290,N_991,N_2038);
nand U3291 (N_3291,N_33,N_1086);
nand U3292 (N_3292,N_1920,N_2948);
nand U3293 (N_3293,N_146,N_2563);
and U3294 (N_3294,N_2957,N_1283);
nand U3295 (N_3295,N_1968,N_567);
or U3296 (N_3296,N_2867,N_3119);
or U3297 (N_3297,N_284,N_1302);
nand U3298 (N_3298,N_2593,N_412);
and U3299 (N_3299,N_640,N_732);
and U3300 (N_3300,N_2597,N_650);
nor U3301 (N_3301,N_1098,N_422);
or U3302 (N_3302,N_720,N_1378);
nor U3303 (N_3303,N_1318,N_1462);
or U3304 (N_3304,N_1681,N_738);
nor U3305 (N_3305,N_1142,N_2817);
and U3306 (N_3306,N_1323,N_1598);
and U3307 (N_3307,N_647,N_2437);
xnor U3308 (N_3308,N_1905,N_377);
or U3309 (N_3309,N_1203,N_1985);
nand U3310 (N_3310,N_2024,N_2697);
nand U3311 (N_3311,N_1179,N_1393);
nand U3312 (N_3312,N_2807,N_2327);
nand U3313 (N_3313,N_16,N_2320);
or U3314 (N_3314,N_678,N_600);
and U3315 (N_3315,N_3040,N_1915);
xnor U3316 (N_3316,N_1334,N_595);
and U3317 (N_3317,N_1478,N_862);
nand U3318 (N_3318,N_521,N_2687);
or U3319 (N_3319,N_2241,N_3054);
nand U3320 (N_3320,N_786,N_1821);
xnor U3321 (N_3321,N_2120,N_1280);
or U3322 (N_3322,N_333,N_194);
nor U3323 (N_3323,N_940,N_3116);
and U3324 (N_3324,N_2754,N_1494);
nand U3325 (N_3325,N_1267,N_2854);
or U3326 (N_3326,N_160,N_2553);
and U3327 (N_3327,N_118,N_1856);
nor U3328 (N_3328,N_2770,N_287);
nor U3329 (N_3329,N_258,N_1274);
nand U3330 (N_3330,N_2371,N_256);
xnor U3331 (N_3331,N_857,N_3033);
nor U3332 (N_3332,N_224,N_1287);
nor U3333 (N_3333,N_2461,N_797);
nand U3334 (N_3334,N_937,N_894);
xor U3335 (N_3335,N_997,N_2868);
nand U3336 (N_3336,N_2325,N_2037);
xor U3337 (N_3337,N_2056,N_1775);
and U3338 (N_3338,N_1306,N_2923);
and U3339 (N_3339,N_607,N_2902);
nand U3340 (N_3340,N_1183,N_889);
or U3341 (N_3341,N_0,N_1769);
nand U3342 (N_3342,N_693,N_1545);
xnor U3343 (N_3343,N_1830,N_2551);
nor U3344 (N_3344,N_2227,N_1143);
nor U3345 (N_3345,N_2846,N_2251);
nand U3346 (N_3346,N_1451,N_2405);
and U3347 (N_3347,N_1618,N_2565);
xnor U3348 (N_3348,N_877,N_3032);
xor U3349 (N_3349,N_2634,N_1296);
or U3350 (N_3350,N_2177,N_2451);
nand U3351 (N_3351,N_1249,N_1864);
nor U3352 (N_3352,N_1138,N_1796);
xor U3353 (N_3353,N_1212,N_445);
nor U3354 (N_3354,N_1809,N_565);
nor U3355 (N_3355,N_2618,N_291);
nor U3356 (N_3356,N_802,N_361);
nand U3357 (N_3357,N_1810,N_2123);
nand U3358 (N_3358,N_1526,N_1476);
nor U3359 (N_3359,N_2132,N_2435);
or U3360 (N_3360,N_1333,N_2007);
nand U3361 (N_3361,N_1401,N_1930);
nand U3362 (N_3362,N_392,N_1717);
and U3363 (N_3363,N_1305,N_1929);
nand U3364 (N_3364,N_821,N_1133);
and U3365 (N_3365,N_2142,N_2316);
and U3366 (N_3366,N_1112,N_30);
xnor U3367 (N_3367,N_2598,N_2450);
nor U3368 (N_3368,N_1246,N_116);
nor U3369 (N_3369,N_2480,N_834);
or U3370 (N_3370,N_460,N_3087);
or U3371 (N_3371,N_1997,N_2804);
or U3372 (N_3372,N_2091,N_662);
xnor U3373 (N_3373,N_2891,N_2178);
xor U3374 (N_3374,N_2353,N_102);
xnor U3375 (N_3375,N_1783,N_3123);
and U3376 (N_3376,N_2122,N_23);
xnor U3377 (N_3377,N_211,N_2481);
nor U3378 (N_3378,N_346,N_1723);
nand U3379 (N_3379,N_1927,N_1017);
nor U3380 (N_3380,N_1315,N_2972);
and U3381 (N_3381,N_1660,N_2562);
or U3382 (N_3382,N_2507,N_1977);
and U3383 (N_3383,N_1527,N_955);
xnor U3384 (N_3384,N_2166,N_2337);
nor U3385 (N_3385,N_2870,N_2375);
or U3386 (N_3386,N_639,N_578);
nand U3387 (N_3387,N_1234,N_94);
xnor U3388 (N_3388,N_781,N_866);
and U3389 (N_3389,N_238,N_1782);
or U3390 (N_3390,N_393,N_3012);
nor U3391 (N_3391,N_2601,N_2647);
xnor U3392 (N_3392,N_1685,N_229);
or U3393 (N_3393,N_1344,N_863);
xnor U3394 (N_3394,N_1419,N_1615);
or U3395 (N_3395,N_1268,N_274);
nor U3396 (N_3396,N_1826,N_1792);
xor U3397 (N_3397,N_2305,N_1388);
and U3398 (N_3398,N_329,N_450);
nor U3399 (N_3399,N_3083,N_574);
xor U3400 (N_3400,N_2205,N_267);
nor U3401 (N_3401,N_2383,N_702);
xor U3402 (N_3402,N_594,N_2408);
nand U3403 (N_3403,N_1627,N_2654);
and U3404 (N_3404,N_897,N_924);
and U3405 (N_3405,N_2254,N_1438);
xnor U3406 (N_3406,N_1192,N_2761);
and U3407 (N_3407,N_1121,N_2729);
or U3408 (N_3408,N_2361,N_444);
xor U3409 (N_3409,N_1114,N_1559);
and U3410 (N_3410,N_2637,N_1331);
and U3411 (N_3411,N_838,N_1343);
or U3412 (N_3412,N_751,N_2930);
and U3413 (N_3413,N_915,N_1962);
or U3414 (N_3414,N_2727,N_1722);
nand U3415 (N_3415,N_2537,N_237);
nor U3416 (N_3416,N_1295,N_1576);
nor U3417 (N_3417,N_1197,N_2530);
nand U3418 (N_3418,N_2349,N_1689);
and U3419 (N_3419,N_228,N_1761);
or U3420 (N_3420,N_363,N_2358);
xor U3421 (N_3421,N_2615,N_2498);
nor U3422 (N_3422,N_384,N_1349);
nor U3423 (N_3423,N_1982,N_1095);
or U3424 (N_3424,N_2061,N_1412);
nand U3425 (N_3425,N_1372,N_2040);
nand U3426 (N_3426,N_2221,N_2222);
nand U3427 (N_3427,N_186,N_2396);
xnor U3428 (N_3428,N_1879,N_625);
nand U3429 (N_3429,N_2228,N_2347);
or U3430 (N_3430,N_1237,N_458);
or U3431 (N_3431,N_629,N_2777);
xnor U3432 (N_3432,N_2610,N_2993);
and U3433 (N_3433,N_2586,N_2448);
nor U3434 (N_3434,N_1668,N_2155);
xnor U3435 (N_3435,N_2313,N_1411);
and U3436 (N_3436,N_2938,N_1354);
nand U3437 (N_3437,N_2156,N_1322);
or U3438 (N_3438,N_1518,N_1934);
xnor U3439 (N_3439,N_1122,N_2857);
and U3440 (N_3440,N_2999,N_398);
and U3441 (N_3441,N_993,N_2146);
or U3442 (N_3442,N_1051,N_1849);
xnor U3443 (N_3443,N_2875,N_547);
or U3444 (N_3444,N_871,N_1321);
and U3445 (N_3445,N_782,N_1415);
nor U3446 (N_3446,N_3105,N_2031);
nand U3447 (N_3447,N_2022,N_1648);
nand U3448 (N_3448,N_2663,N_3106);
nand U3449 (N_3449,N_366,N_579);
or U3450 (N_3450,N_1284,N_2995);
xor U3451 (N_3451,N_2556,N_1898);
nand U3452 (N_3452,N_1595,N_2963);
nor U3453 (N_3453,N_2855,N_1484);
nor U3454 (N_3454,N_487,N_184);
and U3455 (N_3455,N_3052,N_1846);
nand U3456 (N_3456,N_2608,N_1734);
nand U3457 (N_3457,N_1611,N_419);
nand U3458 (N_3458,N_1466,N_2886);
and U3459 (N_3459,N_562,N_2063);
nor U3460 (N_3460,N_502,N_369);
nor U3461 (N_3461,N_3063,N_36);
nor U3462 (N_3462,N_2785,N_2812);
and U3463 (N_3463,N_1759,N_1475);
and U3464 (N_3464,N_263,N_1776);
or U3465 (N_3465,N_1345,N_1159);
nand U3466 (N_3466,N_903,N_1693);
and U3467 (N_3467,N_1510,N_962);
and U3468 (N_3468,N_707,N_1079);
and U3469 (N_3469,N_712,N_973);
or U3470 (N_3470,N_2628,N_1632);
and U3471 (N_3471,N_2749,N_1189);
or U3472 (N_3472,N_929,N_1431);
nor U3473 (N_3473,N_519,N_1998);
nand U3474 (N_3474,N_176,N_1675);
nor U3475 (N_3475,N_451,N_1666);
xor U3476 (N_3476,N_1706,N_421);
xnor U3477 (N_3477,N_1779,N_2356);
or U3478 (N_3478,N_415,N_1087);
xnor U3479 (N_3479,N_182,N_1379);
xor U3480 (N_3480,N_1694,N_76);
nand U3481 (N_3481,N_1316,N_1464);
nand U3482 (N_3482,N_172,N_1413);
xnor U3483 (N_3483,N_628,N_2896);
xnor U3484 (N_3484,N_254,N_1450);
xor U3485 (N_3485,N_410,N_2924);
nor U3486 (N_3486,N_2390,N_2624);
nand U3487 (N_3487,N_1842,N_899);
or U3488 (N_3488,N_12,N_2984);
and U3489 (N_3489,N_85,N_1902);
nor U3490 (N_3490,N_2939,N_2602);
or U3491 (N_3491,N_2906,N_529);
or U3492 (N_3492,N_2872,N_2744);
and U3493 (N_3493,N_271,N_1037);
xnor U3494 (N_3494,N_1590,N_2763);
xor U3495 (N_3495,N_1878,N_402);
and U3496 (N_3496,N_1680,N_2192);
nand U3497 (N_3497,N_710,N_767);
and U3498 (N_3498,N_2443,N_2286);
nor U3499 (N_3499,N_340,N_1195);
and U3500 (N_3500,N_2367,N_811);
or U3501 (N_3501,N_676,N_497);
nor U3502 (N_3502,N_972,N_1990);
nor U3503 (N_3503,N_47,N_2874);
nand U3504 (N_3504,N_908,N_1885);
or U3505 (N_3505,N_2425,N_286);
nand U3506 (N_3506,N_2137,N_1802);
nand U3507 (N_3507,N_1755,N_986);
and U3508 (N_3508,N_1700,N_1044);
xor U3509 (N_3509,N_619,N_2831);
nand U3510 (N_3510,N_2118,N_120);
nor U3511 (N_3511,N_1926,N_2738);
or U3512 (N_3512,N_1391,N_1721);
or U3513 (N_3513,N_888,N_1007);
nor U3514 (N_3514,N_2136,N_1487);
nand U3515 (N_3515,N_2332,N_288);
or U3516 (N_3516,N_705,N_2008);
or U3517 (N_3517,N_2552,N_165);
and U3518 (N_3518,N_646,N_1736);
and U3519 (N_3519,N_1422,N_2696);
nor U3520 (N_3520,N_1210,N_2173);
nand U3521 (N_3521,N_1572,N_1848);
nand U3522 (N_3522,N_1708,N_1376);
xor U3523 (N_3523,N_2417,N_2300);
or U3524 (N_3524,N_2404,N_2255);
or U3525 (N_3525,N_482,N_356);
or U3526 (N_3526,N_3081,N_2101);
and U3527 (N_3527,N_569,N_1084);
xnor U3528 (N_3528,N_1912,N_1144);
xor U3529 (N_3529,N_2020,N_2774);
nand U3530 (N_3530,N_1871,N_1078);
and U3531 (N_3531,N_1400,N_31);
xnor U3532 (N_3532,N_1840,N_2247);
or U3533 (N_3533,N_2324,N_2168);
xnor U3534 (N_3534,N_455,N_191);
or U3535 (N_3535,N_1022,N_1724);
nor U3536 (N_3536,N_2062,N_2740);
nand U3537 (N_3537,N_1630,N_317);
xor U3538 (N_3538,N_2764,N_3099);
nand U3539 (N_3539,N_1904,N_128);
and U3540 (N_3540,N_1277,N_2438);
or U3541 (N_3541,N_2728,N_1719);
and U3542 (N_3542,N_1063,N_1161);
xnor U3543 (N_3543,N_1958,N_1528);
nand U3544 (N_3544,N_2385,N_2871);
nor U3545 (N_3545,N_41,N_2152);
and U3546 (N_3546,N_2926,N_2527);
or U3547 (N_3547,N_1099,N_2622);
and U3548 (N_3548,N_2059,N_1107);
xor U3549 (N_3549,N_1973,N_3);
xnor U3550 (N_3550,N_759,N_2077);
or U3551 (N_3551,N_1554,N_2220);
nor U3552 (N_3552,N_510,N_931);
nor U3553 (N_3553,N_1034,N_2603);
or U3554 (N_3554,N_837,N_2196);
nand U3555 (N_3555,N_1822,N_987);
nand U3556 (N_3556,N_1988,N_246);
or U3557 (N_3557,N_1134,N_669);
and U3558 (N_3558,N_2202,N_1895);
nor U3559 (N_3559,N_1900,N_3066);
and U3560 (N_3560,N_2755,N_1485);
nor U3561 (N_3561,N_1377,N_2837);
nor U3562 (N_3562,N_2246,N_928);
xnor U3563 (N_3563,N_370,N_2395);
xnor U3564 (N_3564,N_795,N_2828);
or U3565 (N_3565,N_2632,N_1916);
or U3566 (N_3566,N_1617,N_515);
or U3567 (N_3567,N_1263,N_1628);
nand U3568 (N_3568,N_1360,N_2787);
or U3569 (N_3569,N_840,N_2204);
or U3570 (N_3570,N_2589,N_1861);
or U3571 (N_3571,N_1654,N_1188);
nand U3572 (N_3572,N_2830,N_1823);
or U3573 (N_3573,N_394,N_3097);
nor U3574 (N_3574,N_1024,N_1432);
or U3575 (N_3575,N_2508,N_1006);
and U3576 (N_3576,N_2277,N_2102);
and U3577 (N_3577,N_2636,N_1647);
nand U3578 (N_3578,N_107,N_2611);
nand U3579 (N_3579,N_1945,N_824);
nor U3580 (N_3580,N_2950,N_1229);
and U3581 (N_3581,N_2546,N_91);
or U3582 (N_3582,N_1430,N_2030);
or U3583 (N_3583,N_2893,N_2167);
nor U3584 (N_3584,N_1616,N_733);
xnor U3585 (N_3585,N_2330,N_1383);
nand U3586 (N_3586,N_1062,N_2491);
and U3587 (N_3587,N_685,N_2033);
nor U3588 (N_3588,N_531,N_2892);
or U3589 (N_3589,N_2372,N_401);
or U3590 (N_3590,N_1153,N_201);
or U3591 (N_3591,N_3027,N_835);
or U3592 (N_3592,N_2680,N_2702);
and U3593 (N_3593,N_1993,N_295);
nor U3594 (N_3594,N_374,N_2111);
nor U3595 (N_3595,N_1458,N_1065);
nand U3596 (N_3596,N_719,N_942);
and U3597 (N_3597,N_2472,N_3108);
xor U3598 (N_3598,N_3046,N_1778);
or U3599 (N_3599,N_1715,N_1955);
or U3600 (N_3600,N_1794,N_293);
xor U3601 (N_3601,N_3095,N_3028);
nand U3602 (N_3602,N_390,N_2065);
xnor U3603 (N_3603,N_2531,N_1502);
nor U3604 (N_3604,N_1981,N_3077);
nor U3605 (N_3605,N_1606,N_108);
or U3606 (N_3606,N_2821,N_72);
and U3607 (N_3607,N_566,N_1937);
and U3608 (N_3608,N_1967,N_2661);
or U3609 (N_3609,N_2420,N_1172);
nor U3610 (N_3610,N_691,N_2224);
xor U3611 (N_3611,N_2130,N_703);
nand U3612 (N_3612,N_272,N_161);
or U3613 (N_3613,N_239,N_2429);
xnor U3614 (N_3614,N_2458,N_1808);
nor U3615 (N_3615,N_70,N_1398);
xnor U3616 (N_3616,N_1852,N_1402);
xor U3617 (N_3617,N_1552,N_2824);
and U3618 (N_3618,N_2713,N_413);
nand U3619 (N_3619,N_1655,N_2581);
and U3620 (N_3620,N_709,N_2894);
and U3621 (N_3621,N_2767,N_3004);
nand U3622 (N_3622,N_2584,N_2907);
and U3623 (N_3623,N_1850,N_28);
nand U3624 (N_3624,N_2662,N_372);
nor U3625 (N_3625,N_2055,N_1353);
nand U3626 (N_3626,N_2271,N_252);
nand U3627 (N_3627,N_551,N_2057);
xor U3628 (N_3628,N_2499,N_1317);
nand U3629 (N_3629,N_1233,N_1182);
xnor U3630 (N_3630,N_1493,N_2841);
and U3631 (N_3631,N_1566,N_2683);
nand U3632 (N_3632,N_2105,N_1049);
xor U3633 (N_3633,N_2818,N_469);
or U3634 (N_3634,N_1367,N_1053);
and U3635 (N_3635,N_311,N_1589);
nor U3636 (N_3636,N_2469,N_486);
or U3637 (N_3637,N_1247,N_716);
xnor U3638 (N_3638,N_2523,N_819);
nor U3639 (N_3639,N_243,N_1417);
or U3640 (N_3640,N_1932,N_427);
or U3641 (N_3641,N_2447,N_2028);
xor U3642 (N_3642,N_15,N_2141);
nand U3643 (N_3643,N_2034,N_1140);
xor U3644 (N_3644,N_1497,N_1674);
or U3645 (N_3645,N_1948,N_2758);
nor U3646 (N_3646,N_2793,N_730);
nand U3647 (N_3647,N_727,N_203);
nand U3648 (N_3648,N_1370,N_3076);
or U3649 (N_3649,N_416,N_2026);
nor U3650 (N_3650,N_2319,N_735);
nand U3651 (N_3651,N_2509,N_2306);
or U3652 (N_3652,N_1591,N_860);
xnor U3653 (N_3653,N_1711,N_1667);
and U3654 (N_3654,N_453,N_1865);
xnor U3655 (N_3655,N_627,N_2036);
nand U3656 (N_3656,N_659,N_1781);
or U3657 (N_3657,N_537,N_2769);
and U3658 (N_3658,N_183,N_2183);
or U3659 (N_3659,N_265,N_1340);
nand U3660 (N_3660,N_18,N_2525);
and U3661 (N_3661,N_99,N_2715);
and U3662 (N_3662,N_221,N_20);
xnor U3663 (N_3663,N_2138,N_407);
or U3664 (N_3664,N_2809,N_777);
and U3665 (N_3665,N_2600,N_1908);
or U3666 (N_3666,N_1480,N_437);
xor U3667 (N_3667,N_534,N_1407);
and U3668 (N_3668,N_1479,N_432);
nor U3669 (N_3669,N_190,N_2550);
nor U3670 (N_3670,N_2164,N_2842);
xnor U3671 (N_3671,N_820,N_130);
nor U3672 (N_3672,N_2099,N_3002);
nor U3673 (N_3673,N_2329,N_2266);
and U3674 (N_3674,N_1368,N_554);
or U3675 (N_3675,N_1683,N_2840);
or U3676 (N_3676,N_1108,N_477);
nor U3677 (N_3677,N_1762,N_2019);
xor U3678 (N_3678,N_2387,N_1449);
nand U3679 (N_3679,N_7,N_2025);
nand U3680 (N_3680,N_1060,N_804);
nand U3681 (N_3681,N_97,N_2717);
or U3682 (N_3682,N_829,N_606);
nand U3683 (N_3683,N_1529,N_216);
and U3684 (N_3684,N_2253,N_1088);
nor U3685 (N_3685,N_589,N_2170);
nor U3686 (N_3686,N_1240,N_1067);
nor U3687 (N_3687,N_75,N_2526);
xnor U3688 (N_3688,N_2545,N_616);
xnor U3689 (N_3689,N_1298,N_1585);
nand U3690 (N_3690,N_1285,N_892);
xor U3691 (N_3691,N_608,N_1339);
xor U3692 (N_3692,N_2920,N_543);
nor U3693 (N_3693,N_431,N_1012);
xnor U3694 (N_3694,N_2182,N_3092);
xnor U3695 (N_3695,N_3088,N_2722);
nor U3696 (N_3696,N_1866,N_957);
and U3697 (N_3697,N_1950,N_1116);
and U3698 (N_3698,N_2445,N_1477);
nor U3699 (N_3699,N_2350,N_3056);
or U3700 (N_3700,N_2412,N_197);
and U3701 (N_3701,N_813,N_328);
or U3702 (N_3702,N_1482,N_2653);
or U3703 (N_3703,N_1046,N_2159);
or U3704 (N_3704,N_788,N_2716);
or U3705 (N_3705,N_3017,N_2236);
or U3706 (N_3706,N_2078,N_144);
xor U3707 (N_3707,N_558,N_494);
and U3708 (N_3708,N_943,N_2465);
nor U3709 (N_3709,N_736,N_2188);
xor U3710 (N_3710,N_1010,N_2161);
nor U3711 (N_3711,N_2287,N_651);
xor U3712 (N_3712,N_269,N_2011);
nor U3713 (N_3713,N_1922,N_1102);
nand U3714 (N_3714,N_2592,N_2684);
or U3715 (N_3715,N_2452,N_699);
nor U3716 (N_3716,N_977,N_273);
xor U3717 (N_3717,N_1726,N_1709);
or U3718 (N_3718,N_2493,N_301);
xnor U3719 (N_3719,N_1405,N_1137);
nor U3720 (N_3720,N_556,N_397);
and U3721 (N_3721,N_2200,N_1358);
xor U3722 (N_3722,N_830,N_725);
nor U3723 (N_3723,N_1437,N_2235);
and U3724 (N_3724,N_2540,N_230);
or U3725 (N_3725,N_1365,N_109);
or U3726 (N_3726,N_2656,N_1784);
or U3727 (N_3727,N_1938,N_2261);
nor U3728 (N_3728,N_2726,N_816);
or U3729 (N_3729,N_1186,N_960);
nor U3730 (N_3730,N_1947,N_2175);
or U3731 (N_3731,N_1669,N_2256);
xor U3732 (N_3732,N_836,N_2016);
nor U3733 (N_3733,N_2765,N_2516);
or U3734 (N_3734,N_971,N_1961);
nor U3735 (N_3735,N_2272,N_1266);
and U3736 (N_3736,N_3078,N_461);
or U3737 (N_3737,N_248,N_389);
or U3738 (N_3738,N_530,N_796);
nor U3739 (N_3739,N_262,N_405);
and U3740 (N_3740,N_35,N_2561);
nand U3741 (N_3741,N_2298,N_40);
and U3742 (N_3742,N_2069,N_2265);
nor U3743 (N_3743,N_247,N_2505);
nand U3744 (N_3744,N_2583,N_1714);
and U3745 (N_3745,N_2604,N_1521);
nand U3746 (N_3746,N_2606,N_193);
and U3747 (N_3747,N_2756,N_1499);
nor U3748 (N_3748,N_1106,N_479);
and U3749 (N_3749,N_1738,N_893);
and U3750 (N_3750,N_1352,N_717);
nor U3751 (N_3751,N_135,N_2964);
nor U3752 (N_3752,N_2958,N_842);
nor U3753 (N_3753,N_2149,N_1470);
or U3754 (N_3754,N_586,N_1303);
xnor U3755 (N_3755,N_2668,N_332);
nand U3756 (N_3756,N_1128,N_48);
nor U3757 (N_3757,N_2967,N_2751);
and U3758 (N_3758,N_909,N_2888);
and U3759 (N_3759,N_1699,N_3103);
nor U3760 (N_3760,N_1505,N_1757);
or U3761 (N_3761,N_902,N_2810);
or U3762 (N_3762,N_1868,N_1939);
nand U3763 (N_3763,N_3080,N_1765);
nand U3764 (N_3764,N_668,N_2097);
nor U3765 (N_3765,N_1956,N_2153);
and U3766 (N_3766,N_2933,N_2039);
nor U3767 (N_3767,N_1805,N_778);
xor U3768 (N_3768,N_2724,N_1254);
xnor U3769 (N_3769,N_2479,N_1818);
or U3770 (N_3770,N_841,N_2922);
nor U3771 (N_3771,N_794,N_2143);
and U3772 (N_3772,N_1544,N_612);
or U3773 (N_3773,N_1819,N_61);
nand U3774 (N_3774,N_2945,N_689);
nor U3775 (N_3775,N_1536,N_2252);
or U3776 (N_3776,N_1141,N_2619);
nor U3777 (N_3777,N_158,N_418);
or U3778 (N_3778,N_1844,N_2557);
nor U3779 (N_3779,N_2106,N_2685);
or U3780 (N_3780,N_121,N_2865);
nor U3781 (N_3781,N_978,N_1211);
nand U3782 (N_3782,N_1057,N_1886);
xnor U3783 (N_3783,N_1242,N_2079);
nand U3784 (N_3784,N_1773,N_952);
and U3785 (N_3785,N_2544,N_1041);
xor U3786 (N_3786,N_917,N_2960);
nand U3787 (N_3787,N_2862,N_1336);
or U3788 (N_3788,N_2230,N_1687);
and U3789 (N_3789,N_655,N_1678);
nor U3790 (N_3790,N_1991,N_1255);
nor U3791 (N_3791,N_1015,N_2436);
nand U3792 (N_3792,N_1256,N_2431);
nand U3793 (N_3793,N_125,N_641);
or U3794 (N_3794,N_14,N_653);
xnor U3795 (N_3795,N_887,N_481);
nand U3796 (N_3796,N_2833,N_3084);
or U3797 (N_3797,N_1341,N_101);
and U3798 (N_3798,N_93,N_2836);
nand U3799 (N_3799,N_587,N_3006);
nor U3800 (N_3800,N_2085,N_3016);
and U3801 (N_3801,N_1691,N_850);
nand U3802 (N_3802,N_2899,N_1130);
nor U3803 (N_3803,N_2303,N_2370);
xor U3804 (N_3804,N_188,N_104);
nand U3805 (N_3805,N_2207,N_1767);
nand U3806 (N_3806,N_2794,N_86);
or U3807 (N_3807,N_2691,N_583);
xnor U3808 (N_3808,N_1350,N_858);
nor U3809 (N_3809,N_856,N_3098);
xnor U3810 (N_3810,N_1546,N_459);
or U3811 (N_3811,N_1665,N_1066);
nor U3812 (N_3812,N_1828,N_1863);
xnor U3813 (N_3813,N_1887,N_1395);
and U3814 (N_3814,N_467,N_768);
xnor U3815 (N_3815,N_695,N_1749);
xnor U3816 (N_3816,N_1160,N_259);
nand U3817 (N_3817,N_623,N_223);
or U3818 (N_3818,N_2631,N_2186);
or U3819 (N_3819,N_2197,N_1335);
xor U3820 (N_3820,N_1297,N_2905);
or U3821 (N_3821,N_3115,N_1157);
nor U3822 (N_3822,N_3020,N_1329);
nand U3823 (N_3823,N_1096,N_2968);
nand U3824 (N_3824,N_2991,N_3102);
and U3825 (N_3825,N_2386,N_2547);
and U3826 (N_3826,N_610,N_2240);
and U3827 (N_3827,N_1512,N_1168);
nand U3828 (N_3828,N_1202,N_1909);
and U3829 (N_3829,N_2244,N_2955);
xnor U3830 (N_3830,N_505,N_1059);
nor U3831 (N_3831,N_2802,N_1539);
and U3832 (N_3832,N_226,N_1733);
nor U3833 (N_3833,N_2304,N_3118);
or U3834 (N_3834,N_2943,N_1357);
xor U3835 (N_3835,N_2638,N_1790);
nor U3836 (N_3836,N_1741,N_1906);
nor U3837 (N_3837,N_2116,N_954);
nor U3838 (N_3838,N_2482,N_645);
nand U3839 (N_3839,N_718,N_2718);
nor U3840 (N_3840,N_544,N_553);
nand U3841 (N_3841,N_52,N_2989);
nand U3842 (N_3842,N_489,N_2075);
nor U3843 (N_3843,N_2492,N_514);
or U3844 (N_3844,N_171,N_2962);
nand U3845 (N_3845,N_1995,N_1979);
or U3846 (N_3846,N_2771,N_3048);
or U3847 (N_3847,N_2780,N_1313);
nand U3848 (N_3848,N_522,N_2301);
nor U3849 (N_3849,N_1440,N_2534);
nand U3850 (N_3850,N_2876,N_50);
nand U3851 (N_3851,N_1085,N_1292);
or U3852 (N_3852,N_2357,N_387);
or U3853 (N_3853,N_2210,N_665);
or U3854 (N_3854,N_1293,N_1807);
or U3855 (N_3855,N_2500,N_139);
xor U3856 (N_3856,N_1394,N_847);
nor U3857 (N_3857,N_1917,N_1443);
and U3858 (N_3858,N_309,N_167);
xnor U3859 (N_3859,N_1226,N_2921);
or U3860 (N_3860,N_2421,N_2665);
nor U3861 (N_3861,N_2736,N_365);
and U3862 (N_3862,N_1231,N_688);
nand U3863 (N_3863,N_1414,N_1009);
and U3864 (N_3864,N_464,N_2911);
nand U3865 (N_3865,N_2532,N_1446);
nor U3866 (N_3866,N_2904,N_1614);
or U3867 (N_3867,N_2422,N_2935);
and U3868 (N_3868,N_2981,N_1201);
or U3869 (N_3869,N_2376,N_1543);
or U3870 (N_3870,N_2049,N_473);
nand U3871 (N_3871,N_2843,N_992);
nor U3872 (N_3872,N_2659,N_375);
xnor U3873 (N_3873,N_706,N_1704);
xnor U3874 (N_3874,N_3111,N_898);
nand U3875 (N_3875,N_219,N_2791);
and U3876 (N_3876,N_80,N_3030);
nand U3877 (N_3877,N_1307,N_721);
nand U3878 (N_3878,N_513,N_1486);
nor U3879 (N_3879,N_302,N_2879);
nand U3880 (N_3880,N_349,N_404);
nand U3881 (N_3881,N_1047,N_585);
and U3882 (N_3882,N_1523,N_480);
xnor U3883 (N_3883,N_2851,N_1897);
xnor U3884 (N_3884,N_2988,N_442);
nor U3885 (N_3885,N_1608,N_2714);
nand U3886 (N_3886,N_3062,N_2160);
or U3887 (N_3887,N_2570,N_1574);
nand U3888 (N_3888,N_2399,N_1798);
nor U3889 (N_3889,N_2135,N_1152);
nor U3890 (N_3890,N_1797,N_1126);
nor U3891 (N_3891,N_584,N_2712);
or U3892 (N_3892,N_2695,N_348);
nand U3893 (N_3893,N_2826,N_2743);
nor U3894 (N_3894,N_2660,N_1014);
nand U3895 (N_3895,N_2463,N_199);
nand U3896 (N_3896,N_362,N_1200);
nand U3897 (N_3897,N_3029,N_1185);
nor U3898 (N_3898,N_1404,N_3074);
nor U3899 (N_3899,N_414,N_910);
and U3900 (N_3900,N_812,N_2384);
xnor U3901 (N_3901,N_298,N_456);
nand U3902 (N_3902,N_1504,N_745);
and U3903 (N_3903,N_2071,N_1971);
and U3904 (N_3904,N_1960,N_1101);
xor U3905 (N_3905,N_2762,N_2733);
or U3906 (N_3906,N_376,N_2820);
xnor U3907 (N_3907,N_961,N_590);
xnor U3908 (N_3908,N_1461,N_1568);
nand U3909 (N_3909,N_1003,N_1214);
nor U3910 (N_3910,N_1613,N_1241);
and U3911 (N_3911,N_166,N_793);
or U3912 (N_3912,N_3041,N_424);
nand U3913 (N_3913,N_1725,N_2772);
nand U3914 (N_3914,N_791,N_557);
or U3915 (N_3915,N_1582,N_1649);
nor U3916 (N_3916,N_698,N_1332);
and U3917 (N_3917,N_2987,N_2206);
xnor U3918 (N_3918,N_66,N_895);
nand U3919 (N_3919,N_2318,N_1841);
nor U3920 (N_3920,N_1671,N_926);
nand U3921 (N_3921,N_2426,N_289);
xor U3922 (N_3922,N_2524,N_2737);
xnor U3923 (N_3923,N_2310,N_1530);
xnor U3924 (N_3924,N_1170,N_2209);
xor U3925 (N_3925,N_2110,N_2778);
and U3926 (N_3926,N_2198,N_933);
xnor U3927 (N_3927,N_27,N_1677);
or U3928 (N_3928,N_282,N_3060);
or U3929 (N_3929,N_922,N_818);
nor U3930 (N_3930,N_814,N_1005);
xnor U3931 (N_3931,N_439,N_1963);
and U3932 (N_3932,N_331,N_989);
nand U3933 (N_3933,N_173,N_1592);
or U3934 (N_3934,N_436,N_2503);
xnor U3935 (N_3935,N_2502,N_1596);
and U3936 (N_3936,N_1000,N_339);
or U3937 (N_3937,N_140,N_2154);
and U3938 (N_3938,N_2800,N_84);
and U3939 (N_3939,N_1118,N_1278);
xnor U3940 (N_3940,N_1198,N_22);
nor U3941 (N_3941,N_3045,N_1944);
nor U3942 (N_3942,N_490,N_949);
xnor U3943 (N_3943,N_3085,N_2822);
or U3944 (N_3944,N_2368,N_723);
xor U3945 (N_3945,N_1004,N_523);
xnor U3946 (N_3946,N_575,N_980);
xor U3947 (N_3947,N_423,N_1491);
nor U3948 (N_3948,N_2474,N_2259);
nand U3949 (N_3949,N_105,N_1433);
nand U3950 (N_3950,N_2335,N_1753);
xor U3951 (N_3951,N_1974,N_2229);
nand U3952 (N_3952,N_351,N_1695);
and U3953 (N_3953,N_1883,N_843);
or U3954 (N_3954,N_54,N_345);
nand U3955 (N_3955,N_2979,N_2646);
nor U3956 (N_3956,N_1382,N_2863);
nand U3957 (N_3957,N_2699,N_498);
and U3958 (N_3958,N_261,N_2373);
or U3959 (N_3959,N_2956,N_2211);
nor U3960 (N_3960,N_3025,N_2798);
nor U3961 (N_3961,N_694,N_831);
xnor U3962 (N_3962,N_354,N_2449);
nand U3963 (N_3963,N_1801,N_2575);
xor U3964 (N_3964,N_2409,N_2566);
nand U3965 (N_3965,N_2076,N_1520);
nor U3966 (N_3966,N_2982,N_511);
and U3967 (N_3967,N_632,N_2978);
and U3968 (N_3968,N_1517,N_1213);
xnor U3969 (N_3969,N_1562,N_1940);
xnor U3970 (N_3970,N_1073,N_2486);
nand U3971 (N_3971,N_2250,N_1739);
nand U3972 (N_3972,N_68,N_527);
nand U3973 (N_3973,N_499,N_3015);
or U3974 (N_3974,N_2340,N_483);
nor U3975 (N_3975,N_2739,N_3124);
xor U3976 (N_3976,N_1094,N_371);
or U3977 (N_3977,N_2908,N_988);
or U3978 (N_3978,N_1039,N_1641);
xor U3979 (N_3979,N_2342,N_493);
xor U3980 (N_3980,N_1330,N_1999);
and U3981 (N_3981,N_815,N_2151);
nor U3982 (N_3982,N_2901,N_792);
xnor U3983 (N_3983,N_883,N_687);
nand U3984 (N_3984,N_212,N_1489);
xor U3985 (N_3985,N_142,N_1230);
xnor U3986 (N_3986,N_2973,N_891);
nand U3987 (N_3987,N_2710,N_1881);
nor U3988 (N_3988,N_938,N_2657);
xnor U3989 (N_3989,N_3000,N_2009);
xnor U3990 (N_3990,N_944,N_64);
or U3991 (N_3991,N_470,N_1732);
nor U3992 (N_3992,N_3069,N_3039);
nor U3993 (N_3993,N_2679,N_1252);
xor U3994 (N_3994,N_1270,N_2578);
nor U3995 (N_3995,N_1204,N_868);
xnor U3996 (N_3996,N_1232,N_457);
and U3997 (N_3997,N_1374,N_278);
nand U3998 (N_3998,N_1558,N_115);
nor U3999 (N_3999,N_1439,N_56);
and U4000 (N_4000,N_2873,N_89);
xor U4001 (N_4001,N_2070,N_746);
xor U4002 (N_4002,N_1980,N_2884);
nand U4003 (N_4003,N_2709,N_3086);
and U4004 (N_4004,N_2633,N_1789);
or U4005 (N_4005,N_501,N_1253);
xor U4006 (N_4006,N_1356,N_1756);
xor U4007 (N_4007,N_2466,N_1055);
or U4008 (N_4008,N_2776,N_1525);
and U4009 (N_4009,N_1847,N_2279);
xor U4010 (N_4010,N_1279,N_2887);
nor U4011 (N_4011,N_618,N_800);
or U4012 (N_4012,N_34,N_1058);
or U4013 (N_4013,N_1804,N_1342);
and U4014 (N_4014,N_1786,N_187);
nand U4015 (N_4015,N_642,N_196);
xnor U4016 (N_4016,N_1867,N_2157);
nand U4017 (N_4017,N_2620,N_429);
xor U4018 (N_4018,N_1166,N_2514);
nand U4019 (N_4019,N_2214,N_1894);
xnor U4020 (N_4020,N_622,N_148);
nor U4021 (N_4021,N_1215,N_2354);
xor U4022 (N_4022,N_1503,N_2434);
and U4023 (N_4023,N_1710,N_1556);
and U4024 (N_4024,N_2418,N_205);
or U4025 (N_4025,N_388,N_1097);
and U4026 (N_4026,N_2218,N_2441);
or U4027 (N_4027,N_1483,N_2936);
or U4028 (N_4028,N_2089,N_1635);
or U4029 (N_4029,N_552,N_236);
xor U4030 (N_4030,N_1171,N_44);
or U4031 (N_4031,N_1875,N_2457);
nand U4032 (N_4032,N_2323,N_2219);
or U4033 (N_4033,N_2021,N_3101);
nor U4034 (N_4034,N_825,N_1452);
nor U4035 (N_4035,N_1877,N_180);
nand U4036 (N_4036,N_1652,N_1946);
xnor U4037 (N_4037,N_1387,N_3026);
and U4038 (N_4038,N_1129,N_2932);
nor U4039 (N_4039,N_433,N_1780);
or U4040 (N_4040,N_1727,N_2595);
nand U4041 (N_4041,N_1540,N_496);
and U4042 (N_4042,N_250,N_3031);
nand U4043 (N_4043,N_381,N_602);
nor U4044 (N_4044,N_2308,N_2934);
or U4045 (N_4045,N_1838,N_996);
nand U4046 (N_4046,N_525,N_1173);
nand U4047 (N_4047,N_1071,N_2667);
xor U4048 (N_4048,N_2344,N_283);
nor U4049 (N_4049,N_766,N_630);
and U4050 (N_4050,N_2245,N_2217);
and U4051 (N_4051,N_1626,N_900);
and U4052 (N_4052,N_2195,N_2134);
xor U4053 (N_4053,N_2834,N_1703);
or U4054 (N_4054,N_1903,N_621);
xnor U4055 (N_4055,N_2098,N_1987);
nor U4056 (N_4056,N_1474,N_739);
or U4057 (N_4057,N_2649,N_382);
or U4058 (N_4058,N_2092,N_2928);
nor U4059 (N_4059,N_463,N_2510);
xnor U4060 (N_4060,N_2814,N_948);
or U4061 (N_4061,N_65,N_3094);
nor U4062 (N_4062,N_1359,N_2723);
nand U4063 (N_4063,N_2706,N_1766);
nand U4064 (N_4064,N_303,N_1371);
or U4065 (N_4065,N_2393,N_448);
or U4066 (N_4066,N_714,N_677);
or U4067 (N_4067,N_152,N_1758);
nand U4068 (N_4068,N_1964,N_861);
nand U4069 (N_4069,N_2571,N_568);
or U4070 (N_4070,N_1036,N_2513);
or U4071 (N_4071,N_1275,N_2407);
and U4072 (N_4072,N_1206,N_45);
nand U4073 (N_4073,N_2671,N_1220);
nor U4074 (N_4074,N_1573,N_96);
xor U4075 (N_4075,N_1410,N_637);
nor U4076 (N_4076,N_1396,N_1456);
nor U4077 (N_4077,N_1645,N_1501);
xnor U4078 (N_4078,N_851,N_1825);
nand U4079 (N_4079,N_1111,N_1115);
xnor U4080 (N_4080,N_1465,N_2360);
xnor U4081 (N_4081,N_896,N_743);
or U4082 (N_4082,N_2704,N_446);
or U4083 (N_4083,N_1441,N_296);
and U4084 (N_4084,N_1860,N_2816);
or U4085 (N_4085,N_3009,N_1406);
and U4086 (N_4086,N_2478,N_1835);
and U4087 (N_4087,N_435,N_1445);
nor U4088 (N_4088,N_1272,N_2616);
nor U4089 (N_4089,N_1567,N_2835);
and U4090 (N_4090,N_2107,N_400);
nor U4091 (N_4091,N_2380,N_1656);
xnor U4092 (N_4092,N_1953,N_1911);
nor U4093 (N_4093,N_3065,N_2060);
xor U4094 (N_4094,N_593,N_1820);
nor U4095 (N_4095,N_604,N_930);
nand U4096 (N_4096,N_1208,N_77);
xor U4097 (N_4097,N_1629,N_1324);
nor U4098 (N_4098,N_1175,N_1599);
or U4099 (N_4099,N_845,N_890);
nand U4100 (N_4100,N_1770,N_1038);
or U4101 (N_4101,N_1533,N_875);
xor U4102 (N_4102,N_1839,N_2609);
xnor U4103 (N_4103,N_2364,N_1748);
nand U4104 (N_4104,N_1570,N_914);
nor U4105 (N_4105,N_3109,N_1327);
xnor U4106 (N_4106,N_1508,N_395);
nand U4107 (N_4107,N_1467,N_772);
and U4108 (N_4108,N_1221,N_2864);
nor U4109 (N_4109,N_2003,N_1702);
or U4110 (N_4110,N_1403,N_26);
and U4111 (N_4111,N_1320,N_911);
or U4112 (N_4112,N_1774,N_62);
or U4113 (N_4113,N_654,N_2959);
xnor U4114 (N_4114,N_1752,N_953);
nand U4115 (N_4115,N_2735,N_982);
nor U4116 (N_4116,N_3021,N_1448);
or U4117 (N_4117,N_2470,N_1672);
xor U4118 (N_4118,N_2567,N_264);
and U4119 (N_4119,N_2927,N_779);
or U4120 (N_4120,N_1560,N_2700);
and U4121 (N_4121,N_2543,N_886);
and U4122 (N_4122,N_1870,N_1442);
and U4123 (N_4123,N_1924,N_855);
nor U4124 (N_4124,N_2262,N_1673);
xnor U4125 (N_4125,N_701,N_2760);
nand U4126 (N_4126,N_1083,N_1896);
and U4127 (N_4127,N_2898,N_337);
nor U4128 (N_4128,N_292,N_1742);
nand U4129 (N_4129,N_1286,N_1650);
and U4130 (N_4130,N_963,N_675);
or U4131 (N_4131,N_1045,N_1787);
or U4132 (N_4132,N_995,N_1361);
and U4133 (N_4133,N_2374,N_170);
or U4134 (N_4134,N_631,N_1271);
nand U4135 (N_4135,N_2747,N_90);
xnor U4136 (N_4136,N_1077,N_555);
and U4137 (N_4137,N_2915,N_1216);
and U4138 (N_4138,N_214,N_2994);
and U4139 (N_4139,N_682,N_1743);
nor U4140 (N_4140,N_1061,N_1720);
nand U4141 (N_4141,N_2940,N_492);
and U4142 (N_4142,N_2859,N_964);
and U4143 (N_4143,N_2977,N_1859);
and U4144 (N_4144,N_1507,N_1338);
nand U4145 (N_4145,N_2000,N_2803);
nand U4146 (N_4146,N_359,N_1209);
or U4147 (N_4147,N_3064,N_1224);
nor U4148 (N_4148,N_1532,N_686);
xnor U4149 (N_4149,N_24,N_1768);
nor U4150 (N_4150,N_1471,N_2121);
nand U4151 (N_4151,N_1548,N_2415);
or U4152 (N_4152,N_2365,N_2520);
or U4153 (N_4153,N_2919,N_2811);
and U4154 (N_4154,N_2237,N_2961);
or U4155 (N_4155,N_1519,N_2162);
or U4156 (N_4156,N_342,N_60);
nand U4157 (N_4157,N_1425,N_2238);
and U4158 (N_4158,N_1698,N_13);
nor U4159 (N_4159,N_1132,N_2275);
and U4160 (N_4160,N_760,N_1799);
or U4161 (N_4161,N_1728,N_872);
nand U4162 (N_4162,N_218,N_2288);
or U4163 (N_4163,N_304,N_2827);
nand U4164 (N_4164,N_3121,N_378);
and U4165 (N_4165,N_1131,N_1290);
xor U4166 (N_4166,N_1584,N_2788);
and U4167 (N_4167,N_867,N_2402);
and U4168 (N_4168,N_1219,N_103);
xnor U4169 (N_4169,N_592,N_327);
nor U4170 (N_4170,N_652,N_1355);
nand U4171 (N_4171,N_1610,N_3082);
and U4172 (N_4172,N_974,N_1646);
nand U4173 (N_4173,N_985,N_1537);
xor U4174 (N_4174,N_2512,N_2260);
xnor U4175 (N_4175,N_927,N_2046);
or U4176 (N_4176,N_150,N_2);
xor U4177 (N_4177,N_2270,N_1918);
and U4178 (N_4178,N_1369,N_1105);
and U4179 (N_4179,N_1607,N_2847);
and U4180 (N_4180,N_3035,N_443);
nand U4181 (N_4181,N_1264,N_649);
and U4182 (N_4182,N_3071,N_611);
xnor U4183 (N_4183,N_100,N_343);
or U4184 (N_4184,N_671,N_305);
nor U4185 (N_4185,N_2269,N_1976);
nand U4186 (N_4186,N_1972,N_1541);
xnor U4187 (N_4187,N_1978,N_2048);
and U4188 (N_4188,N_994,N_2067);
nor U4189 (N_4189,N_320,N_2397);
or U4190 (N_4190,N_1190,N_2233);
and U4191 (N_4191,N_1604,N_1688);
and U4192 (N_4192,N_2651,N_1837);
or U4193 (N_4193,N_260,N_965);
and U4194 (N_4194,N_1104,N_1542);
and U4195 (N_4195,N_1346,N_2066);
nand U4196 (N_4196,N_67,N_3091);
and U4197 (N_4197,N_1248,N_1436);
and U4198 (N_4198,N_2655,N_2456);
nor U4199 (N_4199,N_2133,N_1035);
xor U4200 (N_4200,N_1460,N_2018);
nor U4201 (N_4201,N_765,N_2239);
xnor U4202 (N_4202,N_2058,N_876);
nand U4203 (N_4203,N_2440,N_2012);
or U4204 (N_4204,N_1994,N_925);
and U4205 (N_4205,N_1579,N_4);
nor U4206 (N_4206,N_2171,N_1925);
and U4207 (N_4207,N_1565,N_2766);
xnor U4208 (N_4208,N_2705,N_3007);
or U4209 (N_4209,N_2095,N_210);
nand U4210 (N_4210,N_57,N_1891);
nor U4211 (N_4211,N_1954,N_1434);
nor U4212 (N_4212,N_524,N_2381);
xnor U4213 (N_4213,N_1957,N_149);
and U4214 (N_4214,N_1636,N_620);
and U4215 (N_4215,N_1156,N_2912);
xnor U4216 (N_4216,N_2005,N_2231);
or U4217 (N_4217,N_2355,N_1984);
xnor U4218 (N_4218,N_2853,N_853);
xnor U4219 (N_4219,N_1273,N_520);
and U4220 (N_4220,N_2293,N_2346);
or U4221 (N_4221,N_2391,N_1763);
and U4222 (N_4222,N_1594,N_1609);
xor U4223 (N_4223,N_2669,N_1869);
and U4224 (N_4224,N_752,N_1244);
nand U4225 (N_4225,N_2549,N_2083);
or U4226 (N_4226,N_3019,N_2109);
or U4227 (N_4227,N_3090,N_2627);
xor U4228 (N_4228,N_1731,N_1772);
and U4229 (N_4229,N_912,N_1392);
and U4230 (N_4230,N_538,N_2720);
and U4231 (N_4231,N_2084,N_854);
nand U4232 (N_4232,N_2856,N_648);
or U4233 (N_4233,N_2890,N_906);
or U4234 (N_4234,N_2650,N_2273);
or U4235 (N_4235,N_758,N_2232);
xnor U4236 (N_4236,N_2223,N_2023);
nor U4237 (N_4237,N_1764,N_2741);
xnor U4238 (N_4238,N_2797,N_3114);
xor U4239 (N_4239,N_1076,N_1531);
nand U4240 (N_4240,N_63,N_2317);
xor U4241 (N_4241,N_1030,N_2483);
and U4242 (N_4242,N_1553,N_2328);
nand U4243 (N_4243,N_503,N_380);
nand U4244 (N_4244,N_117,N_1492);
nand U4245 (N_4245,N_966,N_2903);
nand U4246 (N_4246,N_2476,N_1707);
and U4247 (N_4247,N_1481,N_1109);
nand U4248 (N_4248,N_3010,N_1569);
and U4249 (N_4249,N_1193,N_485);
nor U4250 (N_4250,N_3117,N_2292);
or U4251 (N_4251,N_2388,N_318);
and U4252 (N_4252,N_484,N_462);
xnor U4253 (N_4253,N_1663,N_1364);
nor U4254 (N_4254,N_379,N_2555);
nor U4255 (N_4255,N_681,N_2302);
or U4256 (N_4256,N_1149,N_975);
nor U4257 (N_4257,N_3057,N_1427);
nand U4258 (N_4258,N_454,N_644);
xor U4259 (N_4259,N_582,N_728);
and U4260 (N_4260,N_1914,N_310);
nor U4261 (N_4261,N_3043,N_1637);
xnor U4262 (N_4262,N_1843,N_129);
nand U4263 (N_4263,N_2533,N_306);
nand U4264 (N_4264,N_958,N_2895);
or U4265 (N_4265,N_471,N_2439);
nor U4266 (N_4266,N_724,N_1884);
and U4267 (N_4267,N_1803,N_546);
and U4268 (N_4268,N_1969,N_59);
xor U4269 (N_4269,N_192,N_882);
or U4270 (N_4270,N_1262,N_979);
xor U4271 (N_4271,N_1424,N_6);
or U4272 (N_4272,N_2382,N_1827);
nor U4273 (N_4273,N_21,N_939);
or U4274 (N_4274,N_1228,N_757);
or U4275 (N_4275,N_1243,N_934);
nand U4276 (N_4276,N_1547,N_2336);
and U4277 (N_4277,N_2949,N_3079);
and U4278 (N_4278,N_2630,N_1588);
nor U4279 (N_4279,N_2446,N_1815);
and U4280 (N_4280,N_1048,N_1180);
nand U4281 (N_4281,N_2194,N_1888);
or U4282 (N_4282,N_697,N_2635);
xor U4283 (N_4283,N_2282,N_2591);
xor U4284 (N_4284,N_1311,N_2464);
or U4285 (N_4285,N_313,N_2080);
xnor U4286 (N_4286,N_1522,N_1686);
or U4287 (N_4287,N_1580,N_1633);
nand U4288 (N_4288,N_598,N_334);
and U4289 (N_4289,N_1301,N_2554);
xnor U4290 (N_4290,N_2511,N_2773);
nor U4291 (N_4291,N_2489,N_846);
xor U4292 (N_4292,N_826,N_88);
or U4293 (N_4293,N_2163,N_2613);
or U4294 (N_4294,N_279,N_1169);
xnor U4295 (N_4295,N_2990,N_1033);
nand U4296 (N_4296,N_2366,N_2535);
nor U4297 (N_4297,N_918,N_3107);
or U4298 (N_4298,N_2805,N_2053);
and U4299 (N_4299,N_1205,N_2433);
nand U4300 (N_4300,N_805,N_1550);
or U4301 (N_4301,N_2052,N_873);
and U4302 (N_4302,N_2913,N_1375);
nor U4303 (N_4303,N_1154,N_3034);
or U4304 (N_4304,N_1639,N_881);
nand U4305 (N_4305,N_561,N_658);
and U4306 (N_4306,N_1513,N_1587);
nand U4307 (N_4307,N_2181,N_1389);
or U4308 (N_4308,N_870,N_2212);
nor U4309 (N_4309,N_2419,N_2880);
nand U4310 (N_4310,N_200,N_428);
nor U4311 (N_4311,N_2249,N_385);
and U4312 (N_4312,N_2176,N_69);
or U4313 (N_4313,N_2732,N_98);
and U4314 (N_4314,N_2129,N_2746);
and U4315 (N_4315,N_106,N_10);
nand U4316 (N_4316,N_154,N_801);
xor U4317 (N_4317,N_1075,N_1294);
and U4318 (N_4318,N_245,N_2569);
nand U4319 (N_4319,N_1718,N_1581);
nor U4320 (N_4320,N_2542,N_2799);
xnor U4321 (N_4321,N_2042,N_2423);
and U4322 (N_4322,N_680,N_2676);
xnor U4323 (N_4323,N_3014,N_1676);
and U4324 (N_4324,N_2389,N_1225);
and U4325 (N_4325,N_1135,N_1269);
or U4326 (N_4326,N_2297,N_386);
or U4327 (N_4327,N_599,N_2682);
xnor U4328 (N_4328,N_1750,N_1258);
nor U4329 (N_4329,N_1072,N_124);
and U4330 (N_4330,N_3067,N_810);
xor U4331 (N_4331,N_2017,N_1239);
nand U4332 (N_4332,N_1409,N_884);
nor U4333 (N_4333,N_3011,N_1251);
and U4334 (N_4334,N_1309,N_270);
and U4335 (N_4335,N_488,N_74);
nand U4336 (N_4336,N_1966,N_2742);
and U4337 (N_4337,N_2688,N_42);
or U4338 (N_4338,N_157,N_2035);
or U4339 (N_4339,N_257,N_603);
xor U4340 (N_4340,N_71,N_2392);
nor U4341 (N_4341,N_3053,N_731);
or U4342 (N_4342,N_2191,N_784);
or U4343 (N_4343,N_1538,N_1091);
and U4344 (N_4344,N_251,N_2529);
nor U4345 (N_4345,N_2707,N_1235);
or U4346 (N_4346,N_1139,N_748);
nor U4347 (N_4347,N_2299,N_2640);
xnor U4348 (N_4348,N_1824,N_3089);
nand U4349 (N_4349,N_2594,N_83);
and U4350 (N_4350,N_2032,N_839);
xnor U4351 (N_4351,N_833,N_1390);
nor U4352 (N_4352,N_807,N_2580);
nor U4353 (N_4353,N_1194,N_2126);
or U4354 (N_4354,N_1735,N_528);
or U4355 (N_4355,N_1468,N_163);
xor U4356 (N_4356,N_87,N_2086);
or U4357 (N_4357,N_1622,N_3036);
xnor U4358 (N_4358,N_2264,N_360);
or U4359 (N_4359,N_2698,N_968);
and U4360 (N_4360,N_2750,N_2243);
xnor U4361 (N_4361,N_1136,N_3008);
or U4362 (N_4362,N_2664,N_195);
or U4363 (N_4363,N_225,N_2792);
nor U4364 (N_4364,N_1578,N_2484);
and U4365 (N_4365,N_1970,N_2752);
or U4366 (N_4366,N_38,N_111);
or U4367 (N_4367,N_726,N_1148);
nand U4368 (N_4368,N_114,N_1746);
nor U4369 (N_4369,N_1167,N_2013);
and U4370 (N_4370,N_545,N_2496);
nand U4371 (N_4371,N_1420,N_780);
xnor U4372 (N_4372,N_2641,N_2087);
and U4373 (N_4373,N_2866,N_3068);
and U4374 (N_4374,N_3075,N_2730);
or U4375 (N_4375,N_2455,N_391);
and U4376 (N_4376,N_1495,N_1090);
nor U4377 (N_4377,N_1276,N_1001);
and U4378 (N_4378,N_2002,N_2568);
and U4379 (N_4379,N_2073,N_2858);
xor U4380 (N_4380,N_2165,N_729);
xor U4381 (N_4381,N_232,N_1601);
or U4382 (N_4382,N_947,N_2910);
nor U4383 (N_4383,N_2104,N_1855);
xor U4384 (N_4384,N_55,N_2941);
and U4385 (N_4385,N_95,N_2257);
xor U4386 (N_4386,N_2263,N_440);
and U4387 (N_4387,N_970,N_1366);
or U4388 (N_4388,N_1310,N_1624);
xor U4389 (N_4389,N_1643,N_2861);
nor U4390 (N_4390,N_548,N_692);
and U4391 (N_4391,N_2432,N_2112);
nor U4392 (N_4392,N_2331,N_1638);
or U4393 (N_4393,N_2471,N_447);
xnor U4394 (N_4394,N_1227,N_2454);
nand U4395 (N_4395,N_1651,N_2775);
and U4396 (N_4396,N_2768,N_73);
and U4397 (N_4397,N_1217,N_2617);
nand U4398 (N_4398,N_588,N_905);
or U4399 (N_4399,N_572,N_1081);
or U4400 (N_4400,N_715,N_823);
and U4401 (N_4401,N_134,N_2199);
or U4402 (N_4402,N_147,N_2128);
nand U4403 (N_4403,N_336,N_1103);
or U4404 (N_4404,N_1653,N_49);
xor U4405 (N_4405,N_1696,N_299);
nor U4406 (N_4406,N_1928,N_1236);
nand U4407 (N_4407,N_2072,N_1788);
nand U4408 (N_4408,N_2784,N_2579);
xnor U4409 (N_4409,N_2703,N_1534);
xnor U4410 (N_4410,N_126,N_2248);
nand U4411 (N_4411,N_1535,N_1089);
and U4412 (N_4412,N_253,N_700);
xor U4413 (N_4413,N_1701,N_2944);
xnor U4414 (N_4414,N_1851,N_1814);
nor U4415 (N_4415,N_2980,N_754);
or U4416 (N_4416,N_749,N_2113);
and U4417 (N_4417,N_799,N_822);
or U4418 (N_4418,N_2759,N_2185);
nor U4419 (N_4419,N_540,N_3018);
nor U4420 (N_4420,N_517,N_2225);
nand U4421 (N_4421,N_2201,N_110);
and U4422 (N_4422,N_2315,N_1716);
and U4423 (N_4423,N_2401,N_409);
or U4424 (N_4424,N_2029,N_133);
and U4425 (N_4425,N_1040,N_2280);
nor U4426 (N_4426,N_2644,N_1811);
nand U4427 (N_4427,N_1640,N_1747);
nand U4428 (N_4428,N_1561,N_2639);
and U4429 (N_4429,N_2648,N_275);
nor U4430 (N_4430,N_2521,N_679);
or U4431 (N_4431,N_1600,N_1326);
or U4432 (N_4432,N_1829,N_1056);
and U4433 (N_4433,N_466,N_2345);
nor U4434 (N_4434,N_2100,N_3051);
nand U4435 (N_4435,N_2522,N_217);
and U4436 (N_4436,N_817,N_1093);
nor U4437 (N_4437,N_2307,N_2954);
or U4438 (N_4438,N_945,N_179);
nor U4439 (N_4439,N_2587,N_2678);
xnor U4440 (N_4440,N_1245,N_2477);
nor U4441 (N_4441,N_308,N_753);
xor U4442 (N_4442,N_2914,N_2808);
nand U4443 (N_4443,N_2734,N_643);
xor U4444 (N_4444,N_155,N_532);
nand U4445 (N_4445,N_2213,N_406);
nand U4446 (N_4446,N_2947,N_2813);
nor U4447 (N_4447,N_2789,N_2082);
nor U4448 (N_4448,N_2596,N_2605);
or U4449 (N_4449,N_2453,N_156);
xor U4450 (N_4450,N_119,N_168);
nand U4451 (N_4451,N_591,N_2314);
and U4452 (N_4452,N_1705,N_2541);
xor U4453 (N_4453,N_1191,N_1418);
or U4454 (N_4454,N_314,N_1751);
nand U4455 (N_4455,N_3005,N_2400);
and U4456 (N_4456,N_920,N_1373);
nor U4457 (N_4457,N_268,N_2588);
xnor U4458 (N_4458,N_785,N_636);
and U4459 (N_4459,N_2623,N_2689);
or U4460 (N_4460,N_79,N_1261);
nand U4461 (N_4461,N_2674,N_789);
nor U4462 (N_4462,N_1812,N_3113);
and U4463 (N_4463,N_1381,N_2090);
xnor U4464 (N_4464,N_2114,N_2917);
xor U4465 (N_4465,N_3001,N_541);
and U4466 (N_4466,N_869,N_1509);
nand U4467 (N_4467,N_1575,N_2369);
and U4468 (N_4468,N_198,N_281);
or U4469 (N_4469,N_1423,N_2460);
nand U4470 (N_4470,N_2673,N_3044);
or U4471 (N_4471,N_1018,N_1496);
or U4472 (N_4472,N_2694,N_683);
or U4473 (N_4473,N_667,N_1901);
or U4474 (N_4474,N_2819,N_367);
nor U4475 (N_4475,N_1935,N_533);
nand U4476 (N_4476,N_742,N_879);
nand U4477 (N_4477,N_708,N_1551);
or U4478 (N_4478,N_1257,N_2585);
xor U4479 (N_4479,N_2093,N_1959);
nand U4480 (N_4480,N_1921,N_512);
or U4481 (N_4481,N_615,N_2897);
or U4482 (N_4482,N_901,N_3022);
xor U4483 (N_4483,N_769,N_2779);
nor U4484 (N_4484,N_2929,N_1026);
xnor U4485 (N_4485,N_2539,N_2564);
or U4486 (N_4486,N_2416,N_2190);
nand U4487 (N_4487,N_1740,N_2883);
or U4488 (N_4488,N_983,N_1658);
and U4489 (N_4489,N_613,N_1989);
nand U4490 (N_4490,N_2577,N_2572);
xnor U4491 (N_4491,N_1199,N_2626);
nand U4492 (N_4492,N_2403,N_941);
nor U4493 (N_4493,N_2590,N_2672);
or U4494 (N_4494,N_2786,N_1222);
xnor U4495 (N_4495,N_1127,N_2996);
and U4496 (N_4496,N_1670,N_1027);
nor U4497 (N_4497,N_2139,N_2748);
nand U4498 (N_4498,N_865,N_828);
nor U4499 (N_4499,N_2180,N_1054);
and U4500 (N_4500,N_1949,N_2559);
nor U4501 (N_4501,N_2311,N_1021);
nand U4502 (N_4502,N_2321,N_316);
xor U4503 (N_4503,N_506,N_1919);
nor U4504 (N_4504,N_1429,N_2900);
or U4505 (N_4505,N_235,N_153);
nand U4506 (N_4506,N_1050,N_859);
nand U4507 (N_4507,N_1068,N_1936);
nor U4508 (N_4508,N_465,N_1612);
or U4509 (N_4509,N_2643,N_92);
or U4510 (N_4510,N_1308,N_923);
nand U4511 (N_4511,N_771,N_2362);
nand U4512 (N_4512,N_2179,N_2148);
nand U4513 (N_4513,N_185,N_2410);
nor U4514 (N_4514,N_326,N_885);
or U4515 (N_4515,N_127,N_2701);
nor U4516 (N_4516,N_2538,N_2878);
xor U4517 (N_4517,N_3024,N_2174);
nand U4518 (N_4518,N_1416,N_2398);
xnor U4519 (N_4519,N_773,N_53);
and U4520 (N_4520,N_1793,N_1836);
xnor U4521 (N_4521,N_1421,N_1923);
nand U4522 (N_4522,N_1899,N_2150);
and U4523 (N_4523,N_426,N_2334);
and U4524 (N_4524,N_2285,N_664);
or U4525 (N_4525,N_2599,N_276);
nor U4526 (N_4526,N_674,N_770);
or U4527 (N_4527,N_208,N_1023);
xor U4528 (N_4528,N_1454,N_1892);
or U4529 (N_4529,N_626,N_672);
nand U4530 (N_4530,N_132,N_3100);
or U4531 (N_4531,N_663,N_1833);
and U4532 (N_4532,N_500,N_3110);
xor U4533 (N_4533,N_277,N_2333);
and U4534 (N_4534,N_2339,N_169);
nand U4535 (N_4535,N_2909,N_1016);
and U4536 (N_4536,N_357,N_472);
nor U4537 (N_4537,N_189,N_1880);
or U4538 (N_4538,N_559,N_2829);
nand U4539 (N_4539,N_624,N_2652);
xnor U4540 (N_4540,N_1013,N_2215);
nor U4541 (N_4541,N_734,N_2848);
and U4542 (N_4542,N_605,N_756);
or U4543 (N_4543,N_2096,N_3120);
and U4544 (N_4544,N_1164,N_255);
nand U4545 (N_4545,N_776,N_495);
nand U4546 (N_4546,N_206,N_880);
nand U4547 (N_4547,N_536,N_633);
xor U4548 (N_4548,N_1603,N_138);
nor U4549 (N_4549,N_976,N_2145);
or U4550 (N_4550,N_300,N_1754);
nor U4551 (N_4551,N_2187,N_1435);
or U4552 (N_4552,N_1907,N_1941);
nand U4553 (N_4553,N_2832,N_204);
and U4554 (N_4554,N_242,N_921);
and U4555 (N_4555,N_560,N_280);
or U4556 (N_4556,N_2147,N_2497);
or U4557 (N_4557,N_1874,N_1952);
nand U4558 (N_4558,N_1490,N_452);
and U4559 (N_4559,N_2158,N_1362);
nor U4560 (N_4560,N_1123,N_2612);
and U4561 (N_4561,N_1469,N_3112);
nand U4562 (N_4562,N_1177,N_438);
nand U4563 (N_4563,N_1488,N_2326);
or U4564 (N_4564,N_1386,N_1028);
xor U4565 (N_4565,N_3104,N_2953);
and U4566 (N_4566,N_1020,N_2745);
xnor U4567 (N_4567,N_352,N_1319);
or U4568 (N_4568,N_1082,N_1380);
or U4569 (N_4569,N_11,N_266);
xnor U4570 (N_4570,N_1265,N_213);
and U4571 (N_4571,N_2504,N_790);
or U4572 (N_4572,N_956,N_2815);
or U4573 (N_4573,N_2338,N_827);
and U4574 (N_4574,N_3093,N_3049);
nand U4575 (N_4575,N_2414,N_1162);
nor U4576 (N_4576,N_2103,N_1597);
nand U4577 (N_4577,N_234,N_516);
or U4578 (N_4578,N_741,N_2115);
nor U4579 (N_4579,N_1184,N_775);
nor U4580 (N_4580,N_2184,N_2444);
nor U4581 (N_4581,N_744,N_143);
xnor U4582 (N_4582,N_803,N_350);
or U4583 (N_4583,N_864,N_1684);
nand U4584 (N_4584,N_596,N_2290);
nor U4585 (N_4585,N_1621,N_434);
nand U4586 (N_4586,N_1942,N_137);
xnor U4587 (N_4587,N_1745,N_1145);
nor U4588 (N_4588,N_1549,N_1125);
and U4589 (N_4589,N_504,N_713);
or U4590 (N_4590,N_3058,N_330);
or U4591 (N_4591,N_1785,N_1817);
and U4592 (N_4592,N_2041,N_1657);
or U4593 (N_4593,N_2294,N_430);
or U4594 (N_4594,N_175,N_1873);
nand U4595 (N_4595,N_1150,N_1593);
or U4596 (N_4596,N_1661,N_798);
xnor U4597 (N_4597,N_2781,N_399);
nand U4598 (N_4598,N_2536,N_131);
nor U4599 (N_4599,N_2291,N_2951);
xnor U4600 (N_4600,N_1777,N_177);
nor U4601 (N_4601,N_1730,N_932);
and U4602 (N_4602,N_81,N_2172);
or U4603 (N_4603,N_2378,N_417);
or U4604 (N_4604,N_3096,N_2193);
nor U4605 (N_4605,N_1289,N_2983);
xor U4606 (N_4606,N_17,N_571);
nor U4607 (N_4607,N_491,N_1052);
and U4608 (N_4608,N_2969,N_684);
or U4609 (N_4609,N_2043,N_2363);
or U4610 (N_4610,N_476,N_82);
nor U4611 (N_4611,N_358,N_1325);
or U4612 (N_4612,N_151,N_1176);
nand U4613 (N_4613,N_2074,N_174);
and U4614 (N_4614,N_1889,N_231);
or U4615 (N_4615,N_1951,N_1328);
xor U4616 (N_4616,N_661,N_215);
nor U4617 (N_4617,N_8,N_1092);
or U4618 (N_4618,N_518,N_1516);
nand U4619 (N_4619,N_353,N_2952);
nor U4620 (N_4620,N_1146,N_1858);
nand U4621 (N_4621,N_2351,N_2975);
nand U4622 (N_4622,N_420,N_750);
xor U4623 (N_4623,N_2242,N_2394);
and U4624 (N_4624,N_478,N_2666);
xor U4625 (N_4625,N_2068,N_1165);
or U4626 (N_4626,N_1514,N_325);
nand U4627 (N_4627,N_123,N_2693);
and U4628 (N_4628,N_2108,N_2006);
xor U4629 (N_4629,N_3122,N_2281);
nand U4630 (N_4630,N_32,N_740);
nor U4631 (N_4631,N_3050,N_2001);
and U4632 (N_4632,N_1515,N_51);
and U4633 (N_4633,N_2430,N_145);
xor U4634 (N_4634,N_1348,N_2309);
and U4635 (N_4635,N_1008,N_1605);
and U4636 (N_4636,N_178,N_507);
nand U4637 (N_4637,N_1744,N_1498);
or U4638 (N_4638,N_2015,N_2468);
nor U4639 (N_4639,N_2518,N_2625);
and U4640 (N_4640,N_737,N_656);
or U4641 (N_4641,N_297,N_711);
nor U4642 (N_4642,N_2849,N_581);
nand U4643 (N_4643,N_601,N_570);
nor U4644 (N_4644,N_3023,N_2971);
and U4645 (N_4645,N_1831,N_1119);
xor U4646 (N_4646,N_2377,N_2267);
and U4647 (N_4647,N_539,N_2081);
or U4648 (N_4648,N_341,N_2757);
or U4649 (N_4649,N_1500,N_227);
nor U4650 (N_4650,N_564,N_2027);
nand U4651 (N_4651,N_1207,N_338);
or U4652 (N_4652,N_2284,N_1453);
or U4653 (N_4653,N_2054,N_181);
and U4654 (N_4654,N_2998,N_1644);
nand U4655 (N_4655,N_1384,N_2467);
xor U4656 (N_4656,N_2413,N_722);
and U4657 (N_4657,N_1259,N_1642);
and U4658 (N_4658,N_2411,N_441);
or U4659 (N_4659,N_1737,N_468);
nor U4660 (N_4660,N_2558,N_1178);
nor U4661 (N_4661,N_1845,N_580);
or U4662 (N_4662,N_2885,N_761);
nand U4663 (N_4663,N_1260,N_2916);
nor U4664 (N_4664,N_319,N_39);
nor U4665 (N_4665,N_1623,N_222);
xnor U4666 (N_4666,N_1965,N_2731);
nor U4667 (N_4667,N_2711,N_1304);
nor U4668 (N_4668,N_787,N_959);
and U4669 (N_4669,N_1557,N_2790);
nand U4670 (N_4670,N_2782,N_1155);
and U4671 (N_4671,N_2424,N_1117);
and U4672 (N_4672,N_913,N_852);
nor U4673 (N_4673,N_2845,N_364);
nand U4674 (N_4674,N_25,N_1163);
nand U4675 (N_4675,N_1147,N_1151);
nor U4676 (N_4676,N_2992,N_1291);
and U4677 (N_4677,N_244,N_141);
xnor U4678 (N_4678,N_904,N_2140);
nor U4679 (N_4679,N_373,N_1069);
nor U4680 (N_4680,N_808,N_763);
or U4681 (N_4681,N_2234,N_1853);
nor U4682 (N_4682,N_1890,N_657);
nor U4683 (N_4683,N_2877,N_2216);
or U4684 (N_4684,N_542,N_509);
nor U4685 (N_4685,N_294,N_1110);
and U4686 (N_4686,N_2495,N_1124);
xor U4687 (N_4687,N_2576,N_903);
nand U4688 (N_4688,N_1428,N_676);
xnor U4689 (N_4689,N_2069,N_2068);
or U4690 (N_4690,N_1761,N_3060);
or U4691 (N_4691,N_2137,N_1561);
xor U4692 (N_4692,N_1354,N_421);
or U4693 (N_4693,N_414,N_1404);
nor U4694 (N_4694,N_591,N_353);
and U4695 (N_4695,N_2628,N_707);
nand U4696 (N_4696,N_352,N_1856);
nand U4697 (N_4697,N_2152,N_829);
xnor U4698 (N_4698,N_1887,N_1396);
nand U4699 (N_4699,N_246,N_976);
nor U4700 (N_4700,N_1227,N_1605);
xnor U4701 (N_4701,N_767,N_938);
xor U4702 (N_4702,N_540,N_2003);
nor U4703 (N_4703,N_2554,N_2191);
nand U4704 (N_4704,N_1918,N_2763);
nand U4705 (N_4705,N_760,N_747);
xnor U4706 (N_4706,N_882,N_1858);
xnor U4707 (N_4707,N_214,N_2176);
or U4708 (N_4708,N_2438,N_2369);
or U4709 (N_4709,N_1637,N_845);
or U4710 (N_4710,N_1123,N_366);
nand U4711 (N_4711,N_2034,N_349);
or U4712 (N_4712,N_1571,N_1122);
or U4713 (N_4713,N_1419,N_792);
nand U4714 (N_4714,N_1728,N_2606);
xnor U4715 (N_4715,N_1818,N_1875);
and U4716 (N_4716,N_1384,N_292);
and U4717 (N_4717,N_1536,N_2613);
and U4718 (N_4718,N_1068,N_2249);
and U4719 (N_4719,N_500,N_114);
and U4720 (N_4720,N_1191,N_2792);
nand U4721 (N_4721,N_1391,N_18);
or U4722 (N_4722,N_1777,N_1853);
and U4723 (N_4723,N_1004,N_1382);
nand U4724 (N_4724,N_2725,N_1866);
nand U4725 (N_4725,N_764,N_1384);
and U4726 (N_4726,N_709,N_742);
nor U4727 (N_4727,N_975,N_17);
and U4728 (N_4728,N_687,N_463);
or U4729 (N_4729,N_499,N_2760);
xnor U4730 (N_4730,N_2609,N_769);
or U4731 (N_4731,N_2828,N_1991);
nand U4732 (N_4732,N_241,N_2321);
and U4733 (N_4733,N_2350,N_828);
nor U4734 (N_4734,N_1063,N_1228);
and U4735 (N_4735,N_193,N_474);
and U4736 (N_4736,N_1757,N_2834);
nand U4737 (N_4737,N_333,N_91);
nand U4738 (N_4738,N_597,N_918);
nand U4739 (N_4739,N_376,N_2131);
or U4740 (N_4740,N_1389,N_1814);
and U4741 (N_4741,N_2979,N_1033);
and U4742 (N_4742,N_1961,N_1207);
or U4743 (N_4743,N_1393,N_571);
xnor U4744 (N_4744,N_1706,N_298);
xnor U4745 (N_4745,N_314,N_2066);
xor U4746 (N_4746,N_2138,N_1700);
or U4747 (N_4747,N_1022,N_636);
and U4748 (N_4748,N_403,N_377);
and U4749 (N_4749,N_1212,N_832);
or U4750 (N_4750,N_1201,N_2113);
xnor U4751 (N_4751,N_2614,N_911);
nand U4752 (N_4752,N_1436,N_2997);
nor U4753 (N_4753,N_2429,N_2979);
nor U4754 (N_4754,N_1700,N_29);
or U4755 (N_4755,N_1187,N_1813);
nor U4756 (N_4756,N_1402,N_2049);
xor U4757 (N_4757,N_2637,N_2526);
nand U4758 (N_4758,N_392,N_954);
nor U4759 (N_4759,N_1814,N_2745);
nand U4760 (N_4760,N_890,N_1213);
xnor U4761 (N_4761,N_857,N_2194);
xor U4762 (N_4762,N_1938,N_218);
nor U4763 (N_4763,N_2296,N_1393);
and U4764 (N_4764,N_2346,N_2122);
or U4765 (N_4765,N_1365,N_1456);
nand U4766 (N_4766,N_2571,N_286);
xor U4767 (N_4767,N_1476,N_452);
nor U4768 (N_4768,N_2778,N_1765);
or U4769 (N_4769,N_2988,N_2869);
nor U4770 (N_4770,N_1434,N_551);
or U4771 (N_4771,N_1987,N_619);
nor U4772 (N_4772,N_926,N_1474);
nand U4773 (N_4773,N_154,N_1264);
nor U4774 (N_4774,N_2179,N_2037);
nand U4775 (N_4775,N_2186,N_888);
xor U4776 (N_4776,N_734,N_530);
nand U4777 (N_4777,N_1651,N_1452);
and U4778 (N_4778,N_2413,N_907);
or U4779 (N_4779,N_1086,N_2607);
or U4780 (N_4780,N_125,N_2263);
nand U4781 (N_4781,N_3117,N_5);
and U4782 (N_4782,N_3058,N_2345);
and U4783 (N_4783,N_796,N_813);
nor U4784 (N_4784,N_2114,N_1545);
xnor U4785 (N_4785,N_29,N_2869);
and U4786 (N_4786,N_3049,N_1739);
and U4787 (N_4787,N_2173,N_696);
xnor U4788 (N_4788,N_678,N_1148);
nand U4789 (N_4789,N_184,N_1337);
and U4790 (N_4790,N_1202,N_612);
xor U4791 (N_4791,N_1837,N_732);
and U4792 (N_4792,N_2458,N_445);
or U4793 (N_4793,N_716,N_1900);
xor U4794 (N_4794,N_937,N_2789);
xnor U4795 (N_4795,N_3075,N_984);
or U4796 (N_4796,N_426,N_1868);
and U4797 (N_4797,N_1267,N_255);
xor U4798 (N_4798,N_763,N_1337);
nor U4799 (N_4799,N_2997,N_2851);
or U4800 (N_4800,N_1864,N_3030);
or U4801 (N_4801,N_411,N_3094);
xor U4802 (N_4802,N_2412,N_1400);
nor U4803 (N_4803,N_76,N_2723);
or U4804 (N_4804,N_1648,N_2151);
and U4805 (N_4805,N_2575,N_312);
and U4806 (N_4806,N_6,N_3102);
nor U4807 (N_4807,N_17,N_798);
nor U4808 (N_4808,N_1630,N_2707);
xnor U4809 (N_4809,N_242,N_1102);
nor U4810 (N_4810,N_2082,N_837);
xnor U4811 (N_4811,N_1361,N_2077);
nor U4812 (N_4812,N_211,N_253);
nor U4813 (N_4813,N_1134,N_2988);
and U4814 (N_4814,N_954,N_2162);
nor U4815 (N_4815,N_2494,N_2053);
nor U4816 (N_4816,N_2205,N_2070);
nand U4817 (N_4817,N_3042,N_1975);
nor U4818 (N_4818,N_1124,N_1509);
or U4819 (N_4819,N_1680,N_1040);
nand U4820 (N_4820,N_1546,N_378);
or U4821 (N_4821,N_2567,N_2724);
or U4822 (N_4822,N_280,N_620);
or U4823 (N_4823,N_1689,N_2576);
nor U4824 (N_4824,N_722,N_2067);
or U4825 (N_4825,N_2231,N_3111);
nand U4826 (N_4826,N_1318,N_1787);
nand U4827 (N_4827,N_624,N_2441);
and U4828 (N_4828,N_3010,N_1150);
xnor U4829 (N_4829,N_254,N_2879);
or U4830 (N_4830,N_2103,N_1038);
xnor U4831 (N_4831,N_1919,N_422);
nand U4832 (N_4832,N_2531,N_2634);
xnor U4833 (N_4833,N_2616,N_1887);
nor U4834 (N_4834,N_72,N_3013);
nor U4835 (N_4835,N_2518,N_1733);
nand U4836 (N_4836,N_1861,N_953);
and U4837 (N_4837,N_1694,N_840);
nand U4838 (N_4838,N_779,N_1604);
nor U4839 (N_4839,N_1196,N_2462);
or U4840 (N_4840,N_899,N_1362);
nand U4841 (N_4841,N_2887,N_2655);
or U4842 (N_4842,N_2123,N_726);
and U4843 (N_4843,N_1924,N_1825);
nand U4844 (N_4844,N_2862,N_1230);
nand U4845 (N_4845,N_21,N_1363);
and U4846 (N_4846,N_2766,N_1839);
or U4847 (N_4847,N_2854,N_57);
or U4848 (N_4848,N_701,N_2135);
and U4849 (N_4849,N_2650,N_194);
and U4850 (N_4850,N_163,N_2480);
nor U4851 (N_4851,N_2584,N_1391);
and U4852 (N_4852,N_2507,N_2470);
nand U4853 (N_4853,N_1209,N_1328);
nor U4854 (N_4854,N_2262,N_2644);
nand U4855 (N_4855,N_1604,N_2);
xor U4856 (N_4856,N_2492,N_961);
nand U4857 (N_4857,N_1294,N_687);
xor U4858 (N_4858,N_2707,N_1923);
and U4859 (N_4859,N_536,N_3103);
or U4860 (N_4860,N_1535,N_2724);
nor U4861 (N_4861,N_1510,N_3117);
or U4862 (N_4862,N_970,N_2410);
nand U4863 (N_4863,N_799,N_896);
nor U4864 (N_4864,N_2601,N_9);
nor U4865 (N_4865,N_221,N_1641);
xor U4866 (N_4866,N_1874,N_1094);
nor U4867 (N_4867,N_1678,N_3081);
nor U4868 (N_4868,N_574,N_1274);
xnor U4869 (N_4869,N_2229,N_745);
xnor U4870 (N_4870,N_2520,N_613);
nand U4871 (N_4871,N_1188,N_2393);
nor U4872 (N_4872,N_2138,N_2093);
and U4873 (N_4873,N_1840,N_1381);
or U4874 (N_4874,N_1057,N_1149);
nor U4875 (N_4875,N_2472,N_1414);
and U4876 (N_4876,N_1635,N_1006);
or U4877 (N_4877,N_3114,N_2386);
or U4878 (N_4878,N_981,N_2696);
or U4879 (N_4879,N_827,N_28);
xor U4880 (N_4880,N_1136,N_978);
or U4881 (N_4881,N_1758,N_2720);
and U4882 (N_4882,N_1208,N_418);
and U4883 (N_4883,N_1826,N_2628);
xnor U4884 (N_4884,N_1601,N_1999);
nand U4885 (N_4885,N_1976,N_458);
nor U4886 (N_4886,N_918,N_429);
or U4887 (N_4887,N_1212,N_2846);
and U4888 (N_4888,N_2384,N_69);
xnor U4889 (N_4889,N_2975,N_2340);
nor U4890 (N_4890,N_1238,N_1370);
or U4891 (N_4891,N_2197,N_943);
and U4892 (N_4892,N_2595,N_1501);
or U4893 (N_4893,N_2116,N_548);
xor U4894 (N_4894,N_2271,N_1554);
xor U4895 (N_4895,N_2295,N_1582);
nand U4896 (N_4896,N_1916,N_2834);
nand U4897 (N_4897,N_2435,N_814);
and U4898 (N_4898,N_1387,N_802);
xnor U4899 (N_4899,N_2857,N_532);
nand U4900 (N_4900,N_1713,N_2446);
xor U4901 (N_4901,N_1558,N_2387);
xor U4902 (N_4902,N_1382,N_606);
or U4903 (N_4903,N_418,N_1411);
and U4904 (N_4904,N_1052,N_2115);
and U4905 (N_4905,N_650,N_522);
xor U4906 (N_4906,N_2373,N_787);
nor U4907 (N_4907,N_214,N_1069);
nand U4908 (N_4908,N_717,N_974);
or U4909 (N_4909,N_2241,N_536);
nand U4910 (N_4910,N_1386,N_2265);
nor U4911 (N_4911,N_1573,N_1251);
and U4912 (N_4912,N_2019,N_2803);
and U4913 (N_4913,N_1357,N_1553);
and U4914 (N_4914,N_708,N_709);
or U4915 (N_4915,N_720,N_1068);
and U4916 (N_4916,N_2117,N_1755);
nand U4917 (N_4917,N_2732,N_2310);
nor U4918 (N_4918,N_2713,N_1997);
or U4919 (N_4919,N_2306,N_2512);
xor U4920 (N_4920,N_1617,N_162);
and U4921 (N_4921,N_2811,N_1928);
or U4922 (N_4922,N_1518,N_1505);
nor U4923 (N_4923,N_2375,N_2679);
nand U4924 (N_4924,N_2112,N_1519);
nor U4925 (N_4925,N_1497,N_2765);
xnor U4926 (N_4926,N_482,N_3054);
or U4927 (N_4927,N_2623,N_384);
and U4928 (N_4928,N_2605,N_2248);
nand U4929 (N_4929,N_891,N_975);
and U4930 (N_4930,N_768,N_486);
nand U4931 (N_4931,N_2263,N_1560);
and U4932 (N_4932,N_459,N_352);
nor U4933 (N_4933,N_447,N_1536);
nand U4934 (N_4934,N_1687,N_2403);
nor U4935 (N_4935,N_2862,N_1711);
xnor U4936 (N_4936,N_714,N_1810);
nand U4937 (N_4937,N_3108,N_2625);
or U4938 (N_4938,N_1279,N_587);
nand U4939 (N_4939,N_2558,N_2223);
xnor U4940 (N_4940,N_247,N_2572);
and U4941 (N_4941,N_115,N_2807);
nor U4942 (N_4942,N_19,N_1728);
xor U4943 (N_4943,N_2088,N_1830);
or U4944 (N_4944,N_1535,N_2047);
nand U4945 (N_4945,N_400,N_1100);
and U4946 (N_4946,N_1704,N_1709);
or U4947 (N_4947,N_2413,N_1192);
nand U4948 (N_4948,N_2368,N_182);
nand U4949 (N_4949,N_1233,N_2921);
or U4950 (N_4950,N_742,N_434);
and U4951 (N_4951,N_1869,N_713);
nand U4952 (N_4952,N_798,N_2611);
and U4953 (N_4953,N_2276,N_1328);
xor U4954 (N_4954,N_2535,N_2092);
or U4955 (N_4955,N_267,N_508);
nor U4956 (N_4956,N_230,N_2353);
nand U4957 (N_4957,N_1875,N_2760);
xor U4958 (N_4958,N_1386,N_2497);
xnor U4959 (N_4959,N_1719,N_512);
nand U4960 (N_4960,N_1630,N_2402);
xor U4961 (N_4961,N_426,N_619);
or U4962 (N_4962,N_946,N_2121);
nand U4963 (N_4963,N_270,N_1626);
nor U4964 (N_4964,N_177,N_1677);
xor U4965 (N_4965,N_2861,N_1914);
nand U4966 (N_4966,N_314,N_2470);
xor U4967 (N_4967,N_1582,N_1670);
or U4968 (N_4968,N_956,N_1987);
or U4969 (N_4969,N_1199,N_695);
xnor U4970 (N_4970,N_1112,N_45);
nor U4971 (N_4971,N_1475,N_2440);
or U4972 (N_4972,N_2481,N_267);
xnor U4973 (N_4973,N_2622,N_388);
nand U4974 (N_4974,N_1213,N_1927);
or U4975 (N_4975,N_995,N_495);
and U4976 (N_4976,N_3073,N_1979);
or U4977 (N_4977,N_2745,N_659);
and U4978 (N_4978,N_1002,N_1296);
nor U4979 (N_4979,N_862,N_23);
or U4980 (N_4980,N_2333,N_2380);
and U4981 (N_4981,N_264,N_2389);
and U4982 (N_4982,N_194,N_2204);
and U4983 (N_4983,N_469,N_2101);
and U4984 (N_4984,N_1361,N_1601);
nor U4985 (N_4985,N_2684,N_1887);
xor U4986 (N_4986,N_2689,N_712);
and U4987 (N_4987,N_2180,N_673);
or U4988 (N_4988,N_2062,N_757);
nand U4989 (N_4989,N_234,N_2355);
xor U4990 (N_4990,N_824,N_2970);
and U4991 (N_4991,N_2063,N_1981);
xor U4992 (N_4992,N_2483,N_1749);
nand U4993 (N_4993,N_792,N_1846);
nor U4994 (N_4994,N_2544,N_2276);
nor U4995 (N_4995,N_594,N_2522);
and U4996 (N_4996,N_1415,N_16);
nand U4997 (N_4997,N_722,N_713);
nor U4998 (N_4998,N_2039,N_1012);
xnor U4999 (N_4999,N_1440,N_465);
nor U5000 (N_5000,N_2490,N_2714);
and U5001 (N_5001,N_396,N_1749);
and U5002 (N_5002,N_646,N_741);
and U5003 (N_5003,N_1106,N_2263);
xor U5004 (N_5004,N_2188,N_2375);
and U5005 (N_5005,N_960,N_1227);
xor U5006 (N_5006,N_2637,N_925);
nand U5007 (N_5007,N_1573,N_691);
nand U5008 (N_5008,N_2100,N_1095);
or U5009 (N_5009,N_2874,N_1832);
xor U5010 (N_5010,N_1523,N_565);
and U5011 (N_5011,N_1264,N_2876);
and U5012 (N_5012,N_2117,N_1337);
xnor U5013 (N_5013,N_15,N_1707);
or U5014 (N_5014,N_1900,N_2765);
nor U5015 (N_5015,N_3050,N_798);
xor U5016 (N_5016,N_451,N_874);
xor U5017 (N_5017,N_942,N_2418);
nor U5018 (N_5018,N_2005,N_2818);
or U5019 (N_5019,N_2120,N_893);
and U5020 (N_5020,N_2414,N_2146);
nor U5021 (N_5021,N_2435,N_128);
and U5022 (N_5022,N_2274,N_1624);
nand U5023 (N_5023,N_35,N_861);
xor U5024 (N_5024,N_457,N_2846);
nand U5025 (N_5025,N_2591,N_120);
xor U5026 (N_5026,N_2895,N_2014);
or U5027 (N_5027,N_311,N_469);
and U5028 (N_5028,N_542,N_1034);
and U5029 (N_5029,N_1643,N_2176);
or U5030 (N_5030,N_2602,N_2790);
and U5031 (N_5031,N_2097,N_622);
nand U5032 (N_5032,N_394,N_3052);
xnor U5033 (N_5033,N_1949,N_1242);
nor U5034 (N_5034,N_914,N_1396);
nand U5035 (N_5035,N_463,N_490);
and U5036 (N_5036,N_124,N_2663);
or U5037 (N_5037,N_2829,N_2828);
nor U5038 (N_5038,N_2585,N_47);
nand U5039 (N_5039,N_1270,N_1782);
and U5040 (N_5040,N_3072,N_1150);
nand U5041 (N_5041,N_142,N_959);
or U5042 (N_5042,N_1395,N_396);
nor U5043 (N_5043,N_1491,N_1147);
nor U5044 (N_5044,N_1570,N_1697);
nand U5045 (N_5045,N_1784,N_1285);
nor U5046 (N_5046,N_1075,N_2808);
or U5047 (N_5047,N_2691,N_1348);
and U5048 (N_5048,N_772,N_2822);
and U5049 (N_5049,N_2400,N_2616);
nand U5050 (N_5050,N_1221,N_1430);
xnor U5051 (N_5051,N_2254,N_29);
nor U5052 (N_5052,N_115,N_1523);
xnor U5053 (N_5053,N_1232,N_973);
or U5054 (N_5054,N_1232,N_2941);
or U5055 (N_5055,N_1877,N_875);
nor U5056 (N_5056,N_1906,N_2794);
and U5057 (N_5057,N_199,N_1096);
or U5058 (N_5058,N_2456,N_963);
or U5059 (N_5059,N_703,N_2261);
or U5060 (N_5060,N_515,N_1471);
nor U5061 (N_5061,N_661,N_554);
nand U5062 (N_5062,N_1679,N_2102);
nand U5063 (N_5063,N_3026,N_1974);
or U5064 (N_5064,N_633,N_2964);
nor U5065 (N_5065,N_3010,N_2864);
or U5066 (N_5066,N_1739,N_2651);
nor U5067 (N_5067,N_804,N_2090);
nor U5068 (N_5068,N_2990,N_1499);
nand U5069 (N_5069,N_842,N_85);
or U5070 (N_5070,N_1289,N_2301);
nor U5071 (N_5071,N_864,N_1596);
nor U5072 (N_5072,N_482,N_2614);
nand U5073 (N_5073,N_1387,N_841);
nor U5074 (N_5074,N_0,N_1121);
nor U5075 (N_5075,N_2663,N_2481);
xor U5076 (N_5076,N_2670,N_323);
and U5077 (N_5077,N_2504,N_1950);
nand U5078 (N_5078,N_789,N_2749);
and U5079 (N_5079,N_2278,N_2075);
or U5080 (N_5080,N_315,N_649);
nor U5081 (N_5081,N_603,N_1944);
nor U5082 (N_5082,N_2409,N_2935);
and U5083 (N_5083,N_2565,N_1669);
nand U5084 (N_5084,N_1440,N_1594);
nor U5085 (N_5085,N_30,N_586);
nor U5086 (N_5086,N_2274,N_732);
or U5087 (N_5087,N_3092,N_2638);
or U5088 (N_5088,N_1358,N_2405);
and U5089 (N_5089,N_889,N_1610);
and U5090 (N_5090,N_2032,N_482);
nor U5091 (N_5091,N_3118,N_2711);
nand U5092 (N_5092,N_2877,N_3009);
nand U5093 (N_5093,N_739,N_1953);
xor U5094 (N_5094,N_2922,N_2615);
or U5095 (N_5095,N_545,N_992);
or U5096 (N_5096,N_2673,N_1073);
or U5097 (N_5097,N_3112,N_1163);
nand U5098 (N_5098,N_2304,N_1990);
nand U5099 (N_5099,N_1235,N_437);
nand U5100 (N_5100,N_1121,N_2188);
or U5101 (N_5101,N_862,N_1954);
nor U5102 (N_5102,N_1247,N_1790);
and U5103 (N_5103,N_2407,N_429);
or U5104 (N_5104,N_2448,N_2508);
nand U5105 (N_5105,N_2804,N_1808);
nor U5106 (N_5106,N_1453,N_2115);
nor U5107 (N_5107,N_2990,N_1832);
xnor U5108 (N_5108,N_2611,N_135);
and U5109 (N_5109,N_2136,N_1051);
nand U5110 (N_5110,N_1982,N_1559);
xnor U5111 (N_5111,N_232,N_2235);
nand U5112 (N_5112,N_1842,N_2155);
xnor U5113 (N_5113,N_417,N_1818);
xor U5114 (N_5114,N_539,N_1186);
and U5115 (N_5115,N_2930,N_159);
xnor U5116 (N_5116,N_2314,N_325);
nor U5117 (N_5117,N_1489,N_1538);
nand U5118 (N_5118,N_1606,N_2058);
and U5119 (N_5119,N_1146,N_1098);
xor U5120 (N_5120,N_2680,N_1396);
nor U5121 (N_5121,N_782,N_1056);
and U5122 (N_5122,N_1226,N_683);
and U5123 (N_5123,N_2910,N_2144);
and U5124 (N_5124,N_706,N_2853);
xnor U5125 (N_5125,N_551,N_1220);
or U5126 (N_5126,N_1835,N_319);
and U5127 (N_5127,N_2450,N_1206);
xor U5128 (N_5128,N_1625,N_960);
xor U5129 (N_5129,N_2160,N_101);
nor U5130 (N_5130,N_2817,N_2545);
and U5131 (N_5131,N_3009,N_357);
nor U5132 (N_5132,N_1703,N_595);
and U5133 (N_5133,N_991,N_2397);
or U5134 (N_5134,N_236,N_1378);
nor U5135 (N_5135,N_1818,N_297);
and U5136 (N_5136,N_564,N_1084);
and U5137 (N_5137,N_1110,N_2280);
nand U5138 (N_5138,N_1011,N_163);
nor U5139 (N_5139,N_2342,N_970);
xor U5140 (N_5140,N_967,N_2905);
xnor U5141 (N_5141,N_2512,N_1995);
nand U5142 (N_5142,N_1386,N_1941);
and U5143 (N_5143,N_2767,N_2060);
nor U5144 (N_5144,N_2073,N_680);
nand U5145 (N_5145,N_2827,N_1020);
nand U5146 (N_5146,N_1237,N_1811);
or U5147 (N_5147,N_2803,N_512);
or U5148 (N_5148,N_825,N_978);
xor U5149 (N_5149,N_1539,N_1633);
nand U5150 (N_5150,N_3003,N_1342);
nand U5151 (N_5151,N_621,N_1595);
nor U5152 (N_5152,N_1483,N_636);
or U5153 (N_5153,N_1656,N_2625);
xnor U5154 (N_5154,N_3067,N_1192);
xor U5155 (N_5155,N_2583,N_1421);
nand U5156 (N_5156,N_228,N_898);
and U5157 (N_5157,N_2486,N_2367);
xor U5158 (N_5158,N_2201,N_2696);
nand U5159 (N_5159,N_2170,N_2714);
xnor U5160 (N_5160,N_1064,N_288);
nor U5161 (N_5161,N_2688,N_1543);
or U5162 (N_5162,N_406,N_1241);
nand U5163 (N_5163,N_2356,N_2253);
and U5164 (N_5164,N_1844,N_973);
and U5165 (N_5165,N_767,N_327);
nor U5166 (N_5166,N_2636,N_2095);
nand U5167 (N_5167,N_1851,N_444);
nand U5168 (N_5168,N_879,N_1989);
nand U5169 (N_5169,N_1140,N_264);
nor U5170 (N_5170,N_66,N_2450);
or U5171 (N_5171,N_2763,N_2952);
and U5172 (N_5172,N_1798,N_2407);
xor U5173 (N_5173,N_2568,N_579);
xor U5174 (N_5174,N_1255,N_3007);
or U5175 (N_5175,N_3056,N_953);
nand U5176 (N_5176,N_428,N_994);
xor U5177 (N_5177,N_1166,N_38);
nand U5178 (N_5178,N_19,N_2675);
or U5179 (N_5179,N_2812,N_2077);
nand U5180 (N_5180,N_3034,N_2101);
xor U5181 (N_5181,N_332,N_1258);
and U5182 (N_5182,N_2658,N_2525);
nor U5183 (N_5183,N_2487,N_800);
nor U5184 (N_5184,N_2994,N_208);
nor U5185 (N_5185,N_2313,N_712);
and U5186 (N_5186,N_1378,N_2524);
and U5187 (N_5187,N_2623,N_2017);
and U5188 (N_5188,N_1979,N_924);
xnor U5189 (N_5189,N_2261,N_2369);
or U5190 (N_5190,N_839,N_1383);
xor U5191 (N_5191,N_582,N_1155);
nand U5192 (N_5192,N_1853,N_1647);
nor U5193 (N_5193,N_577,N_2409);
xnor U5194 (N_5194,N_954,N_739);
nor U5195 (N_5195,N_839,N_2573);
and U5196 (N_5196,N_19,N_1803);
or U5197 (N_5197,N_1879,N_2311);
xnor U5198 (N_5198,N_1614,N_523);
nand U5199 (N_5199,N_1073,N_2342);
or U5200 (N_5200,N_135,N_2461);
xor U5201 (N_5201,N_652,N_2967);
nand U5202 (N_5202,N_1755,N_1552);
and U5203 (N_5203,N_456,N_338);
nor U5204 (N_5204,N_2537,N_360);
or U5205 (N_5205,N_471,N_1312);
or U5206 (N_5206,N_2615,N_1932);
or U5207 (N_5207,N_208,N_2976);
and U5208 (N_5208,N_426,N_82);
nor U5209 (N_5209,N_1276,N_3105);
nor U5210 (N_5210,N_2201,N_2761);
nor U5211 (N_5211,N_635,N_3035);
nand U5212 (N_5212,N_2468,N_35);
and U5213 (N_5213,N_866,N_2698);
nor U5214 (N_5214,N_2249,N_2442);
and U5215 (N_5215,N_956,N_2580);
xnor U5216 (N_5216,N_83,N_843);
xnor U5217 (N_5217,N_246,N_1499);
nand U5218 (N_5218,N_138,N_1668);
or U5219 (N_5219,N_614,N_2149);
or U5220 (N_5220,N_1224,N_2245);
or U5221 (N_5221,N_2833,N_748);
xnor U5222 (N_5222,N_1334,N_408);
xnor U5223 (N_5223,N_1811,N_2212);
and U5224 (N_5224,N_1514,N_302);
nor U5225 (N_5225,N_770,N_3037);
nand U5226 (N_5226,N_2555,N_1097);
nor U5227 (N_5227,N_2801,N_2733);
nor U5228 (N_5228,N_2206,N_1814);
nand U5229 (N_5229,N_578,N_3037);
nor U5230 (N_5230,N_741,N_43);
xnor U5231 (N_5231,N_2699,N_2610);
or U5232 (N_5232,N_1220,N_1939);
nor U5233 (N_5233,N_2045,N_872);
nor U5234 (N_5234,N_2521,N_1330);
nor U5235 (N_5235,N_2622,N_1573);
nor U5236 (N_5236,N_606,N_1916);
nand U5237 (N_5237,N_779,N_2173);
and U5238 (N_5238,N_535,N_371);
or U5239 (N_5239,N_3039,N_1687);
or U5240 (N_5240,N_2040,N_1004);
nand U5241 (N_5241,N_511,N_1969);
and U5242 (N_5242,N_1647,N_561);
nand U5243 (N_5243,N_2460,N_2089);
or U5244 (N_5244,N_1702,N_916);
nor U5245 (N_5245,N_500,N_674);
nand U5246 (N_5246,N_2649,N_2488);
nand U5247 (N_5247,N_1765,N_585);
or U5248 (N_5248,N_1546,N_3025);
xnor U5249 (N_5249,N_1097,N_1509);
or U5250 (N_5250,N_2982,N_1661);
nand U5251 (N_5251,N_941,N_619);
xnor U5252 (N_5252,N_2412,N_2341);
or U5253 (N_5253,N_2279,N_2058);
nor U5254 (N_5254,N_1322,N_160);
or U5255 (N_5255,N_2372,N_161);
xnor U5256 (N_5256,N_1486,N_2244);
and U5257 (N_5257,N_1396,N_1906);
nor U5258 (N_5258,N_2190,N_2146);
and U5259 (N_5259,N_737,N_658);
xnor U5260 (N_5260,N_1681,N_1033);
xor U5261 (N_5261,N_398,N_2617);
and U5262 (N_5262,N_2561,N_237);
nor U5263 (N_5263,N_1764,N_1062);
or U5264 (N_5264,N_1966,N_12);
nor U5265 (N_5265,N_2654,N_149);
xnor U5266 (N_5266,N_1730,N_2710);
or U5267 (N_5267,N_1226,N_2647);
nand U5268 (N_5268,N_1868,N_1644);
and U5269 (N_5269,N_2989,N_527);
and U5270 (N_5270,N_2784,N_190);
nor U5271 (N_5271,N_713,N_54);
nor U5272 (N_5272,N_551,N_969);
nor U5273 (N_5273,N_1893,N_1629);
or U5274 (N_5274,N_2623,N_2966);
or U5275 (N_5275,N_108,N_1035);
xor U5276 (N_5276,N_156,N_2029);
and U5277 (N_5277,N_888,N_2566);
and U5278 (N_5278,N_3111,N_2701);
nor U5279 (N_5279,N_2768,N_302);
and U5280 (N_5280,N_285,N_1140);
nand U5281 (N_5281,N_1918,N_2556);
xor U5282 (N_5282,N_1037,N_572);
nand U5283 (N_5283,N_332,N_1799);
or U5284 (N_5284,N_2213,N_2442);
nand U5285 (N_5285,N_1609,N_3001);
nor U5286 (N_5286,N_307,N_2945);
nand U5287 (N_5287,N_2241,N_769);
xor U5288 (N_5288,N_345,N_2942);
and U5289 (N_5289,N_1623,N_1477);
or U5290 (N_5290,N_2844,N_2972);
xnor U5291 (N_5291,N_1661,N_1512);
nand U5292 (N_5292,N_1634,N_2326);
or U5293 (N_5293,N_1213,N_781);
and U5294 (N_5294,N_2660,N_2480);
and U5295 (N_5295,N_2265,N_2931);
nand U5296 (N_5296,N_538,N_3059);
or U5297 (N_5297,N_779,N_687);
or U5298 (N_5298,N_1883,N_2817);
nor U5299 (N_5299,N_2906,N_849);
nand U5300 (N_5300,N_2086,N_2620);
xor U5301 (N_5301,N_1000,N_2714);
nand U5302 (N_5302,N_277,N_624);
xor U5303 (N_5303,N_2315,N_2839);
or U5304 (N_5304,N_577,N_2118);
xor U5305 (N_5305,N_1005,N_3045);
nor U5306 (N_5306,N_36,N_2851);
xnor U5307 (N_5307,N_1626,N_151);
or U5308 (N_5308,N_249,N_1220);
or U5309 (N_5309,N_1812,N_2493);
xor U5310 (N_5310,N_713,N_352);
and U5311 (N_5311,N_234,N_2562);
xnor U5312 (N_5312,N_2614,N_382);
nand U5313 (N_5313,N_2430,N_2616);
xor U5314 (N_5314,N_2882,N_1966);
nor U5315 (N_5315,N_1046,N_583);
xor U5316 (N_5316,N_1839,N_3087);
or U5317 (N_5317,N_1567,N_2531);
nor U5318 (N_5318,N_699,N_533);
xnor U5319 (N_5319,N_370,N_1742);
or U5320 (N_5320,N_1117,N_3085);
xor U5321 (N_5321,N_1598,N_1075);
or U5322 (N_5322,N_2856,N_2922);
nor U5323 (N_5323,N_1375,N_1884);
and U5324 (N_5324,N_1667,N_1182);
or U5325 (N_5325,N_456,N_2596);
nor U5326 (N_5326,N_505,N_1225);
and U5327 (N_5327,N_838,N_1109);
nand U5328 (N_5328,N_1688,N_3104);
nor U5329 (N_5329,N_893,N_1518);
nor U5330 (N_5330,N_1672,N_808);
and U5331 (N_5331,N_3017,N_1204);
xnor U5332 (N_5332,N_2159,N_1973);
xor U5333 (N_5333,N_141,N_2295);
and U5334 (N_5334,N_1386,N_2145);
nor U5335 (N_5335,N_300,N_1967);
xnor U5336 (N_5336,N_1821,N_1520);
nor U5337 (N_5337,N_1258,N_1531);
and U5338 (N_5338,N_1768,N_679);
nand U5339 (N_5339,N_712,N_1317);
or U5340 (N_5340,N_1583,N_1833);
or U5341 (N_5341,N_2637,N_3045);
xor U5342 (N_5342,N_1831,N_2287);
nand U5343 (N_5343,N_1180,N_1311);
or U5344 (N_5344,N_2643,N_614);
nand U5345 (N_5345,N_2774,N_2761);
xor U5346 (N_5346,N_884,N_2163);
xor U5347 (N_5347,N_2574,N_2017);
and U5348 (N_5348,N_546,N_1500);
or U5349 (N_5349,N_1295,N_1484);
nand U5350 (N_5350,N_866,N_1926);
nor U5351 (N_5351,N_328,N_57);
nand U5352 (N_5352,N_133,N_2259);
nand U5353 (N_5353,N_362,N_686);
nor U5354 (N_5354,N_1941,N_2449);
and U5355 (N_5355,N_1714,N_2841);
or U5356 (N_5356,N_2315,N_847);
nor U5357 (N_5357,N_2368,N_2301);
nor U5358 (N_5358,N_1367,N_1180);
or U5359 (N_5359,N_1947,N_878);
and U5360 (N_5360,N_2994,N_2343);
and U5361 (N_5361,N_2959,N_2336);
and U5362 (N_5362,N_2025,N_1731);
and U5363 (N_5363,N_2811,N_3000);
and U5364 (N_5364,N_1026,N_1778);
or U5365 (N_5365,N_226,N_2606);
nor U5366 (N_5366,N_1120,N_1987);
nor U5367 (N_5367,N_3084,N_1389);
nand U5368 (N_5368,N_671,N_1848);
or U5369 (N_5369,N_411,N_162);
nor U5370 (N_5370,N_405,N_1095);
or U5371 (N_5371,N_264,N_2118);
nor U5372 (N_5372,N_392,N_1604);
or U5373 (N_5373,N_2396,N_2380);
xor U5374 (N_5374,N_765,N_2054);
or U5375 (N_5375,N_2043,N_1504);
and U5376 (N_5376,N_465,N_328);
nand U5377 (N_5377,N_302,N_1376);
and U5378 (N_5378,N_2712,N_2081);
or U5379 (N_5379,N_705,N_2746);
or U5380 (N_5380,N_1603,N_3065);
xor U5381 (N_5381,N_2112,N_1862);
nand U5382 (N_5382,N_2431,N_2389);
xor U5383 (N_5383,N_1473,N_1232);
xor U5384 (N_5384,N_554,N_1574);
and U5385 (N_5385,N_1644,N_108);
xor U5386 (N_5386,N_2625,N_2404);
xor U5387 (N_5387,N_2793,N_2524);
nand U5388 (N_5388,N_1762,N_2358);
nand U5389 (N_5389,N_1141,N_2396);
and U5390 (N_5390,N_2365,N_1515);
and U5391 (N_5391,N_143,N_2546);
and U5392 (N_5392,N_2067,N_2286);
or U5393 (N_5393,N_867,N_752);
or U5394 (N_5394,N_2399,N_257);
nor U5395 (N_5395,N_1936,N_137);
and U5396 (N_5396,N_567,N_1579);
xnor U5397 (N_5397,N_131,N_2496);
or U5398 (N_5398,N_2169,N_426);
xnor U5399 (N_5399,N_394,N_333);
xor U5400 (N_5400,N_1385,N_97);
or U5401 (N_5401,N_1740,N_1951);
or U5402 (N_5402,N_426,N_1685);
or U5403 (N_5403,N_2062,N_2229);
and U5404 (N_5404,N_86,N_2249);
and U5405 (N_5405,N_2554,N_131);
or U5406 (N_5406,N_1318,N_1341);
nor U5407 (N_5407,N_471,N_1149);
or U5408 (N_5408,N_879,N_1104);
nor U5409 (N_5409,N_2148,N_2954);
and U5410 (N_5410,N_1922,N_2360);
nor U5411 (N_5411,N_1979,N_974);
nand U5412 (N_5412,N_1355,N_986);
nand U5413 (N_5413,N_2368,N_1113);
or U5414 (N_5414,N_2876,N_1707);
xor U5415 (N_5415,N_2516,N_1586);
or U5416 (N_5416,N_2161,N_2513);
and U5417 (N_5417,N_1736,N_373);
or U5418 (N_5418,N_1608,N_129);
nor U5419 (N_5419,N_842,N_2356);
and U5420 (N_5420,N_605,N_1993);
or U5421 (N_5421,N_2923,N_1567);
nor U5422 (N_5422,N_3003,N_1140);
or U5423 (N_5423,N_2999,N_620);
nand U5424 (N_5424,N_2969,N_874);
xnor U5425 (N_5425,N_335,N_575);
nand U5426 (N_5426,N_2890,N_2603);
and U5427 (N_5427,N_2004,N_869);
nor U5428 (N_5428,N_1980,N_838);
nand U5429 (N_5429,N_2274,N_1550);
nand U5430 (N_5430,N_1124,N_1670);
nor U5431 (N_5431,N_2847,N_407);
and U5432 (N_5432,N_1792,N_937);
and U5433 (N_5433,N_2149,N_1745);
nand U5434 (N_5434,N_1638,N_1618);
nor U5435 (N_5435,N_2006,N_2550);
and U5436 (N_5436,N_1588,N_835);
and U5437 (N_5437,N_1411,N_696);
nand U5438 (N_5438,N_1512,N_2653);
nand U5439 (N_5439,N_374,N_1612);
nor U5440 (N_5440,N_2632,N_2689);
and U5441 (N_5441,N_2447,N_2773);
nor U5442 (N_5442,N_2663,N_2434);
nor U5443 (N_5443,N_193,N_2345);
nand U5444 (N_5444,N_1609,N_1533);
nand U5445 (N_5445,N_890,N_2244);
nor U5446 (N_5446,N_1906,N_1994);
xor U5447 (N_5447,N_2040,N_796);
xnor U5448 (N_5448,N_2961,N_2154);
or U5449 (N_5449,N_420,N_987);
nor U5450 (N_5450,N_2495,N_2519);
and U5451 (N_5451,N_2797,N_1402);
or U5452 (N_5452,N_1969,N_2370);
or U5453 (N_5453,N_2283,N_1342);
and U5454 (N_5454,N_376,N_2673);
xnor U5455 (N_5455,N_2382,N_1070);
nand U5456 (N_5456,N_635,N_1465);
or U5457 (N_5457,N_2257,N_2213);
and U5458 (N_5458,N_2079,N_1920);
nor U5459 (N_5459,N_464,N_2440);
xor U5460 (N_5460,N_1616,N_325);
nand U5461 (N_5461,N_2876,N_2324);
nor U5462 (N_5462,N_466,N_2278);
xnor U5463 (N_5463,N_1792,N_1045);
nand U5464 (N_5464,N_11,N_158);
and U5465 (N_5465,N_20,N_1773);
nor U5466 (N_5466,N_763,N_1667);
xor U5467 (N_5467,N_2197,N_2875);
and U5468 (N_5468,N_2815,N_51);
nor U5469 (N_5469,N_2811,N_1950);
nand U5470 (N_5470,N_2902,N_1726);
nor U5471 (N_5471,N_2930,N_54);
nor U5472 (N_5472,N_227,N_1900);
xor U5473 (N_5473,N_426,N_698);
and U5474 (N_5474,N_2528,N_84);
and U5475 (N_5475,N_866,N_899);
or U5476 (N_5476,N_2879,N_22);
and U5477 (N_5477,N_2374,N_902);
xor U5478 (N_5478,N_1312,N_2144);
and U5479 (N_5479,N_1435,N_2340);
and U5480 (N_5480,N_2588,N_1771);
or U5481 (N_5481,N_1948,N_1162);
nor U5482 (N_5482,N_265,N_1586);
xor U5483 (N_5483,N_1434,N_2753);
xor U5484 (N_5484,N_133,N_2453);
or U5485 (N_5485,N_1325,N_3005);
xnor U5486 (N_5486,N_2165,N_822);
nor U5487 (N_5487,N_1128,N_1425);
nor U5488 (N_5488,N_2820,N_1554);
or U5489 (N_5489,N_1624,N_872);
nand U5490 (N_5490,N_1815,N_367);
nand U5491 (N_5491,N_3122,N_737);
nor U5492 (N_5492,N_868,N_162);
nand U5493 (N_5493,N_1517,N_2737);
and U5494 (N_5494,N_493,N_2711);
nand U5495 (N_5495,N_1151,N_1725);
nor U5496 (N_5496,N_1392,N_886);
or U5497 (N_5497,N_2833,N_2010);
and U5498 (N_5498,N_2610,N_227);
nand U5499 (N_5499,N_2372,N_2402);
nor U5500 (N_5500,N_1453,N_310);
xor U5501 (N_5501,N_2898,N_1796);
nor U5502 (N_5502,N_2194,N_2443);
or U5503 (N_5503,N_1362,N_1183);
xnor U5504 (N_5504,N_1976,N_294);
and U5505 (N_5505,N_1807,N_1913);
xor U5506 (N_5506,N_1105,N_1270);
or U5507 (N_5507,N_1595,N_2691);
or U5508 (N_5508,N_2497,N_15);
xor U5509 (N_5509,N_677,N_583);
xor U5510 (N_5510,N_1105,N_749);
xor U5511 (N_5511,N_1370,N_534);
nand U5512 (N_5512,N_41,N_183);
nand U5513 (N_5513,N_520,N_1116);
nand U5514 (N_5514,N_3101,N_2620);
xnor U5515 (N_5515,N_2737,N_2069);
nand U5516 (N_5516,N_2883,N_1785);
and U5517 (N_5517,N_1135,N_1633);
nand U5518 (N_5518,N_772,N_1075);
nand U5519 (N_5519,N_2026,N_365);
xor U5520 (N_5520,N_1157,N_1435);
or U5521 (N_5521,N_1131,N_2647);
nor U5522 (N_5522,N_2153,N_2707);
xnor U5523 (N_5523,N_2467,N_1168);
or U5524 (N_5524,N_2182,N_2981);
xor U5525 (N_5525,N_936,N_2187);
nor U5526 (N_5526,N_1977,N_631);
or U5527 (N_5527,N_1974,N_2789);
nor U5528 (N_5528,N_2801,N_1509);
and U5529 (N_5529,N_1838,N_1716);
nor U5530 (N_5530,N_327,N_198);
nand U5531 (N_5531,N_309,N_1194);
nor U5532 (N_5532,N_1087,N_2126);
nor U5533 (N_5533,N_1672,N_2068);
xor U5534 (N_5534,N_2308,N_2673);
xor U5535 (N_5535,N_956,N_1927);
nor U5536 (N_5536,N_8,N_525);
nand U5537 (N_5537,N_1563,N_2291);
xor U5538 (N_5538,N_1565,N_731);
nor U5539 (N_5539,N_304,N_2908);
and U5540 (N_5540,N_982,N_2089);
or U5541 (N_5541,N_512,N_896);
nand U5542 (N_5542,N_1989,N_2741);
nor U5543 (N_5543,N_931,N_660);
nor U5544 (N_5544,N_880,N_1236);
nand U5545 (N_5545,N_2158,N_620);
xnor U5546 (N_5546,N_2122,N_1278);
xor U5547 (N_5547,N_3011,N_2281);
and U5548 (N_5548,N_147,N_1254);
nor U5549 (N_5549,N_286,N_593);
and U5550 (N_5550,N_2916,N_2615);
xnor U5551 (N_5551,N_1006,N_2783);
nand U5552 (N_5552,N_1068,N_2456);
nor U5553 (N_5553,N_629,N_2302);
or U5554 (N_5554,N_1444,N_2463);
xor U5555 (N_5555,N_1043,N_2279);
and U5556 (N_5556,N_1810,N_1967);
or U5557 (N_5557,N_1822,N_1788);
and U5558 (N_5558,N_528,N_187);
or U5559 (N_5559,N_205,N_1760);
and U5560 (N_5560,N_363,N_1910);
nor U5561 (N_5561,N_2093,N_402);
xnor U5562 (N_5562,N_352,N_251);
and U5563 (N_5563,N_1625,N_3079);
nor U5564 (N_5564,N_2558,N_1050);
or U5565 (N_5565,N_248,N_2910);
or U5566 (N_5566,N_231,N_1274);
nor U5567 (N_5567,N_734,N_2124);
or U5568 (N_5568,N_1231,N_1279);
and U5569 (N_5569,N_2001,N_1268);
nor U5570 (N_5570,N_1784,N_941);
nor U5571 (N_5571,N_1556,N_578);
xnor U5572 (N_5572,N_1554,N_2882);
nor U5573 (N_5573,N_2361,N_2427);
xnor U5574 (N_5574,N_1906,N_1276);
xor U5575 (N_5575,N_1220,N_232);
or U5576 (N_5576,N_257,N_2942);
nor U5577 (N_5577,N_2365,N_2188);
nand U5578 (N_5578,N_100,N_2241);
nor U5579 (N_5579,N_1006,N_1485);
xor U5580 (N_5580,N_2335,N_2787);
nor U5581 (N_5581,N_1882,N_732);
nand U5582 (N_5582,N_116,N_1129);
nor U5583 (N_5583,N_2186,N_2646);
nor U5584 (N_5584,N_2566,N_2348);
xnor U5585 (N_5585,N_517,N_3108);
or U5586 (N_5586,N_1711,N_1565);
and U5587 (N_5587,N_586,N_1858);
nor U5588 (N_5588,N_595,N_2624);
nand U5589 (N_5589,N_2241,N_2404);
xor U5590 (N_5590,N_590,N_2732);
nand U5591 (N_5591,N_218,N_2021);
nand U5592 (N_5592,N_1586,N_1512);
xnor U5593 (N_5593,N_956,N_58);
nor U5594 (N_5594,N_3072,N_2189);
and U5595 (N_5595,N_3119,N_2472);
nand U5596 (N_5596,N_2680,N_2035);
and U5597 (N_5597,N_1543,N_2255);
xnor U5598 (N_5598,N_529,N_128);
and U5599 (N_5599,N_2077,N_1982);
xnor U5600 (N_5600,N_58,N_1086);
nand U5601 (N_5601,N_199,N_2580);
nor U5602 (N_5602,N_1008,N_2716);
and U5603 (N_5603,N_1968,N_831);
xor U5604 (N_5604,N_856,N_2886);
xnor U5605 (N_5605,N_632,N_2794);
nand U5606 (N_5606,N_1893,N_635);
xnor U5607 (N_5607,N_1557,N_2758);
or U5608 (N_5608,N_808,N_439);
and U5609 (N_5609,N_1994,N_2227);
or U5610 (N_5610,N_1528,N_3105);
xnor U5611 (N_5611,N_1238,N_529);
and U5612 (N_5612,N_947,N_982);
or U5613 (N_5613,N_2635,N_160);
and U5614 (N_5614,N_597,N_1196);
and U5615 (N_5615,N_1152,N_93);
nand U5616 (N_5616,N_1398,N_2102);
or U5617 (N_5617,N_1708,N_2563);
or U5618 (N_5618,N_463,N_1739);
or U5619 (N_5619,N_3118,N_828);
xor U5620 (N_5620,N_1000,N_8);
xor U5621 (N_5621,N_216,N_3117);
nand U5622 (N_5622,N_1140,N_1709);
nand U5623 (N_5623,N_1294,N_1090);
nor U5624 (N_5624,N_2311,N_2573);
nor U5625 (N_5625,N_3072,N_909);
or U5626 (N_5626,N_2190,N_2052);
and U5627 (N_5627,N_1511,N_2108);
nor U5628 (N_5628,N_2274,N_1799);
or U5629 (N_5629,N_1606,N_811);
nor U5630 (N_5630,N_2314,N_755);
nor U5631 (N_5631,N_112,N_1084);
and U5632 (N_5632,N_3069,N_133);
nor U5633 (N_5633,N_127,N_1162);
or U5634 (N_5634,N_948,N_2831);
xnor U5635 (N_5635,N_1395,N_945);
nand U5636 (N_5636,N_803,N_2292);
xnor U5637 (N_5637,N_488,N_1744);
nand U5638 (N_5638,N_2053,N_492);
or U5639 (N_5639,N_1975,N_1077);
and U5640 (N_5640,N_1998,N_1818);
or U5641 (N_5641,N_2888,N_2128);
xor U5642 (N_5642,N_1552,N_1119);
xnor U5643 (N_5643,N_2830,N_2218);
nor U5644 (N_5644,N_2462,N_1189);
and U5645 (N_5645,N_464,N_2504);
or U5646 (N_5646,N_905,N_3046);
or U5647 (N_5647,N_2276,N_2359);
and U5648 (N_5648,N_2406,N_281);
nand U5649 (N_5649,N_2274,N_1307);
xnor U5650 (N_5650,N_554,N_562);
or U5651 (N_5651,N_399,N_1005);
nand U5652 (N_5652,N_2178,N_1995);
nand U5653 (N_5653,N_1615,N_3029);
nor U5654 (N_5654,N_1705,N_665);
nor U5655 (N_5655,N_1780,N_1905);
and U5656 (N_5656,N_2846,N_1872);
nand U5657 (N_5657,N_1692,N_2962);
or U5658 (N_5658,N_2171,N_1985);
and U5659 (N_5659,N_345,N_1241);
or U5660 (N_5660,N_2606,N_1865);
nor U5661 (N_5661,N_2680,N_1996);
and U5662 (N_5662,N_3014,N_1112);
nor U5663 (N_5663,N_1961,N_3116);
and U5664 (N_5664,N_1066,N_1908);
and U5665 (N_5665,N_564,N_2118);
nor U5666 (N_5666,N_1665,N_1108);
and U5667 (N_5667,N_2199,N_2963);
and U5668 (N_5668,N_2807,N_676);
xor U5669 (N_5669,N_1340,N_1353);
and U5670 (N_5670,N_1532,N_2223);
nand U5671 (N_5671,N_1024,N_1408);
nand U5672 (N_5672,N_536,N_2277);
nor U5673 (N_5673,N_1517,N_676);
or U5674 (N_5674,N_914,N_997);
nor U5675 (N_5675,N_1517,N_206);
nand U5676 (N_5676,N_3082,N_952);
or U5677 (N_5677,N_1408,N_765);
nor U5678 (N_5678,N_2676,N_3122);
xnor U5679 (N_5679,N_1749,N_2099);
or U5680 (N_5680,N_140,N_1396);
xor U5681 (N_5681,N_572,N_1814);
nand U5682 (N_5682,N_3056,N_373);
xor U5683 (N_5683,N_1617,N_9);
xor U5684 (N_5684,N_1012,N_2868);
or U5685 (N_5685,N_2379,N_2695);
nor U5686 (N_5686,N_2278,N_462);
xor U5687 (N_5687,N_2624,N_1704);
xnor U5688 (N_5688,N_2126,N_995);
nand U5689 (N_5689,N_228,N_97);
xnor U5690 (N_5690,N_1584,N_1653);
nor U5691 (N_5691,N_766,N_2768);
and U5692 (N_5692,N_2795,N_1965);
and U5693 (N_5693,N_383,N_99);
xnor U5694 (N_5694,N_1422,N_1160);
xor U5695 (N_5695,N_2746,N_1749);
or U5696 (N_5696,N_1277,N_1578);
and U5697 (N_5697,N_1934,N_1073);
xor U5698 (N_5698,N_1107,N_2930);
xor U5699 (N_5699,N_1491,N_2846);
or U5700 (N_5700,N_2175,N_22);
and U5701 (N_5701,N_1516,N_2569);
and U5702 (N_5702,N_3100,N_1946);
nor U5703 (N_5703,N_809,N_974);
nand U5704 (N_5704,N_1300,N_3068);
nor U5705 (N_5705,N_951,N_1913);
nand U5706 (N_5706,N_2865,N_2233);
and U5707 (N_5707,N_390,N_1181);
nand U5708 (N_5708,N_223,N_2395);
nand U5709 (N_5709,N_1798,N_1406);
xnor U5710 (N_5710,N_2383,N_1317);
nor U5711 (N_5711,N_2755,N_953);
or U5712 (N_5712,N_1209,N_213);
nor U5713 (N_5713,N_559,N_25);
nor U5714 (N_5714,N_1516,N_1021);
nor U5715 (N_5715,N_1718,N_639);
nand U5716 (N_5716,N_2284,N_2706);
or U5717 (N_5717,N_1059,N_3041);
xnor U5718 (N_5718,N_223,N_2984);
xnor U5719 (N_5719,N_3,N_2780);
xor U5720 (N_5720,N_1742,N_2183);
xnor U5721 (N_5721,N_1713,N_1546);
or U5722 (N_5722,N_2631,N_2280);
nor U5723 (N_5723,N_1181,N_2786);
xnor U5724 (N_5724,N_753,N_1789);
or U5725 (N_5725,N_873,N_937);
nor U5726 (N_5726,N_2343,N_452);
xor U5727 (N_5727,N_664,N_2578);
nor U5728 (N_5728,N_1801,N_1158);
nor U5729 (N_5729,N_459,N_1145);
xnor U5730 (N_5730,N_3045,N_2378);
and U5731 (N_5731,N_2783,N_2311);
or U5732 (N_5732,N_1036,N_2949);
xor U5733 (N_5733,N_2958,N_2227);
nand U5734 (N_5734,N_2061,N_2527);
xor U5735 (N_5735,N_1766,N_1326);
xnor U5736 (N_5736,N_2461,N_923);
xor U5737 (N_5737,N_212,N_2405);
xnor U5738 (N_5738,N_670,N_99);
and U5739 (N_5739,N_2330,N_2480);
and U5740 (N_5740,N_2263,N_2369);
xnor U5741 (N_5741,N_81,N_1654);
or U5742 (N_5742,N_1484,N_2278);
nand U5743 (N_5743,N_1773,N_2211);
or U5744 (N_5744,N_2630,N_2560);
nand U5745 (N_5745,N_871,N_1867);
nor U5746 (N_5746,N_1922,N_627);
and U5747 (N_5747,N_1162,N_1998);
nor U5748 (N_5748,N_157,N_2428);
or U5749 (N_5749,N_2757,N_588);
nor U5750 (N_5750,N_2914,N_1910);
or U5751 (N_5751,N_657,N_91);
nand U5752 (N_5752,N_2713,N_2480);
xor U5753 (N_5753,N_1355,N_2973);
nand U5754 (N_5754,N_1207,N_1003);
and U5755 (N_5755,N_967,N_2345);
or U5756 (N_5756,N_193,N_2313);
and U5757 (N_5757,N_2471,N_2336);
xnor U5758 (N_5758,N_453,N_985);
nand U5759 (N_5759,N_497,N_1777);
nor U5760 (N_5760,N_608,N_2645);
and U5761 (N_5761,N_276,N_2939);
nor U5762 (N_5762,N_2889,N_1987);
or U5763 (N_5763,N_1406,N_2177);
xor U5764 (N_5764,N_669,N_784);
nor U5765 (N_5765,N_1833,N_1400);
xnor U5766 (N_5766,N_1617,N_781);
nand U5767 (N_5767,N_2255,N_1143);
xnor U5768 (N_5768,N_2110,N_1341);
nand U5769 (N_5769,N_598,N_1347);
xor U5770 (N_5770,N_1892,N_1952);
nand U5771 (N_5771,N_540,N_2484);
nor U5772 (N_5772,N_909,N_2183);
and U5773 (N_5773,N_2547,N_1366);
nor U5774 (N_5774,N_1972,N_2658);
and U5775 (N_5775,N_728,N_2555);
or U5776 (N_5776,N_2925,N_1138);
and U5777 (N_5777,N_1498,N_3097);
nand U5778 (N_5778,N_1708,N_216);
nor U5779 (N_5779,N_1063,N_1478);
nor U5780 (N_5780,N_1605,N_1259);
nand U5781 (N_5781,N_789,N_1399);
xnor U5782 (N_5782,N_1744,N_462);
nand U5783 (N_5783,N_346,N_2740);
and U5784 (N_5784,N_1692,N_1576);
and U5785 (N_5785,N_2705,N_557);
or U5786 (N_5786,N_989,N_2385);
nor U5787 (N_5787,N_1603,N_1506);
xor U5788 (N_5788,N_2404,N_1030);
xor U5789 (N_5789,N_612,N_2999);
nand U5790 (N_5790,N_1323,N_710);
nand U5791 (N_5791,N_2167,N_49);
and U5792 (N_5792,N_1277,N_1410);
and U5793 (N_5793,N_611,N_1256);
or U5794 (N_5794,N_2535,N_2540);
nand U5795 (N_5795,N_317,N_3107);
xor U5796 (N_5796,N_30,N_2174);
nand U5797 (N_5797,N_211,N_992);
and U5798 (N_5798,N_1341,N_1421);
nand U5799 (N_5799,N_250,N_2067);
nand U5800 (N_5800,N_2623,N_608);
and U5801 (N_5801,N_2510,N_2058);
and U5802 (N_5802,N_2627,N_2647);
xor U5803 (N_5803,N_2137,N_1268);
nand U5804 (N_5804,N_111,N_2885);
and U5805 (N_5805,N_1848,N_985);
or U5806 (N_5806,N_2617,N_364);
nand U5807 (N_5807,N_2737,N_3123);
and U5808 (N_5808,N_617,N_2922);
nor U5809 (N_5809,N_99,N_170);
nor U5810 (N_5810,N_911,N_1476);
or U5811 (N_5811,N_2539,N_2331);
nand U5812 (N_5812,N_2788,N_2872);
nor U5813 (N_5813,N_338,N_625);
and U5814 (N_5814,N_2183,N_3114);
and U5815 (N_5815,N_1533,N_1712);
or U5816 (N_5816,N_2442,N_789);
xnor U5817 (N_5817,N_1005,N_1578);
and U5818 (N_5818,N_1647,N_1286);
nor U5819 (N_5819,N_1574,N_450);
xor U5820 (N_5820,N_2694,N_1516);
or U5821 (N_5821,N_2867,N_1600);
nand U5822 (N_5822,N_2657,N_123);
or U5823 (N_5823,N_376,N_1625);
nand U5824 (N_5824,N_3080,N_2199);
and U5825 (N_5825,N_2045,N_2700);
nor U5826 (N_5826,N_691,N_1769);
or U5827 (N_5827,N_1984,N_1122);
xor U5828 (N_5828,N_199,N_2412);
xor U5829 (N_5829,N_1903,N_2447);
or U5830 (N_5830,N_2059,N_1671);
xor U5831 (N_5831,N_3053,N_2038);
nor U5832 (N_5832,N_2276,N_453);
xnor U5833 (N_5833,N_2941,N_1138);
nand U5834 (N_5834,N_155,N_1017);
nand U5835 (N_5835,N_1389,N_417);
nand U5836 (N_5836,N_1405,N_2612);
nor U5837 (N_5837,N_1505,N_365);
nor U5838 (N_5838,N_1521,N_2914);
nand U5839 (N_5839,N_2015,N_1226);
and U5840 (N_5840,N_1575,N_1279);
or U5841 (N_5841,N_2039,N_2907);
xor U5842 (N_5842,N_1422,N_718);
and U5843 (N_5843,N_1791,N_1257);
and U5844 (N_5844,N_2556,N_1868);
and U5845 (N_5845,N_2227,N_1339);
nor U5846 (N_5846,N_1853,N_1671);
nor U5847 (N_5847,N_2479,N_240);
and U5848 (N_5848,N_1888,N_660);
nand U5849 (N_5849,N_604,N_3099);
nor U5850 (N_5850,N_1354,N_2802);
and U5851 (N_5851,N_1610,N_2573);
nand U5852 (N_5852,N_705,N_942);
and U5853 (N_5853,N_1834,N_460);
or U5854 (N_5854,N_1580,N_1814);
nor U5855 (N_5855,N_1366,N_2463);
and U5856 (N_5856,N_2170,N_1166);
nor U5857 (N_5857,N_856,N_804);
nor U5858 (N_5858,N_222,N_2455);
nor U5859 (N_5859,N_1090,N_2560);
or U5860 (N_5860,N_2859,N_1275);
xnor U5861 (N_5861,N_136,N_2836);
and U5862 (N_5862,N_2501,N_2768);
and U5863 (N_5863,N_1533,N_2741);
nand U5864 (N_5864,N_2859,N_1790);
nand U5865 (N_5865,N_719,N_3064);
nand U5866 (N_5866,N_1397,N_2639);
or U5867 (N_5867,N_2405,N_2844);
and U5868 (N_5868,N_2803,N_168);
and U5869 (N_5869,N_1447,N_1426);
nor U5870 (N_5870,N_2542,N_2762);
or U5871 (N_5871,N_2644,N_565);
xnor U5872 (N_5872,N_1032,N_1727);
xor U5873 (N_5873,N_870,N_1783);
xor U5874 (N_5874,N_2444,N_2877);
or U5875 (N_5875,N_1367,N_1176);
and U5876 (N_5876,N_929,N_618);
or U5877 (N_5877,N_1878,N_2272);
nor U5878 (N_5878,N_736,N_347);
and U5879 (N_5879,N_227,N_2725);
nand U5880 (N_5880,N_2810,N_2415);
nand U5881 (N_5881,N_165,N_463);
or U5882 (N_5882,N_1673,N_1381);
and U5883 (N_5883,N_2924,N_1856);
and U5884 (N_5884,N_84,N_555);
nor U5885 (N_5885,N_2490,N_824);
or U5886 (N_5886,N_1240,N_1944);
and U5887 (N_5887,N_1617,N_1847);
nand U5888 (N_5888,N_464,N_867);
nand U5889 (N_5889,N_1862,N_2653);
or U5890 (N_5890,N_1083,N_3119);
and U5891 (N_5891,N_296,N_3075);
xor U5892 (N_5892,N_1867,N_2511);
and U5893 (N_5893,N_2078,N_23);
nor U5894 (N_5894,N_768,N_3030);
nor U5895 (N_5895,N_892,N_2095);
nand U5896 (N_5896,N_2396,N_36);
or U5897 (N_5897,N_1098,N_2316);
and U5898 (N_5898,N_3040,N_1940);
nand U5899 (N_5899,N_1876,N_1393);
or U5900 (N_5900,N_2028,N_1529);
nand U5901 (N_5901,N_64,N_1507);
nand U5902 (N_5902,N_2258,N_721);
xnor U5903 (N_5903,N_286,N_2174);
nor U5904 (N_5904,N_2283,N_2859);
nand U5905 (N_5905,N_1993,N_2009);
and U5906 (N_5906,N_319,N_487);
nand U5907 (N_5907,N_1010,N_286);
or U5908 (N_5908,N_356,N_1228);
or U5909 (N_5909,N_994,N_2977);
nor U5910 (N_5910,N_2607,N_1685);
nand U5911 (N_5911,N_2448,N_1326);
nand U5912 (N_5912,N_1238,N_1557);
and U5913 (N_5913,N_679,N_90);
and U5914 (N_5914,N_670,N_1723);
and U5915 (N_5915,N_1959,N_1230);
and U5916 (N_5916,N_96,N_13);
nand U5917 (N_5917,N_2039,N_3078);
xnor U5918 (N_5918,N_1541,N_2029);
nand U5919 (N_5919,N_2771,N_1835);
nor U5920 (N_5920,N_275,N_659);
xnor U5921 (N_5921,N_2426,N_1776);
or U5922 (N_5922,N_2820,N_1531);
xor U5923 (N_5923,N_1440,N_1763);
nor U5924 (N_5924,N_1868,N_2960);
nand U5925 (N_5925,N_1800,N_2806);
nor U5926 (N_5926,N_824,N_390);
or U5927 (N_5927,N_3069,N_262);
xor U5928 (N_5928,N_551,N_157);
and U5929 (N_5929,N_1881,N_1362);
xor U5930 (N_5930,N_1819,N_1486);
nor U5931 (N_5931,N_238,N_2849);
and U5932 (N_5932,N_3044,N_2344);
nor U5933 (N_5933,N_2738,N_2057);
xor U5934 (N_5934,N_1880,N_657);
xor U5935 (N_5935,N_2578,N_381);
xnor U5936 (N_5936,N_2925,N_3009);
nand U5937 (N_5937,N_473,N_1409);
nor U5938 (N_5938,N_973,N_1421);
or U5939 (N_5939,N_2439,N_2566);
xor U5940 (N_5940,N_576,N_1294);
and U5941 (N_5941,N_333,N_2642);
or U5942 (N_5942,N_1426,N_46);
and U5943 (N_5943,N_895,N_624);
xor U5944 (N_5944,N_2353,N_2115);
or U5945 (N_5945,N_2404,N_1672);
xor U5946 (N_5946,N_2550,N_1898);
nor U5947 (N_5947,N_2235,N_2540);
nand U5948 (N_5948,N_1434,N_3036);
or U5949 (N_5949,N_614,N_2746);
nand U5950 (N_5950,N_1578,N_1522);
or U5951 (N_5951,N_1488,N_1836);
and U5952 (N_5952,N_1536,N_552);
xnor U5953 (N_5953,N_643,N_487);
xnor U5954 (N_5954,N_1475,N_2515);
xor U5955 (N_5955,N_1075,N_833);
xnor U5956 (N_5956,N_2092,N_2936);
nand U5957 (N_5957,N_437,N_2045);
or U5958 (N_5958,N_2040,N_2193);
xnor U5959 (N_5959,N_715,N_1187);
nor U5960 (N_5960,N_1390,N_1329);
xor U5961 (N_5961,N_2994,N_2926);
and U5962 (N_5962,N_1757,N_1264);
and U5963 (N_5963,N_33,N_2559);
nor U5964 (N_5964,N_737,N_151);
and U5965 (N_5965,N_1828,N_2184);
nor U5966 (N_5966,N_208,N_326);
nand U5967 (N_5967,N_162,N_974);
or U5968 (N_5968,N_2406,N_172);
xor U5969 (N_5969,N_628,N_2130);
or U5970 (N_5970,N_589,N_2518);
or U5971 (N_5971,N_1331,N_839);
and U5972 (N_5972,N_2826,N_1218);
nor U5973 (N_5973,N_449,N_2177);
nand U5974 (N_5974,N_1639,N_1385);
nor U5975 (N_5975,N_3031,N_3025);
nor U5976 (N_5976,N_1937,N_423);
or U5977 (N_5977,N_2209,N_1577);
and U5978 (N_5978,N_2787,N_474);
xnor U5979 (N_5979,N_1795,N_1449);
nor U5980 (N_5980,N_2139,N_1708);
nor U5981 (N_5981,N_1390,N_747);
xor U5982 (N_5982,N_1520,N_2381);
xor U5983 (N_5983,N_2544,N_738);
xor U5984 (N_5984,N_377,N_294);
nor U5985 (N_5985,N_2950,N_1193);
or U5986 (N_5986,N_899,N_1255);
xor U5987 (N_5987,N_3085,N_681);
and U5988 (N_5988,N_1753,N_428);
xor U5989 (N_5989,N_2433,N_120);
nand U5990 (N_5990,N_1400,N_2533);
xnor U5991 (N_5991,N_574,N_1628);
or U5992 (N_5992,N_1252,N_360);
and U5993 (N_5993,N_1173,N_1475);
xor U5994 (N_5994,N_1516,N_2973);
xnor U5995 (N_5995,N_2565,N_818);
xor U5996 (N_5996,N_3083,N_475);
xnor U5997 (N_5997,N_1823,N_2602);
or U5998 (N_5998,N_692,N_1330);
nand U5999 (N_5999,N_1368,N_3037);
and U6000 (N_6000,N_1065,N_1371);
and U6001 (N_6001,N_2798,N_661);
and U6002 (N_6002,N_2562,N_1520);
or U6003 (N_6003,N_75,N_2110);
nor U6004 (N_6004,N_2064,N_331);
or U6005 (N_6005,N_3002,N_1046);
or U6006 (N_6006,N_1919,N_1977);
nor U6007 (N_6007,N_1905,N_1772);
nor U6008 (N_6008,N_1267,N_1885);
nor U6009 (N_6009,N_290,N_1039);
or U6010 (N_6010,N_263,N_2325);
or U6011 (N_6011,N_1340,N_2233);
nand U6012 (N_6012,N_119,N_2433);
or U6013 (N_6013,N_2183,N_3098);
nand U6014 (N_6014,N_2296,N_43);
or U6015 (N_6015,N_2131,N_2988);
xor U6016 (N_6016,N_110,N_2927);
nor U6017 (N_6017,N_86,N_2518);
xor U6018 (N_6018,N_589,N_2680);
and U6019 (N_6019,N_1664,N_696);
nand U6020 (N_6020,N_2740,N_2202);
or U6021 (N_6021,N_547,N_2691);
and U6022 (N_6022,N_746,N_2146);
or U6023 (N_6023,N_1263,N_1579);
nand U6024 (N_6024,N_2849,N_837);
nor U6025 (N_6025,N_1131,N_1339);
and U6026 (N_6026,N_2167,N_196);
and U6027 (N_6027,N_1669,N_1405);
nand U6028 (N_6028,N_1859,N_1796);
or U6029 (N_6029,N_1229,N_2481);
xor U6030 (N_6030,N_1026,N_2460);
and U6031 (N_6031,N_2237,N_1978);
and U6032 (N_6032,N_95,N_1925);
or U6033 (N_6033,N_146,N_864);
or U6034 (N_6034,N_2857,N_1295);
nand U6035 (N_6035,N_293,N_489);
nand U6036 (N_6036,N_191,N_320);
nor U6037 (N_6037,N_3104,N_1265);
and U6038 (N_6038,N_66,N_306);
xor U6039 (N_6039,N_954,N_1554);
or U6040 (N_6040,N_915,N_1380);
nand U6041 (N_6041,N_534,N_952);
and U6042 (N_6042,N_1447,N_2540);
or U6043 (N_6043,N_839,N_1908);
nor U6044 (N_6044,N_1820,N_1362);
xor U6045 (N_6045,N_679,N_1564);
and U6046 (N_6046,N_1583,N_569);
and U6047 (N_6047,N_1805,N_1736);
or U6048 (N_6048,N_84,N_1875);
and U6049 (N_6049,N_1423,N_1373);
xor U6050 (N_6050,N_2280,N_2880);
nor U6051 (N_6051,N_3118,N_1349);
nand U6052 (N_6052,N_2967,N_2657);
xor U6053 (N_6053,N_2751,N_507);
nand U6054 (N_6054,N_1333,N_1647);
nand U6055 (N_6055,N_2001,N_2534);
or U6056 (N_6056,N_1992,N_1649);
or U6057 (N_6057,N_248,N_2539);
nand U6058 (N_6058,N_138,N_322);
nor U6059 (N_6059,N_1930,N_680);
nand U6060 (N_6060,N_1524,N_991);
or U6061 (N_6061,N_1550,N_1685);
nor U6062 (N_6062,N_180,N_2903);
or U6063 (N_6063,N_281,N_2727);
and U6064 (N_6064,N_821,N_3078);
nand U6065 (N_6065,N_534,N_69);
xor U6066 (N_6066,N_1569,N_174);
and U6067 (N_6067,N_2486,N_2928);
or U6068 (N_6068,N_2018,N_937);
nand U6069 (N_6069,N_3053,N_2940);
nand U6070 (N_6070,N_1202,N_2402);
nor U6071 (N_6071,N_2886,N_2487);
and U6072 (N_6072,N_1914,N_816);
xor U6073 (N_6073,N_2720,N_351);
nand U6074 (N_6074,N_723,N_1921);
nor U6075 (N_6075,N_837,N_494);
nand U6076 (N_6076,N_2330,N_1863);
and U6077 (N_6077,N_1318,N_2310);
and U6078 (N_6078,N_1874,N_1502);
xor U6079 (N_6079,N_2537,N_3093);
nand U6080 (N_6080,N_2267,N_2455);
nand U6081 (N_6081,N_2522,N_947);
or U6082 (N_6082,N_1090,N_2417);
nand U6083 (N_6083,N_2932,N_1337);
xnor U6084 (N_6084,N_1794,N_1252);
nand U6085 (N_6085,N_1293,N_930);
and U6086 (N_6086,N_1814,N_1112);
xor U6087 (N_6087,N_1654,N_2716);
nand U6088 (N_6088,N_333,N_2698);
or U6089 (N_6089,N_1113,N_768);
xnor U6090 (N_6090,N_1205,N_1016);
xnor U6091 (N_6091,N_900,N_1630);
xor U6092 (N_6092,N_1544,N_1096);
nor U6093 (N_6093,N_1029,N_2298);
or U6094 (N_6094,N_1236,N_2629);
nor U6095 (N_6095,N_2571,N_2681);
or U6096 (N_6096,N_2497,N_832);
xor U6097 (N_6097,N_2384,N_1187);
nand U6098 (N_6098,N_1319,N_3051);
or U6099 (N_6099,N_1613,N_2142);
nand U6100 (N_6100,N_685,N_1919);
xor U6101 (N_6101,N_1420,N_1918);
or U6102 (N_6102,N_915,N_1801);
nor U6103 (N_6103,N_403,N_2451);
nand U6104 (N_6104,N_2984,N_2192);
or U6105 (N_6105,N_267,N_1871);
nand U6106 (N_6106,N_2672,N_2045);
nand U6107 (N_6107,N_1755,N_143);
or U6108 (N_6108,N_1152,N_2048);
xor U6109 (N_6109,N_2911,N_2346);
nand U6110 (N_6110,N_415,N_1528);
nand U6111 (N_6111,N_2736,N_2877);
nand U6112 (N_6112,N_2218,N_2536);
or U6113 (N_6113,N_2408,N_1358);
xnor U6114 (N_6114,N_2176,N_620);
nor U6115 (N_6115,N_3029,N_231);
and U6116 (N_6116,N_1742,N_702);
nor U6117 (N_6117,N_1262,N_1710);
nor U6118 (N_6118,N_1963,N_1868);
nand U6119 (N_6119,N_418,N_1175);
nand U6120 (N_6120,N_1780,N_2350);
nor U6121 (N_6121,N_200,N_829);
xnor U6122 (N_6122,N_2090,N_59);
and U6123 (N_6123,N_651,N_455);
nand U6124 (N_6124,N_1552,N_833);
xnor U6125 (N_6125,N_662,N_112);
and U6126 (N_6126,N_996,N_1579);
nand U6127 (N_6127,N_2886,N_1778);
xnor U6128 (N_6128,N_357,N_316);
nor U6129 (N_6129,N_556,N_525);
or U6130 (N_6130,N_2110,N_2558);
xor U6131 (N_6131,N_2022,N_430);
xnor U6132 (N_6132,N_664,N_486);
nand U6133 (N_6133,N_2779,N_1050);
nand U6134 (N_6134,N_154,N_709);
nand U6135 (N_6135,N_2837,N_662);
or U6136 (N_6136,N_872,N_296);
or U6137 (N_6137,N_2994,N_1286);
and U6138 (N_6138,N_1237,N_300);
nor U6139 (N_6139,N_2689,N_630);
nor U6140 (N_6140,N_835,N_1403);
xnor U6141 (N_6141,N_2777,N_2242);
or U6142 (N_6142,N_2389,N_1070);
nor U6143 (N_6143,N_2304,N_2400);
or U6144 (N_6144,N_3040,N_1129);
nor U6145 (N_6145,N_2550,N_328);
or U6146 (N_6146,N_47,N_2216);
nor U6147 (N_6147,N_2995,N_2460);
xnor U6148 (N_6148,N_1186,N_3020);
or U6149 (N_6149,N_2958,N_940);
or U6150 (N_6150,N_2685,N_2273);
nor U6151 (N_6151,N_1765,N_1873);
or U6152 (N_6152,N_406,N_1563);
or U6153 (N_6153,N_2062,N_2386);
nor U6154 (N_6154,N_1071,N_1668);
xor U6155 (N_6155,N_497,N_1608);
and U6156 (N_6156,N_2846,N_425);
and U6157 (N_6157,N_1589,N_1776);
xnor U6158 (N_6158,N_1881,N_862);
and U6159 (N_6159,N_2084,N_1076);
or U6160 (N_6160,N_2600,N_837);
and U6161 (N_6161,N_3072,N_2304);
and U6162 (N_6162,N_420,N_2787);
xnor U6163 (N_6163,N_1005,N_1141);
xnor U6164 (N_6164,N_992,N_1855);
or U6165 (N_6165,N_2248,N_1809);
nor U6166 (N_6166,N_971,N_1921);
nor U6167 (N_6167,N_2055,N_2854);
xor U6168 (N_6168,N_1196,N_368);
nand U6169 (N_6169,N_351,N_2367);
and U6170 (N_6170,N_135,N_1326);
nand U6171 (N_6171,N_1003,N_1768);
and U6172 (N_6172,N_173,N_1120);
or U6173 (N_6173,N_1093,N_1492);
nor U6174 (N_6174,N_1922,N_2826);
nand U6175 (N_6175,N_167,N_2130);
nor U6176 (N_6176,N_1337,N_1958);
nor U6177 (N_6177,N_2297,N_644);
xor U6178 (N_6178,N_2171,N_510);
xor U6179 (N_6179,N_1561,N_1079);
xor U6180 (N_6180,N_2686,N_220);
nand U6181 (N_6181,N_49,N_2543);
or U6182 (N_6182,N_1992,N_1477);
nor U6183 (N_6183,N_2201,N_2321);
or U6184 (N_6184,N_743,N_741);
xor U6185 (N_6185,N_858,N_2043);
and U6186 (N_6186,N_603,N_122);
nand U6187 (N_6187,N_292,N_1608);
xnor U6188 (N_6188,N_199,N_2850);
and U6189 (N_6189,N_1717,N_1310);
nand U6190 (N_6190,N_2675,N_1363);
xnor U6191 (N_6191,N_2993,N_2363);
or U6192 (N_6192,N_631,N_341);
xnor U6193 (N_6193,N_1221,N_1804);
and U6194 (N_6194,N_733,N_170);
or U6195 (N_6195,N_1716,N_2210);
xor U6196 (N_6196,N_2610,N_1239);
nand U6197 (N_6197,N_1243,N_3120);
and U6198 (N_6198,N_819,N_2423);
nor U6199 (N_6199,N_1503,N_341);
nand U6200 (N_6200,N_2896,N_2262);
xor U6201 (N_6201,N_769,N_787);
nor U6202 (N_6202,N_830,N_2380);
or U6203 (N_6203,N_1155,N_1785);
and U6204 (N_6204,N_2133,N_3014);
xor U6205 (N_6205,N_269,N_2927);
or U6206 (N_6206,N_2697,N_821);
nor U6207 (N_6207,N_487,N_483);
xor U6208 (N_6208,N_2177,N_2889);
or U6209 (N_6209,N_1250,N_790);
nand U6210 (N_6210,N_1758,N_1529);
nand U6211 (N_6211,N_2208,N_152);
nand U6212 (N_6212,N_1024,N_47);
nor U6213 (N_6213,N_3057,N_942);
and U6214 (N_6214,N_718,N_1684);
nor U6215 (N_6215,N_2904,N_2430);
and U6216 (N_6216,N_745,N_1105);
nand U6217 (N_6217,N_1183,N_2011);
and U6218 (N_6218,N_1933,N_1074);
nor U6219 (N_6219,N_2998,N_2614);
nand U6220 (N_6220,N_2550,N_2036);
xnor U6221 (N_6221,N_933,N_1279);
nand U6222 (N_6222,N_937,N_1107);
or U6223 (N_6223,N_2027,N_1395);
nand U6224 (N_6224,N_368,N_1576);
nand U6225 (N_6225,N_824,N_468);
xor U6226 (N_6226,N_1259,N_2082);
nand U6227 (N_6227,N_2007,N_1497);
nor U6228 (N_6228,N_2606,N_2317);
nand U6229 (N_6229,N_2675,N_408);
or U6230 (N_6230,N_3090,N_555);
nand U6231 (N_6231,N_1416,N_37);
nor U6232 (N_6232,N_630,N_2413);
or U6233 (N_6233,N_483,N_2503);
xor U6234 (N_6234,N_1505,N_1017);
xor U6235 (N_6235,N_531,N_305);
or U6236 (N_6236,N_550,N_1351);
or U6237 (N_6237,N_999,N_254);
and U6238 (N_6238,N_1410,N_2241);
or U6239 (N_6239,N_1106,N_2887);
and U6240 (N_6240,N_1019,N_1389);
nor U6241 (N_6241,N_1093,N_1718);
or U6242 (N_6242,N_1132,N_425);
or U6243 (N_6243,N_1162,N_1079);
or U6244 (N_6244,N_1915,N_2459);
nor U6245 (N_6245,N_511,N_2555);
and U6246 (N_6246,N_2099,N_584);
xnor U6247 (N_6247,N_16,N_1183);
or U6248 (N_6248,N_785,N_57);
nand U6249 (N_6249,N_2407,N_2995);
or U6250 (N_6250,N_3463,N_5663);
and U6251 (N_6251,N_5045,N_4555);
xnor U6252 (N_6252,N_6149,N_5390);
xnor U6253 (N_6253,N_4982,N_3848);
or U6254 (N_6254,N_5312,N_5531);
nor U6255 (N_6255,N_5183,N_5159);
nand U6256 (N_6256,N_5788,N_5616);
nor U6257 (N_6257,N_4691,N_4227);
and U6258 (N_6258,N_4729,N_3269);
or U6259 (N_6259,N_4315,N_4815);
nor U6260 (N_6260,N_4138,N_3907);
or U6261 (N_6261,N_4610,N_5562);
nand U6262 (N_6262,N_5011,N_6076);
xor U6263 (N_6263,N_5017,N_3270);
nor U6264 (N_6264,N_5711,N_5622);
xor U6265 (N_6265,N_3179,N_3916);
xnor U6266 (N_6266,N_5796,N_3716);
or U6267 (N_6267,N_3444,N_3814);
nor U6268 (N_6268,N_3898,N_5386);
and U6269 (N_6269,N_5684,N_5307);
and U6270 (N_6270,N_5119,N_4583);
or U6271 (N_6271,N_4503,N_5803);
xor U6272 (N_6272,N_5191,N_3903);
and U6273 (N_6273,N_4410,N_3671);
and U6274 (N_6274,N_5362,N_5528);
nor U6275 (N_6275,N_3466,N_5012);
nor U6276 (N_6276,N_4762,N_3494);
and U6277 (N_6277,N_4591,N_3316);
nand U6278 (N_6278,N_4553,N_4398);
xnor U6279 (N_6279,N_3180,N_3835);
nand U6280 (N_6280,N_6093,N_3993);
nand U6281 (N_6281,N_4873,N_4977);
xor U6282 (N_6282,N_3794,N_5423);
and U6283 (N_6283,N_5300,N_4329);
xnor U6284 (N_6284,N_3811,N_5624);
or U6285 (N_6285,N_6161,N_5908);
xnor U6286 (N_6286,N_5083,N_5403);
xor U6287 (N_6287,N_5208,N_3265);
nand U6288 (N_6288,N_5199,N_4884);
nand U6289 (N_6289,N_5617,N_4914);
nor U6290 (N_6290,N_4737,N_5626);
and U6291 (N_6291,N_6197,N_3820);
or U6292 (N_6292,N_5072,N_5543);
nor U6293 (N_6293,N_5727,N_5775);
or U6294 (N_6294,N_3951,N_4724);
nor U6295 (N_6295,N_5217,N_5063);
xnor U6296 (N_6296,N_3507,N_3165);
nor U6297 (N_6297,N_5211,N_4627);
xnor U6298 (N_6298,N_4129,N_4303);
xnor U6299 (N_6299,N_5640,N_4387);
xor U6300 (N_6300,N_4931,N_6067);
or U6301 (N_6301,N_4402,N_4870);
nand U6302 (N_6302,N_5227,N_5858);
xor U6303 (N_6303,N_5736,N_5262);
nor U6304 (N_6304,N_5077,N_5849);
or U6305 (N_6305,N_6145,N_4214);
nor U6306 (N_6306,N_3302,N_6237);
or U6307 (N_6307,N_5621,N_4996);
and U6308 (N_6308,N_5888,N_5221);
and U6309 (N_6309,N_4649,N_4516);
or U6310 (N_6310,N_3550,N_3245);
nand U6311 (N_6311,N_3796,N_5339);
xnor U6312 (N_6312,N_4279,N_5461);
xor U6313 (N_6313,N_3578,N_5482);
nor U6314 (N_6314,N_3896,N_4442);
or U6315 (N_6315,N_4656,N_5857);
or U6316 (N_6316,N_5812,N_5299);
xnor U6317 (N_6317,N_4060,N_6057);
nor U6318 (N_6318,N_5039,N_5365);
and U6319 (N_6319,N_5337,N_4812);
nor U6320 (N_6320,N_3497,N_5376);
nor U6321 (N_6321,N_4484,N_3751);
xor U6322 (N_6322,N_5925,N_3196);
or U6323 (N_6323,N_3859,N_5181);
nor U6324 (N_6324,N_5085,N_5443);
nand U6325 (N_6325,N_3281,N_5658);
nor U6326 (N_6326,N_6162,N_4789);
xnor U6327 (N_6327,N_3556,N_4770);
and U6328 (N_6328,N_4108,N_5723);
nor U6329 (N_6329,N_4180,N_3944);
or U6330 (N_6330,N_5308,N_3504);
or U6331 (N_6331,N_3523,N_4290);
nand U6332 (N_6332,N_6113,N_4527);
nor U6333 (N_6333,N_4013,N_5468);
xnor U6334 (N_6334,N_6177,N_4838);
nand U6335 (N_6335,N_4694,N_5281);
or U6336 (N_6336,N_4961,N_3841);
nor U6337 (N_6337,N_5135,N_4550);
nor U6338 (N_6338,N_5848,N_5374);
and U6339 (N_6339,N_4302,N_4069);
nor U6340 (N_6340,N_4598,N_3709);
nor U6341 (N_6341,N_5476,N_3478);
and U6342 (N_6342,N_5909,N_5741);
and U6343 (N_6343,N_6074,N_3838);
or U6344 (N_6344,N_6114,N_5398);
and U6345 (N_6345,N_5559,N_4209);
nor U6346 (N_6346,N_5263,N_3276);
or U6347 (N_6347,N_4787,N_3605);
nor U6348 (N_6348,N_5941,N_3666);
xor U6349 (N_6349,N_4744,N_4952);
or U6350 (N_6350,N_5947,N_5876);
and U6351 (N_6351,N_6059,N_5918);
nor U6352 (N_6352,N_4678,N_3579);
nor U6353 (N_6353,N_4839,N_5037);
or U6354 (N_6354,N_5031,N_5514);
or U6355 (N_6355,N_5273,N_3219);
and U6356 (N_6356,N_4029,N_3129);
nor U6357 (N_6357,N_5132,N_4558);
or U6358 (N_6358,N_5597,N_4431);
nand U6359 (N_6359,N_3166,N_3768);
or U6360 (N_6360,N_3503,N_5016);
nand U6361 (N_6361,N_3668,N_3192);
or U6362 (N_6362,N_4505,N_3187);
and U6363 (N_6363,N_4603,N_4749);
nand U6364 (N_6364,N_4507,N_4096);
and U6365 (N_6365,N_4473,N_4814);
nor U6366 (N_6366,N_3942,N_6083);
xor U6367 (N_6367,N_5363,N_4933);
or U6368 (N_6368,N_5146,N_5413);
xnor U6369 (N_6369,N_4418,N_4208);
nor U6370 (N_6370,N_5634,N_5896);
nor U6371 (N_6371,N_3839,N_4150);
xnor U6372 (N_6372,N_3686,N_6196);
or U6373 (N_6373,N_6117,N_6118);
and U6374 (N_6374,N_6061,N_3149);
nor U6375 (N_6375,N_5394,N_4276);
xnor U6376 (N_6376,N_5573,N_3905);
nand U6377 (N_6377,N_5393,N_5831);
xor U6378 (N_6378,N_4490,N_3570);
and U6379 (N_6379,N_3665,N_4712);
xnor U6380 (N_6380,N_5767,N_5582);
or U6381 (N_6381,N_4561,N_3663);
xnor U6382 (N_6382,N_4545,N_3202);
xor U6383 (N_6383,N_4606,N_4786);
nand U6384 (N_6384,N_4761,N_4778);
and U6385 (N_6385,N_3418,N_3986);
or U6386 (N_6386,N_5529,N_4396);
and U6387 (N_6387,N_3296,N_4485);
or U6388 (N_6388,N_3856,N_4187);
and U6389 (N_6389,N_5501,N_3705);
nand U6390 (N_6390,N_3627,N_3528);
or U6391 (N_6391,N_4859,N_5681);
nor U6392 (N_6392,N_5652,N_4014);
nand U6393 (N_6393,N_4270,N_4697);
xnor U6394 (N_6394,N_5030,N_5608);
nor U6395 (N_6395,N_3341,N_4244);
nand U6396 (N_6396,N_5959,N_6070);
and U6397 (N_6397,N_3761,N_5133);
nor U6398 (N_6398,N_5537,N_4866);
nor U6399 (N_6399,N_4582,N_5533);
nor U6400 (N_6400,N_3195,N_5677);
nor U6401 (N_6401,N_3628,N_3176);
xnor U6402 (N_6402,N_4206,N_3152);
and U6403 (N_6403,N_5689,N_5615);
or U6404 (N_6404,N_5752,N_4991);
xor U6405 (N_6405,N_4680,N_4097);
nor U6406 (N_6406,N_6190,N_3130);
nand U6407 (N_6407,N_4532,N_6035);
nor U6408 (N_6408,N_4463,N_4768);
nor U6409 (N_6409,N_6228,N_4035);
nand U6410 (N_6410,N_6064,N_5370);
xor U6411 (N_6411,N_3161,N_5444);
xnor U6412 (N_6412,N_4774,N_5725);
and U6413 (N_6413,N_5309,N_4658);
or U6414 (N_6414,N_4200,N_5686);
or U6415 (N_6415,N_6231,N_6003);
nand U6416 (N_6416,N_3591,N_3428);
xor U6417 (N_6417,N_5619,N_5553);
nand U6418 (N_6418,N_4891,N_4574);
or U6419 (N_6419,N_5259,N_5271);
and U6420 (N_6420,N_4628,N_4347);
and U6421 (N_6421,N_4454,N_3874);
xor U6422 (N_6422,N_4158,N_5161);
and U6423 (N_6423,N_3707,N_4482);
nor U6424 (N_6424,N_4647,N_6096);
and U6425 (N_6425,N_4089,N_5598);
nand U6426 (N_6426,N_3647,N_5167);
xnor U6427 (N_6427,N_3381,N_5983);
nor U6428 (N_6428,N_3831,N_6183);
or U6429 (N_6429,N_4681,N_3810);
nor U6430 (N_6430,N_6198,N_4433);
or U6431 (N_6431,N_4769,N_4047);
nand U6432 (N_6432,N_3800,N_3694);
nand U6433 (N_6433,N_3416,N_4856);
xnor U6434 (N_6434,N_4364,N_3173);
xnor U6435 (N_6435,N_3448,N_5136);
nand U6436 (N_6436,N_5510,N_3978);
nor U6437 (N_6437,N_4183,N_5593);
xor U6438 (N_6438,N_3985,N_4862);
nand U6439 (N_6439,N_3486,N_4515);
xor U6440 (N_6440,N_4900,N_4311);
nand U6441 (N_6441,N_5570,N_3725);
nand U6442 (N_6442,N_3755,N_4796);
nand U6443 (N_6443,N_3169,N_4664);
and U6444 (N_6444,N_3710,N_5743);
and U6445 (N_6445,N_5838,N_3363);
and U6446 (N_6446,N_3894,N_4704);
nor U6447 (N_6447,N_5241,N_4701);
xor U6448 (N_6448,N_4168,N_5919);
xor U6449 (N_6449,N_3275,N_4827);
xor U6450 (N_6450,N_4675,N_3509);
xor U6451 (N_6451,N_5242,N_3759);
nor U6452 (N_6452,N_3357,N_5794);
xor U6453 (N_6453,N_3912,N_3337);
and U6454 (N_6454,N_3421,N_3634);
xnor U6455 (N_6455,N_4995,N_3857);
and U6456 (N_6456,N_3818,N_4058);
or U6457 (N_6457,N_3867,N_5986);
xnor U6458 (N_6458,N_6156,N_5236);
nor U6459 (N_6459,N_3758,N_4958);
and U6460 (N_6460,N_4993,N_4887);
nor U6461 (N_6461,N_4400,N_6013);
or U6462 (N_6462,N_4855,N_4457);
and U6463 (N_6463,N_4167,N_3997);
and U6464 (N_6464,N_5994,N_5409);
nor U6465 (N_6465,N_3359,N_6136);
nand U6466 (N_6466,N_5499,N_3190);
and U6467 (N_6467,N_4243,N_4460);
nand U6468 (N_6468,N_4412,N_6014);
nand U6469 (N_6469,N_5773,N_6009);
nor U6470 (N_6470,N_4381,N_4237);
nand U6471 (N_6471,N_5284,N_4940);
and U6472 (N_6472,N_3368,N_3735);
nand U6473 (N_6473,N_4091,N_5034);
and U6474 (N_6474,N_5556,N_3511);
and U6475 (N_6475,N_4909,N_4772);
nor U6476 (N_6476,N_4001,N_5216);
nand U6477 (N_6477,N_3949,N_4468);
nand U6478 (N_6478,N_5193,N_5505);
nand U6479 (N_6479,N_5209,N_3212);
nand U6480 (N_6480,N_5620,N_5068);
nand U6481 (N_6481,N_3624,N_3536);
and U6482 (N_6482,N_5926,N_3879);
and U6483 (N_6483,N_3643,N_4359);
nor U6484 (N_6484,N_4282,N_4423);
and U6485 (N_6485,N_3954,N_5086);
nor U6486 (N_6486,N_4602,N_5789);
nand U6487 (N_6487,N_6055,N_3910);
and U6488 (N_6488,N_3775,N_3955);
or U6489 (N_6489,N_4084,N_3893);
nor U6490 (N_6490,N_5350,N_3564);
nand U6491 (N_6491,N_4963,N_3351);
nand U6492 (N_6492,N_4126,N_4061);
xor U6493 (N_6493,N_4450,N_3524);
nand U6494 (N_6494,N_4333,N_5430);
and U6495 (N_6495,N_5138,N_3324);
and U6496 (N_6496,N_5157,N_3481);
nor U6497 (N_6497,N_4175,N_4038);
xnor U6498 (N_6498,N_6058,N_5928);
nor U6499 (N_6499,N_3979,N_3322);
xnor U6500 (N_6500,N_4960,N_4984);
nand U6501 (N_6501,N_5279,N_3318);
nand U6502 (N_6502,N_5538,N_3505);
or U6503 (N_6503,N_5998,N_5878);
or U6504 (N_6504,N_5740,N_5306);
or U6505 (N_6505,N_5387,N_6075);
xnor U6506 (N_6506,N_3653,N_4074);
and U6507 (N_6507,N_4893,N_5134);
xor U6508 (N_6508,N_5870,N_5781);
nor U6509 (N_6509,N_6008,N_4703);
nand U6510 (N_6510,N_4078,N_6215);
or U6511 (N_6511,N_4925,N_4103);
xor U6512 (N_6512,N_5934,N_3516);
nand U6513 (N_6513,N_3726,N_5046);
nor U6514 (N_6514,N_4998,N_3155);
or U6515 (N_6515,N_4144,N_3892);
or U6516 (N_6516,N_4434,N_3392);
xor U6517 (N_6517,N_5400,N_5297);
and U6518 (N_6518,N_3430,N_5759);
xor U6519 (N_6519,N_5890,N_3610);
nand U6520 (N_6520,N_5534,N_4453);
or U6521 (N_6521,N_3805,N_3684);
nand U6522 (N_6522,N_5601,N_3870);
nor U6523 (N_6523,N_4586,N_4917);
xnor U6524 (N_6524,N_5111,N_4945);
or U6525 (N_6525,N_5687,N_5318);
or U6526 (N_6526,N_4504,N_3128);
nand U6527 (N_6527,N_5401,N_4759);
or U6528 (N_6528,N_5575,N_4009);
nand U6529 (N_6529,N_5807,N_3264);
and U6530 (N_6530,N_4916,N_3537);
nand U6531 (N_6531,N_4926,N_4077);
xor U6532 (N_6532,N_3642,N_3883);
or U6533 (N_6533,N_4405,N_4853);
xor U6534 (N_6534,N_4910,N_4562);
and U6535 (N_6535,N_5912,N_4110);
nor U6536 (N_6536,N_3221,N_4639);
nor U6537 (N_6537,N_4593,N_4957);
and U6538 (N_6538,N_5153,N_5753);
nand U6539 (N_6539,N_5048,N_3555);
nor U6540 (N_6540,N_3354,N_3387);
and U6541 (N_6541,N_3257,N_5612);
nor U6542 (N_6542,N_3635,N_4406);
nor U6543 (N_6543,N_3355,N_5218);
xor U6544 (N_6544,N_3297,N_4050);
and U6545 (N_6545,N_5706,N_6240);
xor U6546 (N_6546,N_6242,N_3808);
nand U6547 (N_6547,N_6031,N_5825);
xor U6548 (N_6548,N_3571,N_3968);
or U6549 (N_6549,N_4030,N_3443);
and U6550 (N_6550,N_5219,N_5602);
nand U6551 (N_6551,N_3482,N_5483);
nand U6552 (N_6552,N_5666,N_6176);
nor U6553 (N_6553,N_5006,N_5572);
and U6554 (N_6554,N_3498,N_5715);
xnor U6555 (N_6555,N_4436,N_5478);
and U6556 (N_6556,N_3329,N_4189);
and U6557 (N_6557,N_5253,N_4548);
xor U6558 (N_6558,N_5574,N_4717);
nand U6559 (N_6559,N_4010,N_4927);
xor U6560 (N_6560,N_3479,N_3607);
nor U6561 (N_6561,N_3521,N_3230);
and U6562 (N_6562,N_5627,N_5411);
xor U6563 (N_6563,N_5859,N_5019);
nand U6564 (N_6564,N_5013,N_5373);
and U6565 (N_6565,N_4261,N_5320);
or U6566 (N_6566,N_4155,N_3215);
and U6567 (N_6567,N_4266,N_3849);
nand U6568 (N_6568,N_5645,N_3287);
nand U6569 (N_6569,N_5388,N_4751);
or U6570 (N_6570,N_5007,N_4732);
xnor U6571 (N_6571,N_4756,N_3361);
nor U6572 (N_6572,N_3433,N_3791);
and U6573 (N_6573,N_5707,N_6106);
or U6574 (N_6574,N_5101,N_3178);
or U6575 (N_6575,N_5455,N_4806);
nand U6576 (N_6576,N_5557,N_3972);
or U6577 (N_6577,N_5254,N_5229);
nor U6578 (N_6578,N_4057,N_3236);
nor U6579 (N_6579,N_6092,N_4713);
xor U6580 (N_6580,N_6179,N_5830);
and U6581 (N_6581,N_3563,N_4792);
or U6582 (N_6582,N_4317,N_5366);
xnor U6583 (N_6583,N_3691,N_3734);
xor U6584 (N_6584,N_4157,N_3931);
or U6585 (N_6585,N_4617,N_4992);
nand U6586 (N_6586,N_5600,N_5577);
and U6587 (N_6587,N_4849,N_3621);
nor U6588 (N_6588,N_4489,N_3895);
or U6589 (N_6589,N_4559,N_3721);
xor U6590 (N_6590,N_5171,N_3706);
or U6591 (N_6591,N_5359,N_5778);
xnor U6592 (N_6592,N_3899,N_5438);
xnor U6593 (N_6593,N_4878,N_5780);
or U6594 (N_6594,N_4590,N_5755);
nand U6595 (N_6595,N_4544,N_4518);
nor U6596 (N_6596,N_3732,N_5603);
or U6597 (N_6597,N_4948,N_3658);
xnor U6598 (N_6598,N_4219,N_5569);
xnor U6599 (N_6599,N_3175,N_5614);
xnor U6600 (N_6600,N_5021,N_4576);
and U6601 (N_6601,N_5202,N_6226);
nand U6602 (N_6602,N_4066,N_4369);
or U6603 (N_6603,N_3941,N_5493);
or U6604 (N_6604,N_5814,N_4903);
nor U6605 (N_6605,N_3366,N_6018);
and U6606 (N_6606,N_4249,N_4677);
nor U6607 (N_6607,N_4336,N_3286);
and U6608 (N_6608,N_4832,N_3817);
and U6609 (N_6609,N_4746,N_3823);
or U6610 (N_6610,N_6159,N_3746);
xnor U6611 (N_6611,N_5408,N_4819);
xor U6612 (N_6612,N_4292,N_4300);
nand U6613 (N_6613,N_5642,N_4525);
or U6614 (N_6614,N_3325,N_3623);
or U6615 (N_6615,N_3675,N_3590);
or U6616 (N_6616,N_5892,N_3339);
or U6617 (N_6617,N_3364,N_3600);
or U6618 (N_6618,N_4018,N_5594);
and U6619 (N_6619,N_3868,N_6154);
xor U6620 (N_6620,N_4882,N_3971);
nand U6621 (N_6621,N_4896,N_3452);
xor U6622 (N_6622,N_3304,N_6109);
or U6623 (N_6623,N_5886,N_3223);
and U6624 (N_6624,N_5028,N_3826);
or U6625 (N_6625,N_6168,N_4966);
nor U6626 (N_6626,N_5804,N_5964);
nand U6627 (N_6627,N_6023,N_5421);
xnor U6628 (N_6628,N_3778,N_4465);
nand U6629 (N_6629,N_3163,N_4655);
nor U6630 (N_6630,N_4065,N_4173);
xnor U6631 (N_6631,N_3415,N_6097);
or U6632 (N_6632,N_5798,N_5996);
and U6633 (N_6633,N_4908,N_4784);
and U6634 (N_6634,N_5516,N_3695);
nor U6635 (N_6635,N_5850,N_3789);
nand U6636 (N_6636,N_5173,N_5987);
nor U6637 (N_6637,N_5567,N_3777);
xnor U6638 (N_6638,N_3834,N_5315);
xnor U6639 (N_6639,N_5922,N_5846);
nor U6640 (N_6640,N_4002,N_5014);
or U6641 (N_6641,N_3143,N_4835);
nand U6642 (N_6642,N_6206,N_3568);
nand U6643 (N_6643,N_4962,N_5980);
nor U6644 (N_6644,N_5795,N_5671);
and U6645 (N_6645,N_4625,N_6110);
and U6646 (N_6646,N_4384,N_6028);
nor U6647 (N_6647,N_3307,N_3784);
nor U6648 (N_6648,N_5875,N_4528);
and U6649 (N_6649,N_4459,N_5322);
nand U6650 (N_6650,N_5226,N_6088);
nand U6651 (N_6651,N_3501,N_3657);
nor U6652 (N_6652,N_4139,N_4698);
or U6653 (N_6653,N_3154,N_4274);
nand U6654 (N_6654,N_4725,N_3455);
and U6655 (N_6655,N_4134,N_4372);
nand U6656 (N_6656,N_4714,N_6165);
or U6657 (N_6657,N_4913,N_5901);
and U6658 (N_6658,N_5233,N_4930);
and U6659 (N_6659,N_3765,N_5523);
xor U6660 (N_6660,N_6232,N_3239);
and U6661 (N_6661,N_3168,N_3674);
or U6662 (N_6662,N_5917,N_4342);
nand U6663 (N_6663,N_6172,N_4679);
nor U6664 (N_6664,N_3923,N_3365);
nor U6665 (N_6665,N_3177,N_5240);
xor U6666 (N_6666,N_5722,N_6184);
xnor U6667 (N_6667,N_5842,N_3153);
and U6668 (N_6668,N_5295,N_5847);
nand U6669 (N_6669,N_5823,N_6025);
xnor U6670 (N_6670,N_5385,N_4332);
nand U6671 (N_6671,N_3240,N_3661);
nand U6672 (N_6672,N_3667,N_4973);
and U6673 (N_6673,N_5566,N_4673);
nand U6674 (N_6674,N_4990,N_5852);
nor U6675 (N_6675,N_5784,N_4255);
nand U6676 (N_6676,N_4529,N_6062);
nand U6677 (N_6677,N_5940,N_5881);
nor U6678 (N_6678,N_3447,N_3301);
nand U6679 (N_6679,N_4154,N_3908);
and U6680 (N_6680,N_5731,N_4217);
xor U6681 (N_6681,N_5460,N_5436);
nand U6682 (N_6682,N_3996,N_5674);
or U6683 (N_6683,N_6225,N_4165);
or U6684 (N_6684,N_3850,N_3829);
xnor U6685 (N_6685,N_4685,N_5345);
or U6686 (N_6686,N_6148,N_5296);
nand U6687 (N_6687,N_3188,N_3790);
nor U6688 (N_6688,N_3699,N_4809);
or U6689 (N_6689,N_3587,N_4204);
nor U6690 (N_6690,N_3937,N_3427);
nor U6691 (N_6691,N_4757,N_5333);
nand U6692 (N_6692,N_5225,N_4760);
nor U6693 (N_6693,N_5613,N_6020);
nand U6694 (N_6694,N_6006,N_5431);
nand U6695 (N_6695,N_5180,N_3529);
nor U6696 (N_6696,N_4512,N_3306);
nand U6697 (N_6697,N_3224,N_6208);
or U6698 (N_6698,N_6111,N_4825);
xnor U6699 (N_6699,N_5989,N_3827);
or U6700 (N_6700,N_3538,N_5889);
nand U6701 (N_6701,N_3891,N_3945);
xnor U6702 (N_6702,N_5456,N_6244);
xor U6703 (N_6703,N_5592,N_3201);
nor U6704 (N_6704,N_4833,N_3526);
nor U6705 (N_6705,N_5827,N_4880);
nor U6706 (N_6706,N_3442,N_3927);
nand U6707 (N_6707,N_4689,N_4580);
nand U6708 (N_6708,N_4624,N_3340);
xnor U6709 (N_6709,N_5285,N_5916);
xor U6710 (N_6710,N_4182,N_5503);
xor U6711 (N_6711,N_3491,N_4161);
nor U6712 (N_6712,N_5192,N_3876);
nor U6713 (N_6713,N_5412,N_5950);
or U6714 (N_6714,N_3338,N_3483);
or U6715 (N_6715,N_4538,N_5486);
or U6716 (N_6716,N_4517,N_5156);
or U6717 (N_6717,N_4808,N_4104);
and U6718 (N_6718,N_4147,N_4798);
nand U6719 (N_6719,N_5972,N_5787);
nand U6720 (N_6720,N_4813,N_3546);
nor U6721 (N_6721,N_6128,N_5962);
or U6722 (N_6722,N_5527,N_5507);
and U6723 (N_6723,N_4011,N_5949);
xor U6724 (N_6724,N_3251,N_6134);
or U6725 (N_6725,N_4389,N_5022);
xnor U6726 (N_6726,N_4535,N_3396);
nand U6727 (N_6727,N_3825,N_5774);
or U6728 (N_6728,N_5231,N_4592);
xor U6729 (N_6729,N_4318,N_4631);
xor U6730 (N_6730,N_4337,N_4376);
xor U6731 (N_6731,N_4199,N_4193);
and U6732 (N_6732,N_3648,N_3693);
nor U6733 (N_6733,N_5854,N_5667);
and U6734 (N_6734,N_3393,N_3872);
nand U6735 (N_6735,N_3901,N_4543);
nand U6736 (N_6736,N_3999,N_6038);
xnor U6737 (N_6737,N_3147,N_5047);
nor U6738 (N_6738,N_3394,N_5267);
or U6739 (N_6739,N_6121,N_4083);
nor U6740 (N_6740,N_3283,N_3559);
or U6741 (N_6741,N_3654,N_6175);
or U6742 (N_6742,N_5049,N_4470);
or U6743 (N_6743,N_4291,N_3137);
nand U6744 (N_6744,N_5628,N_5368);
xnor U6745 (N_6745,N_4191,N_4857);
nor U6746 (N_6746,N_5414,N_5150);
and U6747 (N_6747,N_4728,N_4171);
xor U6748 (N_6748,N_3853,N_4031);
nor U6749 (N_6749,N_3744,N_3636);
and U6750 (N_6750,N_5139,N_5002);
nand U6751 (N_6751,N_3461,N_5129);
and U6752 (N_6752,N_5407,N_4136);
or U6753 (N_6753,N_5657,N_5884);
xor U6754 (N_6754,N_5439,N_5265);
nor U6755 (N_6755,N_5383,N_4956);
and U6756 (N_6756,N_5147,N_6142);
nand U6757 (N_6757,N_3450,N_5094);
xor U6758 (N_6758,N_5948,N_3860);
and U6759 (N_6759,N_3608,N_4863);
nor U6760 (N_6760,N_4229,N_3664);
and U6761 (N_6761,N_3399,N_4401);
and U6762 (N_6762,N_3268,N_3947);
or U6763 (N_6763,N_3343,N_4539);
xor U6764 (N_6764,N_4386,N_4026);
and U6765 (N_6765,N_3182,N_3244);
and U6766 (N_6766,N_4840,N_3689);
nand U6767 (N_6767,N_5340,N_4186);
nand U6768 (N_6768,N_5801,N_3961);
xnor U6769 (N_6769,N_3500,N_3770);
nor U6770 (N_6770,N_3631,N_3209);
xnor U6771 (N_6771,N_4779,N_4107);
nand U6772 (N_6772,N_3754,N_4994);
and U6773 (N_6773,N_4430,N_3438);
xnor U6774 (N_6774,N_3878,N_4289);
and U6775 (N_6775,N_4563,N_4321);
nand U6776 (N_6776,N_4601,N_4661);
nand U6777 (N_6777,N_3577,N_3822);
and U6778 (N_6778,N_4817,N_3830);
or U6779 (N_6779,N_6241,N_4847);
or U6780 (N_6780,N_5480,N_4526);
or U6781 (N_6781,N_5777,N_5355);
nand U6782 (N_6782,N_4669,N_4411);
nand U6783 (N_6783,N_5286,N_6140);
or U6784 (N_6784,N_4017,N_4742);
or U6785 (N_6785,N_4810,N_5797);
nor U6786 (N_6786,N_3513,N_3719);
nand U6787 (N_6787,N_3806,N_4600);
xor U6788 (N_6788,N_3983,N_4745);
nor U6789 (N_6789,N_6194,N_5920);
or U6790 (N_6790,N_5897,N_5554);
or U6791 (N_6791,N_5951,N_5548);
and U6792 (N_6792,N_5939,N_5539);
or U6793 (N_6793,N_4063,N_4027);
or U6794 (N_6794,N_3909,N_5705);
or U6795 (N_6795,N_5437,N_5893);
xnor U6796 (N_6796,N_4020,N_5954);
xnor U6797 (N_6797,N_4095,N_3254);
xnor U6798 (N_6798,N_3400,N_5703);
or U6799 (N_6799,N_4972,N_5343);
and U6800 (N_6800,N_6169,N_3217);
nand U6801 (N_6801,N_5489,N_5163);
nor U6802 (N_6802,N_6201,N_3159);
or U6803 (N_6803,N_3484,N_3522);
and U6804 (N_6804,N_4415,N_4801);
nand U6805 (N_6805,N_4455,N_5032);
xnor U6806 (N_6806,N_3973,N_3476);
nor U6807 (N_6807,N_4928,N_3678);
nand U6808 (N_6808,N_5377,N_4803);
or U6809 (N_6809,N_4604,N_3701);
xnor U6810 (N_6810,N_4361,N_6210);
nor U6811 (N_6811,N_5498,N_5329);
and U6812 (N_6812,N_4034,N_3962);
nor U6813 (N_6813,N_4458,N_5690);
and U6814 (N_6814,N_4898,N_4672);
and U6815 (N_6815,N_5571,N_3552);
or U6816 (N_6816,N_3708,N_4842);
xor U6817 (N_6817,N_5301,N_5982);
nor U6818 (N_6818,N_3943,N_4348);
xnor U6819 (N_6819,N_6063,N_5026);
nand U6820 (N_6820,N_3267,N_5609);
nor U6821 (N_6821,N_5269,N_5128);
xnor U6822 (N_6822,N_3298,N_5003);
nand U6823 (N_6823,N_4286,N_4246);
nor U6824 (N_6824,N_3844,N_4722);
or U6825 (N_6825,N_4667,N_6135);
and U6826 (N_6826,N_5641,N_3843);
xnor U6827 (N_6827,N_4312,N_4382);
xor U6828 (N_6828,N_5517,N_5335);
and U6829 (N_6829,N_4942,N_3875);
and U6830 (N_6830,N_5033,N_5230);
or U6831 (N_6831,N_5079,N_4397);
or U6832 (N_6832,N_5905,N_3423);
xor U6833 (N_6833,N_3781,N_5625);
nand U6834 (N_6834,N_4552,N_4439);
nand U6835 (N_6835,N_5334,N_3629);
nand U6836 (N_6836,N_3633,N_5915);
and U6837 (N_6837,N_4651,N_5898);
or U6838 (N_6838,N_6214,N_6245);
and U6839 (N_6839,N_5452,N_5255);
and U6840 (N_6840,N_5702,N_4605);
nand U6841 (N_6841,N_3345,N_3253);
xor U6842 (N_6842,N_4986,N_4152);
xnor U6843 (N_6843,N_5541,N_3897);
and U6844 (N_6844,N_3210,N_6238);
nor U6845 (N_6845,N_4273,N_3326);
and U6846 (N_6846,N_6126,N_5692);
or U6847 (N_6847,N_3604,N_5971);
or U6848 (N_6848,N_4287,N_5813);
nand U6849 (N_6849,N_5038,N_4076);
or U6850 (N_6850,N_4752,N_4936);
xnor U6851 (N_6851,N_5970,N_5168);
or U6852 (N_6852,N_6205,N_5805);
or U6853 (N_6853,N_4632,N_5237);
and U6854 (N_6854,N_3651,N_4146);
nand U6855 (N_6855,N_3956,N_3262);
xor U6856 (N_6856,N_4119,N_4585);
xor U6857 (N_6857,N_4487,N_4499);
or U6858 (N_6858,N_4595,N_4619);
xnor U6859 (N_6859,N_4905,N_4185);
or U6860 (N_6860,N_5595,N_5053);
or U6861 (N_6861,N_6191,N_5351);
or U6862 (N_6862,N_3692,N_5165);
or U6863 (N_6863,N_5508,N_3353);
xnor U6864 (N_6864,N_5863,N_4448);
and U6865 (N_6865,N_4881,N_5494);
or U6866 (N_6866,N_4015,N_4895);
xor U6867 (N_6867,N_4125,N_3291);
or U6868 (N_6868,N_5389,N_4626);
xor U6869 (N_6869,N_5332,N_4500);
nand U6870 (N_6870,N_6141,N_4693);
nand U6871 (N_6871,N_5342,N_4894);
xor U6872 (N_6872,N_3402,N_5874);
or U6873 (N_6873,N_5471,N_5109);
xnor U6874 (N_6874,N_3238,N_5290);
nand U6875 (N_6875,N_5885,N_5542);
xnor U6876 (N_6876,N_4688,N_4758);
or U6877 (N_6877,N_4794,N_5367);
or U6878 (N_6878,N_4533,N_6227);
and U6879 (N_6879,N_5304,N_3683);
and U6880 (N_6880,N_3540,N_3728);
nor U6881 (N_6881,N_4920,N_3519);
xor U6882 (N_6882,N_4016,N_5891);
nor U6883 (N_6883,N_5141,N_5170);
nand U6884 (N_6884,N_4172,N_4976);
nor U6885 (N_6885,N_6024,N_4299);
xor U6886 (N_6886,N_5025,N_5535);
xor U6887 (N_6887,N_3589,N_4646);
nand U6888 (N_6888,N_5344,N_3184);
nand U6889 (N_6889,N_6173,N_5590);
nor U6890 (N_6890,N_4888,N_5440);
nand U6891 (N_6891,N_5585,N_3273);
nor U6892 (N_6892,N_3809,N_3771);
nor U6893 (N_6893,N_6181,N_4805);
nor U6894 (N_6894,N_6163,N_4723);
xor U6895 (N_6895,N_5442,N_4320);
or U6896 (N_6896,N_5636,N_3696);
nor U6897 (N_6897,N_5938,N_4524);
or U6898 (N_6898,N_4338,N_3711);
nor U6899 (N_6899,N_4236,N_3347);
nand U6900 (N_6900,N_5201,N_3385);
nor U6901 (N_6901,N_5700,N_5293);
and U6902 (N_6902,N_3824,N_4250);
and U6903 (N_6903,N_4368,N_3200);
or U6904 (N_6904,N_3681,N_5008);
nand U6905 (N_6905,N_5429,N_3890);
and U6906 (N_6906,N_5137,N_3193);
and U6907 (N_6907,N_5130,N_5070);
or U6908 (N_6908,N_3641,N_4028);
and U6909 (N_6909,N_5509,N_4059);
and U6910 (N_6910,N_4776,N_5287);
or U6911 (N_6911,N_3518,N_4051);
nand U6912 (N_6912,N_5637,N_5502);
nand U6913 (N_6913,N_6107,N_3930);
or U6914 (N_6914,N_4939,N_3389);
xnor U6915 (N_6915,N_3406,N_6108);
nor U6916 (N_6916,N_3742,N_5462);
xnor U6917 (N_6917,N_3852,N_3950);
nor U6918 (N_6918,N_6138,N_3807);
xor U6919 (N_6919,N_3309,N_3618);
and U6920 (N_6920,N_5646,N_6187);
xnor U6921 (N_6921,N_4864,N_5762);
or U6922 (N_6922,N_4417,N_5589);
or U6923 (N_6923,N_3851,N_5675);
nand U6924 (N_6924,N_4143,N_4753);
nor U6925 (N_6925,N_5764,N_5190);
or U6926 (N_6926,N_3299,N_3871);
or U6927 (N_6927,N_5010,N_5779);
and U6928 (N_6928,N_4392,N_3186);
nand U6929 (N_6929,N_5757,N_6219);
or U6930 (N_6930,N_5903,N_5708);
xor U6931 (N_6931,N_3456,N_5867);
nor U6932 (N_6932,N_3572,N_3547);
xnor U6933 (N_6933,N_3214,N_4309);
or U6934 (N_6934,N_6022,N_4718);
nand U6935 (N_6935,N_5511,N_6017);
and U6936 (N_6936,N_4834,N_5606);
or U6937 (N_6937,N_5417,N_3388);
and U6938 (N_6938,N_5268,N_3639);
nor U6939 (N_6939,N_3939,N_5699);
nand U6940 (N_6940,N_5744,N_6000);
nand U6941 (N_6941,N_3232,N_4174);
xnor U6942 (N_6942,N_5249,N_4919);
or U6943 (N_6943,N_4964,N_4709);
or U6944 (N_6944,N_4429,N_5685);
xnor U6945 (N_6945,N_3785,N_3376);
and U6946 (N_6946,N_4974,N_5212);
xor U6947 (N_6947,N_3126,N_4164);
xor U6948 (N_6948,N_3391,N_4985);
or U6949 (N_6949,N_4506,N_5145);
nand U6950 (N_6950,N_3205,N_3420);
nor U6951 (N_6951,N_4462,N_5746);
xnor U6952 (N_6952,N_4213,N_4304);
and U6953 (N_6953,N_3864,N_3987);
nor U6954 (N_6954,N_5993,N_5172);
nor U6955 (N_6955,N_4686,N_6101);
nand U6956 (N_6956,N_5005,N_5448);
or U6957 (N_6957,N_6098,N_3798);
nor U6958 (N_6958,N_4464,N_4159);
xnor U6959 (N_6959,N_5742,N_3609);
nand U6960 (N_6960,N_4633,N_5203);
nor U6961 (N_6961,N_4668,N_4629);
xnor U6962 (N_6962,N_4692,N_5467);
nand U6963 (N_6963,N_4350,N_3981);
or U6964 (N_6964,N_5821,N_5406);
nor U6965 (N_6965,N_5035,N_4510);
and U6966 (N_6966,N_5840,N_5069);
or U6967 (N_6967,N_5151,N_5623);
or U6968 (N_6968,N_4989,N_4427);
nand U6969 (N_6969,N_3740,N_5182);
or U6970 (N_6970,N_4087,N_4589);
and U6971 (N_6971,N_3670,N_5808);
nand U6972 (N_6972,N_3289,N_4570);
xnor U6973 (N_6973,N_4935,N_6056);
and U6974 (N_6974,N_6167,N_3360);
or U6975 (N_6975,N_4380,N_5245);
and U6976 (N_6976,N_3592,N_5693);
and U6977 (N_6977,N_3233,N_3774);
nand U6978 (N_6978,N_5953,N_4612);
nand U6979 (N_6979,N_5904,N_5824);
xnor U6980 (N_6980,N_3471,N_4740);
xor U6981 (N_6981,N_5105,N_5327);
and U6982 (N_6982,N_5451,N_6192);
nand U6983 (N_6983,N_5149,N_3714);
nor U6984 (N_6984,N_6202,N_5520);
or U6985 (N_6985,N_4223,N_4356);
xnor U6986 (N_6986,N_4263,N_5961);
nor U6987 (N_6987,N_4488,N_4636);
nand U6988 (N_6988,N_5361,N_4682);
xor U6989 (N_6989,N_3204,N_5937);
nand U6990 (N_6990,N_5524,N_6034);
nor U6991 (N_6991,N_3548,N_5247);
xnor U6992 (N_6992,N_6166,N_4005);
or U6993 (N_6993,N_3926,N_6103);
nor U6994 (N_6994,N_5266,N_6048);
or U6995 (N_6995,N_4599,N_5294);
and U6996 (N_6996,N_4541,N_6002);
and U6997 (N_6997,N_4269,N_4620);
xnor U6998 (N_6998,N_4220,N_4075);
and U6999 (N_6999,N_4100,N_4256);
nand U7000 (N_7000,N_3562,N_3328);
and U7001 (N_7001,N_4271,N_6130);
nand U7002 (N_7002,N_4088,N_5766);
nor U7003 (N_7003,N_5694,N_5923);
xor U7004 (N_7004,N_5732,N_6004);
nand U7005 (N_7005,N_4652,N_5311);
and U7006 (N_7006,N_4298,N_5536);
xnor U7007 (N_7007,N_3317,N_6041);
xor U7008 (N_7008,N_6072,N_4637);
or U7009 (N_7009,N_4816,N_3611);
xor U7010 (N_7010,N_5465,N_3869);
nand U7011 (N_7011,N_4106,N_5472);
or U7012 (N_7012,N_4226,N_5481);
xnor U7013 (N_7013,N_3917,N_3649);
xnor U7014 (N_7014,N_6012,N_4440);
xnor U7015 (N_7015,N_3982,N_5113);
or U7016 (N_7016,N_5174,N_3144);
xor U7017 (N_7017,N_3373,N_5449);
nor U7018 (N_7018,N_5341,N_5745);
xor U7019 (N_7019,N_4642,N_5257);
nor U7020 (N_7020,N_6164,N_3372);
or U7021 (N_7021,N_5073,N_5942);
nor U7022 (N_7022,N_4242,N_3226);
nand U7023 (N_7023,N_3462,N_6127);
xor U7024 (N_7024,N_3398,N_4366);
xnor U7025 (N_7025,N_3139,N_4536);
nor U7026 (N_7026,N_3127,N_4259);
nand U7027 (N_7027,N_5356,N_6112);
or U7028 (N_7028,N_5252,N_5000);
or U7029 (N_7029,N_5833,N_5424);
nand U7030 (N_7030,N_4841,N_4741);
nand U7031 (N_7031,N_4184,N_6049);
or U7032 (N_7032,N_6132,N_3880);
and U7033 (N_7033,N_5222,N_4616);
nand U7034 (N_7034,N_3531,N_3348);
and U7035 (N_7035,N_5464,N_5580);
xor U7036 (N_7036,N_5721,N_5596);
nor U7037 (N_7037,N_5506,N_5347);
or U7038 (N_7038,N_3736,N_5475);
xnor U7039 (N_7039,N_3576,N_4132);
nand U7040 (N_7040,N_6077,N_4551);
or U7041 (N_7041,N_4491,N_4253);
nor U7042 (N_7042,N_5988,N_4793);
nand U7043 (N_7043,N_4877,N_5913);
xor U7044 (N_7044,N_5581,N_4764);
or U7045 (N_7045,N_4979,N_3603);
and U7046 (N_7046,N_5115,N_5453);
or U7047 (N_7047,N_4306,N_3352);
nor U7048 (N_7048,N_5419,N_5738);
and U7049 (N_7049,N_5793,N_3704);
nand U7050 (N_7050,N_5810,N_5630);
and U7051 (N_7051,N_3756,N_3677);
nor U7052 (N_7052,N_3208,N_4296);
nand U7053 (N_7053,N_4780,N_5712);
and U7054 (N_7054,N_5120,N_5836);
or U7055 (N_7055,N_3409,N_3832);
nand U7056 (N_7056,N_4367,N_4666);
nand U7057 (N_7057,N_5631,N_4128);
nor U7058 (N_7058,N_4195,N_5369);
nor U7059 (N_7059,N_3295,N_3225);
and U7060 (N_7060,N_3762,N_5080);
nand U7061 (N_7061,N_5899,N_5052);
or U7062 (N_7062,N_3162,N_3989);
nand U7063 (N_7063,N_3248,N_6178);
xnor U7064 (N_7064,N_4225,N_5588);
and U7065 (N_7065,N_5256,N_3718);
nand U7066 (N_7066,N_5043,N_5761);
nand U7067 (N_7067,N_3646,N_5415);
nand U7068 (N_7068,N_5871,N_5326);
xor U7069 (N_7069,N_4360,N_5118);
nand U7070 (N_7070,N_5095,N_6084);
or U7071 (N_7071,N_4695,N_3783);
xor U7072 (N_7072,N_4643,N_4444);
xor U7073 (N_7073,N_5660,N_5958);
or U7074 (N_7074,N_3320,N_3924);
and U7075 (N_7075,N_3637,N_3969);
and U7076 (N_7076,N_3473,N_4177);
nor U7077 (N_7077,N_4471,N_4763);
and U7078 (N_7078,N_4943,N_3492);
or U7079 (N_7079,N_4521,N_4212);
xnor U7080 (N_7080,N_3349,N_4141);
and U7081 (N_7081,N_5716,N_4054);
or U7082 (N_7082,N_5635,N_3588);
nor U7083 (N_7083,N_5164,N_4301);
nor U7084 (N_7084,N_4564,N_5783);
and U7085 (N_7085,N_5023,N_3992);
or U7086 (N_7086,N_4283,N_3769);
and U7087 (N_7087,N_3242,N_3614);
or U7088 (N_7088,N_3183,N_3913);
nand U7089 (N_7089,N_3414,N_4352);
xor U7090 (N_7090,N_3679,N_3723);
xor U7091 (N_7091,N_4706,N_3581);
nor U7092 (N_7092,N_6050,N_5189);
nor U7093 (N_7093,N_4004,N_4767);
and U7094 (N_7094,N_5457,N_4999);
or U7095 (N_7095,N_5059,N_5098);
or U7096 (N_7096,N_5215,N_6223);
nand U7097 (N_7097,N_5860,N_5470);
and U7098 (N_7098,N_6129,N_4008);
and U7099 (N_7099,N_4120,N_5375);
xnor U7100 (N_7100,N_5127,N_4665);
and U7101 (N_7101,N_6221,N_6033);
and U7102 (N_7102,N_4892,N_5330);
nand U7103 (N_7103,N_4824,N_5747);
or U7104 (N_7104,N_3902,N_5058);
and U7105 (N_7105,N_3279,N_4093);
nand U7106 (N_7106,N_3496,N_5491);
and U7107 (N_7107,N_3862,N_4314);
xor U7108 (N_7108,N_4573,N_5364);
nand U7109 (N_7109,N_5274,N_4876);
nor U7110 (N_7110,N_5914,N_6015);
nor U7111 (N_7111,N_3227,N_4684);
nor U7112 (N_7112,N_5321,N_5586);
xor U7113 (N_7113,N_5545,N_3911);
xnor U7114 (N_7114,N_4923,N_3918);
and U7115 (N_7115,N_3314,N_5124);
and U7116 (N_7116,N_5446,N_5428);
and U7117 (N_7117,N_5261,N_3197);
xor U7118 (N_7118,N_4469,N_3866);
nor U7119 (N_7119,N_3469,N_3953);
xor U7120 (N_7120,N_5697,N_4608);
or U7121 (N_7121,N_3551,N_6069);
xnor U7122 (N_7122,N_3656,N_5015);
or U7123 (N_7123,N_3411,N_5936);
or U7124 (N_7124,N_4334,N_4775);
and U7125 (N_7125,N_5090,N_3228);
nor U7126 (N_7126,N_5790,N_3963);
xor U7127 (N_7127,N_5894,N_5244);
nor U7128 (N_7128,N_5643,N_4135);
nand U7129 (N_7129,N_3199,N_3487);
xnor U7130 (N_7130,N_4568,N_6087);
nor U7131 (N_7131,N_5071,N_3506);
and U7132 (N_7132,N_6122,N_3288);
xor U7133 (N_7133,N_4477,N_5841);
xor U7134 (N_7134,N_5305,N_4085);
or U7135 (N_7135,N_5116,N_4121);
nor U7136 (N_7136,N_4911,N_5205);
nor U7137 (N_7137,N_3764,N_3440);
and U7138 (N_7138,N_5930,N_5981);
xnor U7139 (N_7139,N_4850,N_5051);
nor U7140 (N_7140,N_4247,N_4766);
or U7141 (N_7141,N_3619,N_3207);
and U7142 (N_7142,N_4216,N_3445);
nand U7143 (N_7143,N_5868,N_5220);
and U7144 (N_7144,N_3220,N_4922);
xnor U7145 (N_7145,N_4519,N_5162);
and U7146 (N_7146,N_4113,N_3994);
nor U7147 (N_7147,N_3271,N_5123);
xnor U7148 (N_7148,N_5837,N_3964);
nand U7149 (N_7149,N_4540,N_5027);
nand U7150 (N_7150,N_4330,N_5188);
nor U7151 (N_7151,N_3544,N_5662);
or U7152 (N_7152,N_4391,N_3194);
nand U7153 (N_7153,N_5733,N_3294);
nor U7154 (N_7154,N_3206,N_5661);
nand U7155 (N_7155,N_5963,N_5075);
nor U7156 (N_7156,N_3237,N_4511);
and U7157 (N_7157,N_4211,N_3460);
and U7158 (N_7158,N_5647,N_4435);
nand U7159 (N_7159,N_4452,N_4239);
nor U7160 (N_7160,N_5504,N_5062);
nor U7161 (N_7161,N_4426,N_3138);
or U7162 (N_7162,N_5142,N_4351);
xor U7163 (N_7163,N_5317,N_5834);
xnor U7164 (N_7164,N_3715,N_5018);
nor U7165 (N_7165,N_4566,N_5410);
xnor U7166 (N_7166,N_4048,N_4820);
xor U7167 (N_7167,N_5040,N_5477);
nand U7168 (N_7168,N_4578,N_3858);
nor U7169 (N_7169,N_6030,N_4033);
nor U7170 (N_7170,N_5397,N_3965);
and U7171 (N_7171,N_3310,N_4613);
nand U7172 (N_7172,N_3191,N_4522);
xnor U7173 (N_7173,N_5758,N_3266);
xnor U7174 (N_7174,N_3554,N_4325);
and U7175 (N_7175,N_6082,N_4443);
nor U7176 (N_7176,N_4307,N_5578);
and U7177 (N_7177,N_4080,N_4498);
or U7178 (N_7178,N_3408,N_5735);
and U7179 (N_7179,N_5820,N_5664);
nor U7180 (N_7180,N_3601,N_5055);
and U7181 (N_7181,N_3698,N_3842);
nor U7182 (N_7182,N_6204,N_5782);
nor U7183 (N_7183,N_5298,N_4248);
or U7184 (N_7184,N_3370,N_5653);
xnor U7185 (N_7185,N_4886,N_3599);
nor U7186 (N_7186,N_4374,N_4316);
nor U7187 (N_7187,N_4163,N_5944);
or U7188 (N_7188,N_4019,N_4822);
nor U7189 (N_7189,N_4040,N_4305);
or U7190 (N_7190,N_4441,N_5198);
xnor U7191 (N_7191,N_5492,N_4133);
nand U7192 (N_7192,N_4858,N_5067);
xor U7193 (N_7193,N_4370,N_6213);
or U7194 (N_7194,N_4650,N_4782);
nor U7195 (N_7195,N_3311,N_3371);
xor U7196 (N_7196,N_4388,N_3375);
xnor U7197 (N_7197,N_3231,N_5303);
nand U7198 (N_7198,N_5422,N_6185);
or U7199 (N_7199,N_4837,N_4983);
and U7200 (N_7200,N_5288,N_5818);
nor U7201 (N_7201,N_4556,N_5082);
nor U7202 (N_7202,N_6124,N_4071);
or U7203 (N_7203,N_5526,N_5089);
or U7204 (N_7204,N_4587,N_3146);
and U7205 (N_7205,N_6203,N_4331);
nor U7206 (N_7206,N_3877,N_4735);
xnor U7207 (N_7207,N_4032,N_4170);
and U7208 (N_7208,N_5313,N_4007);
xnor U7209 (N_7209,N_5945,N_6234);
xor U7210 (N_7210,N_6239,N_5490);
nand U7211 (N_7211,N_3261,N_3431);
xor U7212 (N_7212,N_5346,N_3750);
nor U7213 (N_7213,N_4224,N_4596);
and U7214 (N_7214,N_5270,N_3904);
nor U7215 (N_7215,N_4043,N_3134);
and U7216 (N_7216,N_4201,N_5599);
or U7217 (N_7217,N_3255,N_3612);
and U7218 (N_7218,N_3125,N_3472);
and U7219 (N_7219,N_5084,N_5488);
or U7220 (N_7220,N_4501,N_5425);
or U7221 (N_7221,N_5822,N_4747);
nand U7222 (N_7222,N_5995,N_3258);
xnor U7223 (N_7223,N_5066,N_4571);
nor U7224 (N_7224,N_3763,N_3467);
or U7225 (N_7225,N_6212,N_4474);
xnor U7226 (N_7226,N_4821,N_6174);
and U7227 (N_7227,N_5432,N_4875);
nand U7228 (N_7228,N_3495,N_5404);
nand U7229 (N_7229,N_5544,N_5078);
nor U7230 (N_7230,N_3410,N_5103);
xnor U7231 (N_7231,N_3672,N_3948);
nor U7232 (N_7232,N_3229,N_4687);
xor U7233 (N_7233,N_3613,N_5324);
and U7234 (N_7234,N_4508,N_6153);
xnor U7235 (N_7235,N_4257,N_6230);
nand U7236 (N_7236,N_4284,N_5734);
and U7237 (N_7237,N_4581,N_5968);
or U7238 (N_7238,N_6222,N_4978);
nor U7239 (N_7239,N_3799,N_4082);
and U7240 (N_7240,N_5887,N_4365);
xor U7241 (N_7241,N_5447,N_5328);
xor U7242 (N_7242,N_4799,N_5372);
nor U7243 (N_7243,N_4476,N_5319);
nor U7244 (N_7244,N_4987,N_3222);
and U7245 (N_7245,N_4614,N_4988);
and U7246 (N_7246,N_4294,N_5131);
xnor U7247 (N_7247,N_3720,N_6026);
and U7248 (N_7248,N_6066,N_5546);
nand U7249 (N_7249,N_5770,N_3527);
and U7250 (N_7250,N_5029,N_6079);
nor U7251 (N_7251,N_3474,N_3573);
xor U7252 (N_7252,N_6158,N_5004);
xor U7253 (N_7253,N_4055,N_3757);
nand U7254 (N_7254,N_4449,N_3865);
nand U7255 (N_7255,N_4938,N_3802);
nor U7256 (N_7256,N_3847,N_3574);
and U7257 (N_7257,N_4188,N_5806);
and U7258 (N_7258,N_4494,N_4327);
nor U7259 (N_7259,N_5391,N_6248);
nor U7260 (N_7260,N_5974,N_4790);
or U7261 (N_7261,N_5973,N_4281);
or U7262 (N_7262,N_5772,N_3626);
nor U7263 (N_7263,N_5024,N_4379);
xor U7264 (N_7264,N_6151,N_4451);
nor U7265 (N_7265,N_3510,N_5607);
xor U7266 (N_7266,N_3386,N_3887);
nor U7267 (N_7267,N_4495,N_5519);
xor U7268 (N_7268,N_5338,N_5112);
nor U7269 (N_7269,N_3136,N_5463);
nor U7270 (N_7270,N_5353,N_5074);
and U7271 (N_7271,N_5076,N_4807);
nor U7272 (N_7272,N_4293,N_4733);
and U7273 (N_7273,N_5907,N_6125);
and U7274 (N_7274,N_4148,N_4959);
nor U7275 (N_7275,N_4149,N_4549);
or U7276 (N_7276,N_5696,N_4618);
or U7277 (N_7277,N_4268,N_5633);
or U7278 (N_7278,N_4377,N_5769);
or U7279 (N_7279,N_3401,N_4073);
xnor U7280 (N_7280,N_6037,N_5855);
or U7281 (N_7281,N_3975,N_3454);
xnor U7282 (N_7282,N_3906,N_5275);
xnor U7283 (N_7283,N_4319,N_4042);
or U7284 (N_7284,N_6090,N_5882);
or U7285 (N_7285,N_4218,N_4690);
nor U7286 (N_7286,N_5547,N_5496);
xnor U7287 (N_7287,N_3952,N_5380);
nor U7288 (N_7288,N_6243,N_5178);
xnor U7289 (N_7289,N_4865,N_5659);
and U7290 (N_7290,N_3697,N_4915);
or U7291 (N_7291,N_4781,N_5289);
and U7292 (N_7292,N_6247,N_4657);
xor U7293 (N_7293,N_5358,N_5969);
nor U7294 (N_7294,N_5618,N_3660);
nand U7295 (N_7295,N_4044,N_6019);
xor U7296 (N_7296,N_4860,N_5644);
and U7297 (N_7297,N_3747,N_5100);
xnor U7298 (N_7298,N_4262,N_3786);
or U7299 (N_7299,N_4955,N_3247);
xor U7300 (N_7300,N_5668,N_3739);
xnor U7301 (N_7301,N_3390,N_5927);
xnor U7302 (N_7302,N_4280,N_3863);
and U7303 (N_7303,N_3700,N_3426);
nor U7304 (N_7304,N_4413,N_4240);
xor U7305 (N_7305,N_3845,N_5371);
nand U7306 (N_7306,N_5750,N_5832);
nand U7307 (N_7307,N_3933,N_5728);
nor U7308 (N_7308,N_4447,N_3412);
and U7309 (N_7309,N_3914,N_3246);
and U7310 (N_7310,N_3569,N_5484);
xor U7311 (N_7311,N_5900,N_3940);
or U7312 (N_7312,N_5420,N_4232);
and U7313 (N_7313,N_4192,N_5061);
xor U7314 (N_7314,N_3333,N_5565);
nor U7315 (N_7315,N_5196,N_5967);
nor U7316 (N_7316,N_5276,N_5551);
or U7317 (N_7317,N_3470,N_3335);
or U7318 (N_7318,N_4739,N_5576);
xnor U7319 (N_7319,N_4934,N_3313);
or U7320 (N_7320,N_6073,N_3437);
nand U7321 (N_7321,N_4068,N_5416);
nand U7322 (N_7322,N_6091,N_3724);
and U7323 (N_7323,N_6147,N_3760);
or U7324 (N_7324,N_5179,N_5800);
or U7325 (N_7325,N_4285,N_5177);
xnor U7326 (N_7326,N_4953,N_4634);
or U7327 (N_7327,N_4137,N_5906);
or U7328 (N_7328,N_5186,N_5246);
or U7329 (N_7329,N_4344,N_3819);
and U7330 (N_7330,N_3748,N_3422);
nor U7331 (N_7331,N_4140,N_4609);
nor U7332 (N_7332,N_4944,N_4575);
nand U7333 (N_7333,N_3533,N_4569);
and U7334 (N_7334,N_4313,N_5924);
nor U7335 (N_7335,N_6131,N_5042);
nor U7336 (N_7336,N_3929,N_5065);
and U7337 (N_7337,N_3160,N_4403);
nor U7338 (N_7338,N_4674,N_6043);
nand U7339 (N_7339,N_5250,N_6104);
and U7340 (N_7340,N_3729,N_6086);
xor U7341 (N_7341,N_4502,N_5610);
or U7342 (N_7342,N_5977,N_3932);
nand U7343 (N_7343,N_3650,N_5921);
or U7344 (N_7344,N_5864,N_4970);
nor U7345 (N_7345,N_5495,N_3625);
nand U7346 (N_7346,N_5771,N_5354);
nand U7347 (N_7347,N_4902,N_3767);
xnor U7348 (N_7348,N_4341,N_5650);
xnor U7349 (N_7349,N_5272,N_3995);
or U7350 (N_7350,N_5865,N_5719);
nor U7351 (N_7351,N_5991,N_5092);
nand U7352 (N_7352,N_5862,N_5251);
and U7353 (N_7353,N_5088,N_3170);
xor U7354 (N_7354,N_4981,N_3712);
or U7355 (N_7355,N_5932,N_5960);
and U7356 (N_7356,N_3350,N_4736);
xor U7357 (N_7357,N_5673,N_4130);
nor U7358 (N_7358,N_4630,N_4811);
nor U7359 (N_7359,N_3813,N_4362);
xor U7360 (N_7360,N_4467,N_4052);
and U7361 (N_7361,N_6042,N_3417);
nand U7362 (N_7362,N_3216,N_3957);
and U7363 (N_7363,N_5175,N_5054);
nand U7364 (N_7364,N_5243,N_5160);
and U7365 (N_7365,N_5009,N_3584);
or U7366 (N_7366,N_3586,N_5861);
nand U7367 (N_7367,N_4867,N_4520);
or U7368 (N_7368,N_3582,N_5816);
nor U7369 (N_7369,N_3151,N_5185);
nor U7370 (N_7370,N_6217,N_3545);
nor U7371 (N_7371,N_3713,N_3171);
or U7372 (N_7372,N_5979,N_3512);
and U7373 (N_7373,N_3703,N_4053);
or U7374 (N_7374,N_4092,N_4475);
nand U7375 (N_7375,N_3812,N_5144);
and U7376 (N_7376,N_4202,N_6133);
and U7377 (N_7377,N_5656,N_5760);
and U7378 (N_7378,N_5473,N_6105);
nor U7379 (N_7379,N_4203,N_5228);
and U7380 (N_7380,N_5639,N_5264);
xor U7381 (N_7381,N_3733,N_5126);
or U7382 (N_7382,N_4021,N_3330);
nand U7383 (N_7383,N_3441,N_3377);
and U7384 (N_7384,N_3549,N_4390);
and U7385 (N_7385,N_5213,N_5931);
nor U7386 (N_7386,N_3425,N_5223);
or U7387 (N_7387,N_4707,N_3308);
nor U7388 (N_7388,N_4696,N_5564);
or U7389 (N_7389,N_3413,N_5698);
nor U7390 (N_7390,N_4969,N_5560);
or U7391 (N_7391,N_3935,N_4178);
and U7392 (N_7392,N_5087,N_4683);
or U7393 (N_7393,N_4012,N_4791);
nor U7394 (N_7394,N_3886,N_3583);
and U7395 (N_7395,N_4486,N_3158);
nor U7396 (N_7396,N_4339,N_4094);
and U7397 (N_7397,N_3779,N_3630);
and U7398 (N_7398,N_5785,N_3815);
and U7399 (N_7399,N_4355,N_4830);
xor U7400 (N_7400,N_5041,N_3673);
xor U7401 (N_7401,N_5512,N_6152);
nor U7402 (N_7402,N_4421,N_5091);
xnor U7403 (N_7403,N_4190,N_3397);
xnor U7404 (N_7404,N_3717,N_4710);
nor U7405 (N_7405,N_4480,N_5395);
nand U7406 (N_7406,N_4221,N_6081);
and U7407 (N_7407,N_4831,N_3640);
nand U7408 (N_7408,N_5672,N_5194);
or U7409 (N_7409,N_5902,N_4641);
nor U7410 (N_7410,N_5445,N_4514);
nand U7411 (N_7411,N_4324,N_4479);
nand U7412 (N_7412,N_3676,N_6170);
and U7413 (N_7413,N_5302,N_3384);
and U7414 (N_7414,N_4238,N_6200);
nor U7415 (N_7415,N_5649,N_4105);
or U7416 (N_7416,N_4425,N_4006);
and U7417 (N_7417,N_3429,N_4771);
nand U7418 (N_7418,N_4699,N_4607);
nor U7419 (N_7419,N_5336,N_3888);
nor U7420 (N_7420,N_4345,N_5278);
or U7421 (N_7421,N_4797,N_4275);
xor U7422 (N_7422,N_5809,N_3788);
and U7423 (N_7423,N_5314,N_3543);
or U7424 (N_7424,N_5197,N_6102);
and U7425 (N_7425,N_3727,N_4497);
xor U7426 (N_7426,N_3743,N_4000);
xor U7427 (N_7427,N_4492,N_4743);
xor U7428 (N_7428,N_3234,N_4176);
and U7429 (N_7429,N_4335,N_5125);
nand U7430 (N_7430,N_4868,N_3530);
xnor U7431 (N_7431,N_4929,N_4879);
and U7432 (N_7432,N_4111,N_4565);
nor U7433 (N_7433,N_5352,N_4231);
and U7434 (N_7434,N_3383,N_4912);
nor U7435 (N_7435,N_3382,N_6186);
nand U7436 (N_7436,N_3285,N_5239);
or U7437 (N_7437,N_4523,N_3966);
or U7438 (N_7438,N_4278,N_3203);
nand U7439 (N_7439,N_4049,N_4907);
or U7440 (N_7440,N_3277,N_4621);
nand U7441 (N_7441,N_4424,N_4727);
or U7442 (N_7442,N_4937,N_5763);
and U7443 (N_7443,N_5638,N_4422);
or U7444 (N_7444,N_4788,N_5382);
or U7445 (N_7445,N_4023,N_3967);
xnor U7446 (N_7446,N_4615,N_4836);
nand U7447 (N_7447,N_4363,N_5605);
and U7448 (N_7448,N_4064,N_3766);
xor U7449 (N_7449,N_3535,N_4322);
or U7450 (N_7450,N_4941,N_4951);
xnor U7451 (N_7451,N_3854,N_5532);
or U7452 (N_7452,N_6236,N_3922);
nor U7453 (N_7453,N_4949,N_5096);
xnor U7454 (N_7454,N_3362,N_3480);
nand U7455 (N_7455,N_4230,N_4676);
nor U7456 (N_7456,N_3374,N_4950);
xor U7457 (N_7457,N_5561,N_5730);
xor U7458 (N_7458,N_4160,N_4481);
and U7459 (N_7459,N_4597,N_5655);
xor U7460 (N_7460,N_3731,N_5695);
nand U7461 (N_7461,N_3566,N_4181);
xor U7462 (N_7462,N_5282,N_4546);
nor U7463 (N_7463,N_5985,N_3833);
or U7464 (N_7464,N_3620,N_3682);
xor U7465 (N_7465,N_4258,N_3991);
or U7466 (N_7466,N_6211,N_3131);
xor U7467 (N_7467,N_6099,N_5877);
nand U7468 (N_7468,N_6157,N_4648);
nor U7469 (N_7469,N_5665,N_3133);
nand U7470 (N_7470,N_4947,N_3502);
nand U7471 (N_7471,N_3959,N_5568);
and U7472 (N_7472,N_5555,N_5396);
nor U7473 (N_7473,N_3787,N_3457);
xor U7474 (N_7474,N_4162,N_4196);
and U7475 (N_7475,N_3702,N_4968);
or U7476 (N_7476,N_4730,N_6045);
nand U7477 (N_7477,N_5515,N_3632);
nor U7478 (N_7478,N_3342,N_5992);
and U7479 (N_7479,N_4461,N_5152);
and U7480 (N_7480,N_5513,N_4251);
xor U7481 (N_7481,N_3439,N_3135);
xnor U7482 (N_7482,N_4117,N_3446);
or U7483 (N_7483,N_3315,N_6044);
and U7484 (N_7484,N_5957,N_5469);
and U7485 (N_7485,N_5399,N_4980);
nor U7486 (N_7486,N_4131,N_3565);
and U7487 (N_7487,N_3585,N_5102);
and U7488 (N_7488,N_5873,N_3776);
and U7489 (N_7489,N_5768,N_5786);
nand U7490 (N_7490,N_4472,N_4557);
nor U7491 (N_7491,N_5117,N_4635);
xor U7492 (N_7492,N_6032,N_3745);
nor U7493 (N_7493,N_6047,N_3278);
nor U7494 (N_7494,N_3970,N_3459);
nor U7495 (N_7495,N_3616,N_3984);
xnor U7496 (N_7496,N_3958,N_4123);
and U7497 (N_7497,N_5819,N_5584);
or U7498 (N_7498,N_4663,N_5811);
nand U7499 (N_7499,N_5121,N_4537);
or U7500 (N_7500,N_3432,N_6021);
and U7501 (N_7501,N_5384,N_4395);
nand U7502 (N_7502,N_3164,N_3243);
nor U7503 (N_7503,N_6180,N_4228);
or U7504 (N_7504,N_3998,N_6249);
xnor U7505 (N_7505,N_4530,N_5258);
xnor U7506 (N_7506,N_4478,N_4885);
xor U7507 (N_7507,N_5169,N_3580);
nor U7508 (N_7508,N_6233,N_5717);
xor U7509 (N_7509,N_3380,N_5844);
nand U7510 (N_7510,N_5357,N_4826);
nand U7511 (N_7511,N_3508,N_3615);
or U7512 (N_7512,N_3174,N_5688);
nor U7513 (N_7513,N_4288,N_4383);
or U7514 (N_7514,N_5316,N_6150);
xnor U7515 (N_7515,N_4638,N_5349);
nor U7516 (N_7516,N_5872,N_5799);
nor U7517 (N_7517,N_4897,N_3960);
xnor U7518 (N_7518,N_3356,N_4777);
nor U7519 (N_7519,N_3140,N_3558);
nand U7520 (N_7520,N_3344,N_6001);
nand U7521 (N_7521,N_3881,N_5479);
xnor U7522 (N_7522,N_5521,N_3685);
xor U7523 (N_7523,N_4845,N_4965);
xor U7524 (N_7524,N_5866,N_5155);
xnor U7525 (N_7525,N_4906,N_3218);
or U7526 (N_7526,N_5791,N_4326);
nor U7527 (N_7527,N_5158,N_4804);
or U7528 (N_7528,N_5701,N_3980);
nand U7529 (N_7529,N_5911,N_4260);
xor U7530 (N_7530,N_5176,N_3284);
nand U7531 (N_7531,N_4829,N_5418);
and U7532 (N_7532,N_5474,N_6144);
nand U7533 (N_7533,N_4584,N_3889);
nand U7534 (N_7534,N_5990,N_3274);
or U7535 (N_7535,N_4046,N_3539);
or U7536 (N_7536,N_5459,N_3157);
nand U7537 (N_7537,N_5976,N_3148);
xor U7538 (N_7538,N_3606,N_3836);
and U7539 (N_7539,N_4323,N_3598);
or U7540 (N_7540,N_4967,N_5835);
and U7541 (N_7541,N_5726,N_4755);
nand U7542 (N_7542,N_4419,N_3925);
xor U7543 (N_7543,N_4640,N_5851);
nor U7544 (N_7544,N_5522,N_5670);
and U7545 (N_7545,N_4918,N_5497);
nor U7546 (N_7546,N_4207,N_5579);
nand U7547 (N_7547,N_5817,N_5965);
nand U7548 (N_7548,N_3782,N_4067);
nand U7549 (N_7549,N_3542,N_5232);
nand U7550 (N_7550,N_4509,N_6005);
and U7551 (N_7551,N_4720,N_3534);
nand U7552 (N_7552,N_6054,N_5207);
nand U7553 (N_7553,N_3921,N_5036);
and U7554 (N_7554,N_4715,N_4437);
nor U7555 (N_7555,N_4205,N_3644);
nand U7556 (N_7556,N_5632,N_4711);
xor U7557 (N_7557,N_4726,N_4721);
xnor U7558 (N_7558,N_3465,N_3235);
and U7559 (N_7559,N_4846,N_3662);
and U7560 (N_7560,N_5323,N_3451);
nand U7561 (N_7561,N_4234,N_4070);
or U7562 (N_7562,N_3690,N_3167);
xnor U7563 (N_7563,N_3263,N_4371);
or U7564 (N_7564,N_5935,N_4235);
nand U7565 (N_7565,N_5802,N_5187);
xnor U7566 (N_7566,N_4975,N_4765);
nor U7567 (N_7567,N_4861,N_5714);
nand U7568 (N_7568,N_3792,N_5654);
xnor U7569 (N_7569,N_3435,N_3557);
and U7570 (N_7570,N_6016,N_3885);
nand U7571 (N_7571,N_4124,N_5099);
xnor U7572 (N_7572,N_4101,N_5143);
nand U7573 (N_7573,N_3900,N_4802);
nor U7574 (N_7574,N_3334,N_3655);
xor U7575 (N_7575,N_4127,N_3525);
and U7576 (N_7576,N_4890,N_3319);
xnor U7577 (N_7577,N_3560,N_4252);
or U7578 (N_7578,N_3659,N_4024);
nand U7579 (N_7579,N_5737,N_6119);
nor U7580 (N_7580,N_5392,N_5378);
or U7581 (N_7581,N_5880,N_6216);
or U7582 (N_7582,N_3602,N_4671);
and U7583 (N_7583,N_3293,N_4818);
and U7584 (N_7584,N_5057,N_5235);
and U7585 (N_7585,N_5828,N_5108);
or U7586 (N_7586,N_4233,N_5454);
xor U7587 (N_7587,N_3150,N_5277);
and U7588 (N_7588,N_3321,N_5402);
or U7589 (N_7589,N_5910,N_3974);
xor U7590 (N_7590,N_5815,N_5093);
nand U7591 (N_7591,N_3142,N_3332);
and U7592 (N_7592,N_3489,N_4662);
or U7593 (N_7593,N_3305,N_4102);
xor U7594 (N_7594,N_4210,N_4754);
nand U7595 (N_7595,N_6051,N_3532);
nand U7596 (N_7596,N_4852,N_4844);
xor U7597 (N_7597,N_6080,N_3928);
and U7598 (N_7598,N_6246,N_4946);
or U7599 (N_7599,N_6100,N_5792);
nor U7600 (N_7600,N_3424,N_3593);
and U7601 (N_7601,N_5943,N_5682);
xor U7602 (N_7602,N_3141,N_4883);
nand U7603 (N_7603,N_4109,N_5978);
nand U7604 (N_7604,N_6193,N_5999);
or U7605 (N_7605,N_4062,N_6143);
nand U7606 (N_7606,N_5756,N_4750);
or U7607 (N_7607,N_6146,N_3541);
nor U7608 (N_7608,N_4924,N_5563);
xor U7609 (N_7609,N_6235,N_5500);
xor U7610 (N_7610,N_5678,N_5853);
or U7611 (N_7611,N_4098,N_5587);
nand U7612 (N_7612,N_5748,N_6068);
nand U7613 (N_7613,N_5933,N_3145);
xnor U7614 (N_7614,N_3741,N_5195);
and U7615 (N_7615,N_5280,N_4534);
xnor U7616 (N_7616,N_6137,N_6207);
nor U7617 (N_7617,N_5845,N_5975);
nand U7618 (N_7618,N_4554,N_4438);
and U7619 (N_7619,N_5434,N_3795);
nand U7620 (N_7620,N_5427,N_4854);
and U7621 (N_7621,N_3804,N_6007);
or U7622 (N_7622,N_5485,N_5360);
xnor U7623 (N_7623,N_5540,N_5044);
or U7624 (N_7624,N_4432,N_3976);
or U7625 (N_7625,N_4115,N_3595);
or U7626 (N_7626,N_4899,N_3517);
or U7627 (N_7627,N_3617,N_3300);
or U7628 (N_7628,N_5883,N_5238);
xor U7629 (N_7629,N_4738,N_4349);
nor U7630 (N_7630,N_6027,N_5552);
xor U7631 (N_7631,N_3181,N_4731);
nand U7632 (N_7632,N_3737,N_5458);
or U7633 (N_7633,N_4773,N_3597);
nand U7634 (N_7634,N_3249,N_4346);
nor U7635 (N_7635,N_4385,N_5709);
xor U7636 (N_7636,N_5683,N_6189);
xnor U7637 (N_7637,N_3449,N_5435);
nor U7638 (N_7638,N_3934,N_6123);
xnor U7639 (N_7639,N_4645,N_3801);
xnor U7640 (N_7640,N_5946,N_4297);
xnor U7641 (N_7641,N_3407,N_4874);
and U7642 (N_7642,N_4393,N_4513);
nand U7643 (N_7643,N_4399,N_6089);
xnor U7644 (N_7644,N_4653,N_4145);
nand U7645 (N_7645,N_5966,N_6046);
xnor U7646 (N_7646,N_5518,N_5348);
xnor U7647 (N_7647,N_3553,N_4375);
xnor U7648 (N_7648,N_5754,N_4156);
or U7649 (N_7649,N_4037,N_4241);
or U7650 (N_7650,N_3499,N_4003);
and U7651 (N_7651,N_4493,N_3596);
nor U7652 (N_7652,N_3468,N_3453);
nor U7653 (N_7653,N_6094,N_3990);
xnor U7654 (N_7654,N_3730,N_3485);
nor U7655 (N_7655,N_4222,N_5929);
and U7656 (N_7656,N_3936,N_5680);
nand U7657 (N_7657,N_5056,N_4404);
or U7658 (N_7658,N_3198,N_6011);
or U7659 (N_7659,N_4708,N_4623);
nand U7660 (N_7660,N_3213,N_5106);
xor U7661 (N_7661,N_5114,N_4428);
or U7662 (N_7662,N_4358,N_3821);
xor U7663 (N_7663,N_4783,N_3358);
and U7664 (N_7664,N_4378,N_3645);
nand U7665 (N_7665,N_3336,N_4112);
xor U7666 (N_7666,N_4198,N_4267);
nand U7667 (N_7667,N_4654,N_3738);
xnor U7668 (N_7668,N_3515,N_4446);
nand U7669 (N_7669,N_5331,N_6078);
xnor U7670 (N_7670,N_3488,N_5234);
nor U7671 (N_7671,N_3837,N_6182);
nor U7672 (N_7672,N_4932,N_4483);
nand U7673 (N_7673,N_6036,N_3490);
nand U7674 (N_7674,N_3369,N_5713);
nand U7675 (N_7675,N_4056,N_4045);
nor U7676 (N_7676,N_5765,N_5104);
xor U7677 (N_7677,N_6224,N_6195);
nor U7678 (N_7678,N_4445,N_4343);
or U7679 (N_7679,N_5450,N_3780);
nand U7680 (N_7680,N_6218,N_4194);
nor U7681 (N_7681,N_3828,N_4354);
nor U7682 (N_7682,N_5248,N_4179);
and U7683 (N_7683,N_5718,N_3652);
nand U7684 (N_7684,N_6095,N_4142);
nor U7685 (N_7685,N_5669,N_3594);
or U7686 (N_7686,N_4277,N_4843);
nand U7687 (N_7687,N_4072,N_5648);
xor U7688 (N_7688,N_5206,N_5829);
and U7689 (N_7689,N_4579,N_3280);
nor U7690 (N_7690,N_4245,N_4357);
and U7691 (N_7691,N_6029,N_6220);
nor U7692 (N_7692,N_5433,N_6065);
or U7693 (N_7693,N_4118,N_5064);
nor U7694 (N_7694,N_5122,N_4547);
and U7695 (N_7695,N_5749,N_6010);
nand U7696 (N_7696,N_4572,N_5148);
nor U7697 (N_7697,N_5583,N_4660);
nor U7698 (N_7698,N_6053,N_4036);
or U7699 (N_7699,N_3919,N_4308);
xnor U7700 (N_7700,N_3312,N_3172);
nor U7701 (N_7701,N_5869,N_4748);
and U7702 (N_7702,N_3464,N_4800);
or U7703 (N_7703,N_4997,N_4122);
nor U7704 (N_7704,N_3493,N_3323);
nor U7705 (N_7705,N_4169,N_5676);
and U7706 (N_7706,N_4705,N_5466);
or U7707 (N_7707,N_4328,N_3688);
nand U7708 (N_7708,N_4588,N_5050);
or U7709 (N_7709,N_3680,N_4254);
nor U7710 (N_7710,N_4670,N_5110);
xnor U7711 (N_7711,N_4025,N_6040);
nor U7712 (N_7712,N_5729,N_5097);
nor U7713 (N_7713,N_4197,N_4039);
nand U7714 (N_7714,N_4828,N_4265);
nor U7715 (N_7715,N_4531,N_5955);
or U7716 (N_7716,N_6085,N_5710);
xor U7717 (N_7717,N_5604,N_5081);
nor U7718 (N_7718,N_5691,N_5107);
nand U7719 (N_7719,N_4785,N_3938);
nor U7720 (N_7720,N_3561,N_3434);
xor U7721 (N_7721,N_3211,N_5310);
nand U7722 (N_7722,N_5550,N_4719);
nand U7723 (N_7723,N_4700,N_3669);
nand U7724 (N_7724,N_4567,N_3773);
or U7725 (N_7725,N_5629,N_4416);
nor U7726 (N_7726,N_4099,N_3520);
or U7727 (N_7727,N_4456,N_4577);
nor U7728 (N_7728,N_4409,N_3303);
and U7729 (N_7729,N_4971,N_3946);
or U7730 (N_7730,N_3346,N_5739);
and U7731 (N_7731,N_5060,N_4921);
and U7732 (N_7732,N_4407,N_3567);
nand U7733 (N_7733,N_6139,N_3458);
nand U7734 (N_7734,N_5843,N_5530);
or U7735 (N_7735,N_4272,N_4560);
xnor U7736 (N_7736,N_4542,N_3327);
nor U7737 (N_7737,N_5724,N_3840);
nand U7738 (N_7738,N_3803,N_3331);
or U7739 (N_7739,N_4611,N_4869);
nor U7740 (N_7740,N_5214,N_3749);
or U7741 (N_7741,N_4848,N_3752);
nand U7742 (N_7742,N_4823,N_4310);
nand U7743 (N_7743,N_4116,N_3882);
and U7744 (N_7744,N_4901,N_5879);
nor U7745 (N_7745,N_6039,N_4496);
or U7746 (N_7746,N_3419,N_3378);
xnor U7747 (N_7747,N_4889,N_3920);
nand U7748 (N_7748,N_4394,N_5379);
xor U7749 (N_7749,N_5487,N_3622);
nor U7750 (N_7750,N_4151,N_6155);
nand U7751 (N_7751,N_5210,N_6229);
nand U7752 (N_7752,N_5381,N_3241);
and U7753 (N_7753,N_6120,N_5839);
and U7754 (N_7754,N_6071,N_5224);
xnor U7755 (N_7755,N_4716,N_6199);
or U7756 (N_7756,N_4954,N_4264);
nor U7757 (N_7757,N_4702,N_3256);
or U7758 (N_7758,N_3250,N_4041);
or U7759 (N_7759,N_5140,N_3475);
nor U7760 (N_7760,N_3797,N_4872);
nand U7761 (N_7761,N_3189,N_5591);
or U7762 (N_7762,N_3753,N_5704);
nor U7763 (N_7763,N_6160,N_5154);
xnor U7764 (N_7764,N_3977,N_4851);
or U7765 (N_7765,N_3132,N_4414);
or U7766 (N_7766,N_3292,N_4644);
xor U7767 (N_7767,N_5525,N_5895);
nand U7768 (N_7768,N_3252,N_5720);
nand U7769 (N_7769,N_5283,N_4353);
and U7770 (N_7770,N_3884,N_3575);
nor U7771 (N_7771,N_5984,N_4340);
xor U7772 (N_7772,N_3156,N_4166);
nand U7773 (N_7773,N_3272,N_3290);
nor U7774 (N_7774,N_5776,N_4594);
nor U7775 (N_7775,N_3861,N_3260);
and U7776 (N_7776,N_4086,N_6171);
and U7777 (N_7777,N_4622,N_3793);
xor U7778 (N_7778,N_3404,N_5204);
and U7779 (N_7779,N_3514,N_3638);
and U7780 (N_7780,N_5651,N_5751);
and U7781 (N_7781,N_3722,N_5549);
and U7782 (N_7782,N_6115,N_4659);
nand U7783 (N_7783,N_3687,N_5405);
nand U7784 (N_7784,N_5291,N_5611);
nor U7785 (N_7785,N_4734,N_5166);
xor U7786 (N_7786,N_3436,N_4022);
and U7787 (N_7787,N_5020,N_5200);
or U7788 (N_7788,N_3816,N_3403);
nand U7789 (N_7789,N_3915,N_3185);
or U7790 (N_7790,N_5292,N_5260);
nor U7791 (N_7791,N_3988,N_6116);
xnor U7792 (N_7792,N_4408,N_5679);
xnor U7793 (N_7793,N_4081,N_3846);
and U7794 (N_7794,N_3259,N_3873);
xnor U7795 (N_7795,N_3477,N_3379);
nand U7796 (N_7796,N_4795,N_6188);
and U7797 (N_7797,N_4904,N_6209);
or U7798 (N_7798,N_5441,N_4373);
xor U7799 (N_7799,N_5184,N_5856);
or U7800 (N_7800,N_3405,N_4090);
nor U7801 (N_7801,N_5997,N_4420);
or U7802 (N_7802,N_4466,N_5001);
xnor U7803 (N_7803,N_6060,N_4295);
nor U7804 (N_7804,N_4871,N_4114);
or U7805 (N_7805,N_5426,N_5956);
nand U7806 (N_7806,N_5826,N_4079);
or U7807 (N_7807,N_3395,N_5952);
nand U7808 (N_7808,N_4215,N_5558);
and U7809 (N_7809,N_6052,N_3772);
nand U7810 (N_7810,N_3367,N_3282);
nand U7811 (N_7811,N_5325,N_3855);
and U7812 (N_7812,N_4153,N_4060);
nor U7813 (N_7813,N_3750,N_3437);
xnor U7814 (N_7814,N_6011,N_4567);
or U7815 (N_7815,N_5655,N_4121);
and U7816 (N_7816,N_5708,N_4478);
or U7817 (N_7817,N_3847,N_4823);
and U7818 (N_7818,N_5059,N_3865);
nor U7819 (N_7819,N_4897,N_4487);
xor U7820 (N_7820,N_4666,N_3689);
or U7821 (N_7821,N_6088,N_3684);
or U7822 (N_7822,N_3665,N_6138);
xnor U7823 (N_7823,N_4021,N_4686);
nor U7824 (N_7824,N_5016,N_4602);
or U7825 (N_7825,N_5791,N_5105);
xor U7826 (N_7826,N_3134,N_4923);
and U7827 (N_7827,N_3281,N_4180);
nand U7828 (N_7828,N_6030,N_3349);
nor U7829 (N_7829,N_5553,N_4881);
nand U7830 (N_7830,N_5737,N_3306);
nand U7831 (N_7831,N_4119,N_3770);
nor U7832 (N_7832,N_5724,N_6020);
and U7833 (N_7833,N_4727,N_5328);
nor U7834 (N_7834,N_6115,N_4829);
or U7835 (N_7835,N_4910,N_3231);
nand U7836 (N_7836,N_5849,N_5806);
and U7837 (N_7837,N_3295,N_5693);
nor U7838 (N_7838,N_5033,N_5469);
or U7839 (N_7839,N_3691,N_5196);
nand U7840 (N_7840,N_5961,N_5128);
xnor U7841 (N_7841,N_3879,N_4945);
and U7842 (N_7842,N_5464,N_3591);
xor U7843 (N_7843,N_3317,N_5315);
nor U7844 (N_7844,N_4477,N_5236);
or U7845 (N_7845,N_5217,N_4764);
nor U7846 (N_7846,N_5307,N_4499);
or U7847 (N_7847,N_5045,N_5146);
or U7848 (N_7848,N_3529,N_5105);
and U7849 (N_7849,N_5328,N_4959);
nor U7850 (N_7850,N_3737,N_4168);
nor U7851 (N_7851,N_5400,N_4158);
or U7852 (N_7852,N_3935,N_3229);
xor U7853 (N_7853,N_4413,N_6114);
nor U7854 (N_7854,N_3240,N_3210);
or U7855 (N_7855,N_4377,N_5342);
and U7856 (N_7856,N_6117,N_5113);
xor U7857 (N_7857,N_4976,N_4551);
nand U7858 (N_7858,N_5638,N_4891);
and U7859 (N_7859,N_3660,N_5345);
nor U7860 (N_7860,N_5144,N_5322);
or U7861 (N_7861,N_4913,N_5587);
or U7862 (N_7862,N_5966,N_4236);
nand U7863 (N_7863,N_5303,N_4121);
or U7864 (N_7864,N_3858,N_4682);
and U7865 (N_7865,N_4157,N_3142);
nand U7866 (N_7866,N_5594,N_6244);
nor U7867 (N_7867,N_5898,N_4305);
nand U7868 (N_7868,N_3372,N_5178);
nand U7869 (N_7869,N_3746,N_4817);
nand U7870 (N_7870,N_4103,N_3740);
and U7871 (N_7871,N_4463,N_4507);
or U7872 (N_7872,N_4147,N_4395);
and U7873 (N_7873,N_4884,N_4559);
xnor U7874 (N_7874,N_3928,N_5271);
xor U7875 (N_7875,N_5209,N_5681);
nand U7876 (N_7876,N_3559,N_3747);
or U7877 (N_7877,N_4552,N_4972);
or U7878 (N_7878,N_4949,N_5753);
nand U7879 (N_7879,N_3437,N_5027);
or U7880 (N_7880,N_5175,N_3633);
or U7881 (N_7881,N_5970,N_3932);
xnor U7882 (N_7882,N_5237,N_3606);
nor U7883 (N_7883,N_3336,N_5440);
and U7884 (N_7884,N_3291,N_5512);
nand U7885 (N_7885,N_4975,N_3461);
xor U7886 (N_7886,N_4218,N_4318);
and U7887 (N_7887,N_3617,N_4342);
nand U7888 (N_7888,N_5053,N_5783);
nor U7889 (N_7889,N_5026,N_4323);
xnor U7890 (N_7890,N_4205,N_4390);
nor U7891 (N_7891,N_3369,N_3562);
and U7892 (N_7892,N_5273,N_4389);
nor U7893 (N_7893,N_4967,N_4841);
xnor U7894 (N_7894,N_4004,N_5369);
nand U7895 (N_7895,N_5443,N_3308);
or U7896 (N_7896,N_4579,N_3579);
nand U7897 (N_7897,N_6101,N_5712);
nand U7898 (N_7898,N_5931,N_6084);
and U7899 (N_7899,N_6207,N_3204);
xnor U7900 (N_7900,N_5043,N_3143);
and U7901 (N_7901,N_5229,N_4026);
nor U7902 (N_7902,N_4298,N_5023);
nand U7903 (N_7903,N_5179,N_3813);
and U7904 (N_7904,N_4069,N_3602);
or U7905 (N_7905,N_4909,N_5874);
xor U7906 (N_7906,N_6235,N_4536);
nor U7907 (N_7907,N_4881,N_6165);
nor U7908 (N_7908,N_5111,N_4801);
xor U7909 (N_7909,N_6206,N_4254);
nand U7910 (N_7910,N_5448,N_5882);
or U7911 (N_7911,N_3134,N_3388);
and U7912 (N_7912,N_6098,N_3211);
xor U7913 (N_7913,N_5049,N_6135);
or U7914 (N_7914,N_4583,N_5950);
and U7915 (N_7915,N_4472,N_5575);
xnor U7916 (N_7916,N_4180,N_6242);
nor U7917 (N_7917,N_4514,N_4439);
or U7918 (N_7918,N_5505,N_5351);
and U7919 (N_7919,N_3927,N_3353);
or U7920 (N_7920,N_5592,N_3557);
or U7921 (N_7921,N_4638,N_5361);
and U7922 (N_7922,N_5642,N_4602);
or U7923 (N_7923,N_4284,N_4514);
and U7924 (N_7924,N_4175,N_4785);
nand U7925 (N_7925,N_4922,N_4068);
or U7926 (N_7926,N_5759,N_6116);
and U7927 (N_7927,N_4134,N_3718);
xor U7928 (N_7928,N_4653,N_6099);
or U7929 (N_7929,N_3173,N_4932);
or U7930 (N_7930,N_5636,N_5174);
nor U7931 (N_7931,N_5029,N_5048);
or U7932 (N_7932,N_3381,N_4407);
and U7933 (N_7933,N_4486,N_4081);
or U7934 (N_7934,N_5385,N_5562);
nand U7935 (N_7935,N_5965,N_5784);
or U7936 (N_7936,N_3677,N_3586);
or U7937 (N_7937,N_4728,N_3923);
nor U7938 (N_7938,N_3518,N_6052);
nand U7939 (N_7939,N_3338,N_4610);
xor U7940 (N_7940,N_4610,N_4715);
xnor U7941 (N_7941,N_5992,N_3732);
or U7942 (N_7942,N_3534,N_4780);
or U7943 (N_7943,N_4047,N_4252);
or U7944 (N_7944,N_5530,N_4114);
nor U7945 (N_7945,N_3669,N_5649);
nand U7946 (N_7946,N_3979,N_4121);
nor U7947 (N_7947,N_4320,N_3770);
or U7948 (N_7948,N_4938,N_4200);
and U7949 (N_7949,N_5970,N_5816);
xnor U7950 (N_7950,N_4361,N_5167);
or U7951 (N_7951,N_5636,N_5810);
or U7952 (N_7952,N_5009,N_6229);
nand U7953 (N_7953,N_4904,N_6157);
xor U7954 (N_7954,N_4550,N_5137);
or U7955 (N_7955,N_3238,N_5426);
and U7956 (N_7956,N_5387,N_3683);
nand U7957 (N_7957,N_5777,N_6130);
nand U7958 (N_7958,N_3807,N_3186);
nor U7959 (N_7959,N_4092,N_5980);
and U7960 (N_7960,N_5744,N_6247);
and U7961 (N_7961,N_3331,N_4188);
nand U7962 (N_7962,N_3411,N_6221);
nand U7963 (N_7963,N_6141,N_6177);
nor U7964 (N_7964,N_3370,N_3360);
nand U7965 (N_7965,N_5583,N_4693);
or U7966 (N_7966,N_4140,N_3990);
xor U7967 (N_7967,N_4580,N_5023);
nor U7968 (N_7968,N_5071,N_5592);
nor U7969 (N_7969,N_3276,N_4353);
nor U7970 (N_7970,N_3704,N_5263);
nor U7971 (N_7971,N_3946,N_3901);
or U7972 (N_7972,N_3665,N_3251);
xor U7973 (N_7973,N_4813,N_6100);
xor U7974 (N_7974,N_4287,N_5766);
xnor U7975 (N_7975,N_4925,N_3533);
and U7976 (N_7976,N_5928,N_5190);
and U7977 (N_7977,N_6089,N_5001);
nand U7978 (N_7978,N_6119,N_3935);
and U7979 (N_7979,N_5409,N_5958);
nor U7980 (N_7980,N_5612,N_4295);
and U7981 (N_7981,N_3656,N_4899);
or U7982 (N_7982,N_4892,N_5211);
nor U7983 (N_7983,N_4964,N_3447);
nor U7984 (N_7984,N_4858,N_4818);
nor U7985 (N_7985,N_3933,N_3342);
and U7986 (N_7986,N_4772,N_3589);
nor U7987 (N_7987,N_3256,N_4932);
and U7988 (N_7988,N_3918,N_4030);
xor U7989 (N_7989,N_3743,N_5441);
and U7990 (N_7990,N_4969,N_4155);
nand U7991 (N_7991,N_3136,N_6247);
xnor U7992 (N_7992,N_4588,N_3970);
and U7993 (N_7993,N_3153,N_4310);
nor U7994 (N_7994,N_3604,N_3575);
or U7995 (N_7995,N_4266,N_6031);
or U7996 (N_7996,N_3670,N_4537);
nor U7997 (N_7997,N_3931,N_4665);
nand U7998 (N_7998,N_4932,N_5952);
xor U7999 (N_7999,N_5744,N_3703);
xor U8000 (N_8000,N_5360,N_3455);
or U8001 (N_8001,N_4629,N_3186);
or U8002 (N_8002,N_3981,N_4843);
nor U8003 (N_8003,N_4222,N_4718);
xor U8004 (N_8004,N_3542,N_5123);
nor U8005 (N_8005,N_5317,N_3364);
nand U8006 (N_8006,N_5993,N_4085);
nand U8007 (N_8007,N_5246,N_4334);
or U8008 (N_8008,N_4164,N_3338);
xor U8009 (N_8009,N_5219,N_4823);
nor U8010 (N_8010,N_4204,N_6247);
nand U8011 (N_8011,N_3533,N_5909);
nor U8012 (N_8012,N_3902,N_4603);
nand U8013 (N_8013,N_3142,N_3842);
nor U8014 (N_8014,N_5290,N_3140);
or U8015 (N_8015,N_4019,N_5186);
and U8016 (N_8016,N_3859,N_4922);
nor U8017 (N_8017,N_5218,N_3857);
nor U8018 (N_8018,N_4471,N_3412);
or U8019 (N_8019,N_4328,N_5272);
xnor U8020 (N_8020,N_5738,N_4513);
and U8021 (N_8021,N_4742,N_5662);
and U8022 (N_8022,N_4944,N_3853);
and U8023 (N_8023,N_4988,N_4168);
nor U8024 (N_8024,N_3862,N_3990);
nor U8025 (N_8025,N_6150,N_4498);
and U8026 (N_8026,N_4448,N_4429);
and U8027 (N_8027,N_5635,N_3607);
nor U8028 (N_8028,N_3616,N_5083);
or U8029 (N_8029,N_4432,N_5539);
and U8030 (N_8030,N_5152,N_6191);
and U8031 (N_8031,N_6170,N_5393);
nand U8032 (N_8032,N_3869,N_3549);
or U8033 (N_8033,N_3315,N_3204);
nand U8034 (N_8034,N_3933,N_6047);
nand U8035 (N_8035,N_3746,N_5318);
xnor U8036 (N_8036,N_5238,N_3268);
nor U8037 (N_8037,N_3923,N_4517);
xnor U8038 (N_8038,N_3674,N_5067);
xnor U8039 (N_8039,N_4020,N_5966);
nand U8040 (N_8040,N_6176,N_3496);
xor U8041 (N_8041,N_5479,N_5277);
nor U8042 (N_8042,N_4364,N_6135);
nor U8043 (N_8043,N_3438,N_3666);
nand U8044 (N_8044,N_4416,N_5378);
nand U8045 (N_8045,N_4368,N_3921);
nor U8046 (N_8046,N_5893,N_6249);
xnor U8047 (N_8047,N_5808,N_4593);
and U8048 (N_8048,N_5304,N_5102);
or U8049 (N_8049,N_6030,N_6061);
nand U8050 (N_8050,N_6222,N_3666);
xor U8051 (N_8051,N_4393,N_5341);
nand U8052 (N_8052,N_3355,N_3126);
or U8053 (N_8053,N_3355,N_4611);
nand U8054 (N_8054,N_3965,N_3867);
and U8055 (N_8055,N_3726,N_4408);
nand U8056 (N_8056,N_5264,N_5223);
or U8057 (N_8057,N_3559,N_3681);
and U8058 (N_8058,N_6080,N_5377);
nor U8059 (N_8059,N_5983,N_3382);
or U8060 (N_8060,N_5365,N_4373);
or U8061 (N_8061,N_3270,N_5555);
nand U8062 (N_8062,N_3960,N_5010);
or U8063 (N_8063,N_5484,N_3773);
and U8064 (N_8064,N_4994,N_4425);
xnor U8065 (N_8065,N_5345,N_3798);
nand U8066 (N_8066,N_4632,N_4427);
nand U8067 (N_8067,N_4089,N_3755);
nor U8068 (N_8068,N_3824,N_5032);
xor U8069 (N_8069,N_5556,N_3665);
nand U8070 (N_8070,N_4150,N_3875);
xnor U8071 (N_8071,N_6223,N_5187);
xnor U8072 (N_8072,N_5327,N_3522);
or U8073 (N_8073,N_5120,N_4110);
and U8074 (N_8074,N_3383,N_4516);
nand U8075 (N_8075,N_3988,N_6184);
and U8076 (N_8076,N_6079,N_5648);
and U8077 (N_8077,N_5592,N_5422);
nand U8078 (N_8078,N_5941,N_4965);
nor U8079 (N_8079,N_3251,N_4834);
and U8080 (N_8080,N_3728,N_5379);
nor U8081 (N_8081,N_3748,N_3764);
nand U8082 (N_8082,N_4482,N_6083);
nor U8083 (N_8083,N_5645,N_4269);
and U8084 (N_8084,N_3739,N_3647);
and U8085 (N_8085,N_5688,N_4550);
xor U8086 (N_8086,N_3470,N_5501);
nand U8087 (N_8087,N_5419,N_3323);
nor U8088 (N_8088,N_5328,N_3202);
nand U8089 (N_8089,N_3694,N_4086);
nand U8090 (N_8090,N_5688,N_4492);
nor U8091 (N_8091,N_5582,N_5659);
and U8092 (N_8092,N_4122,N_4256);
or U8093 (N_8093,N_5100,N_4321);
and U8094 (N_8094,N_4159,N_4473);
or U8095 (N_8095,N_4946,N_4131);
nor U8096 (N_8096,N_5173,N_5745);
nand U8097 (N_8097,N_3328,N_4323);
or U8098 (N_8098,N_4339,N_5297);
nor U8099 (N_8099,N_6005,N_5211);
nor U8100 (N_8100,N_5847,N_5099);
nand U8101 (N_8101,N_3546,N_3666);
or U8102 (N_8102,N_4985,N_6051);
and U8103 (N_8103,N_5682,N_6106);
nand U8104 (N_8104,N_4240,N_3880);
nor U8105 (N_8105,N_5813,N_4281);
xor U8106 (N_8106,N_4764,N_5952);
or U8107 (N_8107,N_5565,N_3538);
nand U8108 (N_8108,N_6148,N_3982);
and U8109 (N_8109,N_4732,N_6204);
xnor U8110 (N_8110,N_4122,N_3612);
nor U8111 (N_8111,N_3416,N_4779);
xnor U8112 (N_8112,N_4657,N_6076);
xor U8113 (N_8113,N_4872,N_4633);
or U8114 (N_8114,N_4797,N_5771);
and U8115 (N_8115,N_5092,N_4010);
nor U8116 (N_8116,N_3339,N_5684);
nand U8117 (N_8117,N_5309,N_3746);
or U8118 (N_8118,N_4130,N_5530);
xnor U8119 (N_8119,N_5110,N_5038);
nor U8120 (N_8120,N_5654,N_3813);
nor U8121 (N_8121,N_5126,N_4510);
or U8122 (N_8122,N_4653,N_5572);
nand U8123 (N_8123,N_4947,N_4466);
nor U8124 (N_8124,N_4779,N_4382);
xor U8125 (N_8125,N_5648,N_5824);
nor U8126 (N_8126,N_5323,N_5302);
and U8127 (N_8127,N_3613,N_5931);
xnor U8128 (N_8128,N_3805,N_4781);
xnor U8129 (N_8129,N_6187,N_4426);
or U8130 (N_8130,N_4960,N_5680);
nor U8131 (N_8131,N_4244,N_4251);
xor U8132 (N_8132,N_5158,N_3416);
xnor U8133 (N_8133,N_3872,N_4415);
xnor U8134 (N_8134,N_3956,N_5594);
and U8135 (N_8135,N_6073,N_3773);
or U8136 (N_8136,N_3274,N_4052);
xor U8137 (N_8137,N_3617,N_5572);
or U8138 (N_8138,N_5810,N_3385);
xor U8139 (N_8139,N_4302,N_4059);
or U8140 (N_8140,N_5790,N_6183);
and U8141 (N_8141,N_6187,N_5434);
nor U8142 (N_8142,N_5374,N_5392);
and U8143 (N_8143,N_3501,N_5263);
xnor U8144 (N_8144,N_5551,N_4313);
or U8145 (N_8145,N_3378,N_4055);
nand U8146 (N_8146,N_5534,N_5198);
or U8147 (N_8147,N_3339,N_4664);
and U8148 (N_8148,N_3785,N_3788);
and U8149 (N_8149,N_3419,N_6184);
nand U8150 (N_8150,N_3156,N_5303);
nor U8151 (N_8151,N_4904,N_3841);
xor U8152 (N_8152,N_5408,N_3261);
or U8153 (N_8153,N_4838,N_4724);
nand U8154 (N_8154,N_5233,N_5605);
and U8155 (N_8155,N_4996,N_5528);
nor U8156 (N_8156,N_5396,N_4340);
nand U8157 (N_8157,N_4168,N_5296);
nor U8158 (N_8158,N_3389,N_4844);
and U8159 (N_8159,N_4127,N_3393);
and U8160 (N_8160,N_5171,N_3628);
nand U8161 (N_8161,N_3366,N_6093);
nand U8162 (N_8162,N_5873,N_5104);
and U8163 (N_8163,N_5387,N_4333);
nand U8164 (N_8164,N_4235,N_3670);
or U8165 (N_8165,N_3141,N_4878);
nor U8166 (N_8166,N_5678,N_5562);
or U8167 (N_8167,N_4080,N_3885);
nand U8168 (N_8168,N_4267,N_4664);
or U8169 (N_8169,N_6033,N_3846);
or U8170 (N_8170,N_4244,N_4354);
and U8171 (N_8171,N_3581,N_5417);
nor U8172 (N_8172,N_5409,N_4884);
xnor U8173 (N_8173,N_5613,N_4086);
nand U8174 (N_8174,N_4753,N_4300);
nor U8175 (N_8175,N_4304,N_5399);
xnor U8176 (N_8176,N_4679,N_4630);
nand U8177 (N_8177,N_4007,N_4967);
and U8178 (N_8178,N_5443,N_4756);
xor U8179 (N_8179,N_5646,N_4488);
xor U8180 (N_8180,N_4949,N_4389);
nand U8181 (N_8181,N_4597,N_5815);
nor U8182 (N_8182,N_4792,N_5328);
and U8183 (N_8183,N_4852,N_3225);
and U8184 (N_8184,N_4643,N_6120);
xor U8185 (N_8185,N_5398,N_5636);
or U8186 (N_8186,N_4399,N_6179);
and U8187 (N_8187,N_5447,N_3163);
xor U8188 (N_8188,N_4358,N_4004);
nor U8189 (N_8189,N_6217,N_5343);
xor U8190 (N_8190,N_3337,N_4399);
nor U8191 (N_8191,N_5809,N_6159);
nand U8192 (N_8192,N_5605,N_3477);
nand U8193 (N_8193,N_3675,N_6162);
nand U8194 (N_8194,N_5109,N_4263);
and U8195 (N_8195,N_5681,N_5268);
nand U8196 (N_8196,N_3502,N_4804);
or U8197 (N_8197,N_5563,N_6105);
nor U8198 (N_8198,N_3474,N_3277);
xor U8199 (N_8199,N_5165,N_4506);
xor U8200 (N_8200,N_4116,N_5153);
nor U8201 (N_8201,N_3275,N_5505);
and U8202 (N_8202,N_5962,N_5052);
or U8203 (N_8203,N_3804,N_4716);
and U8204 (N_8204,N_5736,N_4144);
xnor U8205 (N_8205,N_6049,N_3916);
nor U8206 (N_8206,N_5065,N_3351);
and U8207 (N_8207,N_3330,N_5635);
nand U8208 (N_8208,N_4930,N_4313);
or U8209 (N_8209,N_5121,N_3142);
nor U8210 (N_8210,N_5263,N_4582);
xnor U8211 (N_8211,N_4583,N_6121);
nand U8212 (N_8212,N_4644,N_6009);
nor U8213 (N_8213,N_5504,N_3472);
nand U8214 (N_8214,N_5090,N_5350);
and U8215 (N_8215,N_4675,N_3759);
nand U8216 (N_8216,N_5096,N_3504);
nand U8217 (N_8217,N_5745,N_6169);
or U8218 (N_8218,N_4002,N_4906);
or U8219 (N_8219,N_5392,N_3455);
and U8220 (N_8220,N_3979,N_3985);
nand U8221 (N_8221,N_6002,N_6056);
and U8222 (N_8222,N_4084,N_5731);
and U8223 (N_8223,N_4829,N_3685);
nor U8224 (N_8224,N_5032,N_4053);
xor U8225 (N_8225,N_3193,N_3501);
and U8226 (N_8226,N_4312,N_4501);
and U8227 (N_8227,N_3953,N_5266);
xnor U8228 (N_8228,N_4215,N_3598);
nor U8229 (N_8229,N_4664,N_5146);
and U8230 (N_8230,N_5883,N_5133);
nand U8231 (N_8231,N_4625,N_4615);
xnor U8232 (N_8232,N_5607,N_5353);
and U8233 (N_8233,N_4000,N_4429);
nor U8234 (N_8234,N_5994,N_4652);
or U8235 (N_8235,N_6002,N_6061);
nand U8236 (N_8236,N_4717,N_4520);
or U8237 (N_8237,N_3157,N_6205);
nand U8238 (N_8238,N_4503,N_5645);
nand U8239 (N_8239,N_3211,N_4429);
nor U8240 (N_8240,N_5481,N_3428);
nand U8241 (N_8241,N_3482,N_4574);
and U8242 (N_8242,N_3954,N_4940);
or U8243 (N_8243,N_5968,N_3950);
and U8244 (N_8244,N_6132,N_5866);
and U8245 (N_8245,N_4342,N_3329);
nor U8246 (N_8246,N_4261,N_3685);
nor U8247 (N_8247,N_4197,N_3415);
or U8248 (N_8248,N_6137,N_5767);
nand U8249 (N_8249,N_3233,N_5098);
nor U8250 (N_8250,N_6108,N_5749);
nand U8251 (N_8251,N_4371,N_5287);
and U8252 (N_8252,N_5522,N_4633);
nand U8253 (N_8253,N_4123,N_5383);
nand U8254 (N_8254,N_5937,N_4577);
xnor U8255 (N_8255,N_4714,N_3360);
xnor U8256 (N_8256,N_5774,N_6114);
nand U8257 (N_8257,N_4211,N_3685);
and U8258 (N_8258,N_6159,N_4754);
nand U8259 (N_8259,N_4673,N_5845);
nand U8260 (N_8260,N_3765,N_4543);
xor U8261 (N_8261,N_5135,N_3371);
xnor U8262 (N_8262,N_4625,N_3258);
xnor U8263 (N_8263,N_5390,N_3796);
or U8264 (N_8264,N_5055,N_5554);
or U8265 (N_8265,N_4507,N_6083);
nand U8266 (N_8266,N_6115,N_5345);
xor U8267 (N_8267,N_5181,N_5899);
or U8268 (N_8268,N_4101,N_4214);
nand U8269 (N_8269,N_3859,N_3872);
xor U8270 (N_8270,N_3789,N_3376);
and U8271 (N_8271,N_3534,N_5114);
xor U8272 (N_8272,N_4917,N_4647);
or U8273 (N_8273,N_3953,N_5877);
and U8274 (N_8274,N_4554,N_4678);
nand U8275 (N_8275,N_3319,N_3687);
or U8276 (N_8276,N_4219,N_4727);
and U8277 (N_8277,N_3311,N_4776);
xor U8278 (N_8278,N_4586,N_5662);
or U8279 (N_8279,N_5206,N_5997);
and U8280 (N_8280,N_5234,N_4052);
nand U8281 (N_8281,N_6198,N_3239);
xor U8282 (N_8282,N_5190,N_4676);
nor U8283 (N_8283,N_4909,N_4133);
or U8284 (N_8284,N_4739,N_6035);
nor U8285 (N_8285,N_3879,N_5310);
nor U8286 (N_8286,N_5474,N_4689);
nor U8287 (N_8287,N_3987,N_4617);
or U8288 (N_8288,N_6078,N_6016);
nand U8289 (N_8289,N_5051,N_3348);
and U8290 (N_8290,N_5519,N_3890);
or U8291 (N_8291,N_5146,N_4451);
and U8292 (N_8292,N_6223,N_6158);
or U8293 (N_8293,N_5546,N_3931);
and U8294 (N_8294,N_5251,N_3882);
or U8295 (N_8295,N_3799,N_3526);
xnor U8296 (N_8296,N_3656,N_5428);
and U8297 (N_8297,N_5619,N_5106);
nor U8298 (N_8298,N_3956,N_5183);
or U8299 (N_8299,N_4924,N_6201);
xor U8300 (N_8300,N_4030,N_3820);
and U8301 (N_8301,N_5040,N_4645);
nor U8302 (N_8302,N_4673,N_3542);
and U8303 (N_8303,N_4091,N_4002);
nor U8304 (N_8304,N_5743,N_5940);
nand U8305 (N_8305,N_5911,N_4452);
nand U8306 (N_8306,N_4630,N_5194);
nor U8307 (N_8307,N_4342,N_5462);
nor U8308 (N_8308,N_5129,N_3630);
or U8309 (N_8309,N_3490,N_4920);
or U8310 (N_8310,N_6162,N_6144);
nand U8311 (N_8311,N_5592,N_4754);
nor U8312 (N_8312,N_4581,N_5160);
xnor U8313 (N_8313,N_3723,N_4385);
nor U8314 (N_8314,N_5945,N_4539);
nor U8315 (N_8315,N_3550,N_5207);
nor U8316 (N_8316,N_3327,N_3866);
nand U8317 (N_8317,N_3696,N_4957);
nor U8318 (N_8318,N_3255,N_3195);
or U8319 (N_8319,N_3216,N_4473);
xor U8320 (N_8320,N_5822,N_3794);
nor U8321 (N_8321,N_4736,N_3613);
nand U8322 (N_8322,N_3462,N_5391);
or U8323 (N_8323,N_4401,N_3572);
or U8324 (N_8324,N_3365,N_5817);
xnor U8325 (N_8325,N_5438,N_6156);
xnor U8326 (N_8326,N_5617,N_4940);
nand U8327 (N_8327,N_4147,N_5927);
nor U8328 (N_8328,N_3332,N_4676);
and U8329 (N_8329,N_6223,N_5697);
and U8330 (N_8330,N_3351,N_3315);
xnor U8331 (N_8331,N_3359,N_3822);
or U8332 (N_8332,N_3280,N_3652);
or U8333 (N_8333,N_3799,N_4184);
nand U8334 (N_8334,N_5323,N_3465);
nor U8335 (N_8335,N_3953,N_4207);
nand U8336 (N_8336,N_6015,N_3195);
nor U8337 (N_8337,N_4072,N_5582);
and U8338 (N_8338,N_3291,N_4267);
nand U8339 (N_8339,N_5317,N_4748);
xor U8340 (N_8340,N_3712,N_4349);
or U8341 (N_8341,N_5899,N_4651);
and U8342 (N_8342,N_5300,N_3541);
and U8343 (N_8343,N_3529,N_5659);
nor U8344 (N_8344,N_4015,N_5344);
nand U8345 (N_8345,N_3786,N_4099);
or U8346 (N_8346,N_3962,N_3704);
xnor U8347 (N_8347,N_4644,N_6101);
nor U8348 (N_8348,N_3765,N_4572);
nand U8349 (N_8349,N_3565,N_4571);
or U8350 (N_8350,N_4764,N_4164);
nor U8351 (N_8351,N_4580,N_6161);
xor U8352 (N_8352,N_4963,N_5487);
nor U8353 (N_8353,N_6139,N_4401);
nand U8354 (N_8354,N_4996,N_5976);
nor U8355 (N_8355,N_4318,N_4041);
nor U8356 (N_8356,N_6088,N_3987);
and U8357 (N_8357,N_3841,N_3753);
nand U8358 (N_8358,N_3551,N_5982);
or U8359 (N_8359,N_6177,N_5371);
and U8360 (N_8360,N_3967,N_4435);
or U8361 (N_8361,N_6185,N_5658);
and U8362 (N_8362,N_6161,N_5762);
xor U8363 (N_8363,N_4825,N_3464);
nor U8364 (N_8364,N_3909,N_5914);
nor U8365 (N_8365,N_3768,N_5646);
nand U8366 (N_8366,N_4979,N_4271);
or U8367 (N_8367,N_3699,N_5354);
nor U8368 (N_8368,N_4009,N_4267);
nand U8369 (N_8369,N_5559,N_4790);
and U8370 (N_8370,N_5401,N_4228);
nor U8371 (N_8371,N_4471,N_4248);
nor U8372 (N_8372,N_4793,N_5762);
nor U8373 (N_8373,N_6037,N_5897);
or U8374 (N_8374,N_5175,N_3659);
or U8375 (N_8375,N_5851,N_4509);
nand U8376 (N_8376,N_3626,N_4074);
xor U8377 (N_8377,N_5367,N_5887);
or U8378 (N_8378,N_3438,N_5154);
xnor U8379 (N_8379,N_3361,N_3945);
xnor U8380 (N_8380,N_3687,N_4059);
and U8381 (N_8381,N_3968,N_4095);
xor U8382 (N_8382,N_5007,N_4670);
xnor U8383 (N_8383,N_4897,N_5644);
and U8384 (N_8384,N_4638,N_3381);
and U8385 (N_8385,N_3418,N_3254);
and U8386 (N_8386,N_3441,N_5033);
nand U8387 (N_8387,N_3381,N_3302);
or U8388 (N_8388,N_5345,N_4765);
nand U8389 (N_8389,N_3393,N_4406);
or U8390 (N_8390,N_3261,N_4505);
nand U8391 (N_8391,N_5539,N_5819);
nor U8392 (N_8392,N_4884,N_4821);
nor U8393 (N_8393,N_3284,N_5395);
or U8394 (N_8394,N_4104,N_4260);
and U8395 (N_8395,N_3570,N_4652);
and U8396 (N_8396,N_5776,N_6035);
nand U8397 (N_8397,N_6215,N_3884);
nand U8398 (N_8398,N_5811,N_4698);
xnor U8399 (N_8399,N_4142,N_4296);
nand U8400 (N_8400,N_4822,N_6121);
and U8401 (N_8401,N_4147,N_4207);
nor U8402 (N_8402,N_4255,N_5385);
and U8403 (N_8403,N_3930,N_6009);
xnor U8404 (N_8404,N_4584,N_5979);
nor U8405 (N_8405,N_6143,N_6093);
or U8406 (N_8406,N_6026,N_4574);
xor U8407 (N_8407,N_3457,N_5727);
nor U8408 (N_8408,N_5536,N_4695);
and U8409 (N_8409,N_4562,N_5402);
nor U8410 (N_8410,N_3867,N_3859);
or U8411 (N_8411,N_5468,N_3966);
and U8412 (N_8412,N_5374,N_3416);
and U8413 (N_8413,N_6011,N_3701);
nor U8414 (N_8414,N_5567,N_4387);
and U8415 (N_8415,N_3204,N_4658);
nand U8416 (N_8416,N_3357,N_4358);
xor U8417 (N_8417,N_5777,N_3892);
and U8418 (N_8418,N_5432,N_4820);
or U8419 (N_8419,N_5910,N_5935);
and U8420 (N_8420,N_4102,N_4151);
or U8421 (N_8421,N_4139,N_3194);
nand U8422 (N_8422,N_6153,N_5537);
and U8423 (N_8423,N_6197,N_3335);
and U8424 (N_8424,N_4997,N_5737);
and U8425 (N_8425,N_5352,N_3840);
nand U8426 (N_8426,N_4275,N_4636);
nand U8427 (N_8427,N_5825,N_3961);
or U8428 (N_8428,N_5399,N_4244);
nand U8429 (N_8429,N_4126,N_3825);
and U8430 (N_8430,N_4558,N_5035);
xor U8431 (N_8431,N_3392,N_3474);
or U8432 (N_8432,N_4343,N_6244);
and U8433 (N_8433,N_3327,N_3789);
nand U8434 (N_8434,N_3653,N_5416);
xor U8435 (N_8435,N_3198,N_5043);
xor U8436 (N_8436,N_3869,N_5277);
or U8437 (N_8437,N_3984,N_5474);
and U8438 (N_8438,N_5781,N_5391);
and U8439 (N_8439,N_5964,N_3547);
nand U8440 (N_8440,N_6075,N_4334);
xor U8441 (N_8441,N_5726,N_4907);
and U8442 (N_8442,N_3701,N_4697);
nor U8443 (N_8443,N_4033,N_3518);
xor U8444 (N_8444,N_5102,N_3604);
nand U8445 (N_8445,N_4257,N_3301);
xnor U8446 (N_8446,N_3689,N_4365);
nand U8447 (N_8447,N_5334,N_3195);
and U8448 (N_8448,N_4815,N_5563);
nand U8449 (N_8449,N_6169,N_4479);
and U8450 (N_8450,N_5133,N_4152);
nand U8451 (N_8451,N_5992,N_4504);
nand U8452 (N_8452,N_3624,N_3885);
or U8453 (N_8453,N_5538,N_5101);
and U8454 (N_8454,N_5247,N_3503);
xor U8455 (N_8455,N_5874,N_3910);
nor U8456 (N_8456,N_6059,N_4767);
or U8457 (N_8457,N_3550,N_4760);
and U8458 (N_8458,N_4877,N_6056);
nand U8459 (N_8459,N_5231,N_4930);
xor U8460 (N_8460,N_5927,N_3798);
nand U8461 (N_8461,N_5223,N_5138);
xnor U8462 (N_8462,N_3590,N_4060);
nand U8463 (N_8463,N_4209,N_5316);
and U8464 (N_8464,N_5675,N_4380);
or U8465 (N_8465,N_3428,N_4276);
nand U8466 (N_8466,N_5698,N_5823);
xor U8467 (N_8467,N_3520,N_6153);
or U8468 (N_8468,N_5655,N_5270);
and U8469 (N_8469,N_4475,N_4345);
or U8470 (N_8470,N_4065,N_5818);
and U8471 (N_8471,N_5841,N_4064);
xnor U8472 (N_8472,N_6100,N_3806);
nand U8473 (N_8473,N_5528,N_5987);
and U8474 (N_8474,N_4721,N_6013);
xnor U8475 (N_8475,N_3481,N_3521);
xor U8476 (N_8476,N_3995,N_3916);
xor U8477 (N_8477,N_3149,N_3529);
and U8478 (N_8478,N_4994,N_5265);
and U8479 (N_8479,N_3496,N_4983);
or U8480 (N_8480,N_5234,N_4365);
and U8481 (N_8481,N_4534,N_4515);
and U8482 (N_8482,N_4169,N_5047);
xnor U8483 (N_8483,N_5226,N_5090);
xor U8484 (N_8484,N_4872,N_4115);
or U8485 (N_8485,N_4531,N_5021);
nand U8486 (N_8486,N_4761,N_5982);
xor U8487 (N_8487,N_3148,N_4109);
and U8488 (N_8488,N_4041,N_3213);
nor U8489 (N_8489,N_5064,N_5810);
nor U8490 (N_8490,N_6057,N_4648);
nand U8491 (N_8491,N_4888,N_3125);
xor U8492 (N_8492,N_4723,N_3548);
xnor U8493 (N_8493,N_3684,N_4753);
nand U8494 (N_8494,N_4667,N_4717);
nand U8495 (N_8495,N_4592,N_3480);
or U8496 (N_8496,N_5788,N_6213);
nand U8497 (N_8497,N_3314,N_6222);
nand U8498 (N_8498,N_4950,N_5958);
nand U8499 (N_8499,N_3854,N_3141);
and U8500 (N_8500,N_5722,N_5050);
nor U8501 (N_8501,N_4940,N_4628);
xnor U8502 (N_8502,N_5921,N_4563);
xor U8503 (N_8503,N_4751,N_5823);
nor U8504 (N_8504,N_4199,N_3950);
xnor U8505 (N_8505,N_6006,N_3173);
or U8506 (N_8506,N_5322,N_5819);
xor U8507 (N_8507,N_5968,N_5904);
xnor U8508 (N_8508,N_5965,N_4603);
nand U8509 (N_8509,N_4893,N_3648);
nor U8510 (N_8510,N_4424,N_3337);
or U8511 (N_8511,N_4796,N_5760);
nand U8512 (N_8512,N_6194,N_5256);
nand U8513 (N_8513,N_3879,N_3663);
nand U8514 (N_8514,N_3586,N_6164);
xor U8515 (N_8515,N_4329,N_3687);
nand U8516 (N_8516,N_4782,N_4225);
xnor U8517 (N_8517,N_5891,N_3872);
nor U8518 (N_8518,N_5493,N_6199);
or U8519 (N_8519,N_4950,N_4665);
and U8520 (N_8520,N_3397,N_3816);
xnor U8521 (N_8521,N_4813,N_4107);
xor U8522 (N_8522,N_3970,N_5303);
xnor U8523 (N_8523,N_5151,N_4481);
nand U8524 (N_8524,N_5098,N_6136);
or U8525 (N_8525,N_3177,N_4887);
and U8526 (N_8526,N_5414,N_4986);
xnor U8527 (N_8527,N_4044,N_4943);
and U8528 (N_8528,N_3806,N_5896);
xor U8529 (N_8529,N_6137,N_3729);
and U8530 (N_8530,N_5053,N_4174);
and U8531 (N_8531,N_5673,N_3838);
or U8532 (N_8532,N_5883,N_5887);
xnor U8533 (N_8533,N_4186,N_3747);
or U8534 (N_8534,N_3422,N_5145);
nand U8535 (N_8535,N_4937,N_6045);
or U8536 (N_8536,N_4831,N_5173);
nand U8537 (N_8537,N_4449,N_4330);
xnor U8538 (N_8538,N_3643,N_4666);
xnor U8539 (N_8539,N_6145,N_5700);
nand U8540 (N_8540,N_6046,N_4430);
xor U8541 (N_8541,N_4122,N_3243);
xnor U8542 (N_8542,N_4254,N_5151);
or U8543 (N_8543,N_3207,N_5201);
nand U8544 (N_8544,N_5298,N_4116);
nand U8545 (N_8545,N_5510,N_5104);
and U8546 (N_8546,N_6222,N_5102);
nand U8547 (N_8547,N_5843,N_4664);
nand U8548 (N_8548,N_5089,N_4473);
and U8549 (N_8549,N_4232,N_3888);
nand U8550 (N_8550,N_4288,N_6008);
and U8551 (N_8551,N_3700,N_4079);
and U8552 (N_8552,N_5660,N_3650);
xor U8553 (N_8553,N_4184,N_4415);
nor U8554 (N_8554,N_4164,N_5900);
and U8555 (N_8555,N_5838,N_6128);
nor U8556 (N_8556,N_5460,N_3287);
nand U8557 (N_8557,N_5981,N_5445);
xnor U8558 (N_8558,N_4679,N_4566);
or U8559 (N_8559,N_3669,N_4467);
nand U8560 (N_8560,N_5539,N_3360);
nand U8561 (N_8561,N_4829,N_3410);
or U8562 (N_8562,N_4933,N_4382);
xor U8563 (N_8563,N_3515,N_4349);
nand U8564 (N_8564,N_4329,N_5282);
xor U8565 (N_8565,N_5001,N_4089);
nor U8566 (N_8566,N_3214,N_3442);
and U8567 (N_8567,N_3397,N_4930);
nor U8568 (N_8568,N_5437,N_5895);
and U8569 (N_8569,N_3343,N_4544);
nor U8570 (N_8570,N_3898,N_3689);
nand U8571 (N_8571,N_4965,N_6066);
nor U8572 (N_8572,N_3883,N_5780);
or U8573 (N_8573,N_5886,N_5682);
xor U8574 (N_8574,N_5716,N_6146);
nand U8575 (N_8575,N_3190,N_6157);
nor U8576 (N_8576,N_6227,N_4665);
or U8577 (N_8577,N_5306,N_3873);
and U8578 (N_8578,N_5203,N_3912);
xnor U8579 (N_8579,N_5550,N_4001);
nor U8580 (N_8580,N_4925,N_3327);
and U8581 (N_8581,N_5419,N_3340);
xor U8582 (N_8582,N_5325,N_3347);
and U8583 (N_8583,N_5032,N_4997);
nand U8584 (N_8584,N_3906,N_3375);
or U8585 (N_8585,N_4664,N_4822);
and U8586 (N_8586,N_4274,N_3140);
nor U8587 (N_8587,N_4765,N_5526);
xor U8588 (N_8588,N_3249,N_4612);
nand U8589 (N_8589,N_5736,N_5255);
nand U8590 (N_8590,N_5209,N_5376);
nor U8591 (N_8591,N_4630,N_3460);
or U8592 (N_8592,N_4060,N_3971);
nor U8593 (N_8593,N_4920,N_4397);
nand U8594 (N_8594,N_4816,N_5221);
and U8595 (N_8595,N_5897,N_5446);
nand U8596 (N_8596,N_3486,N_5958);
nor U8597 (N_8597,N_4319,N_4857);
and U8598 (N_8598,N_3386,N_3248);
nor U8599 (N_8599,N_5471,N_3501);
or U8600 (N_8600,N_6107,N_5420);
xor U8601 (N_8601,N_4284,N_6017);
nor U8602 (N_8602,N_3533,N_3723);
nand U8603 (N_8603,N_6079,N_4031);
xnor U8604 (N_8604,N_4588,N_4310);
xor U8605 (N_8605,N_3644,N_4490);
and U8606 (N_8606,N_3248,N_5578);
nand U8607 (N_8607,N_4239,N_4520);
xnor U8608 (N_8608,N_4019,N_3526);
or U8609 (N_8609,N_6002,N_4063);
or U8610 (N_8610,N_5081,N_5847);
nor U8611 (N_8611,N_3602,N_5854);
or U8612 (N_8612,N_6118,N_3827);
nand U8613 (N_8613,N_3140,N_5608);
nand U8614 (N_8614,N_3265,N_5013);
or U8615 (N_8615,N_6220,N_6030);
nor U8616 (N_8616,N_5570,N_5769);
and U8617 (N_8617,N_5558,N_4701);
nand U8618 (N_8618,N_5776,N_4093);
nor U8619 (N_8619,N_4857,N_6192);
nor U8620 (N_8620,N_5677,N_3964);
nand U8621 (N_8621,N_4867,N_3362);
or U8622 (N_8622,N_3293,N_4114);
or U8623 (N_8623,N_5030,N_3208);
and U8624 (N_8624,N_3690,N_3671);
xnor U8625 (N_8625,N_5865,N_5631);
nor U8626 (N_8626,N_3887,N_5561);
xor U8627 (N_8627,N_5254,N_5874);
xor U8628 (N_8628,N_5167,N_5483);
nor U8629 (N_8629,N_4679,N_6239);
and U8630 (N_8630,N_3137,N_6083);
nand U8631 (N_8631,N_4637,N_4438);
or U8632 (N_8632,N_4031,N_4709);
nor U8633 (N_8633,N_4243,N_5944);
or U8634 (N_8634,N_3699,N_5063);
nand U8635 (N_8635,N_5735,N_4657);
xnor U8636 (N_8636,N_4208,N_5051);
and U8637 (N_8637,N_3750,N_6173);
xnor U8638 (N_8638,N_4061,N_3310);
or U8639 (N_8639,N_3271,N_6216);
nor U8640 (N_8640,N_4542,N_5721);
nand U8641 (N_8641,N_3694,N_4100);
nor U8642 (N_8642,N_5362,N_4763);
xnor U8643 (N_8643,N_5833,N_5856);
xnor U8644 (N_8644,N_3937,N_5522);
and U8645 (N_8645,N_5283,N_4090);
or U8646 (N_8646,N_3452,N_4214);
xor U8647 (N_8647,N_6139,N_5692);
nand U8648 (N_8648,N_3239,N_3976);
xnor U8649 (N_8649,N_5357,N_4342);
or U8650 (N_8650,N_4792,N_5237);
xnor U8651 (N_8651,N_4201,N_5404);
or U8652 (N_8652,N_3809,N_5277);
nand U8653 (N_8653,N_5881,N_4111);
nand U8654 (N_8654,N_5247,N_5764);
or U8655 (N_8655,N_4919,N_5854);
and U8656 (N_8656,N_5940,N_4385);
and U8657 (N_8657,N_4023,N_5153);
xor U8658 (N_8658,N_3681,N_5579);
nor U8659 (N_8659,N_6050,N_3126);
and U8660 (N_8660,N_5826,N_5415);
and U8661 (N_8661,N_5652,N_5745);
nor U8662 (N_8662,N_6196,N_4545);
nor U8663 (N_8663,N_4102,N_4368);
nand U8664 (N_8664,N_6232,N_4779);
nand U8665 (N_8665,N_4917,N_4175);
and U8666 (N_8666,N_5648,N_3135);
nand U8667 (N_8667,N_4953,N_5804);
nor U8668 (N_8668,N_3433,N_3641);
or U8669 (N_8669,N_6233,N_5718);
and U8670 (N_8670,N_4177,N_3652);
nand U8671 (N_8671,N_4688,N_5499);
nor U8672 (N_8672,N_3589,N_3668);
xnor U8673 (N_8673,N_3190,N_4926);
nor U8674 (N_8674,N_4886,N_3701);
and U8675 (N_8675,N_3517,N_5599);
xnor U8676 (N_8676,N_5967,N_5952);
xnor U8677 (N_8677,N_5283,N_5246);
nand U8678 (N_8678,N_4734,N_5912);
or U8679 (N_8679,N_4188,N_5087);
and U8680 (N_8680,N_3604,N_4695);
nand U8681 (N_8681,N_5477,N_3539);
xnor U8682 (N_8682,N_5862,N_5583);
or U8683 (N_8683,N_4919,N_4295);
xnor U8684 (N_8684,N_4703,N_3847);
xnor U8685 (N_8685,N_5525,N_3605);
nor U8686 (N_8686,N_3398,N_3664);
nor U8687 (N_8687,N_6035,N_5097);
nand U8688 (N_8688,N_4291,N_4998);
or U8689 (N_8689,N_3195,N_4536);
or U8690 (N_8690,N_5204,N_3629);
nand U8691 (N_8691,N_5688,N_3405);
and U8692 (N_8692,N_5761,N_5659);
nand U8693 (N_8693,N_5613,N_3664);
xnor U8694 (N_8694,N_6052,N_3987);
and U8695 (N_8695,N_3873,N_3460);
nor U8696 (N_8696,N_6037,N_4396);
and U8697 (N_8697,N_3184,N_3949);
nor U8698 (N_8698,N_3915,N_3652);
or U8699 (N_8699,N_3658,N_3273);
and U8700 (N_8700,N_5360,N_6231);
and U8701 (N_8701,N_3157,N_5190);
or U8702 (N_8702,N_3719,N_5907);
xor U8703 (N_8703,N_3625,N_5066);
xor U8704 (N_8704,N_4221,N_5894);
or U8705 (N_8705,N_3859,N_6076);
or U8706 (N_8706,N_4982,N_4692);
nand U8707 (N_8707,N_3626,N_3135);
xnor U8708 (N_8708,N_4450,N_4399);
nand U8709 (N_8709,N_4389,N_5975);
nand U8710 (N_8710,N_4538,N_5049);
nor U8711 (N_8711,N_3731,N_4699);
nor U8712 (N_8712,N_4959,N_5185);
nand U8713 (N_8713,N_5593,N_3900);
nor U8714 (N_8714,N_5155,N_4581);
and U8715 (N_8715,N_4897,N_3218);
and U8716 (N_8716,N_3483,N_5345);
and U8717 (N_8717,N_3392,N_4785);
nand U8718 (N_8718,N_5314,N_3522);
xor U8719 (N_8719,N_6144,N_4275);
xnor U8720 (N_8720,N_3251,N_4919);
nand U8721 (N_8721,N_4386,N_3541);
nand U8722 (N_8722,N_3252,N_4158);
xor U8723 (N_8723,N_4355,N_4714);
or U8724 (N_8724,N_4337,N_5695);
and U8725 (N_8725,N_5706,N_5933);
and U8726 (N_8726,N_3758,N_3591);
and U8727 (N_8727,N_4921,N_5753);
and U8728 (N_8728,N_3992,N_3434);
nor U8729 (N_8729,N_4126,N_3871);
nor U8730 (N_8730,N_4068,N_3353);
and U8731 (N_8731,N_3609,N_4758);
and U8732 (N_8732,N_3746,N_3219);
or U8733 (N_8733,N_5418,N_3813);
xnor U8734 (N_8734,N_5355,N_3510);
or U8735 (N_8735,N_5613,N_5573);
or U8736 (N_8736,N_3929,N_4722);
xor U8737 (N_8737,N_5160,N_3204);
nand U8738 (N_8738,N_5509,N_5129);
nor U8739 (N_8739,N_3736,N_5326);
xor U8740 (N_8740,N_5107,N_3314);
nand U8741 (N_8741,N_6109,N_4772);
and U8742 (N_8742,N_3656,N_5430);
xor U8743 (N_8743,N_4285,N_4086);
and U8744 (N_8744,N_5788,N_3995);
nand U8745 (N_8745,N_5380,N_3858);
nor U8746 (N_8746,N_3271,N_5819);
xnor U8747 (N_8747,N_4843,N_5939);
nand U8748 (N_8748,N_4886,N_3938);
nor U8749 (N_8749,N_6087,N_3941);
nand U8750 (N_8750,N_6016,N_3361);
and U8751 (N_8751,N_3898,N_4613);
and U8752 (N_8752,N_6172,N_3215);
and U8753 (N_8753,N_4492,N_3405);
nand U8754 (N_8754,N_3822,N_5129);
nor U8755 (N_8755,N_4971,N_4654);
xor U8756 (N_8756,N_4674,N_5479);
nor U8757 (N_8757,N_4614,N_5824);
nand U8758 (N_8758,N_3813,N_3540);
nor U8759 (N_8759,N_3876,N_5219);
or U8760 (N_8760,N_5702,N_4689);
and U8761 (N_8761,N_4289,N_5643);
nor U8762 (N_8762,N_3434,N_5132);
nand U8763 (N_8763,N_3696,N_4601);
and U8764 (N_8764,N_3236,N_4109);
nor U8765 (N_8765,N_4278,N_5050);
and U8766 (N_8766,N_4970,N_5540);
and U8767 (N_8767,N_3517,N_4923);
or U8768 (N_8768,N_4561,N_4851);
or U8769 (N_8769,N_3470,N_5952);
and U8770 (N_8770,N_5828,N_6139);
or U8771 (N_8771,N_6038,N_4849);
nor U8772 (N_8772,N_3550,N_6068);
nor U8773 (N_8773,N_3174,N_6173);
nand U8774 (N_8774,N_3448,N_5525);
nand U8775 (N_8775,N_6058,N_5323);
xnor U8776 (N_8776,N_5972,N_3166);
nor U8777 (N_8777,N_5665,N_5937);
and U8778 (N_8778,N_5313,N_5774);
nand U8779 (N_8779,N_4255,N_5379);
and U8780 (N_8780,N_5304,N_6059);
nand U8781 (N_8781,N_4900,N_5498);
and U8782 (N_8782,N_5712,N_5518);
or U8783 (N_8783,N_5278,N_3533);
or U8784 (N_8784,N_5433,N_4159);
and U8785 (N_8785,N_4804,N_4284);
or U8786 (N_8786,N_5750,N_5771);
and U8787 (N_8787,N_5949,N_4497);
xnor U8788 (N_8788,N_4455,N_3949);
or U8789 (N_8789,N_5321,N_5758);
nor U8790 (N_8790,N_4206,N_5248);
nand U8791 (N_8791,N_6134,N_4670);
or U8792 (N_8792,N_5018,N_3964);
and U8793 (N_8793,N_5325,N_4205);
and U8794 (N_8794,N_4688,N_4982);
xnor U8795 (N_8795,N_4307,N_3983);
nor U8796 (N_8796,N_4724,N_5332);
nand U8797 (N_8797,N_5427,N_3354);
nand U8798 (N_8798,N_5236,N_5682);
xor U8799 (N_8799,N_5992,N_4547);
nand U8800 (N_8800,N_3293,N_6091);
nor U8801 (N_8801,N_4810,N_6051);
and U8802 (N_8802,N_4702,N_4049);
nor U8803 (N_8803,N_3302,N_3515);
and U8804 (N_8804,N_4111,N_5234);
and U8805 (N_8805,N_4002,N_5311);
or U8806 (N_8806,N_3825,N_3254);
or U8807 (N_8807,N_3620,N_3632);
nand U8808 (N_8808,N_3817,N_5864);
or U8809 (N_8809,N_3906,N_4789);
nor U8810 (N_8810,N_3826,N_5739);
xor U8811 (N_8811,N_5314,N_3450);
xnor U8812 (N_8812,N_5669,N_3947);
xnor U8813 (N_8813,N_4228,N_3870);
and U8814 (N_8814,N_3236,N_3269);
nor U8815 (N_8815,N_3392,N_4460);
and U8816 (N_8816,N_6124,N_5796);
nor U8817 (N_8817,N_5786,N_5005);
xor U8818 (N_8818,N_3638,N_4093);
xnor U8819 (N_8819,N_3373,N_3411);
and U8820 (N_8820,N_6236,N_5969);
and U8821 (N_8821,N_3272,N_5480);
or U8822 (N_8822,N_5915,N_3209);
or U8823 (N_8823,N_5239,N_3356);
nand U8824 (N_8824,N_4393,N_3254);
nor U8825 (N_8825,N_6217,N_3364);
or U8826 (N_8826,N_4655,N_4844);
xor U8827 (N_8827,N_3183,N_5325);
nor U8828 (N_8828,N_5556,N_5926);
or U8829 (N_8829,N_3272,N_4783);
nand U8830 (N_8830,N_4618,N_6195);
or U8831 (N_8831,N_3704,N_3815);
nor U8832 (N_8832,N_3717,N_5313);
nor U8833 (N_8833,N_5788,N_4335);
and U8834 (N_8834,N_3607,N_4625);
or U8835 (N_8835,N_4155,N_3295);
xnor U8836 (N_8836,N_4027,N_3351);
and U8837 (N_8837,N_6079,N_4411);
and U8838 (N_8838,N_4394,N_3903);
or U8839 (N_8839,N_3365,N_5185);
nand U8840 (N_8840,N_4737,N_4910);
xnor U8841 (N_8841,N_5600,N_3845);
xnor U8842 (N_8842,N_3355,N_3963);
nor U8843 (N_8843,N_4090,N_5859);
xor U8844 (N_8844,N_4670,N_3730);
and U8845 (N_8845,N_5549,N_4098);
xnor U8846 (N_8846,N_5445,N_5183);
nand U8847 (N_8847,N_5831,N_5080);
nand U8848 (N_8848,N_4900,N_4137);
or U8849 (N_8849,N_4924,N_3691);
and U8850 (N_8850,N_4711,N_4863);
or U8851 (N_8851,N_4830,N_5142);
or U8852 (N_8852,N_3873,N_4552);
nand U8853 (N_8853,N_4580,N_4684);
and U8854 (N_8854,N_3875,N_6049);
nor U8855 (N_8855,N_4493,N_4745);
xor U8856 (N_8856,N_4839,N_5305);
or U8857 (N_8857,N_5560,N_4121);
or U8858 (N_8858,N_5557,N_3641);
nand U8859 (N_8859,N_5539,N_5063);
nand U8860 (N_8860,N_3787,N_3271);
nor U8861 (N_8861,N_4030,N_3496);
nand U8862 (N_8862,N_5061,N_5554);
xnor U8863 (N_8863,N_3317,N_6146);
and U8864 (N_8864,N_4253,N_6176);
nand U8865 (N_8865,N_4981,N_3534);
nor U8866 (N_8866,N_4420,N_4430);
xnor U8867 (N_8867,N_4634,N_4107);
or U8868 (N_8868,N_6031,N_6057);
or U8869 (N_8869,N_4909,N_3804);
nand U8870 (N_8870,N_4140,N_3625);
xor U8871 (N_8871,N_6051,N_5154);
nand U8872 (N_8872,N_4012,N_3818);
nor U8873 (N_8873,N_5631,N_4593);
nand U8874 (N_8874,N_6201,N_3168);
and U8875 (N_8875,N_5733,N_4473);
or U8876 (N_8876,N_3909,N_5482);
xor U8877 (N_8877,N_3820,N_4453);
or U8878 (N_8878,N_4856,N_4652);
or U8879 (N_8879,N_4901,N_3329);
or U8880 (N_8880,N_4347,N_5748);
xor U8881 (N_8881,N_5473,N_4263);
nand U8882 (N_8882,N_4033,N_4350);
and U8883 (N_8883,N_3369,N_4136);
xnor U8884 (N_8884,N_4193,N_5076);
nor U8885 (N_8885,N_4948,N_5849);
or U8886 (N_8886,N_3910,N_3564);
nand U8887 (N_8887,N_4492,N_5330);
or U8888 (N_8888,N_6115,N_3384);
xor U8889 (N_8889,N_3805,N_5921);
nor U8890 (N_8890,N_5471,N_4131);
nand U8891 (N_8891,N_5637,N_4550);
nor U8892 (N_8892,N_5180,N_4219);
and U8893 (N_8893,N_4880,N_4440);
nor U8894 (N_8894,N_5360,N_4251);
and U8895 (N_8895,N_5600,N_4933);
nor U8896 (N_8896,N_3754,N_5495);
xnor U8897 (N_8897,N_5606,N_5504);
and U8898 (N_8898,N_5983,N_4830);
nand U8899 (N_8899,N_5554,N_5814);
and U8900 (N_8900,N_3572,N_5273);
nor U8901 (N_8901,N_5879,N_6030);
nor U8902 (N_8902,N_6009,N_4007);
or U8903 (N_8903,N_5364,N_4283);
and U8904 (N_8904,N_3320,N_6087);
and U8905 (N_8905,N_4378,N_5611);
nor U8906 (N_8906,N_5084,N_6029);
xor U8907 (N_8907,N_4315,N_4467);
xnor U8908 (N_8908,N_3787,N_5088);
nand U8909 (N_8909,N_4587,N_5323);
nor U8910 (N_8910,N_6155,N_3606);
nor U8911 (N_8911,N_5843,N_4034);
xnor U8912 (N_8912,N_4714,N_5780);
or U8913 (N_8913,N_4222,N_5560);
nor U8914 (N_8914,N_4559,N_5845);
nand U8915 (N_8915,N_5560,N_5179);
or U8916 (N_8916,N_4516,N_4896);
and U8917 (N_8917,N_4419,N_5313);
xnor U8918 (N_8918,N_4651,N_4164);
nand U8919 (N_8919,N_5436,N_5006);
nor U8920 (N_8920,N_5932,N_4791);
and U8921 (N_8921,N_5385,N_5054);
nor U8922 (N_8922,N_3696,N_4321);
nor U8923 (N_8923,N_5847,N_6075);
and U8924 (N_8924,N_4201,N_5228);
nand U8925 (N_8925,N_5314,N_5281);
nor U8926 (N_8926,N_5676,N_5927);
nand U8927 (N_8927,N_3269,N_3579);
or U8928 (N_8928,N_6223,N_5377);
or U8929 (N_8929,N_4969,N_5202);
xor U8930 (N_8930,N_3572,N_5621);
xor U8931 (N_8931,N_3613,N_5627);
nand U8932 (N_8932,N_5581,N_4264);
nor U8933 (N_8933,N_3306,N_3294);
nand U8934 (N_8934,N_5052,N_6073);
or U8935 (N_8935,N_3321,N_5156);
or U8936 (N_8936,N_5153,N_6095);
nand U8937 (N_8937,N_6222,N_5686);
nand U8938 (N_8938,N_6115,N_5129);
nor U8939 (N_8939,N_3712,N_5016);
and U8940 (N_8940,N_3701,N_3907);
xor U8941 (N_8941,N_5026,N_3999);
and U8942 (N_8942,N_5897,N_5440);
nor U8943 (N_8943,N_4367,N_4007);
nor U8944 (N_8944,N_5650,N_4760);
nor U8945 (N_8945,N_3758,N_5805);
or U8946 (N_8946,N_5472,N_4792);
or U8947 (N_8947,N_3248,N_4586);
and U8948 (N_8948,N_3495,N_5075);
or U8949 (N_8949,N_6047,N_4907);
xnor U8950 (N_8950,N_5928,N_6088);
nor U8951 (N_8951,N_5206,N_3332);
nor U8952 (N_8952,N_3491,N_4762);
and U8953 (N_8953,N_4642,N_4123);
nand U8954 (N_8954,N_4382,N_3494);
nor U8955 (N_8955,N_3580,N_5987);
nand U8956 (N_8956,N_5531,N_3688);
xnor U8957 (N_8957,N_4498,N_5389);
or U8958 (N_8958,N_5412,N_4404);
nand U8959 (N_8959,N_3399,N_5264);
and U8960 (N_8960,N_5106,N_5863);
xnor U8961 (N_8961,N_5112,N_3433);
nand U8962 (N_8962,N_4032,N_5309);
nor U8963 (N_8963,N_5420,N_4469);
nand U8964 (N_8964,N_5973,N_5440);
and U8965 (N_8965,N_5655,N_5379);
xor U8966 (N_8966,N_5886,N_5706);
nand U8967 (N_8967,N_5529,N_3621);
nor U8968 (N_8968,N_3348,N_5299);
nand U8969 (N_8969,N_4229,N_5329);
nor U8970 (N_8970,N_4556,N_4755);
xnor U8971 (N_8971,N_3428,N_5894);
nand U8972 (N_8972,N_4196,N_5440);
nor U8973 (N_8973,N_4830,N_5429);
or U8974 (N_8974,N_5973,N_4372);
xnor U8975 (N_8975,N_4699,N_4822);
xnor U8976 (N_8976,N_3356,N_4511);
xnor U8977 (N_8977,N_5693,N_4518);
xnor U8978 (N_8978,N_4346,N_3643);
and U8979 (N_8979,N_4139,N_6244);
nand U8980 (N_8980,N_5008,N_5097);
or U8981 (N_8981,N_5214,N_5382);
nand U8982 (N_8982,N_5314,N_3293);
and U8983 (N_8983,N_5309,N_3260);
nor U8984 (N_8984,N_4508,N_4513);
xnor U8985 (N_8985,N_6174,N_5033);
or U8986 (N_8986,N_3691,N_3745);
xnor U8987 (N_8987,N_6156,N_6226);
and U8988 (N_8988,N_3613,N_3403);
xnor U8989 (N_8989,N_4866,N_5158);
and U8990 (N_8990,N_3255,N_5136);
nor U8991 (N_8991,N_3785,N_5131);
or U8992 (N_8992,N_4370,N_6216);
nor U8993 (N_8993,N_5324,N_4540);
xnor U8994 (N_8994,N_6186,N_5985);
nor U8995 (N_8995,N_3273,N_3492);
and U8996 (N_8996,N_3489,N_5344);
xor U8997 (N_8997,N_4611,N_5369);
nand U8998 (N_8998,N_3707,N_5720);
xor U8999 (N_8999,N_5051,N_4514);
and U9000 (N_9000,N_5262,N_5671);
or U9001 (N_9001,N_3236,N_3978);
nor U9002 (N_9002,N_5135,N_5823);
or U9003 (N_9003,N_4025,N_4453);
or U9004 (N_9004,N_4054,N_4942);
and U9005 (N_9005,N_4222,N_5129);
xor U9006 (N_9006,N_5293,N_4888);
xor U9007 (N_9007,N_4245,N_5093);
or U9008 (N_9008,N_3747,N_4273);
nand U9009 (N_9009,N_6020,N_3187);
xor U9010 (N_9010,N_5974,N_4751);
or U9011 (N_9011,N_5471,N_4432);
or U9012 (N_9012,N_6082,N_4733);
or U9013 (N_9013,N_5397,N_4301);
nor U9014 (N_9014,N_5379,N_4696);
or U9015 (N_9015,N_5974,N_6094);
nand U9016 (N_9016,N_5938,N_3587);
nand U9017 (N_9017,N_3993,N_5718);
xnor U9018 (N_9018,N_5829,N_5298);
nand U9019 (N_9019,N_3347,N_3832);
nor U9020 (N_9020,N_4630,N_3404);
or U9021 (N_9021,N_4931,N_5689);
nor U9022 (N_9022,N_6094,N_3837);
xor U9023 (N_9023,N_4175,N_5405);
and U9024 (N_9024,N_4258,N_3411);
nand U9025 (N_9025,N_5495,N_5462);
and U9026 (N_9026,N_5972,N_4994);
nor U9027 (N_9027,N_4521,N_5620);
xnor U9028 (N_9028,N_5739,N_4001);
and U9029 (N_9029,N_3198,N_5733);
or U9030 (N_9030,N_5297,N_5223);
xor U9031 (N_9031,N_5183,N_5594);
xnor U9032 (N_9032,N_3506,N_5311);
nand U9033 (N_9033,N_3564,N_4878);
and U9034 (N_9034,N_5843,N_5393);
xor U9035 (N_9035,N_3790,N_5207);
nor U9036 (N_9036,N_3473,N_4195);
or U9037 (N_9037,N_5107,N_3591);
or U9038 (N_9038,N_5558,N_5426);
nand U9039 (N_9039,N_5549,N_4649);
and U9040 (N_9040,N_3328,N_5218);
xor U9041 (N_9041,N_4837,N_5465);
and U9042 (N_9042,N_3392,N_3460);
nor U9043 (N_9043,N_4365,N_4840);
and U9044 (N_9044,N_4399,N_3306);
xnor U9045 (N_9045,N_5437,N_5180);
nor U9046 (N_9046,N_4281,N_5308);
nand U9047 (N_9047,N_3800,N_3791);
or U9048 (N_9048,N_5508,N_5249);
or U9049 (N_9049,N_3818,N_5055);
and U9050 (N_9050,N_5673,N_5435);
nor U9051 (N_9051,N_4144,N_4814);
nor U9052 (N_9052,N_3456,N_5155);
or U9053 (N_9053,N_5008,N_5384);
or U9054 (N_9054,N_4562,N_4889);
nand U9055 (N_9055,N_4658,N_5721);
nand U9056 (N_9056,N_3286,N_5285);
nor U9057 (N_9057,N_3455,N_5575);
nor U9058 (N_9058,N_5236,N_5205);
or U9059 (N_9059,N_5818,N_5528);
xor U9060 (N_9060,N_3820,N_4326);
and U9061 (N_9061,N_5423,N_4203);
or U9062 (N_9062,N_5350,N_5178);
xnor U9063 (N_9063,N_5380,N_3542);
or U9064 (N_9064,N_5159,N_4046);
nor U9065 (N_9065,N_6008,N_3584);
and U9066 (N_9066,N_4409,N_4569);
nand U9067 (N_9067,N_5577,N_6056);
and U9068 (N_9068,N_3429,N_5484);
and U9069 (N_9069,N_5343,N_3324);
xor U9070 (N_9070,N_4081,N_5285);
nor U9071 (N_9071,N_5124,N_5173);
nand U9072 (N_9072,N_4206,N_3172);
or U9073 (N_9073,N_5724,N_4039);
and U9074 (N_9074,N_4560,N_3885);
nand U9075 (N_9075,N_4821,N_5153);
nand U9076 (N_9076,N_4459,N_5790);
and U9077 (N_9077,N_6118,N_6223);
nand U9078 (N_9078,N_5765,N_5766);
nor U9079 (N_9079,N_6107,N_4154);
nand U9080 (N_9080,N_3211,N_4539);
nand U9081 (N_9081,N_4867,N_3314);
nor U9082 (N_9082,N_3249,N_4077);
and U9083 (N_9083,N_3682,N_5315);
nor U9084 (N_9084,N_3271,N_5588);
and U9085 (N_9085,N_3848,N_4661);
nor U9086 (N_9086,N_6186,N_5291);
xnor U9087 (N_9087,N_4282,N_5802);
nor U9088 (N_9088,N_5135,N_4740);
or U9089 (N_9089,N_4829,N_5929);
or U9090 (N_9090,N_4623,N_4275);
nor U9091 (N_9091,N_5321,N_5118);
nor U9092 (N_9092,N_3279,N_6200);
and U9093 (N_9093,N_5260,N_5688);
xor U9094 (N_9094,N_3439,N_5386);
and U9095 (N_9095,N_6157,N_5300);
or U9096 (N_9096,N_5376,N_4123);
xnor U9097 (N_9097,N_5184,N_3968);
nand U9098 (N_9098,N_6046,N_5405);
nor U9099 (N_9099,N_4835,N_4395);
xnor U9100 (N_9100,N_5906,N_3347);
nand U9101 (N_9101,N_5942,N_3245);
and U9102 (N_9102,N_5538,N_4285);
nor U9103 (N_9103,N_4867,N_5300);
nand U9104 (N_9104,N_4207,N_3667);
nor U9105 (N_9105,N_3848,N_5212);
and U9106 (N_9106,N_5627,N_6003);
and U9107 (N_9107,N_6233,N_3587);
xor U9108 (N_9108,N_6021,N_5589);
nor U9109 (N_9109,N_5545,N_6004);
or U9110 (N_9110,N_3357,N_4170);
nand U9111 (N_9111,N_3163,N_6174);
nor U9112 (N_9112,N_5878,N_4074);
nor U9113 (N_9113,N_5582,N_5836);
or U9114 (N_9114,N_4598,N_5232);
or U9115 (N_9115,N_4139,N_4798);
xor U9116 (N_9116,N_3755,N_6212);
or U9117 (N_9117,N_5516,N_5639);
nor U9118 (N_9118,N_4973,N_3616);
nand U9119 (N_9119,N_4644,N_4171);
xnor U9120 (N_9120,N_5287,N_3587);
and U9121 (N_9121,N_3344,N_4266);
or U9122 (N_9122,N_6038,N_3655);
or U9123 (N_9123,N_3319,N_6116);
or U9124 (N_9124,N_5938,N_3579);
nand U9125 (N_9125,N_3540,N_3576);
nand U9126 (N_9126,N_5636,N_5878);
nand U9127 (N_9127,N_5008,N_5630);
nor U9128 (N_9128,N_6096,N_3661);
nand U9129 (N_9129,N_5983,N_4065);
nand U9130 (N_9130,N_5679,N_4513);
or U9131 (N_9131,N_4493,N_3195);
xnor U9132 (N_9132,N_4957,N_3587);
nor U9133 (N_9133,N_3972,N_4706);
nand U9134 (N_9134,N_5204,N_3326);
nor U9135 (N_9135,N_4462,N_3134);
xor U9136 (N_9136,N_5819,N_5593);
nand U9137 (N_9137,N_5279,N_3254);
nand U9138 (N_9138,N_6188,N_5192);
nor U9139 (N_9139,N_3845,N_3473);
and U9140 (N_9140,N_5897,N_6094);
or U9141 (N_9141,N_5432,N_3163);
nand U9142 (N_9142,N_5402,N_4401);
nor U9143 (N_9143,N_3748,N_3227);
and U9144 (N_9144,N_5583,N_6055);
or U9145 (N_9145,N_3704,N_4311);
and U9146 (N_9146,N_3335,N_3781);
nor U9147 (N_9147,N_4697,N_4582);
xnor U9148 (N_9148,N_3321,N_4078);
and U9149 (N_9149,N_3712,N_3446);
and U9150 (N_9150,N_4060,N_4006);
xor U9151 (N_9151,N_4351,N_3864);
or U9152 (N_9152,N_4285,N_4088);
xor U9153 (N_9153,N_6086,N_3404);
nand U9154 (N_9154,N_5106,N_4613);
xnor U9155 (N_9155,N_3450,N_3157);
and U9156 (N_9156,N_4001,N_5356);
xor U9157 (N_9157,N_4896,N_4707);
nand U9158 (N_9158,N_4937,N_5490);
or U9159 (N_9159,N_4912,N_5411);
xor U9160 (N_9160,N_4250,N_4797);
xor U9161 (N_9161,N_3692,N_4923);
xnor U9162 (N_9162,N_4103,N_3334);
nor U9163 (N_9163,N_3337,N_5636);
or U9164 (N_9164,N_5441,N_4244);
nor U9165 (N_9165,N_4673,N_5696);
nor U9166 (N_9166,N_4461,N_3594);
and U9167 (N_9167,N_4971,N_5224);
or U9168 (N_9168,N_4411,N_5920);
nor U9169 (N_9169,N_5404,N_5971);
nor U9170 (N_9170,N_3959,N_5574);
xor U9171 (N_9171,N_3923,N_3141);
and U9172 (N_9172,N_3758,N_3881);
nand U9173 (N_9173,N_5301,N_4504);
or U9174 (N_9174,N_5490,N_5108);
xor U9175 (N_9175,N_3137,N_5618);
xnor U9176 (N_9176,N_5266,N_4861);
and U9177 (N_9177,N_3182,N_4988);
nand U9178 (N_9178,N_4202,N_4940);
nand U9179 (N_9179,N_3873,N_4382);
xor U9180 (N_9180,N_6121,N_5618);
and U9181 (N_9181,N_6092,N_4900);
nand U9182 (N_9182,N_5747,N_5715);
xnor U9183 (N_9183,N_5180,N_4258);
xnor U9184 (N_9184,N_3915,N_6176);
or U9185 (N_9185,N_5537,N_5569);
or U9186 (N_9186,N_3523,N_5568);
nor U9187 (N_9187,N_5607,N_4681);
or U9188 (N_9188,N_5447,N_5276);
nand U9189 (N_9189,N_5896,N_4736);
nand U9190 (N_9190,N_4372,N_3892);
nand U9191 (N_9191,N_3936,N_3235);
nor U9192 (N_9192,N_5709,N_5916);
nand U9193 (N_9193,N_3426,N_4658);
or U9194 (N_9194,N_5756,N_4418);
or U9195 (N_9195,N_6038,N_4386);
xor U9196 (N_9196,N_4433,N_3524);
nand U9197 (N_9197,N_6136,N_3367);
nor U9198 (N_9198,N_5082,N_5337);
xor U9199 (N_9199,N_5305,N_3446);
and U9200 (N_9200,N_5419,N_3708);
xnor U9201 (N_9201,N_4752,N_3864);
nor U9202 (N_9202,N_4251,N_5113);
or U9203 (N_9203,N_4909,N_5081);
nand U9204 (N_9204,N_4418,N_3851);
and U9205 (N_9205,N_5646,N_4406);
and U9206 (N_9206,N_3735,N_5672);
nand U9207 (N_9207,N_5220,N_5136);
xnor U9208 (N_9208,N_5080,N_3231);
or U9209 (N_9209,N_4465,N_5288);
xnor U9210 (N_9210,N_5344,N_5472);
or U9211 (N_9211,N_4539,N_3971);
and U9212 (N_9212,N_3534,N_5872);
nand U9213 (N_9213,N_5683,N_4099);
and U9214 (N_9214,N_6197,N_5149);
nor U9215 (N_9215,N_3725,N_3917);
and U9216 (N_9216,N_4678,N_3209);
nor U9217 (N_9217,N_3181,N_3993);
or U9218 (N_9218,N_3242,N_5425);
and U9219 (N_9219,N_6149,N_5710);
or U9220 (N_9220,N_5801,N_6177);
or U9221 (N_9221,N_4957,N_3773);
nand U9222 (N_9222,N_4416,N_5572);
and U9223 (N_9223,N_3998,N_5343);
or U9224 (N_9224,N_3479,N_5356);
xor U9225 (N_9225,N_3773,N_3252);
nor U9226 (N_9226,N_4951,N_3141);
or U9227 (N_9227,N_5169,N_3302);
nor U9228 (N_9228,N_4598,N_4331);
and U9229 (N_9229,N_3345,N_4825);
nor U9230 (N_9230,N_5124,N_4907);
nand U9231 (N_9231,N_3996,N_4737);
nand U9232 (N_9232,N_5970,N_4068);
xnor U9233 (N_9233,N_3438,N_3153);
nand U9234 (N_9234,N_4934,N_4685);
xor U9235 (N_9235,N_5532,N_5206);
nor U9236 (N_9236,N_3155,N_5771);
nand U9237 (N_9237,N_3152,N_4195);
nand U9238 (N_9238,N_3663,N_4469);
and U9239 (N_9239,N_4311,N_4894);
and U9240 (N_9240,N_4156,N_5024);
and U9241 (N_9241,N_4600,N_5777);
nor U9242 (N_9242,N_5472,N_5140);
or U9243 (N_9243,N_5358,N_6103);
or U9244 (N_9244,N_4042,N_5024);
nor U9245 (N_9245,N_5122,N_6244);
nor U9246 (N_9246,N_3333,N_5785);
or U9247 (N_9247,N_3626,N_5418);
and U9248 (N_9248,N_5301,N_4708);
xor U9249 (N_9249,N_4903,N_4583);
nor U9250 (N_9250,N_3539,N_6207);
nand U9251 (N_9251,N_3635,N_5197);
nand U9252 (N_9252,N_3695,N_4949);
nor U9253 (N_9253,N_3604,N_4791);
nand U9254 (N_9254,N_6233,N_4096);
nor U9255 (N_9255,N_6020,N_5139);
and U9256 (N_9256,N_5275,N_4942);
nand U9257 (N_9257,N_6036,N_3952);
nand U9258 (N_9258,N_3952,N_3904);
nor U9259 (N_9259,N_5386,N_4451);
and U9260 (N_9260,N_4318,N_5262);
nand U9261 (N_9261,N_6047,N_5770);
nand U9262 (N_9262,N_3574,N_5973);
nand U9263 (N_9263,N_5454,N_5583);
or U9264 (N_9264,N_3935,N_3927);
nor U9265 (N_9265,N_3861,N_4639);
xor U9266 (N_9266,N_5248,N_5797);
nor U9267 (N_9267,N_5500,N_5645);
nand U9268 (N_9268,N_3881,N_5153);
nor U9269 (N_9269,N_4222,N_3995);
or U9270 (N_9270,N_5034,N_4182);
nor U9271 (N_9271,N_3910,N_3715);
xor U9272 (N_9272,N_4843,N_4940);
and U9273 (N_9273,N_3522,N_3589);
and U9274 (N_9274,N_5737,N_4903);
nor U9275 (N_9275,N_3888,N_4496);
xor U9276 (N_9276,N_4954,N_4587);
and U9277 (N_9277,N_3380,N_4997);
and U9278 (N_9278,N_5889,N_4088);
nand U9279 (N_9279,N_5983,N_4685);
nor U9280 (N_9280,N_3471,N_3714);
and U9281 (N_9281,N_4429,N_6083);
and U9282 (N_9282,N_5783,N_4533);
nand U9283 (N_9283,N_5453,N_3310);
and U9284 (N_9284,N_4350,N_3188);
nor U9285 (N_9285,N_5199,N_3200);
nor U9286 (N_9286,N_5929,N_5845);
nand U9287 (N_9287,N_5157,N_3861);
nor U9288 (N_9288,N_4365,N_4800);
or U9289 (N_9289,N_4592,N_5453);
nor U9290 (N_9290,N_3395,N_3766);
and U9291 (N_9291,N_5551,N_3915);
xnor U9292 (N_9292,N_5353,N_4719);
or U9293 (N_9293,N_5097,N_4505);
nand U9294 (N_9294,N_5789,N_5512);
and U9295 (N_9295,N_3713,N_4807);
xnor U9296 (N_9296,N_5887,N_5420);
nor U9297 (N_9297,N_3753,N_3953);
nand U9298 (N_9298,N_5473,N_3945);
xor U9299 (N_9299,N_4139,N_4172);
nor U9300 (N_9300,N_5387,N_4440);
or U9301 (N_9301,N_4014,N_5812);
nand U9302 (N_9302,N_5404,N_5273);
or U9303 (N_9303,N_4978,N_5376);
or U9304 (N_9304,N_3540,N_4327);
and U9305 (N_9305,N_3745,N_4630);
xor U9306 (N_9306,N_3972,N_3533);
nand U9307 (N_9307,N_4899,N_3438);
xnor U9308 (N_9308,N_5420,N_4744);
nor U9309 (N_9309,N_4216,N_5521);
or U9310 (N_9310,N_5601,N_3874);
nor U9311 (N_9311,N_4970,N_4186);
or U9312 (N_9312,N_5590,N_3671);
or U9313 (N_9313,N_4584,N_3834);
or U9314 (N_9314,N_5863,N_4439);
nor U9315 (N_9315,N_4398,N_5638);
nand U9316 (N_9316,N_6219,N_4600);
nand U9317 (N_9317,N_3371,N_3713);
xnor U9318 (N_9318,N_6024,N_5932);
or U9319 (N_9319,N_5538,N_5559);
xnor U9320 (N_9320,N_5483,N_3857);
and U9321 (N_9321,N_3902,N_4914);
xnor U9322 (N_9322,N_3763,N_4941);
nor U9323 (N_9323,N_3959,N_5358);
nand U9324 (N_9324,N_4490,N_3187);
nor U9325 (N_9325,N_6043,N_4590);
xnor U9326 (N_9326,N_6104,N_3401);
or U9327 (N_9327,N_4012,N_3526);
nor U9328 (N_9328,N_5701,N_3188);
and U9329 (N_9329,N_3879,N_3965);
and U9330 (N_9330,N_4127,N_4749);
nor U9331 (N_9331,N_4498,N_4721);
and U9332 (N_9332,N_3228,N_4867);
nor U9333 (N_9333,N_5856,N_4324);
nor U9334 (N_9334,N_4215,N_3415);
or U9335 (N_9335,N_3246,N_5992);
xor U9336 (N_9336,N_5549,N_5461);
and U9337 (N_9337,N_5408,N_4393);
nand U9338 (N_9338,N_5056,N_3153);
and U9339 (N_9339,N_3181,N_4941);
or U9340 (N_9340,N_4502,N_3324);
or U9341 (N_9341,N_5122,N_4651);
or U9342 (N_9342,N_3433,N_3987);
nand U9343 (N_9343,N_5270,N_4780);
nand U9344 (N_9344,N_3255,N_4690);
xnor U9345 (N_9345,N_6136,N_4497);
nand U9346 (N_9346,N_5760,N_3814);
nand U9347 (N_9347,N_3502,N_6112);
or U9348 (N_9348,N_5380,N_4516);
or U9349 (N_9349,N_5010,N_4125);
or U9350 (N_9350,N_3413,N_6235);
and U9351 (N_9351,N_4034,N_4491);
nand U9352 (N_9352,N_3998,N_6142);
nor U9353 (N_9353,N_5083,N_4012);
nor U9354 (N_9354,N_3260,N_4797);
xor U9355 (N_9355,N_3364,N_4220);
or U9356 (N_9356,N_3641,N_5181);
xor U9357 (N_9357,N_6040,N_6063);
and U9358 (N_9358,N_4891,N_3701);
or U9359 (N_9359,N_6222,N_4165);
and U9360 (N_9360,N_5095,N_3946);
or U9361 (N_9361,N_5904,N_3954);
nand U9362 (N_9362,N_5471,N_5068);
nand U9363 (N_9363,N_5479,N_3869);
xor U9364 (N_9364,N_3804,N_5121);
or U9365 (N_9365,N_4942,N_4204);
xor U9366 (N_9366,N_4145,N_5382);
nor U9367 (N_9367,N_4748,N_3567);
nand U9368 (N_9368,N_5680,N_4214);
xor U9369 (N_9369,N_5368,N_3802);
xnor U9370 (N_9370,N_4189,N_5336);
nor U9371 (N_9371,N_5647,N_5095);
nor U9372 (N_9372,N_3438,N_4071);
xnor U9373 (N_9373,N_5471,N_5310);
or U9374 (N_9374,N_5048,N_5565);
and U9375 (N_9375,N_6557,N_6829);
nor U9376 (N_9376,N_6635,N_6296);
nor U9377 (N_9377,N_8569,N_8909);
and U9378 (N_9378,N_8166,N_6560);
nand U9379 (N_9379,N_6492,N_6422);
or U9380 (N_9380,N_9141,N_8000);
nor U9381 (N_9381,N_7790,N_7216);
xnor U9382 (N_9382,N_8769,N_7448);
nor U9383 (N_9383,N_8915,N_8177);
or U9384 (N_9384,N_6441,N_6938);
xnor U9385 (N_9385,N_6715,N_6723);
nand U9386 (N_9386,N_6523,N_9190);
and U9387 (N_9387,N_7999,N_8237);
or U9388 (N_9388,N_7012,N_6291);
and U9389 (N_9389,N_8581,N_8115);
xnor U9390 (N_9390,N_9068,N_9136);
xnor U9391 (N_9391,N_7891,N_9284);
nand U9392 (N_9392,N_9101,N_7478);
or U9393 (N_9393,N_8524,N_7146);
or U9394 (N_9394,N_8351,N_9123);
or U9395 (N_9395,N_6538,N_7271);
nor U9396 (N_9396,N_8251,N_6848);
and U9397 (N_9397,N_6720,N_7415);
nor U9398 (N_9398,N_6596,N_8656);
xnor U9399 (N_9399,N_8650,N_7477);
nor U9400 (N_9400,N_6565,N_8389);
nor U9401 (N_9401,N_7578,N_6937);
and U9402 (N_9402,N_9307,N_6475);
nand U9403 (N_9403,N_7688,N_6782);
and U9404 (N_9404,N_6924,N_6618);
or U9405 (N_9405,N_6373,N_9134);
nor U9406 (N_9406,N_6571,N_7876);
and U9407 (N_9407,N_7858,N_9237);
nor U9408 (N_9408,N_7436,N_7453);
xnor U9409 (N_9409,N_8175,N_8978);
xor U9410 (N_9410,N_7276,N_8357);
and U9411 (N_9411,N_6554,N_6935);
and U9412 (N_9412,N_7340,N_9099);
xnor U9413 (N_9413,N_6941,N_9130);
xnor U9414 (N_9414,N_9162,N_9070);
nand U9415 (N_9415,N_9370,N_8970);
nor U9416 (N_9416,N_7615,N_8813);
and U9417 (N_9417,N_9100,N_7856);
and U9418 (N_9418,N_7614,N_7768);
xor U9419 (N_9419,N_6709,N_7752);
nor U9420 (N_9420,N_8655,N_7665);
and U9421 (N_9421,N_9183,N_7230);
nor U9422 (N_9422,N_8661,N_9102);
nand U9423 (N_9423,N_7612,N_7016);
nand U9424 (N_9424,N_7729,N_6951);
xnor U9425 (N_9425,N_7481,N_9228);
xor U9426 (N_9426,N_7795,N_6402);
nand U9427 (N_9427,N_6983,N_6408);
or U9428 (N_9428,N_8510,N_9327);
xor U9429 (N_9429,N_7906,N_7849);
nand U9430 (N_9430,N_7402,N_8766);
nor U9431 (N_9431,N_7308,N_7474);
and U9432 (N_9432,N_6790,N_6696);
nor U9433 (N_9433,N_7541,N_9089);
and U9434 (N_9434,N_7242,N_6477);
nand U9435 (N_9435,N_7452,N_7869);
or U9436 (N_9436,N_7324,N_9251);
nor U9437 (N_9437,N_8875,N_7489);
nand U9438 (N_9438,N_7420,N_8490);
nand U9439 (N_9439,N_6687,N_6942);
nand U9440 (N_9440,N_6359,N_6777);
nor U9441 (N_9441,N_8937,N_6494);
nor U9442 (N_9442,N_8283,N_7401);
and U9443 (N_9443,N_6989,N_6621);
xnor U9444 (N_9444,N_7585,N_8538);
and U9445 (N_9445,N_7034,N_8022);
or U9446 (N_9446,N_8838,N_8688);
xor U9447 (N_9447,N_7653,N_9249);
xor U9448 (N_9448,N_6730,N_6251);
xor U9449 (N_9449,N_7260,N_7766);
xor U9450 (N_9450,N_9244,N_9314);
nand U9451 (N_9451,N_8300,N_8780);
and U9452 (N_9452,N_8025,N_7936);
xor U9453 (N_9453,N_8741,N_8206);
or U9454 (N_9454,N_6774,N_8602);
xnor U9455 (N_9455,N_8028,N_8527);
xnor U9456 (N_9456,N_6916,N_6310);
or U9457 (N_9457,N_9172,N_8094);
or U9458 (N_9458,N_6614,N_8042);
and U9459 (N_9459,N_7123,N_6511);
nor U9460 (N_9460,N_7218,N_7113);
and U9461 (N_9461,N_7093,N_8522);
or U9462 (N_9462,N_9337,N_8111);
nor U9463 (N_9463,N_8185,N_6431);
or U9464 (N_9464,N_7544,N_8667);
nand U9465 (N_9465,N_7832,N_9185);
nand U9466 (N_9466,N_7997,N_8020);
xor U9467 (N_9467,N_8475,N_8248);
nor U9468 (N_9468,N_7721,N_9230);
and U9469 (N_9469,N_8267,N_7964);
or U9470 (N_9470,N_8823,N_6481);
nor U9471 (N_9471,N_8224,N_7560);
or U9472 (N_9472,N_6800,N_9161);
and U9473 (N_9473,N_6946,N_7442);
xor U9474 (N_9474,N_8596,N_8827);
xnor U9475 (N_9475,N_7470,N_8165);
nor U9476 (N_9476,N_7839,N_7536);
xor U9477 (N_9477,N_6595,N_7433);
xnor U9478 (N_9478,N_8247,N_7733);
nand U9479 (N_9479,N_7460,N_8414);
or U9480 (N_9480,N_7645,N_6430);
nand U9481 (N_9481,N_9084,N_8200);
nor U9482 (N_9482,N_8988,N_6284);
xor U9483 (N_9483,N_8782,N_6742);
nor U9484 (N_9484,N_6352,N_6269);
and U9485 (N_9485,N_6954,N_7755);
or U9486 (N_9486,N_8545,N_8217);
nand U9487 (N_9487,N_9143,N_6758);
or U9488 (N_9488,N_6378,N_8412);
or U9489 (N_9489,N_7026,N_8822);
or U9490 (N_9490,N_7746,N_8256);
nor U9491 (N_9491,N_7138,N_7055);
and U9492 (N_9492,N_7728,N_8019);
or U9493 (N_9493,N_8274,N_7919);
or U9494 (N_9494,N_6889,N_6690);
nor U9495 (N_9495,N_7036,N_8726);
and U9496 (N_9496,N_6705,N_8110);
nor U9497 (N_9497,N_8755,N_7791);
xnor U9498 (N_9498,N_7343,N_8464);
and U9499 (N_9499,N_6607,N_9202);
xor U9500 (N_9500,N_6905,N_7675);
and U9501 (N_9501,N_8621,N_8039);
nor U9502 (N_9502,N_6823,N_8333);
or U9503 (N_9503,N_8506,N_7457);
or U9504 (N_9504,N_6520,N_8393);
nand U9505 (N_9505,N_9242,N_6780);
or U9506 (N_9506,N_7062,N_7852);
xnor U9507 (N_9507,N_7387,N_8745);
nand U9508 (N_9508,N_9164,N_6473);
nor U9509 (N_9509,N_6318,N_8752);
nor U9510 (N_9510,N_8530,N_6336);
nand U9511 (N_9511,N_8117,N_9177);
and U9512 (N_9512,N_7185,N_6770);
and U9513 (N_9513,N_9279,N_7792);
xor U9514 (N_9514,N_9232,N_7559);
nand U9515 (N_9515,N_8129,N_6713);
nor U9516 (N_9516,N_7030,N_6645);
xor U9517 (N_9517,N_7043,N_8600);
xor U9518 (N_9518,N_6526,N_7465);
or U9519 (N_9519,N_7933,N_8365);
xor U9520 (N_9520,N_7804,N_7313);
xor U9521 (N_9521,N_8941,N_8724);
nand U9522 (N_9522,N_6587,N_7890);
nand U9523 (N_9523,N_8382,N_7178);
or U9524 (N_9524,N_9306,N_8531);
nand U9525 (N_9525,N_8829,N_7473);
or U9526 (N_9526,N_7732,N_8114);
nor U9527 (N_9527,N_7318,N_9049);
and U9528 (N_9528,N_6399,N_7899);
and U9529 (N_9529,N_9085,N_8555);
xor U9530 (N_9530,N_7667,N_8358);
or U9531 (N_9531,N_9080,N_7562);
nor U9532 (N_9532,N_9151,N_6710);
xor U9533 (N_9533,N_7520,N_8448);
nand U9534 (N_9534,N_6558,N_8196);
xor U9535 (N_9535,N_8372,N_7785);
or U9536 (N_9536,N_6650,N_9153);
or U9537 (N_9537,N_7526,N_8265);
or U9538 (N_9538,N_6641,N_6578);
nand U9539 (N_9539,N_6325,N_8260);
or U9540 (N_9540,N_7683,N_9215);
or U9541 (N_9541,N_7014,N_6451);
and U9542 (N_9542,N_6436,N_8092);
xor U9543 (N_9543,N_6866,N_6302);
nand U9544 (N_9544,N_7846,N_6572);
and U9545 (N_9545,N_8168,N_8164);
nand U9546 (N_9546,N_8669,N_6369);
nor U9547 (N_9547,N_8529,N_8950);
nor U9548 (N_9548,N_6959,N_7788);
xnor U9549 (N_9549,N_7598,N_8367);
nand U9550 (N_9550,N_8904,N_8394);
or U9551 (N_9551,N_6410,N_7820);
and U9552 (N_9552,N_9260,N_8402);
or U9553 (N_9553,N_6366,N_8622);
xnor U9554 (N_9554,N_7987,N_6298);
nand U9555 (N_9555,N_6277,N_8677);
nor U9556 (N_9556,N_7764,N_8613);
and U9557 (N_9557,N_8606,N_9347);
xnor U9558 (N_9558,N_7082,N_8477);
nand U9559 (N_9559,N_7525,N_8913);
nor U9560 (N_9560,N_9131,N_7061);
and U9561 (N_9561,N_7912,N_7961);
nand U9562 (N_9562,N_6750,N_9175);
or U9563 (N_9563,N_8882,N_6737);
nand U9564 (N_9564,N_7747,N_7468);
nand U9565 (N_9565,N_9341,N_7753);
and U9566 (N_9566,N_8582,N_8031);
nor U9567 (N_9567,N_6514,N_7145);
xor U9568 (N_9568,N_7148,N_7704);
nor U9569 (N_9569,N_6842,N_7022);
or U9570 (N_9570,N_8816,N_6348);
xor U9571 (N_9571,N_6839,N_7068);
or U9572 (N_9572,N_8027,N_8630);
nor U9573 (N_9573,N_8681,N_8304);
nor U9574 (N_9574,N_7861,N_9112);
or U9575 (N_9575,N_6948,N_9308);
nor U9576 (N_9576,N_6731,N_7265);
or U9577 (N_9577,N_8002,N_8349);
nor U9578 (N_9578,N_8905,N_7582);
nor U9579 (N_9579,N_8443,N_7505);
xor U9580 (N_9580,N_9047,N_9028);
and U9581 (N_9581,N_9331,N_8705);
nand U9582 (N_9582,N_6341,N_9004);
nor U9583 (N_9583,N_9247,N_7840);
xnor U9584 (N_9584,N_6884,N_7648);
and U9585 (N_9585,N_8936,N_7706);
nor U9586 (N_9586,N_7802,N_8996);
and U9587 (N_9587,N_7736,N_7199);
xnor U9588 (N_9588,N_6552,N_9108);
nand U9589 (N_9589,N_6757,N_9147);
or U9590 (N_9590,N_7893,N_8364);
and U9591 (N_9591,N_6631,N_7639);
and U9592 (N_9592,N_7817,N_9304);
nand U9593 (N_9593,N_8785,N_9142);
and U9594 (N_9594,N_7716,N_7122);
xnor U9595 (N_9595,N_7682,N_7441);
and U9596 (N_9596,N_7603,N_8362);
and U9597 (N_9597,N_6784,N_7118);
nor U9598 (N_9598,N_7794,N_8303);
or U9599 (N_9599,N_8084,N_7715);
nand U9600 (N_9600,N_7516,N_7263);
xnor U9601 (N_9601,N_7257,N_6677);
and U9602 (N_9602,N_8760,N_8878);
and U9603 (N_9603,N_8906,N_6364);
or U9604 (N_9604,N_6575,N_9193);
xnor U9605 (N_9605,N_8733,N_8892);
nand U9606 (N_9606,N_6390,N_6427);
or U9607 (N_9607,N_8809,N_8326);
or U9608 (N_9608,N_7135,N_8979);
nand U9609 (N_9609,N_8654,N_8857);
and U9610 (N_9610,N_7634,N_8439);
xor U9611 (N_9611,N_6400,N_7713);
nand U9612 (N_9612,N_9173,N_8790);
nand U9613 (N_9613,N_7393,N_6796);
and U9614 (N_9614,N_7397,N_9201);
and U9615 (N_9615,N_7835,N_8282);
nor U9616 (N_9616,N_7259,N_8986);
xnor U9617 (N_9617,N_7540,N_6684);
nor U9618 (N_9618,N_8585,N_8016);
or U9619 (N_9619,N_7215,N_6654);
xor U9620 (N_9620,N_6857,N_8750);
or U9621 (N_9621,N_7895,N_8848);
nor U9622 (N_9622,N_8890,N_8102);
nand U9623 (N_9623,N_8231,N_6764);
and U9624 (N_9624,N_7017,N_9007);
nor U9625 (N_9625,N_7142,N_7613);
and U9626 (N_9626,N_8607,N_6998);
nor U9627 (N_9627,N_8471,N_9313);
and U9628 (N_9628,N_8536,N_6890);
xor U9629 (N_9629,N_8280,N_6319);
or U9630 (N_9630,N_8220,N_7357);
and U9631 (N_9631,N_6944,N_7344);
nand U9632 (N_9632,N_7314,N_8948);
nand U9633 (N_9633,N_7815,N_6389);
or U9634 (N_9634,N_8048,N_7002);
xor U9635 (N_9635,N_8170,N_6748);
and U9636 (N_9636,N_6483,N_6426);
nand U9637 (N_9637,N_8526,N_7444);
nand U9638 (N_9638,N_7927,N_6642);
nor U9639 (N_9639,N_8122,N_6980);
nand U9640 (N_9640,N_8850,N_8063);
and U9641 (N_9641,N_6566,N_6556);
nand U9642 (N_9642,N_8145,N_7326);
xnor U9643 (N_9643,N_8325,N_9234);
nand U9644 (N_9644,N_6535,N_6879);
nor U9645 (N_9645,N_8473,N_8077);
nor U9646 (N_9646,N_7623,N_8198);
or U9647 (N_9647,N_8184,N_7480);
nand U9648 (N_9648,N_6920,N_6919);
xor U9649 (N_9649,N_7647,N_9008);
nor U9650 (N_9650,N_9043,N_7696);
xor U9651 (N_9651,N_8884,N_9223);
xnor U9652 (N_9652,N_8873,N_7793);
nor U9653 (N_9653,N_7725,N_7549);
nor U9654 (N_9654,N_8101,N_8043);
and U9655 (N_9655,N_8203,N_9350);
and U9656 (N_9656,N_6733,N_8078);
nor U9657 (N_9657,N_8993,N_7008);
or U9658 (N_9658,N_9252,N_8955);
and U9659 (N_9659,N_9038,N_8381);
xor U9660 (N_9660,N_6599,N_8431);
or U9661 (N_9661,N_8194,N_8479);
or U9662 (N_9662,N_8589,N_8916);
nand U9663 (N_9663,N_7131,N_6855);
xor U9664 (N_9664,N_6409,N_6472);
xnor U9665 (N_9665,N_7984,N_9319);
or U9666 (N_9666,N_7396,N_8371);
nor U9667 (N_9667,N_8587,N_7134);
and U9668 (N_9668,N_7015,N_7312);
nand U9669 (N_9669,N_9066,N_9081);
nand U9670 (N_9670,N_7167,N_7518);
nor U9671 (N_9671,N_9148,N_8710);
xor U9672 (N_9672,N_8434,N_8109);
xor U9673 (N_9673,N_7205,N_7085);
or U9674 (N_9674,N_8449,N_6945);
and U9675 (N_9675,N_8685,N_9297);
xnor U9676 (N_9676,N_8014,N_8794);
nand U9677 (N_9677,N_7405,N_6736);
xnor U9678 (N_9678,N_9034,N_7952);
xor U9679 (N_9679,N_7757,N_6798);
nand U9680 (N_9680,N_6322,N_8962);
xor U9681 (N_9681,N_6491,N_9364);
or U9682 (N_9682,N_7500,N_8007);
and U9683 (N_9683,N_7173,N_6747);
or U9684 (N_9684,N_8923,N_8321);
or U9685 (N_9685,N_6281,N_8968);
and U9686 (N_9686,N_8784,N_8727);
nand U9687 (N_9687,N_7702,N_8824);
xor U9688 (N_9688,N_7574,N_8963);
nor U9689 (N_9689,N_6909,N_8577);
xor U9690 (N_9690,N_8821,N_8008);
nor U9691 (N_9691,N_8953,N_6868);
nor U9692 (N_9692,N_8957,N_9051);
or U9693 (N_9693,N_7070,N_9310);
nand U9694 (N_9694,N_6913,N_9061);
and U9695 (N_9695,N_7970,N_7132);
xnor U9696 (N_9696,N_7154,N_6931);
and U9697 (N_9697,N_6676,N_7864);
nor U9698 (N_9698,N_7718,N_6775);
xnor U9699 (N_9699,N_8843,N_6809);
nand U9700 (N_9700,N_7333,N_7556);
or U9701 (N_9701,N_7749,N_9361);
nand U9702 (N_9702,N_7780,N_6656);
nor U9703 (N_9703,N_6267,N_7954);
nor U9704 (N_9704,N_7141,N_8627);
nor U9705 (N_9705,N_6387,N_7158);
or U9706 (N_9706,N_6679,N_6972);
and U9707 (N_9707,N_9217,N_8480);
xnor U9708 (N_9708,N_7483,N_7310);
and U9709 (N_9709,N_8299,N_7741);
xnor U9710 (N_9710,N_7367,N_6382);
and U9711 (N_9711,N_8751,N_6772);
nand U9712 (N_9712,N_8392,N_8792);
nand U9713 (N_9713,N_6873,N_6285);
nand U9714 (N_9714,N_7059,N_7214);
and U9715 (N_9715,N_6689,N_7922);
and U9716 (N_9716,N_8478,N_8975);
xnor U9717 (N_9717,N_6338,N_8348);
nand U9718 (N_9718,N_6900,N_7910);
nand U9719 (N_9719,N_7924,N_6286);
xnor U9720 (N_9720,N_9285,N_7646);
nor U9721 (N_9721,N_8350,N_7868);
or U9722 (N_9722,N_6957,N_7088);
nand U9723 (N_9723,N_8861,N_7969);
xnor U9724 (N_9724,N_8492,N_8447);
nor U9725 (N_9725,N_8297,N_7399);
or U9726 (N_9726,N_8328,N_7807);
and U9727 (N_9727,N_8868,N_6636);
and U9728 (N_9728,N_7193,N_8052);
or U9729 (N_9729,N_7884,N_9330);
and U9730 (N_9730,N_6647,N_8637);
nand U9731 (N_9731,N_7476,N_7917);
or U9732 (N_9732,N_6693,N_8897);
or U9733 (N_9733,N_6849,N_8659);
nand U9734 (N_9734,N_8097,N_7748);
xnor U9735 (N_9735,N_8099,N_7772);
nor U9736 (N_9736,N_6996,N_7001);
nand U9737 (N_9737,N_8263,N_6425);
xor U9738 (N_9738,N_9082,N_8199);
or U9739 (N_9739,N_7384,N_7903);
nor U9740 (N_9740,N_6643,N_8663);
or U9741 (N_9741,N_8429,N_8773);
nand U9742 (N_9742,N_8812,N_6760);
nand U9743 (N_9743,N_7596,N_8893);
or U9744 (N_9744,N_9255,N_8134);
or U9745 (N_9745,N_7763,N_8635);
nor U9746 (N_9746,N_9261,N_8140);
nor U9747 (N_9747,N_8568,N_8649);
xnor U9748 (N_9748,N_8819,N_7504);
nor U9749 (N_9749,N_8307,N_8512);
xor U9750 (N_9750,N_9321,N_7883);
or U9751 (N_9751,N_7213,N_7601);
nor U9752 (N_9752,N_7092,N_7509);
xor U9753 (N_9753,N_7934,N_7362);
and U9754 (N_9754,N_8396,N_6486);
or U9755 (N_9755,N_7838,N_6977);
nor U9756 (N_9756,N_7617,N_7121);
nand U9757 (N_9757,N_6613,N_7963);
nor U9758 (N_9758,N_8846,N_8514);
xor U9759 (N_9759,N_7353,N_8003);
nand U9760 (N_9760,N_7488,N_6531);
and U9761 (N_9761,N_6651,N_8011);
or U9762 (N_9762,N_7278,N_6982);
xnor U9763 (N_9763,N_7102,N_7611);
or U9764 (N_9764,N_6343,N_9086);
or U9765 (N_9765,N_7463,N_7188);
xnor U9766 (N_9766,N_8682,N_6708);
and U9767 (N_9767,N_8754,N_6567);
xor U9768 (N_9768,N_7427,N_6739);
xnor U9769 (N_9769,N_6569,N_7607);
nand U9770 (N_9770,N_8156,N_8665);
nand U9771 (N_9771,N_8051,N_7000);
or U9772 (N_9772,N_8863,N_6898);
nor U9773 (N_9773,N_7060,N_8591);
nor U9774 (N_9774,N_6907,N_6470);
and U9775 (N_9775,N_6887,N_9294);
xnor U9776 (N_9776,N_7009,N_9317);
and U9777 (N_9777,N_8273,N_8922);
xnor U9778 (N_9778,N_9189,N_9023);
nand U9779 (N_9779,N_6601,N_9322);
and U9780 (N_9780,N_8742,N_8684);
xor U9781 (N_9781,N_8422,N_8167);
or U9782 (N_9782,N_8666,N_8130);
nand U9783 (N_9783,N_8229,N_9096);
or U9784 (N_9784,N_6949,N_8559);
or U9785 (N_9785,N_8867,N_7352);
nor U9786 (N_9786,N_7777,N_6850);
and U9787 (N_9787,N_7641,N_9290);
and U9788 (N_9788,N_7425,N_7886);
nor U9789 (N_9789,N_8418,N_6461);
nand U9790 (N_9790,N_6530,N_9140);
nor U9791 (N_9791,N_8958,N_6947);
or U9792 (N_9792,N_7447,N_9240);
nor U9793 (N_9793,N_7323,N_8121);
nand U9794 (N_9794,N_8789,N_8646);
or U9795 (N_9795,N_8050,N_6518);
nand U9796 (N_9796,N_8417,N_6542);
or U9797 (N_9797,N_7281,N_7108);
nor U9798 (N_9798,N_7466,N_9011);
xnor U9799 (N_9799,N_8450,N_6858);
and U9800 (N_9800,N_6391,N_7649);
nor U9801 (N_9801,N_7222,N_7942);
nand U9802 (N_9802,N_8391,N_7104);
nand U9803 (N_9803,N_6633,N_9132);
nor U9804 (N_9804,N_7065,N_8015);
nand U9805 (N_9805,N_7773,N_8066);
or U9806 (N_9806,N_8605,N_7117);
nand U9807 (N_9807,N_7437,N_6619);
nand U9808 (N_9808,N_7827,N_7956);
nor U9809 (N_9809,N_8136,N_6648);
and U9810 (N_9810,N_6672,N_7527);
or U9811 (N_9811,N_8706,N_8058);
and U9812 (N_9812,N_7317,N_9137);
xnor U9813 (N_9813,N_7176,N_7244);
xnor U9814 (N_9814,N_9093,N_8271);
nand U9815 (N_9815,N_8067,N_9336);
nand U9816 (N_9816,N_9125,N_7179);
nand U9817 (N_9817,N_6406,N_7191);
nor U9818 (N_9818,N_9312,N_7255);
or U9819 (N_9819,N_7854,N_7169);
or U9820 (N_9820,N_6906,N_7050);
nor U9821 (N_9821,N_7047,N_8947);
xnor U9822 (N_9822,N_9257,N_6927);
nand U9823 (N_9823,N_6471,N_6314);
nor U9824 (N_9824,N_6810,N_6702);
or U9825 (N_9825,N_8528,N_7564);
or U9826 (N_9826,N_8833,N_7159);
nand U9827 (N_9827,N_8610,N_8999);
or U9828 (N_9828,N_6719,N_6344);
xnor U9829 (N_9829,N_8776,N_8346);
and U9830 (N_9830,N_7053,N_8240);
or U9831 (N_9831,N_8148,N_7041);
or U9832 (N_9832,N_7859,N_7745);
nor U9833 (N_9833,N_8075,N_6262);
nor U9834 (N_9834,N_9267,N_9262);
or U9835 (N_9835,N_7621,N_8151);
nand U9836 (N_9836,N_8376,N_9362);
or U9837 (N_9837,N_7524,N_7586);
nor U9838 (N_9838,N_8715,N_6999);
xnor U9839 (N_9839,N_8871,N_9318);
xnor U9840 (N_9840,N_7039,N_9064);
and U9841 (N_9841,N_8090,N_8842);
xnor U9842 (N_9842,N_8990,N_7045);
nor U9843 (N_9843,N_6661,N_7666);
and U9844 (N_9844,N_6564,N_7708);
nand U9845 (N_9845,N_8930,N_6712);
and U9846 (N_9846,N_7422,N_7482);
xnor U9847 (N_9847,N_6266,N_6724);
xor U9848 (N_9848,N_8690,N_8289);
or U9849 (N_9849,N_8366,N_8633);
or U9850 (N_9850,N_6707,N_6423);
and U9851 (N_9851,N_7049,N_7915);
xor U9852 (N_9852,N_7904,N_9358);
or U9853 (N_9853,N_9349,N_9369);
or U9854 (N_9854,N_9091,N_7440);
nor U9855 (N_9855,N_7731,N_9316);
nand U9856 (N_9856,N_8533,N_7207);
and U9857 (N_9857,N_7558,N_6934);
nor U9858 (N_9858,N_9243,N_7739);
and U9859 (N_9859,N_7822,N_8513);
and U9860 (N_9860,N_6479,N_6392);
nor U9861 (N_9861,N_7398,N_7200);
xnor U9862 (N_9862,N_7988,N_8811);
nand U9863 (N_9863,N_8214,N_6700);
xnor U9864 (N_9864,N_8686,N_8716);
xnor U9865 (N_9865,N_9014,N_6274);
and U9866 (N_9866,N_8876,N_7825);
or U9867 (N_9867,N_7687,N_7537);
and U9868 (N_9868,N_7386,N_9299);
nand U9869 (N_9869,N_9045,N_6603);
xor U9870 (N_9870,N_9345,N_6467);
nand U9871 (N_9871,N_6482,N_9374);
nand U9872 (N_9872,N_8500,N_6447);
xnor U9873 (N_9873,N_7051,N_8195);
xor U9874 (N_9874,N_8898,N_9114);
nand U9875 (N_9875,N_8721,N_6718);
nand U9876 (N_9876,N_8180,N_7629);
nand U9877 (N_9877,N_6804,N_7403);
and U9878 (N_9878,N_7863,N_7974);
nand U9879 (N_9879,N_7349,N_8446);
nand U9880 (N_9880,N_6265,N_8169);
and U9881 (N_9881,N_7511,N_7303);
or U9882 (N_9882,N_6657,N_8764);
and U9883 (N_9883,N_8614,N_6590);
or U9884 (N_9884,N_9135,N_8565);
or U9885 (N_9885,N_6697,N_6740);
and U9886 (N_9886,N_8012,N_9216);
nor U9887 (N_9887,N_8074,N_8687);
or U9888 (N_9888,N_7125,N_8657);
nand U9889 (N_9889,N_9032,N_8250);
nor U9890 (N_9890,N_8758,N_8172);
or U9891 (N_9891,N_9254,N_8820);
or U9892 (N_9892,N_7373,N_9155);
nand U9893 (N_9893,N_8415,N_8983);
and U9894 (N_9894,N_8507,N_6489);
and U9895 (N_9895,N_7127,N_8211);
nand U9896 (N_9896,N_7584,N_7074);
and U9897 (N_9897,N_9344,N_7156);
nand U9898 (N_9898,N_6914,N_6658);
and U9899 (N_9899,N_7760,N_7319);
or U9900 (N_9900,N_6956,N_8330);
or U9901 (N_9901,N_6312,N_7407);
nor U9902 (N_9902,N_7069,N_9144);
xor U9903 (N_9903,N_7421,N_7633);
nand U9904 (N_9904,N_8221,N_6308);
or U9905 (N_9905,N_6749,N_6717);
xnor U9906 (N_9906,N_7982,N_7532);
nor U9907 (N_9907,N_7913,N_6598);
nand U9908 (N_9908,N_7048,N_8647);
and U9909 (N_9909,N_8047,N_8452);
nand U9910 (N_9910,N_8205,N_7395);
nand U9911 (N_9911,N_8190,N_6685);
or U9912 (N_9912,N_6428,N_8576);
nor U9913 (N_9913,N_7411,N_6550);
nor U9914 (N_9914,N_8803,N_7486);
and U9915 (N_9915,N_8149,N_9300);
and U9916 (N_9916,N_6321,N_8759);
nor U9917 (N_9917,N_8746,N_8738);
nand U9918 (N_9918,N_7563,N_8294);
or U9919 (N_9919,N_8311,N_8860);
or U9920 (N_9920,N_8547,N_6334);
nand U9921 (N_9921,N_6987,N_8262);
xor U9922 (N_9922,N_6506,N_7046);
nor U9923 (N_9923,N_8009,N_6860);
and U9924 (N_9924,N_7487,N_7233);
nor U9925 (N_9925,N_6439,N_7266);
nand U9926 (N_9926,N_7581,N_9323);
or U9927 (N_9927,N_8845,N_6540);
xnor U9928 (N_9928,N_7932,N_8128);
nor U9929 (N_9929,N_8227,N_9103);
nor U9930 (N_9930,N_7003,N_6541);
or U9931 (N_9931,N_6453,N_6616);
xor U9932 (N_9932,N_6449,N_9181);
and U9933 (N_9933,N_7371,N_7388);
nand U9934 (N_9934,N_6617,N_7622);
nor U9935 (N_9935,N_7106,N_8894);
nand U9936 (N_9936,N_8594,N_6754);
xor U9937 (N_9937,N_9040,N_9133);
or U9938 (N_9938,N_7161,N_8660);
nor U9939 (N_9939,N_9033,N_7262);
xnor U9940 (N_9940,N_8481,N_8036);
nor U9941 (N_9941,N_8086,N_7947);
and U9942 (N_9942,N_8632,N_9059);
xor U9943 (N_9943,N_8154,N_8964);
and U9944 (N_9944,N_6899,N_6683);
nand U9945 (N_9945,N_9124,N_7429);
or U9946 (N_9946,N_9292,N_8839);
nor U9947 (N_9947,N_7810,N_6939);
and U9948 (N_9948,N_6831,N_7162);
xor U9949 (N_9949,N_8176,N_8786);
nand U9950 (N_9950,N_6250,N_8055);
xor U9951 (N_9951,N_7618,N_7986);
xor U9952 (N_9952,N_7898,N_6289);
xnor U9953 (N_9953,N_9276,N_8918);
or U9954 (N_9954,N_7261,N_6502);
nor U9955 (N_9955,N_7252,N_8013);
nor U9956 (N_9956,N_7090,N_7812);
and U9957 (N_9957,N_7655,N_8332);
and U9958 (N_9958,N_8495,N_6856);
and U9959 (N_9959,N_8489,N_6875);
nor U9960 (N_9960,N_6877,N_9315);
and U9961 (N_9961,N_8834,N_8841);
nand U9962 (N_9962,N_8319,N_8815);
nor U9963 (N_9963,N_6891,N_8295);
xor U9964 (N_9964,N_6820,N_9139);
xnor U9965 (N_9965,N_7661,N_8472);
xor U9966 (N_9966,N_8980,N_8926);
xor U9967 (N_9967,N_8085,N_9270);
nor U9968 (N_9968,N_6252,N_7406);
nand U9969 (N_9969,N_8939,N_7140);
xnor U9970 (N_9970,N_8032,N_6403);
xnor U9971 (N_9971,N_7921,N_6586);
nor U9972 (N_9972,N_8763,N_6474);
and U9973 (N_9973,N_9002,N_6930);
and U9974 (N_9974,N_8261,N_6978);
xor U9975 (N_9975,N_9069,N_6952);
nand U9976 (N_9976,N_7608,N_7990);
nand U9977 (N_9977,N_9338,N_8157);
and U9978 (N_9978,N_8232,N_8053);
or U9979 (N_9979,N_7454,N_9063);
xnor U9980 (N_9980,N_7996,N_8562);
nor U9981 (N_9981,N_6503,N_6304);
and U9982 (N_9982,N_6505,N_8411);
xor U9983 (N_9983,N_9166,N_7375);
nor U9984 (N_9984,N_7184,N_7459);
or U9985 (N_9985,N_8679,N_9365);
or U9986 (N_9986,N_7669,N_7241);
xor U9987 (N_9987,N_8836,N_7105);
and U9988 (N_9988,N_7192,N_6434);
nor U9989 (N_9989,N_8911,N_7013);
nor U9990 (N_9990,N_6433,N_6527);
or U9991 (N_9991,N_8539,N_7336);
xnor U9992 (N_9992,N_6744,N_9233);
or U9993 (N_9993,N_6283,N_6287);
xor U9994 (N_9994,N_7848,N_6501);
or U9995 (N_9995,N_8451,N_8228);
or U9996 (N_9996,N_7703,N_7366);
xor U9997 (N_9997,N_8380,N_8521);
nand U9998 (N_9998,N_8689,N_6955);
and U9999 (N_9999,N_7926,N_7519);
nand U10000 (N_10000,N_6573,N_8831);
and U10001 (N_10001,N_7350,N_7779);
nand U10002 (N_10002,N_8044,N_7451);
nand U10003 (N_10003,N_7330,N_8586);
and U10004 (N_10004,N_8397,N_9289);
nand U10005 (N_10005,N_8219,N_6933);
or U10006 (N_10006,N_6911,N_9018);
nand U10007 (N_10007,N_7624,N_6801);
nand U10008 (N_10008,N_7499,N_6385);
nor U10009 (N_10009,N_6979,N_7727);
nor U10010 (N_10010,N_7991,N_8409);
and U10011 (N_10011,N_6771,N_8756);
nor U10012 (N_10012,N_6563,N_6317);
or U10013 (N_10013,N_9226,N_7183);
nand U10014 (N_10014,N_8501,N_8076);
and U10015 (N_10015,N_8096,N_7517);
xor U10016 (N_10016,N_6260,N_8830);
or U10017 (N_10017,N_8942,N_8268);
or U10018 (N_10018,N_7889,N_9303);
or U10019 (N_10019,N_6583,N_8441);
xnor U10020 (N_10020,N_8054,N_7150);
and U10021 (N_10021,N_8814,N_7605);
nor U10022 (N_10022,N_7139,N_7204);
nand U10023 (N_10023,N_8187,N_6836);
or U10024 (N_10024,N_8474,N_9204);
nor U10025 (N_10025,N_8801,N_8611);
or U10026 (N_10026,N_8720,N_7325);
xnor U10027 (N_10027,N_7744,N_9212);
nor U10028 (N_10028,N_8491,N_7250);
nor U10029 (N_10029,N_8989,N_7507);
nor U10030 (N_10030,N_9359,N_8761);
nor U10031 (N_10031,N_7652,N_8108);
nor U10032 (N_10032,N_6812,N_8574);
or U10033 (N_10033,N_9246,N_7850);
or U10034 (N_10034,N_7689,N_7369);
or U10035 (N_10035,N_7738,N_7844);
nand U10036 (N_10036,N_6299,N_7700);
nand U10037 (N_10037,N_7025,N_9180);
nand U10038 (N_10038,N_8191,N_8388);
and U10039 (N_10039,N_6324,N_8877);
and U10040 (N_10040,N_7723,N_7533);
and U10041 (N_10041,N_7637,N_8927);
nand U10042 (N_10042,N_7076,N_8281);
or U10043 (N_10043,N_6463,N_8879);
xor U10044 (N_10044,N_9296,N_8608);
or U10045 (N_10045,N_7056,N_9015);
or U10046 (N_10046,N_8954,N_9170);
nand U10047 (N_10047,N_8564,N_6918);
nor U10048 (N_10048,N_6524,N_7124);
nor U10049 (N_10049,N_8112,N_7797);
nand U10050 (N_10050,N_9325,N_7998);
nor U10051 (N_10051,N_6863,N_7109);
and U10052 (N_10052,N_7888,N_8971);
or U10053 (N_10053,N_7809,N_8694);
nand U10054 (N_10054,N_7650,N_9035);
xor U10055 (N_10055,N_8515,N_7803);
or U10056 (N_10056,N_6841,N_6703);
xnor U10057 (N_10057,N_9055,N_8347);
nor U10058 (N_10058,N_8554,N_8504);
nand U10059 (N_10059,N_7264,N_6673);
nand U10060 (N_10060,N_8735,N_6574);
nor U10061 (N_10061,N_8302,N_8925);
nor U10062 (N_10062,N_9271,N_8639);
nand U10063 (N_10063,N_9238,N_7994);
xnor U10064 (N_10064,N_6340,N_7307);
xor U10065 (N_10065,N_8468,N_7575);
nand U10066 (N_10066,N_8287,N_6834);
nand U10067 (N_10067,N_6681,N_7163);
nand U10068 (N_10068,N_6293,N_8425);
nand U10069 (N_10069,N_8082,N_6484);
and U10070 (N_10070,N_8236,N_7591);
nand U10071 (N_10071,N_9253,N_8731);
or U10072 (N_10072,N_6495,N_7272);
and U10073 (N_10073,N_9104,N_8672);
nor U10074 (N_10074,N_6735,N_7701);
nand U10075 (N_10075,N_6362,N_9118);
xor U10076 (N_10076,N_6429,N_9348);
nand U10077 (N_10077,N_8625,N_6786);
or U10078 (N_10078,N_6487,N_8344);
nand U10079 (N_10079,N_6545,N_7098);
xnor U10080 (N_10080,N_6692,N_6646);
nand U10081 (N_10081,N_8931,N_9129);
nor U10082 (N_10082,N_7029,N_6383);
xor U10083 (N_10083,N_7496,N_7946);
or U10084 (N_10084,N_7761,N_7950);
or U10085 (N_10085,N_8004,N_9058);
nor U10086 (N_10086,N_8116,N_7843);
and U10087 (N_10087,N_6675,N_6594);
and U10088 (N_10088,N_8178,N_8127);
nor U10089 (N_10089,N_7692,N_6943);
xnor U10090 (N_10090,N_7767,N_9280);
nand U10091 (N_10091,N_6917,N_9211);
xnor U10092 (N_10092,N_7928,N_9057);
xor U10093 (N_10093,N_7418,N_7038);
and U10094 (N_10094,N_8313,N_8327);
nor U10095 (N_10095,N_6851,N_7223);
xor U10096 (N_10096,N_7710,N_6349);
nand U10097 (N_10097,N_9121,N_7112);
xnor U10098 (N_10098,N_6975,N_6926);
nor U10099 (N_10099,N_8341,N_6534);
and U10100 (N_10100,N_8340,N_7095);
nand U10101 (N_10101,N_6626,N_6468);
xor U10102 (N_10102,N_8316,N_7172);
nor U10103 (N_10103,N_7931,N_6803);
and U10104 (N_10104,N_8525,N_6756);
nor U10105 (N_10105,N_7668,N_6342);
nand U10106 (N_10106,N_7654,N_9044);
nor U10107 (N_10107,N_8486,N_8234);
nand U10108 (N_10108,N_6981,N_7279);
or U10109 (N_10109,N_6711,N_7842);
and U10110 (N_10110,N_8673,N_6753);
xnor U10111 (N_10111,N_6837,N_7590);
and U10112 (N_10112,N_6398,N_7805);
and U10113 (N_10113,N_6806,N_6570);
or U10114 (N_10114,N_8387,N_7680);
and U10115 (N_10115,N_7879,N_7058);
and U10116 (N_10116,N_7294,N_7329);
xnor U10117 (N_10117,N_6290,N_7730);
and U10118 (N_10118,N_6716,N_7240);
nand U10119 (N_10119,N_9025,N_9309);
nor U10120 (N_10120,N_6568,N_6787);
and U10121 (N_10121,N_6445,N_7337);
or U10122 (N_10122,N_7320,N_6883);
and U10123 (N_10123,N_7677,N_8264);
or U10124 (N_10124,N_7147,N_7164);
nor U10125 (N_10125,N_9053,N_7079);
nand U10126 (N_10126,N_7828,N_9198);
nand U10127 (N_10127,N_7446,N_8883);
nor U10128 (N_10128,N_7857,N_8712);
nor U10129 (N_10129,N_8997,N_8623);
and U10130 (N_10130,N_7714,N_8966);
nor U10131 (N_10131,N_8643,N_8826);
nand U10132 (N_10132,N_8137,N_9241);
and U10133 (N_10133,N_9343,N_7908);
nor U10134 (N_10134,N_8567,N_6827);
nand U10135 (N_10135,N_8965,N_7945);
nor U10136 (N_10136,N_6874,N_8359);
nand U10137 (N_10137,N_7837,N_7566);
xnor U10138 (N_10138,N_6872,N_7450);
nor U10139 (N_10139,N_8428,N_8998);
or U10140 (N_10140,N_8023,N_7456);
nand U10141 (N_10141,N_8534,N_7506);
or U10142 (N_10142,N_8360,N_6480);
nor U10143 (N_10143,N_8641,N_7547);
or U10144 (N_10144,N_7722,N_6878);
xor U10145 (N_10145,N_6818,N_8571);
or U10146 (N_10146,N_9017,N_8832);
xnor U10147 (N_10147,N_8255,N_6490);
nand U10148 (N_10148,N_8609,N_9158);
xor U10149 (N_10149,N_8105,N_8992);
and U10150 (N_10150,N_9278,N_9199);
and U10151 (N_10151,N_6859,N_8006);
nand U10152 (N_10152,N_8557,N_7734);
and U10153 (N_10153,N_7332,N_8976);
or U10154 (N_10154,N_7285,N_7662);
xnor U10155 (N_10155,N_7180,N_8532);
xor U10156 (N_10156,N_8147,N_8511);
nand U10157 (N_10157,N_6902,N_8290);
or U10158 (N_10158,N_8005,N_6622);
and U10159 (N_10159,N_7589,N_9165);
and U10160 (N_10160,N_7197,N_9001);
nor U10161 (N_10161,N_8584,N_8125);
xor U10162 (N_10162,N_7128,N_9113);
nand U10163 (N_10163,N_8723,N_8767);
nor U10164 (N_10164,N_7005,N_6404);
nand U10165 (N_10165,N_9186,N_6354);
nand U10166 (N_10166,N_9016,N_8865);
nand U10167 (N_10167,N_6498,N_6640);
nand U10168 (N_10168,N_8046,N_8335);
or U10169 (N_10169,N_7249,N_7830);
xnor U10170 (N_10170,N_7028,N_7672);
and U10171 (N_10171,N_6327,N_8799);
or U10172 (N_10172,N_7569,N_8698);
nor U10173 (N_10173,N_8578,N_7331);
xnor U10174 (N_10174,N_9024,N_6743);
or U10175 (N_10175,N_8544,N_6665);
and U10176 (N_10176,N_7737,N_8091);
nand U10177 (N_10177,N_6691,N_7659);
xnor U10178 (N_10178,N_7202,N_8343);
and U10179 (N_10179,N_7979,N_6372);
nand U10180 (N_10180,N_8943,N_6746);
or U10181 (N_10181,N_6414,N_9200);
nor U10182 (N_10182,N_6592,N_7811);
xnor U10183 (N_10183,N_6805,N_9239);
nor U10184 (N_10184,N_8748,N_8523);
xor U10185 (N_10185,N_7115,N_7006);
and U10186 (N_10186,N_6350,N_7322);
nand U10187 (N_10187,N_7960,N_8384);
nand U10188 (N_10188,N_7953,N_9005);
or U10189 (N_10189,N_6254,N_8717);
nand U10190 (N_10190,N_6699,N_8308);
and U10191 (N_10191,N_8144,N_8161);
nor U10192 (N_10192,N_7801,N_8269);
and U10193 (N_10193,N_7238,N_9231);
nor U10194 (N_10194,N_8035,N_8699);
and U10195 (N_10195,N_7301,N_9191);
and U10196 (N_10196,N_8695,N_8597);
and U10197 (N_10197,N_7561,N_8919);
xnor U10198 (N_10198,N_7513,N_8088);
or U10199 (N_10199,N_6300,N_6808);
nor U10200 (N_10200,N_6353,N_7054);
nor U10201 (N_10201,N_7885,N_7531);
and U10202 (N_10202,N_7243,N_7693);
and U10203 (N_10203,N_8089,N_8323);
nor U10204 (N_10204,N_6662,N_7973);
xnor U10205 (N_10205,N_8379,N_9146);
nand U10206 (N_10206,N_6966,N_8378);
and U10207 (N_10207,N_9062,N_7103);
and U10208 (N_10208,N_7379,N_7686);
nand U10209 (N_10209,N_8887,N_8664);
nor U10210 (N_10210,N_8369,N_6496);
nand U10211 (N_10211,N_8062,N_8615);
xnor U10212 (N_10212,N_6865,N_6497);
xor U10213 (N_10213,N_6517,N_6867);
nor U10214 (N_10214,N_6311,N_8152);
or U10215 (N_10215,N_7471,N_8095);
xnor U10216 (N_10216,N_7775,N_6706);
nand U10217 (N_10217,N_8375,N_6813);
nand U10218 (N_10218,N_8001,N_8579);
and U10219 (N_10219,N_9072,N_7799);
and U10220 (N_10220,N_8683,N_6303);
or U10221 (N_10221,N_7236,N_9355);
xnor U10222 (N_10222,N_7171,N_8493);
and U10223 (N_10223,N_6751,N_9353);
xnor U10224 (N_10224,N_9229,N_8142);
and U10225 (N_10225,N_7120,N_9340);
or U10226 (N_10226,N_6815,N_6854);
nor U10227 (N_10227,N_6579,N_7248);
or U10228 (N_10228,N_6417,N_6921);
nand U10229 (N_10229,N_7671,N_9167);
nor U10230 (N_10230,N_8652,N_6360);
and U10231 (N_10231,N_8696,N_7394);
xor U10232 (N_10232,N_6896,N_9013);
or U10233 (N_10233,N_8601,N_8420);
xor U10234 (N_10234,N_8404,N_9075);
nor U10235 (N_10235,N_6728,N_8740);
nand U10236 (N_10236,N_8692,N_7309);
nor U10237 (N_10237,N_8862,N_8222);
nor U10238 (N_10238,N_6799,N_7091);
and U10239 (N_10239,N_8550,N_6761);
xnor U10240 (N_10240,N_6537,N_8235);
and U10241 (N_10241,N_7529,N_7153);
xnor U10242 (N_10242,N_7063,N_6929);
and U10243 (N_10243,N_7295,N_7656);
and U10244 (N_10244,N_8153,N_8104);
nand U10245 (N_10245,N_6411,N_8060);
or U10246 (N_10246,N_9168,N_7841);
and U10247 (N_10247,N_8064,N_8558);
nand U10248 (N_10248,N_6376,N_6415);
xnor U10249 (N_10249,N_6932,N_6288);
and U10250 (N_10250,N_6280,N_6292);
or U10251 (N_10251,N_7435,N_6830);
or U10252 (N_10252,N_7631,N_9250);
xor U10253 (N_10253,N_7865,N_9346);
nor U10254 (N_10254,N_9265,N_8329);
or U10255 (N_10255,N_6438,N_6822);
xor U10256 (N_10256,N_8642,N_6628);
nand U10257 (N_10257,N_7040,N_9109);
xor U10258 (N_10258,N_8383,N_7286);
nor U10259 (N_10259,N_7101,N_8542);
nand U10260 (N_10260,N_7078,N_7455);
nand U10261 (N_10261,N_9293,N_9078);
or U10262 (N_10262,N_7186,N_8886);
nand U10263 (N_10263,N_9149,N_7774);
and U10264 (N_10264,N_8259,N_6781);
nor U10265 (N_10265,N_8291,N_8079);
or U10266 (N_10266,N_8120,N_6843);
or U10267 (N_10267,N_9248,N_8588);
xnor U10268 (N_10268,N_7679,N_6272);
nor U10269 (N_10269,N_6405,N_7365);
nor U10270 (N_10270,N_6315,N_8080);
and U10271 (N_10271,N_6499,N_6512);
xor U10272 (N_10272,N_7769,N_8938);
xnor U10273 (N_10273,N_6418,N_8580);
and U10274 (N_10274,N_6835,N_6962);
nor U10275 (N_10275,N_7632,N_9029);
nor U10276 (N_10276,N_8870,N_8593);
or U10277 (N_10277,N_7514,N_8061);
xnor U10278 (N_10278,N_8355,N_6732);
or U10279 (N_10279,N_7602,N_7663);
and U10280 (N_10280,N_8466,N_8693);
xor U10281 (N_10281,N_7208,N_9356);
xnor U10282 (N_10282,N_7847,N_9156);
and U10283 (N_10283,N_8276,N_8995);
nand U10284 (N_10284,N_9222,N_7576);
xnor U10285 (N_10285,N_6559,N_8783);
xnor U10286 (N_10286,N_7592,N_8208);
xor U10287 (N_10287,N_7735,N_9090);
xor U10288 (N_10288,N_8889,N_7151);
or U10289 (N_10289,N_8945,N_6768);
nand U10290 (N_10290,N_7583,N_6638);
xor U10291 (N_10291,N_9203,N_7874);
nor U10292 (N_10292,N_7907,N_8810);
nand U10293 (N_10293,N_6844,N_7035);
nand U10294 (N_10294,N_6653,N_7705);
nor U10295 (N_10295,N_8802,N_6725);
nor U10296 (N_10296,N_6632,N_7289);
nand U10297 (N_10297,N_8073,N_7400);
and U10298 (N_10298,N_7995,N_7327);
xor U10299 (N_10299,N_8624,N_7609);
nand U10300 (N_10300,N_7409,N_6864);
nand U10301 (N_10301,N_6670,N_6773);
or U10302 (N_10302,N_6329,N_8818);
and U10303 (N_10303,N_7497,N_8852);
or U10304 (N_10304,N_8093,N_8520);
or U10305 (N_10305,N_6620,N_8640);
and U10306 (N_10306,N_7989,N_8847);
xor U10307 (N_10307,N_7360,N_7833);
xor U10308 (N_10308,N_9372,N_7699);
and U10309 (N_10309,N_7443,N_9335);
nor U10310 (N_10310,N_8462,N_9095);
nand U10311 (N_10311,N_7503,N_7867);
nand U10312 (N_10312,N_7720,N_7075);
nor U10313 (N_10313,N_8174,N_8940);
and U10314 (N_10314,N_8057,N_7978);
nor U10315 (N_10315,N_7413,N_8775);
or U10316 (N_10316,N_7638,N_6316);
and U10317 (N_10317,N_7458,N_8935);
or U10318 (N_10318,N_8575,N_7305);
nand U10319 (N_10319,N_8284,N_8286);
nand U10320 (N_10320,N_8293,N_8403);
and U10321 (N_10321,N_6762,N_6270);
nor U10322 (N_10322,N_8910,N_8363);
nand U10323 (N_10323,N_7410,N_7464);
xnor U10324 (N_10324,N_7548,N_7695);
or U10325 (N_10325,N_6992,N_8561);
nor U10326 (N_10326,N_7348,N_9182);
xor U10327 (N_10327,N_7182,N_7545);
and U10328 (N_10328,N_7152,N_7940);
and U10329 (N_10329,N_6432,N_8146);
nand U10330 (N_10330,N_8853,N_6279);
or U10331 (N_10331,N_6840,N_7168);
or U10332 (N_10332,N_7967,N_8709);
xnor U10333 (N_10333,N_8336,N_7224);
or U10334 (N_10334,N_8985,N_8201);
xor U10335 (N_10335,N_7196,N_7758);
or U10336 (N_10336,N_9220,N_6729);
and U10337 (N_10337,N_8225,N_7116);
or U10338 (N_10338,N_7479,N_6547);
and U10339 (N_10339,N_8793,N_6612);
xor U10340 (N_10340,N_7834,N_7228);
nor U10341 (N_10341,N_7894,N_8467);
xnor U10342 (N_10342,N_8160,N_8257);
or U10343 (N_10343,N_9116,N_8702);
or U10344 (N_10344,N_8192,N_7742);
nand U10345 (N_10345,N_7144,N_6807);
nand U10346 (N_10346,N_8470,N_7111);
and U10347 (N_10347,N_8150,N_7980);
nor U10348 (N_10348,N_8258,N_6307);
and U10349 (N_10349,N_8849,N_6663);
xor U10350 (N_10350,N_7992,N_8900);
xnor U10351 (N_10351,N_7382,N_7083);
and U10352 (N_10352,N_7086,N_7258);
nor U10353 (N_10353,N_8496,N_9012);
and U10354 (N_10354,N_8312,N_6551);
xor U10355 (N_10355,N_7126,N_7143);
nand U10356 (N_10356,N_6332,N_7300);
nor U10357 (N_10357,N_8173,N_7291);
or U10358 (N_10358,N_9079,N_8653);
and U10359 (N_10359,N_6893,N_6339);
and U10360 (N_10360,N_8419,N_8049);
and U10361 (N_10361,N_7770,N_6794);
nand U10362 (N_10362,N_8320,N_6255);
and U10363 (N_10363,N_6386,N_7674);
xnor U10364 (N_10364,N_8680,N_6306);
nand U10365 (N_10365,N_7251,N_7316);
and U10366 (N_10366,N_8245,N_8618);
nor U10367 (N_10367,N_6257,N_8238);
nor U10368 (N_10368,N_8087,N_7782);
nand U10369 (N_10369,N_7845,N_6256);
xnor U10370 (N_10370,N_8636,N_6792);
nor U10371 (N_10371,N_8433,N_7137);
xor U10372 (N_10372,N_7472,N_7808);
nor U10373 (N_10373,N_7080,N_7993);
nor U10374 (N_10374,N_7897,N_6516);
xnor U10375 (N_10375,N_8453,N_9019);
xnor U10376 (N_10376,N_9106,N_8987);
nor U10377 (N_10377,N_9366,N_7133);
or U10378 (N_10378,N_6797,N_7905);
xor U10379 (N_10379,N_7916,N_9060);
xor U10380 (N_10380,N_6345,N_9218);
and U10381 (N_10381,N_7751,N_8804);
nand U10382 (N_10382,N_7873,N_6509);
xor U10383 (N_10383,N_8408,N_7750);
and U10384 (N_10384,N_6961,N_7552);
nor U10385 (N_10385,N_6462,N_8476);
or U10386 (N_10386,N_7203,N_8241);
nor U10387 (N_10387,N_7892,N_8932);
and U10388 (N_10388,N_6847,N_6597);
and U10389 (N_10389,N_8458,N_6995);
and U10390 (N_10390,N_9324,N_6448);
nand U10391 (N_10391,N_9157,N_6763);
and U10392 (N_10392,N_8552,N_7201);
and U10393 (N_10393,N_8400,N_8944);
xnor U10394 (N_10394,N_7198,N_6553);
or U10395 (N_10395,N_6817,N_7475);
nor U10396 (N_10396,N_8499,N_7521);
nor U10397 (N_10397,N_8406,N_6845);
nand U10398 (N_10398,N_6500,N_6894);
xor U10399 (N_10399,N_9036,N_6611);
xnor U10400 (N_10400,N_7311,N_7170);
nor U10401 (N_10401,N_6420,N_9021);
nand U10402 (N_10402,N_7971,N_8018);
nor U10403 (N_10403,N_7719,N_7096);
and U10404 (N_10404,N_7784,N_9119);
nand U10405 (N_10405,N_6824,N_7381);
xnor U10406 (N_10406,N_7818,N_6637);
nand U10407 (N_10407,N_8516,N_7024);
nor U10408 (N_10408,N_8427,N_7855);
nor U10409 (N_10409,N_7959,N_8212);
xnor U10410 (N_10410,N_6630,N_8732);
nor U10411 (N_10411,N_8197,N_9213);
nor U10412 (N_10412,N_8126,N_8498);
and U10413 (N_10413,N_8851,N_8675);
xor U10414 (N_10414,N_8730,N_6625);
and U10415 (N_10415,N_7328,N_8278);
nand U10416 (N_10416,N_9277,N_6440);
xnor U10417 (N_10417,N_8920,N_8155);
xnor U10418 (N_10418,N_7538,N_7110);
nand U10419 (N_10419,N_6828,N_8233);
nand U10420 (N_10420,N_6936,N_7887);
nor U10421 (N_10421,N_6644,N_7951);
xnor U10422 (N_10422,N_6370,N_6904);
nor U10423 (N_10423,N_9150,N_8310);
xor U10424 (N_10424,N_8171,N_6602);
or U10425 (N_10425,N_6985,N_6388);
or U10426 (N_10426,N_7431,N_6660);
nand U10427 (N_10427,N_8209,N_7573);
nand U10428 (N_10428,N_6666,N_7539);
xnor U10429 (N_10429,N_6669,N_9264);
nor U10430 (N_10430,N_7968,N_7502);
xnor U10431 (N_10431,N_8322,N_9368);
or U10432 (N_10432,N_8482,N_8924);
and U10433 (N_10433,N_7306,N_8885);
or U10434 (N_10434,N_7315,N_8956);
and U10435 (N_10435,N_7358,N_8795);
xnor U10436 (N_10436,N_7819,N_7492);
or U10437 (N_10437,N_7626,N_9352);
xnor U10438 (N_10438,N_9126,N_9067);
nand U10439 (N_10439,N_6671,N_8455);
or U10440 (N_10440,N_8386,N_7190);
nand U10441 (N_10441,N_6546,N_9077);
xor U10442 (N_10442,N_8410,N_9054);
or U10443 (N_10443,N_8158,N_7372);
and U10444 (N_10444,N_8540,N_9363);
nor U10445 (N_10445,N_8292,N_8436);
nor U10446 (N_10446,N_6444,N_8368);
nand U10447 (N_10447,N_8902,N_8509);
or U10448 (N_10448,N_7789,N_8318);
or U10449 (N_10449,N_7099,N_8182);
or U10450 (N_10450,N_6833,N_9041);
nand U10451 (N_10451,N_9110,N_7929);
xnor U10452 (N_10452,N_6582,N_9288);
or U10453 (N_10453,N_8807,N_6380);
or U10454 (N_10454,N_9311,N_8298);
or U10455 (N_10455,N_7019,N_8432);
or U10456 (N_10456,N_9128,N_6892);
xor U10457 (N_10457,N_9159,N_8543);
or U10458 (N_10458,N_8072,N_6923);
nand U10459 (N_10459,N_8399,N_6688);
nor U10460 (N_10460,N_6493,N_7616);
or U10461 (N_10461,N_8124,N_8714);
or U10462 (N_10462,N_7643,N_8405);
and U10463 (N_10463,N_6458,N_7829);
xor U10464 (N_10464,N_8572,N_7935);
nor U10465 (N_10465,N_7670,N_6912);
nand U10466 (N_10466,N_6412,N_7335);
and U10467 (N_10467,N_7957,N_7067);
nor U10468 (N_10468,N_8488,N_7597);
or U10469 (N_10469,N_7870,N_8395);
nand U10470 (N_10470,N_8747,N_7726);
or U10471 (N_10471,N_7157,N_8266);
xnor U10472 (N_10472,N_7685,N_7189);
nand U10473 (N_10473,N_8034,N_7339);
and U10474 (N_10474,N_7087,N_7211);
or U10475 (N_10475,N_6533,N_8306);
nor U10476 (N_10476,N_7522,N_8361);
xor U10477 (N_10477,N_8030,N_8729);
or U10478 (N_10478,N_6488,N_9192);
and U10479 (N_10479,N_8546,N_9174);
or U10480 (N_10480,N_7018,N_8872);
and U10481 (N_10481,N_7640,N_8352);
or U10482 (N_10482,N_8519,N_8903);
xor U10483 (N_10483,N_6888,N_6320);
and U10484 (N_10484,N_8207,N_8788);
or U10485 (N_10485,N_7781,N_8186);
or U10486 (N_10486,N_6968,N_6986);
xor U10487 (N_10487,N_8017,N_8239);
nor U10488 (N_10488,N_6543,N_6532);
nand U10489 (N_10489,N_6584,N_9042);
and U10490 (N_10490,N_7206,N_6585);
or U10491 (N_10491,N_7094,N_7826);
and U10492 (N_10492,N_8969,N_8356);
or U10493 (N_10493,N_7361,N_7246);
nand U10494 (N_10494,N_6396,N_8891);
nor U10495 (N_10495,N_8617,N_9373);
nor U10496 (N_10496,N_7851,N_8503);
or U10497 (N_10497,N_6734,N_7878);
xor U10498 (N_10498,N_7273,N_7364);
nand U10499 (N_10499,N_8296,N_7221);
nand U10500 (N_10500,N_6783,N_7981);
and U10501 (N_10501,N_8560,N_7195);
xnor U10502 (N_10502,N_6593,N_7944);
nor U10503 (N_10503,N_7302,N_9236);
or U10504 (N_10504,N_9357,N_7535);
nor U10505 (N_10505,N_6330,N_6323);
xor U10506 (N_10506,N_7918,N_8440);
nor U10507 (N_10507,N_9076,N_8796);
nor U10508 (N_10508,N_7493,N_6778);
or U10509 (N_10509,N_8244,N_7253);
and U10510 (N_10510,N_6485,N_7642);
or U10511 (N_10511,N_6368,N_8272);
nor U10512 (N_10512,N_8768,N_8435);
or U10513 (N_10513,N_8123,N_7690);
nor U10514 (N_10514,N_7580,N_7587);
and U10515 (N_10515,N_8753,N_7523);
xnor U10516 (N_10516,N_8374,N_8570);
nand U10517 (N_10517,N_8162,N_7786);
or U10518 (N_10518,N_6958,N_7299);
or U10519 (N_10519,N_9259,N_6925);
or U10520 (N_10520,N_7321,N_6394);
nor U10521 (N_10521,N_7510,N_8483);
and U10522 (N_10522,N_9245,N_8071);
nand U10523 (N_10523,N_7037,N_8825);
or U10524 (N_10524,N_6928,N_7939);
xnor U10525 (N_10525,N_9339,N_7800);
or U10526 (N_10526,N_7684,N_8010);
or U10527 (N_10527,N_9176,N_7604);
or U10528 (N_10528,N_7965,N_6375);
and U10529 (N_10529,N_7697,N_9268);
or U10530 (N_10530,N_8141,N_6832);
nor U10531 (N_10531,N_9065,N_8737);
and U10532 (N_10532,N_8798,N_6791);
nor U10533 (N_10533,N_7412,N_8619);
nor U10534 (N_10534,N_7491,N_6609);
nor U10535 (N_10535,N_6419,N_7557);
or U10536 (N_10536,N_9050,N_7280);
and U10537 (N_10537,N_7821,N_9027);
xor U10538 (N_10538,N_7495,N_6667);
or U10539 (N_10539,N_9274,N_6969);
and U10540 (N_10540,N_7762,N_9000);
and U10541 (N_10541,N_7347,N_8179);
and U10542 (N_10542,N_6421,N_9026);
or U10543 (N_10543,N_8331,N_8638);
or U10544 (N_10544,N_7274,N_8991);
and U10545 (N_10545,N_6738,N_6970);
nand U10546 (N_10546,N_7334,N_7644);
nand U10547 (N_10547,N_9291,N_6377);
and U10548 (N_10548,N_7543,N_9263);
nand U10549 (N_10549,N_7042,N_7976);
nand U10550 (N_10550,N_6363,N_8188);
xor U10551 (N_10551,N_6588,N_8460);
nor U10552 (N_10552,N_8739,N_8285);
nand U10553 (N_10553,N_6401,N_7966);
nand U10554 (N_10554,N_7467,N_8744);
xor U10555 (N_10555,N_9273,N_8620);
and U10556 (N_10556,N_9003,N_9197);
xnor U10557 (N_10557,N_8648,N_9046);
nand U10558 (N_10558,N_6897,N_8736);
and U10559 (N_10559,N_6722,N_7177);
and U10560 (N_10560,N_9171,N_9098);
and U10561 (N_10561,N_6513,N_6649);
nor U10562 (N_10562,N_6963,N_8858);
nor U10563 (N_10563,N_6991,N_6726);
nor U10564 (N_10564,N_7247,N_8828);
and U10565 (N_10565,N_7606,N_7100);
nor U10566 (N_10566,N_9214,N_7925);
xnor U10567 (N_10567,N_7836,N_7417);
nand U10568 (N_10568,N_7237,N_6263);
or U10569 (N_10569,N_8338,N_9210);
xnor U10570 (N_10570,N_9163,N_9088);
and U10571 (N_10571,N_7293,N_8583);
nor U10572 (N_10572,N_6686,N_7376);
nand U10573 (N_10573,N_6846,N_7428);
nand U10574 (N_10574,N_6682,N_6357);
or U10575 (N_10575,N_6301,N_9122);
xnor U10576 (N_10576,N_8045,N_7711);
or U10577 (N_10577,N_9208,N_6634);
and U10578 (N_10578,N_8502,N_8901);
or U10579 (N_10579,N_6337,N_7268);
and U10580 (N_10580,N_7709,N_8676);
or U10581 (N_10581,N_6437,N_6456);
nand U10582 (N_10582,N_7077,N_7342);
nand U10583 (N_10583,N_8083,N_7392);
or U10584 (N_10584,N_6652,N_6515);
xor U10585 (N_10585,N_6767,N_8972);
nor U10586 (N_10586,N_8324,N_8671);
nand U10587 (N_10587,N_8370,N_7756);
nand U10588 (N_10588,N_8880,N_8106);
xnor U10589 (N_10589,N_8213,N_7955);
nor U10590 (N_10590,N_7033,N_8024);
or U10591 (N_10591,N_7920,N_6600);
or U10592 (N_10592,N_7554,N_9037);
or U10593 (N_10593,N_8549,N_8631);
nor U10594 (N_10594,N_8339,N_8713);
or U10595 (N_10595,N_8416,N_9225);
or U10596 (N_10596,N_8202,N_8469);
nor U10597 (N_10597,N_9020,N_7902);
nor U10598 (N_10598,N_8065,N_8951);
and U10599 (N_10599,N_8390,N_8377);
or U10600 (N_10600,N_6793,N_8131);
xnor U10601 (N_10601,N_6776,N_9286);
nand U10602 (N_10602,N_7972,N_7114);
and U10603 (N_10603,N_8774,N_8967);
xor U10604 (N_10604,N_7383,N_7949);
nand U10605 (N_10605,N_6581,N_6755);
xnor U10606 (N_10606,N_6876,N_6668);
nand U10607 (N_10607,N_6454,N_8438);
or U10608 (N_10608,N_8301,N_6825);
or U10609 (N_10609,N_6779,N_6273);
and U10610 (N_10610,N_7871,N_7798);
xor U10611 (N_10611,N_7004,N_6561);
nand U10612 (N_10612,N_8139,N_7234);
and U10613 (N_10613,N_7862,N_7227);
and U10614 (N_10614,N_6371,N_6278);
or U10615 (N_10615,N_6659,N_9329);
and U10616 (N_10616,N_8703,N_8563);
or U10617 (N_10617,N_8143,N_8487);
and U10618 (N_10618,N_6871,N_6465);
nand U10619 (N_10619,N_8770,N_6727);
and U10620 (N_10620,N_7565,N_6384);
and U10621 (N_10621,N_8163,N_6536);
xnor U10622 (N_10622,N_6606,N_7194);
nand U10623 (N_10623,N_7181,N_9039);
nor U10624 (N_10624,N_7776,N_7484);
nand U10625 (N_10625,N_6457,N_7304);
and U10626 (N_10626,N_7245,N_7508);
and U10627 (N_10627,N_9302,N_7882);
xor U10628 (N_10628,N_8888,N_6960);
xnor U10629 (N_10629,N_8038,N_7423);
xor U10630 (N_10630,N_6604,N_7635);
nand U10631 (N_10631,N_8505,N_8442);
nor U10632 (N_10632,N_7380,N_7219);
xnor U10633 (N_10633,N_8835,N_6974);
xor U10634 (N_10634,N_8722,N_8728);
nor U10635 (N_10635,N_7256,N_6529);
xnor U10636 (N_10636,N_6549,N_7351);
xnor U10637 (N_10637,N_9332,N_6698);
xnor U10638 (N_10638,N_6788,N_7368);
nor U10639 (N_10639,N_7129,N_9105);
xnor U10640 (N_10640,N_9071,N_8806);
or U10641 (N_10641,N_8734,N_9031);
or U10642 (N_10642,N_8634,N_8242);
or U10643 (N_10643,N_8612,N_9326);
or U10644 (N_10644,N_8921,N_8385);
nand U10645 (N_10645,N_6821,N_8107);
xnor U10646 (N_10646,N_8494,N_9009);
nor U10647 (N_10647,N_8204,N_8765);
or U10648 (N_10648,N_7625,N_6424);
or U10649 (N_10649,N_9188,N_6608);
and U10650 (N_10650,N_8946,N_8749);
xnor U10651 (N_10651,N_7010,N_6346);
nor U10652 (N_10652,N_8701,N_9196);
or U10653 (N_10653,N_7149,N_6940);
or U10654 (N_10654,N_6367,N_7619);
or U10655 (N_10655,N_9184,N_7107);
and U10656 (N_10656,N_7783,N_6853);
and U10657 (N_10657,N_7901,N_7853);
and U10658 (N_10658,N_7064,N_8463);
and U10659 (N_10659,N_6605,N_7610);
or U10660 (N_10660,N_7174,N_8103);
or U10661 (N_10661,N_8787,N_6264);
nor U10662 (N_10662,N_7187,N_6922);
or U10663 (N_10663,N_7555,N_8781);
and U10664 (N_10664,N_8644,N_8537);
or U10665 (N_10665,N_8456,N_6365);
or U10666 (N_10666,N_9010,N_8628);
and U10667 (N_10667,N_8697,N_7284);
nor U10668 (N_10668,N_7462,N_7930);
nand U10669 (N_10669,N_6309,N_8777);
or U10670 (N_10670,N_6903,N_9354);
nand U10671 (N_10671,N_9287,N_7390);
or U10672 (N_10672,N_6741,N_8864);
xnor U10673 (N_10673,N_8026,N_8626);
and U10674 (N_10674,N_7269,N_6965);
nor U10675 (N_10675,N_6347,N_7977);
and U10676 (N_10676,N_7130,N_6544);
or U10677 (N_10677,N_7359,N_6869);
nand U10678 (N_10678,N_6355,N_6752);
nor U10679 (N_10679,N_7155,N_7212);
nand U10680 (N_10680,N_8573,N_8461);
or U10681 (N_10681,N_9227,N_7628);
or U10682 (N_10682,N_7027,N_9205);
or U10683 (N_10683,N_8135,N_8933);
or U10684 (N_10684,N_6990,N_6886);
or U10685 (N_10685,N_6395,N_7754);
or U10686 (N_10686,N_8881,N_6826);
or U10687 (N_10687,N_7160,N_8896);
nand U10688 (N_10688,N_6589,N_7806);
or U10689 (N_10689,N_7941,N_6476);
xor U10690 (N_10690,N_6510,N_9256);
nor U10691 (N_10691,N_6881,N_8138);
xnor U10692 (N_10692,N_7627,N_9107);
or U10693 (N_10693,N_8859,N_7469);
and U10694 (N_10694,N_9006,N_7724);
nand U10695 (N_10695,N_7282,N_8484);
nand U10696 (N_10696,N_7530,N_7175);
or U10697 (N_10697,N_8556,N_6331);
nor U10698 (N_10698,N_9074,N_9094);
xor U10699 (N_10699,N_6268,N_8407);
and U10700 (N_10700,N_6548,N_8254);
xnor U10701 (N_10701,N_6994,N_7553);
or U10702 (N_10702,N_8949,N_7707);
xnor U10703 (N_10703,N_7717,N_7044);
nand U10704 (N_10704,N_9127,N_6258);
or U10705 (N_10705,N_8658,N_6459);
nor U10706 (N_10706,N_9367,N_7210);
or U10707 (N_10707,N_6276,N_6294);
or U10708 (N_10708,N_7658,N_7232);
xor U10709 (N_10709,N_8373,N_6519);
or U10710 (N_10710,N_7498,N_8454);
xor U10711 (N_10711,N_6450,N_7073);
and U10712 (N_10712,N_7209,N_9048);
or U10713 (N_10713,N_6393,N_8805);
or U10714 (N_10714,N_7231,N_6795);
xor U10715 (N_10715,N_7287,N_8725);
or U10716 (N_10716,N_6862,N_8797);
nor U10717 (N_10717,N_7020,N_7288);
and U10718 (N_10718,N_7363,N_6623);
or U10719 (N_10719,N_8249,N_6680);
or U10720 (N_10720,N_7636,N_7220);
and U10721 (N_10721,N_7066,N_7136);
nor U10722 (N_10722,N_6997,N_8223);
nor U10723 (N_10723,N_8437,N_6577);
nand U10724 (N_10724,N_8629,N_7983);
and U10725 (N_10725,N_7948,N_7866);
and U10726 (N_10726,N_8994,N_6701);
nand U10727 (N_10727,N_8743,N_8899);
and U10728 (N_10728,N_7515,N_8719);
and U10729 (N_10729,N_6356,N_8708);
nand U10730 (N_10730,N_7439,N_6335);
xor U10731 (N_10731,N_6664,N_7408);
and U10732 (N_10732,N_7881,N_6464);
nand U10733 (N_10733,N_8275,N_6381);
nand U10734 (N_10734,N_7007,N_8081);
xnor U10735 (N_10735,N_7346,N_7385);
or U10736 (N_10736,N_8840,N_8465);
or U10737 (N_10737,N_7461,N_9258);
or U10738 (N_10738,N_8800,N_6639);
or U10739 (N_10739,N_7426,N_8934);
or U10740 (N_10740,N_8973,N_8668);
xor U10741 (N_10741,N_8961,N_7593);
and U10742 (N_10742,N_8314,N_6971);
or U10743 (N_10743,N_6769,N_8662);
xnor U10744 (N_10744,N_7943,N_8981);
nor U10745 (N_10745,N_8423,N_8553);
nor U10746 (N_10746,N_8771,N_8678);
and U10747 (N_10747,N_8974,N_7290);
and U10748 (N_10748,N_7542,N_6615);
nor U10749 (N_10749,N_7057,N_7424);
nand U10750 (N_10750,N_8056,N_6950);
nand U10751 (N_10751,N_6282,N_6460);
or U10752 (N_10752,N_7226,N_9282);
and U10753 (N_10753,N_7490,N_7267);
nor U10754 (N_10754,N_9269,N_6695);
or U10755 (N_10755,N_9022,N_8691);
and U10756 (N_10756,N_6880,N_8033);
or U10757 (N_10757,N_6508,N_7778);
or U10758 (N_10758,N_9178,N_8029);
xnor U10759 (N_10759,N_6452,N_7528);
or U10760 (N_10760,N_8844,N_8551);
or U10761 (N_10761,N_7567,N_7023);
nor U10762 (N_10762,N_8908,N_6721);
or U10763 (N_10763,N_7072,N_7217);
and U10764 (N_10764,N_9283,N_7694);
and U10765 (N_10765,N_7097,N_8132);
and U10766 (N_10766,N_7923,N_9115);
nor U10767 (N_10767,N_6397,N_7341);
nand U10768 (N_10768,N_6988,N_9281);
xnor U10769 (N_10769,N_9111,N_9298);
xnor U10770 (N_10770,N_7571,N_8159);
nand U10771 (N_10771,N_6789,N_6525);
nor U10772 (N_10772,N_7089,N_8216);
or U10773 (N_10773,N_7430,N_7449);
nor U10774 (N_10774,N_7434,N_9160);
xnor U10775 (N_10775,N_7743,N_9360);
or U10776 (N_10776,N_6507,N_6361);
and U10777 (N_10777,N_8541,N_6627);
xor U10778 (N_10778,N_9138,N_9328);
or U10779 (N_10779,N_8914,N_8984);
and U10780 (N_10780,N_7298,N_7740);
and U10781 (N_10781,N_8421,N_9187);
or U10782 (N_10782,N_8430,N_8700);
xnor U10783 (N_10783,N_9169,N_7630);
nand U10784 (N_10784,N_7937,N_8315);
or U10785 (N_10785,N_8779,N_6261);
xor U10786 (N_10786,N_6967,N_7229);
xor U10787 (N_10787,N_7416,N_6759);
nor U10788 (N_10788,N_7877,N_7938);
nand U10789 (N_10789,N_8704,N_8059);
or U10790 (N_10790,N_7550,N_7165);
nand U10791 (N_10791,N_7595,N_6326);
xor U10792 (N_10792,N_6816,N_7771);
xnor U10793 (N_10793,N_7896,N_9097);
nand U10794 (N_10794,N_7119,N_8401);
xnor U10795 (N_10795,N_8535,N_6313);
nor U10796 (N_10796,N_7071,N_7432);
nor U10797 (N_10797,N_7796,N_8590);
and U10798 (N_10798,N_8424,N_6852);
nand U10799 (N_10799,N_8595,N_7052);
xor U10800 (N_10800,N_8068,N_9120);
or U10801 (N_10801,N_7270,N_8866);
xnor U10802 (N_10802,N_6704,N_6466);
nand U10803 (N_10803,N_6576,N_8670);
and U10804 (N_10804,N_7880,N_9266);
nor U10805 (N_10805,N_7011,N_8246);
nand U10806 (N_10806,N_8874,N_8566);
xnor U10807 (N_10807,N_6678,N_7691);
nand U10808 (N_10808,N_8855,N_8895);
nor U10809 (N_10809,N_8907,N_8243);
nand U10810 (N_10810,N_7277,N_8398);
or U10811 (N_10811,N_7599,N_7600);
or U10812 (N_10812,N_8041,N_9305);
nor U10813 (N_10813,N_8021,N_6674);
or U10814 (N_10814,N_7678,N_6407);
nand U10815 (N_10815,N_9194,N_6870);
and U10816 (N_10816,N_6885,N_8959);
or U10817 (N_10817,N_7283,N_7909);
nor U10818 (N_10818,N_7445,N_7501);
nor U10819 (N_10819,N_9219,N_8778);
nor U10820 (N_10820,N_8952,N_7594);
nand U10821 (N_10821,N_7084,N_7681);
nor U10822 (N_10822,N_8808,N_7389);
and U10823 (N_10823,N_7759,N_8599);
nand U10824 (N_10824,N_6819,N_9154);
nand U10825 (N_10825,N_6379,N_7275);
nand U10826 (N_10826,N_8345,N_6901);
nand U10827 (N_10827,N_9179,N_9301);
xor U10828 (N_10828,N_7419,N_8230);
and U10829 (N_10829,N_6802,N_8119);
nor U10830 (N_10830,N_6528,N_6908);
or U10831 (N_10831,N_6785,N_7438);
xnor U10832 (N_10832,N_7814,N_8982);
xnor U10833 (N_10833,N_8645,N_6295);
nor U10834 (N_10834,N_7494,N_7577);
and U10835 (N_10835,N_7914,N_7823);
and U10836 (N_10836,N_8288,N_6993);
or U10837 (N_10837,N_8854,N_7534);
nand U10838 (N_10838,N_7860,N_8100);
nor U10839 (N_10839,N_6766,N_8037);
or U10840 (N_10840,N_8604,N_8837);
or U10841 (N_10841,N_7485,N_9272);
nand U10842 (N_10842,N_7414,N_6333);
xnor U10843 (N_10843,N_8133,N_7345);
xor U10844 (N_10844,N_7166,N_9334);
nor U10845 (N_10845,N_7570,N_9351);
xor U10846 (N_10846,N_8711,N_8317);
or U10847 (N_10847,N_8426,N_8040);
and U10848 (N_10848,N_6915,N_7657);
nor U10849 (N_10849,N_6973,N_8189);
and U10850 (N_10850,N_6443,N_8210);
nor U10851 (N_10851,N_6442,N_7765);
xor U10852 (N_10852,N_6374,N_9152);
or U10853 (N_10853,N_6275,N_7824);
nand U10854 (N_10854,N_7254,N_7712);
xor U10855 (N_10855,N_7651,N_8252);
xor U10856 (N_10856,N_9295,N_6882);
and U10857 (N_10857,N_7374,N_9206);
nand U10858 (N_10858,N_9342,N_7032);
or U10859 (N_10859,N_8444,N_6745);
xnor U10860 (N_10860,N_9209,N_6413);
nor U10861 (N_10861,N_7356,N_6624);
and U10862 (N_10862,N_9221,N_6416);
or U10863 (N_10863,N_9195,N_7021);
xnor U10864 (N_10864,N_8497,N_8342);
and U10865 (N_10865,N_7551,N_6521);
xor U10866 (N_10866,N_9092,N_6655);
nor U10867 (N_10867,N_8856,N_8309);
xnor U10868 (N_10868,N_6297,N_6358);
and U10869 (N_10869,N_8912,N_7081);
or U10870 (N_10870,N_6811,N_8457);
or U10871 (N_10871,N_6714,N_6629);
nor U10872 (N_10872,N_7660,N_6861);
and U10873 (N_10873,N_7588,N_7875);
nor U10874 (N_10874,N_8772,N_8279);
and U10875 (N_10875,N_8869,N_7404);
nand U10876 (N_10876,N_9117,N_9275);
and U10877 (N_10877,N_6522,N_7911);
nand U10878 (N_10878,N_8598,N_8929);
nor U10879 (N_10879,N_6964,N_7355);
or U10880 (N_10880,N_8218,N_7975);
or U10881 (N_10881,N_9224,N_8548);
and U10882 (N_10882,N_7572,N_8817);
nor U10883 (N_10883,N_8069,N_8070);
and U10884 (N_10884,N_8334,N_7813);
nand U10885 (N_10885,N_6562,N_6328);
or U10886 (N_10886,N_9371,N_6555);
or U10887 (N_10887,N_7962,N_8193);
nor U10888 (N_10888,N_7239,N_8762);
xnor U10889 (N_10889,N_8226,N_7568);
nor U10890 (N_10890,N_9207,N_7354);
nand U10891 (N_10891,N_8354,N_6351);
and U10892 (N_10892,N_7620,N_9235);
nor U10893 (N_10893,N_6591,N_8098);
or U10894 (N_10894,N_8603,N_6253);
nand U10895 (N_10895,N_8353,N_8413);
nor U10896 (N_10896,N_6765,N_7370);
nor U10897 (N_10897,N_6455,N_7225);
nand U10898 (N_10898,N_8592,N_7787);
and U10899 (N_10899,N_6895,N_8616);
or U10900 (N_10900,N_7673,N_8757);
xor U10901 (N_10901,N_9056,N_7872);
or U10902 (N_10902,N_8791,N_7378);
nand U10903 (N_10903,N_6976,N_7292);
nand U10904 (N_10904,N_7338,N_7698);
nor U10905 (N_10905,N_6539,N_8305);
and U10906 (N_10906,N_7235,N_8960);
and U10907 (N_10907,N_6580,N_8518);
nor U10908 (N_10908,N_7831,N_6259);
and U10909 (N_10909,N_8508,N_7900);
nor U10910 (N_10910,N_8928,N_8674);
nor U10911 (N_10911,N_8181,N_7296);
or U10912 (N_10912,N_7297,N_8459);
or U10913 (N_10913,N_8445,N_8917);
or U10914 (N_10914,N_7377,N_6610);
and U10915 (N_10915,N_9333,N_6984);
nand U10916 (N_10916,N_7816,N_6305);
and U10917 (N_10917,N_6469,N_6435);
nor U10918 (N_10918,N_7546,N_8977);
nand U10919 (N_10919,N_8337,N_7512);
and U10920 (N_10920,N_9145,N_8651);
nand U10921 (N_10921,N_7676,N_8113);
xnor U10922 (N_10922,N_8118,N_8277);
and U10923 (N_10923,N_8485,N_6446);
and U10924 (N_10924,N_6953,N_8707);
nand U10925 (N_10925,N_8270,N_9052);
or U10926 (N_10926,N_8718,N_9320);
nor U10927 (N_10927,N_9073,N_7391);
nor U10928 (N_10928,N_6271,N_7664);
and U10929 (N_10929,N_6838,N_7031);
xnor U10930 (N_10930,N_6910,N_7985);
nand U10931 (N_10931,N_9087,N_6814);
nand U10932 (N_10932,N_9030,N_8215);
or U10933 (N_10933,N_6478,N_6694);
and U10934 (N_10934,N_8517,N_8183);
or U10935 (N_10935,N_9083,N_6504);
or U10936 (N_10936,N_7579,N_7958);
xor U10937 (N_10937,N_8253,N_8870);
nand U10938 (N_10938,N_9243,N_7847);
nand U10939 (N_10939,N_7292,N_7293);
and U10940 (N_10940,N_8646,N_7515);
and U10941 (N_10941,N_7180,N_8187);
and U10942 (N_10942,N_8560,N_8456);
or U10943 (N_10943,N_8889,N_8048);
xor U10944 (N_10944,N_8788,N_7941);
or U10945 (N_10945,N_6844,N_7480);
nor U10946 (N_10946,N_8241,N_8293);
xnor U10947 (N_10947,N_8842,N_7336);
xor U10948 (N_10948,N_7817,N_7333);
or U10949 (N_10949,N_7792,N_8764);
or U10950 (N_10950,N_7165,N_7503);
nand U10951 (N_10951,N_7490,N_6533);
or U10952 (N_10952,N_8791,N_8096);
and U10953 (N_10953,N_8115,N_6948);
xnor U10954 (N_10954,N_6583,N_6836);
nor U10955 (N_10955,N_7798,N_6574);
or U10956 (N_10956,N_7307,N_6439);
and U10957 (N_10957,N_7850,N_6861);
and U10958 (N_10958,N_7341,N_9194);
nand U10959 (N_10959,N_7223,N_8571);
nand U10960 (N_10960,N_7520,N_6728);
and U10961 (N_10961,N_9341,N_7892);
and U10962 (N_10962,N_7870,N_6421);
and U10963 (N_10963,N_6736,N_7420);
nand U10964 (N_10964,N_7473,N_9076);
xor U10965 (N_10965,N_7749,N_6687);
and U10966 (N_10966,N_8045,N_7183);
and U10967 (N_10967,N_6429,N_7422);
nor U10968 (N_10968,N_8476,N_7884);
nor U10969 (N_10969,N_7869,N_9358);
nor U10970 (N_10970,N_7317,N_7906);
xor U10971 (N_10971,N_7591,N_6982);
nor U10972 (N_10972,N_7561,N_8835);
nor U10973 (N_10973,N_6456,N_7656);
nor U10974 (N_10974,N_7706,N_7542);
nand U10975 (N_10975,N_6961,N_7680);
xnor U10976 (N_10976,N_9119,N_7278);
or U10977 (N_10977,N_8695,N_6557);
nand U10978 (N_10978,N_6632,N_8078);
nor U10979 (N_10979,N_6454,N_7515);
and U10980 (N_10980,N_8194,N_8046);
or U10981 (N_10981,N_7354,N_8766);
or U10982 (N_10982,N_9085,N_8845);
or U10983 (N_10983,N_6373,N_6531);
nand U10984 (N_10984,N_6528,N_8058);
or U10985 (N_10985,N_9044,N_9229);
nand U10986 (N_10986,N_8776,N_8774);
and U10987 (N_10987,N_7125,N_8310);
nor U10988 (N_10988,N_7688,N_8505);
nand U10989 (N_10989,N_9288,N_7097);
nand U10990 (N_10990,N_7426,N_9155);
nand U10991 (N_10991,N_6562,N_7001);
nor U10992 (N_10992,N_9289,N_7747);
nor U10993 (N_10993,N_9191,N_8463);
and U10994 (N_10994,N_7619,N_7836);
nand U10995 (N_10995,N_8861,N_6916);
nor U10996 (N_10996,N_6450,N_8602);
nor U10997 (N_10997,N_6795,N_8700);
or U10998 (N_10998,N_8625,N_8987);
nand U10999 (N_10999,N_6611,N_9316);
xnor U11000 (N_11000,N_6416,N_6697);
nand U11001 (N_11001,N_7079,N_9258);
nand U11002 (N_11002,N_8900,N_6358);
and U11003 (N_11003,N_8100,N_8257);
or U11004 (N_11004,N_8363,N_8719);
or U11005 (N_11005,N_8654,N_9374);
nor U11006 (N_11006,N_6881,N_9242);
or U11007 (N_11007,N_8658,N_7644);
xnor U11008 (N_11008,N_8043,N_7063);
or U11009 (N_11009,N_8497,N_6850);
xnor U11010 (N_11010,N_9361,N_6308);
nand U11011 (N_11011,N_6765,N_9028);
or U11012 (N_11012,N_8005,N_8089);
and U11013 (N_11013,N_9354,N_8486);
nor U11014 (N_11014,N_7482,N_8327);
nand U11015 (N_11015,N_6532,N_6861);
and U11016 (N_11016,N_6958,N_6855);
or U11017 (N_11017,N_6973,N_7265);
nand U11018 (N_11018,N_8641,N_8883);
xnor U11019 (N_11019,N_8953,N_8775);
nor U11020 (N_11020,N_7686,N_8473);
nor U11021 (N_11021,N_7299,N_8502);
nor U11022 (N_11022,N_9049,N_6568);
xor U11023 (N_11023,N_6861,N_7178);
and U11024 (N_11024,N_8650,N_7339);
nor U11025 (N_11025,N_6442,N_8648);
or U11026 (N_11026,N_6785,N_9194);
or U11027 (N_11027,N_7620,N_6334);
or U11028 (N_11028,N_8529,N_7419);
or U11029 (N_11029,N_8333,N_6552);
nand U11030 (N_11030,N_7705,N_9215);
and U11031 (N_11031,N_6664,N_7046);
and U11032 (N_11032,N_7707,N_8429);
or U11033 (N_11033,N_7380,N_8855);
and U11034 (N_11034,N_7945,N_9173);
and U11035 (N_11035,N_8784,N_7144);
or U11036 (N_11036,N_9273,N_8507);
nor U11037 (N_11037,N_8264,N_8199);
nand U11038 (N_11038,N_6844,N_8776);
and U11039 (N_11039,N_6524,N_6759);
nor U11040 (N_11040,N_7312,N_8365);
xnor U11041 (N_11041,N_9314,N_7430);
or U11042 (N_11042,N_6821,N_8191);
and U11043 (N_11043,N_9190,N_8202);
nand U11044 (N_11044,N_8783,N_8506);
nand U11045 (N_11045,N_9046,N_8858);
xor U11046 (N_11046,N_6347,N_6927);
and U11047 (N_11047,N_7606,N_9106);
nor U11048 (N_11048,N_8427,N_7619);
and U11049 (N_11049,N_7621,N_8834);
and U11050 (N_11050,N_6718,N_8638);
or U11051 (N_11051,N_8474,N_7757);
nor U11052 (N_11052,N_9147,N_8451);
nor U11053 (N_11053,N_7413,N_6850);
and U11054 (N_11054,N_8442,N_8998);
nor U11055 (N_11055,N_8737,N_8304);
or U11056 (N_11056,N_8704,N_6297);
nor U11057 (N_11057,N_7479,N_7015);
xor U11058 (N_11058,N_7574,N_6942);
or U11059 (N_11059,N_6253,N_8763);
nand U11060 (N_11060,N_9024,N_6307);
nor U11061 (N_11061,N_6719,N_8817);
nand U11062 (N_11062,N_9233,N_8760);
nor U11063 (N_11063,N_8053,N_8882);
or U11064 (N_11064,N_7053,N_8996);
xor U11065 (N_11065,N_7643,N_9065);
and U11066 (N_11066,N_9262,N_7053);
or U11067 (N_11067,N_6292,N_8099);
nor U11068 (N_11068,N_6605,N_7914);
and U11069 (N_11069,N_8153,N_8366);
or U11070 (N_11070,N_9151,N_8503);
nor U11071 (N_11071,N_6551,N_6768);
or U11072 (N_11072,N_7965,N_9124);
nor U11073 (N_11073,N_7919,N_7739);
nor U11074 (N_11074,N_9204,N_7132);
nor U11075 (N_11075,N_8393,N_9100);
or U11076 (N_11076,N_6766,N_8076);
and U11077 (N_11077,N_8436,N_7413);
xnor U11078 (N_11078,N_6444,N_9266);
xor U11079 (N_11079,N_8611,N_6325);
or U11080 (N_11080,N_7753,N_7551);
nor U11081 (N_11081,N_6589,N_9366);
and U11082 (N_11082,N_8371,N_8612);
nor U11083 (N_11083,N_8695,N_7249);
nand U11084 (N_11084,N_7877,N_7740);
nand U11085 (N_11085,N_9247,N_7293);
nand U11086 (N_11086,N_8107,N_7558);
and U11087 (N_11087,N_7233,N_8435);
and U11088 (N_11088,N_7877,N_7634);
or U11089 (N_11089,N_6743,N_7525);
or U11090 (N_11090,N_8511,N_6276);
xor U11091 (N_11091,N_9163,N_8405);
and U11092 (N_11092,N_8111,N_7932);
and U11093 (N_11093,N_8464,N_7075);
nand U11094 (N_11094,N_7217,N_9044);
or U11095 (N_11095,N_7944,N_9089);
xor U11096 (N_11096,N_7391,N_7916);
nand U11097 (N_11097,N_6915,N_7332);
or U11098 (N_11098,N_7801,N_7617);
xor U11099 (N_11099,N_8206,N_9065);
nor U11100 (N_11100,N_9223,N_7158);
nor U11101 (N_11101,N_9057,N_9206);
and U11102 (N_11102,N_9230,N_7636);
nand U11103 (N_11103,N_8492,N_8149);
nand U11104 (N_11104,N_8878,N_8316);
xnor U11105 (N_11105,N_9149,N_7085);
nor U11106 (N_11106,N_6912,N_8415);
nor U11107 (N_11107,N_9093,N_7261);
xor U11108 (N_11108,N_8865,N_6768);
xor U11109 (N_11109,N_7029,N_8415);
or U11110 (N_11110,N_8239,N_7701);
nor U11111 (N_11111,N_7335,N_9073);
xnor U11112 (N_11112,N_7476,N_6969);
or U11113 (N_11113,N_6630,N_7121);
nor U11114 (N_11114,N_6904,N_8624);
or U11115 (N_11115,N_7522,N_9023);
and U11116 (N_11116,N_8734,N_8850);
nor U11117 (N_11117,N_8263,N_6846);
and U11118 (N_11118,N_7793,N_6744);
and U11119 (N_11119,N_8375,N_8896);
nand U11120 (N_11120,N_8984,N_8097);
or U11121 (N_11121,N_8666,N_9048);
nand U11122 (N_11122,N_9300,N_7039);
nand U11123 (N_11123,N_8950,N_7305);
xor U11124 (N_11124,N_9122,N_6386);
nor U11125 (N_11125,N_8419,N_8034);
or U11126 (N_11126,N_7500,N_6933);
nor U11127 (N_11127,N_8189,N_7214);
nand U11128 (N_11128,N_6991,N_8913);
or U11129 (N_11129,N_7035,N_8647);
or U11130 (N_11130,N_6823,N_6487);
or U11131 (N_11131,N_7634,N_7689);
and U11132 (N_11132,N_8863,N_7598);
or U11133 (N_11133,N_6743,N_9299);
or U11134 (N_11134,N_6891,N_8598);
xor U11135 (N_11135,N_7289,N_7374);
and U11136 (N_11136,N_7026,N_6947);
xnor U11137 (N_11137,N_7885,N_6978);
nor U11138 (N_11138,N_7777,N_8084);
and U11139 (N_11139,N_9308,N_8628);
nor U11140 (N_11140,N_8104,N_6868);
nor U11141 (N_11141,N_7304,N_8286);
xor U11142 (N_11142,N_8835,N_8052);
xor U11143 (N_11143,N_6499,N_8672);
xor U11144 (N_11144,N_8823,N_8336);
or U11145 (N_11145,N_7478,N_7886);
nor U11146 (N_11146,N_7962,N_7756);
and U11147 (N_11147,N_7153,N_8251);
nor U11148 (N_11148,N_7868,N_7687);
nand U11149 (N_11149,N_7035,N_7884);
nor U11150 (N_11150,N_7228,N_6831);
or U11151 (N_11151,N_6414,N_8602);
or U11152 (N_11152,N_8892,N_8899);
xor U11153 (N_11153,N_6475,N_7703);
nand U11154 (N_11154,N_7778,N_7366);
and U11155 (N_11155,N_8890,N_9177);
and U11156 (N_11156,N_7260,N_7123);
nand U11157 (N_11157,N_8292,N_6699);
nand U11158 (N_11158,N_7977,N_7502);
nand U11159 (N_11159,N_6659,N_9325);
nand U11160 (N_11160,N_8259,N_8662);
nor U11161 (N_11161,N_9215,N_8789);
nand U11162 (N_11162,N_6366,N_8096);
and U11163 (N_11163,N_7825,N_8384);
nand U11164 (N_11164,N_7842,N_7597);
or U11165 (N_11165,N_8207,N_6635);
xnor U11166 (N_11166,N_7704,N_6800);
xnor U11167 (N_11167,N_8706,N_8100);
or U11168 (N_11168,N_6515,N_6724);
nor U11169 (N_11169,N_9103,N_6661);
xor U11170 (N_11170,N_7713,N_6668);
nand U11171 (N_11171,N_8460,N_7360);
nand U11172 (N_11172,N_8638,N_6522);
or U11173 (N_11173,N_8779,N_7200);
and U11174 (N_11174,N_8683,N_8624);
nor U11175 (N_11175,N_8457,N_7732);
nor U11176 (N_11176,N_6703,N_7654);
and U11177 (N_11177,N_8035,N_8131);
nand U11178 (N_11178,N_6646,N_8526);
and U11179 (N_11179,N_8285,N_8126);
nand U11180 (N_11180,N_6869,N_6617);
nor U11181 (N_11181,N_7058,N_8689);
and U11182 (N_11182,N_9052,N_8596);
or U11183 (N_11183,N_6866,N_7392);
or U11184 (N_11184,N_7831,N_6536);
or U11185 (N_11185,N_8936,N_6962);
nor U11186 (N_11186,N_8121,N_8452);
nor U11187 (N_11187,N_6528,N_7558);
and U11188 (N_11188,N_8536,N_8844);
xor U11189 (N_11189,N_6639,N_9226);
xnor U11190 (N_11190,N_7558,N_8328);
or U11191 (N_11191,N_7934,N_7408);
or U11192 (N_11192,N_6619,N_7405);
nand U11193 (N_11193,N_9035,N_6394);
nor U11194 (N_11194,N_8498,N_8712);
and U11195 (N_11195,N_8751,N_8678);
or U11196 (N_11196,N_6314,N_8689);
nor U11197 (N_11197,N_7257,N_9373);
or U11198 (N_11198,N_6770,N_7524);
or U11199 (N_11199,N_7415,N_8528);
or U11200 (N_11200,N_8193,N_8069);
xnor U11201 (N_11201,N_7008,N_9032);
and U11202 (N_11202,N_8617,N_7415);
nand U11203 (N_11203,N_9173,N_7656);
or U11204 (N_11204,N_8048,N_8616);
nand U11205 (N_11205,N_8187,N_6910);
and U11206 (N_11206,N_8557,N_8788);
nor U11207 (N_11207,N_8111,N_6293);
and U11208 (N_11208,N_7941,N_8371);
xor U11209 (N_11209,N_8981,N_8224);
nand U11210 (N_11210,N_7739,N_6499);
or U11211 (N_11211,N_8512,N_8266);
or U11212 (N_11212,N_8059,N_7153);
nand U11213 (N_11213,N_8517,N_8712);
nor U11214 (N_11214,N_6374,N_6418);
or U11215 (N_11215,N_8788,N_8448);
and U11216 (N_11216,N_8395,N_6509);
and U11217 (N_11217,N_8773,N_8593);
nor U11218 (N_11218,N_8861,N_7294);
and U11219 (N_11219,N_9074,N_8602);
xnor U11220 (N_11220,N_7424,N_7394);
or U11221 (N_11221,N_8993,N_6354);
nor U11222 (N_11222,N_6601,N_8468);
nor U11223 (N_11223,N_8647,N_6750);
or U11224 (N_11224,N_7093,N_8987);
xor U11225 (N_11225,N_7341,N_8541);
nand U11226 (N_11226,N_7710,N_8511);
nand U11227 (N_11227,N_7180,N_6901);
nor U11228 (N_11228,N_9084,N_7182);
and U11229 (N_11229,N_9074,N_9057);
or U11230 (N_11230,N_6997,N_8620);
nand U11231 (N_11231,N_6854,N_6879);
and U11232 (N_11232,N_7583,N_8098);
and U11233 (N_11233,N_8349,N_8085);
xor U11234 (N_11234,N_8142,N_7367);
nor U11235 (N_11235,N_7837,N_8025);
nand U11236 (N_11236,N_8328,N_8329);
and U11237 (N_11237,N_8290,N_6596);
xor U11238 (N_11238,N_6775,N_8727);
and U11239 (N_11239,N_6673,N_9275);
or U11240 (N_11240,N_7891,N_6475);
and U11241 (N_11241,N_8686,N_6957);
nand U11242 (N_11242,N_7386,N_7046);
or U11243 (N_11243,N_9100,N_8818);
xnor U11244 (N_11244,N_9305,N_8809);
xor U11245 (N_11245,N_8314,N_8155);
or U11246 (N_11246,N_7980,N_7757);
nor U11247 (N_11247,N_8437,N_7410);
xnor U11248 (N_11248,N_7794,N_6414);
nand U11249 (N_11249,N_7862,N_6910);
nand U11250 (N_11250,N_9165,N_8463);
xnor U11251 (N_11251,N_6354,N_7928);
nand U11252 (N_11252,N_7969,N_6671);
nor U11253 (N_11253,N_7151,N_7077);
and U11254 (N_11254,N_6705,N_8969);
xnor U11255 (N_11255,N_7568,N_6303);
xor U11256 (N_11256,N_7297,N_6633);
or U11257 (N_11257,N_8369,N_9134);
and U11258 (N_11258,N_8275,N_8159);
nor U11259 (N_11259,N_9206,N_7645);
xnor U11260 (N_11260,N_6788,N_6318);
xnor U11261 (N_11261,N_6744,N_7987);
nor U11262 (N_11262,N_7539,N_6900);
nand U11263 (N_11263,N_9193,N_9177);
or U11264 (N_11264,N_7665,N_9003);
and U11265 (N_11265,N_7625,N_9213);
and U11266 (N_11266,N_8652,N_8896);
nor U11267 (N_11267,N_8206,N_8133);
nor U11268 (N_11268,N_8704,N_8741);
and U11269 (N_11269,N_7172,N_7046);
nor U11270 (N_11270,N_8001,N_8605);
nor U11271 (N_11271,N_9331,N_6367);
or U11272 (N_11272,N_6723,N_6981);
or U11273 (N_11273,N_8200,N_8482);
xor U11274 (N_11274,N_8847,N_7996);
nor U11275 (N_11275,N_7766,N_8987);
and U11276 (N_11276,N_9069,N_6337);
xnor U11277 (N_11277,N_9267,N_8672);
and U11278 (N_11278,N_7735,N_6958);
nor U11279 (N_11279,N_9297,N_7235);
nand U11280 (N_11280,N_8124,N_6509);
nand U11281 (N_11281,N_6647,N_7551);
and U11282 (N_11282,N_6870,N_6368);
or U11283 (N_11283,N_7814,N_6976);
nor U11284 (N_11284,N_8021,N_7630);
and U11285 (N_11285,N_7718,N_7109);
or U11286 (N_11286,N_8266,N_8389);
xnor U11287 (N_11287,N_8267,N_7853);
nand U11288 (N_11288,N_7469,N_8843);
nand U11289 (N_11289,N_7701,N_6679);
and U11290 (N_11290,N_6943,N_7018);
xnor U11291 (N_11291,N_7154,N_8732);
or U11292 (N_11292,N_8843,N_8306);
xnor U11293 (N_11293,N_7286,N_7951);
and U11294 (N_11294,N_8313,N_7372);
or U11295 (N_11295,N_7874,N_7005);
nor U11296 (N_11296,N_6802,N_7720);
xor U11297 (N_11297,N_9046,N_6327);
and U11298 (N_11298,N_8006,N_6633);
nand U11299 (N_11299,N_8065,N_7690);
xor U11300 (N_11300,N_8709,N_9329);
nand U11301 (N_11301,N_9288,N_9103);
and U11302 (N_11302,N_7345,N_9317);
nand U11303 (N_11303,N_8171,N_7973);
or U11304 (N_11304,N_7918,N_9160);
or U11305 (N_11305,N_7626,N_7115);
xnor U11306 (N_11306,N_6858,N_9089);
or U11307 (N_11307,N_9329,N_6958);
and U11308 (N_11308,N_8326,N_6411);
nor U11309 (N_11309,N_8801,N_6869);
and U11310 (N_11310,N_6689,N_9233);
xor U11311 (N_11311,N_7756,N_6568);
nand U11312 (N_11312,N_6697,N_7140);
nor U11313 (N_11313,N_6698,N_8865);
nor U11314 (N_11314,N_6585,N_7669);
nor U11315 (N_11315,N_6576,N_7322);
and U11316 (N_11316,N_8464,N_6617);
nor U11317 (N_11317,N_8918,N_7301);
xor U11318 (N_11318,N_7926,N_8413);
xor U11319 (N_11319,N_9302,N_9184);
or U11320 (N_11320,N_7470,N_7962);
nand U11321 (N_11321,N_7875,N_8676);
or U11322 (N_11322,N_8450,N_7783);
or U11323 (N_11323,N_8433,N_8589);
or U11324 (N_11324,N_8445,N_7986);
nand U11325 (N_11325,N_8809,N_8296);
xnor U11326 (N_11326,N_8706,N_7892);
nor U11327 (N_11327,N_8487,N_8313);
nand U11328 (N_11328,N_7872,N_8640);
nand U11329 (N_11329,N_7306,N_8457);
nor U11330 (N_11330,N_8379,N_7932);
xor U11331 (N_11331,N_8900,N_7796);
nor U11332 (N_11332,N_8023,N_9296);
and U11333 (N_11333,N_7063,N_9361);
or U11334 (N_11334,N_8112,N_8126);
xnor U11335 (N_11335,N_8631,N_8208);
or U11336 (N_11336,N_6798,N_9040);
nor U11337 (N_11337,N_9337,N_9280);
nand U11338 (N_11338,N_7645,N_8512);
or U11339 (N_11339,N_7399,N_9097);
or U11340 (N_11340,N_8881,N_7789);
or U11341 (N_11341,N_8381,N_8573);
or U11342 (N_11342,N_7798,N_9090);
and U11343 (N_11343,N_7499,N_7019);
xnor U11344 (N_11344,N_6372,N_8765);
xnor U11345 (N_11345,N_7383,N_8021);
and U11346 (N_11346,N_7833,N_7973);
nor U11347 (N_11347,N_8860,N_7448);
and U11348 (N_11348,N_6573,N_8327);
nand U11349 (N_11349,N_8759,N_6485);
xnor U11350 (N_11350,N_7413,N_6698);
and U11351 (N_11351,N_9132,N_7562);
nor U11352 (N_11352,N_6938,N_7158);
nand U11353 (N_11353,N_7687,N_7611);
and U11354 (N_11354,N_8245,N_8104);
nand U11355 (N_11355,N_8255,N_8595);
xor U11356 (N_11356,N_7099,N_6627);
and U11357 (N_11357,N_7712,N_8885);
and U11358 (N_11358,N_7339,N_9129);
nor U11359 (N_11359,N_7516,N_6878);
nor U11360 (N_11360,N_9368,N_6899);
nand U11361 (N_11361,N_6974,N_7260);
and U11362 (N_11362,N_6373,N_7074);
xnor U11363 (N_11363,N_7999,N_6824);
xnor U11364 (N_11364,N_7536,N_8748);
and U11365 (N_11365,N_7549,N_8958);
xnor U11366 (N_11366,N_7633,N_8902);
xor U11367 (N_11367,N_6826,N_8986);
xnor U11368 (N_11368,N_6714,N_7286);
xnor U11369 (N_11369,N_7252,N_8672);
or U11370 (N_11370,N_7101,N_6713);
nand U11371 (N_11371,N_9114,N_9240);
nand U11372 (N_11372,N_8709,N_9363);
and U11373 (N_11373,N_9090,N_6544);
and U11374 (N_11374,N_7464,N_8600);
xnor U11375 (N_11375,N_8067,N_7508);
nor U11376 (N_11376,N_9325,N_6499);
or U11377 (N_11377,N_8972,N_9203);
or U11378 (N_11378,N_6700,N_8434);
nand U11379 (N_11379,N_9036,N_6926);
or U11380 (N_11380,N_7187,N_6701);
and U11381 (N_11381,N_8399,N_7644);
nor U11382 (N_11382,N_7162,N_6528);
nor U11383 (N_11383,N_7059,N_7484);
nand U11384 (N_11384,N_9199,N_9115);
nor U11385 (N_11385,N_7900,N_6398);
xnor U11386 (N_11386,N_6508,N_8226);
and U11387 (N_11387,N_7074,N_6850);
nor U11388 (N_11388,N_6256,N_6403);
nand U11389 (N_11389,N_6843,N_8339);
or U11390 (N_11390,N_8819,N_7617);
or U11391 (N_11391,N_8362,N_7081);
or U11392 (N_11392,N_7635,N_8844);
nand U11393 (N_11393,N_6480,N_7885);
xnor U11394 (N_11394,N_8804,N_6418);
nand U11395 (N_11395,N_6864,N_8722);
nand U11396 (N_11396,N_6899,N_6460);
nand U11397 (N_11397,N_7867,N_7444);
nand U11398 (N_11398,N_7058,N_8327);
or U11399 (N_11399,N_9338,N_9261);
xnor U11400 (N_11400,N_9015,N_8863);
and U11401 (N_11401,N_7433,N_6341);
or U11402 (N_11402,N_9247,N_7197);
or U11403 (N_11403,N_7285,N_6394);
nor U11404 (N_11404,N_8547,N_7049);
or U11405 (N_11405,N_6432,N_8369);
xnor U11406 (N_11406,N_8251,N_7987);
and U11407 (N_11407,N_6496,N_7987);
nor U11408 (N_11408,N_6319,N_6477);
or U11409 (N_11409,N_6570,N_7099);
nand U11410 (N_11410,N_6356,N_6623);
and U11411 (N_11411,N_7619,N_7844);
nand U11412 (N_11412,N_6997,N_8434);
nand U11413 (N_11413,N_9305,N_9373);
or U11414 (N_11414,N_8608,N_7053);
nor U11415 (N_11415,N_7866,N_8922);
or U11416 (N_11416,N_6562,N_9126);
or U11417 (N_11417,N_8659,N_6428);
or U11418 (N_11418,N_9125,N_8498);
or U11419 (N_11419,N_9027,N_9169);
nor U11420 (N_11420,N_6684,N_6331);
nor U11421 (N_11421,N_7821,N_8828);
nand U11422 (N_11422,N_9306,N_9058);
nor U11423 (N_11423,N_7716,N_6538);
or U11424 (N_11424,N_8431,N_7110);
or U11425 (N_11425,N_7474,N_8479);
nand U11426 (N_11426,N_7908,N_8304);
or U11427 (N_11427,N_6463,N_8539);
nor U11428 (N_11428,N_8335,N_6902);
nand U11429 (N_11429,N_9289,N_8321);
and U11430 (N_11430,N_7756,N_7118);
and U11431 (N_11431,N_8915,N_7959);
or U11432 (N_11432,N_6351,N_8910);
and U11433 (N_11433,N_8535,N_8215);
nor U11434 (N_11434,N_6610,N_8866);
nor U11435 (N_11435,N_8915,N_6343);
xnor U11436 (N_11436,N_7171,N_6597);
and U11437 (N_11437,N_6380,N_7151);
nor U11438 (N_11438,N_7083,N_8528);
nor U11439 (N_11439,N_6766,N_6442);
xor U11440 (N_11440,N_7278,N_6695);
xnor U11441 (N_11441,N_7681,N_7538);
or U11442 (N_11442,N_7074,N_6617);
xnor U11443 (N_11443,N_6611,N_7512);
or U11444 (N_11444,N_8449,N_7209);
xnor U11445 (N_11445,N_8613,N_8519);
and U11446 (N_11446,N_7051,N_7583);
nor U11447 (N_11447,N_8704,N_6543);
and U11448 (N_11448,N_6252,N_8202);
nand U11449 (N_11449,N_7036,N_7211);
xnor U11450 (N_11450,N_8455,N_7561);
nor U11451 (N_11451,N_8977,N_8292);
nor U11452 (N_11452,N_8793,N_8961);
and U11453 (N_11453,N_7421,N_8699);
xor U11454 (N_11454,N_8531,N_6819);
xor U11455 (N_11455,N_6253,N_6480);
and U11456 (N_11456,N_6550,N_6743);
and U11457 (N_11457,N_8378,N_8787);
nor U11458 (N_11458,N_7577,N_6797);
and U11459 (N_11459,N_7753,N_7933);
nand U11460 (N_11460,N_8779,N_7476);
nor U11461 (N_11461,N_8573,N_7734);
nor U11462 (N_11462,N_7819,N_6479);
and U11463 (N_11463,N_6624,N_6988);
nor U11464 (N_11464,N_8242,N_8972);
or U11465 (N_11465,N_7393,N_7161);
nand U11466 (N_11466,N_6276,N_7002);
nand U11467 (N_11467,N_7345,N_7223);
nor U11468 (N_11468,N_8914,N_8896);
and U11469 (N_11469,N_7399,N_7897);
xnor U11470 (N_11470,N_8530,N_7462);
nor U11471 (N_11471,N_7387,N_8103);
nor U11472 (N_11472,N_8805,N_7476);
xor U11473 (N_11473,N_8427,N_6633);
xnor U11474 (N_11474,N_7234,N_6423);
nor U11475 (N_11475,N_8539,N_8054);
nand U11476 (N_11476,N_7428,N_6762);
and U11477 (N_11477,N_8997,N_7493);
or U11478 (N_11478,N_7016,N_8032);
xnor U11479 (N_11479,N_8774,N_7573);
and U11480 (N_11480,N_8385,N_8225);
and U11481 (N_11481,N_7532,N_7665);
or U11482 (N_11482,N_8518,N_8809);
and U11483 (N_11483,N_6499,N_7534);
nor U11484 (N_11484,N_7746,N_8835);
or U11485 (N_11485,N_8796,N_6798);
xor U11486 (N_11486,N_6739,N_7402);
and U11487 (N_11487,N_6657,N_8056);
nor U11488 (N_11488,N_6979,N_8527);
or U11489 (N_11489,N_6272,N_8164);
xnor U11490 (N_11490,N_8035,N_8529);
or U11491 (N_11491,N_8763,N_9257);
nor U11492 (N_11492,N_9111,N_7627);
xor U11493 (N_11493,N_7218,N_7261);
nand U11494 (N_11494,N_6777,N_6395);
nor U11495 (N_11495,N_7334,N_8609);
nor U11496 (N_11496,N_8478,N_7591);
xor U11497 (N_11497,N_6931,N_8851);
and U11498 (N_11498,N_7595,N_7980);
nor U11499 (N_11499,N_7597,N_9069);
and U11500 (N_11500,N_9004,N_8709);
and U11501 (N_11501,N_9334,N_8973);
nor U11502 (N_11502,N_8243,N_6967);
xor U11503 (N_11503,N_9143,N_9097);
nor U11504 (N_11504,N_8202,N_8787);
or U11505 (N_11505,N_7534,N_7559);
nor U11506 (N_11506,N_6436,N_6892);
and U11507 (N_11507,N_8986,N_6389);
nand U11508 (N_11508,N_6670,N_7221);
xnor U11509 (N_11509,N_6475,N_7190);
and U11510 (N_11510,N_7737,N_8503);
nand U11511 (N_11511,N_8414,N_8446);
nand U11512 (N_11512,N_9081,N_6637);
and U11513 (N_11513,N_9012,N_9137);
nand U11514 (N_11514,N_8016,N_7657);
or U11515 (N_11515,N_7226,N_8811);
nor U11516 (N_11516,N_7965,N_8024);
or U11517 (N_11517,N_7748,N_6613);
nor U11518 (N_11518,N_6792,N_7544);
nand U11519 (N_11519,N_7212,N_7250);
and U11520 (N_11520,N_8662,N_7901);
and U11521 (N_11521,N_6651,N_6674);
nand U11522 (N_11522,N_8462,N_7721);
and U11523 (N_11523,N_7176,N_6936);
and U11524 (N_11524,N_8306,N_7103);
xnor U11525 (N_11525,N_8387,N_7224);
and U11526 (N_11526,N_6634,N_6989);
and U11527 (N_11527,N_9352,N_7112);
nor U11528 (N_11528,N_7018,N_9048);
and U11529 (N_11529,N_7197,N_7231);
xnor U11530 (N_11530,N_6729,N_7588);
and U11531 (N_11531,N_7643,N_6422);
or U11532 (N_11532,N_7494,N_8326);
and U11533 (N_11533,N_8655,N_6418);
xnor U11534 (N_11534,N_8527,N_7863);
and U11535 (N_11535,N_6706,N_6776);
nor U11536 (N_11536,N_9220,N_8089);
or U11537 (N_11537,N_7220,N_8466);
nand U11538 (N_11538,N_6701,N_6570);
or U11539 (N_11539,N_9308,N_8378);
nor U11540 (N_11540,N_9002,N_8569);
nor U11541 (N_11541,N_6723,N_7114);
xor U11542 (N_11542,N_8292,N_8105);
nor U11543 (N_11543,N_8392,N_9331);
and U11544 (N_11544,N_7247,N_8829);
nand U11545 (N_11545,N_9015,N_8709);
xor U11546 (N_11546,N_7277,N_6564);
xnor U11547 (N_11547,N_7439,N_7718);
nor U11548 (N_11548,N_8479,N_7941);
or U11549 (N_11549,N_6460,N_6831);
nor U11550 (N_11550,N_8118,N_7017);
xnor U11551 (N_11551,N_7097,N_7224);
nand U11552 (N_11552,N_7052,N_7162);
nor U11553 (N_11553,N_7808,N_7156);
or U11554 (N_11554,N_8575,N_7887);
or U11555 (N_11555,N_6299,N_7510);
xnor U11556 (N_11556,N_7907,N_7885);
nor U11557 (N_11557,N_9033,N_9058);
and U11558 (N_11558,N_7080,N_7399);
nor U11559 (N_11559,N_8195,N_7587);
or U11560 (N_11560,N_8508,N_6386);
nor U11561 (N_11561,N_8235,N_6898);
xor U11562 (N_11562,N_7660,N_7307);
nand U11563 (N_11563,N_7903,N_8958);
nand U11564 (N_11564,N_7377,N_6921);
nand U11565 (N_11565,N_8163,N_8627);
nand U11566 (N_11566,N_7846,N_6711);
nand U11567 (N_11567,N_7827,N_8116);
and U11568 (N_11568,N_7242,N_6355);
xor U11569 (N_11569,N_8683,N_7918);
nand U11570 (N_11570,N_8099,N_6634);
nand U11571 (N_11571,N_8552,N_8014);
or U11572 (N_11572,N_6430,N_7952);
nand U11573 (N_11573,N_6979,N_9071);
nand U11574 (N_11574,N_7151,N_8670);
nand U11575 (N_11575,N_7199,N_7840);
or U11576 (N_11576,N_7217,N_6531);
nand U11577 (N_11577,N_6304,N_8037);
and U11578 (N_11578,N_8335,N_8029);
and U11579 (N_11579,N_6854,N_6754);
or U11580 (N_11580,N_8644,N_7917);
nand U11581 (N_11581,N_7339,N_6317);
nor U11582 (N_11582,N_6255,N_8256);
nand U11583 (N_11583,N_8101,N_9256);
and U11584 (N_11584,N_8921,N_7931);
nor U11585 (N_11585,N_6610,N_7184);
or U11586 (N_11586,N_8373,N_6605);
nand U11587 (N_11587,N_8406,N_6775);
or U11588 (N_11588,N_7602,N_7783);
and U11589 (N_11589,N_6659,N_7978);
xor U11590 (N_11590,N_8012,N_8448);
xnor U11591 (N_11591,N_8661,N_8591);
nor U11592 (N_11592,N_6484,N_8554);
or U11593 (N_11593,N_6971,N_8789);
and U11594 (N_11594,N_6860,N_7190);
nand U11595 (N_11595,N_6665,N_7394);
xor U11596 (N_11596,N_8594,N_8887);
nor U11597 (N_11597,N_8461,N_8460);
nand U11598 (N_11598,N_6818,N_7354);
or U11599 (N_11599,N_7678,N_8900);
nand U11600 (N_11600,N_8393,N_6344);
and U11601 (N_11601,N_8275,N_6633);
or U11602 (N_11602,N_6694,N_6339);
or U11603 (N_11603,N_7204,N_7371);
nand U11604 (N_11604,N_8221,N_6515);
nand U11605 (N_11605,N_7214,N_9304);
xor U11606 (N_11606,N_6305,N_7334);
nor U11607 (N_11607,N_7043,N_6477);
and U11608 (N_11608,N_9210,N_9206);
or U11609 (N_11609,N_8827,N_7407);
nor U11610 (N_11610,N_8874,N_8760);
nor U11611 (N_11611,N_7633,N_6323);
xnor U11612 (N_11612,N_7928,N_8263);
or U11613 (N_11613,N_8779,N_6981);
or U11614 (N_11614,N_6901,N_6833);
xor U11615 (N_11615,N_7383,N_8476);
or U11616 (N_11616,N_6371,N_9074);
nand U11617 (N_11617,N_8675,N_8748);
or U11618 (N_11618,N_9272,N_7297);
xor U11619 (N_11619,N_7372,N_9208);
or U11620 (N_11620,N_7613,N_7942);
xnor U11621 (N_11621,N_7245,N_6985);
nor U11622 (N_11622,N_8546,N_9123);
nand U11623 (N_11623,N_6536,N_8030);
nand U11624 (N_11624,N_8024,N_8790);
and U11625 (N_11625,N_6480,N_8105);
nand U11626 (N_11626,N_6690,N_8755);
nand U11627 (N_11627,N_6635,N_6769);
nand U11628 (N_11628,N_8211,N_6548);
and U11629 (N_11629,N_6429,N_7313);
or U11630 (N_11630,N_8225,N_6666);
xnor U11631 (N_11631,N_7620,N_7094);
nand U11632 (N_11632,N_7167,N_9250);
nand U11633 (N_11633,N_8645,N_7816);
and U11634 (N_11634,N_6546,N_6756);
nand U11635 (N_11635,N_7712,N_7524);
and U11636 (N_11636,N_7674,N_9258);
or U11637 (N_11637,N_8333,N_6797);
xor U11638 (N_11638,N_8759,N_6896);
nand U11639 (N_11639,N_6847,N_7072);
nor U11640 (N_11640,N_7600,N_7994);
nand U11641 (N_11641,N_7445,N_8829);
and U11642 (N_11642,N_7364,N_8270);
xor U11643 (N_11643,N_7188,N_8238);
or U11644 (N_11644,N_8155,N_7824);
nor U11645 (N_11645,N_9139,N_7057);
xor U11646 (N_11646,N_7364,N_8262);
nand U11647 (N_11647,N_9030,N_6486);
or U11648 (N_11648,N_9011,N_6844);
or U11649 (N_11649,N_8751,N_8118);
and U11650 (N_11650,N_8797,N_8536);
xor U11651 (N_11651,N_7594,N_7146);
nor U11652 (N_11652,N_7280,N_7905);
or U11653 (N_11653,N_7696,N_9205);
and U11654 (N_11654,N_6706,N_7212);
xor U11655 (N_11655,N_7665,N_8682);
nand U11656 (N_11656,N_7401,N_9232);
xor U11657 (N_11657,N_7814,N_6690);
nor U11658 (N_11658,N_7146,N_9263);
nor U11659 (N_11659,N_8374,N_8098);
xnor U11660 (N_11660,N_6920,N_9182);
xor U11661 (N_11661,N_6520,N_8646);
nor U11662 (N_11662,N_7738,N_7187);
nor U11663 (N_11663,N_6512,N_7273);
nor U11664 (N_11664,N_7321,N_7204);
and U11665 (N_11665,N_9057,N_6545);
or U11666 (N_11666,N_9201,N_7762);
nand U11667 (N_11667,N_8521,N_7043);
or U11668 (N_11668,N_7003,N_6418);
nor U11669 (N_11669,N_8907,N_7776);
and U11670 (N_11670,N_6991,N_6485);
nand U11671 (N_11671,N_7007,N_6772);
nor U11672 (N_11672,N_8325,N_8612);
and U11673 (N_11673,N_9306,N_6470);
or U11674 (N_11674,N_9070,N_7283);
nand U11675 (N_11675,N_8067,N_8270);
nand U11676 (N_11676,N_6603,N_9187);
and U11677 (N_11677,N_8631,N_8711);
or U11678 (N_11678,N_8438,N_6678);
nand U11679 (N_11679,N_7514,N_9352);
or U11680 (N_11680,N_8681,N_6456);
and U11681 (N_11681,N_8294,N_8646);
or U11682 (N_11682,N_8704,N_8524);
or U11683 (N_11683,N_9143,N_7172);
nand U11684 (N_11684,N_7125,N_7685);
or U11685 (N_11685,N_8370,N_8427);
and U11686 (N_11686,N_6265,N_8660);
nand U11687 (N_11687,N_7768,N_8623);
nor U11688 (N_11688,N_7690,N_8627);
nor U11689 (N_11689,N_8864,N_7060);
nand U11690 (N_11690,N_6557,N_8275);
nor U11691 (N_11691,N_9112,N_6627);
and U11692 (N_11692,N_7189,N_6973);
xnor U11693 (N_11693,N_6658,N_8792);
xor U11694 (N_11694,N_7516,N_7350);
or U11695 (N_11695,N_7483,N_8583);
nand U11696 (N_11696,N_9323,N_8868);
nor U11697 (N_11697,N_7106,N_8789);
nand U11698 (N_11698,N_6801,N_6979);
xor U11699 (N_11699,N_7911,N_6779);
nor U11700 (N_11700,N_6870,N_9331);
nand U11701 (N_11701,N_8338,N_7170);
xor U11702 (N_11702,N_8587,N_6286);
xor U11703 (N_11703,N_9264,N_8301);
and U11704 (N_11704,N_6576,N_9171);
nand U11705 (N_11705,N_7343,N_7360);
xnor U11706 (N_11706,N_8584,N_8819);
and U11707 (N_11707,N_8883,N_8964);
nor U11708 (N_11708,N_8168,N_9260);
nor U11709 (N_11709,N_6753,N_7670);
and U11710 (N_11710,N_6917,N_6478);
or U11711 (N_11711,N_7398,N_8981);
nor U11712 (N_11712,N_8547,N_7521);
or U11713 (N_11713,N_6529,N_8774);
xor U11714 (N_11714,N_7970,N_6556);
and U11715 (N_11715,N_7410,N_6771);
xor U11716 (N_11716,N_7210,N_6954);
xnor U11717 (N_11717,N_6509,N_8350);
or U11718 (N_11718,N_6875,N_8054);
nor U11719 (N_11719,N_6522,N_8941);
or U11720 (N_11720,N_9295,N_8255);
nor U11721 (N_11721,N_8113,N_8655);
and U11722 (N_11722,N_7213,N_6377);
nand U11723 (N_11723,N_8070,N_6368);
and U11724 (N_11724,N_6854,N_8474);
and U11725 (N_11725,N_8066,N_8379);
and U11726 (N_11726,N_7727,N_8123);
xnor U11727 (N_11727,N_7955,N_7216);
nand U11728 (N_11728,N_7608,N_6933);
nor U11729 (N_11729,N_9050,N_7975);
and U11730 (N_11730,N_8839,N_8709);
xor U11731 (N_11731,N_7628,N_8982);
nor U11732 (N_11732,N_8234,N_7116);
nor U11733 (N_11733,N_6827,N_7368);
nand U11734 (N_11734,N_8860,N_8526);
nand U11735 (N_11735,N_6757,N_8137);
xnor U11736 (N_11736,N_7059,N_9115);
nor U11737 (N_11737,N_8879,N_6471);
xnor U11738 (N_11738,N_9041,N_9157);
xnor U11739 (N_11739,N_6745,N_7664);
and U11740 (N_11740,N_8262,N_8689);
nor U11741 (N_11741,N_7848,N_8999);
nand U11742 (N_11742,N_8035,N_8698);
and U11743 (N_11743,N_7695,N_7130);
or U11744 (N_11744,N_8038,N_6665);
nor U11745 (N_11745,N_8320,N_8038);
xor U11746 (N_11746,N_8267,N_7839);
nand U11747 (N_11747,N_7544,N_8413);
nand U11748 (N_11748,N_8708,N_7259);
and U11749 (N_11749,N_6580,N_7334);
or U11750 (N_11750,N_8735,N_7335);
or U11751 (N_11751,N_8907,N_7706);
xnor U11752 (N_11752,N_7046,N_8950);
and U11753 (N_11753,N_6495,N_6618);
nand U11754 (N_11754,N_6705,N_9057);
and U11755 (N_11755,N_8118,N_7134);
xnor U11756 (N_11756,N_9137,N_6367);
nand U11757 (N_11757,N_7270,N_8126);
and U11758 (N_11758,N_6828,N_7036);
or U11759 (N_11759,N_7234,N_8116);
nand U11760 (N_11760,N_8454,N_8864);
xor U11761 (N_11761,N_6510,N_9077);
and U11762 (N_11762,N_7156,N_7769);
xnor U11763 (N_11763,N_7571,N_6294);
xor U11764 (N_11764,N_6931,N_9361);
nand U11765 (N_11765,N_8759,N_6663);
xnor U11766 (N_11766,N_7604,N_7415);
nor U11767 (N_11767,N_9060,N_8045);
or U11768 (N_11768,N_7154,N_7568);
and U11769 (N_11769,N_6379,N_8299);
nand U11770 (N_11770,N_7976,N_7813);
nand U11771 (N_11771,N_7813,N_6885);
nor U11772 (N_11772,N_6979,N_8461);
or U11773 (N_11773,N_7349,N_7054);
nor U11774 (N_11774,N_9294,N_6915);
and U11775 (N_11775,N_9226,N_8239);
nor U11776 (N_11776,N_6423,N_7852);
and U11777 (N_11777,N_6263,N_7209);
or U11778 (N_11778,N_9269,N_7128);
nand U11779 (N_11779,N_8854,N_7265);
nor U11780 (N_11780,N_7694,N_8402);
nand U11781 (N_11781,N_7520,N_7450);
nand U11782 (N_11782,N_8605,N_7271);
and U11783 (N_11783,N_8303,N_7332);
nand U11784 (N_11784,N_8695,N_9060);
and U11785 (N_11785,N_9101,N_8314);
or U11786 (N_11786,N_6500,N_7308);
and U11787 (N_11787,N_9159,N_6870);
and U11788 (N_11788,N_7430,N_6921);
and U11789 (N_11789,N_7410,N_8370);
xor U11790 (N_11790,N_7154,N_6945);
nor U11791 (N_11791,N_7451,N_7338);
or U11792 (N_11792,N_7778,N_7126);
xor U11793 (N_11793,N_7921,N_6331);
nand U11794 (N_11794,N_9136,N_7391);
nand U11795 (N_11795,N_9129,N_6993);
xor U11796 (N_11796,N_7922,N_7434);
or U11797 (N_11797,N_8185,N_6714);
xor U11798 (N_11798,N_7991,N_6941);
and U11799 (N_11799,N_8967,N_7076);
or U11800 (N_11800,N_8057,N_7723);
nand U11801 (N_11801,N_6876,N_6295);
nor U11802 (N_11802,N_7865,N_7309);
nand U11803 (N_11803,N_7746,N_6925);
nor U11804 (N_11804,N_8845,N_6483);
and U11805 (N_11805,N_7269,N_8802);
or U11806 (N_11806,N_8773,N_7450);
nand U11807 (N_11807,N_7289,N_7972);
nand U11808 (N_11808,N_6403,N_6901);
or U11809 (N_11809,N_7021,N_9240);
nand U11810 (N_11810,N_8562,N_8492);
nand U11811 (N_11811,N_7307,N_6809);
and U11812 (N_11812,N_9108,N_7920);
nor U11813 (N_11813,N_7332,N_8799);
and U11814 (N_11814,N_8152,N_7856);
and U11815 (N_11815,N_7908,N_8170);
and U11816 (N_11816,N_6566,N_6504);
nor U11817 (N_11817,N_8773,N_9241);
and U11818 (N_11818,N_7788,N_7184);
nand U11819 (N_11819,N_8641,N_8444);
xor U11820 (N_11820,N_8829,N_8132);
or U11821 (N_11821,N_8434,N_7252);
nand U11822 (N_11822,N_7902,N_8629);
and U11823 (N_11823,N_8956,N_9071);
xor U11824 (N_11824,N_7096,N_8882);
xor U11825 (N_11825,N_6315,N_8698);
or U11826 (N_11826,N_7939,N_6865);
xor U11827 (N_11827,N_7651,N_6356);
and U11828 (N_11828,N_7633,N_9365);
nor U11829 (N_11829,N_8100,N_7552);
and U11830 (N_11830,N_9307,N_6803);
or U11831 (N_11831,N_7951,N_8616);
nand U11832 (N_11832,N_8505,N_6699);
nor U11833 (N_11833,N_7580,N_7895);
nor U11834 (N_11834,N_6489,N_8878);
and U11835 (N_11835,N_8085,N_8712);
nor U11836 (N_11836,N_8732,N_7790);
xor U11837 (N_11837,N_6433,N_8017);
or U11838 (N_11838,N_8529,N_7023);
nor U11839 (N_11839,N_7360,N_8225);
nand U11840 (N_11840,N_7173,N_7054);
and U11841 (N_11841,N_6636,N_7345);
nor U11842 (N_11842,N_8830,N_8528);
and U11843 (N_11843,N_7992,N_7154);
and U11844 (N_11844,N_8708,N_9216);
or U11845 (N_11845,N_8412,N_7857);
or U11846 (N_11846,N_8505,N_7766);
nand U11847 (N_11847,N_6465,N_6355);
xor U11848 (N_11848,N_7900,N_7871);
nor U11849 (N_11849,N_8489,N_8195);
or U11850 (N_11850,N_9112,N_7259);
or U11851 (N_11851,N_8351,N_9161);
and U11852 (N_11852,N_9240,N_7444);
or U11853 (N_11853,N_6385,N_8143);
and U11854 (N_11854,N_6793,N_8432);
xor U11855 (N_11855,N_7825,N_6623);
nand U11856 (N_11856,N_9252,N_7782);
nor U11857 (N_11857,N_7055,N_8087);
or U11858 (N_11858,N_7791,N_7961);
nor U11859 (N_11859,N_6569,N_6987);
xor U11860 (N_11860,N_7709,N_8223);
nand U11861 (N_11861,N_8280,N_7501);
nand U11862 (N_11862,N_6425,N_6410);
nor U11863 (N_11863,N_6536,N_8837);
xor U11864 (N_11864,N_8592,N_7250);
xor U11865 (N_11865,N_9309,N_8522);
or U11866 (N_11866,N_7495,N_7412);
nor U11867 (N_11867,N_9197,N_7700);
or U11868 (N_11868,N_8654,N_7104);
nor U11869 (N_11869,N_6339,N_8709);
and U11870 (N_11870,N_6747,N_6697);
xnor U11871 (N_11871,N_8842,N_7606);
nor U11872 (N_11872,N_7006,N_7691);
xor U11873 (N_11873,N_6523,N_8564);
or U11874 (N_11874,N_6942,N_8962);
xnor U11875 (N_11875,N_7421,N_6697);
or U11876 (N_11876,N_7329,N_7780);
xnor U11877 (N_11877,N_7698,N_6626);
xor U11878 (N_11878,N_8973,N_6874);
xnor U11879 (N_11879,N_6842,N_7760);
nand U11880 (N_11880,N_8290,N_6340);
or U11881 (N_11881,N_7509,N_6892);
or U11882 (N_11882,N_8244,N_7185);
and U11883 (N_11883,N_7528,N_8700);
xor U11884 (N_11884,N_8186,N_8652);
xor U11885 (N_11885,N_8203,N_7242);
nand U11886 (N_11886,N_8758,N_7807);
and U11887 (N_11887,N_7162,N_8522);
nor U11888 (N_11888,N_8120,N_8938);
and U11889 (N_11889,N_8065,N_6304);
nor U11890 (N_11890,N_7112,N_7844);
xnor U11891 (N_11891,N_6970,N_8730);
nor U11892 (N_11892,N_9249,N_9001);
nand U11893 (N_11893,N_8321,N_9069);
xnor U11894 (N_11894,N_6811,N_8551);
nor U11895 (N_11895,N_8919,N_6917);
xor U11896 (N_11896,N_7279,N_7166);
and U11897 (N_11897,N_8225,N_7508);
nand U11898 (N_11898,N_8993,N_7237);
and U11899 (N_11899,N_6532,N_8042);
or U11900 (N_11900,N_7596,N_8057);
or U11901 (N_11901,N_9114,N_6520);
or U11902 (N_11902,N_7905,N_8261);
nand U11903 (N_11903,N_8377,N_8717);
nand U11904 (N_11904,N_8662,N_8648);
or U11905 (N_11905,N_8325,N_7510);
xnor U11906 (N_11906,N_9090,N_6997);
nor U11907 (N_11907,N_6734,N_6924);
or U11908 (N_11908,N_7107,N_7052);
nand U11909 (N_11909,N_6357,N_7087);
nor U11910 (N_11910,N_8626,N_6618);
xnor U11911 (N_11911,N_6720,N_6405);
nand U11912 (N_11912,N_7679,N_8892);
nand U11913 (N_11913,N_7145,N_8039);
xnor U11914 (N_11914,N_6774,N_9101);
or U11915 (N_11915,N_7329,N_7530);
nor U11916 (N_11916,N_9122,N_8740);
or U11917 (N_11917,N_7075,N_7788);
nor U11918 (N_11918,N_7946,N_6862);
nor U11919 (N_11919,N_6604,N_8879);
nor U11920 (N_11920,N_6423,N_7387);
and U11921 (N_11921,N_6644,N_8295);
and U11922 (N_11922,N_9268,N_8448);
nor U11923 (N_11923,N_8670,N_8633);
and U11924 (N_11924,N_8699,N_7777);
nor U11925 (N_11925,N_6934,N_7466);
or U11926 (N_11926,N_7884,N_6569);
nor U11927 (N_11927,N_8262,N_7634);
nand U11928 (N_11928,N_8384,N_8709);
and U11929 (N_11929,N_6927,N_7783);
and U11930 (N_11930,N_8031,N_8055);
xor U11931 (N_11931,N_7279,N_6838);
xnor U11932 (N_11932,N_8729,N_6978);
nand U11933 (N_11933,N_7954,N_8869);
nand U11934 (N_11934,N_7106,N_7249);
nor U11935 (N_11935,N_7495,N_7241);
xnor U11936 (N_11936,N_9170,N_6523);
xnor U11937 (N_11937,N_7623,N_7071);
xor U11938 (N_11938,N_6627,N_9251);
or U11939 (N_11939,N_6267,N_8051);
nor U11940 (N_11940,N_8787,N_8213);
nand U11941 (N_11941,N_7451,N_9246);
nand U11942 (N_11942,N_7936,N_7081);
or U11943 (N_11943,N_9180,N_8809);
nand U11944 (N_11944,N_6975,N_8767);
or U11945 (N_11945,N_9174,N_9281);
nor U11946 (N_11946,N_8956,N_6337);
nand U11947 (N_11947,N_9040,N_7348);
nor U11948 (N_11948,N_7109,N_8756);
xor U11949 (N_11949,N_7030,N_7636);
and U11950 (N_11950,N_8782,N_8785);
nand U11951 (N_11951,N_7981,N_8863);
xnor U11952 (N_11952,N_7087,N_8448);
nand U11953 (N_11953,N_7622,N_7603);
or U11954 (N_11954,N_9330,N_8373);
xnor U11955 (N_11955,N_6718,N_6466);
xor U11956 (N_11956,N_9198,N_6793);
xor U11957 (N_11957,N_6468,N_6475);
and U11958 (N_11958,N_8151,N_7120);
or U11959 (N_11959,N_7900,N_7768);
or U11960 (N_11960,N_8364,N_8955);
nand U11961 (N_11961,N_6791,N_7653);
or U11962 (N_11962,N_7613,N_8687);
xnor U11963 (N_11963,N_6960,N_8607);
xor U11964 (N_11964,N_9276,N_7300);
and U11965 (N_11965,N_6988,N_8409);
xor U11966 (N_11966,N_6833,N_8328);
or U11967 (N_11967,N_8930,N_9183);
xor U11968 (N_11968,N_7982,N_8431);
or U11969 (N_11969,N_7984,N_7676);
and U11970 (N_11970,N_8879,N_8668);
xor U11971 (N_11971,N_8971,N_7277);
and U11972 (N_11972,N_6861,N_6620);
xor U11973 (N_11973,N_7945,N_8884);
xor U11974 (N_11974,N_6551,N_8461);
and U11975 (N_11975,N_8843,N_7518);
and U11976 (N_11976,N_8386,N_7081);
nor U11977 (N_11977,N_7009,N_9004);
nand U11978 (N_11978,N_6262,N_8183);
or U11979 (N_11979,N_6911,N_8833);
or U11980 (N_11980,N_7272,N_7184);
or U11981 (N_11981,N_6456,N_9053);
and U11982 (N_11982,N_6747,N_8313);
xnor U11983 (N_11983,N_6996,N_9032);
nor U11984 (N_11984,N_7764,N_8806);
and U11985 (N_11985,N_8324,N_6852);
xnor U11986 (N_11986,N_7873,N_6311);
nand U11987 (N_11987,N_8784,N_8993);
nor U11988 (N_11988,N_9078,N_7145);
xor U11989 (N_11989,N_8490,N_6603);
xor U11990 (N_11990,N_7023,N_7865);
nand U11991 (N_11991,N_8052,N_7148);
nor U11992 (N_11992,N_8350,N_7832);
and U11993 (N_11993,N_9219,N_8732);
nor U11994 (N_11994,N_6442,N_6856);
and U11995 (N_11995,N_7322,N_7145);
nor U11996 (N_11996,N_6274,N_9114);
nand U11997 (N_11997,N_8870,N_9028);
or U11998 (N_11998,N_7826,N_9243);
and U11999 (N_11999,N_7570,N_9348);
and U12000 (N_12000,N_8811,N_9041);
nor U12001 (N_12001,N_6451,N_8206);
xor U12002 (N_12002,N_6368,N_8793);
or U12003 (N_12003,N_7011,N_7631);
or U12004 (N_12004,N_6287,N_8423);
nor U12005 (N_12005,N_7704,N_6684);
xnor U12006 (N_12006,N_8089,N_8316);
or U12007 (N_12007,N_7889,N_7311);
and U12008 (N_12008,N_9001,N_8369);
and U12009 (N_12009,N_8875,N_6750);
xnor U12010 (N_12010,N_9151,N_7136);
xnor U12011 (N_12011,N_6283,N_7789);
xor U12012 (N_12012,N_7079,N_7036);
nand U12013 (N_12013,N_8889,N_7086);
or U12014 (N_12014,N_8837,N_7221);
nor U12015 (N_12015,N_8014,N_8028);
and U12016 (N_12016,N_7179,N_8760);
nand U12017 (N_12017,N_7191,N_8226);
and U12018 (N_12018,N_8284,N_6560);
nor U12019 (N_12019,N_6709,N_8875);
or U12020 (N_12020,N_6972,N_7011);
or U12021 (N_12021,N_8337,N_6573);
and U12022 (N_12022,N_8596,N_6297);
nand U12023 (N_12023,N_6964,N_6658);
xor U12024 (N_12024,N_6413,N_9004);
xor U12025 (N_12025,N_7358,N_7763);
or U12026 (N_12026,N_8739,N_8098);
or U12027 (N_12027,N_9348,N_6838);
nor U12028 (N_12028,N_9216,N_9128);
or U12029 (N_12029,N_7201,N_6291);
nor U12030 (N_12030,N_6874,N_8767);
and U12031 (N_12031,N_6650,N_8596);
xor U12032 (N_12032,N_7653,N_6827);
nand U12033 (N_12033,N_9044,N_7749);
nand U12034 (N_12034,N_8688,N_7424);
xor U12035 (N_12035,N_6803,N_7553);
or U12036 (N_12036,N_8555,N_6944);
and U12037 (N_12037,N_7732,N_8244);
xnor U12038 (N_12038,N_8923,N_8605);
or U12039 (N_12039,N_6711,N_6261);
or U12040 (N_12040,N_9296,N_8452);
or U12041 (N_12041,N_8344,N_8206);
nor U12042 (N_12042,N_7077,N_8669);
xnor U12043 (N_12043,N_8367,N_8523);
nand U12044 (N_12044,N_8030,N_8902);
nor U12045 (N_12045,N_7070,N_8467);
and U12046 (N_12046,N_6921,N_8136);
and U12047 (N_12047,N_8623,N_8422);
xor U12048 (N_12048,N_9092,N_8123);
nand U12049 (N_12049,N_7980,N_6442);
nor U12050 (N_12050,N_8963,N_8489);
xor U12051 (N_12051,N_7401,N_8040);
or U12052 (N_12052,N_7491,N_6424);
or U12053 (N_12053,N_6351,N_6490);
nor U12054 (N_12054,N_7441,N_7833);
xnor U12055 (N_12055,N_9076,N_6868);
nand U12056 (N_12056,N_7790,N_8450);
or U12057 (N_12057,N_8774,N_8734);
xnor U12058 (N_12058,N_6663,N_7595);
and U12059 (N_12059,N_7202,N_7228);
or U12060 (N_12060,N_6842,N_8009);
or U12061 (N_12061,N_7489,N_8509);
xnor U12062 (N_12062,N_8779,N_7077);
nand U12063 (N_12063,N_8093,N_6325);
nand U12064 (N_12064,N_6528,N_7613);
nand U12065 (N_12065,N_7801,N_7145);
or U12066 (N_12066,N_8697,N_7307);
nand U12067 (N_12067,N_9356,N_9098);
nor U12068 (N_12068,N_7139,N_8195);
or U12069 (N_12069,N_6257,N_6762);
or U12070 (N_12070,N_9078,N_8075);
nand U12071 (N_12071,N_8644,N_8693);
xnor U12072 (N_12072,N_7583,N_6936);
and U12073 (N_12073,N_9277,N_8094);
and U12074 (N_12074,N_7860,N_8011);
xnor U12075 (N_12075,N_9180,N_8196);
nor U12076 (N_12076,N_6809,N_6308);
xor U12077 (N_12077,N_8605,N_8162);
and U12078 (N_12078,N_7617,N_7828);
or U12079 (N_12079,N_8565,N_8732);
nand U12080 (N_12080,N_8417,N_6722);
xnor U12081 (N_12081,N_8294,N_9052);
and U12082 (N_12082,N_8661,N_6461);
or U12083 (N_12083,N_7143,N_7318);
and U12084 (N_12084,N_6488,N_8272);
and U12085 (N_12085,N_6510,N_8847);
xnor U12086 (N_12086,N_7856,N_9086);
nand U12087 (N_12087,N_7182,N_6956);
or U12088 (N_12088,N_7347,N_7746);
nor U12089 (N_12089,N_7330,N_6537);
xor U12090 (N_12090,N_6580,N_6433);
or U12091 (N_12091,N_6477,N_8892);
xnor U12092 (N_12092,N_9133,N_6296);
or U12093 (N_12093,N_6901,N_9024);
nor U12094 (N_12094,N_9202,N_9155);
nand U12095 (N_12095,N_6578,N_6952);
nor U12096 (N_12096,N_6639,N_7871);
and U12097 (N_12097,N_7116,N_8458);
xnor U12098 (N_12098,N_8641,N_7936);
or U12099 (N_12099,N_6366,N_6513);
and U12100 (N_12100,N_7433,N_6693);
nand U12101 (N_12101,N_6831,N_7206);
xnor U12102 (N_12102,N_8692,N_8566);
nor U12103 (N_12103,N_9017,N_8254);
or U12104 (N_12104,N_8511,N_6956);
and U12105 (N_12105,N_6749,N_6855);
or U12106 (N_12106,N_6884,N_8539);
or U12107 (N_12107,N_6378,N_6465);
xnor U12108 (N_12108,N_8457,N_7501);
nand U12109 (N_12109,N_6954,N_8723);
and U12110 (N_12110,N_6510,N_6729);
nand U12111 (N_12111,N_9364,N_7410);
or U12112 (N_12112,N_8529,N_7952);
nor U12113 (N_12113,N_7522,N_6282);
xnor U12114 (N_12114,N_6682,N_8146);
nand U12115 (N_12115,N_8218,N_9117);
nor U12116 (N_12116,N_8870,N_9212);
xor U12117 (N_12117,N_7919,N_6852);
nand U12118 (N_12118,N_9015,N_9036);
and U12119 (N_12119,N_6693,N_9246);
xnor U12120 (N_12120,N_6555,N_6893);
nor U12121 (N_12121,N_8820,N_7282);
xor U12122 (N_12122,N_8093,N_7180);
xor U12123 (N_12123,N_6914,N_8437);
xor U12124 (N_12124,N_6802,N_6361);
nand U12125 (N_12125,N_9194,N_6301);
and U12126 (N_12126,N_8078,N_9114);
and U12127 (N_12127,N_8098,N_6912);
xnor U12128 (N_12128,N_6854,N_7165);
xnor U12129 (N_12129,N_9008,N_6700);
xor U12130 (N_12130,N_9185,N_7822);
nand U12131 (N_12131,N_7092,N_7320);
nand U12132 (N_12132,N_8443,N_8433);
or U12133 (N_12133,N_6391,N_7832);
or U12134 (N_12134,N_7336,N_8357);
nor U12135 (N_12135,N_8903,N_8256);
nand U12136 (N_12136,N_9292,N_8113);
xnor U12137 (N_12137,N_6890,N_8905);
nor U12138 (N_12138,N_9054,N_7813);
and U12139 (N_12139,N_7398,N_7434);
xor U12140 (N_12140,N_9226,N_6981);
xnor U12141 (N_12141,N_7398,N_9284);
and U12142 (N_12142,N_9166,N_8912);
xor U12143 (N_12143,N_9237,N_8693);
xor U12144 (N_12144,N_9317,N_7921);
nor U12145 (N_12145,N_8618,N_8948);
or U12146 (N_12146,N_8573,N_7829);
nand U12147 (N_12147,N_7440,N_6343);
xor U12148 (N_12148,N_6849,N_7464);
xor U12149 (N_12149,N_6452,N_6326);
nor U12150 (N_12150,N_8908,N_8754);
nand U12151 (N_12151,N_7100,N_8520);
or U12152 (N_12152,N_9097,N_8912);
nor U12153 (N_12153,N_9270,N_7368);
nor U12154 (N_12154,N_9301,N_7606);
and U12155 (N_12155,N_7596,N_8663);
nor U12156 (N_12156,N_9089,N_7539);
nand U12157 (N_12157,N_8922,N_8477);
nand U12158 (N_12158,N_8236,N_6950);
or U12159 (N_12159,N_6329,N_7665);
xnor U12160 (N_12160,N_8271,N_7130);
and U12161 (N_12161,N_8246,N_8720);
and U12162 (N_12162,N_7706,N_7662);
xnor U12163 (N_12163,N_9283,N_7833);
xnor U12164 (N_12164,N_6463,N_6626);
and U12165 (N_12165,N_9062,N_7346);
or U12166 (N_12166,N_8686,N_8121);
nor U12167 (N_12167,N_9150,N_8122);
nor U12168 (N_12168,N_9026,N_7149);
and U12169 (N_12169,N_8222,N_6315);
nand U12170 (N_12170,N_7976,N_6343);
xnor U12171 (N_12171,N_8764,N_9351);
xor U12172 (N_12172,N_8315,N_6912);
nor U12173 (N_12173,N_7761,N_8891);
or U12174 (N_12174,N_7446,N_8707);
nor U12175 (N_12175,N_7972,N_8443);
or U12176 (N_12176,N_9145,N_6837);
or U12177 (N_12177,N_7984,N_8435);
nor U12178 (N_12178,N_7009,N_6862);
nand U12179 (N_12179,N_6951,N_9285);
nor U12180 (N_12180,N_7325,N_6301);
and U12181 (N_12181,N_7428,N_7434);
and U12182 (N_12182,N_8288,N_7203);
nand U12183 (N_12183,N_6596,N_6531);
and U12184 (N_12184,N_7750,N_9225);
and U12185 (N_12185,N_8198,N_7559);
nor U12186 (N_12186,N_7083,N_6419);
and U12187 (N_12187,N_6442,N_8483);
or U12188 (N_12188,N_8038,N_7933);
and U12189 (N_12189,N_7402,N_7004);
or U12190 (N_12190,N_8535,N_8248);
xor U12191 (N_12191,N_7651,N_6545);
and U12192 (N_12192,N_7118,N_6714);
nand U12193 (N_12193,N_8682,N_6490);
and U12194 (N_12194,N_7297,N_6838);
nand U12195 (N_12195,N_8639,N_6629);
xnor U12196 (N_12196,N_7052,N_6524);
or U12197 (N_12197,N_9087,N_6432);
and U12198 (N_12198,N_6658,N_6522);
nand U12199 (N_12199,N_6820,N_8168);
nor U12200 (N_12200,N_9197,N_8332);
xor U12201 (N_12201,N_8565,N_6755);
or U12202 (N_12202,N_6923,N_7661);
xor U12203 (N_12203,N_8218,N_7502);
nor U12204 (N_12204,N_6314,N_6349);
xor U12205 (N_12205,N_6733,N_7011);
and U12206 (N_12206,N_8599,N_8207);
or U12207 (N_12207,N_7557,N_8229);
and U12208 (N_12208,N_6671,N_6654);
xnor U12209 (N_12209,N_7844,N_8787);
nand U12210 (N_12210,N_7414,N_7427);
xor U12211 (N_12211,N_9131,N_6461);
xnor U12212 (N_12212,N_8562,N_7414);
nand U12213 (N_12213,N_7753,N_9141);
nor U12214 (N_12214,N_8422,N_7810);
nor U12215 (N_12215,N_7119,N_7164);
xor U12216 (N_12216,N_7554,N_7267);
xnor U12217 (N_12217,N_8014,N_7142);
nor U12218 (N_12218,N_8658,N_8897);
xnor U12219 (N_12219,N_9105,N_7815);
and U12220 (N_12220,N_7990,N_6384);
nand U12221 (N_12221,N_6563,N_6468);
or U12222 (N_12222,N_7969,N_8875);
nor U12223 (N_12223,N_8179,N_7298);
xnor U12224 (N_12224,N_7805,N_8934);
nand U12225 (N_12225,N_8820,N_8216);
xnor U12226 (N_12226,N_6505,N_8441);
nand U12227 (N_12227,N_7060,N_8687);
and U12228 (N_12228,N_7966,N_9263);
or U12229 (N_12229,N_6355,N_8427);
nor U12230 (N_12230,N_8327,N_7844);
or U12231 (N_12231,N_6669,N_7211);
nand U12232 (N_12232,N_7953,N_8183);
nand U12233 (N_12233,N_9065,N_7808);
nor U12234 (N_12234,N_7119,N_6984);
nand U12235 (N_12235,N_8449,N_7145);
nor U12236 (N_12236,N_6733,N_6668);
xor U12237 (N_12237,N_9092,N_9211);
xor U12238 (N_12238,N_7376,N_8978);
nor U12239 (N_12239,N_9261,N_8152);
and U12240 (N_12240,N_6859,N_7446);
xor U12241 (N_12241,N_8172,N_8658);
nand U12242 (N_12242,N_6447,N_6465);
and U12243 (N_12243,N_8487,N_8057);
and U12244 (N_12244,N_6931,N_8297);
or U12245 (N_12245,N_8522,N_9312);
nand U12246 (N_12246,N_7604,N_7812);
and U12247 (N_12247,N_8470,N_6319);
nand U12248 (N_12248,N_7382,N_8037);
or U12249 (N_12249,N_7961,N_8136);
and U12250 (N_12250,N_6644,N_6789);
nor U12251 (N_12251,N_6257,N_8718);
nand U12252 (N_12252,N_9020,N_6664);
xor U12253 (N_12253,N_6553,N_7212);
and U12254 (N_12254,N_7765,N_9193);
xnor U12255 (N_12255,N_8363,N_7383);
xnor U12256 (N_12256,N_7373,N_8236);
nand U12257 (N_12257,N_6334,N_8942);
nand U12258 (N_12258,N_8746,N_7078);
or U12259 (N_12259,N_9119,N_6649);
nor U12260 (N_12260,N_6431,N_8801);
or U12261 (N_12261,N_6480,N_6344);
and U12262 (N_12262,N_8574,N_7193);
nor U12263 (N_12263,N_6525,N_8447);
nor U12264 (N_12264,N_8956,N_6929);
or U12265 (N_12265,N_7268,N_7233);
xor U12266 (N_12266,N_6741,N_9253);
and U12267 (N_12267,N_7257,N_8229);
nand U12268 (N_12268,N_6947,N_8098);
or U12269 (N_12269,N_8833,N_7784);
and U12270 (N_12270,N_6454,N_8409);
or U12271 (N_12271,N_7991,N_7077);
nor U12272 (N_12272,N_7595,N_8869);
and U12273 (N_12273,N_8060,N_8218);
nor U12274 (N_12274,N_8925,N_8992);
nor U12275 (N_12275,N_7766,N_8724);
and U12276 (N_12276,N_7046,N_6521);
and U12277 (N_12277,N_6962,N_6720);
nor U12278 (N_12278,N_7243,N_9165);
xnor U12279 (N_12279,N_7765,N_8954);
and U12280 (N_12280,N_9075,N_8509);
xor U12281 (N_12281,N_7303,N_7022);
nor U12282 (N_12282,N_7920,N_6732);
and U12283 (N_12283,N_6483,N_7470);
nor U12284 (N_12284,N_7419,N_9022);
nand U12285 (N_12285,N_9051,N_6872);
or U12286 (N_12286,N_8765,N_7926);
and U12287 (N_12287,N_6488,N_7255);
and U12288 (N_12288,N_6471,N_7455);
nor U12289 (N_12289,N_6778,N_8181);
xor U12290 (N_12290,N_7115,N_7960);
nand U12291 (N_12291,N_7333,N_6788);
and U12292 (N_12292,N_6281,N_7190);
nand U12293 (N_12293,N_6754,N_7491);
nand U12294 (N_12294,N_9181,N_7717);
xnor U12295 (N_12295,N_8762,N_8095);
nand U12296 (N_12296,N_9041,N_8748);
and U12297 (N_12297,N_8389,N_9160);
or U12298 (N_12298,N_7539,N_6815);
and U12299 (N_12299,N_6975,N_8617);
nand U12300 (N_12300,N_9246,N_8926);
nand U12301 (N_12301,N_6768,N_8981);
or U12302 (N_12302,N_6907,N_8060);
nand U12303 (N_12303,N_7990,N_8284);
nand U12304 (N_12304,N_8130,N_7414);
or U12305 (N_12305,N_6416,N_6332);
and U12306 (N_12306,N_8572,N_8762);
or U12307 (N_12307,N_6450,N_7223);
nand U12308 (N_12308,N_9260,N_6569);
nand U12309 (N_12309,N_8982,N_8357);
nand U12310 (N_12310,N_8197,N_7953);
nor U12311 (N_12311,N_6709,N_6423);
or U12312 (N_12312,N_8389,N_8366);
xor U12313 (N_12313,N_7639,N_8637);
and U12314 (N_12314,N_8361,N_6357);
and U12315 (N_12315,N_7858,N_9024);
and U12316 (N_12316,N_9020,N_8194);
nand U12317 (N_12317,N_9044,N_7012);
xnor U12318 (N_12318,N_7968,N_7260);
and U12319 (N_12319,N_8092,N_9116);
nand U12320 (N_12320,N_8553,N_7758);
nand U12321 (N_12321,N_9355,N_8269);
nand U12322 (N_12322,N_9177,N_8150);
xnor U12323 (N_12323,N_7936,N_8777);
xnor U12324 (N_12324,N_7014,N_6859);
nand U12325 (N_12325,N_7950,N_7471);
nand U12326 (N_12326,N_6824,N_9235);
or U12327 (N_12327,N_9336,N_6786);
nor U12328 (N_12328,N_7964,N_8729);
nor U12329 (N_12329,N_8960,N_8352);
or U12330 (N_12330,N_8216,N_6962);
xnor U12331 (N_12331,N_8548,N_8514);
nand U12332 (N_12332,N_7238,N_6625);
xor U12333 (N_12333,N_8245,N_8430);
xnor U12334 (N_12334,N_7584,N_7243);
and U12335 (N_12335,N_8175,N_6888);
nand U12336 (N_12336,N_8435,N_6860);
and U12337 (N_12337,N_9321,N_6907);
nor U12338 (N_12338,N_7649,N_9178);
and U12339 (N_12339,N_6832,N_6648);
or U12340 (N_12340,N_7245,N_7110);
xnor U12341 (N_12341,N_8968,N_8882);
nand U12342 (N_12342,N_7048,N_7733);
nor U12343 (N_12343,N_9245,N_8849);
nor U12344 (N_12344,N_8559,N_9088);
and U12345 (N_12345,N_7840,N_7018);
nand U12346 (N_12346,N_6926,N_7232);
and U12347 (N_12347,N_7530,N_8771);
xor U12348 (N_12348,N_8166,N_6306);
nor U12349 (N_12349,N_8937,N_7434);
xnor U12350 (N_12350,N_7149,N_7276);
nor U12351 (N_12351,N_9207,N_8737);
nor U12352 (N_12352,N_9249,N_6696);
and U12353 (N_12353,N_9013,N_7697);
nor U12354 (N_12354,N_6745,N_8463);
and U12355 (N_12355,N_7770,N_7868);
or U12356 (N_12356,N_9136,N_9227);
xnor U12357 (N_12357,N_7834,N_6673);
or U12358 (N_12358,N_8314,N_7442);
xor U12359 (N_12359,N_7493,N_8010);
nor U12360 (N_12360,N_8186,N_8004);
or U12361 (N_12361,N_8844,N_8988);
and U12362 (N_12362,N_6915,N_8921);
or U12363 (N_12363,N_8536,N_6741);
nand U12364 (N_12364,N_6627,N_6531);
nand U12365 (N_12365,N_8586,N_8602);
nand U12366 (N_12366,N_6531,N_7266);
or U12367 (N_12367,N_9337,N_8756);
xnor U12368 (N_12368,N_7757,N_8064);
nor U12369 (N_12369,N_7731,N_6709);
nor U12370 (N_12370,N_6658,N_7254);
xnor U12371 (N_12371,N_6923,N_8370);
nand U12372 (N_12372,N_9146,N_9268);
nor U12373 (N_12373,N_6603,N_8243);
nor U12374 (N_12374,N_7598,N_7485);
xor U12375 (N_12375,N_8949,N_6348);
nor U12376 (N_12376,N_7054,N_9231);
xor U12377 (N_12377,N_7661,N_8262);
xor U12378 (N_12378,N_8034,N_9003);
or U12379 (N_12379,N_8136,N_6329);
nand U12380 (N_12380,N_8862,N_6289);
nand U12381 (N_12381,N_9058,N_7395);
xor U12382 (N_12382,N_7152,N_7397);
and U12383 (N_12383,N_7612,N_8731);
nor U12384 (N_12384,N_9239,N_7665);
and U12385 (N_12385,N_7915,N_8441);
xor U12386 (N_12386,N_7799,N_6706);
nand U12387 (N_12387,N_8261,N_6549);
nand U12388 (N_12388,N_8782,N_9319);
nor U12389 (N_12389,N_8515,N_8640);
nor U12390 (N_12390,N_7254,N_7530);
xor U12391 (N_12391,N_8572,N_8793);
nor U12392 (N_12392,N_7962,N_6412);
nand U12393 (N_12393,N_9087,N_7536);
xnor U12394 (N_12394,N_7637,N_6577);
or U12395 (N_12395,N_6370,N_8030);
xor U12396 (N_12396,N_6337,N_6860);
or U12397 (N_12397,N_6385,N_6884);
and U12398 (N_12398,N_7711,N_7272);
nand U12399 (N_12399,N_7741,N_8892);
nor U12400 (N_12400,N_7953,N_6876);
nand U12401 (N_12401,N_7975,N_7924);
or U12402 (N_12402,N_8567,N_8130);
nand U12403 (N_12403,N_8804,N_8642);
or U12404 (N_12404,N_7943,N_7293);
nor U12405 (N_12405,N_6260,N_6954);
xnor U12406 (N_12406,N_8979,N_6456);
and U12407 (N_12407,N_7718,N_9241);
nor U12408 (N_12408,N_8016,N_8256);
nor U12409 (N_12409,N_8233,N_7465);
xnor U12410 (N_12410,N_6675,N_6281);
nor U12411 (N_12411,N_9103,N_6685);
nor U12412 (N_12412,N_6438,N_8374);
nand U12413 (N_12413,N_6830,N_7236);
and U12414 (N_12414,N_6550,N_6359);
and U12415 (N_12415,N_7152,N_9112);
or U12416 (N_12416,N_6271,N_7804);
nand U12417 (N_12417,N_9065,N_8729);
nand U12418 (N_12418,N_7855,N_8574);
and U12419 (N_12419,N_7901,N_6532);
and U12420 (N_12420,N_6547,N_7979);
or U12421 (N_12421,N_7273,N_8065);
nor U12422 (N_12422,N_9361,N_7367);
and U12423 (N_12423,N_9371,N_6329);
nand U12424 (N_12424,N_9113,N_8409);
xnor U12425 (N_12425,N_6711,N_7460);
nor U12426 (N_12426,N_6901,N_9027);
nor U12427 (N_12427,N_7189,N_7945);
nand U12428 (N_12428,N_6694,N_8352);
nor U12429 (N_12429,N_9181,N_9293);
or U12430 (N_12430,N_8087,N_7384);
or U12431 (N_12431,N_7332,N_7403);
nand U12432 (N_12432,N_7885,N_6373);
and U12433 (N_12433,N_7430,N_8698);
and U12434 (N_12434,N_7471,N_6862);
and U12435 (N_12435,N_9134,N_7075);
nor U12436 (N_12436,N_8012,N_7361);
xor U12437 (N_12437,N_6643,N_7694);
xnor U12438 (N_12438,N_7469,N_8665);
nor U12439 (N_12439,N_6553,N_8593);
or U12440 (N_12440,N_8827,N_7754);
and U12441 (N_12441,N_8372,N_6637);
nand U12442 (N_12442,N_7712,N_8407);
nand U12443 (N_12443,N_6723,N_7868);
xnor U12444 (N_12444,N_6469,N_6639);
or U12445 (N_12445,N_8083,N_9037);
xnor U12446 (N_12446,N_8171,N_7974);
nand U12447 (N_12447,N_8850,N_8881);
or U12448 (N_12448,N_6636,N_9080);
or U12449 (N_12449,N_7696,N_6761);
or U12450 (N_12450,N_6895,N_7868);
xor U12451 (N_12451,N_7297,N_8772);
nand U12452 (N_12452,N_9343,N_9216);
or U12453 (N_12453,N_9088,N_6852);
nand U12454 (N_12454,N_8321,N_8050);
and U12455 (N_12455,N_8836,N_9072);
nand U12456 (N_12456,N_7761,N_6513);
xnor U12457 (N_12457,N_9280,N_8814);
or U12458 (N_12458,N_7905,N_9143);
and U12459 (N_12459,N_6640,N_7207);
or U12460 (N_12460,N_7736,N_8522);
nand U12461 (N_12461,N_9215,N_7922);
xor U12462 (N_12462,N_8570,N_9169);
nor U12463 (N_12463,N_7337,N_6363);
nor U12464 (N_12464,N_8829,N_8768);
or U12465 (N_12465,N_8069,N_6697);
nand U12466 (N_12466,N_8063,N_7816);
xor U12467 (N_12467,N_7823,N_8836);
nor U12468 (N_12468,N_8493,N_8945);
xor U12469 (N_12469,N_7789,N_7679);
nor U12470 (N_12470,N_8803,N_6903);
nor U12471 (N_12471,N_6476,N_8184);
nor U12472 (N_12472,N_8236,N_8830);
nor U12473 (N_12473,N_6985,N_8335);
or U12474 (N_12474,N_8543,N_6458);
xor U12475 (N_12475,N_7900,N_9275);
xor U12476 (N_12476,N_8658,N_6943);
nor U12477 (N_12477,N_9355,N_8103);
nor U12478 (N_12478,N_9198,N_6282);
nand U12479 (N_12479,N_7955,N_7616);
or U12480 (N_12480,N_7196,N_8668);
and U12481 (N_12481,N_6601,N_7912);
nor U12482 (N_12482,N_9036,N_7470);
nand U12483 (N_12483,N_9214,N_8085);
and U12484 (N_12484,N_7790,N_6328);
or U12485 (N_12485,N_6761,N_6615);
xor U12486 (N_12486,N_8731,N_9331);
nor U12487 (N_12487,N_6425,N_7888);
nand U12488 (N_12488,N_6428,N_6654);
nand U12489 (N_12489,N_8721,N_8700);
and U12490 (N_12490,N_7679,N_8418);
or U12491 (N_12491,N_7544,N_7818);
nor U12492 (N_12492,N_7850,N_6803);
nor U12493 (N_12493,N_7295,N_6355);
or U12494 (N_12494,N_9148,N_6323);
xnor U12495 (N_12495,N_7314,N_6864);
nor U12496 (N_12496,N_7781,N_7503);
nor U12497 (N_12497,N_9031,N_7737);
nand U12498 (N_12498,N_6768,N_7817);
nand U12499 (N_12499,N_7871,N_7238);
nor U12500 (N_12500,N_11629,N_11367);
nor U12501 (N_12501,N_12132,N_9604);
or U12502 (N_12502,N_10908,N_10256);
or U12503 (N_12503,N_10891,N_10332);
xor U12504 (N_12504,N_12483,N_10921);
and U12505 (N_12505,N_11091,N_11806);
nor U12506 (N_12506,N_10063,N_12148);
or U12507 (N_12507,N_12313,N_10077);
nor U12508 (N_12508,N_10638,N_10854);
nor U12509 (N_12509,N_12238,N_9881);
nor U12510 (N_12510,N_10468,N_11914);
xor U12511 (N_12511,N_9468,N_9544);
nand U12512 (N_12512,N_9754,N_10033);
nor U12513 (N_12513,N_11606,N_11744);
nand U12514 (N_12514,N_9847,N_11167);
xnor U12515 (N_12515,N_10973,N_10103);
and U12516 (N_12516,N_9417,N_11920);
nand U12517 (N_12517,N_10678,N_11880);
xor U12518 (N_12518,N_11359,N_12149);
nand U12519 (N_12519,N_10090,N_12112);
and U12520 (N_12520,N_10858,N_11430);
nor U12521 (N_12521,N_10054,N_10494);
and U12522 (N_12522,N_9711,N_12154);
nor U12523 (N_12523,N_12284,N_12374);
nand U12524 (N_12524,N_10152,N_12330);
or U12525 (N_12525,N_10706,N_12038);
xor U12526 (N_12526,N_11390,N_10842);
nand U12527 (N_12527,N_10965,N_9966);
or U12528 (N_12528,N_10221,N_12256);
or U12529 (N_12529,N_10113,N_10338);
and U12530 (N_12530,N_9786,N_10093);
and U12531 (N_12531,N_11712,N_10329);
nor U12532 (N_12532,N_9992,N_9545);
or U12533 (N_12533,N_12053,N_11174);
and U12534 (N_12534,N_10775,N_12480);
xor U12535 (N_12535,N_10347,N_9902);
nand U12536 (N_12536,N_12066,N_9515);
nand U12537 (N_12537,N_9645,N_11849);
nor U12538 (N_12538,N_11533,N_10450);
or U12539 (N_12539,N_11959,N_9858);
or U12540 (N_12540,N_11345,N_11297);
nor U12541 (N_12541,N_11679,N_10506);
xnor U12542 (N_12542,N_12447,N_10198);
and U12543 (N_12543,N_11395,N_11871);
nand U12544 (N_12544,N_10281,N_9542);
or U12545 (N_12545,N_11609,N_12479);
xnor U12546 (N_12546,N_11069,N_11076);
xor U12547 (N_12547,N_10607,N_10396);
nor U12548 (N_12548,N_11696,N_11272);
nor U12549 (N_12549,N_12065,N_11011);
or U12550 (N_12550,N_10668,N_11984);
nor U12551 (N_12551,N_10110,N_10645);
xnor U12552 (N_12552,N_10625,N_11885);
xnor U12553 (N_12553,N_10618,N_10685);
xor U12554 (N_12554,N_11136,N_12080);
or U12555 (N_12555,N_9827,N_11465);
nor U12556 (N_12556,N_12410,N_11888);
and U12557 (N_12557,N_12225,N_12365);
nand U12558 (N_12558,N_10791,N_9698);
nor U12559 (N_12559,N_10736,N_11342);
nor U12560 (N_12560,N_10774,N_12120);
nand U12561 (N_12561,N_12122,N_12451);
nor U12562 (N_12562,N_9581,N_11455);
nand U12563 (N_12563,N_10749,N_11128);
and U12564 (N_12564,N_9565,N_11713);
or U12565 (N_12565,N_10314,N_11701);
nand U12566 (N_12566,N_9998,N_9427);
or U12567 (N_12567,N_11692,N_12147);
nand U12568 (N_12568,N_11540,N_12312);
xor U12569 (N_12569,N_12308,N_11596);
xor U12570 (N_12570,N_9891,N_11036);
nor U12571 (N_12571,N_11265,N_9602);
or U12572 (N_12572,N_11886,N_12474);
or U12573 (N_12573,N_10700,N_9843);
or U12574 (N_12574,N_10265,N_9957);
and U12575 (N_12575,N_11073,N_10885);
nand U12576 (N_12576,N_11799,N_11057);
nor U12577 (N_12577,N_12357,N_12119);
nor U12578 (N_12578,N_12071,N_9480);
nand U12579 (N_12579,N_9636,N_11633);
nor U12580 (N_12580,N_10980,N_11018);
nand U12581 (N_12581,N_11224,N_11550);
xnor U12582 (N_12582,N_11163,N_11574);
xor U12583 (N_12583,N_9696,N_9913);
xnor U12584 (N_12584,N_11809,N_12243);
nor U12585 (N_12585,N_10301,N_12487);
or U12586 (N_12586,N_10853,N_12187);
and U12587 (N_12587,N_9936,N_10401);
nand U12588 (N_12588,N_12145,N_11241);
nor U12589 (N_12589,N_12353,N_10298);
or U12590 (N_12590,N_11226,N_10280);
nand U12591 (N_12591,N_12437,N_12342);
nand U12592 (N_12592,N_9747,N_9755);
nand U12593 (N_12593,N_10500,N_11741);
and U12594 (N_12594,N_11068,N_9407);
nand U12595 (N_12595,N_10560,N_12459);
xor U12596 (N_12596,N_11437,N_10955);
xnor U12597 (N_12597,N_9730,N_10830);
xor U12598 (N_12598,N_11321,N_10336);
or U12599 (N_12599,N_12272,N_10691);
xnor U12600 (N_12600,N_11129,N_9970);
nor U12601 (N_12601,N_9620,N_9430);
or U12602 (N_12602,N_10828,N_10349);
or U12603 (N_12603,N_9394,N_10303);
nor U12604 (N_12604,N_11992,N_11577);
and U12605 (N_12605,N_10931,N_10391);
nand U12606 (N_12606,N_9731,N_9988);
and U12607 (N_12607,N_12029,N_10809);
xnor U12608 (N_12608,N_10631,N_11471);
nand U12609 (N_12609,N_11147,N_11832);
xnor U12610 (N_12610,N_12265,N_11737);
xor U12611 (N_12611,N_10271,N_10553);
nor U12612 (N_12612,N_11893,N_10894);
xor U12613 (N_12613,N_12213,N_10750);
nand U12614 (N_12614,N_10133,N_9493);
nor U12615 (N_12615,N_11710,N_9382);
xnor U12616 (N_12616,N_11721,N_10174);
nand U12617 (N_12617,N_11054,N_11085);
nor U12618 (N_12618,N_9651,N_10808);
nand U12619 (N_12619,N_11676,N_12129);
and U12620 (N_12620,N_11594,N_9705);
or U12621 (N_12621,N_11458,N_12267);
nor U12622 (N_12622,N_10367,N_9533);
and U12623 (N_12623,N_12244,N_9664);
nor U12624 (N_12624,N_9953,N_10065);
nor U12625 (N_12625,N_12060,N_11267);
xor U12626 (N_12626,N_9802,N_9765);
or U12627 (N_12627,N_11515,N_12061);
or U12628 (N_12628,N_10386,N_10493);
nand U12629 (N_12629,N_11989,N_10657);
or U12630 (N_12630,N_9376,N_11851);
and U12631 (N_12631,N_11995,N_11301);
nor U12632 (N_12632,N_10439,N_10240);
xor U12633 (N_12633,N_10489,N_10377);
or U12634 (N_12634,N_11923,N_11523);
xnor U12635 (N_12635,N_11909,N_10855);
and U12636 (N_12636,N_9749,N_9816);
nor U12637 (N_12637,N_10169,N_9693);
and U12638 (N_12638,N_10532,N_12102);
or U12639 (N_12639,N_11690,N_11333);
nand U12640 (N_12640,N_11474,N_9815);
nand U12641 (N_12641,N_10173,N_9785);
or U12642 (N_12642,N_12363,N_12124);
or U12643 (N_12643,N_10252,N_12005);
or U12644 (N_12644,N_10909,N_11199);
or U12645 (N_12645,N_9605,N_10730);
nand U12646 (N_12646,N_11137,N_12223);
xor U12647 (N_12647,N_10041,N_11930);
nand U12648 (N_12648,N_10109,N_12171);
xor U12649 (N_12649,N_9483,N_10202);
nor U12650 (N_12650,N_12428,N_11542);
xnor U12651 (N_12651,N_12017,N_9836);
nand U12652 (N_12652,N_10988,N_11431);
xor U12653 (N_12653,N_11470,N_11440);
nand U12654 (N_12654,N_12042,N_9505);
xor U12655 (N_12655,N_11557,N_11111);
xnor U12656 (N_12656,N_10036,N_11065);
nor U12657 (N_12657,N_10130,N_9844);
nand U12658 (N_12658,N_12345,N_9535);
or U12659 (N_12659,N_9388,N_9593);
and U12660 (N_12660,N_12260,N_11309);
nand U12661 (N_12661,N_9642,N_12442);
xnor U12662 (N_12662,N_10938,N_11269);
nand U12663 (N_12663,N_10264,N_10187);
nand U12664 (N_12664,N_10902,N_9674);
or U12665 (N_12665,N_11035,N_11452);
nor U12666 (N_12666,N_12489,N_10515);
or U12667 (N_12667,N_12209,N_10559);
or U12668 (N_12668,N_9395,N_12302);
nand U12669 (N_12669,N_9796,N_10001);
xnor U12670 (N_12670,N_11578,N_12221);
nand U12671 (N_12671,N_11276,N_10942);
or U12672 (N_12672,N_11489,N_12138);
nand U12673 (N_12673,N_12463,N_11289);
or U12674 (N_12674,N_12264,N_11869);
xnor U12675 (N_12675,N_12032,N_10870);
nand U12676 (N_12676,N_12297,N_9889);
nor U12677 (N_12677,N_12116,N_12384);
nand U12678 (N_12678,N_9810,N_11154);
xor U12679 (N_12679,N_9848,N_9912);
or U12680 (N_12680,N_10008,N_10954);
or U12681 (N_12681,N_10667,N_10370);
and U12682 (N_12682,N_11102,N_9510);
xor U12683 (N_12683,N_12299,N_9562);
nor U12684 (N_12684,N_9590,N_11268);
nor U12685 (N_12685,N_9962,N_10584);
nand U12686 (N_12686,N_11376,N_9431);
nor U12687 (N_12687,N_11170,N_9672);
or U12688 (N_12688,N_9979,N_12462);
xnor U12689 (N_12689,N_11165,N_11948);
nor U12690 (N_12690,N_10312,N_9877);
and U12691 (N_12691,N_10565,N_12433);
or U12692 (N_12692,N_11161,N_11564);
nor U12693 (N_12693,N_10918,N_11666);
xor U12694 (N_12694,N_10260,N_12052);
and U12695 (N_12695,N_9484,N_9647);
nand U12696 (N_12696,N_10470,N_9787);
xor U12697 (N_12697,N_11013,N_11108);
nor U12698 (N_12698,N_9863,N_11598);
xor U12699 (N_12699,N_10897,N_10320);
and U12700 (N_12700,N_11897,N_9668);
xor U12701 (N_12701,N_10801,N_11411);
nor U12702 (N_12702,N_9514,N_12091);
nor U12703 (N_12703,N_9426,N_10154);
nor U12704 (N_12704,N_10195,N_10434);
nand U12705 (N_12705,N_10718,N_9435);
xnor U12706 (N_12706,N_11778,N_10175);
and U12707 (N_12707,N_12290,N_11983);
or U12708 (N_12708,N_10724,N_10640);
nand U12709 (N_12709,N_11106,N_9952);
nor U12710 (N_12710,N_9971,N_12099);
xnor U12711 (N_12711,N_10756,N_9767);
xor U12712 (N_12712,N_11435,N_9540);
nand U12713 (N_12713,N_12494,N_11244);
or U12714 (N_12714,N_10142,N_11976);
and U12715 (N_12715,N_9718,N_10940);
xnor U12716 (N_12716,N_11957,N_10040);
nand U12717 (N_12717,N_11355,N_9539);
nor U12718 (N_12718,N_12310,N_10785);
nand U12719 (N_12719,N_12300,N_11934);
xnor U12720 (N_12720,N_9673,N_11481);
and U12721 (N_12721,N_9829,N_10816);
and U12722 (N_12722,N_11787,N_11233);
or U12723 (N_12723,N_10458,N_10058);
nor U12724 (N_12724,N_9723,N_10210);
and U12725 (N_12725,N_12204,N_9830);
nand U12726 (N_12726,N_11965,N_10917);
or U12727 (N_12727,N_11563,N_11991);
or U12728 (N_12728,N_12126,N_9671);
nor U12729 (N_12729,N_10135,N_12003);
nor U12730 (N_12730,N_10714,N_10636);
xor U12731 (N_12731,N_10185,N_11543);
nor U12732 (N_12732,N_11829,N_9563);
nor U12733 (N_12733,N_10527,N_12224);
nand U12734 (N_12734,N_10160,N_11225);
nor U12735 (N_12735,N_11191,N_10744);
xnor U12736 (N_12736,N_11780,N_10936);
nor U12737 (N_12737,N_9455,N_10232);
or U12738 (N_12738,N_10658,N_10177);
and U12739 (N_12739,N_11801,N_11931);
xor U12740 (N_12740,N_10779,N_11266);
and U12741 (N_12741,N_11447,N_11232);
nand U12742 (N_12742,N_11653,N_11682);
nor U12743 (N_12743,N_11777,N_12283);
or U12744 (N_12744,N_12020,N_11652);
and U12745 (N_12745,N_11705,N_11617);
xor U12746 (N_12746,N_11718,N_9446);
nand U12747 (N_12747,N_11047,N_11605);
nand U12748 (N_12748,N_12379,N_10117);
nor U12749 (N_12749,N_9584,N_12389);
nor U12750 (N_12750,N_10603,N_12320);
and U12751 (N_12751,N_11545,N_9919);
or U12752 (N_12752,N_10148,N_10294);
nor U12753 (N_12753,N_11332,N_11944);
xor U12754 (N_12754,N_10953,N_11962);
nand U12755 (N_12755,N_10086,N_9783);
or U12756 (N_12756,N_10806,N_10547);
or U12757 (N_12757,N_9413,N_10015);
nand U12758 (N_12758,N_11981,N_10964);
nor U12759 (N_12759,N_9649,N_10698);
xor U12760 (N_12760,N_10318,N_10097);
nand U12761 (N_12761,N_9949,N_11726);
nor U12762 (N_12762,N_10963,N_12324);
nor U12763 (N_12763,N_11381,N_10592);
xor U12764 (N_12764,N_11240,N_11130);
xnor U12765 (N_12765,N_10328,N_12180);
or U12766 (N_12766,N_11811,N_12291);
xor U12767 (N_12767,N_11348,N_10926);
and U12768 (N_12768,N_12018,N_12359);
xor U12769 (N_12769,N_11887,N_11260);
and U12770 (N_12770,N_10395,N_11518);
xor U12771 (N_12771,N_11369,N_9965);
or U12772 (N_12772,N_12048,N_10792);
or U12773 (N_12773,N_10143,N_12134);
nor U12774 (N_12774,N_10932,N_9381);
xnor U12775 (N_12775,N_10514,N_11398);
nor U12776 (N_12776,N_10100,N_11002);
or U12777 (N_12777,N_12387,N_12226);
nand U12778 (N_12778,N_11910,N_9987);
and U12779 (N_12779,N_10793,N_12248);
and U12780 (N_12780,N_9842,N_11502);
nor U12781 (N_12781,N_12047,N_12239);
xor U12782 (N_12782,N_10136,N_11305);
nand U12783 (N_12783,N_9485,N_12054);
xor U12784 (N_12784,N_10882,N_11133);
nand U12785 (N_12785,N_10188,N_11322);
nand U12786 (N_12786,N_11649,N_10453);
nand U12787 (N_12787,N_10689,N_11422);
xor U12788 (N_12788,N_10781,N_10569);
and U12789 (N_12789,N_12306,N_11256);
and U12790 (N_12790,N_10326,N_9894);
and U12791 (N_12791,N_10052,N_10423);
nor U12792 (N_12792,N_9692,N_9405);
and U12793 (N_12793,N_10272,N_10333);
nor U12794 (N_12794,N_12208,N_11750);
or U12795 (N_12795,N_9610,N_10087);
nand U12796 (N_12796,N_11038,N_11214);
nand U12797 (N_12797,N_10956,N_10299);
nand U12798 (N_12798,N_10012,N_10522);
xnor U12799 (N_12799,N_11439,N_9733);
or U12800 (N_12800,N_10504,N_11288);
and U12801 (N_12801,N_9550,N_12081);
nor U12802 (N_12802,N_10536,N_11253);
xor U12803 (N_12803,N_11354,N_10270);
nand U12804 (N_12804,N_11501,N_11115);
or U12805 (N_12805,N_9702,N_12216);
nor U12806 (N_12806,N_12070,N_11402);
and U12807 (N_12807,N_9530,N_12163);
xnor U12808 (N_12808,N_9414,N_9613);
and U12809 (N_12809,N_11042,N_10368);
nand U12810 (N_12810,N_12377,N_11053);
and U12811 (N_12811,N_11060,N_10179);
xnor U12812 (N_12812,N_10002,N_10192);
nor U12813 (N_12813,N_12152,N_10279);
nand U12814 (N_12814,N_10805,N_12343);
xor U12815 (N_12815,N_10880,N_9956);
and U12816 (N_12816,N_10523,N_11584);
and U12817 (N_12817,N_11017,N_12482);
and U12818 (N_12818,N_9699,N_9429);
nand U12819 (N_12819,N_9888,N_9884);
nor U12820 (N_12820,N_10151,N_11669);
xor U12821 (N_12821,N_10311,N_9764);
xor U12822 (N_12822,N_9448,N_10913);
and U12823 (N_12823,N_11123,N_11784);
xor U12824 (N_12824,N_9474,N_11215);
nand U12825 (N_12825,N_12161,N_9527);
nor U12826 (N_12826,N_11670,N_12250);
and U12827 (N_12827,N_11979,N_11528);
or U12828 (N_12828,N_12013,N_9502);
nand U12829 (N_12829,N_12215,N_10482);
xor U12830 (N_12830,N_12318,N_12034);
nand U12831 (N_12831,N_9954,N_10751);
nand U12832 (N_12832,N_11377,N_9589);
nand U12833 (N_12833,N_9890,N_11374);
or U12834 (N_12834,N_10984,N_11343);
nor U12835 (N_12835,N_9701,N_9909);
nand U12836 (N_12836,N_12491,N_10836);
nand U12837 (N_12837,N_12309,N_12103);
nor U12838 (N_12838,N_10771,N_11547);
xor U12839 (N_12839,N_10732,N_11138);
or U12840 (N_12840,N_10692,N_9577);
nor U12841 (N_12841,N_12142,N_11158);
nor U12842 (N_12842,N_11634,N_11330);
or U12843 (N_12843,N_11392,N_10933);
nor U12844 (N_12844,N_10905,N_11166);
nor U12845 (N_12845,N_12222,N_12454);
nor U12846 (N_12846,N_9985,N_10042);
or U12847 (N_12847,N_9803,N_10284);
xnor U12848 (N_12848,N_12490,N_9857);
or U12849 (N_12849,N_11541,N_11835);
or U12850 (N_12850,N_11001,N_9721);
xnor U12851 (N_12851,N_12174,N_10826);
nand U12852 (N_12852,N_9421,N_11691);
nor U12853 (N_12853,N_9408,N_10627);
xor U12854 (N_12854,N_9757,N_11906);
and U12855 (N_12855,N_11865,N_9820);
or U12856 (N_12856,N_9396,N_11025);
or U12857 (N_12857,N_11293,N_12485);
or U12858 (N_12858,N_10379,N_11278);
or U12859 (N_12859,N_11824,N_11996);
and U12860 (N_12860,N_11109,N_9406);
or U12861 (N_12861,N_12408,N_9839);
nor U12862 (N_12862,N_10167,N_9986);
xnor U12863 (N_12863,N_10501,N_10297);
xnor U12864 (N_12864,N_10170,N_11234);
and U12865 (N_12865,N_9716,N_9742);
xor U12866 (N_12866,N_10034,N_11867);
and U12867 (N_12867,N_10420,N_12476);
and U12868 (N_12868,N_10823,N_12123);
nor U12869 (N_12869,N_11071,N_11254);
and U12870 (N_12870,N_10197,N_9801);
xor U12871 (N_12871,N_10021,N_12347);
and U12872 (N_12872,N_10542,N_12402);
xor U12873 (N_12873,N_9492,N_11681);
nand U12874 (N_12874,N_9631,N_10674);
nor U12875 (N_12875,N_9797,N_10991);
xor U12876 (N_12876,N_11586,N_11107);
or U12877 (N_12877,N_9831,N_11998);
xor U12878 (N_12878,N_11347,N_10017);
or U12879 (N_12879,N_12155,N_9459);
and U12880 (N_12880,N_9425,N_11913);
xnor U12881 (N_12881,N_11074,N_9740);
nand U12882 (N_12882,N_10121,N_12259);
xnor U12883 (N_12883,N_11049,N_12167);
nor U12884 (N_12884,N_9882,N_11206);
nand U12885 (N_12885,N_9977,N_10101);
nor U12886 (N_12886,N_11506,N_11766);
or U12887 (N_12887,N_12405,N_10381);
or U12888 (N_12888,N_9553,N_11717);
nor U12889 (N_12889,N_11480,N_10189);
or U12890 (N_12890,N_10587,N_9466);
xnor U12891 (N_12891,N_12380,N_11988);
and U12892 (N_12892,N_11704,N_12004);
nor U12893 (N_12893,N_11426,N_12268);
and U12894 (N_12894,N_9823,N_10459);
nand U12895 (N_12895,N_9532,N_11461);
nand U12896 (N_12896,N_10947,N_12196);
and U12897 (N_12897,N_11724,N_10208);
nor U12898 (N_12898,N_11615,N_10731);
nor U12899 (N_12899,N_10355,N_11040);
xnor U12900 (N_12900,N_9805,N_11929);
or U12901 (N_12901,N_11418,N_12094);
or U12902 (N_12902,N_11834,N_10235);
nand U12903 (N_12903,N_12214,N_10739);
xnor U12904 (N_12904,N_9519,N_11488);
nor U12905 (N_12905,N_11507,N_11202);
and U12906 (N_12906,N_11546,N_10306);
and U12907 (N_12907,N_10865,N_10056);
and U12908 (N_12908,N_12218,N_10448);
xor U12909 (N_12909,N_12464,N_9851);
or U12910 (N_12910,N_11671,N_11132);
and U12911 (N_12911,N_11524,N_9729);
nor U12912 (N_12912,N_11493,N_11771);
nor U12913 (N_12913,N_10398,N_9561);
and U12914 (N_12914,N_11486,N_10228);
nand U12915 (N_12915,N_9488,N_11514);
nand U12916 (N_12916,N_10230,N_10180);
nand U12917 (N_12917,N_11641,N_9402);
xor U12918 (N_12918,N_9508,N_9451);
or U12919 (N_12919,N_11595,N_11818);
nand U12920 (N_12920,N_9903,N_10372);
xor U12921 (N_12921,N_11101,N_9849);
xor U12922 (N_12922,N_10959,N_9378);
nand U12923 (N_12923,N_10159,N_12486);
xor U12924 (N_12924,N_12461,N_11654);
nor U12925 (N_12925,N_12366,N_11796);
nand U12926 (N_12926,N_10752,N_11762);
nor U12927 (N_12927,N_11841,N_12432);
nand U12928 (N_12928,N_12114,N_11194);
or U12929 (N_12929,N_10075,N_10665);
nand U12930 (N_12930,N_10654,N_10886);
and U12931 (N_12931,N_12354,N_9416);
nor U12932 (N_12932,N_9548,N_11261);
nor U12933 (N_12933,N_11296,N_12253);
xnor U12934 (N_12934,N_10262,N_11052);
and U12935 (N_12935,N_10581,N_11328);
nor U12936 (N_12936,N_10122,N_11419);
and U12937 (N_12937,N_11490,N_11868);
and U12938 (N_12938,N_9481,N_11770);
nand U12939 (N_12939,N_10912,N_11993);
and U12940 (N_12940,N_9895,N_9697);
xnor U12941 (N_12941,N_11243,N_10519);
nand U12942 (N_12942,N_11714,N_10877);
nand U12943 (N_12943,N_9436,N_10044);
nand U12944 (N_12944,N_11110,N_12139);
nand U12945 (N_12945,N_10994,N_12372);
nand U12946 (N_12946,N_10009,N_12059);
xor U12947 (N_12947,N_10551,N_9683);
nand U12948 (N_12948,N_11695,N_11459);
nand U12949 (N_12949,N_11856,N_11838);
and U12950 (N_12950,N_9790,N_10137);
nand U12951 (N_12951,N_11366,N_10487);
or U12952 (N_12952,N_10900,N_10105);
nor U12953 (N_12953,N_10027,N_10119);
xor U12954 (N_12954,N_12311,N_12275);
nand U12955 (N_12955,N_11902,N_11250);
xnor U12956 (N_12956,N_11416,N_10778);
xor U12957 (N_12957,N_9569,N_11927);
nor U12958 (N_12958,N_12160,N_9558);
or U12959 (N_12959,N_10903,N_12092);
or U12960 (N_12960,N_11980,N_10701);
nand U12961 (N_12961,N_10330,N_10629);
or U12962 (N_12962,N_10127,N_10211);
xor U12963 (N_12963,N_11631,N_11697);
xor U12964 (N_12964,N_10558,N_12315);
nor U12965 (N_12965,N_12173,N_9552);
xor U12966 (N_12966,N_10800,N_9753);
nor U12967 (N_12967,N_9989,N_11326);
nand U12968 (N_12968,N_9497,N_10025);
or U12969 (N_12969,N_11208,N_11284);
or U12970 (N_12970,N_9925,N_12176);
nor U12971 (N_12971,N_10971,N_11401);
nand U12972 (N_12972,N_10418,N_11952);
and U12973 (N_12973,N_11121,N_12037);
nand U12974 (N_12974,N_10300,N_12475);
or U12975 (N_12975,N_11092,N_11884);
or U12976 (N_12976,N_12427,N_11555);
nor U12977 (N_12977,N_11125,N_12230);
nand U12978 (N_12978,N_10089,N_10796);
or U12979 (N_12979,N_9564,N_12137);
or U12980 (N_12980,N_11498,N_10096);
nand U12981 (N_12981,N_9513,N_11951);
nor U12982 (N_12982,N_12327,N_9748);
nand U12983 (N_12983,N_9969,N_11752);
and U12984 (N_12984,N_11361,N_12189);
and U12985 (N_12985,N_12322,N_9415);
or U12986 (N_12986,N_9661,N_10406);
or U12987 (N_12987,N_10986,N_9546);
and U12988 (N_12988,N_11664,N_9799);
nand U12989 (N_12989,N_9591,N_10941);
nand U12990 (N_12990,N_12007,N_9997);
nand U12991 (N_12991,N_10864,N_11259);
nor U12992 (N_12992,N_11142,N_9727);
xor U12993 (N_12993,N_11687,N_10411);
or U12994 (N_12994,N_10943,N_12232);
xnor U12995 (N_12995,N_12009,N_9499);
and U12996 (N_12996,N_10219,N_11292);
and U12997 (N_12997,N_9720,N_10374);
xor U12998 (N_12998,N_12328,N_10850);
nor U12999 (N_12999,N_11279,N_12014);
or U13000 (N_13000,N_12407,N_9585);
nor U13001 (N_13001,N_9964,N_11745);
and U13002 (N_13002,N_9943,N_9469);
xor U13003 (N_13003,N_12068,N_11080);
and U13004 (N_13004,N_10521,N_11316);
nor U13005 (N_13005,N_11114,N_10073);
nor U13006 (N_13006,N_10702,N_9401);
nor U13007 (N_13007,N_12397,N_10490);
or U13008 (N_13008,N_11593,N_12287);
nand U13009 (N_13009,N_12266,N_12105);
or U13010 (N_13010,N_10859,N_9410);
nand U13011 (N_13011,N_10145,N_11499);
or U13012 (N_13012,N_10076,N_11892);
nor U13013 (N_13013,N_10513,N_10492);
nand U13014 (N_13014,N_11067,N_11707);
nand U13015 (N_13015,N_10408,N_11448);
xnor U13016 (N_13016,N_12495,N_12301);
or U13017 (N_13017,N_11467,N_11335);
and U13018 (N_13018,N_10223,N_11876);
or U13019 (N_13019,N_11875,N_10049);
and U13020 (N_13020,N_10004,N_12211);
or U13021 (N_13021,N_9486,N_10660);
nand U13022 (N_13022,N_11790,N_9665);
and U13023 (N_13023,N_11753,N_12041);
and U13024 (N_13024,N_9475,N_11183);
nor U13025 (N_13025,N_11580,N_10417);
and U13026 (N_13026,N_9901,N_12335);
and U13027 (N_13027,N_9686,N_9773);
or U13028 (N_13028,N_9471,N_12064);
nand U13029 (N_13029,N_9942,N_10608);
and U13030 (N_13030,N_9726,N_11949);
nor U13031 (N_13031,N_11131,N_9746);
nor U13032 (N_13032,N_10829,N_11383);
nor U13033 (N_13033,N_9886,N_9489);
and U13034 (N_13034,N_9526,N_9399);
nor U13035 (N_13035,N_11314,N_11665);
or U13036 (N_13036,N_12111,N_11220);
nor U13037 (N_13037,N_11187,N_10144);
xor U13038 (N_13038,N_10380,N_12172);
nand U13039 (N_13039,N_11294,N_12415);
or U13040 (N_13040,N_12496,N_9559);
and U13041 (N_13041,N_10376,N_10035);
xnor U13042 (N_13042,N_11227,N_9419);
or U13043 (N_13043,N_10181,N_9918);
nor U13044 (N_13044,N_9719,N_12125);
nand U13045 (N_13045,N_10150,N_10031);
or U13046 (N_13046,N_9932,N_12458);
xor U13047 (N_13047,N_12039,N_10907);
or U13048 (N_13048,N_11807,N_10139);
and U13049 (N_13049,N_10725,N_11907);
nand U13050 (N_13050,N_11020,N_9538);
and U13051 (N_13051,N_10769,N_11616);
xor U13052 (N_13052,N_12035,N_12245);
xnor U13053 (N_13053,N_11650,N_9892);
or U13054 (N_13054,N_10883,N_10747);
nand U13055 (N_13055,N_11325,N_9732);
and U13056 (N_13056,N_11496,N_11351);
and U13057 (N_13057,N_9972,N_10115);
nand U13058 (N_13058,N_10840,N_12206);
and U13059 (N_13059,N_10575,N_12140);
or U13060 (N_13060,N_12192,N_12376);
nor U13061 (N_13061,N_12336,N_11472);
nor U13062 (N_13062,N_11891,N_10098);
and U13063 (N_13063,N_9614,N_10839);
nor U13064 (N_13064,N_9959,N_10243);
and U13065 (N_13065,N_10969,N_12077);
or U13066 (N_13066,N_10182,N_9769);
nand U13067 (N_13067,N_11743,N_11733);
xor U13068 (N_13068,N_9400,N_9814);
nand U13069 (N_13069,N_12242,N_9660);
xor U13070 (N_13070,N_11487,N_11928);
nor U13071 (N_13071,N_11221,N_9834);
and U13072 (N_13072,N_10764,N_11638);
or U13073 (N_13073,N_10837,N_11715);
nand U13074 (N_13074,N_9961,N_11608);
xnor U13075 (N_13075,N_11432,N_10589);
nor U13076 (N_13076,N_9397,N_11193);
nand U13077 (N_13077,N_10768,N_11010);
xnor U13078 (N_13078,N_10588,N_11444);
and U13079 (N_13079,N_10535,N_10772);
xor U13080 (N_13080,N_9656,N_10365);
nand U13081 (N_13081,N_9494,N_9700);
nor U13082 (N_13082,N_12382,N_10441);
nand U13083 (N_13083,N_10019,N_12130);
nand U13084 (N_13084,N_12453,N_12416);
nor U13085 (N_13085,N_9758,N_10707);
xor U13086 (N_13086,N_11912,N_9867);
nor U13087 (N_13087,N_12079,N_10485);
or U13088 (N_13088,N_11573,N_12375);
nor U13089 (N_13089,N_10600,N_10172);
or U13090 (N_13090,N_12278,N_10615);
nor U13091 (N_13091,N_10595,N_9930);
or U13092 (N_13092,N_12423,N_11084);
and U13093 (N_13093,N_11096,N_11083);
xnor U13094 (N_13094,N_11075,N_9873);
nor U13095 (N_13095,N_10383,N_10814);
or U13096 (N_13096,N_12036,N_10321);
nor U13097 (N_13097,N_11409,N_10066);
nor U13098 (N_13098,N_10295,N_10533);
xor U13099 (N_13099,N_11521,N_9626);
and U13100 (N_13100,N_10893,N_10078);
and U13101 (N_13101,N_11331,N_10617);
nor U13102 (N_13102,N_11558,N_10313);
xor U13103 (N_13103,N_10647,N_11291);
nand U13104 (N_13104,N_9464,N_11693);
or U13105 (N_13105,N_11148,N_12233);
or U13106 (N_13106,N_10231,N_10716);
nand U13107 (N_13107,N_12016,N_12084);
and U13108 (N_13108,N_12295,N_11093);
nand U13109 (N_13109,N_10898,N_9691);
or U13110 (N_13110,N_10037,N_10023);
nor U13111 (N_13111,N_10857,N_9662);
nor U13112 (N_13112,N_11776,N_11900);
or U13113 (N_13113,N_11720,N_11719);
and U13114 (N_13114,N_10782,N_12178);
xor U13115 (N_13115,N_10471,N_12279);
or U13116 (N_13116,N_11860,N_10534);
nor U13117 (N_13117,N_11532,N_9776);
nand U13118 (N_13118,N_9615,N_10200);
xor U13119 (N_13119,N_11249,N_10479);
or U13120 (N_13120,N_10876,N_10304);
xnor U13121 (N_13121,N_11014,N_10104);
or U13122 (N_13122,N_9387,N_11986);
nor U13123 (N_13123,N_10266,N_12236);
nor U13124 (N_13124,N_10292,N_9905);
xnor U13125 (N_13125,N_9412,N_11700);
nand U13126 (N_13126,N_9573,N_10373);
nor U13127 (N_13127,N_11955,N_10438);
or U13128 (N_13128,N_11565,N_10350);
or U13129 (N_13129,N_12056,N_11162);
nand U13130 (N_13130,N_10540,N_10602);
nand U13131 (N_13131,N_10717,N_10102);
and U13132 (N_13132,N_9637,N_10989);
nand U13133 (N_13133,N_12110,N_9588);
xor U13134 (N_13134,N_11723,N_12399);
nor U13135 (N_13135,N_10360,N_12460);
or U13136 (N_13136,N_12456,N_9438);
and U13137 (N_13137,N_10951,N_11097);
xor U13138 (N_13138,N_9509,N_11635);
and U13139 (N_13139,N_10799,N_10720);
xor U13140 (N_13140,N_11972,N_10454);
xnor U13141 (N_13141,N_11273,N_11006);
and U13142 (N_13142,N_9770,N_11747);
and U13143 (N_13143,N_10112,N_10810);
and U13144 (N_13144,N_12072,N_11689);
and U13145 (N_13145,N_11275,N_11236);
and U13146 (N_13146,N_10227,N_10573);
nand U13147 (N_13147,N_10426,N_10590);
nand U13148 (N_13148,N_9375,N_10126);
nand U13149 (N_13149,N_10246,N_10663);
or U13150 (N_13150,N_10591,N_10435);
nand U13151 (N_13151,N_10339,N_10797);
or U13152 (N_13152,N_11883,N_9617);
or U13153 (N_13153,N_9926,N_11019);
or U13154 (N_13154,N_10359,N_10916);
nand U13155 (N_13155,N_11100,N_9898);
nor U13156 (N_13156,N_9951,N_10798);
nor U13157 (N_13157,N_10568,N_11285);
xor U13158 (N_13158,N_10018,N_10307);
or U13159 (N_13159,N_11731,N_9460);
or U13160 (N_13160,N_11389,N_9940);
nor U13161 (N_13161,N_11870,N_10813);
nand U13162 (N_13162,N_10709,N_11245);
and U13163 (N_13163,N_10815,N_10704);
or U13164 (N_13164,N_11384,N_10003);
xnor U13165 (N_13165,N_11530,N_11966);
nand U13166 (N_13166,N_12373,N_10464);
xor U13167 (N_13167,N_11552,N_11798);
xnor U13168 (N_13168,N_11621,N_10337);
or U13169 (N_13169,N_10345,N_12434);
xnor U13170 (N_13170,N_9845,N_11442);
nand U13171 (N_13171,N_10676,N_10444);
or U13172 (N_13172,N_11622,N_10164);
or U13173 (N_13173,N_12378,N_9874);
and U13174 (N_13174,N_11009,N_12426);
xor U13175 (N_13175,N_10888,N_11642);
and U13176 (N_13176,N_9960,N_12231);
or U13177 (N_13177,N_12292,N_10026);
or U13178 (N_13178,N_10788,N_9938);
or U13179 (N_13179,N_10116,N_10465);
or U13180 (N_13180,N_12277,N_11896);
and U13181 (N_13181,N_9479,N_9596);
nand U13182 (N_13182,N_12286,N_10664);
or U13183 (N_13183,N_10168,N_9784);
or U13184 (N_13184,N_9929,N_10682);
and U13185 (N_13185,N_10789,N_10648);
or U13186 (N_13186,N_10686,N_10118);
xor U13187 (N_13187,N_9630,N_9928);
xor U13188 (N_13188,N_9958,N_11800);
and U13189 (N_13189,N_12191,N_11511);
and U13190 (N_13190,N_11808,N_11270);
nand U13191 (N_13191,N_12089,N_10422);
nor U13192 (N_13192,N_9751,N_10650);
xnor U13193 (N_13193,N_12468,N_9608);
nor U13194 (N_13194,N_9864,N_10711);
nand U13195 (N_13195,N_11117,N_9690);
nand U13196 (N_13196,N_12356,N_11620);
or U13197 (N_13197,N_9878,N_10447);
or U13198 (N_13198,N_10924,N_10476);
nor U13199 (N_13199,N_12106,N_10432);
xnor U13200 (N_13200,N_10509,N_10111);
xor U13201 (N_13201,N_9984,N_9817);
or U13202 (N_13202,N_11300,N_10503);
nor U13203 (N_13203,N_11504,N_11373);
xnor U13204 (N_13204,N_10050,N_11522);
xnor U13205 (N_13205,N_10609,N_9795);
and U13206 (N_13206,N_11247,N_11391);
nor U13207 (N_13207,N_11589,N_10672);
and U13208 (N_13208,N_11571,N_9666);
nor U13209 (N_13209,N_12057,N_10250);
and U13210 (N_13210,N_10022,N_12296);
or U13211 (N_13211,N_10529,N_9808);
xor U13212 (N_13212,N_11767,N_10194);
and U13213 (N_13213,N_11201,N_11850);
nand U13214 (N_13214,N_11196,N_10906);
xnor U13215 (N_13215,N_9380,N_11947);
xnor U13216 (N_13216,N_11549,N_11727);
nand U13217 (N_13217,N_11607,N_9871);
nor U13218 (N_13218,N_9384,N_10719);
nor U13219 (N_13219,N_11567,N_11181);
and U13220 (N_13220,N_10652,N_9525);
xnor U13221 (N_13221,N_10178,N_11556);
xnor U13222 (N_13222,N_10765,N_10237);
and U13223 (N_13223,N_12240,N_11982);
xor U13224 (N_13224,N_11684,N_12201);
nand U13225 (N_13225,N_12212,N_12101);
xnor U13226 (N_13226,N_12141,N_10445);
and U13227 (N_13227,N_10047,N_10433);
and U13228 (N_13228,N_10545,N_10741);
and U13229 (N_13229,N_9915,N_11862);
nor U13230 (N_13230,N_10275,N_9452);
and U13231 (N_13231,N_10011,N_12383);
and U13232 (N_13232,N_10163,N_11258);
and U13233 (N_13233,N_11271,N_9433);
or U13234 (N_13234,N_10758,N_9995);
nor U13235 (N_13235,N_12252,N_10053);
or U13236 (N_13236,N_10875,N_10414);
nand U13237 (N_13237,N_9735,N_9579);
nand U13238 (N_13238,N_9440,N_10171);
xnor U13239 (N_13239,N_10308,N_11945);
nand U13240 (N_13240,N_9789,N_9679);
nand U13241 (N_13241,N_9423,N_9739);
nor U13242 (N_13242,N_10157,N_10911);
nand U13243 (N_13243,N_12457,N_10550);
nand U13244 (N_13244,N_10043,N_10451);
xor U13245 (N_13245,N_9663,N_9571);
or U13246 (N_13246,N_10759,N_10846);
nor U13247 (N_13247,N_10945,N_11171);
or U13248 (N_13248,N_11674,N_10653);
xor U13249 (N_13249,N_12391,N_10512);
nor U13250 (N_13250,N_11623,N_10344);
nand U13251 (N_13251,N_11788,N_10269);
or U13252 (N_13252,N_9506,N_11842);
or U13253 (N_13253,N_10477,N_11407);
nand U13254 (N_13254,N_9556,N_10123);
nor U13255 (N_13255,N_10935,N_10184);
nand U13256 (N_13256,N_11150,N_10474);
or U13257 (N_13257,N_11420,N_12107);
and U13258 (N_13258,N_10728,N_10425);
and U13259 (N_13259,N_11323,N_9922);
xnor U13260 (N_13260,N_10985,N_10310);
and U13261 (N_13261,N_11730,N_11899);
and U13262 (N_13262,N_12144,N_9741);
nand U13263 (N_13263,N_11802,N_9744);
nand U13264 (N_13264,N_11677,N_9422);
and U13265 (N_13265,N_10958,N_10675);
or U13266 (N_13266,N_11015,N_10261);
or U13267 (N_13267,N_10156,N_11317);
nand U13268 (N_13268,N_9463,N_11803);
nand U13269 (N_13269,N_11099,N_11823);
and U13270 (N_13270,N_12165,N_10580);
or U13271 (N_13271,N_11706,N_10939);
nor U13272 (N_13272,N_9876,N_9462);
and U13273 (N_13273,N_12076,N_11703);
nand U13274 (N_13274,N_11313,N_10394);
nor U13275 (N_13275,N_10234,N_11938);
or U13276 (N_13276,N_9973,N_9528);
nand U13277 (N_13277,N_10334,N_12393);
xor U13278 (N_13278,N_11151,N_11368);
nand U13279 (N_13279,N_12069,N_10599);
xor U13280 (N_13280,N_10429,N_10502);
nor U13281 (N_13281,N_11456,N_9576);
and U13282 (N_13282,N_12455,N_12085);
nor U13283 (N_13283,N_9937,N_11344);
and U13284 (N_13284,N_9738,N_12033);
and U13285 (N_13285,N_9780,N_11242);
and U13286 (N_13286,N_10841,N_11307);
and U13287 (N_13287,N_10624,N_11237);
xor U13288 (N_13288,N_11263,N_12219);
nor U13289 (N_13289,N_10346,N_10578);
xor U13290 (N_13290,N_11667,N_11544);
xnor U13291 (N_13291,N_10874,N_10263);
or U13292 (N_13292,N_11352,N_12118);
or U13293 (N_13293,N_11852,N_9567);
nor U13294 (N_13294,N_9933,N_10045);
or U13295 (N_13295,N_10378,N_11414);
xor U13296 (N_13296,N_10267,N_11554);
and U13297 (N_13297,N_12395,N_10072);
nand U13298 (N_13298,N_10745,N_10612);
xor U13299 (N_13299,N_10934,N_10404);
xnor U13300 (N_13300,N_11535,N_10081);
or U13301 (N_13301,N_11469,N_12414);
nor U13302 (N_13302,N_9618,N_12028);
and U13303 (N_13303,N_9712,N_10622);
xnor U13304 (N_13304,N_9503,N_11423);
and U13305 (N_13305,N_11559,N_9714);
and U13306 (N_13306,N_11126,N_9728);
and U13307 (N_13307,N_9612,N_11937);
nor U13308 (N_13308,N_11548,N_12499);
nand U13309 (N_13309,N_11327,N_10046);
or U13310 (N_13310,N_9914,N_10006);
nor U13311 (N_13311,N_11646,N_10511);
nor U13312 (N_13312,N_12194,N_9897);
nor U13313 (N_13313,N_9869,N_11579);
or U13314 (N_13314,N_10566,N_10776);
xor U13315 (N_13315,N_12096,N_9772);
and U13316 (N_13316,N_11274,N_11618);
nor U13317 (N_13317,N_10585,N_11843);
or U13318 (N_13318,N_9616,N_11772);
nand U13319 (N_13319,N_11211,N_10804);
and U13320 (N_13320,N_10000,N_12197);
or U13321 (N_13321,N_9875,N_12097);
or U13322 (N_13322,N_10204,N_10606);
or U13323 (N_13323,N_12073,N_10403);
or U13324 (N_13324,N_10833,N_10389);
xor U13325 (N_13325,N_12188,N_12255);
or U13326 (N_13326,N_12289,N_10852);
nand U13327 (N_13327,N_11306,N_11686);
and U13328 (N_13328,N_11742,N_12261);
or U13329 (N_13329,N_11387,N_10259);
and U13330 (N_13330,N_11779,N_11310);
nor U13331 (N_13331,N_11890,N_9541);
xnor U13332 (N_13332,N_10218,N_11393);
xnor U13333 (N_13333,N_12040,N_11879);
nor U13334 (N_13334,N_9543,N_12294);
and U13335 (N_13335,N_11662,N_12229);
or U13336 (N_13336,N_9648,N_10363);
xor U13337 (N_13337,N_10213,N_9657);
nor U13338 (N_13338,N_10209,N_10095);
xnor U13339 (N_13339,N_11277,N_9885);
and U13340 (N_13340,N_10998,N_11246);
xnor U13341 (N_13341,N_12390,N_10697);
nor U13342 (N_13342,N_11184,N_10293);
xnor U13343 (N_13343,N_12030,N_11610);
nor U13344 (N_13344,N_9507,N_10987);
xor U13345 (N_13345,N_10552,N_10248);
xor U13346 (N_13346,N_12471,N_11454);
or U13347 (N_13347,N_9779,N_9638);
nand U13348 (N_13348,N_12104,N_11815);
or U13349 (N_13349,N_11415,N_11881);
and U13350 (N_13350,N_12472,N_10315);
or U13351 (N_13351,N_10992,N_11064);
or U13352 (N_13352,N_11198,N_9443);
nand U13353 (N_13353,N_9482,N_11877);
or U13354 (N_13354,N_9920,N_9924);
nand U13355 (N_13355,N_10974,N_10190);
xor U13356 (N_13356,N_12364,N_10071);
or U13357 (N_13357,N_12237,N_10795);
nor U13358 (N_13358,N_12371,N_9597);
nor U13359 (N_13359,N_9955,N_11238);
nand U13360 (N_13360,N_11819,N_12170);
xnor U13361 (N_13361,N_12158,N_10217);
or U13362 (N_13362,N_12135,N_10079);
nor U13363 (N_13363,N_12417,N_12350);
or U13364 (N_13364,N_11757,N_9907);
nor U13365 (N_13365,N_11385,N_10528);
nand U13366 (N_13366,N_9389,N_11283);
nand U13367 (N_13367,N_9709,N_10525);
nor U13368 (N_13368,N_11751,N_11494);
nor U13369 (N_13369,N_11817,N_11820);
and U13370 (N_13370,N_10892,N_11954);
and U13371 (N_13371,N_10092,N_11477);
xnor U13372 (N_13372,N_11089,N_10656);
and U13373 (N_13373,N_9516,N_10574);
and U13374 (N_13374,N_9859,N_11725);
or U13375 (N_13375,N_12401,N_11141);
or U13376 (N_13376,N_11831,N_10325);
or U13377 (N_13377,N_9453,N_11026);
nand U13378 (N_13378,N_11795,N_9743);
and U13379 (N_13379,N_9689,N_12305);
and U13380 (N_13380,N_10531,N_12043);
xnor U13381 (N_13381,N_9981,N_9996);
and U13382 (N_13382,N_10134,N_11836);
nand U13383 (N_13383,N_12045,N_11953);
nor U13384 (N_13384,N_10597,N_10922);
or U13385 (N_13385,N_11412,N_9491);
xnor U13386 (N_13386,N_10863,N_11781);
nor U13387 (N_13387,N_10586,N_12431);
nor U13388 (N_13388,N_9684,N_11604);
and U13389 (N_13389,N_10322,N_10428);
and U13390 (N_13390,N_10611,N_9768);
nand U13391 (N_13391,N_9611,N_10461);
nor U13392 (N_13392,N_10452,N_10193);
xor U13393 (N_13393,N_10544,N_9404);
nand U13394 (N_13394,N_12497,N_10361);
nand U13395 (N_13395,N_12153,N_9975);
and U13396 (N_13396,N_11632,N_10484);
nor U13397 (N_13397,N_11087,N_11190);
xor U13398 (N_13398,N_9599,N_9500);
nor U13399 (N_13399,N_11866,N_11421);
xor U13400 (N_13400,N_12273,N_12063);
or U13401 (N_13401,N_11103,N_11135);
or U13402 (N_13402,N_10366,N_11847);
xnor U13403 (N_13403,N_11783,N_12258);
and U13404 (N_13404,N_9641,N_9658);
nand U13405 (N_13405,N_10419,N_12168);
or U13406 (N_13406,N_10510,N_11822);
or U13407 (N_13407,N_11613,N_12484);
or U13408 (N_13408,N_9771,N_9628);
nand U13409 (N_13409,N_11967,N_9794);
or U13410 (N_13410,N_11003,N_12331);
nand U13411 (N_13411,N_11318,N_10556);
nand U13412 (N_13412,N_11529,N_12409);
or U13413 (N_13413,N_10684,N_11839);
nor U13414 (N_13414,N_11702,N_12422);
and U13415 (N_13415,N_10901,N_9467);
nand U13416 (N_13416,N_12281,N_10968);
or U13417 (N_13417,N_10623,N_11000);
nand U13418 (N_13418,N_12438,N_10253);
xnor U13419 (N_13419,N_9855,N_10961);
xnor U13420 (N_13420,N_9825,N_10436);
or U13421 (N_13421,N_12012,N_11797);
xnor U13422 (N_13422,N_11814,N_11756);
nor U13423 (N_13423,N_12108,N_11561);
nand U13424 (N_13424,N_9557,N_9473);
xnor U13425 (N_13425,N_11044,N_11840);
nand U13426 (N_13426,N_10662,N_12429);
nor U13427 (N_13427,N_9603,N_10710);
nor U13428 (N_13428,N_10928,N_9379);
nor U13429 (N_13429,N_10726,N_12205);
xor U13430 (N_13430,N_9837,N_10084);
xor U13431 (N_13431,N_10106,N_9441);
xnor U13432 (N_13432,N_10966,N_12021);
nor U13433 (N_13433,N_9454,N_10794);
and U13434 (N_13434,N_10919,N_11680);
nand U13435 (N_13435,N_12276,N_10239);
xnor U13436 (N_13436,N_10753,N_10895);
and U13437 (N_13437,N_10524,N_11773);
nor U13438 (N_13438,N_11189,N_11863);
or U13439 (N_13439,N_11531,N_11188);
or U13440 (N_13440,N_11177,N_12062);
nor U13441 (N_13441,N_11505,N_11397);
or U13442 (N_13442,N_10405,N_12203);
or U13443 (N_13443,N_11207,N_11231);
xnor U13444 (N_13444,N_9520,N_10496);
or U13445 (N_13445,N_11468,N_10896);
nor U13446 (N_13446,N_11922,N_10074);
nor U13447 (N_13447,N_12115,N_9537);
nand U13448 (N_13448,N_10449,N_11977);
or U13449 (N_13449,N_9518,N_10060);
and U13450 (N_13450,N_10520,N_11527);
nand U13451 (N_13451,N_12082,N_10283);
xor U13452 (N_13452,N_12000,N_9945);
or U13453 (N_13453,N_11637,N_10767);
xnor U13454 (N_13454,N_9840,N_9852);
nand U13455 (N_13455,N_10099,N_10690);
nand U13456 (N_13456,N_9675,N_11360);
nand U13457 (N_13457,N_12090,N_11627);
or U13458 (N_13458,N_10186,N_9643);
nor U13459 (N_13459,N_9644,N_12314);
or U13460 (N_13460,N_11732,N_10166);
nor U13461 (N_13461,N_11086,N_11519);
nand U13462 (N_13462,N_9601,N_9908);
xor U13463 (N_13463,N_9465,N_10149);
nand U13464 (N_13464,N_12321,N_10605);
xnor U13465 (N_13465,N_11157,N_11736);
nor U13466 (N_13466,N_10777,N_9910);
xor U13467 (N_13467,N_11223,N_11936);
xor U13468 (N_13468,N_10491,N_10466);
xnor U13469 (N_13469,N_11908,N_11059);
nor U13470 (N_13470,N_12086,N_10291);
and U13471 (N_13471,N_10371,N_11337);
or U13472 (N_13472,N_9941,N_12166);
or U13473 (N_13473,N_9570,N_10548);
or U13474 (N_13474,N_11655,N_9826);
xnor U13475 (N_13475,N_9669,N_10669);
nand U13476 (N_13476,N_10203,N_9627);
and U13477 (N_13477,N_11143,N_9916);
or U13478 (N_13478,N_10356,N_12058);
nand U13479 (N_13479,N_11525,N_11063);
xor U13480 (N_13480,N_10305,N_11248);
xnor U13481 (N_13481,N_12326,N_9854);
and U13482 (N_13482,N_10146,N_10708);
and U13483 (N_13483,N_11643,N_9893);
nor U13484 (N_13484,N_9832,N_11460);
xor U13485 (N_13485,N_11363,N_10131);
nand U13486 (N_13486,N_9521,N_9498);
or U13487 (N_13487,N_11479,N_11678);
and U13488 (N_13488,N_11716,N_10069);
nor U13489 (N_13489,N_10323,N_12087);
nand U13490 (N_13490,N_9841,N_10462);
or U13491 (N_13491,N_11941,N_9781);
xnor U13492 (N_13492,N_11364,N_9420);
and U13493 (N_13493,N_10499,N_11061);
or U13494 (N_13494,N_9999,N_10677);
nand U13495 (N_13495,N_11985,N_9704);
and U13496 (N_13496,N_9819,N_10273);
or U13497 (N_13497,N_9450,N_10392);
or U13498 (N_13498,N_10646,N_11916);
nand U13499 (N_13499,N_10244,N_10460);
xor U13500 (N_13500,N_12465,N_9621);
nor U13501 (N_13501,N_11657,N_12235);
xnor U13502 (N_13502,N_11786,N_9517);
nand U13503 (N_13503,N_9578,N_11462);
and U13504 (N_13504,N_11255,N_10207);
xor U13505 (N_13505,N_11536,N_11262);
and U13506 (N_13506,N_9403,N_10153);
xor U13507 (N_13507,N_11950,N_9646);
xor U13508 (N_13508,N_12334,N_11628);
and U13509 (N_13509,N_11789,N_11282);
nor U13510 (N_13510,N_12441,N_11827);
and U13511 (N_13511,N_9980,N_9424);
nand U13512 (N_13512,N_10561,N_10757);
and U13513 (N_13513,N_11340,N_10993);
nor U13514 (N_13514,N_12049,N_11295);
nor U13515 (N_13515,N_11758,N_10415);
xor U13516 (N_13516,N_9653,N_9994);
or U13517 (N_13517,N_10442,N_11882);
nand U13518 (N_13518,N_9990,N_11463);
nand U13519 (N_13519,N_11873,N_10541);
or U13520 (N_13520,N_11324,N_9687);
nor U13521 (N_13521,N_10670,N_9670);
xnor U13522 (N_13522,N_10610,N_10039);
xor U13523 (N_13523,N_11740,N_10242);
nand U13524 (N_13524,N_10443,N_9624);
or U13525 (N_13525,N_12337,N_10324);
nor U13526 (N_13526,N_11619,N_11095);
nor U13527 (N_13527,N_9457,N_10427);
nor U13528 (N_13528,N_11590,N_10201);
nand U13529 (N_13529,N_12210,N_12303);
and U13530 (N_13530,N_11152,N_11090);
nand U13531 (N_13531,N_9522,N_10596);
nand U13532 (N_13532,N_10108,N_11738);
nand U13533 (N_13533,N_11576,N_10890);
nand U13534 (N_13534,N_9706,N_11855);
nor U13535 (N_13535,N_10770,N_11445);
xnor U13536 (N_13536,N_11630,N_11878);
or U13537 (N_13537,N_9676,N_10402);
nor U13538 (N_13538,N_10080,N_11030);
and U13539 (N_13539,N_9523,N_10245);
or U13540 (N_13540,N_11754,N_12398);
nor U13541 (N_13541,N_12157,N_10787);
or U13542 (N_13542,N_11358,N_11329);
nor U13543 (N_13543,N_11551,N_12386);
xor U13544 (N_13544,N_12338,N_12443);
nor U13545 (N_13545,N_11763,N_12271);
nand U13546 (N_13546,N_10790,N_11012);
nand U13547 (N_13547,N_11785,N_12420);
or U13548 (N_13548,N_12492,N_12293);
and U13549 (N_13549,N_9606,N_9512);
and U13550 (N_13550,N_10930,N_11235);
or U13551 (N_13551,N_10735,N_10821);
nand U13552 (N_13552,N_11539,N_10970);
nor U13553 (N_13553,N_10410,N_12341);
xnor U13554 (N_13554,N_12418,N_11864);
or U13555 (N_13555,N_11492,N_10120);
or U13556 (N_13556,N_11168,N_10390);
or U13557 (N_13557,N_10655,N_10620);
and U13558 (N_13558,N_12340,N_11999);
nor U13559 (N_13559,N_9487,N_10327);
nand U13560 (N_13560,N_11008,N_11037);
and U13561 (N_13561,N_11386,N_12128);
nand U13562 (N_13562,N_10165,N_9383);
xnor U13563 (N_13563,N_11854,N_10743);
xnor U13564 (N_13564,N_10282,N_10884);
nor U13565 (N_13565,N_10400,N_11122);
or U13566 (N_13566,N_10673,N_10226);
nand U13567 (N_13567,N_11640,N_10844);
nor U13568 (N_13568,N_11940,N_10680);
and U13569 (N_13569,N_11186,N_10681);
nor U13570 (N_13570,N_11925,N_9860);
nor U13571 (N_13571,N_9428,N_10601);
and U13572 (N_13572,N_10915,N_12362);
and U13573 (N_13573,N_10357,N_9560);
or U13574 (N_13574,N_11264,N_12002);
nor U13575 (N_13575,N_10457,N_11185);
or U13576 (N_13576,N_10424,N_10848);
xnor U13577 (N_13577,N_11178,N_10729);
or U13578 (N_13578,N_9391,N_9736);
or U13579 (N_13579,N_10538,N_9880);
or U13580 (N_13580,N_10539,N_11739);
nor U13581 (N_13581,N_10316,N_11711);
nand U13582 (N_13582,N_11491,N_10140);
xor U13583 (N_13583,N_11961,N_9575);
nor U13584 (N_13584,N_11859,N_12027);
xnor U13585 (N_13585,N_9445,N_10899);
nor U13586 (N_13586,N_11175,N_9568);
nand U13587 (N_13587,N_10887,N_11424);
xnor U13588 (N_13588,N_10666,N_10555);
nor U13589 (N_13589,N_10981,N_9715);
nand U13590 (N_13590,N_10114,N_9722);
nand U13591 (N_13591,N_11372,N_11394);
xnor U13592 (N_13592,N_11833,N_10683);
nor U13593 (N_13593,N_12051,N_10319);
nand U13594 (N_13594,N_11434,N_11476);
nand U13595 (N_13595,N_11405,N_10290);
nor U13596 (N_13596,N_10013,N_11495);
nor U13597 (N_13597,N_11280,N_12067);
nand U13598 (N_13598,N_10354,N_12195);
nor U13599 (N_13599,N_11287,N_11810);
xor U13600 (N_13600,N_11774,N_9639);
or U13601 (N_13601,N_10091,N_11503);
or U13602 (N_13602,N_11639,N_9931);
xnor U13603 (N_13603,N_10695,N_12074);
or U13604 (N_13604,N_10925,N_12050);
and U13605 (N_13605,N_11517,N_12136);
xnor U13606 (N_13606,N_9778,N_11082);
or U13607 (N_13607,N_9948,N_10176);
xor U13608 (N_13608,N_10024,N_9756);
nor U13609 (N_13609,N_9818,N_10014);
or U13610 (N_13610,N_10904,N_9504);
or U13611 (N_13611,N_10995,N_10977);
nand U13612 (N_13612,N_11651,N_11222);
nand U13613 (N_13613,N_10687,N_12411);
nand U13614 (N_13614,N_10412,N_10948);
nand U13615 (N_13615,N_10351,N_11172);
xnor U13616 (N_13616,N_11960,N_10214);
nor U13617 (N_13617,N_12424,N_9566);
nand U13618 (N_13618,N_11560,N_12182);
or U13619 (N_13619,N_10997,N_9572);
xor U13620 (N_13620,N_12394,N_9833);
xnor U13621 (N_13621,N_11990,N_12282);
nor U13622 (N_13622,N_11582,N_11566);
xor U13623 (N_13623,N_10085,N_12179);
nand U13624 (N_13624,N_10571,N_12481);
and U13625 (N_13625,N_11813,N_10820);
xnor U13626 (N_13626,N_10633,N_10742);
or U13627 (N_13627,N_10051,N_10616);
nor U13628 (N_13628,N_12288,N_11663);
xor U13629 (N_13629,N_9439,N_11905);
xnor U13630 (N_13630,N_12263,N_10286);
nor U13631 (N_13631,N_11304,N_12228);
xor U13632 (N_13632,N_10413,N_12419);
nand U13633 (N_13633,N_12075,N_10057);
and U13634 (N_13634,N_12421,N_11775);
nor U13635 (N_13635,N_12010,N_11625);
xnor U13636 (N_13636,N_11708,N_11120);
xnor U13637 (N_13637,N_9761,N_9788);
nand U13638 (N_13638,N_11942,N_11228);
xor U13639 (N_13639,N_12450,N_10070);
nand U13640 (N_13640,N_11874,N_12346);
nand U13641 (N_13641,N_11024,N_9782);
nor U13642 (N_13642,N_10914,N_10713);
or U13643 (N_13643,N_10055,N_10766);
nand U13644 (N_13644,N_11749,N_12466);
nor U13645 (N_13645,N_12055,N_9652);
xor U13646 (N_13646,N_11213,N_11371);
nor U13647 (N_13647,N_10463,N_12151);
nand U13648 (N_13648,N_11971,N_10819);
and U13649 (N_13649,N_12270,N_9470);
and U13650 (N_13650,N_11709,N_10802);
nand U13651 (N_13651,N_10480,N_12323);
and U13652 (N_13652,N_10873,N_11895);
and U13653 (N_13653,N_11599,N_11180);
or U13654 (N_13654,N_11769,N_11004);
xnor U13655 (N_13655,N_12478,N_10773);
nand U13656 (N_13656,N_11987,N_10059);
nor U13657 (N_13657,N_9725,N_10543);
nand U13658 (N_13658,N_11298,N_10475);
nand U13659 (N_13659,N_12316,N_9534);
or U13660 (N_13660,N_9461,N_10397);
or U13661 (N_13661,N_11746,N_11164);
nor U13662 (N_13662,N_9680,N_9685);
nand U13663 (N_13663,N_10375,N_12403);
xnor U13664 (N_13664,N_10562,N_11728);
nor U13665 (N_13665,N_9809,N_11648);
nor U13666 (N_13666,N_10593,N_9511);
xnor U13667 (N_13667,N_9806,N_10296);
xor U13668 (N_13668,N_9766,N_11484);
and U13669 (N_13669,N_9632,N_10257);
or U13670 (N_13670,N_10132,N_9835);
and U13671 (N_13671,N_10199,N_11427);
xor U13672 (N_13672,N_10554,N_10598);
nand U13673 (N_13673,N_10212,N_10748);
nor U13674 (N_13674,N_11005,N_11353);
or U13675 (N_13675,N_10982,N_10385);
nor U13676 (N_13676,N_11872,N_12234);
nand U13677 (N_13677,N_11205,N_11520);
nor U13678 (N_13678,N_9555,N_11583);
nor U13679 (N_13679,N_11216,N_10276);
nand U13680 (N_13680,N_10497,N_10688);
nor U13681 (N_13681,N_11978,N_10546);
and U13682 (N_13682,N_10626,N_11022);
or U13683 (N_13683,N_11516,N_9694);
or U13684 (N_13684,N_9442,N_12344);
nand U13685 (N_13685,N_11209,N_12445);
xnor U13686 (N_13686,N_9536,N_9418);
nand U13687 (N_13687,N_11029,N_11281);
xor U13688 (N_13688,N_11079,N_10331);
xor U13689 (N_13689,N_12169,N_10317);
or U13690 (N_13690,N_11915,N_11404);
nor U13691 (N_13691,N_10369,N_11290);
xnor U13692 (N_13692,N_11413,N_10811);
nand U13693 (N_13693,N_9385,N_11428);
nand U13694 (N_13694,N_11144,N_11826);
nor U13695 (N_13695,N_12448,N_12404);
and U13696 (N_13696,N_11685,N_11399);
xor U13697 (N_13697,N_9822,N_11483);
and U13698 (N_13698,N_9792,N_10030);
nor U13699 (N_13699,N_9634,N_11204);
nor U13700 (N_13700,N_10020,N_10868);
nor U13701 (N_13701,N_10225,N_11239);
nand U13702 (N_13702,N_10721,N_10537);
or U13703 (N_13703,N_11858,N_11145);
xor U13704 (N_13704,N_9906,N_12436);
and U13705 (N_13705,N_11597,N_9547);
nor U13706 (N_13706,N_10835,N_9850);
xor U13707 (N_13707,N_11362,N_10088);
nand U13708 (N_13708,N_12006,N_10843);
xnor U13709 (N_13709,N_11837,N_10929);
nor U13710 (N_13710,N_11526,N_9447);
xor U13711 (N_13711,N_11350,N_9377);
nand U13712 (N_13712,N_9944,N_10162);
or U13713 (N_13713,N_10456,N_11698);
nand U13714 (N_13714,N_11118,N_11176);
or U13715 (N_13715,N_10937,N_11601);
nand U13716 (N_13716,N_12280,N_12202);
nand U13717 (N_13717,N_10473,N_12186);
nand U13718 (N_13718,N_12046,N_10343);
or U13719 (N_13719,N_11509,N_9444);
and U13720 (N_13720,N_9654,N_11028);
nand U13721 (N_13721,N_10851,N_11603);
nand U13722 (N_13722,N_10362,N_11210);
xor U13723 (N_13723,N_11812,N_11088);
xnor U13724 (N_13724,N_11636,N_11286);
xor U13725 (N_13725,N_10927,N_11160);
nor U13726 (N_13726,N_10549,N_11735);
or U13727 (N_13727,N_11626,N_10822);
or U13728 (N_13728,N_11041,N_9752);
xnor U13729 (N_13729,N_11830,N_10972);
or U13730 (N_13730,N_11034,N_12473);
nand U13731 (N_13731,N_10818,N_11591);
nor U13732 (N_13732,N_11994,N_10399);
or U13733 (N_13733,N_11969,N_10978);
and U13734 (N_13734,N_11845,N_9762);
or U13735 (N_13735,N_10737,N_12449);
nand U13736 (N_13736,N_9991,N_12117);
xnor U13737 (N_13737,N_11203,N_11443);
and U13738 (N_13738,N_11464,N_10249);
and U13739 (N_13739,N_10358,N_11098);
xnor U13740 (N_13740,N_9640,N_9804);
or U13741 (N_13741,N_9824,N_10478);
nor U13742 (N_13742,N_9870,N_11134);
xnor U13743 (N_13743,N_11339,N_10446);
and U13744 (N_13744,N_10029,N_11970);
nor U13745 (N_13745,N_9607,N_11645);
and U13746 (N_13746,N_12352,N_10866);
or U13747 (N_13747,N_10979,N_12156);
or U13748 (N_13748,N_11585,N_10274);
nor U13749 (N_13749,N_10430,N_10340);
and U13750 (N_13750,N_10083,N_10236);
nor U13751 (N_13751,N_12477,N_11672);
xnor U13752 (N_13752,N_11964,N_11055);
xor U13753 (N_13753,N_10727,N_9707);
nor U13754 (N_13754,N_9724,N_11155);
and U13755 (N_13755,N_11077,N_11156);
or U13756 (N_13756,N_10124,N_11974);
or U13757 (N_13757,N_10158,N_10495);
nor U13758 (N_13758,N_11688,N_11917);
xor U13759 (N_13759,N_11315,N_12251);
or U13760 (N_13760,N_10644,N_9650);
or U13761 (N_13761,N_12444,N_10382);
nand U13762 (N_13762,N_12078,N_9861);
and U13763 (N_13763,N_9623,N_11308);
nor U13764 (N_13764,N_12351,N_11023);
nand U13765 (N_13765,N_10032,N_10247);
xnor U13766 (N_13766,N_10715,N_9434);
or U13767 (N_13767,N_9968,N_10206);
and U13768 (N_13768,N_10582,N_10807);
and U13769 (N_13769,N_10233,N_11946);
nand U13770 (N_13770,N_9856,N_11112);
nand U13771 (N_13771,N_11478,N_10570);
xnor U13772 (N_13772,N_11729,N_12011);
nand U13773 (N_13773,N_10094,N_11039);
nand U13774 (N_13774,N_11375,N_12109);
and U13775 (N_13775,N_10762,N_12274);
nand U13776 (N_13776,N_12093,N_10803);
and U13777 (N_13777,N_10125,N_11311);
or U13778 (N_13778,N_11094,N_11644);
and U13779 (N_13779,N_11572,N_12467);
or U13780 (N_13780,N_10572,N_10881);
or U13781 (N_13781,N_9594,N_11764);
nand U13782 (N_13782,N_12162,N_11661);
and U13783 (N_13783,N_9896,N_11921);
nand U13784 (N_13784,N_10642,N_11919);
nand U13785 (N_13785,N_9501,N_12406);
xor U13786 (N_13786,N_9708,N_11417);
and U13787 (N_13787,N_10867,N_10387);
and U13788 (N_13788,N_9496,N_9667);
xor U13789 (N_13789,N_11334,N_9476);
and U13790 (N_13790,N_10962,N_10254);
xor U13791 (N_13791,N_12150,N_9866);
nor U13792 (N_13792,N_11932,N_10847);
and U13793 (N_13793,N_12392,N_10693);
nand U13794 (N_13794,N_11119,N_10834);
nor U13795 (N_13795,N_9655,N_11197);
nor U13796 (N_13796,N_11453,N_9386);
nor U13797 (N_13797,N_11918,N_11592);
nor U13798 (N_13798,N_9495,N_11312);
nand U13799 (N_13799,N_11846,N_10229);
nor U13800 (N_13800,N_11485,N_10832);
xnor U13801 (N_13801,N_11438,N_9681);
nand U13802 (N_13802,N_10783,N_10838);
nand U13803 (N_13803,N_11760,N_10138);
xor U13804 (N_13804,N_11153,N_12348);
xor U13805 (N_13805,N_10944,N_12127);
and U13806 (N_13806,N_11903,N_9717);
or U13807 (N_13807,N_11346,N_9950);
nand U13808 (N_13808,N_11853,N_10635);
nor U13809 (N_13809,N_10530,N_11958);
or U13810 (N_13810,N_12015,N_10488);
and U13811 (N_13811,N_12190,N_11659);
nand U13812 (N_13812,N_11600,N_11748);
or U13813 (N_13813,N_10576,N_10440);
and U13814 (N_13814,N_9478,N_12370);
xor U13815 (N_13815,N_11512,N_12440);
or U13816 (N_13816,N_10353,N_9737);
nand U13817 (N_13817,N_10746,N_11370);
nor U13818 (N_13818,N_9587,N_11791);
nand U13819 (N_13819,N_12430,N_11257);
and U13820 (N_13820,N_10878,N_11425);
nand U13821 (N_13821,N_9695,N_9458);
xor U13822 (N_13822,N_10335,N_12412);
and U13823 (N_13823,N_10679,N_12200);
nand U13824 (N_13824,N_10409,N_10483);
and U13825 (N_13825,N_12031,N_11081);
nor U13826 (N_13826,N_10388,N_9713);
nand U13827 (N_13827,N_11939,N_11200);
nand U13828 (N_13828,N_11968,N_10564);
nor U13829 (N_13829,N_9549,N_11675);
or U13830 (N_13830,N_12220,N_9838);
nor U13831 (N_13831,N_9574,N_10141);
nand U13832 (N_13832,N_10812,N_10393);
xor U13833 (N_13833,N_9409,N_11179);
xor U13834 (N_13834,N_9775,N_9688);
nor U13835 (N_13835,N_12469,N_9529);
or U13836 (N_13836,N_9659,N_12317);
nor U13837 (N_13837,N_9682,N_9449);
nor U13838 (N_13838,N_10920,N_9967);
nand U13839 (N_13839,N_11408,N_11508);
nand U13840 (N_13840,N_11647,N_12008);
nor U13841 (N_13841,N_10861,N_11336);
nor U13842 (N_13842,N_12367,N_11357);
or U13843 (N_13843,N_12227,N_11534);
or U13844 (N_13844,N_9622,N_9598);
xnor U13845 (N_13845,N_11821,N_10407);
and U13846 (N_13846,N_10289,N_11457);
or U13847 (N_13847,N_12177,N_9582);
xnor U13848 (N_13848,N_10416,N_9879);
nor U13849 (N_13849,N_12133,N_11218);
xor U13850 (N_13850,N_9947,N_10763);
nor U13851 (N_13851,N_9472,N_9554);
and U13852 (N_13852,N_11382,N_10010);
xor U13853 (N_13853,N_12095,N_11804);
nor U13854 (N_13854,N_10082,N_11624);
nand U13855 (N_13855,N_12360,N_11451);
xnor U13856 (N_13856,N_10287,N_10062);
or U13857 (N_13857,N_11319,N_10879);
nand U13858 (N_13858,N_10637,N_9868);
or U13859 (N_13859,N_11683,N_11537);
nor U13860 (N_13860,N_11673,N_10740);
xnor U13861 (N_13861,N_10786,N_10508);
or U13862 (N_13862,N_9976,N_10856);
and U13863 (N_13863,N_12241,N_11792);
nor U13864 (N_13864,N_11299,N_10518);
nand U13865 (N_13865,N_10910,N_9800);
nand U13866 (N_13866,N_10630,N_11538);
xnor U13867 (N_13867,N_10760,N_9437);
xnor U13868 (N_13868,N_12333,N_9865);
and U13869 (N_13869,N_10604,N_10946);
nand U13870 (N_13870,N_11794,N_10028);
or U13871 (N_13871,N_10038,N_12285);
nor U13872 (N_13872,N_12023,N_10952);
or U13873 (N_13873,N_10486,N_10967);
or U13874 (N_13874,N_9490,N_11043);
nand U13875 (N_13875,N_12257,N_10224);
nor U13876 (N_13876,N_10507,N_11699);
nor U13877 (N_13877,N_11553,N_10827);
or U13878 (N_13878,N_10871,N_10277);
or U13879 (N_13879,N_10161,N_9411);
or U13880 (N_13880,N_10632,N_12396);
nand U13881 (N_13881,N_11302,N_9828);
and U13882 (N_13882,N_12358,N_12361);
nor U13883 (N_13883,N_12164,N_9609);
xnor U13884 (N_13884,N_12269,N_10659);
or U13885 (N_13885,N_10628,N_10481);
xnor U13886 (N_13886,N_12304,N_11611);
or U13887 (N_13887,N_10064,N_10621);
or U13888 (N_13888,N_9392,N_11889);
nand U13889 (N_13889,N_11146,N_10215);
and U13890 (N_13890,N_10469,N_10342);
and U13891 (N_13891,N_9390,N_11848);
nand U13892 (N_13892,N_11045,N_10258);
or U13893 (N_13893,N_9853,N_12185);
nor U13894 (N_13894,N_11078,N_11575);
or U13895 (N_13895,N_10498,N_11050);
or U13896 (N_13896,N_12339,N_9813);
or U13897 (N_13897,N_10128,N_10309);
nand U13898 (N_13898,N_10288,N_10516);
xnor U13899 (N_13899,N_10352,N_10784);
nor U13900 (N_13900,N_9974,N_12159);
nor U13901 (N_13901,N_9807,N_11051);
or U13902 (N_13902,N_11027,N_9927);
xor U13903 (N_13903,N_10699,N_11169);
nor U13904 (N_13904,N_12022,N_10705);
nor U13905 (N_13905,N_11997,N_10723);
or U13906 (N_13906,N_11768,N_9812);
nand U13907 (N_13907,N_11926,N_10191);
nor U13908 (N_13908,N_10147,N_11219);
and U13909 (N_13909,N_12262,N_10661);
and U13910 (N_13910,N_9551,N_10238);
nor U13911 (N_13911,N_11033,N_11379);
or U13912 (N_13912,N_10455,N_11032);
nand U13913 (N_13913,N_11497,N_12247);
nor U13914 (N_13914,N_11116,N_11388);
nand U13915 (N_13915,N_9777,N_10634);
and U13916 (N_13916,N_9793,N_9904);
and U13917 (N_13917,N_9477,N_11861);
nand U13918 (N_13918,N_10734,N_9872);
or U13919 (N_13919,N_9619,N_10869);
and U13920 (N_13920,N_11031,N_12146);
nor U13921 (N_13921,N_11612,N_10285);
nand U13922 (N_13922,N_9774,N_9846);
or U13923 (N_13923,N_9946,N_12493);
nor U13924 (N_13924,N_11446,N_10216);
nor U13925 (N_13925,N_10949,N_9887);
nand U13926 (N_13926,N_10671,N_10016);
nand U13927 (N_13927,N_10733,N_11793);
nor U13928 (N_13928,N_12349,N_11602);
or U13929 (N_13929,N_12355,N_11510);
xor U13930 (N_13930,N_12329,N_10950);
nor U13931 (N_13931,N_12026,N_9921);
nor U13932 (N_13932,N_11924,N_10577);
or U13933 (N_13933,N_10613,N_11694);
xor U13934 (N_13934,N_12181,N_12368);
nor U13935 (N_13935,N_11149,N_11429);
xor U13936 (N_13936,N_11056,N_9633);
nor U13937 (N_13937,N_10005,N_10817);
nand U13938 (N_13938,N_11943,N_10738);
xor U13939 (N_13939,N_9586,N_10067);
xor U13940 (N_13940,N_10694,N_9899);
xnor U13941 (N_13941,N_11433,N_10845);
nor U13942 (N_13942,N_10517,N_9934);
or U13943 (N_13943,N_10220,N_11570);
and U13944 (N_13944,N_9734,N_11963);
nor U13945 (N_13945,N_10205,N_11105);
xor U13946 (N_13946,N_11587,N_10268);
nand U13947 (N_13947,N_11072,N_11062);
xor U13948 (N_13948,N_10183,N_10761);
xnor U13949 (N_13949,N_12083,N_11828);
nor U13950 (N_13950,N_12446,N_10712);
xnor U13951 (N_13951,N_12388,N_9883);
xor U13952 (N_13952,N_11473,N_12470);
nor U13953 (N_13953,N_10068,N_12217);
or U13954 (N_13954,N_10594,N_10583);
nor U13955 (N_13955,N_10990,N_10831);
xor U13956 (N_13956,N_10889,N_12024);
and U13957 (N_13957,N_11656,N_11441);
xnor U13958 (N_13958,N_11380,N_11229);
nor U13959 (N_13959,N_11449,N_11365);
or U13960 (N_13960,N_11124,N_10431);
nor U13961 (N_13961,N_10467,N_12001);
and U13962 (N_13962,N_9398,N_12435);
nand U13963 (N_13963,N_11378,N_10579);
nand U13964 (N_13964,N_9745,N_11192);
or U13965 (N_13965,N_12025,N_11562);
or U13966 (N_13966,N_11016,N_12184);
xor U13967 (N_13967,N_11252,N_11159);
xnor U13968 (N_13968,N_9393,N_10975);
or U13969 (N_13969,N_10255,N_12439);
and U13970 (N_13970,N_9531,N_10563);
nor U13971 (N_13971,N_10302,N_11482);
and U13972 (N_13972,N_10557,N_11782);
xnor U13973 (N_13973,N_11356,N_10957);
and U13974 (N_13974,N_11761,N_11396);
or U13975 (N_13975,N_9583,N_12425);
nand U13976 (N_13976,N_10619,N_11614);
nor U13977 (N_13977,N_12332,N_11230);
nand U13978 (N_13978,N_12121,N_12198);
nand U13979 (N_13979,N_12385,N_10364);
or U13980 (N_13980,N_10999,N_11658);
nor U13981 (N_13981,N_10567,N_11182);
xnor U13982 (N_13982,N_11911,N_11212);
nor U13983 (N_13983,N_12199,N_9595);
and U13984 (N_13984,N_12019,N_11140);
xnor U13985 (N_13985,N_11894,N_10754);
nor U13986 (N_13986,N_11400,N_9677);
xor U13987 (N_13987,N_10241,N_11755);
nor U13988 (N_13988,N_10505,N_11765);
nor U13989 (N_13989,N_11217,N_10976);
or U13990 (N_13990,N_10825,N_11251);
xor U13991 (N_13991,N_9963,N_11406);
or U13992 (N_13992,N_9911,N_10437);
nand U13993 (N_13993,N_11857,N_9791);
and U13994 (N_13994,N_10703,N_9939);
and U13995 (N_13995,N_11436,N_11403);
xor U13996 (N_13996,N_12044,N_9798);
xnor U13997 (N_13997,N_12131,N_9821);
nand U13998 (N_13998,N_12249,N_10780);
nor U13999 (N_13999,N_10755,N_11195);
and U14000 (N_14000,N_11070,N_10983);
or U14001 (N_14001,N_10222,N_9710);
nand U14002 (N_14002,N_10526,N_10824);
or U14003 (N_14003,N_10155,N_11046);
nand U14004 (N_14004,N_11410,N_9524);
nand U14005 (N_14005,N_11973,N_10196);
or U14006 (N_14006,N_9917,N_9592);
or U14007 (N_14007,N_11588,N_12143);
xor U14008 (N_14008,N_12183,N_10996);
nor U14009 (N_14009,N_12452,N_10048);
nor U14010 (N_14010,N_9978,N_9811);
xnor U14011 (N_14011,N_9763,N_11825);
xnor U14012 (N_14012,N_10129,N_11450);
nand U14013 (N_14013,N_10614,N_11173);
nor U14014 (N_14014,N_10860,N_9635);
or U14015 (N_14015,N_11349,N_10651);
nor U14016 (N_14016,N_10649,N_12207);
or U14017 (N_14017,N_11338,N_10251);
or U14018 (N_14018,N_11568,N_10348);
or U14019 (N_14019,N_11734,N_9993);
nand U14020 (N_14020,N_12298,N_9625);
nor U14021 (N_14021,N_11844,N_10849);
nand U14022 (N_14022,N_12307,N_12498);
nand U14023 (N_14023,N_11104,N_9750);
nor U14024 (N_14024,N_12319,N_12100);
nor U14025 (N_14025,N_9900,N_11341);
nor U14026 (N_14026,N_11021,N_11975);
xor U14027 (N_14027,N_9456,N_10923);
xnor U14028 (N_14028,N_11569,N_10960);
and U14029 (N_14029,N_12088,N_10862);
and U14030 (N_14030,N_9759,N_11066);
nor U14031 (N_14031,N_11660,N_12413);
nand U14032 (N_14032,N_9923,N_9600);
and U14033 (N_14033,N_10278,N_10696);
or U14034 (N_14034,N_12325,N_10872);
and U14035 (N_14035,N_11722,N_12175);
or U14036 (N_14036,N_10421,N_10107);
or U14037 (N_14037,N_11466,N_12254);
nor U14038 (N_14038,N_11500,N_9760);
and U14039 (N_14039,N_9580,N_11113);
nor U14040 (N_14040,N_11956,N_11805);
xor U14041 (N_14041,N_10641,N_9983);
and U14042 (N_14042,N_9678,N_11320);
nand U14043 (N_14043,N_10341,N_12113);
and U14044 (N_14044,N_10007,N_11048);
nand U14045 (N_14045,N_10722,N_11816);
or U14046 (N_14046,N_12369,N_10643);
or U14047 (N_14047,N_12193,N_9862);
and U14048 (N_14048,N_11668,N_11933);
nor U14049 (N_14049,N_10384,N_9432);
and U14050 (N_14050,N_9935,N_11901);
nand U14051 (N_14051,N_11581,N_11127);
or U14052 (N_14052,N_10061,N_10639);
xor U14053 (N_14053,N_9703,N_9629);
and U14054 (N_14054,N_12381,N_11139);
and U14055 (N_14055,N_12098,N_11935);
and U14056 (N_14056,N_12246,N_11904);
and U14057 (N_14057,N_11759,N_11058);
xor U14058 (N_14058,N_11475,N_11007);
nand U14059 (N_14059,N_10472,N_11898);
and U14060 (N_14060,N_9982,N_11303);
xor U14061 (N_14061,N_12488,N_11513);
or U14062 (N_14062,N_12400,N_11097);
nand U14063 (N_14063,N_10211,N_11601);
nand U14064 (N_14064,N_9542,N_11751);
nand U14065 (N_14065,N_9599,N_9881);
and U14066 (N_14066,N_10117,N_10869);
and U14067 (N_14067,N_10394,N_12427);
nand U14068 (N_14068,N_9720,N_12281);
xor U14069 (N_14069,N_11179,N_9614);
nand U14070 (N_14070,N_11612,N_11018);
or U14071 (N_14071,N_10172,N_10990);
or U14072 (N_14072,N_10573,N_9718);
nor U14073 (N_14073,N_9376,N_11348);
nor U14074 (N_14074,N_10376,N_9451);
or U14075 (N_14075,N_11301,N_9994);
nand U14076 (N_14076,N_10303,N_10431);
and U14077 (N_14077,N_10359,N_11166);
xor U14078 (N_14078,N_9530,N_9552);
and U14079 (N_14079,N_10846,N_10240);
xor U14080 (N_14080,N_10594,N_9890);
or U14081 (N_14081,N_11290,N_10828);
nor U14082 (N_14082,N_10094,N_10606);
or U14083 (N_14083,N_10868,N_11539);
xor U14084 (N_14084,N_11697,N_11970);
nand U14085 (N_14085,N_12074,N_11488);
and U14086 (N_14086,N_12249,N_9514);
xor U14087 (N_14087,N_11442,N_10054);
xor U14088 (N_14088,N_9688,N_12276);
nor U14089 (N_14089,N_10103,N_10523);
nand U14090 (N_14090,N_11226,N_12389);
or U14091 (N_14091,N_10683,N_12398);
nor U14092 (N_14092,N_11102,N_10263);
or U14093 (N_14093,N_9546,N_10693);
nand U14094 (N_14094,N_10534,N_11840);
nand U14095 (N_14095,N_10338,N_10019);
nor U14096 (N_14096,N_10080,N_9884);
nor U14097 (N_14097,N_10161,N_11575);
or U14098 (N_14098,N_9712,N_11092);
or U14099 (N_14099,N_10063,N_12073);
nor U14100 (N_14100,N_10773,N_11535);
nand U14101 (N_14101,N_9689,N_10235);
xnor U14102 (N_14102,N_9426,N_12239);
and U14103 (N_14103,N_9481,N_11186);
nand U14104 (N_14104,N_9772,N_10876);
nor U14105 (N_14105,N_11150,N_9681);
nor U14106 (N_14106,N_9981,N_11917);
and U14107 (N_14107,N_10517,N_11571);
or U14108 (N_14108,N_10269,N_11173);
or U14109 (N_14109,N_10352,N_9492);
xnor U14110 (N_14110,N_9486,N_12330);
or U14111 (N_14111,N_12109,N_12382);
xnor U14112 (N_14112,N_9760,N_12293);
nor U14113 (N_14113,N_9740,N_11649);
and U14114 (N_14114,N_9376,N_12096);
or U14115 (N_14115,N_10482,N_9633);
nor U14116 (N_14116,N_11400,N_11471);
or U14117 (N_14117,N_12349,N_10975);
nor U14118 (N_14118,N_10964,N_11352);
nor U14119 (N_14119,N_10386,N_10459);
xor U14120 (N_14120,N_11667,N_11467);
xnor U14121 (N_14121,N_10620,N_12042);
nand U14122 (N_14122,N_12038,N_10999);
and U14123 (N_14123,N_10092,N_11382);
nor U14124 (N_14124,N_10758,N_10492);
xnor U14125 (N_14125,N_9415,N_11438);
xor U14126 (N_14126,N_10525,N_10930);
nor U14127 (N_14127,N_9544,N_11271);
nor U14128 (N_14128,N_9553,N_12111);
or U14129 (N_14129,N_10581,N_12177);
or U14130 (N_14130,N_11016,N_9646);
nand U14131 (N_14131,N_11666,N_10763);
and U14132 (N_14132,N_9627,N_10870);
nor U14133 (N_14133,N_9610,N_10578);
and U14134 (N_14134,N_9830,N_11921);
nand U14135 (N_14135,N_9988,N_10269);
and U14136 (N_14136,N_10803,N_10343);
and U14137 (N_14137,N_12463,N_10055);
nor U14138 (N_14138,N_12458,N_12361);
nand U14139 (N_14139,N_10651,N_10896);
or U14140 (N_14140,N_9991,N_12372);
or U14141 (N_14141,N_10751,N_11662);
and U14142 (N_14142,N_10764,N_9606);
nor U14143 (N_14143,N_10927,N_11522);
and U14144 (N_14144,N_12247,N_11695);
xnor U14145 (N_14145,N_9951,N_12038);
or U14146 (N_14146,N_10314,N_11444);
or U14147 (N_14147,N_9869,N_11862);
nor U14148 (N_14148,N_12426,N_12267);
nand U14149 (N_14149,N_10357,N_10692);
xor U14150 (N_14150,N_12043,N_10103);
nor U14151 (N_14151,N_9645,N_10899);
nor U14152 (N_14152,N_9378,N_9656);
or U14153 (N_14153,N_11236,N_10226);
nor U14154 (N_14154,N_10948,N_11828);
nand U14155 (N_14155,N_9584,N_9491);
nand U14156 (N_14156,N_10655,N_12436);
nor U14157 (N_14157,N_12461,N_10574);
and U14158 (N_14158,N_11290,N_11099);
xor U14159 (N_14159,N_9999,N_11146);
nor U14160 (N_14160,N_9690,N_10637);
nor U14161 (N_14161,N_11974,N_11786);
or U14162 (N_14162,N_9435,N_11585);
or U14163 (N_14163,N_10412,N_10511);
nor U14164 (N_14164,N_12298,N_10835);
nor U14165 (N_14165,N_12121,N_10886);
nor U14166 (N_14166,N_12194,N_12227);
or U14167 (N_14167,N_9505,N_9427);
xor U14168 (N_14168,N_11476,N_9626);
and U14169 (N_14169,N_10533,N_11362);
and U14170 (N_14170,N_10497,N_9674);
nand U14171 (N_14171,N_9830,N_12249);
and U14172 (N_14172,N_12199,N_9723);
xor U14173 (N_14173,N_10856,N_9666);
nand U14174 (N_14174,N_9405,N_12200);
nand U14175 (N_14175,N_12128,N_11110);
and U14176 (N_14176,N_11430,N_11119);
xnor U14177 (N_14177,N_12391,N_11541);
xnor U14178 (N_14178,N_9915,N_12209);
xnor U14179 (N_14179,N_10809,N_12232);
nor U14180 (N_14180,N_10258,N_12386);
and U14181 (N_14181,N_10908,N_10201);
or U14182 (N_14182,N_11812,N_10395);
nand U14183 (N_14183,N_12401,N_12023);
xnor U14184 (N_14184,N_10164,N_12064);
and U14185 (N_14185,N_12499,N_12182);
or U14186 (N_14186,N_10093,N_10611);
nand U14187 (N_14187,N_10585,N_11646);
nor U14188 (N_14188,N_10197,N_9816);
xnor U14189 (N_14189,N_9884,N_9661);
or U14190 (N_14190,N_10955,N_11438);
and U14191 (N_14191,N_12173,N_11479);
and U14192 (N_14192,N_10575,N_10105);
and U14193 (N_14193,N_10952,N_9764);
nor U14194 (N_14194,N_11283,N_10649);
nand U14195 (N_14195,N_10803,N_11005);
nand U14196 (N_14196,N_10652,N_11935);
xnor U14197 (N_14197,N_9467,N_10880);
or U14198 (N_14198,N_9850,N_9779);
nand U14199 (N_14199,N_12194,N_9869);
or U14200 (N_14200,N_11926,N_11712);
or U14201 (N_14201,N_12206,N_11955);
nor U14202 (N_14202,N_9399,N_9705);
xor U14203 (N_14203,N_11999,N_10323);
nor U14204 (N_14204,N_10009,N_11213);
and U14205 (N_14205,N_9904,N_9508);
xor U14206 (N_14206,N_10460,N_9649);
and U14207 (N_14207,N_11418,N_12193);
and U14208 (N_14208,N_9434,N_9775);
and U14209 (N_14209,N_9387,N_12336);
xor U14210 (N_14210,N_12452,N_10420);
nor U14211 (N_14211,N_11893,N_12196);
and U14212 (N_14212,N_10919,N_11165);
and U14213 (N_14213,N_9680,N_10990);
nor U14214 (N_14214,N_10744,N_11970);
or U14215 (N_14215,N_10952,N_11563);
and U14216 (N_14216,N_12382,N_12031);
and U14217 (N_14217,N_11164,N_10672);
and U14218 (N_14218,N_10976,N_11559);
and U14219 (N_14219,N_11280,N_9388);
nor U14220 (N_14220,N_11950,N_10610);
nor U14221 (N_14221,N_10189,N_11929);
and U14222 (N_14222,N_11896,N_11545);
xnor U14223 (N_14223,N_11389,N_12383);
and U14224 (N_14224,N_10906,N_11941);
and U14225 (N_14225,N_9443,N_10709);
xor U14226 (N_14226,N_10982,N_10117);
nand U14227 (N_14227,N_11893,N_9609);
nand U14228 (N_14228,N_10998,N_10113);
and U14229 (N_14229,N_12283,N_10682);
or U14230 (N_14230,N_11648,N_11646);
or U14231 (N_14231,N_11576,N_10361);
nor U14232 (N_14232,N_11213,N_9397);
nor U14233 (N_14233,N_10779,N_10050);
nand U14234 (N_14234,N_11359,N_11610);
nand U14235 (N_14235,N_10980,N_12169);
xor U14236 (N_14236,N_9409,N_11187);
nor U14237 (N_14237,N_11381,N_10982);
xor U14238 (N_14238,N_10727,N_11919);
xor U14239 (N_14239,N_11532,N_10749);
or U14240 (N_14240,N_11460,N_9837);
and U14241 (N_14241,N_12106,N_10897);
xnor U14242 (N_14242,N_12110,N_11594);
or U14243 (N_14243,N_10513,N_11554);
nand U14244 (N_14244,N_9504,N_12106);
xnor U14245 (N_14245,N_10902,N_10576);
xnor U14246 (N_14246,N_9568,N_11173);
or U14247 (N_14247,N_12065,N_9924);
and U14248 (N_14248,N_10459,N_11050);
and U14249 (N_14249,N_9402,N_12070);
xor U14250 (N_14250,N_11244,N_12206);
nor U14251 (N_14251,N_11811,N_10097);
or U14252 (N_14252,N_10659,N_11646);
nor U14253 (N_14253,N_10530,N_11181);
and U14254 (N_14254,N_11295,N_9441);
or U14255 (N_14255,N_12231,N_9894);
xnor U14256 (N_14256,N_9831,N_12044);
nand U14257 (N_14257,N_11605,N_11856);
xnor U14258 (N_14258,N_10443,N_9518);
or U14259 (N_14259,N_10226,N_10040);
xor U14260 (N_14260,N_11628,N_10334);
nand U14261 (N_14261,N_10504,N_10638);
and U14262 (N_14262,N_12392,N_9409);
and U14263 (N_14263,N_11899,N_11539);
nor U14264 (N_14264,N_10538,N_10046);
or U14265 (N_14265,N_10213,N_11116);
or U14266 (N_14266,N_10916,N_11664);
nand U14267 (N_14267,N_10052,N_10016);
xor U14268 (N_14268,N_10702,N_9548);
or U14269 (N_14269,N_11479,N_10951);
xnor U14270 (N_14270,N_11154,N_12144);
or U14271 (N_14271,N_9710,N_10791);
nand U14272 (N_14272,N_12296,N_10221);
xnor U14273 (N_14273,N_11624,N_10457);
xor U14274 (N_14274,N_9642,N_9565);
and U14275 (N_14275,N_10811,N_11147);
xor U14276 (N_14276,N_12007,N_12254);
nor U14277 (N_14277,N_11799,N_11015);
and U14278 (N_14278,N_11808,N_11181);
nand U14279 (N_14279,N_9559,N_9633);
or U14280 (N_14280,N_12110,N_12246);
xor U14281 (N_14281,N_11731,N_11471);
xnor U14282 (N_14282,N_11443,N_11193);
nand U14283 (N_14283,N_10239,N_9571);
nand U14284 (N_14284,N_11849,N_9886);
nand U14285 (N_14285,N_12071,N_9610);
or U14286 (N_14286,N_9830,N_10531);
nand U14287 (N_14287,N_12033,N_10704);
or U14288 (N_14288,N_11152,N_12070);
or U14289 (N_14289,N_9924,N_12440);
and U14290 (N_14290,N_9885,N_12498);
nor U14291 (N_14291,N_10617,N_10757);
xor U14292 (N_14292,N_9627,N_11774);
nor U14293 (N_14293,N_10085,N_10014);
or U14294 (N_14294,N_10064,N_11498);
and U14295 (N_14295,N_11760,N_11178);
and U14296 (N_14296,N_12219,N_10585);
nand U14297 (N_14297,N_9593,N_9447);
nand U14298 (N_14298,N_10248,N_10920);
xor U14299 (N_14299,N_10172,N_9557);
xnor U14300 (N_14300,N_9960,N_9580);
or U14301 (N_14301,N_12078,N_10608);
and U14302 (N_14302,N_11424,N_12311);
or U14303 (N_14303,N_10388,N_10648);
or U14304 (N_14304,N_9800,N_12049);
nand U14305 (N_14305,N_11208,N_10737);
or U14306 (N_14306,N_9470,N_10559);
and U14307 (N_14307,N_12376,N_10888);
or U14308 (N_14308,N_10825,N_9518);
xnor U14309 (N_14309,N_11965,N_10137);
xor U14310 (N_14310,N_9877,N_10844);
or U14311 (N_14311,N_12242,N_9546);
nand U14312 (N_14312,N_9894,N_10790);
nor U14313 (N_14313,N_10599,N_9568);
nand U14314 (N_14314,N_11011,N_11358);
nor U14315 (N_14315,N_9597,N_11846);
nor U14316 (N_14316,N_12385,N_10606);
nor U14317 (N_14317,N_9528,N_9510);
or U14318 (N_14318,N_11117,N_11390);
or U14319 (N_14319,N_11064,N_11424);
xnor U14320 (N_14320,N_11473,N_12335);
nand U14321 (N_14321,N_12008,N_10604);
and U14322 (N_14322,N_11776,N_9583);
nor U14323 (N_14323,N_10012,N_9594);
nor U14324 (N_14324,N_11595,N_9382);
or U14325 (N_14325,N_10999,N_9589);
or U14326 (N_14326,N_9376,N_11558);
and U14327 (N_14327,N_11355,N_11869);
nand U14328 (N_14328,N_12016,N_9710);
nor U14329 (N_14329,N_12383,N_10129);
and U14330 (N_14330,N_10095,N_10269);
or U14331 (N_14331,N_11599,N_11019);
xnor U14332 (N_14332,N_9694,N_12469);
xnor U14333 (N_14333,N_12377,N_10735);
nor U14334 (N_14334,N_10893,N_12225);
nand U14335 (N_14335,N_10384,N_11034);
or U14336 (N_14336,N_12260,N_11153);
nand U14337 (N_14337,N_10659,N_12378);
and U14338 (N_14338,N_10191,N_9734);
xnor U14339 (N_14339,N_12299,N_10355);
xnor U14340 (N_14340,N_10757,N_10467);
nand U14341 (N_14341,N_11579,N_9948);
or U14342 (N_14342,N_11477,N_11406);
nor U14343 (N_14343,N_10332,N_11312);
or U14344 (N_14344,N_10636,N_10200);
nor U14345 (N_14345,N_9597,N_10311);
nor U14346 (N_14346,N_9420,N_9647);
or U14347 (N_14347,N_10391,N_11380);
nor U14348 (N_14348,N_10595,N_10927);
nor U14349 (N_14349,N_9468,N_11242);
nor U14350 (N_14350,N_11979,N_9714);
nor U14351 (N_14351,N_11947,N_11093);
nor U14352 (N_14352,N_10040,N_10931);
or U14353 (N_14353,N_9437,N_11724);
or U14354 (N_14354,N_12343,N_11630);
and U14355 (N_14355,N_11511,N_10149);
or U14356 (N_14356,N_11265,N_9809);
nor U14357 (N_14357,N_12411,N_11797);
and U14358 (N_14358,N_11325,N_9471);
xor U14359 (N_14359,N_9665,N_9882);
nand U14360 (N_14360,N_10635,N_10796);
xnor U14361 (N_14361,N_12090,N_10515);
or U14362 (N_14362,N_12439,N_11391);
or U14363 (N_14363,N_10919,N_10761);
nand U14364 (N_14364,N_10505,N_9412);
or U14365 (N_14365,N_10226,N_11701);
or U14366 (N_14366,N_9411,N_10444);
xor U14367 (N_14367,N_10566,N_11455);
xnor U14368 (N_14368,N_10497,N_9681);
nor U14369 (N_14369,N_10525,N_9808);
and U14370 (N_14370,N_11139,N_12175);
nand U14371 (N_14371,N_11659,N_9776);
nor U14372 (N_14372,N_11248,N_12202);
and U14373 (N_14373,N_9714,N_10486);
nand U14374 (N_14374,N_10601,N_10783);
nor U14375 (N_14375,N_11882,N_10700);
nand U14376 (N_14376,N_12396,N_10851);
or U14377 (N_14377,N_9718,N_12336);
nand U14378 (N_14378,N_9387,N_10580);
xor U14379 (N_14379,N_10597,N_10268);
xnor U14380 (N_14380,N_10516,N_10896);
nor U14381 (N_14381,N_11756,N_10938);
xor U14382 (N_14382,N_9621,N_12477);
xor U14383 (N_14383,N_11965,N_11578);
nor U14384 (N_14384,N_11632,N_12427);
nand U14385 (N_14385,N_9670,N_12179);
xnor U14386 (N_14386,N_9845,N_10677);
xor U14387 (N_14387,N_11212,N_9382);
or U14388 (N_14388,N_11557,N_11088);
and U14389 (N_14389,N_10129,N_12242);
and U14390 (N_14390,N_10470,N_11093);
nor U14391 (N_14391,N_12419,N_10180);
and U14392 (N_14392,N_12135,N_9754);
nand U14393 (N_14393,N_9882,N_12046);
xnor U14394 (N_14394,N_12240,N_10496);
or U14395 (N_14395,N_10327,N_10172);
xor U14396 (N_14396,N_12017,N_9390);
and U14397 (N_14397,N_9950,N_11326);
nand U14398 (N_14398,N_10359,N_10000);
or U14399 (N_14399,N_11987,N_11530);
nand U14400 (N_14400,N_11473,N_9995);
xnor U14401 (N_14401,N_9574,N_12019);
and U14402 (N_14402,N_11036,N_9937);
or U14403 (N_14403,N_9669,N_11453);
and U14404 (N_14404,N_10642,N_12355);
or U14405 (N_14405,N_10200,N_10901);
or U14406 (N_14406,N_12014,N_9996);
xnor U14407 (N_14407,N_9696,N_11147);
or U14408 (N_14408,N_11350,N_9680);
xnor U14409 (N_14409,N_9643,N_10636);
or U14410 (N_14410,N_11057,N_9917);
nor U14411 (N_14411,N_9584,N_9891);
nor U14412 (N_14412,N_10748,N_10018);
xnor U14413 (N_14413,N_11165,N_9540);
nand U14414 (N_14414,N_11934,N_11730);
nand U14415 (N_14415,N_12024,N_11509);
xnor U14416 (N_14416,N_11370,N_9611);
or U14417 (N_14417,N_10800,N_9448);
or U14418 (N_14418,N_10330,N_9735);
xnor U14419 (N_14419,N_10941,N_10205);
and U14420 (N_14420,N_10830,N_12250);
nand U14421 (N_14421,N_11930,N_12270);
and U14422 (N_14422,N_10236,N_10679);
xnor U14423 (N_14423,N_11753,N_10803);
nand U14424 (N_14424,N_10365,N_9897);
nor U14425 (N_14425,N_9919,N_12116);
and U14426 (N_14426,N_10416,N_11238);
nor U14427 (N_14427,N_11858,N_12428);
nand U14428 (N_14428,N_11383,N_11801);
or U14429 (N_14429,N_9598,N_11500);
xor U14430 (N_14430,N_10076,N_12214);
xnor U14431 (N_14431,N_10471,N_12086);
and U14432 (N_14432,N_11113,N_9576);
nand U14433 (N_14433,N_12232,N_9803);
xnor U14434 (N_14434,N_11984,N_11376);
xor U14435 (N_14435,N_11394,N_11413);
xor U14436 (N_14436,N_11758,N_11074);
and U14437 (N_14437,N_9549,N_10501);
or U14438 (N_14438,N_12052,N_11190);
xor U14439 (N_14439,N_12117,N_11116);
and U14440 (N_14440,N_12022,N_11085);
or U14441 (N_14441,N_9915,N_10597);
or U14442 (N_14442,N_11306,N_10217);
xor U14443 (N_14443,N_9714,N_11636);
xnor U14444 (N_14444,N_10110,N_11329);
or U14445 (N_14445,N_12316,N_11685);
nand U14446 (N_14446,N_10105,N_10007);
or U14447 (N_14447,N_12232,N_9478);
or U14448 (N_14448,N_11485,N_9437);
nand U14449 (N_14449,N_11856,N_10567);
nand U14450 (N_14450,N_12190,N_11703);
nor U14451 (N_14451,N_9918,N_11686);
nand U14452 (N_14452,N_11309,N_9976);
or U14453 (N_14453,N_9947,N_11680);
or U14454 (N_14454,N_12273,N_11712);
or U14455 (N_14455,N_11289,N_12033);
nand U14456 (N_14456,N_10946,N_9876);
nor U14457 (N_14457,N_10690,N_11377);
nand U14458 (N_14458,N_12067,N_11966);
nand U14459 (N_14459,N_10538,N_9854);
or U14460 (N_14460,N_9967,N_12209);
or U14461 (N_14461,N_10495,N_11379);
xor U14462 (N_14462,N_12207,N_12367);
xnor U14463 (N_14463,N_9759,N_11579);
and U14464 (N_14464,N_12128,N_11879);
or U14465 (N_14465,N_10794,N_9774);
xor U14466 (N_14466,N_11688,N_11081);
nand U14467 (N_14467,N_10532,N_9688);
nor U14468 (N_14468,N_11702,N_10728);
nor U14469 (N_14469,N_10281,N_10173);
nor U14470 (N_14470,N_11557,N_11754);
nor U14471 (N_14471,N_11313,N_11387);
or U14472 (N_14472,N_10484,N_12127);
or U14473 (N_14473,N_11377,N_10730);
nor U14474 (N_14474,N_11687,N_12095);
and U14475 (N_14475,N_11152,N_9931);
xor U14476 (N_14476,N_11821,N_10084);
nand U14477 (N_14477,N_12470,N_11562);
nand U14478 (N_14478,N_10713,N_11597);
and U14479 (N_14479,N_12496,N_11580);
xnor U14480 (N_14480,N_11876,N_9534);
or U14481 (N_14481,N_10567,N_12420);
nand U14482 (N_14482,N_9677,N_9885);
and U14483 (N_14483,N_11445,N_9472);
and U14484 (N_14484,N_9385,N_11455);
nand U14485 (N_14485,N_9492,N_11366);
xnor U14486 (N_14486,N_12456,N_10813);
and U14487 (N_14487,N_11486,N_9999);
xnor U14488 (N_14488,N_9562,N_10037);
xor U14489 (N_14489,N_11747,N_9810);
and U14490 (N_14490,N_11783,N_11206);
nor U14491 (N_14491,N_11971,N_9687);
or U14492 (N_14492,N_11203,N_11715);
xor U14493 (N_14493,N_11704,N_9488);
or U14494 (N_14494,N_12082,N_11238);
and U14495 (N_14495,N_10221,N_11603);
nand U14496 (N_14496,N_11402,N_10431);
nand U14497 (N_14497,N_11590,N_11313);
nor U14498 (N_14498,N_10857,N_9566);
nand U14499 (N_14499,N_9751,N_11684);
xnor U14500 (N_14500,N_12113,N_12093);
xor U14501 (N_14501,N_11482,N_12095);
xnor U14502 (N_14502,N_10033,N_10315);
nor U14503 (N_14503,N_12183,N_10228);
xor U14504 (N_14504,N_12032,N_10002);
or U14505 (N_14505,N_10665,N_12469);
or U14506 (N_14506,N_10322,N_9709);
xor U14507 (N_14507,N_11872,N_10967);
nand U14508 (N_14508,N_11262,N_10532);
and U14509 (N_14509,N_12484,N_10746);
or U14510 (N_14510,N_10521,N_10711);
nand U14511 (N_14511,N_10613,N_10085);
or U14512 (N_14512,N_11738,N_11928);
and U14513 (N_14513,N_9414,N_11912);
or U14514 (N_14514,N_11441,N_11491);
and U14515 (N_14515,N_11097,N_9482);
or U14516 (N_14516,N_9847,N_10693);
nor U14517 (N_14517,N_11271,N_10376);
or U14518 (N_14518,N_11863,N_9658);
xnor U14519 (N_14519,N_10920,N_10217);
xnor U14520 (N_14520,N_12488,N_11200);
nand U14521 (N_14521,N_11345,N_11767);
and U14522 (N_14522,N_11248,N_12366);
xnor U14523 (N_14523,N_11545,N_11210);
and U14524 (N_14524,N_11508,N_11666);
nand U14525 (N_14525,N_10629,N_12408);
or U14526 (N_14526,N_9770,N_10747);
xnor U14527 (N_14527,N_9972,N_9765);
xnor U14528 (N_14528,N_10675,N_9723);
and U14529 (N_14529,N_11992,N_11931);
nand U14530 (N_14530,N_10299,N_11994);
and U14531 (N_14531,N_12175,N_10770);
or U14532 (N_14532,N_9475,N_9675);
nor U14533 (N_14533,N_11954,N_12125);
xnor U14534 (N_14534,N_12480,N_10984);
xnor U14535 (N_14535,N_12112,N_12188);
nand U14536 (N_14536,N_10462,N_11397);
xor U14537 (N_14537,N_9616,N_10594);
or U14538 (N_14538,N_11132,N_9896);
or U14539 (N_14539,N_10068,N_12277);
xor U14540 (N_14540,N_9761,N_11888);
or U14541 (N_14541,N_10869,N_11067);
or U14542 (N_14542,N_10006,N_10941);
nand U14543 (N_14543,N_12431,N_9440);
and U14544 (N_14544,N_11861,N_10245);
xor U14545 (N_14545,N_11498,N_11446);
nor U14546 (N_14546,N_9550,N_10929);
nand U14547 (N_14547,N_9776,N_11775);
nor U14548 (N_14548,N_11715,N_11978);
nand U14549 (N_14549,N_12126,N_11280);
and U14550 (N_14550,N_10302,N_12416);
xor U14551 (N_14551,N_9708,N_10585);
nor U14552 (N_14552,N_12474,N_11972);
xnor U14553 (N_14553,N_9563,N_9434);
nor U14554 (N_14554,N_10364,N_9753);
nand U14555 (N_14555,N_10444,N_11531);
and U14556 (N_14556,N_12317,N_12400);
nor U14557 (N_14557,N_12183,N_11975);
and U14558 (N_14558,N_10772,N_12366);
xor U14559 (N_14559,N_11591,N_12078);
nand U14560 (N_14560,N_10643,N_12299);
xor U14561 (N_14561,N_9878,N_10473);
nand U14562 (N_14562,N_11878,N_12444);
nor U14563 (N_14563,N_12289,N_11998);
or U14564 (N_14564,N_10937,N_9891);
xnor U14565 (N_14565,N_11275,N_9972);
nand U14566 (N_14566,N_10313,N_10399);
xnor U14567 (N_14567,N_11725,N_11075);
or U14568 (N_14568,N_11056,N_12149);
and U14569 (N_14569,N_12246,N_10690);
nand U14570 (N_14570,N_12230,N_12228);
nor U14571 (N_14571,N_10489,N_12082);
nand U14572 (N_14572,N_10419,N_11175);
or U14573 (N_14573,N_9737,N_12349);
xnor U14574 (N_14574,N_11126,N_11630);
nor U14575 (N_14575,N_11462,N_10074);
and U14576 (N_14576,N_9784,N_12288);
and U14577 (N_14577,N_12037,N_10014);
or U14578 (N_14578,N_9750,N_9747);
and U14579 (N_14579,N_12269,N_11673);
and U14580 (N_14580,N_10392,N_12375);
or U14581 (N_14581,N_11956,N_9507);
xor U14582 (N_14582,N_11499,N_12103);
or U14583 (N_14583,N_11027,N_12243);
nand U14584 (N_14584,N_9447,N_10192);
or U14585 (N_14585,N_12271,N_12253);
nand U14586 (N_14586,N_9557,N_12424);
xor U14587 (N_14587,N_10789,N_11865);
or U14588 (N_14588,N_11040,N_11245);
or U14589 (N_14589,N_9882,N_12324);
nor U14590 (N_14590,N_11424,N_10215);
nor U14591 (N_14591,N_12230,N_10086);
nand U14592 (N_14592,N_9504,N_11244);
or U14593 (N_14593,N_9709,N_11389);
xnor U14594 (N_14594,N_11671,N_10065);
nor U14595 (N_14595,N_11194,N_12194);
or U14596 (N_14596,N_9541,N_10944);
or U14597 (N_14597,N_10068,N_11748);
xor U14598 (N_14598,N_11007,N_10883);
nor U14599 (N_14599,N_11127,N_10730);
or U14600 (N_14600,N_10098,N_10284);
or U14601 (N_14601,N_11013,N_11938);
nor U14602 (N_14602,N_9500,N_9597);
nor U14603 (N_14603,N_11616,N_11408);
and U14604 (N_14604,N_9873,N_12348);
nand U14605 (N_14605,N_11784,N_11908);
and U14606 (N_14606,N_11821,N_9870);
xnor U14607 (N_14607,N_9758,N_11566);
or U14608 (N_14608,N_10173,N_10388);
or U14609 (N_14609,N_9656,N_11445);
nand U14610 (N_14610,N_10659,N_10044);
nor U14611 (N_14611,N_10655,N_12306);
and U14612 (N_14612,N_11110,N_11746);
nand U14613 (N_14613,N_10717,N_10425);
nor U14614 (N_14614,N_10176,N_11498);
xor U14615 (N_14615,N_12437,N_9905);
xor U14616 (N_14616,N_12002,N_12187);
xor U14617 (N_14617,N_9632,N_9953);
or U14618 (N_14618,N_9483,N_10922);
nor U14619 (N_14619,N_12275,N_10045);
xor U14620 (N_14620,N_9912,N_11795);
nand U14621 (N_14621,N_10677,N_10182);
nand U14622 (N_14622,N_9645,N_11589);
xnor U14623 (N_14623,N_10487,N_11151);
xnor U14624 (N_14624,N_9958,N_12370);
nor U14625 (N_14625,N_10697,N_12105);
xnor U14626 (N_14626,N_9690,N_10794);
nor U14627 (N_14627,N_11311,N_10475);
and U14628 (N_14628,N_10010,N_9401);
and U14629 (N_14629,N_12380,N_11526);
or U14630 (N_14630,N_12132,N_9841);
or U14631 (N_14631,N_11626,N_11957);
nor U14632 (N_14632,N_11606,N_10182);
or U14633 (N_14633,N_11354,N_10911);
xor U14634 (N_14634,N_9525,N_10135);
nand U14635 (N_14635,N_10898,N_10232);
xnor U14636 (N_14636,N_10739,N_10750);
nor U14637 (N_14637,N_9875,N_9474);
or U14638 (N_14638,N_11273,N_11380);
xor U14639 (N_14639,N_11494,N_12335);
nand U14640 (N_14640,N_12430,N_10880);
and U14641 (N_14641,N_11844,N_11339);
and U14642 (N_14642,N_11201,N_10975);
nand U14643 (N_14643,N_10763,N_11189);
nand U14644 (N_14644,N_12446,N_12422);
xnor U14645 (N_14645,N_10045,N_9487);
or U14646 (N_14646,N_10687,N_11197);
nand U14647 (N_14647,N_10251,N_11484);
or U14648 (N_14648,N_10660,N_10701);
or U14649 (N_14649,N_12438,N_9799);
and U14650 (N_14650,N_10408,N_11714);
nand U14651 (N_14651,N_12424,N_11056);
nor U14652 (N_14652,N_11444,N_10425);
xnor U14653 (N_14653,N_10797,N_11857);
xnor U14654 (N_14654,N_9676,N_10463);
xnor U14655 (N_14655,N_9394,N_9731);
nor U14656 (N_14656,N_11068,N_10091);
or U14657 (N_14657,N_12046,N_10794);
xor U14658 (N_14658,N_9826,N_11409);
nand U14659 (N_14659,N_10767,N_10673);
or U14660 (N_14660,N_10427,N_12216);
xnor U14661 (N_14661,N_11552,N_10747);
or U14662 (N_14662,N_10458,N_12308);
nor U14663 (N_14663,N_9689,N_9957);
and U14664 (N_14664,N_10962,N_12028);
and U14665 (N_14665,N_12231,N_10688);
xor U14666 (N_14666,N_10306,N_11950);
nor U14667 (N_14667,N_10685,N_11502);
xor U14668 (N_14668,N_10537,N_11086);
xor U14669 (N_14669,N_9924,N_12307);
or U14670 (N_14670,N_11096,N_10117);
and U14671 (N_14671,N_10582,N_10621);
xor U14672 (N_14672,N_11952,N_11720);
nand U14673 (N_14673,N_11586,N_11268);
or U14674 (N_14674,N_10656,N_12200);
xnor U14675 (N_14675,N_11987,N_10317);
and U14676 (N_14676,N_11756,N_11472);
xnor U14677 (N_14677,N_11402,N_12422);
nand U14678 (N_14678,N_11890,N_10414);
nor U14679 (N_14679,N_10871,N_10033);
or U14680 (N_14680,N_11827,N_12234);
or U14681 (N_14681,N_12221,N_12414);
and U14682 (N_14682,N_9479,N_10025);
xor U14683 (N_14683,N_10302,N_9722);
or U14684 (N_14684,N_10350,N_9539);
and U14685 (N_14685,N_11144,N_11884);
xnor U14686 (N_14686,N_12480,N_10731);
nand U14687 (N_14687,N_9401,N_10647);
or U14688 (N_14688,N_10680,N_10698);
and U14689 (N_14689,N_10151,N_10133);
nor U14690 (N_14690,N_11702,N_10590);
and U14691 (N_14691,N_11823,N_12206);
or U14692 (N_14692,N_10685,N_11774);
and U14693 (N_14693,N_9401,N_10586);
nand U14694 (N_14694,N_10448,N_9764);
or U14695 (N_14695,N_10498,N_9802);
xnor U14696 (N_14696,N_11599,N_9834);
and U14697 (N_14697,N_9765,N_10593);
and U14698 (N_14698,N_12329,N_9390);
xor U14699 (N_14699,N_10952,N_11811);
nand U14700 (N_14700,N_9983,N_9979);
and U14701 (N_14701,N_9794,N_10001);
nand U14702 (N_14702,N_9465,N_12434);
or U14703 (N_14703,N_10563,N_12303);
and U14704 (N_14704,N_9964,N_9834);
nand U14705 (N_14705,N_11102,N_11908);
nand U14706 (N_14706,N_10381,N_11295);
and U14707 (N_14707,N_9904,N_9377);
or U14708 (N_14708,N_10378,N_10858);
or U14709 (N_14709,N_10542,N_9908);
and U14710 (N_14710,N_10869,N_12311);
or U14711 (N_14711,N_9633,N_11205);
xnor U14712 (N_14712,N_10225,N_10233);
nand U14713 (N_14713,N_12397,N_12366);
nand U14714 (N_14714,N_10609,N_11258);
and U14715 (N_14715,N_10497,N_11463);
xnor U14716 (N_14716,N_11852,N_11514);
xor U14717 (N_14717,N_10296,N_10104);
and U14718 (N_14718,N_10882,N_10182);
or U14719 (N_14719,N_11648,N_11240);
and U14720 (N_14720,N_11802,N_9873);
nand U14721 (N_14721,N_10283,N_10207);
and U14722 (N_14722,N_10847,N_10988);
nand U14723 (N_14723,N_10093,N_10017);
nand U14724 (N_14724,N_10601,N_11508);
nor U14725 (N_14725,N_11460,N_10703);
nor U14726 (N_14726,N_9704,N_11392);
nand U14727 (N_14727,N_10095,N_10091);
nor U14728 (N_14728,N_10487,N_9848);
xnor U14729 (N_14729,N_10331,N_9826);
xnor U14730 (N_14730,N_11070,N_12245);
nand U14731 (N_14731,N_10844,N_10085);
and U14732 (N_14732,N_9526,N_11696);
nor U14733 (N_14733,N_9779,N_11030);
nor U14734 (N_14734,N_11942,N_9489);
nor U14735 (N_14735,N_11580,N_10048);
xnor U14736 (N_14736,N_11573,N_12044);
or U14737 (N_14737,N_10233,N_10006);
xor U14738 (N_14738,N_10138,N_12266);
and U14739 (N_14739,N_10781,N_12171);
nor U14740 (N_14740,N_11090,N_10764);
xnor U14741 (N_14741,N_9870,N_11401);
and U14742 (N_14742,N_11141,N_11904);
nor U14743 (N_14743,N_10948,N_11281);
nand U14744 (N_14744,N_9379,N_11510);
or U14745 (N_14745,N_10109,N_11631);
nor U14746 (N_14746,N_11158,N_12335);
xor U14747 (N_14747,N_11475,N_10485);
nor U14748 (N_14748,N_11167,N_11009);
xor U14749 (N_14749,N_9428,N_10389);
nand U14750 (N_14750,N_10946,N_10035);
nand U14751 (N_14751,N_10049,N_12375);
xor U14752 (N_14752,N_9447,N_10743);
or U14753 (N_14753,N_11820,N_11841);
nor U14754 (N_14754,N_9879,N_11945);
or U14755 (N_14755,N_10796,N_11037);
or U14756 (N_14756,N_9636,N_10116);
xnor U14757 (N_14757,N_10339,N_11255);
nor U14758 (N_14758,N_9685,N_9914);
xnor U14759 (N_14759,N_10787,N_11246);
xor U14760 (N_14760,N_11474,N_10165);
and U14761 (N_14761,N_10947,N_10511);
and U14762 (N_14762,N_9554,N_12202);
nor U14763 (N_14763,N_11830,N_10822);
nand U14764 (N_14764,N_9714,N_11873);
xor U14765 (N_14765,N_10467,N_12256);
and U14766 (N_14766,N_10572,N_10500);
nor U14767 (N_14767,N_11689,N_10481);
xor U14768 (N_14768,N_9482,N_11804);
nor U14769 (N_14769,N_10844,N_12006);
or U14770 (N_14770,N_10813,N_10893);
and U14771 (N_14771,N_11454,N_10623);
nand U14772 (N_14772,N_9865,N_11131);
nand U14773 (N_14773,N_11719,N_10120);
or U14774 (N_14774,N_9927,N_11266);
xnor U14775 (N_14775,N_11582,N_10330);
nand U14776 (N_14776,N_9765,N_9646);
nand U14777 (N_14777,N_11475,N_11922);
or U14778 (N_14778,N_10439,N_11464);
xnor U14779 (N_14779,N_10312,N_10220);
nand U14780 (N_14780,N_11525,N_9532);
nand U14781 (N_14781,N_10349,N_10250);
xnor U14782 (N_14782,N_9690,N_12220);
xor U14783 (N_14783,N_10352,N_11827);
xnor U14784 (N_14784,N_9963,N_12156);
nor U14785 (N_14785,N_11180,N_10781);
xnor U14786 (N_14786,N_11372,N_11864);
xnor U14787 (N_14787,N_9870,N_10282);
or U14788 (N_14788,N_9422,N_11370);
nand U14789 (N_14789,N_10110,N_12118);
and U14790 (N_14790,N_9708,N_11132);
and U14791 (N_14791,N_12144,N_10679);
nand U14792 (N_14792,N_9760,N_12335);
or U14793 (N_14793,N_10706,N_10145);
nand U14794 (N_14794,N_12188,N_10864);
and U14795 (N_14795,N_9916,N_12206);
and U14796 (N_14796,N_9865,N_11828);
xor U14797 (N_14797,N_10759,N_10338);
and U14798 (N_14798,N_10065,N_11498);
and U14799 (N_14799,N_10632,N_10912);
nand U14800 (N_14800,N_10436,N_9731);
nand U14801 (N_14801,N_9872,N_10865);
and U14802 (N_14802,N_10712,N_10105);
xor U14803 (N_14803,N_11174,N_10151);
and U14804 (N_14804,N_11585,N_9954);
and U14805 (N_14805,N_10862,N_11116);
nand U14806 (N_14806,N_11833,N_11201);
nand U14807 (N_14807,N_11786,N_12193);
nand U14808 (N_14808,N_11611,N_9522);
nor U14809 (N_14809,N_10113,N_12348);
and U14810 (N_14810,N_11470,N_12128);
and U14811 (N_14811,N_12278,N_11612);
nand U14812 (N_14812,N_12076,N_10754);
and U14813 (N_14813,N_10779,N_11066);
or U14814 (N_14814,N_11852,N_10160);
xnor U14815 (N_14815,N_11702,N_11190);
nor U14816 (N_14816,N_9380,N_11289);
or U14817 (N_14817,N_11394,N_11935);
nor U14818 (N_14818,N_10912,N_11260);
or U14819 (N_14819,N_9467,N_10036);
or U14820 (N_14820,N_10784,N_9724);
and U14821 (N_14821,N_11031,N_10721);
or U14822 (N_14822,N_10169,N_11374);
and U14823 (N_14823,N_12379,N_10460);
nand U14824 (N_14824,N_9669,N_10606);
xor U14825 (N_14825,N_9660,N_12482);
nand U14826 (N_14826,N_10170,N_12156);
nor U14827 (N_14827,N_9605,N_9573);
or U14828 (N_14828,N_9870,N_12138);
nand U14829 (N_14829,N_10914,N_10473);
or U14830 (N_14830,N_11270,N_11693);
or U14831 (N_14831,N_11276,N_12122);
nand U14832 (N_14832,N_11456,N_9805);
xnor U14833 (N_14833,N_12180,N_10166);
xnor U14834 (N_14834,N_10081,N_12298);
and U14835 (N_14835,N_12209,N_10677);
or U14836 (N_14836,N_11494,N_10461);
xor U14837 (N_14837,N_11425,N_9410);
xor U14838 (N_14838,N_10013,N_10633);
nand U14839 (N_14839,N_10042,N_9431);
nor U14840 (N_14840,N_11574,N_11079);
and U14841 (N_14841,N_11423,N_10601);
nor U14842 (N_14842,N_9568,N_9786);
nor U14843 (N_14843,N_11382,N_10253);
and U14844 (N_14844,N_9634,N_10224);
nand U14845 (N_14845,N_9601,N_12085);
xor U14846 (N_14846,N_12286,N_11895);
xor U14847 (N_14847,N_11234,N_10291);
xnor U14848 (N_14848,N_10643,N_12315);
and U14849 (N_14849,N_11335,N_10505);
and U14850 (N_14850,N_9515,N_11416);
or U14851 (N_14851,N_10190,N_12153);
nor U14852 (N_14852,N_12014,N_10410);
nand U14853 (N_14853,N_10801,N_10694);
nand U14854 (N_14854,N_10162,N_11647);
and U14855 (N_14855,N_11612,N_9859);
xnor U14856 (N_14856,N_10247,N_12435);
xor U14857 (N_14857,N_12428,N_10522);
or U14858 (N_14858,N_12419,N_9832);
nand U14859 (N_14859,N_9786,N_12362);
nor U14860 (N_14860,N_10917,N_12299);
xor U14861 (N_14861,N_11398,N_12071);
nor U14862 (N_14862,N_9536,N_12388);
nand U14863 (N_14863,N_9645,N_10413);
xnor U14864 (N_14864,N_12213,N_11480);
and U14865 (N_14865,N_11729,N_10995);
nand U14866 (N_14866,N_9705,N_11449);
xnor U14867 (N_14867,N_11269,N_11110);
or U14868 (N_14868,N_10397,N_11137);
nand U14869 (N_14869,N_9794,N_9908);
nor U14870 (N_14870,N_11608,N_11575);
nand U14871 (N_14871,N_11570,N_11441);
or U14872 (N_14872,N_10923,N_12066);
nor U14873 (N_14873,N_10633,N_11640);
xor U14874 (N_14874,N_10147,N_10971);
nand U14875 (N_14875,N_9730,N_10614);
nor U14876 (N_14876,N_12218,N_11162);
and U14877 (N_14877,N_11607,N_11240);
nor U14878 (N_14878,N_12297,N_12355);
or U14879 (N_14879,N_10554,N_11673);
nand U14880 (N_14880,N_11926,N_11859);
or U14881 (N_14881,N_9509,N_12265);
and U14882 (N_14882,N_12104,N_11756);
nor U14883 (N_14883,N_12147,N_9855);
nand U14884 (N_14884,N_12235,N_11125);
or U14885 (N_14885,N_9564,N_11777);
or U14886 (N_14886,N_11979,N_11917);
or U14887 (N_14887,N_12153,N_12351);
or U14888 (N_14888,N_9823,N_9692);
nor U14889 (N_14889,N_11815,N_10727);
xnor U14890 (N_14890,N_10155,N_9783);
xor U14891 (N_14891,N_10968,N_11889);
xnor U14892 (N_14892,N_9958,N_11423);
xor U14893 (N_14893,N_12151,N_12188);
nor U14894 (N_14894,N_10992,N_11458);
nand U14895 (N_14895,N_10935,N_11237);
xor U14896 (N_14896,N_10616,N_9833);
or U14897 (N_14897,N_9528,N_10736);
or U14898 (N_14898,N_12348,N_9960);
nor U14899 (N_14899,N_12266,N_9598);
or U14900 (N_14900,N_10723,N_12333);
and U14901 (N_14901,N_10640,N_10734);
nor U14902 (N_14902,N_10500,N_10147);
nor U14903 (N_14903,N_12320,N_10009);
xnor U14904 (N_14904,N_10988,N_11682);
or U14905 (N_14905,N_10217,N_10773);
xnor U14906 (N_14906,N_9401,N_9475);
xnor U14907 (N_14907,N_9565,N_12335);
nor U14908 (N_14908,N_12277,N_11518);
and U14909 (N_14909,N_10873,N_11322);
nor U14910 (N_14910,N_9412,N_12312);
or U14911 (N_14911,N_12285,N_11043);
or U14912 (N_14912,N_12455,N_11863);
nand U14913 (N_14913,N_10146,N_10820);
or U14914 (N_14914,N_12420,N_10469);
xnor U14915 (N_14915,N_11555,N_10541);
xor U14916 (N_14916,N_10003,N_9521);
xnor U14917 (N_14917,N_10854,N_11332);
and U14918 (N_14918,N_9707,N_10322);
xor U14919 (N_14919,N_11049,N_10592);
xnor U14920 (N_14920,N_11743,N_9412);
xor U14921 (N_14921,N_11459,N_10186);
nand U14922 (N_14922,N_9449,N_11752);
xor U14923 (N_14923,N_9582,N_10710);
nand U14924 (N_14924,N_10151,N_12156);
nor U14925 (N_14925,N_10617,N_11550);
and U14926 (N_14926,N_10640,N_11634);
nor U14927 (N_14927,N_10786,N_10014);
or U14928 (N_14928,N_12347,N_9956);
nand U14929 (N_14929,N_9439,N_9948);
nand U14930 (N_14930,N_10204,N_9789);
xor U14931 (N_14931,N_9421,N_11382);
xor U14932 (N_14932,N_10149,N_9705);
and U14933 (N_14933,N_9444,N_10802);
and U14934 (N_14934,N_10615,N_11640);
and U14935 (N_14935,N_9898,N_12369);
and U14936 (N_14936,N_9560,N_11875);
and U14937 (N_14937,N_10035,N_10788);
and U14938 (N_14938,N_11040,N_12042);
and U14939 (N_14939,N_9520,N_10335);
and U14940 (N_14940,N_11954,N_9528);
nand U14941 (N_14941,N_10752,N_11788);
nand U14942 (N_14942,N_9901,N_11856);
nor U14943 (N_14943,N_10114,N_10327);
nor U14944 (N_14944,N_11310,N_9594);
xor U14945 (N_14945,N_9910,N_12043);
nor U14946 (N_14946,N_10512,N_10205);
and U14947 (N_14947,N_11905,N_11508);
nor U14948 (N_14948,N_12151,N_12495);
xor U14949 (N_14949,N_10816,N_10341);
nand U14950 (N_14950,N_11503,N_10709);
or U14951 (N_14951,N_12325,N_10763);
or U14952 (N_14952,N_12128,N_10676);
or U14953 (N_14953,N_9769,N_10364);
or U14954 (N_14954,N_10143,N_9913);
or U14955 (N_14955,N_11827,N_10517);
nand U14956 (N_14956,N_10426,N_11683);
nor U14957 (N_14957,N_11677,N_9622);
xnor U14958 (N_14958,N_11686,N_11339);
nand U14959 (N_14959,N_10076,N_11920);
or U14960 (N_14960,N_10084,N_12480);
nor U14961 (N_14961,N_10782,N_10900);
and U14962 (N_14962,N_11203,N_10932);
xor U14963 (N_14963,N_10811,N_11317);
and U14964 (N_14964,N_11627,N_10918);
and U14965 (N_14965,N_12108,N_10932);
nor U14966 (N_14966,N_12069,N_12262);
and U14967 (N_14967,N_12304,N_9766);
xnor U14968 (N_14968,N_9926,N_12074);
and U14969 (N_14969,N_9399,N_9598);
xor U14970 (N_14970,N_9999,N_11100);
and U14971 (N_14971,N_9457,N_11943);
xor U14972 (N_14972,N_11152,N_10289);
xnor U14973 (N_14973,N_9509,N_9741);
and U14974 (N_14974,N_10488,N_12037);
and U14975 (N_14975,N_10210,N_11391);
nor U14976 (N_14976,N_11319,N_9398);
nor U14977 (N_14977,N_11785,N_10728);
xnor U14978 (N_14978,N_10127,N_10618);
xor U14979 (N_14979,N_12010,N_10404);
or U14980 (N_14980,N_9454,N_11179);
or U14981 (N_14981,N_11188,N_11135);
nand U14982 (N_14982,N_9726,N_11471);
and U14983 (N_14983,N_12401,N_9379);
and U14984 (N_14984,N_10546,N_9967);
nor U14985 (N_14985,N_11846,N_10230);
xor U14986 (N_14986,N_10255,N_11708);
or U14987 (N_14987,N_10656,N_9973);
xnor U14988 (N_14988,N_11628,N_10934);
and U14989 (N_14989,N_10545,N_12052);
nor U14990 (N_14990,N_11711,N_12189);
nand U14991 (N_14991,N_9828,N_10026);
or U14992 (N_14992,N_12208,N_9648);
and U14993 (N_14993,N_12325,N_9848);
xnor U14994 (N_14994,N_10531,N_12268);
and U14995 (N_14995,N_11654,N_10646);
nand U14996 (N_14996,N_11659,N_10626);
and U14997 (N_14997,N_12366,N_9461);
nand U14998 (N_14998,N_10686,N_10568);
and U14999 (N_14999,N_11602,N_9523);
nand U15000 (N_15000,N_11985,N_10326);
and U15001 (N_15001,N_10136,N_10846);
xnor U15002 (N_15002,N_11179,N_9778);
or U15003 (N_15003,N_9783,N_10842);
nand U15004 (N_15004,N_9844,N_9602);
xnor U15005 (N_15005,N_11373,N_9910);
or U15006 (N_15006,N_12193,N_10039);
nand U15007 (N_15007,N_9906,N_10946);
nor U15008 (N_15008,N_9441,N_12418);
or U15009 (N_15009,N_9835,N_10958);
and U15010 (N_15010,N_11526,N_10999);
or U15011 (N_15011,N_11179,N_10004);
or U15012 (N_15012,N_10189,N_11326);
and U15013 (N_15013,N_11809,N_10439);
and U15014 (N_15014,N_12123,N_10586);
and U15015 (N_15015,N_10620,N_10385);
xnor U15016 (N_15016,N_12233,N_10302);
xnor U15017 (N_15017,N_11199,N_10843);
xnor U15018 (N_15018,N_12405,N_11453);
or U15019 (N_15019,N_11070,N_9648);
or U15020 (N_15020,N_12317,N_11928);
or U15021 (N_15021,N_10352,N_10714);
and U15022 (N_15022,N_11495,N_10027);
xor U15023 (N_15023,N_11056,N_12043);
nand U15024 (N_15024,N_10851,N_12072);
or U15025 (N_15025,N_11140,N_11877);
or U15026 (N_15026,N_10203,N_10588);
nand U15027 (N_15027,N_11287,N_11992);
xor U15028 (N_15028,N_11436,N_12205);
xor U15029 (N_15029,N_11755,N_11863);
nor U15030 (N_15030,N_10058,N_10229);
and U15031 (N_15031,N_9650,N_11245);
xnor U15032 (N_15032,N_9658,N_9930);
nand U15033 (N_15033,N_10841,N_10990);
xor U15034 (N_15034,N_9628,N_11809);
or U15035 (N_15035,N_11693,N_9940);
nor U15036 (N_15036,N_12122,N_10747);
or U15037 (N_15037,N_12124,N_10111);
nor U15038 (N_15038,N_11652,N_10698);
or U15039 (N_15039,N_10671,N_11824);
nor U15040 (N_15040,N_11041,N_11371);
or U15041 (N_15041,N_9443,N_9830);
nand U15042 (N_15042,N_10894,N_11538);
nor U15043 (N_15043,N_10793,N_11626);
nor U15044 (N_15044,N_11212,N_9872);
nand U15045 (N_15045,N_12494,N_9929);
nor U15046 (N_15046,N_11793,N_11063);
xor U15047 (N_15047,N_12021,N_11559);
nor U15048 (N_15048,N_9406,N_10868);
nor U15049 (N_15049,N_10954,N_12374);
xnor U15050 (N_15050,N_10535,N_9609);
nor U15051 (N_15051,N_12176,N_11619);
nor U15052 (N_15052,N_11250,N_9815);
and U15053 (N_15053,N_9635,N_10405);
and U15054 (N_15054,N_11802,N_11774);
nor U15055 (N_15055,N_11452,N_9994);
nor U15056 (N_15056,N_11257,N_10178);
xor U15057 (N_15057,N_10428,N_11202);
and U15058 (N_15058,N_11445,N_10999);
and U15059 (N_15059,N_9900,N_9853);
nor U15060 (N_15060,N_10051,N_11308);
nor U15061 (N_15061,N_11450,N_10120);
xnor U15062 (N_15062,N_12336,N_12145);
or U15063 (N_15063,N_10089,N_10703);
nand U15064 (N_15064,N_12433,N_9403);
and U15065 (N_15065,N_10329,N_9415);
nand U15066 (N_15066,N_10676,N_11963);
nand U15067 (N_15067,N_9910,N_12311);
or U15068 (N_15068,N_9603,N_11134);
or U15069 (N_15069,N_10439,N_11955);
and U15070 (N_15070,N_12314,N_9647);
and U15071 (N_15071,N_12227,N_9642);
and U15072 (N_15072,N_9949,N_9431);
nor U15073 (N_15073,N_11310,N_11842);
xor U15074 (N_15074,N_11636,N_10656);
xor U15075 (N_15075,N_9633,N_10319);
and U15076 (N_15076,N_9736,N_12460);
nor U15077 (N_15077,N_11545,N_11357);
nand U15078 (N_15078,N_9926,N_9989);
or U15079 (N_15079,N_12211,N_12122);
and U15080 (N_15080,N_9600,N_12134);
and U15081 (N_15081,N_9816,N_11596);
nand U15082 (N_15082,N_10939,N_12080);
xnor U15083 (N_15083,N_11011,N_10416);
xor U15084 (N_15084,N_10992,N_11070);
and U15085 (N_15085,N_9794,N_9813);
nor U15086 (N_15086,N_11267,N_11058);
or U15087 (N_15087,N_9843,N_11306);
xor U15088 (N_15088,N_9381,N_9425);
and U15089 (N_15089,N_10864,N_10880);
and U15090 (N_15090,N_11249,N_11319);
xnor U15091 (N_15091,N_12409,N_9545);
or U15092 (N_15092,N_9464,N_10279);
and U15093 (N_15093,N_11543,N_9993);
nor U15094 (N_15094,N_9733,N_12093);
xor U15095 (N_15095,N_10273,N_11239);
or U15096 (N_15096,N_10644,N_12259);
or U15097 (N_15097,N_10150,N_10074);
nor U15098 (N_15098,N_11231,N_11529);
xnor U15099 (N_15099,N_10939,N_12352);
nor U15100 (N_15100,N_11428,N_12447);
or U15101 (N_15101,N_12339,N_11269);
and U15102 (N_15102,N_12441,N_11023);
nor U15103 (N_15103,N_10272,N_12245);
nand U15104 (N_15104,N_10434,N_11999);
nand U15105 (N_15105,N_12326,N_11327);
or U15106 (N_15106,N_12313,N_9943);
or U15107 (N_15107,N_10353,N_11723);
nand U15108 (N_15108,N_11057,N_12125);
nor U15109 (N_15109,N_12405,N_11875);
or U15110 (N_15110,N_12367,N_9422);
xnor U15111 (N_15111,N_10493,N_11424);
or U15112 (N_15112,N_10360,N_10485);
and U15113 (N_15113,N_11240,N_9905);
nor U15114 (N_15114,N_11627,N_10110);
nand U15115 (N_15115,N_12355,N_11453);
or U15116 (N_15116,N_9900,N_9622);
xnor U15117 (N_15117,N_10148,N_10442);
and U15118 (N_15118,N_11565,N_11809);
nor U15119 (N_15119,N_12077,N_9877);
or U15120 (N_15120,N_10391,N_11342);
xnor U15121 (N_15121,N_10142,N_10133);
xnor U15122 (N_15122,N_11234,N_10226);
or U15123 (N_15123,N_12356,N_10204);
nor U15124 (N_15124,N_12283,N_10106);
nor U15125 (N_15125,N_11565,N_9434);
and U15126 (N_15126,N_10337,N_9877);
xnor U15127 (N_15127,N_12043,N_10394);
xor U15128 (N_15128,N_10393,N_11976);
xor U15129 (N_15129,N_10353,N_11548);
nor U15130 (N_15130,N_11587,N_12427);
xnor U15131 (N_15131,N_11508,N_9375);
nor U15132 (N_15132,N_10052,N_10275);
and U15133 (N_15133,N_11083,N_10325);
nor U15134 (N_15134,N_10421,N_11416);
xnor U15135 (N_15135,N_11693,N_10625);
and U15136 (N_15136,N_11968,N_10774);
xnor U15137 (N_15137,N_11272,N_10529);
and U15138 (N_15138,N_12071,N_12355);
xnor U15139 (N_15139,N_11612,N_12256);
xor U15140 (N_15140,N_9956,N_9701);
and U15141 (N_15141,N_11289,N_10415);
xnor U15142 (N_15142,N_11762,N_11687);
nor U15143 (N_15143,N_10203,N_10021);
nand U15144 (N_15144,N_10192,N_11970);
nor U15145 (N_15145,N_12392,N_11939);
nand U15146 (N_15146,N_11672,N_11343);
nor U15147 (N_15147,N_10697,N_11744);
and U15148 (N_15148,N_10359,N_12437);
or U15149 (N_15149,N_12308,N_9971);
nand U15150 (N_15150,N_11193,N_10048);
nand U15151 (N_15151,N_10959,N_11385);
xor U15152 (N_15152,N_11272,N_9454);
nand U15153 (N_15153,N_10337,N_10978);
or U15154 (N_15154,N_10081,N_11184);
and U15155 (N_15155,N_11822,N_9402);
or U15156 (N_15156,N_11244,N_11713);
xor U15157 (N_15157,N_10787,N_9777);
and U15158 (N_15158,N_11857,N_12448);
nand U15159 (N_15159,N_10309,N_10460);
nor U15160 (N_15160,N_9803,N_10967);
or U15161 (N_15161,N_12254,N_11984);
and U15162 (N_15162,N_10909,N_12303);
or U15163 (N_15163,N_11891,N_10222);
or U15164 (N_15164,N_10384,N_10360);
xor U15165 (N_15165,N_10124,N_9694);
and U15166 (N_15166,N_12120,N_10666);
xnor U15167 (N_15167,N_9581,N_10582);
and U15168 (N_15168,N_11799,N_11555);
nand U15169 (N_15169,N_10187,N_11582);
nor U15170 (N_15170,N_11344,N_9813);
xor U15171 (N_15171,N_12417,N_11791);
or U15172 (N_15172,N_12181,N_10005);
or U15173 (N_15173,N_9631,N_9865);
nand U15174 (N_15174,N_12055,N_12238);
or U15175 (N_15175,N_9814,N_11044);
nand U15176 (N_15176,N_11642,N_9611);
nor U15177 (N_15177,N_10176,N_9969);
nor U15178 (N_15178,N_11158,N_9392);
or U15179 (N_15179,N_12266,N_12134);
xor U15180 (N_15180,N_11132,N_9728);
and U15181 (N_15181,N_11401,N_12164);
and U15182 (N_15182,N_10148,N_10460);
or U15183 (N_15183,N_10753,N_11518);
nor U15184 (N_15184,N_10098,N_10151);
nand U15185 (N_15185,N_10515,N_10245);
xnor U15186 (N_15186,N_10459,N_11605);
nor U15187 (N_15187,N_10234,N_11782);
xnor U15188 (N_15188,N_10019,N_10133);
nor U15189 (N_15189,N_11831,N_9380);
nand U15190 (N_15190,N_9640,N_11924);
and U15191 (N_15191,N_11568,N_10135);
xor U15192 (N_15192,N_12006,N_12326);
or U15193 (N_15193,N_10867,N_11593);
and U15194 (N_15194,N_10048,N_11508);
and U15195 (N_15195,N_9878,N_9866);
or U15196 (N_15196,N_9624,N_11396);
nand U15197 (N_15197,N_11422,N_10311);
and U15198 (N_15198,N_9993,N_11732);
and U15199 (N_15199,N_10258,N_11627);
nor U15200 (N_15200,N_9471,N_9752);
or U15201 (N_15201,N_11508,N_10003);
xor U15202 (N_15202,N_12320,N_11182);
xor U15203 (N_15203,N_12210,N_11116);
nand U15204 (N_15204,N_10212,N_12099);
xor U15205 (N_15205,N_9935,N_11387);
and U15206 (N_15206,N_12041,N_12214);
xnor U15207 (N_15207,N_10823,N_10825);
nand U15208 (N_15208,N_9482,N_11466);
nor U15209 (N_15209,N_11130,N_9660);
nand U15210 (N_15210,N_11393,N_10766);
nand U15211 (N_15211,N_9994,N_9401);
nor U15212 (N_15212,N_10608,N_10702);
or U15213 (N_15213,N_11397,N_10795);
nand U15214 (N_15214,N_9844,N_10659);
xor U15215 (N_15215,N_10570,N_11449);
and U15216 (N_15216,N_9586,N_10655);
or U15217 (N_15217,N_11716,N_11120);
xor U15218 (N_15218,N_10138,N_9935);
xnor U15219 (N_15219,N_11329,N_10474);
and U15220 (N_15220,N_12498,N_9467);
and U15221 (N_15221,N_11890,N_10154);
nor U15222 (N_15222,N_10372,N_11570);
or U15223 (N_15223,N_11776,N_9435);
nor U15224 (N_15224,N_10611,N_9922);
xnor U15225 (N_15225,N_10389,N_12370);
xor U15226 (N_15226,N_11630,N_12206);
or U15227 (N_15227,N_12330,N_10373);
and U15228 (N_15228,N_10708,N_10329);
or U15229 (N_15229,N_9507,N_10962);
or U15230 (N_15230,N_11153,N_10676);
xor U15231 (N_15231,N_10006,N_10497);
xor U15232 (N_15232,N_10431,N_10377);
xor U15233 (N_15233,N_10486,N_11189);
xor U15234 (N_15234,N_9803,N_11721);
xor U15235 (N_15235,N_10109,N_10046);
xnor U15236 (N_15236,N_11372,N_10463);
nor U15237 (N_15237,N_10632,N_12232);
or U15238 (N_15238,N_12425,N_11560);
nand U15239 (N_15239,N_12390,N_10970);
xor U15240 (N_15240,N_10504,N_12204);
xor U15241 (N_15241,N_11633,N_10300);
nand U15242 (N_15242,N_12427,N_12247);
xnor U15243 (N_15243,N_11580,N_9551);
nor U15244 (N_15244,N_10557,N_11150);
nor U15245 (N_15245,N_11633,N_10032);
xor U15246 (N_15246,N_10016,N_9693);
or U15247 (N_15247,N_11254,N_9925);
xnor U15248 (N_15248,N_11231,N_12349);
nand U15249 (N_15249,N_11372,N_10094);
xor U15250 (N_15250,N_10376,N_10807);
xnor U15251 (N_15251,N_9709,N_10798);
nand U15252 (N_15252,N_10929,N_11454);
and U15253 (N_15253,N_10401,N_12440);
nor U15254 (N_15254,N_9805,N_11933);
and U15255 (N_15255,N_12146,N_11965);
xnor U15256 (N_15256,N_11141,N_12024);
and U15257 (N_15257,N_12228,N_9587);
nand U15258 (N_15258,N_11718,N_12364);
and U15259 (N_15259,N_9632,N_10289);
and U15260 (N_15260,N_12355,N_11682);
nor U15261 (N_15261,N_12198,N_10958);
xor U15262 (N_15262,N_9421,N_9402);
nor U15263 (N_15263,N_10232,N_9764);
nor U15264 (N_15264,N_11469,N_11034);
or U15265 (N_15265,N_10894,N_9395);
nand U15266 (N_15266,N_11384,N_11470);
nand U15267 (N_15267,N_11172,N_10907);
nor U15268 (N_15268,N_10924,N_11957);
xor U15269 (N_15269,N_9937,N_11577);
nor U15270 (N_15270,N_10664,N_10333);
and U15271 (N_15271,N_11899,N_10126);
or U15272 (N_15272,N_11931,N_12042);
or U15273 (N_15273,N_11028,N_9703);
or U15274 (N_15274,N_10788,N_11148);
or U15275 (N_15275,N_11245,N_12176);
and U15276 (N_15276,N_11063,N_9706);
nand U15277 (N_15277,N_10188,N_9688);
nand U15278 (N_15278,N_10830,N_11799);
or U15279 (N_15279,N_12274,N_10786);
xor U15280 (N_15280,N_10644,N_11928);
or U15281 (N_15281,N_11930,N_9611);
or U15282 (N_15282,N_10992,N_10463);
or U15283 (N_15283,N_11493,N_9462);
xor U15284 (N_15284,N_12412,N_10635);
and U15285 (N_15285,N_9794,N_12104);
nand U15286 (N_15286,N_11421,N_11490);
nor U15287 (N_15287,N_9899,N_9937);
or U15288 (N_15288,N_11779,N_12009);
xor U15289 (N_15289,N_11426,N_9920);
nor U15290 (N_15290,N_11594,N_10175);
xnor U15291 (N_15291,N_9730,N_10525);
or U15292 (N_15292,N_9773,N_11576);
and U15293 (N_15293,N_11327,N_11251);
and U15294 (N_15294,N_9902,N_12422);
xor U15295 (N_15295,N_11129,N_10405);
nor U15296 (N_15296,N_12388,N_10163);
nor U15297 (N_15297,N_11517,N_9506);
nand U15298 (N_15298,N_12360,N_11153);
and U15299 (N_15299,N_10689,N_11600);
or U15300 (N_15300,N_10060,N_11714);
xnor U15301 (N_15301,N_11339,N_10805);
xor U15302 (N_15302,N_11015,N_11418);
and U15303 (N_15303,N_11136,N_10754);
xnor U15304 (N_15304,N_9795,N_9833);
nor U15305 (N_15305,N_12480,N_12105);
or U15306 (N_15306,N_11530,N_10330);
and U15307 (N_15307,N_11098,N_11333);
or U15308 (N_15308,N_11143,N_11794);
and U15309 (N_15309,N_9826,N_9569);
nor U15310 (N_15310,N_9508,N_10789);
nand U15311 (N_15311,N_10134,N_10609);
or U15312 (N_15312,N_12197,N_11430);
nand U15313 (N_15313,N_11933,N_9739);
and U15314 (N_15314,N_11546,N_11855);
xor U15315 (N_15315,N_10945,N_12100);
xnor U15316 (N_15316,N_10097,N_9948);
xor U15317 (N_15317,N_12264,N_11563);
and U15318 (N_15318,N_11639,N_12498);
and U15319 (N_15319,N_11950,N_9886);
nand U15320 (N_15320,N_11188,N_10403);
xnor U15321 (N_15321,N_12086,N_11528);
xor U15322 (N_15322,N_12232,N_10130);
or U15323 (N_15323,N_11776,N_10403);
xnor U15324 (N_15324,N_11970,N_9604);
nor U15325 (N_15325,N_11739,N_11180);
nor U15326 (N_15326,N_11399,N_10344);
or U15327 (N_15327,N_11506,N_11583);
nor U15328 (N_15328,N_10183,N_10334);
and U15329 (N_15329,N_10174,N_10431);
nand U15330 (N_15330,N_11355,N_11081);
and U15331 (N_15331,N_10199,N_10035);
nor U15332 (N_15332,N_12470,N_9919);
or U15333 (N_15333,N_9781,N_10831);
nand U15334 (N_15334,N_12269,N_10703);
xnor U15335 (N_15335,N_11580,N_9611);
nand U15336 (N_15336,N_10504,N_11054);
xor U15337 (N_15337,N_12316,N_11030);
nor U15338 (N_15338,N_12135,N_10442);
nor U15339 (N_15339,N_9404,N_10293);
nor U15340 (N_15340,N_12495,N_11540);
nand U15341 (N_15341,N_12379,N_10852);
and U15342 (N_15342,N_12324,N_12483);
nor U15343 (N_15343,N_9911,N_12211);
and U15344 (N_15344,N_12465,N_10271);
xor U15345 (N_15345,N_10689,N_11036);
or U15346 (N_15346,N_12028,N_12039);
and U15347 (N_15347,N_11338,N_10197);
nand U15348 (N_15348,N_12292,N_10124);
xnor U15349 (N_15349,N_10253,N_11403);
nand U15350 (N_15350,N_11669,N_11294);
nand U15351 (N_15351,N_11495,N_11929);
xor U15352 (N_15352,N_10822,N_11472);
and U15353 (N_15353,N_12034,N_12268);
or U15354 (N_15354,N_11185,N_9770);
nand U15355 (N_15355,N_10372,N_10220);
nor U15356 (N_15356,N_9880,N_11409);
nor U15357 (N_15357,N_10718,N_11912);
and U15358 (N_15358,N_10823,N_11602);
nor U15359 (N_15359,N_10332,N_11763);
nor U15360 (N_15360,N_12031,N_12054);
or U15361 (N_15361,N_9755,N_10121);
nand U15362 (N_15362,N_10702,N_12497);
nor U15363 (N_15363,N_10913,N_11260);
nor U15364 (N_15364,N_11172,N_12247);
xnor U15365 (N_15365,N_12208,N_9489);
nand U15366 (N_15366,N_11031,N_9659);
nor U15367 (N_15367,N_10883,N_12244);
and U15368 (N_15368,N_10672,N_9536);
and U15369 (N_15369,N_11883,N_12220);
xor U15370 (N_15370,N_9410,N_12324);
and U15371 (N_15371,N_9895,N_9952);
or U15372 (N_15372,N_11916,N_12240);
nand U15373 (N_15373,N_9679,N_10712);
nand U15374 (N_15374,N_10391,N_10684);
and U15375 (N_15375,N_9427,N_12356);
nor U15376 (N_15376,N_10158,N_9425);
nand U15377 (N_15377,N_10088,N_11680);
nand U15378 (N_15378,N_12268,N_12204);
nor U15379 (N_15379,N_10144,N_11421);
nor U15380 (N_15380,N_12487,N_12233);
nor U15381 (N_15381,N_12287,N_12238);
nand U15382 (N_15382,N_12145,N_9464);
nor U15383 (N_15383,N_9412,N_10152);
xnor U15384 (N_15384,N_10932,N_11036);
nor U15385 (N_15385,N_10630,N_11138);
xor U15386 (N_15386,N_12249,N_10278);
xor U15387 (N_15387,N_9469,N_9446);
nor U15388 (N_15388,N_11261,N_12468);
nor U15389 (N_15389,N_11234,N_11508);
nand U15390 (N_15390,N_9851,N_10820);
nor U15391 (N_15391,N_11200,N_9916);
xnor U15392 (N_15392,N_11655,N_11077);
or U15393 (N_15393,N_10476,N_12218);
or U15394 (N_15394,N_10078,N_10670);
or U15395 (N_15395,N_11883,N_10605);
xor U15396 (N_15396,N_9612,N_11854);
and U15397 (N_15397,N_12051,N_11715);
and U15398 (N_15398,N_11718,N_10878);
xnor U15399 (N_15399,N_11337,N_9869);
or U15400 (N_15400,N_9784,N_10616);
nand U15401 (N_15401,N_11804,N_11034);
nor U15402 (N_15402,N_10610,N_12307);
nor U15403 (N_15403,N_9859,N_11770);
or U15404 (N_15404,N_10322,N_10530);
nand U15405 (N_15405,N_10862,N_9393);
nand U15406 (N_15406,N_10780,N_10942);
nand U15407 (N_15407,N_10149,N_10321);
and U15408 (N_15408,N_10116,N_10516);
nand U15409 (N_15409,N_11842,N_10616);
nor U15410 (N_15410,N_11409,N_11966);
nand U15411 (N_15411,N_11842,N_11050);
nand U15412 (N_15412,N_10374,N_10629);
nor U15413 (N_15413,N_11856,N_12470);
nand U15414 (N_15414,N_9536,N_11319);
and U15415 (N_15415,N_12323,N_10915);
nor U15416 (N_15416,N_12207,N_11547);
nand U15417 (N_15417,N_11054,N_11593);
or U15418 (N_15418,N_11580,N_11598);
nand U15419 (N_15419,N_11316,N_11524);
nand U15420 (N_15420,N_11807,N_10248);
or U15421 (N_15421,N_10205,N_9954);
xnor U15422 (N_15422,N_12397,N_12147);
or U15423 (N_15423,N_12329,N_11687);
or U15424 (N_15424,N_11133,N_12373);
nor U15425 (N_15425,N_10426,N_10319);
nand U15426 (N_15426,N_10081,N_12193);
nor U15427 (N_15427,N_10756,N_12394);
nand U15428 (N_15428,N_11325,N_9613);
nor U15429 (N_15429,N_10993,N_11500);
xnor U15430 (N_15430,N_12128,N_11337);
nor U15431 (N_15431,N_11329,N_10517);
xnor U15432 (N_15432,N_9847,N_12477);
nor U15433 (N_15433,N_11916,N_11043);
and U15434 (N_15434,N_10417,N_10168);
nand U15435 (N_15435,N_11583,N_11224);
or U15436 (N_15436,N_12083,N_9513);
nand U15437 (N_15437,N_10450,N_11442);
or U15438 (N_15438,N_10525,N_12331);
and U15439 (N_15439,N_10063,N_10027);
or U15440 (N_15440,N_10383,N_11600);
and U15441 (N_15441,N_11413,N_11503);
nor U15442 (N_15442,N_12322,N_10572);
and U15443 (N_15443,N_10432,N_10710);
and U15444 (N_15444,N_12058,N_11884);
xnor U15445 (N_15445,N_10784,N_11424);
nand U15446 (N_15446,N_12227,N_12163);
or U15447 (N_15447,N_9382,N_9495);
and U15448 (N_15448,N_12480,N_11802);
nand U15449 (N_15449,N_11834,N_10222);
and U15450 (N_15450,N_9635,N_12393);
xnor U15451 (N_15451,N_9956,N_10200);
or U15452 (N_15452,N_11438,N_11504);
or U15453 (N_15453,N_11819,N_11389);
or U15454 (N_15454,N_10303,N_12034);
or U15455 (N_15455,N_11858,N_11638);
or U15456 (N_15456,N_11703,N_10865);
nand U15457 (N_15457,N_10425,N_11698);
nor U15458 (N_15458,N_9708,N_12139);
nand U15459 (N_15459,N_11711,N_11684);
nor U15460 (N_15460,N_10019,N_12238);
or U15461 (N_15461,N_11081,N_11294);
nor U15462 (N_15462,N_10782,N_10713);
or U15463 (N_15463,N_11806,N_9831);
nor U15464 (N_15464,N_10938,N_10826);
xnor U15465 (N_15465,N_11284,N_11614);
nand U15466 (N_15466,N_12163,N_10682);
and U15467 (N_15467,N_10340,N_10487);
or U15468 (N_15468,N_9712,N_12350);
nor U15469 (N_15469,N_11272,N_11658);
xor U15470 (N_15470,N_12289,N_11360);
nand U15471 (N_15471,N_11349,N_11006);
nand U15472 (N_15472,N_11339,N_10811);
xor U15473 (N_15473,N_10511,N_10255);
xor U15474 (N_15474,N_10593,N_12381);
nor U15475 (N_15475,N_12238,N_9454);
and U15476 (N_15476,N_11669,N_11692);
or U15477 (N_15477,N_10667,N_12455);
or U15478 (N_15478,N_10639,N_9527);
xnor U15479 (N_15479,N_12439,N_12295);
and U15480 (N_15480,N_11267,N_11604);
nor U15481 (N_15481,N_12463,N_9888);
or U15482 (N_15482,N_10397,N_11674);
nand U15483 (N_15483,N_10823,N_12166);
and U15484 (N_15484,N_11648,N_11357);
or U15485 (N_15485,N_10543,N_11248);
and U15486 (N_15486,N_11000,N_11014);
nand U15487 (N_15487,N_9407,N_9919);
and U15488 (N_15488,N_11933,N_11926);
nand U15489 (N_15489,N_10694,N_12392);
or U15490 (N_15490,N_10379,N_11653);
or U15491 (N_15491,N_9666,N_11537);
nand U15492 (N_15492,N_12023,N_11177);
and U15493 (N_15493,N_11657,N_11674);
xor U15494 (N_15494,N_11922,N_10381);
or U15495 (N_15495,N_12322,N_11071);
nand U15496 (N_15496,N_10143,N_11350);
or U15497 (N_15497,N_9605,N_12384);
or U15498 (N_15498,N_10557,N_11296);
or U15499 (N_15499,N_10927,N_11125);
nor U15500 (N_15500,N_9619,N_10801);
nand U15501 (N_15501,N_11179,N_12363);
xor U15502 (N_15502,N_9874,N_12430);
nand U15503 (N_15503,N_11253,N_10367);
nor U15504 (N_15504,N_12260,N_12025);
or U15505 (N_15505,N_11859,N_9771);
and U15506 (N_15506,N_10073,N_12299);
nand U15507 (N_15507,N_9516,N_11235);
nor U15508 (N_15508,N_9952,N_9566);
nand U15509 (N_15509,N_11590,N_9970);
nor U15510 (N_15510,N_10645,N_12142);
and U15511 (N_15511,N_9742,N_12491);
and U15512 (N_15512,N_11254,N_10192);
or U15513 (N_15513,N_10280,N_11376);
or U15514 (N_15514,N_12477,N_12304);
nand U15515 (N_15515,N_9858,N_9634);
nor U15516 (N_15516,N_12295,N_9512);
nand U15517 (N_15517,N_11076,N_12177);
nor U15518 (N_15518,N_10955,N_12290);
nor U15519 (N_15519,N_12131,N_10682);
and U15520 (N_15520,N_10164,N_10351);
and U15521 (N_15521,N_10333,N_10931);
nand U15522 (N_15522,N_9922,N_11507);
nand U15523 (N_15523,N_10790,N_10812);
xnor U15524 (N_15524,N_11616,N_11071);
nand U15525 (N_15525,N_11415,N_10412);
nor U15526 (N_15526,N_10406,N_9393);
and U15527 (N_15527,N_11991,N_10016);
nor U15528 (N_15528,N_10506,N_10202);
and U15529 (N_15529,N_10454,N_10494);
xor U15530 (N_15530,N_10973,N_11115);
xor U15531 (N_15531,N_11388,N_11997);
or U15532 (N_15532,N_10363,N_9922);
and U15533 (N_15533,N_9510,N_12469);
and U15534 (N_15534,N_9536,N_10863);
nor U15535 (N_15535,N_11849,N_11604);
and U15536 (N_15536,N_10806,N_10030);
or U15537 (N_15537,N_11396,N_11404);
or U15538 (N_15538,N_11495,N_11371);
nor U15539 (N_15539,N_11815,N_10856);
and U15540 (N_15540,N_11568,N_9614);
xor U15541 (N_15541,N_12327,N_11914);
and U15542 (N_15542,N_10315,N_11837);
xor U15543 (N_15543,N_12249,N_12071);
or U15544 (N_15544,N_11531,N_12139);
or U15545 (N_15545,N_9485,N_9945);
and U15546 (N_15546,N_9684,N_12159);
and U15547 (N_15547,N_9675,N_11288);
and U15548 (N_15548,N_9562,N_10614);
nor U15549 (N_15549,N_12253,N_11779);
and U15550 (N_15550,N_12139,N_12259);
nor U15551 (N_15551,N_12373,N_11998);
or U15552 (N_15552,N_12152,N_11985);
and U15553 (N_15553,N_11942,N_11498);
xnor U15554 (N_15554,N_10636,N_9650);
xor U15555 (N_15555,N_10147,N_9518);
nor U15556 (N_15556,N_12266,N_9816);
nor U15557 (N_15557,N_11297,N_11362);
nand U15558 (N_15558,N_12158,N_10710);
xor U15559 (N_15559,N_12078,N_12437);
xnor U15560 (N_15560,N_9375,N_10424);
xor U15561 (N_15561,N_11099,N_10303);
nand U15562 (N_15562,N_11029,N_10341);
and U15563 (N_15563,N_11184,N_11224);
nor U15564 (N_15564,N_10209,N_10684);
nand U15565 (N_15565,N_9905,N_11868);
nor U15566 (N_15566,N_11119,N_11815);
and U15567 (N_15567,N_11562,N_11285);
nand U15568 (N_15568,N_10276,N_10918);
or U15569 (N_15569,N_10052,N_11806);
xor U15570 (N_15570,N_11745,N_10837);
and U15571 (N_15571,N_12155,N_11167);
and U15572 (N_15572,N_10235,N_10556);
nand U15573 (N_15573,N_12205,N_10674);
xnor U15574 (N_15574,N_10033,N_12436);
and U15575 (N_15575,N_12343,N_10810);
xnor U15576 (N_15576,N_10947,N_9590);
and U15577 (N_15577,N_11112,N_11799);
nand U15578 (N_15578,N_12476,N_11840);
or U15579 (N_15579,N_11704,N_10449);
nand U15580 (N_15580,N_9948,N_11014);
or U15581 (N_15581,N_12280,N_9686);
nand U15582 (N_15582,N_12180,N_10169);
or U15583 (N_15583,N_11024,N_11514);
xor U15584 (N_15584,N_10252,N_11627);
or U15585 (N_15585,N_9639,N_10530);
xor U15586 (N_15586,N_10266,N_10227);
xor U15587 (N_15587,N_11996,N_11596);
or U15588 (N_15588,N_9410,N_11578);
nor U15589 (N_15589,N_9790,N_10706);
or U15590 (N_15590,N_9473,N_11260);
nor U15591 (N_15591,N_9537,N_10431);
nor U15592 (N_15592,N_12303,N_11641);
nand U15593 (N_15593,N_12190,N_12036);
xnor U15594 (N_15594,N_11933,N_12269);
nand U15595 (N_15595,N_11964,N_11898);
nand U15596 (N_15596,N_10154,N_9695);
xor U15597 (N_15597,N_11634,N_11564);
and U15598 (N_15598,N_11768,N_11305);
nor U15599 (N_15599,N_10109,N_12292);
xnor U15600 (N_15600,N_12263,N_12073);
and U15601 (N_15601,N_10985,N_10297);
xor U15602 (N_15602,N_12234,N_10463);
nand U15603 (N_15603,N_9958,N_11861);
or U15604 (N_15604,N_9577,N_10010);
or U15605 (N_15605,N_10538,N_12468);
nor U15606 (N_15606,N_11631,N_10945);
or U15607 (N_15607,N_11265,N_10025);
or U15608 (N_15608,N_11318,N_11841);
or U15609 (N_15609,N_9759,N_11957);
xnor U15610 (N_15610,N_9698,N_11027);
xnor U15611 (N_15611,N_9872,N_10842);
xnor U15612 (N_15612,N_12129,N_10319);
nand U15613 (N_15613,N_10897,N_10795);
nand U15614 (N_15614,N_12149,N_11555);
and U15615 (N_15615,N_9634,N_10040);
nand U15616 (N_15616,N_11015,N_12303);
nand U15617 (N_15617,N_11855,N_11088);
nand U15618 (N_15618,N_9862,N_10183);
xnor U15619 (N_15619,N_9403,N_10618);
or U15620 (N_15620,N_9861,N_11639);
and U15621 (N_15621,N_9913,N_11101);
or U15622 (N_15622,N_11360,N_11661);
nand U15623 (N_15623,N_10735,N_11435);
nand U15624 (N_15624,N_10934,N_10912);
and U15625 (N_15625,N_15051,N_14012);
xor U15626 (N_15626,N_13268,N_15287);
and U15627 (N_15627,N_15313,N_14577);
xor U15628 (N_15628,N_13428,N_12735);
and U15629 (N_15629,N_12754,N_15523);
nor U15630 (N_15630,N_14410,N_12873);
xnor U15631 (N_15631,N_13028,N_14421);
nor U15632 (N_15632,N_12737,N_13102);
or U15633 (N_15633,N_13440,N_14375);
and U15634 (N_15634,N_14814,N_14755);
or U15635 (N_15635,N_14368,N_12609);
and U15636 (N_15636,N_12938,N_14436);
nand U15637 (N_15637,N_12719,N_13622);
nand U15638 (N_15638,N_12631,N_12680);
nand U15639 (N_15639,N_15074,N_15352);
xnor U15640 (N_15640,N_13311,N_13376);
nand U15641 (N_15641,N_15200,N_14936);
or U15642 (N_15642,N_13660,N_15530);
or U15643 (N_15643,N_14294,N_14414);
xor U15644 (N_15644,N_14148,N_13762);
xnor U15645 (N_15645,N_15097,N_12671);
xor U15646 (N_15646,N_13141,N_14205);
and U15647 (N_15647,N_13850,N_13297);
nand U15648 (N_15648,N_13839,N_12545);
xnor U15649 (N_15649,N_13289,N_14056);
nor U15650 (N_15650,N_15138,N_13379);
xnor U15651 (N_15651,N_14550,N_14213);
and U15652 (N_15652,N_14809,N_15435);
nand U15653 (N_15653,N_13121,N_13017);
nand U15654 (N_15654,N_13377,N_14722);
nor U15655 (N_15655,N_14683,N_13306);
nor U15656 (N_15656,N_15285,N_13799);
and U15657 (N_15657,N_12763,N_14861);
xor U15658 (N_15658,N_13555,N_14061);
xor U15659 (N_15659,N_13769,N_14830);
nand U15660 (N_15660,N_13866,N_13795);
and U15661 (N_15661,N_14513,N_15219);
nand U15662 (N_15662,N_14460,N_15562);
xnor U15663 (N_15663,N_12687,N_14155);
nor U15664 (N_15664,N_15465,N_13034);
xor U15665 (N_15665,N_14198,N_13914);
and U15666 (N_15666,N_12562,N_15229);
or U15667 (N_15667,N_14178,N_15373);
nand U15668 (N_15668,N_14200,N_15305);
xnor U15669 (N_15669,N_12862,N_13992);
xnor U15670 (N_15670,N_13919,N_15361);
and U15671 (N_15671,N_13653,N_15568);
nor U15672 (N_15672,N_12667,N_15612);
and U15673 (N_15673,N_14121,N_14542);
and U15674 (N_15674,N_13597,N_13347);
nand U15675 (N_15675,N_14656,N_15316);
and U15676 (N_15676,N_12864,N_13542);
nand U15677 (N_15677,N_15330,N_14299);
and U15678 (N_15678,N_14456,N_12824);
or U15679 (N_15679,N_15593,N_13262);
nor U15680 (N_15680,N_13003,N_14693);
xor U15681 (N_15681,N_15171,N_15077);
or U15682 (N_15682,N_15012,N_14437);
or U15683 (N_15683,N_15588,N_13968);
or U15684 (N_15684,N_13656,N_15036);
or U15685 (N_15685,N_13886,N_12602);
xor U15686 (N_15686,N_14505,N_13265);
and U15687 (N_15687,N_13133,N_12511);
nand U15688 (N_15688,N_15471,N_12663);
or U15689 (N_15689,N_14468,N_14382);
and U15690 (N_15690,N_13537,N_14054);
nor U15691 (N_15691,N_12806,N_12962);
nand U15692 (N_15692,N_15033,N_14063);
nor U15693 (N_15693,N_14699,N_12621);
or U15694 (N_15694,N_13177,N_15223);
and U15695 (N_15695,N_14201,N_14469);
or U15696 (N_15696,N_14122,N_14439);
xor U15697 (N_15697,N_13106,N_12752);
nor U15698 (N_15698,N_14230,N_13420);
nand U15699 (N_15699,N_15600,N_12576);
nand U15700 (N_15700,N_14025,N_13872);
nor U15701 (N_15701,N_12946,N_14029);
or U15702 (N_15702,N_15442,N_14046);
and U15703 (N_15703,N_14268,N_14820);
or U15704 (N_15704,N_15463,N_12733);
nor U15705 (N_15705,N_14831,N_12903);
nand U15706 (N_15706,N_12802,N_15543);
nor U15707 (N_15707,N_13817,N_12986);
or U15708 (N_15708,N_14825,N_15039);
or U15709 (N_15709,N_15151,N_13137);
xnor U15710 (N_15710,N_13517,N_15528);
nand U15711 (N_15711,N_15042,N_15315);
nand U15712 (N_15712,N_13545,N_13745);
nor U15713 (N_15713,N_13549,N_12790);
xnor U15714 (N_15714,N_15495,N_13158);
nor U15715 (N_15715,N_13266,N_15414);
xor U15716 (N_15716,N_15494,N_13867);
nor U15717 (N_15717,N_15355,N_15191);
and U15718 (N_15718,N_13583,N_13337);
nand U15719 (N_15719,N_15337,N_15328);
and U15720 (N_15720,N_14409,N_12693);
xnor U15721 (N_15721,N_15172,N_14694);
nor U15722 (N_15722,N_14625,N_12934);
nand U15723 (N_15723,N_15522,N_12504);
nor U15724 (N_15724,N_14968,N_12894);
and U15725 (N_15725,N_12626,N_12568);
xor U15726 (N_15726,N_12753,N_14775);
nor U15727 (N_15727,N_14765,N_13145);
nor U15728 (N_15728,N_14941,N_15016);
or U15729 (N_15729,N_13305,N_12682);
or U15730 (N_15730,N_15481,N_15620);
and U15731 (N_15731,N_14594,N_15547);
and U15732 (N_15732,N_13334,N_14536);
nand U15733 (N_15733,N_14374,N_14551);
xor U15734 (N_15734,N_12773,N_13544);
or U15735 (N_15735,N_14700,N_15426);
and U15736 (N_15736,N_12703,N_14224);
and U15737 (N_15737,N_12859,N_14071);
and U15738 (N_15738,N_13107,N_14091);
or U15739 (N_15739,N_12973,N_13717);
nor U15740 (N_15740,N_13794,N_13277);
and U15741 (N_15741,N_13815,N_13757);
and U15742 (N_15742,N_13461,N_14979);
xnor U15743 (N_15743,N_14899,N_14959);
xnor U15744 (N_15744,N_14133,N_14558);
nand U15745 (N_15745,N_12821,N_15339);
nand U15746 (N_15746,N_13925,N_13562);
nor U15747 (N_15747,N_15427,N_15607);
nand U15748 (N_15748,N_13512,N_13483);
nor U15749 (N_15749,N_12850,N_12513);
nor U15750 (N_15750,N_13422,N_15121);
nand U15751 (N_15751,N_14754,N_15073);
xnor U15752 (N_15752,N_12724,N_13384);
and U15753 (N_15753,N_13957,N_13326);
xor U15754 (N_15754,N_15059,N_15357);
or U15755 (N_15755,N_14366,N_14254);
or U15756 (N_15756,N_14633,N_15597);
or U15757 (N_15757,N_13009,N_14442);
and U15758 (N_15758,N_14985,N_14772);
nand U15759 (N_15759,N_13294,N_15150);
nor U15760 (N_15760,N_13367,N_12800);
and U15761 (N_15761,N_14392,N_14824);
nand U15762 (N_15762,N_13595,N_13015);
nand U15763 (N_15763,N_15445,N_14270);
nor U15764 (N_15764,N_14078,N_12943);
xor U15765 (N_15765,N_14496,N_12991);
xor U15766 (N_15766,N_13548,N_14065);
nand U15767 (N_15767,N_15533,N_12633);
xnor U15768 (N_15768,N_15224,N_13057);
xnor U15769 (N_15769,N_14829,N_14834);
or U15770 (N_15770,N_13144,N_15381);
or U15771 (N_15771,N_12898,N_13524);
xor U15772 (N_15772,N_13425,N_14690);
or U15773 (N_15773,N_15299,N_14107);
xnor U15774 (N_15774,N_13639,N_13462);
or U15775 (N_15775,N_13458,N_15093);
nand U15776 (N_15776,N_15566,N_13082);
or U15777 (N_15777,N_13976,N_12715);
and U15778 (N_15778,N_14996,N_12662);
nand U15779 (N_15779,N_12637,N_15092);
and U15780 (N_15780,N_14736,N_13218);
nand U15781 (N_15781,N_13680,N_15203);
nand U15782 (N_15782,N_13332,N_13429);
nor U15783 (N_15783,N_12540,N_12531);
nand U15784 (N_15784,N_13569,N_13932);
nand U15785 (N_15785,N_13983,N_14395);
and U15786 (N_15786,N_13155,N_15154);
xnor U15787 (N_15787,N_13331,N_14194);
and U15788 (N_15788,N_13257,N_14913);
nor U15789 (N_15789,N_14889,N_12960);
and U15790 (N_15790,N_13491,N_12811);
nor U15791 (N_15791,N_13971,N_14916);
and U15792 (N_15792,N_12917,N_12830);
xnor U15793 (N_15793,N_13668,N_12926);
or U15794 (N_15794,N_14143,N_13743);
nor U15795 (N_15795,N_13186,N_14803);
xnor U15796 (N_15796,N_15284,N_14650);
nand U15797 (N_15797,N_12672,N_12792);
and U15798 (N_15798,N_13154,N_14971);
nor U15799 (N_15799,N_13818,N_15126);
nor U15800 (N_15800,N_12640,N_13699);
nor U15801 (N_15801,N_15011,N_14614);
xor U15802 (N_15802,N_13798,N_15453);
nand U15803 (N_15803,N_12769,N_13073);
nor U15804 (N_15804,N_13109,N_13059);
or U15805 (N_15805,N_14747,N_13942);
nor U15806 (N_15806,N_13000,N_13263);
and U15807 (N_15807,N_13552,N_13541);
and U15808 (N_15808,N_15181,N_14806);
or U15809 (N_15809,N_14611,N_15590);
nor U15810 (N_15810,N_13802,N_15129);
and U15811 (N_15811,N_12730,N_14204);
and U15812 (N_15812,N_13776,N_15135);
xor U15813 (N_15813,N_14680,N_14557);
nand U15814 (N_15814,N_14886,N_12618);
nand U15815 (N_15815,N_12583,N_13369);
and U15816 (N_15816,N_14651,N_13915);
and U15817 (N_15817,N_14362,N_13536);
and U15818 (N_15818,N_13640,N_15557);
and U15819 (N_15819,N_13270,N_14816);
and U15820 (N_15820,N_13753,N_12598);
or U15821 (N_15821,N_12538,N_13891);
nor U15822 (N_15822,N_15417,N_13070);
nand U15823 (N_15823,N_15133,N_14740);
xor U15824 (N_15824,N_15317,N_12785);
nand U15825 (N_15825,N_14554,N_13400);
and U15826 (N_15826,N_13638,N_15436);
xor U15827 (N_15827,N_12646,N_13267);
xnor U15828 (N_15828,N_13151,N_13558);
nand U15829 (N_15829,N_13972,N_14494);
nand U15830 (N_15830,N_15574,N_13259);
nor U15831 (N_15831,N_12783,N_15581);
xnor U15832 (N_15832,N_14042,N_13286);
nand U15833 (N_15833,N_13196,N_13078);
nand U15834 (N_15834,N_13417,N_13816);
or U15835 (N_15835,N_14473,N_14980);
xnor U15836 (N_15836,N_15282,N_13131);
or U15837 (N_15837,N_15119,N_12689);
and U15838 (N_15838,N_13502,N_14880);
or U15839 (N_15839,N_14216,N_14339);
nand U15840 (N_15840,N_14052,N_13923);
xnor U15841 (N_15841,N_13063,N_15141);
nor U15842 (N_15842,N_13979,N_13862);
nand U15843 (N_15843,N_14055,N_14832);
nor U15844 (N_15844,N_13892,N_13112);
nand U15845 (N_15845,N_15534,N_13823);
nand U15846 (N_15846,N_14447,N_12993);
nand U15847 (N_15847,N_12799,N_15399);
nand U15848 (N_15848,N_14553,N_15437);
or U15849 (N_15849,N_13620,N_13947);
nand U15850 (N_15850,N_12756,N_14432);
or U15851 (N_15851,N_13938,N_14704);
and U15852 (N_15852,N_14329,N_15555);
xnor U15853 (N_15853,N_14463,N_14605);
xnor U15854 (N_15854,N_15237,N_14053);
nor U15855 (N_15855,N_13682,N_15105);
nor U15856 (N_15856,N_13076,N_13404);
nand U15857 (N_15857,N_15623,N_15510);
nor U15858 (N_15858,N_13712,N_12767);
xor U15859 (N_15859,N_14712,N_14303);
nand U15860 (N_15860,N_15390,N_14305);
nand U15861 (N_15861,N_13948,N_13242);
xnor U15862 (N_15862,N_13650,N_14232);
or U15863 (N_15863,N_13026,N_15002);
and U15864 (N_15864,N_14687,N_14434);
and U15865 (N_15865,N_13770,N_12853);
and U15866 (N_15866,N_14644,N_15143);
nand U15867 (N_15867,N_15146,N_14635);
or U15868 (N_15868,N_13088,N_14850);
nand U15869 (N_15869,N_14243,N_13335);
nand U15870 (N_15870,N_14083,N_13501);
nor U15871 (N_15871,N_12679,N_13060);
nor U15872 (N_15872,N_13637,N_15486);
nand U15873 (N_15873,N_14267,N_14086);
or U15874 (N_15874,N_12881,N_13758);
nand U15875 (N_15875,N_13681,N_15006);
nor U15876 (N_15876,N_13204,N_13877);
nand U15877 (N_15877,N_13201,N_13674);
nor U15878 (N_15878,N_12977,N_12665);
and U15879 (N_15879,N_12863,N_14376);
nor U15880 (N_15880,N_14438,N_13345);
nor U15881 (N_15881,N_12819,N_13128);
or U15882 (N_15882,N_13732,N_14621);
nor U15883 (N_15883,N_13223,N_13251);
nand U15884 (N_15884,N_13763,N_15014);
nand U15885 (N_15885,N_14870,N_13910);
xnor U15886 (N_15886,N_13878,N_14620);
nand U15887 (N_15887,N_14292,N_14479);
or U15888 (N_15888,N_14180,N_15103);
nand U15889 (N_15889,N_14271,N_15005);
xor U15890 (N_15890,N_15344,N_15245);
xnor U15891 (N_15891,N_14105,N_14064);
xor U15892 (N_15892,N_14852,N_15478);
nor U15893 (N_15893,N_13178,N_14667);
and U15894 (N_15894,N_14347,N_13415);
nand U15895 (N_15895,N_12615,N_14645);
or U15896 (N_15896,N_13599,N_14813);
or U15897 (N_15897,N_14404,N_15415);
nand U15898 (N_15898,N_13838,N_13184);
and U15899 (N_15899,N_15584,N_13143);
and U15900 (N_15900,N_13846,N_12914);
xnor U15901 (N_15901,N_13711,N_13230);
nor U15902 (N_15902,N_13285,N_14038);
nor U15903 (N_15903,N_13287,N_14835);
nand U15904 (N_15904,N_15548,N_14749);
xnor U15905 (N_15905,N_15243,N_14750);
xnor U15906 (N_15906,N_13330,N_13657);
nand U15907 (N_15907,N_13889,N_15554);
nand U15908 (N_15908,N_15156,N_14480);
nor U15909 (N_15909,N_12720,N_13869);
and U15910 (N_15910,N_15501,N_14856);
nand U15911 (N_15911,N_13631,N_14952);
nor U15912 (N_15912,N_13048,N_15076);
nand U15913 (N_15913,N_13706,N_13629);
nand U15914 (N_15914,N_12913,N_12541);
and U15915 (N_15915,N_15202,N_14365);
or U15916 (N_15916,N_13880,N_14786);
nand U15917 (N_15917,N_14171,N_15576);
or U15918 (N_15918,N_14191,N_15614);
and U15919 (N_15919,N_13737,N_14045);
and U15920 (N_15920,N_14278,N_13963);
and U15921 (N_15921,N_13806,N_13888);
xnor U15922 (N_15922,N_13950,N_12842);
nand U15923 (N_15923,N_12697,N_15428);
nand U15924 (N_15924,N_14930,N_14726);
xnor U15925 (N_15925,N_15411,N_14041);
nand U15926 (N_15926,N_14741,N_14357);
nand U15927 (N_15927,N_14309,N_15132);
nand U15928 (N_15928,N_15159,N_15423);
and U15929 (N_15929,N_13825,N_14206);
xor U15930 (N_15930,N_14603,N_14010);
xnor U15931 (N_15931,N_15541,N_14158);
or U15932 (N_15932,N_15173,N_14015);
xnor U15933 (N_15933,N_15031,N_13350);
and U15934 (N_15934,N_14195,N_15400);
nand U15935 (N_15935,N_12673,N_14067);
nor U15936 (N_15936,N_14839,N_13864);
nand U15937 (N_15937,N_14770,N_15211);
nor U15938 (N_15938,N_13445,N_13397);
nand U15939 (N_15939,N_14169,N_13510);
or U15940 (N_15940,N_14332,N_14239);
and U15941 (N_15941,N_13436,N_12526);
or U15942 (N_15942,N_13744,N_15023);
or U15943 (N_15943,N_13723,N_12625);
and U15944 (N_15944,N_13206,N_12843);
xor U15945 (N_15945,N_15186,N_12711);
xnor U15946 (N_15946,N_14882,N_14773);
xor U15947 (N_15947,N_15101,N_14393);
nand U15948 (N_15948,N_13547,N_13272);
nor U15949 (N_15949,N_12995,N_14273);
nor U15950 (N_15950,N_14972,N_15216);
xnor U15951 (N_15951,N_14819,N_14578);
nor U15952 (N_15952,N_13159,N_12937);
nand U15953 (N_15953,N_13767,N_12525);
nand U15954 (N_15954,N_14337,N_13728);
or U15955 (N_15955,N_14570,N_15456);
nor U15956 (N_15956,N_12869,N_13844);
nor U15957 (N_15957,N_13746,N_12817);
nor U15958 (N_15958,N_14821,N_14665);
nand U15959 (N_15959,N_13514,N_14487);
xor U15960 (N_15960,N_13421,N_14211);
nor U15961 (N_15961,N_15281,N_13577);
nand U15962 (N_15962,N_14288,N_14630);
and U15963 (N_15963,N_13987,N_14845);
nand U15964 (N_15964,N_13307,N_12846);
nor U15965 (N_15965,N_13482,N_15573);
xor U15966 (N_15966,N_14225,N_15450);
xnor U15967 (N_15967,N_14139,N_14785);
or U15968 (N_15968,N_14351,N_12952);
and U15969 (N_15969,N_15379,N_12601);
xnor U15970 (N_15970,N_13093,N_13181);
or U15971 (N_15971,N_13383,N_12981);
xnor U15972 (N_15972,N_12599,N_14710);
nand U15973 (N_15973,N_13520,N_15066);
or U15974 (N_15974,N_15296,N_13909);
or U15975 (N_15975,N_14379,N_13999);
or U15976 (N_15976,N_13454,N_12661);
xor U15977 (N_15977,N_14705,N_14576);
or U15978 (N_15978,N_13085,N_14932);
nor U15979 (N_15979,N_14629,N_13720);
nand U15980 (N_15980,N_13591,N_13228);
nand U15981 (N_15981,N_14818,N_15391);
or U15982 (N_15982,N_15559,N_14793);
or U15983 (N_15983,N_15096,N_14002);
nand U15984 (N_15984,N_13249,N_15158);
and U15985 (N_15985,N_12860,N_13022);
nand U15986 (N_15986,N_13875,N_14836);
xor U15987 (N_15987,N_13601,N_15356);
and U15988 (N_15988,N_12605,N_14440);
and U15989 (N_15989,N_14599,N_13969);
xnor U15990 (N_15990,N_15268,N_13023);
and U15991 (N_15991,N_15246,N_12519);
or U15992 (N_15992,N_13386,N_13451);
or U15993 (N_15993,N_15372,N_15354);
nor U15994 (N_15994,N_13004,N_13139);
or U15995 (N_15995,N_14062,N_12746);
nor U15996 (N_15996,N_13352,N_13361);
nand U15997 (N_15997,N_12809,N_12622);
and U15998 (N_15998,N_14356,N_14566);
xor U15999 (N_15999,N_15371,N_15535);
nand U16000 (N_16000,N_15157,N_14093);
nor U16001 (N_16001,N_12854,N_14142);
or U16002 (N_16002,N_13020,N_14150);
nor U16003 (N_16003,N_13202,N_13813);
nor U16004 (N_16004,N_13792,N_14236);
nand U16005 (N_16005,N_15302,N_14246);
xnor U16006 (N_16006,N_13895,N_13295);
or U16007 (N_16007,N_14573,N_14036);
and U16008 (N_16008,N_14348,N_13760);
and U16009 (N_16009,N_12839,N_13410);
nand U16010 (N_16010,N_12958,N_14745);
and U16011 (N_16011,N_14501,N_14848);
or U16012 (N_16012,N_14364,N_14352);
nand U16013 (N_16013,N_13232,N_14855);
or U16014 (N_16014,N_12970,N_15513);
nand U16015 (N_16015,N_14318,N_15416);
or U16016 (N_16016,N_13724,N_14724);
nand U16017 (N_16017,N_14234,N_14919);
nand U16018 (N_16018,N_12659,N_14343);
and U16019 (N_16019,N_13123,N_14373);
nor U16020 (N_16020,N_13709,N_15113);
nand U16021 (N_16021,N_13027,N_13473);
and U16022 (N_16022,N_14543,N_13310);
xnor U16023 (N_16023,N_12514,N_12566);
xor U16024 (N_16024,N_14871,N_14085);
nor U16025 (N_16025,N_14507,N_14713);
and U16026 (N_16026,N_14151,N_12691);
nor U16027 (N_16027,N_15125,N_13284);
xor U16028 (N_16028,N_13831,N_13325);
nor U16029 (N_16029,N_15419,N_13626);
nor U16030 (N_16030,N_13559,N_15516);
or U16031 (N_16031,N_13667,N_13679);
and U16032 (N_16032,N_13973,N_12904);
nand U16033 (N_16033,N_15155,N_13203);
nand U16034 (N_16034,N_13578,N_15508);
and U16035 (N_16035,N_13086,N_15489);
nor U16036 (N_16036,N_15473,N_13687);
and U16037 (N_16037,N_14826,N_13176);
xnor U16038 (N_16038,N_14259,N_12872);
nand U16039 (N_16039,N_14728,N_13374);
xor U16040 (N_16040,N_12939,N_14094);
nor U16041 (N_16041,N_14792,N_13847);
and U16042 (N_16042,N_15195,N_13897);
and U16043 (N_16043,N_13075,N_15575);
or U16044 (N_16044,N_14827,N_14481);
and U16045 (N_16045,N_14097,N_13546);
xor U16046 (N_16046,N_13628,N_13167);
nor U16047 (N_16047,N_14958,N_12560);
and U16048 (N_16048,N_14281,N_15571);
xnor U16049 (N_16049,N_14622,N_12675);
nor U16050 (N_16050,N_13588,N_12867);
or U16051 (N_16051,N_13654,N_13148);
and U16052 (N_16052,N_13926,N_15329);
and U16053 (N_16053,N_15238,N_14682);
or U16054 (N_16054,N_13393,N_14711);
nand U16055 (N_16055,N_14170,N_13564);
or U16056 (N_16056,N_12517,N_12638);
and U16057 (N_16057,N_12718,N_14341);
nand U16058 (N_16058,N_13234,N_13893);
nor U16059 (N_16059,N_12629,N_15000);
or U16060 (N_16060,N_13871,N_13658);
xor U16061 (N_16061,N_14218,N_14312);
xnor U16062 (N_16062,N_14795,N_14123);
or U16063 (N_16063,N_14237,N_13666);
nand U16064 (N_16064,N_15289,N_12770);
and U16065 (N_16065,N_13635,N_14082);
nor U16066 (N_16066,N_14893,N_12515);
nor U16067 (N_16067,N_13215,N_12861);
nand U16068 (N_16068,N_15053,N_14276);
xnor U16069 (N_16069,N_14961,N_13124);
nand U16070 (N_16070,N_14059,N_15585);
or U16071 (N_16071,N_14815,N_12965);
nor U16072 (N_16072,N_12838,N_14965);
nand U16073 (N_16073,N_12942,N_12796);
xnor U16074 (N_16074,N_14548,N_14129);
nor U16075 (N_16075,N_12816,N_15395);
or U16076 (N_16076,N_14662,N_15212);
nor U16077 (N_16077,N_12955,N_13288);
nor U16078 (N_16078,N_13340,N_13195);
xor U16079 (N_16079,N_12882,N_14152);
nor U16080 (N_16080,N_14954,N_15518);
or U16081 (N_16081,N_14381,N_12921);
or U16082 (N_16082,N_13250,N_14784);
or U16083 (N_16083,N_14529,N_12580);
nand U16084 (N_16084,N_15394,N_14090);
nand U16085 (N_16085,N_15234,N_13317);
nand U16086 (N_16086,N_15192,N_15207);
nand U16087 (N_16087,N_14988,N_15565);
nand U16088 (N_16088,N_14619,N_15545);
xnor U16089 (N_16089,N_14407,N_14114);
or U16090 (N_16090,N_13851,N_12876);
xor U16091 (N_16091,N_14937,N_14677);
and U16092 (N_16092,N_13449,N_13675);
nand U16093 (N_16093,N_15024,N_12964);
and U16094 (N_16094,N_14948,N_15459);
nand U16095 (N_16095,N_13803,N_12906);
and U16096 (N_16096,N_15123,N_12655);
and U16097 (N_16097,N_12757,N_13433);
nor U16098 (N_16098,N_13507,N_15063);
and U16099 (N_16099,N_14873,N_13087);
nor U16100 (N_16100,N_14500,N_13156);
nand U16101 (N_16101,N_12848,N_13296);
nand U16102 (N_16102,N_12664,N_15521);
or U16103 (N_16103,N_13114,N_12933);
xor U16104 (N_16104,N_14058,N_13344);
nand U16105 (N_16105,N_15291,N_15134);
xor U16106 (N_16106,N_15507,N_13241);
nand U16107 (N_16107,N_13375,N_13199);
nor U16108 (N_16108,N_14075,N_12585);
nand U16109 (N_16109,N_13945,N_15235);
nand U16110 (N_16110,N_13104,N_13072);
nor U16111 (N_16111,N_14647,N_15217);
nor U16112 (N_16112,N_14540,N_14304);
nand U16113 (N_16113,N_15512,N_14422);
nor U16114 (N_16114,N_14950,N_15589);
xor U16115 (N_16115,N_14240,N_13633);
or U16116 (N_16116,N_14989,N_12779);
nand U16117 (N_16117,N_13399,N_14517);
or U16118 (N_16118,N_13122,N_13565);
xor U16119 (N_16119,N_14923,N_14966);
nor U16120 (N_16120,N_12738,N_13165);
nand U16121 (N_16121,N_14157,N_13033);
xor U16122 (N_16122,N_13837,N_12858);
and U16123 (N_16123,N_13044,N_13011);
nor U16124 (N_16124,N_12600,N_14401);
or U16125 (N_16125,N_13252,N_12959);
nor U16126 (N_16126,N_13935,N_15264);
nor U16127 (N_16127,N_14787,N_13566);
and U16128 (N_16128,N_14903,N_14092);
xor U16129 (N_16129,N_14691,N_15370);
and U16130 (N_16130,N_14938,N_12919);
nor U16131 (N_16131,N_14156,N_13920);
xor U16132 (N_16132,N_15563,N_13389);
and U16133 (N_16133,N_12974,N_13664);
and U16134 (N_16134,N_13382,N_13006);
xnor U16135 (N_16135,N_13188,N_15263);
nor U16136 (N_16136,N_13890,N_14778);
nor U16137 (N_16137,N_15420,N_14289);
xor U16138 (N_16138,N_14984,N_14951);
or U16139 (N_16139,N_13961,N_14617);
nand U16140 (N_16140,N_15052,N_13854);
and U16141 (N_16141,N_12744,N_13496);
nor U16142 (N_16142,N_15613,N_13539);
nor U16143 (N_16143,N_15412,N_14764);
nand U16144 (N_16144,N_12501,N_13554);
and U16145 (N_16145,N_15531,N_14969);
nand U16146 (N_16146,N_13298,N_14623);
or U16147 (N_16147,N_13119,N_14998);
and U16148 (N_16148,N_14420,N_13600);
xnor U16149 (N_16149,N_15338,N_14399);
xnor U16150 (N_16150,N_13349,N_13171);
nand U16151 (N_16151,N_13677,N_14355);
nor U16152 (N_16152,N_14879,N_13907);
xnor U16153 (N_16153,N_15591,N_15088);
xnor U16154 (N_16154,N_12668,N_15401);
and U16155 (N_16155,N_15083,N_14334);
xnor U16156 (N_16156,N_14096,N_14875);
and U16157 (N_16157,N_13630,N_14302);
nor U16158 (N_16158,N_15147,N_12575);
nand U16159 (N_16159,N_14028,N_13900);
nor U16160 (N_16160,N_15010,N_12578);
or U16161 (N_16161,N_14508,N_14499);
nand U16162 (N_16162,N_13964,N_12826);
nand U16163 (N_16163,N_13814,N_14004);
nand U16164 (N_16164,N_15182,N_14904);
xnor U16165 (N_16165,N_13168,N_13117);
and U16166 (N_16166,N_15477,N_13568);
nor U16167 (N_16167,N_13453,N_15470);
or U16168 (N_16168,N_12503,N_12892);
or U16169 (N_16169,N_13320,N_13538);
or U16170 (N_16170,N_12908,N_12777);
or U16171 (N_16171,N_13498,N_14167);
and U16172 (N_16172,N_13670,N_15439);
or U16173 (N_16173,N_14900,N_13774);
xnor U16174 (N_16174,N_13207,N_12941);
xor U16175 (N_16175,N_12915,N_12516);
or U16176 (N_16176,N_13924,N_13580);
nor U16177 (N_16177,N_12610,N_13025);
nor U16178 (N_16178,N_14185,N_15438);
and U16179 (N_16179,N_15309,N_14549);
and U16180 (N_16180,N_13471,N_15128);
or U16181 (N_16181,N_14450,N_13887);
or U16182 (N_16182,N_14634,N_13081);
and U16183 (N_16183,N_13616,N_15496);
nand U16184 (N_16184,N_14915,N_14780);
nand U16185 (N_16185,N_12976,N_13521);
nand U16186 (N_16186,N_14251,N_14506);
xor U16187 (N_16187,N_13855,N_15221);
nand U16188 (N_16188,N_14222,N_14897);
nor U16189 (N_16189,N_15298,N_14037);
xnor U16190 (N_16190,N_13348,N_15409);
xor U16191 (N_16191,N_13381,N_13777);
and U16192 (N_16192,N_14220,N_14226);
xor U16193 (N_16193,N_15558,N_12570);
nor U16194 (N_16194,N_13455,N_13906);
nand U16195 (N_16195,N_12698,N_14322);
nor U16196 (N_16196,N_14794,N_13254);
xor U16197 (N_16197,N_12916,N_12751);
nand U16198 (N_16198,N_13185,N_15183);
xor U16199 (N_16199,N_14639,N_13705);
or U16200 (N_16200,N_14109,N_13698);
nor U16201 (N_16201,N_14396,N_14949);
or U16202 (N_16202,N_12666,N_13986);
nand U16203 (N_16203,N_13614,N_14646);
nor U16204 (N_16204,N_14202,N_14272);
nor U16205 (N_16205,N_12616,N_12654);
or U16206 (N_16206,N_15350,N_13183);
xnor U16207 (N_16207,N_14674,N_14284);
nand U16208 (N_16208,N_15261,N_14618);
nor U16209 (N_16209,N_13231,N_13820);
nor U16210 (N_16210,N_13590,N_14721);
xnor U16211 (N_16211,N_12741,N_13738);
nor U16212 (N_16212,N_15177,N_13189);
or U16213 (N_16213,N_14477,N_13940);
nor U16214 (N_16214,N_14166,N_14330);
nand U16215 (N_16215,N_13443,N_12967);
xnor U16216 (N_16216,N_15469,N_15067);
nand U16217 (N_16217,N_15152,N_15497);
xor U16218 (N_16218,N_14702,N_15550);
nor U16219 (N_16219,N_14643,N_15429);
or U16220 (N_16220,N_14546,N_13585);
nand U16221 (N_16221,N_13010,N_14569);
or U16222 (N_16222,N_14324,N_13665);
nor U16223 (N_16223,N_14884,N_15278);
nand U16224 (N_16224,N_15467,N_14663);
nor U16225 (N_16225,N_14720,N_12709);
or U16226 (N_16226,N_12608,N_15622);
nand U16227 (N_16227,N_14955,N_13772);
nand U16228 (N_16228,N_14005,N_13450);
or U16229 (N_16229,N_14072,N_14340);
and U16230 (N_16230,N_13759,N_15306);
xor U16231 (N_16231,N_15262,N_14669);
or U16232 (N_16232,N_14858,N_14666);
nor U16233 (N_16233,N_13460,N_15407);
and U16234 (N_16234,N_14891,N_14502);
nor U16235 (N_16235,N_15460,N_14602);
nor U16236 (N_16236,N_13260,N_15225);
nand U16237 (N_16237,N_15250,N_12658);
nand U16238 (N_16238,N_14742,N_15506);
or U16239 (N_16239,N_12528,N_15226);
or U16240 (N_16240,N_15402,N_13162);
xor U16241 (N_16241,N_13647,N_13248);
or U16242 (N_16242,N_14174,N_15218);
and U16243 (N_16243,N_12808,N_12983);
nand U16244 (N_16244,N_14080,N_15322);
and U16245 (N_16245,N_13937,N_12645);
or U16246 (N_16246,N_13655,N_15117);
or U16247 (N_16247,N_15615,N_14986);
or U16248 (N_16248,N_13238,N_14509);
or U16249 (N_16249,N_15085,N_15240);
and U16250 (N_16250,N_15009,N_14026);
xnor U16251 (N_16251,N_13722,N_14087);
and U16252 (N_16252,N_13378,N_15283);
or U16253 (N_16253,N_14520,N_14636);
or U16254 (N_16254,N_14350,N_14698);
nor U16255 (N_16255,N_12831,N_14946);
nand U16256 (N_16256,N_12628,N_13469);
and U16257 (N_16257,N_15027,N_14405);
xor U16258 (N_16258,N_13212,N_15539);
nor U16259 (N_16259,N_13412,N_14476);
and U16260 (N_16260,N_13797,N_14497);
xnor U16261 (N_16261,N_15606,N_14047);
and U16262 (N_16262,N_13066,N_14911);
nand U16263 (N_16263,N_14345,N_15065);
nor U16264 (N_16264,N_14177,N_14582);
and U16265 (N_16265,N_15392,N_13801);
nor U16266 (N_16266,N_15255,N_13214);
nor U16267 (N_16267,N_15114,N_13409);
xor U16268 (N_16268,N_15546,N_12870);
or U16269 (N_16269,N_15454,N_12594);
or U16270 (N_16270,N_14184,N_13586);
nor U16271 (N_16271,N_12739,N_14408);
nand U16272 (N_16272,N_14103,N_14993);
and U16273 (N_16273,N_13634,N_14475);
xor U16274 (N_16274,N_13360,N_13149);
nand U16275 (N_16275,N_14034,N_13691);
xnor U16276 (N_16276,N_14161,N_13080);
xnor U16277 (N_16277,N_15025,N_15118);
or U16278 (N_16278,N_15239,N_13380);
and U16279 (N_16279,N_14162,N_13943);
nand U16280 (N_16280,N_14159,N_13953);
nand U16281 (N_16281,N_14124,N_15505);
and U16282 (N_16282,N_12587,N_14280);
nor U16283 (N_16283,N_12805,N_14715);
xor U16284 (N_16284,N_12586,N_15015);
nor U16285 (N_16285,N_13594,N_14113);
and U16286 (N_16286,N_14905,N_15248);
and U16287 (N_16287,N_12620,N_13570);
and U16288 (N_16288,N_14851,N_12747);
and U16289 (N_16289,N_14279,N_12918);
nand U16290 (N_16290,N_14003,N_14692);
and U16291 (N_16291,N_15193,N_15100);
or U16292 (N_16292,N_13007,N_14217);
and U16293 (N_16293,N_15213,N_13084);
xor U16294 (N_16294,N_15190,N_13314);
nand U16295 (N_16295,N_12644,N_12750);
and U16296 (N_16296,N_12888,N_15116);
or U16297 (N_16297,N_13255,N_13956);
and U16298 (N_16298,N_12884,N_14685);
nand U16299 (N_16299,N_13908,N_13354);
or U16300 (N_16300,N_12814,N_12878);
nand U16301 (N_16301,N_13688,N_14429);
xnor U16302 (N_16302,N_14748,N_15458);
nand U16303 (N_16303,N_13136,N_14197);
and U16304 (N_16304,N_12875,N_13730);
and U16305 (N_16305,N_13993,N_12865);
and U16306 (N_16306,N_13885,N_14371);
nand U16307 (N_16307,N_12900,N_12856);
xnor U16308 (N_16308,N_14631,N_15396);
nand U16309 (N_16309,N_14138,N_13824);
or U16310 (N_16310,N_12542,N_12992);
and U16311 (N_16311,N_14732,N_12732);
or U16312 (N_16312,N_14597,N_14753);
xor U16313 (N_16313,N_14596,N_12889);
and U16314 (N_16314,N_14735,N_13258);
and U16315 (N_16315,N_13689,N_14843);
and U16316 (N_16316,N_14321,N_12998);
nor U16317 (N_16317,N_12911,N_15311);
xor U16318 (N_16318,N_13771,N_14774);
or U16319 (N_16319,N_15341,N_14282);
nand U16320 (N_16320,N_13046,N_14221);
or U16321 (N_16321,N_15537,N_13787);
nor U16322 (N_16322,N_13222,N_13394);
nor U16323 (N_16323,N_12740,N_14613);
and U16324 (N_16324,N_13516,N_12971);
nand U16325 (N_16325,N_13853,N_14737);
or U16326 (N_16326,N_13013,N_13118);
nand U16327 (N_16327,N_13531,N_14907);
and U16328 (N_16328,N_13246,N_15247);
and U16329 (N_16329,N_14076,N_12563);
nand U16330 (N_16330,N_12899,N_14483);
nand U16331 (N_16331,N_12928,N_13550);
nand U16332 (N_16332,N_14388,N_12543);
and U16333 (N_16333,N_12508,N_15230);
or U16334 (N_16334,N_15068,N_13219);
xnor U16335 (N_16335,N_13280,N_13605);
xor U16336 (N_16336,N_14323,N_14039);
xnor U16337 (N_16337,N_14579,N_14563);
or U16338 (N_16338,N_15617,N_15175);
nor U16339 (N_16339,N_13985,N_15410);
nand U16340 (N_16340,N_14307,N_12550);
xnor U16341 (N_16341,N_14196,N_13998);
and U16342 (N_16342,N_14470,N_13977);
nor U16343 (N_16343,N_13276,N_13339);
nor U16344 (N_16344,N_15095,N_14586);
nor U16345 (N_16345,N_15075,N_14590);
xor U16346 (N_16346,N_15343,N_13949);
or U16347 (N_16347,N_12985,N_13828);
nor U16348 (N_16348,N_12590,N_14970);
and U16349 (N_16349,N_13490,N_13556);
nor U16350 (N_16350,N_14909,N_13135);
xor U16351 (N_16351,N_14021,N_14119);
or U16352 (N_16352,N_15131,N_12982);
and U16353 (N_16353,N_13543,N_13200);
and U16354 (N_16354,N_14731,N_12833);
xnor U16355 (N_16355,N_14296,N_15209);
nand U16356 (N_16356,N_15017,N_14233);
nand U16357 (N_16357,N_14616,N_12556);
xnor U16358 (N_16358,N_15111,N_13405);
nand U16359 (N_16359,N_13309,N_14783);
and U16360 (N_16360,N_13511,N_14458);
or U16361 (N_16361,N_12987,N_13508);
xnor U16362 (N_16362,N_14530,N_12807);
xor U16363 (N_16363,N_14927,N_13789);
xnor U16364 (N_16364,N_12852,N_13922);
and U16365 (N_16365,N_12948,N_13161);
xor U16366 (N_16366,N_12567,N_14297);
nand U16367 (N_16367,N_12782,N_14445);
nand U16368 (N_16368,N_12812,N_14455);
nor U16369 (N_16369,N_14591,N_14673);
nand U16370 (N_16370,N_14017,N_13058);
xor U16371 (N_16371,N_15332,N_15072);
nor U16372 (N_16372,N_13731,N_13480);
and U16373 (N_16373,N_15321,N_12890);
or U16374 (N_16374,N_13704,N_14810);
nor U16375 (N_16375,N_15178,N_15487);
or U16376 (N_16376,N_14771,N_13958);
nor U16377 (N_16377,N_14326,N_14696);
xnor U16378 (N_16378,N_13805,N_12879);
and U16379 (N_16379,N_15446,N_13965);
nand U16380 (N_16380,N_15257,N_12573);
and U16381 (N_16381,N_14145,N_14664);
and U16382 (N_16382,N_15028,N_14120);
nor U16383 (N_16383,N_13918,N_12696);
and U16384 (N_16384,N_12743,N_13448);
nand U16385 (N_16385,N_14452,N_12630);
nor U16386 (N_16386,N_14564,N_12546);
xnor U16387 (N_16387,N_14498,N_14263);
nor U16388 (N_16388,N_14176,N_12588);
xnor U16389 (N_16389,N_15232,N_13574);
xor U16390 (N_16390,N_13715,N_13663);
nor U16391 (N_16391,N_12871,N_15293);
nor U16392 (N_16392,N_15140,N_12728);
xnor U16393 (N_16393,N_12536,N_13111);
xnor U16394 (N_16394,N_14854,N_14684);
and U16395 (N_16395,N_13780,N_15272);
nor U16396 (N_16396,N_15385,N_12787);
nor U16397 (N_16397,N_14587,N_14798);
xnor U16398 (N_16398,N_14572,N_13018);
and U16399 (N_16399,N_12736,N_14431);
and U16400 (N_16400,N_12847,N_14583);
and U16401 (N_16401,N_13603,N_14471);
nor U16402 (N_16402,N_14349,N_15504);
and U16403 (N_16403,N_12989,N_12702);
xor U16404 (N_16404,N_13120,N_15418);
or U16405 (N_16405,N_13362,N_13368);
or U16406 (N_16406,N_13990,N_12771);
or U16407 (N_16407,N_15060,N_13624);
nand U16408 (N_16408,N_14207,N_12923);
and U16409 (N_16409,N_13506,N_13463);
nand U16410 (N_16410,N_13573,N_14104);
and U16411 (N_16411,N_14533,N_14921);
nand U16412 (N_16412,N_14523,N_15375);
nand U16413 (N_16413,N_12512,N_14757);
and U16414 (N_16414,N_13607,N_13459);
or U16415 (N_16415,N_14269,N_12502);
and U16416 (N_16416,N_13357,N_15578);
nor U16417 (N_16417,N_13669,N_12552);
and U16418 (N_16418,N_14132,N_15586);
or U16419 (N_16419,N_13921,N_14457);
and U16420 (N_16420,N_12932,N_13396);
or U16421 (N_16421,N_14977,N_12500);
nand U16422 (N_16422,N_13418,N_14857);
nor U16423 (N_16423,N_14920,N_13095);
nand U16424 (N_16424,N_12574,N_13526);
and U16425 (N_16425,N_15382,N_14962);
or U16426 (N_16426,N_14864,N_12534);
nand U16427 (N_16427,N_15187,N_14165);
nand U16428 (N_16428,N_12931,N_14146);
nor U16429 (N_16429,N_13431,N_15022);
or U16430 (N_16430,N_14048,N_15184);
nand U16431 (N_16431,N_14009,N_13134);
and U16432 (N_16432,N_14627,N_12930);
nand U16433 (N_16433,N_15286,N_14526);
and U16434 (N_16434,N_14016,N_13761);
xor U16435 (N_16435,N_12963,N_12619);
nand U16436 (N_16436,N_12940,N_15176);
nand U16437 (N_16437,N_13477,N_13673);
and U16438 (N_16438,N_14102,N_13105);
or U16439 (N_16439,N_14413,N_15274);
xor U16440 (N_16440,N_13229,N_12681);
or U16441 (N_16441,N_13782,N_12840);
and U16442 (N_16442,N_13355,N_13739);
nor U16443 (N_16443,N_14552,N_12597);
nor U16444 (N_16444,N_15366,N_14359);
nor U16445 (N_16445,N_13308,N_15580);
nand U16446 (N_16446,N_15142,N_14495);
or U16447 (N_16447,N_14316,N_14301);
or U16448 (N_16448,N_15304,N_15214);
xnor U16449 (N_16449,N_12910,N_12909);
nor U16450 (N_16450,N_13329,N_12749);
nand U16451 (N_16451,N_15386,N_13800);
nand U16452 (N_16452,N_12726,N_15045);
or U16453 (N_16453,N_13954,N_13696);
xnor U16454 (N_16454,N_15325,N_14182);
nand U16455 (N_16455,N_14400,N_12705);
nand U16456 (N_16456,N_14101,N_15342);
nor U16457 (N_16457,N_13750,N_12897);
xnor U16458 (N_16458,N_13540,N_14545);
xnor U16459 (N_16459,N_13391,N_14914);
or U16460 (N_16460,N_13210,N_13700);
xnor U16461 (N_16461,N_12685,N_13532);
nand U16462 (N_16462,N_13226,N_15080);
nand U16463 (N_16463,N_13359,N_13551);
and U16464 (N_16464,N_15424,N_15043);
nor U16465 (N_16465,N_13372,N_13835);
or U16466 (N_16466,N_15553,N_14890);
nor U16467 (N_16467,N_13321,N_13527);
and U16468 (N_16468,N_13446,N_12868);
nor U16469 (N_16469,N_12945,N_14484);
and U16470 (N_16470,N_15621,N_14199);
or U16471 (N_16471,N_14467,N_13036);
and U16472 (N_16472,N_13067,N_14127);
nand U16473 (N_16473,N_13606,N_13192);
nand U16474 (N_16474,N_13849,N_14556);
and U16475 (N_16475,N_13609,N_13035);
xnor U16476 (N_16476,N_13049,N_14253);
and U16477 (N_16477,N_13695,N_15515);
nand U16478 (N_16478,N_14008,N_14730);
nand U16479 (N_16479,N_13303,N_14902);
or U16480 (N_16480,N_12760,N_13883);
and U16481 (N_16481,N_13646,N_13503);
nand U16482 (N_16482,N_14032,N_14223);
or U16483 (N_16483,N_14423,N_14214);
nand U16484 (N_16484,N_13645,N_14867);
and U16485 (N_16485,N_15340,N_14252);
or U16486 (N_16486,N_14863,N_14917);
xnor U16487 (N_16487,N_14574,N_14844);
nand U16488 (N_16488,N_14689,N_15035);
xor U16489 (N_16489,N_14070,N_12554);
and U16490 (N_16490,N_13575,N_12758);
nand U16491 (N_16491,N_14734,N_13358);
nand U16492 (N_16492,N_13652,N_13221);
xor U16493 (N_16493,N_14228,N_14380);
xor U16494 (N_16494,N_15413,N_13147);
nand U16495 (N_16495,N_14044,N_15029);
nor U16496 (N_16496,N_13416,N_12994);
nor U16497 (N_16497,N_15166,N_14073);
nor U16498 (N_16498,N_15596,N_13478);
nand U16499 (N_16499,N_14718,N_14609);
nand U16500 (N_16500,N_12935,N_13312);
and U16501 (N_16501,N_13742,N_14716);
nand U16502 (N_16502,N_15055,N_12692);
or U16503 (N_16503,N_13982,N_14658);
nand U16504 (N_16504,N_12798,N_14888);
or U16505 (N_16505,N_15180,N_13966);
nor U16506 (N_16506,N_13290,N_13012);
nand U16507 (N_16507,N_14179,N_13205);
nor U16508 (N_16508,N_14027,N_12649);
and U16509 (N_16509,N_15098,N_14390);
and U16510 (N_16510,N_15270,N_14153);
nand U16511 (N_16511,N_14320,N_13233);
and U16512 (N_16512,N_14247,N_14974);
nor U16513 (N_16513,N_15452,N_14173);
nor U16514 (N_16514,N_12694,N_13065);
or U16515 (N_16515,N_14719,N_13385);
or U16516 (N_16516,N_12778,N_15542);
and U16517 (N_16517,N_13518,N_14411);
or U16518 (N_16518,N_13623,N_15253);
nand U16519 (N_16519,N_15479,N_14661);
and U16520 (N_16520,N_13515,N_13829);
or U16521 (N_16521,N_14943,N_12954);
or U16522 (N_16522,N_15349,N_13902);
or U16523 (N_16523,N_13833,N_15242);
nand U16524 (N_16524,N_12835,N_13021);
nand U16525 (N_16525,N_15425,N_14242);
or U16526 (N_16526,N_13113,N_15577);
and U16527 (N_16527,N_12581,N_14725);
and U16528 (N_16528,N_14648,N_14128);
and U16529 (N_16529,N_14531,N_14116);
nand U16530 (N_16530,N_14079,N_12555);
or U16531 (N_16531,N_14369,N_13452);
nor U16532 (N_16532,N_13741,N_14555);
nor U16533 (N_16533,N_14987,N_13530);
and U16534 (N_16534,N_14069,N_14245);
nand U16535 (N_16535,N_15538,N_13485);
xnor U16536 (N_16536,N_13589,N_12521);
nor U16537 (N_16537,N_15388,N_15616);
or U16538 (N_16538,N_15057,N_14111);
and U16539 (N_16539,N_14865,N_13395);
xor U16540 (N_16540,N_12648,N_15162);
xor U16541 (N_16541,N_13127,N_13519);
nand U16542 (N_16542,N_12844,N_12652);
nor U16543 (N_16543,N_13403,N_13611);
nand U16544 (N_16544,N_13781,N_13172);
and U16545 (N_16545,N_14874,N_13437);
xor U16546 (N_16546,N_13729,N_12707);
and U16547 (N_16547,N_15106,N_14361);
nor U16548 (N_16548,N_14628,N_13002);
nor U16549 (N_16549,N_13402,N_12522);
and U16550 (N_16550,N_13662,N_14976);
nand U16551 (N_16551,N_14910,N_14274);
and U16552 (N_16552,N_12669,N_14295);
nor U16553 (N_16553,N_12624,N_13786);
nand U16554 (N_16554,N_14632,N_12896);
xnor U16555 (N_16555,N_13783,N_14007);
xnor U16556 (N_16556,N_14641,N_15602);
nor U16557 (N_16557,N_15347,N_14210);
or U16558 (N_16558,N_14790,N_13643);
nand U16559 (N_16559,N_13882,N_14638);
nor U16560 (N_16560,N_14933,N_15041);
or U16561 (N_16561,N_14981,N_14940);
nor U16562 (N_16562,N_14328,N_15603);
nand U16563 (N_16563,N_15474,N_12549);
nor U16564 (N_16564,N_13504,N_13465);
nand U16565 (N_16565,N_13211,N_13099);
or U16566 (N_16566,N_14446,N_12596);
nor U16567 (N_16567,N_13371,N_13198);
xnor U16568 (N_16568,N_13988,N_15524);
or U16569 (N_16569,N_14125,N_14739);
xor U16570 (N_16570,N_15449,N_15148);
and U16571 (N_16571,N_14807,N_14767);
or U16572 (N_16572,N_15222,N_13870);
xnor U16573 (N_16573,N_12627,N_12657);
xnor U16574 (N_16574,N_14928,N_15001);
and U16575 (N_16575,N_12880,N_15046);
nor U16576 (N_16576,N_13951,N_14887);
xnor U16577 (N_16577,N_15551,N_13500);
and U16578 (N_16578,N_15090,N_13563);
xor U16579 (N_16579,N_13528,N_15169);
nand U16580 (N_16580,N_14802,N_14336);
and U16581 (N_16581,N_12641,N_13055);
xnor U16582 (N_16582,N_12579,N_13708);
nor U16583 (N_16583,N_15300,N_15227);
xor U16584 (N_16584,N_15434,N_13690);
or U16585 (N_16585,N_14192,N_14367);
or U16586 (N_16586,N_15564,N_14285);
and U16587 (N_16587,N_15220,N_13039);
and U16588 (N_16588,N_15488,N_13523);
nor U16589 (N_16589,N_14172,N_13860);
xnor U16590 (N_16590,N_13748,N_13725);
nand U16591 (N_16591,N_14019,N_14402);
xnor U16592 (N_16592,N_13180,N_15231);
nand U16593 (N_16593,N_15364,N_15397);
nor U16594 (N_16594,N_13884,N_13441);
xnor U16595 (N_16595,N_14490,N_12979);
or U16596 (N_16596,N_12925,N_14265);
nor U16597 (N_16597,N_15312,N_13930);
and U16598 (N_16598,N_13721,N_15167);
nand U16599 (N_16599,N_13406,N_13807);
and U16600 (N_16600,N_13901,N_13734);
and U16601 (N_16601,N_14260,N_15174);
nor U16602 (N_16602,N_14606,N_15333);
nand U16603 (N_16603,N_15049,N_14317);
xnor U16604 (N_16604,N_12593,N_15583);
or U16605 (N_16605,N_13408,N_14448);
xor U16606 (N_16606,N_13439,N_12813);
nand U16607 (N_16607,N_14248,N_13939);
and U16608 (N_16608,N_14377,N_14671);
or U16609 (N_16609,N_14637,N_12686);
xor U16610 (N_16610,N_13014,N_12784);
or U16611 (N_16611,N_14559,N_12714);
or U16612 (N_16612,N_13584,N_13045);
xnor U16613 (N_16613,N_15021,N_12690);
or U16614 (N_16614,N_15019,N_14717);
xor U16615 (N_16615,N_12810,N_13430);
nand U16616 (N_16616,N_12818,N_15265);
nand U16617 (N_16617,N_12855,N_14212);
and U16618 (N_16618,N_12907,N_12823);
nor U16619 (N_16619,N_15503,N_14598);
xor U16620 (N_16620,N_15018,N_13271);
or U16621 (N_16621,N_12700,N_13494);
and U16622 (N_16622,N_12762,N_13467);
xnor U16623 (N_16623,N_15443,N_14805);
nor U16624 (N_16624,N_12651,N_13896);
nor U16625 (N_16625,N_13278,N_14398);
nor U16626 (N_16626,N_13300,N_12634);
nand U16627 (N_16627,N_13464,N_14535);
nand U16628 (N_16628,N_13497,N_13130);
xor U16629 (N_16629,N_14901,N_15089);
or U16630 (N_16630,N_13363,N_12613);
or U16631 (N_16631,N_12972,N_12572);
xnor U16632 (N_16632,N_14877,N_14649);
xor U16633 (N_16633,N_15124,N_15109);
nand U16634 (N_16634,N_13525,N_14518);
xor U16635 (N_16635,N_12699,N_14729);
nor U16636 (N_16636,N_14812,N_12676);
nor U16637 (N_16637,N_14383,N_12656);
and U16638 (N_16638,N_13784,N_14600);
nor U16639 (N_16639,N_14241,N_15208);
nor U16640 (N_16640,N_14115,N_12660);
nand U16641 (N_16641,N_15582,N_13917);
or U16642 (N_16642,N_13768,N_12745);
or U16643 (N_16643,N_15319,N_15040);
xor U16644 (N_16644,N_13827,N_12595);
xor U16645 (N_16645,N_13859,N_14939);
or U16646 (N_16646,N_13304,N_15476);
xor U16647 (N_16647,N_14990,N_13043);
xnor U16648 (N_16648,N_13208,N_15351);
and U16649 (N_16649,N_13318,N_13749);
xor U16650 (N_16650,N_14504,N_14657);
xor U16651 (N_16651,N_13492,N_14472);
nor U16652 (N_16652,N_12912,N_13388);
nand U16653 (N_16653,N_15086,N_15034);
and U16654 (N_16654,N_14418,N_13032);
nor U16655 (N_16655,N_15277,N_12557);
or U16656 (N_16656,N_14462,N_14723);
nor U16657 (N_16657,N_15525,N_14929);
nor U16658 (N_16658,N_13092,N_14838);
nor U16659 (N_16659,N_15526,N_12956);
or U16660 (N_16660,N_13175,N_14290);
nor U16661 (N_16661,N_14607,N_14147);
nand U16662 (N_16662,N_12684,N_14776);
nor U16663 (N_16663,N_13153,N_14769);
xor U16664 (N_16664,N_15099,N_15387);
or U16665 (N_16665,N_12523,N_14995);
nor U16666 (N_16666,N_12701,N_13343);
or U16667 (N_16667,N_12717,N_13778);
xnor U16668 (N_16668,N_14817,N_13612);
nor U16669 (N_16669,N_14049,N_15189);
nand U16670 (N_16670,N_12539,N_15210);
or U16671 (N_16671,N_14999,N_13561);
or U16672 (N_16672,N_14601,N_15064);
or U16673 (N_16673,N_15271,N_14136);
xnor U16674 (N_16674,N_13719,N_15102);
or U16675 (N_16675,N_14519,N_15233);
and U16676 (N_16676,N_13356,N_13315);
xnor U16677 (N_16677,N_13996,N_13174);
xor U16678 (N_16678,N_13042,N_13834);
nor U16679 (N_16679,N_14209,N_14743);
nor U16680 (N_16680,N_14707,N_14415);
nor U16681 (N_16681,N_14997,N_15334);
nor U16682 (N_16682,N_15273,N_13571);
or U16683 (N_16683,N_14186,N_15168);
and U16684 (N_16684,N_15084,N_13863);
or U16685 (N_16685,N_14088,N_14511);
or U16686 (N_16686,N_15514,N_14485);
nand U16687 (N_16687,N_15201,N_13819);
and U16688 (N_16688,N_14695,N_13468);
and U16689 (N_16689,N_15466,N_14837);
xor U16690 (N_16690,N_12643,N_13488);
nor U16691 (N_16691,N_13390,N_12565);
nand U16692 (N_16692,N_14040,N_13582);
or U16693 (N_16693,N_15556,N_13299);
or U16694 (N_16694,N_14744,N_15050);
nor U16695 (N_16695,N_13487,N_14099);
or U16696 (N_16696,N_14532,N_13686);
xnor U16697 (N_16697,N_14912,N_12650);
nor U16698 (N_16698,N_15110,N_14797);
and U16699 (N_16699,N_14175,N_14926);
xnor U16700 (N_16700,N_12509,N_13765);
nand U16701 (N_16701,N_15288,N_14678);
and U16702 (N_16702,N_13613,N_14266);
nand U16703 (N_16703,N_13370,N_15389);
nand U16704 (N_16704,N_14525,N_15624);
xor U16705 (N_16705,N_12611,N_13191);
xor U16706 (N_16706,N_12988,N_13736);
and U16707 (N_16707,N_15038,N_15198);
or U16708 (N_16708,N_14541,N_15107);
xnor U16709 (N_16709,N_13903,N_14828);
and U16710 (N_16710,N_12635,N_14892);
or U16711 (N_16711,N_14283,N_13411);
or U16712 (N_16712,N_14746,N_12764);
xnor U16713 (N_16713,N_13581,N_13685);
or U16714 (N_16714,N_14215,N_15003);
and U16715 (N_16715,N_13830,N_14585);
and U16716 (N_16716,N_13793,N_15618);
or U16717 (N_16717,N_15532,N_12966);
xor U16718 (N_16718,N_12755,N_14154);
nand U16719 (N_16719,N_13401,N_14898);
nand U16720 (N_16720,N_12776,N_15363);
nor U16721 (N_16721,N_13110,N_14235);
or U16722 (N_16722,N_13157,N_14942);
xnor U16723 (N_16723,N_12804,N_14168);
or U16724 (N_16724,N_15561,N_12606);
and U16725 (N_16725,N_12849,N_14023);
nor U16726 (N_16726,N_13140,N_13108);
xnor U16727 (N_16727,N_13030,N_14451);
nor U16728 (N_16728,N_14799,N_14135);
or U16729 (N_16729,N_14466,N_14163);
xor U16730 (N_16730,N_14866,N_12524);
and U16731 (N_16731,N_14514,N_14310);
xor U16732 (N_16732,N_15058,N_12564);
xnor U16733 (N_16733,N_14384,N_12891);
nand U16734 (N_16734,N_12727,N_13328);
xnor U16735 (N_16735,N_12953,N_12510);
nor U16736 (N_16736,N_15608,N_15054);
and U16737 (N_16737,N_15464,N_12505);
or U16738 (N_16738,N_14869,N_14760);
nor U16739 (N_16739,N_14013,N_14181);
nor U16740 (N_16740,N_15430,N_14849);
xnor U16741 (N_16741,N_15241,N_13182);
or U16742 (N_16742,N_14672,N_13224);
or U16743 (N_16743,N_15490,N_13499);
xnor U16744 (N_16744,N_13456,N_14626);
and U16745 (N_16745,N_14608,N_14727);
nand U16746 (N_16746,N_12506,N_15493);
or U16747 (N_16747,N_14335,N_15275);
xor U16748 (N_16748,N_15292,N_12949);
xor U16749 (N_16749,N_12922,N_14781);
and U16750 (N_16750,N_14325,N_15380);
or U16751 (N_16751,N_13125,N_14975);
nand U16752 (N_16752,N_14020,N_14112);
xnor U16753 (N_16753,N_12828,N_14001);
or U16754 (N_16754,N_13050,N_15301);
nor U16755 (N_16755,N_13142,N_14534);
xor U16756 (N_16756,N_14022,N_14424);
or U16757 (N_16757,N_13694,N_13672);
or U16758 (N_16758,N_13051,N_12678);
or U16759 (N_16759,N_14354,N_12639);
xor U16760 (N_16760,N_15256,N_12722);
nor U16761 (N_16761,N_13269,N_12887);
or U16762 (N_16762,N_13858,N_13160);
and U16763 (N_16763,N_14706,N_14264);
xnor U16764 (N_16764,N_14208,N_13981);
xor U16765 (N_16765,N_15194,N_12721);
nor U16766 (N_16766,N_13868,N_14187);
or U16767 (N_16767,N_14014,N_15047);
nand U16768 (N_16768,N_12788,N_15408);
or U16769 (N_16769,N_13604,N_13484);
nor U16770 (N_16770,N_13703,N_15228);
or U16771 (N_16771,N_14670,N_13424);
nor U16772 (N_16772,N_14298,N_14654);
and U16773 (N_16773,N_13848,N_15441);
xor U16774 (N_16774,N_13414,N_15323);
nand U16775 (N_16775,N_13173,N_13916);
and U16776 (N_16776,N_12589,N_12734);
xor U16777 (N_16777,N_13427,N_13061);
and U16778 (N_16778,N_14846,N_14676);
or U16779 (N_16779,N_13608,N_12857);
nand U16780 (N_16780,N_15161,N_12591);
and U16781 (N_16781,N_14378,N_15179);
nor U16782 (N_16782,N_14100,N_12558);
and U16783 (N_16783,N_13509,N_12748);
and U16784 (N_16784,N_14249,N_15258);
nor U16785 (N_16785,N_12706,N_14527);
or U16786 (N_16786,N_14425,N_15552);
nor U16787 (N_16787,N_14183,N_13754);
or U16788 (N_16788,N_13090,N_15249);
xor U16789 (N_16789,N_13970,N_13836);
and U16790 (N_16790,N_15013,N_12822);
nand U16791 (N_16791,N_15502,N_13627);
or U16792 (N_16792,N_12537,N_13237);
and U16793 (N_16793,N_12950,N_15290);
and U16794 (N_16794,N_13632,N_14333);
and U16795 (N_16795,N_12527,N_14991);
or U16796 (N_16796,N_15320,N_15601);
nand U16797 (N_16797,N_12944,N_14443);
xnor U16798 (N_16798,N_13617,N_13293);
and U16799 (N_16799,N_12604,N_13324);
nand U16800 (N_16800,N_14595,N_14612);
nor U16801 (N_16801,N_13587,N_14453);
or U16802 (N_16802,N_12795,N_14701);
nand U16803 (N_16803,N_14918,N_15360);
xnor U16804 (N_16804,N_13313,N_14313);
nor U16805 (N_16805,N_12851,N_12775);
nand U16806 (N_16806,N_13649,N_12957);
nor U16807 (N_16807,N_14031,N_13069);
or U16808 (N_16808,N_12544,N_12874);
and U16809 (N_16809,N_15358,N_14709);
and U16810 (N_16810,N_12936,N_14842);
or U16811 (N_16811,N_13098,N_13364);
or U16812 (N_16812,N_13505,N_15030);
nor U16813 (N_16813,N_15204,N_13236);
xor U16814 (N_16814,N_14503,N_12801);
xnor U16815 (N_16815,N_14327,N_14244);
nand U16816 (N_16816,N_14947,N_13077);
nand U16817 (N_16817,N_13567,N_12902);
and U16818 (N_16818,N_13197,N_13138);
and U16819 (N_16819,N_13253,N_13593);
nand U16820 (N_16820,N_12789,N_13785);
nand U16821 (N_16821,N_13693,N_15457);
nor U16822 (N_16822,N_14108,N_13955);
or U16823 (N_16823,N_14256,N_13927);
nor U16824 (N_16824,N_12603,N_13493);
or U16825 (N_16825,N_14782,N_14935);
nor U16826 (N_16826,N_14575,N_13486);
or U16827 (N_16827,N_14896,N_12647);
xnor U16828 (N_16828,N_14615,N_14931);
nor U16829 (N_16829,N_14655,N_15145);
nor U16830 (N_16830,N_13041,N_13852);
or U16831 (N_16831,N_13602,N_13217);
or U16832 (N_16832,N_15071,N_12820);
nand U16833 (N_16833,N_13522,N_13714);
or U16834 (N_16834,N_13684,N_14791);
and U16835 (N_16835,N_13773,N_12614);
xor U16836 (N_16836,N_14311,N_15353);
xnor U16837 (N_16837,N_13273,N_15376);
and U16838 (N_16838,N_14789,N_14751);
and U16839 (N_16839,N_15398,N_14024);
and U16840 (N_16840,N_15498,N_14801);
xnor U16841 (N_16841,N_14963,N_12768);
and U16842 (N_16842,N_14098,N_13811);
or U16843 (N_16843,N_14190,N_14510);
and U16844 (N_16844,N_13432,N_14474);
xnor U16845 (N_16845,N_13865,N_13479);
xor U16846 (N_16846,N_13129,N_13702);
nor U16847 (N_16847,N_13534,N_14675);
or U16848 (N_16848,N_13625,N_12623);
nand U16849 (N_16849,N_15421,N_15007);
and U16850 (N_16850,N_14293,N_13651);
nand U16851 (N_16851,N_13100,N_13994);
xnor U16852 (N_16852,N_15314,N_14291);
nand U16853 (N_16853,N_14994,N_15104);
nand U16854 (N_16854,N_13341,N_15451);
nor U16855 (N_16855,N_15115,N_14763);
and U16856 (N_16856,N_14833,N_15462);
xor U16857 (N_16857,N_15318,N_12553);
xnor U16858 (N_16858,N_12547,N_14095);
nor U16859 (N_16859,N_12786,N_13941);
or U16860 (N_16860,N_13692,N_12729);
or U16861 (N_16861,N_13239,N_13016);
or U16862 (N_16862,N_13659,N_13843);
nor U16863 (N_16863,N_12927,N_13054);
or U16864 (N_16864,N_13083,N_15604);
nand U16865 (N_16865,N_13842,N_15348);
nand U16866 (N_16866,N_15570,N_15599);
nand U16867 (N_16867,N_12548,N_12866);
nor U16868 (N_16868,N_13116,N_13592);
or U16869 (N_16869,N_13470,N_13876);
xor U16870 (N_16870,N_14275,N_14386);
nor U16871 (N_16871,N_14610,N_14521);
and U16872 (N_16872,N_13279,N_13209);
nand U16873 (N_16873,N_12612,N_15144);
xor U16874 (N_16874,N_14756,N_14957);
and U16875 (N_16875,N_13005,N_13618);
xor U16876 (N_16876,N_13755,N_14759);
nor U16877 (N_16877,N_13929,N_14762);
nand U16878 (N_16878,N_13751,N_15091);
and U16879 (N_16879,N_15368,N_14872);
nand U16880 (N_16880,N_15032,N_13115);
xor U16881 (N_16881,N_14389,N_13991);
or U16882 (N_16882,N_13392,N_13423);
nor U16883 (N_16883,N_15569,N_14934);
and U16884 (N_16884,N_15206,N_14652);
or U16885 (N_16885,N_12731,N_13808);
nand U16886 (N_16886,N_14796,N_15345);
or U16887 (N_16887,N_12607,N_12742);
xor U16888 (N_16888,N_15511,N_13365);
nor U16889 (N_16889,N_15056,N_13101);
xor U16890 (N_16890,N_15549,N_13213);
xor U16891 (N_16891,N_13697,N_13038);
xnor U16892 (N_16892,N_12947,N_15480);
or U16893 (N_16893,N_12834,N_15044);
and U16894 (N_16894,N_14117,N_13008);
nand U16895 (N_16895,N_12695,N_14568);
xor U16896 (N_16896,N_14231,N_14435);
xnor U16897 (N_16897,N_15082,N_14766);
nor U16898 (N_16898,N_14344,N_14006);
and U16899 (N_16899,N_15122,N_15367);
nand U16900 (N_16900,N_14433,N_12674);
and U16901 (N_16901,N_15251,N_13052);
xor U16902 (N_16902,N_12642,N_13701);
and U16903 (N_16903,N_13068,N_14358);
and U16904 (N_16904,N_15483,N_15260);
xnor U16905 (N_16905,N_12877,N_14427);
nand U16906 (N_16906,N_14370,N_14084);
xnor U16907 (N_16907,N_13576,N_14881);
xnor U16908 (N_16908,N_13934,N_13946);
and U16909 (N_16909,N_13457,N_15215);
xor U16910 (N_16910,N_13775,N_15544);
xor U16911 (N_16911,N_13740,N_13316);
or U16912 (N_16912,N_14822,N_14051);
nor U16913 (N_16913,N_12759,N_13029);
nand U16914 (N_16914,N_14106,N_15037);
nor U16915 (N_16915,N_13096,N_14262);
nand U16916 (N_16916,N_15440,N_14406);
nor U16917 (N_16917,N_15188,N_13904);
or U16918 (N_16918,N_13959,N_15069);
or U16919 (N_16919,N_15327,N_13553);
nand U16920 (N_16920,N_15422,N_12535);
and U16921 (N_16921,N_14011,N_14512);
nor U16922 (N_16922,N_12704,N_13989);
and U16923 (N_16923,N_14419,N_14571);
xor U16924 (N_16924,N_15567,N_14261);
xor U16925 (N_16925,N_12794,N_13718);
and U16926 (N_16926,N_14547,N_12723);
and U16927 (N_16927,N_13898,N_14708);
nand U16928 (N_16928,N_14050,N_14363);
xnor U16929 (N_16929,N_12584,N_14188);
or U16930 (N_16930,N_15383,N_13856);
or U16931 (N_16931,N_12893,N_13841);
xor U16932 (N_16932,N_12920,N_14659);
xnor U16933 (N_16933,N_15517,N_13170);
nor U16934 (N_16934,N_14459,N_13338);
nand U16935 (N_16935,N_14859,N_13899);
xnor U16936 (N_16936,N_14238,N_12832);
xnor U16937 (N_16937,N_13301,N_13187);
xnor U16938 (N_16938,N_14588,N_13845);
nor U16939 (N_16939,N_14134,N_13475);
and U16940 (N_16940,N_13881,N_14397);
nor U16941 (N_16941,N_12577,N_14493);
nor U16942 (N_16942,N_13244,N_15378);
nand U16943 (N_16943,N_13274,N_13716);
and U16944 (N_16944,N_14808,N_13974);
xnor U16945 (N_16945,N_12571,N_15170);
and U16946 (N_16946,N_14306,N_13240);
nand U16947 (N_16947,N_14287,N_14403);
nor U16948 (N_16948,N_13804,N_15070);
and U16949 (N_16949,N_14219,N_14417);
or U16950 (N_16950,N_14604,N_13281);
or U16951 (N_16951,N_14967,N_14077);
xnor U16952 (N_16952,N_15610,N_12569);
or U16953 (N_16953,N_12712,N_14758);
nand U16954 (N_16954,N_15536,N_15472);
xor U16955 (N_16955,N_14229,N_13535);
nand U16956 (N_16956,N_15455,N_12895);
and U16957 (N_16957,N_12765,N_13062);
or U16958 (N_16958,N_12725,N_13040);
nor U16959 (N_16959,N_15405,N_14883);
nor U16960 (N_16960,N_15529,N_13726);
xor U16961 (N_16961,N_13071,N_14372);
and U16962 (N_16962,N_13727,N_14360);
or U16963 (N_16963,N_15307,N_14924);
xor U16964 (N_16964,N_13995,N_13733);
or U16965 (N_16965,N_13764,N_12617);
nand U16966 (N_16966,N_12997,N_13931);
nor U16967 (N_16967,N_15236,N_14697);
and U16968 (N_16968,N_13001,N_15136);
xor U16969 (N_16969,N_14908,N_14992);
or U16970 (N_16970,N_15406,N_14353);
nand U16971 (N_16971,N_15447,N_12520);
nor U16972 (N_16972,N_14140,N_15120);
or U16973 (N_16973,N_12683,N_13089);
xnor U16974 (N_16974,N_14733,N_13621);
or U16975 (N_16975,N_12841,N_15244);
and U16976 (N_16976,N_13840,N_12905);
nor U16977 (N_16977,N_13366,N_15326);
nand U16978 (N_16978,N_14544,N_14738);
or U16979 (N_16979,N_13074,N_13282);
nand U16980 (N_16980,N_14412,N_13636);
xnor U16981 (N_16981,N_14428,N_14258);
xnor U16982 (N_16982,N_14906,N_13169);
and U16983 (N_16983,N_15587,N_12984);
nor U16984 (N_16984,N_14847,N_13373);
nand U16985 (N_16985,N_15374,N_13912);
or U16986 (N_16986,N_14668,N_13438);
nand U16987 (N_16987,N_15199,N_13447);
xor U16988 (N_16988,N_13152,N_14922);
and U16989 (N_16989,N_12772,N_14925);
and U16990 (N_16990,N_13190,N_13333);
nor U16991 (N_16991,N_15619,N_14060);
nand U16992 (N_16992,N_14853,N_13472);
nor U16993 (N_16993,N_14308,N_13019);
nand U16994 (N_16994,N_14804,N_13810);
nor U16995 (N_16995,N_13529,N_14516);
or U16996 (N_16996,N_13678,N_12518);
nor U16997 (N_16997,N_14338,N_14681);
xnor U16998 (N_16998,N_12996,N_15269);
or U16999 (N_16999,N_15335,N_13962);
xnor U17000 (N_17000,N_13489,N_12716);
nand U17001 (N_17001,N_12713,N_14640);
nor U17002 (N_17002,N_14068,N_14018);
nor U17003 (N_17003,N_14581,N_14567);
or U17004 (N_17004,N_14688,N_14823);
or U17005 (N_17005,N_14057,N_14488);
nand U17006 (N_17006,N_13980,N_14944);
nand U17007 (N_17007,N_13126,N_14686);
xnor U17008 (N_17008,N_14110,N_14257);
nor U17009 (N_17009,N_14144,N_12797);
or U17010 (N_17010,N_14391,N_12774);
xnor U17011 (N_17011,N_13879,N_12901);
or U17012 (N_17012,N_13193,N_13413);
xnor U17013 (N_17013,N_13163,N_14387);
or U17014 (N_17014,N_12815,N_13821);
or U17015 (N_17015,N_15280,N_14811);
nand U17016 (N_17016,N_14030,N_15492);
or U17017 (N_17017,N_13132,N_13533);
xor U17018 (N_17018,N_13094,N_15595);
or U17019 (N_17019,N_14956,N_13557);
or U17020 (N_17020,N_13225,N_12837);
and U17021 (N_17021,N_12883,N_15266);
and U17022 (N_17022,N_14346,N_13398);
xor U17023 (N_17023,N_14679,N_13435);
nor U17024 (N_17024,N_14227,N_13936);
and U17025 (N_17025,N_14876,N_15482);
xnor U17026 (N_17026,N_14478,N_12636);
and U17027 (N_17027,N_15267,N_14537);
and U17028 (N_17028,N_13319,N_15598);
and U17029 (N_17029,N_12924,N_15020);
and U17030 (N_17030,N_15196,N_15579);
or U17031 (N_17031,N_13261,N_12968);
nor U17032 (N_17032,N_13960,N_15061);
xnor U17033 (N_17033,N_14426,N_14800);
xor U17034 (N_17034,N_14964,N_12781);
and U17035 (N_17035,N_15149,N_15432);
xnor U17036 (N_17036,N_15468,N_13292);
and U17037 (N_17037,N_13978,N_14035);
xor U17038 (N_17038,N_13220,N_14777);
xor U17039 (N_17039,N_14642,N_15087);
nand U17040 (N_17040,N_12978,N_13476);
xor U17041 (N_17041,N_15252,N_14164);
nand U17042 (N_17042,N_13047,N_12791);
xor U17043 (N_17043,N_14565,N_15139);
xor U17044 (N_17044,N_13747,N_14524);
nor U17045 (N_17045,N_12990,N_15308);
or U17046 (N_17046,N_15393,N_13166);
or U17047 (N_17047,N_15475,N_13164);
and U17048 (N_17048,N_15279,N_14953);
xnor U17049 (N_17049,N_13146,N_15359);
or U17050 (N_17050,N_15509,N_14461);
or U17051 (N_17051,N_14385,N_15276);
nor U17052 (N_17052,N_14862,N_13387);
nand U17053 (N_17053,N_14522,N_14868);
and U17054 (N_17054,N_15609,N_14454);
nand U17055 (N_17055,N_15303,N_15519);
xor U17056 (N_17056,N_15520,N_13642);
xor U17057 (N_17057,N_13788,N_15254);
xnor U17058 (N_17058,N_13809,N_14277);
and U17059 (N_17059,N_13434,N_14538);
nand U17060 (N_17060,N_13905,N_13466);
nand U17061 (N_17061,N_15259,N_13766);
nor U17062 (N_17062,N_14319,N_12710);
xnor U17063 (N_17063,N_14089,N_12670);
xor U17064 (N_17064,N_13444,N_15404);
nand U17065 (N_17065,N_13579,N_14945);
nand U17066 (N_17066,N_13275,N_13812);
nor U17067 (N_17067,N_14714,N_13247);
nand U17068 (N_17068,N_13407,N_14492);
nand U17069 (N_17069,N_13975,N_13103);
nor U17070 (N_17070,N_12975,N_13873);
nand U17071 (N_17071,N_15048,N_14560);
nor U17072 (N_17072,N_14653,N_14465);
and U17073 (N_17073,N_14300,N_13832);
nand U17074 (N_17074,N_14860,N_12677);
or U17075 (N_17075,N_14430,N_15540);
or U17076 (N_17076,N_15369,N_15594);
nor U17077 (N_17077,N_14203,N_13037);
or U17078 (N_17078,N_14193,N_15403);
nand U17079 (N_17079,N_13091,N_14464);
and U17080 (N_17080,N_13323,N_13861);
or U17081 (N_17081,N_15112,N_12845);
nand U17082 (N_17082,N_12885,N_13327);
nand U17083 (N_17083,N_15433,N_14255);
or U17084 (N_17084,N_13150,N_15484);
xor U17085 (N_17085,N_15127,N_14768);
xnor U17086 (N_17086,N_14342,N_15324);
and U17087 (N_17087,N_14043,N_15137);
nand U17088 (N_17088,N_12766,N_14444);
or U17089 (N_17089,N_14160,N_13779);
and U17090 (N_17090,N_13671,N_12708);
or U17091 (N_17091,N_12951,N_13302);
or U17092 (N_17092,N_12980,N_13346);
nor U17093 (N_17093,N_14315,N_13911);
nand U17094 (N_17094,N_14761,N_13641);
nor U17095 (N_17095,N_13874,N_13598);
or U17096 (N_17096,N_12836,N_15346);
or U17097 (N_17097,N_15384,N_15004);
or U17098 (N_17098,N_15165,N_15444);
nor U17099 (N_17099,N_13256,N_14489);
xor U17100 (N_17100,N_15485,N_13619);
and U17101 (N_17101,N_12688,N_13648);
xor U17102 (N_17102,N_14130,N_15108);
and U17103 (N_17103,N_13610,N_14978);
nand U17104 (N_17104,N_14394,N_14482);
or U17105 (N_17105,N_14314,N_13791);
or U17106 (N_17106,N_14593,N_13442);
nor U17107 (N_17107,N_12886,N_14416);
nand U17108 (N_17108,N_14561,N_12829);
nor U17109 (N_17109,N_13707,N_14491);
nor U17110 (N_17110,N_14983,N_15611);
and U17111 (N_17111,N_14539,N_15310);
nor U17112 (N_17112,N_12803,N_15094);
xnor U17113 (N_17113,N_14562,N_13952);
or U17114 (N_17114,N_13513,N_12530);
xnor U17115 (N_17115,N_15163,N_13179);
or U17116 (N_17116,N_13713,N_13031);
nor U17117 (N_17117,N_14752,N_13056);
nand U17118 (N_17118,N_14081,N_14118);
nor U17119 (N_17119,N_14189,N_14250);
nor U17120 (N_17120,N_12592,N_12561);
and U17121 (N_17121,N_13481,N_15572);
nand U17122 (N_17122,N_15197,N_15062);
and U17123 (N_17123,N_15605,N_14141);
xnor U17124 (N_17124,N_13064,N_13495);
xor U17125 (N_17125,N_12793,N_12827);
and U17126 (N_17126,N_14515,N_14286);
and U17127 (N_17127,N_14580,N_15026);
or U17128 (N_17128,N_13243,N_15560);
and U17129 (N_17129,N_12969,N_12761);
nor U17130 (N_17130,N_13967,N_14960);
nor U17131 (N_17131,N_15431,N_12632);
nor U17132 (N_17132,N_15185,N_14074);
and U17133 (N_17133,N_13283,N_14066);
nor U17134 (N_17134,N_12532,N_13615);
and U17135 (N_17135,N_13194,N_15500);
and U17136 (N_17136,N_14126,N_15294);
xor U17137 (N_17137,N_15377,N_13710);
nor U17138 (N_17138,N_14486,N_13596);
xor U17139 (N_17139,N_15336,N_12507);
or U17140 (N_17140,N_14660,N_13933);
nor U17141 (N_17141,N_12825,N_14894);
nor U17142 (N_17142,N_15297,N_13426);
and U17143 (N_17143,N_13322,N_12582);
or U17144 (N_17144,N_14528,N_14703);
nand U17145 (N_17145,N_15160,N_14584);
and U17146 (N_17146,N_13984,N_13079);
and U17147 (N_17147,N_15331,N_13572);
xnor U17148 (N_17148,N_12929,N_15461);
nand U17149 (N_17149,N_14441,N_13264);
or U17150 (N_17150,N_13291,N_13944);
or U17151 (N_17151,N_15491,N_15081);
nand U17152 (N_17152,N_15295,N_15527);
xor U17153 (N_17153,N_12533,N_13752);
and U17154 (N_17154,N_13053,N_12551);
nand U17155 (N_17155,N_12999,N_13913);
and U17156 (N_17156,N_14137,N_14331);
nor U17157 (N_17157,N_14885,N_13353);
xnor U17158 (N_17158,N_13216,N_15130);
xor U17159 (N_17159,N_15164,N_15008);
nand U17160 (N_17160,N_14895,N_14624);
and U17161 (N_17161,N_13661,N_14982);
xnor U17162 (N_17162,N_13683,N_14149);
nand U17163 (N_17163,N_13928,N_13894);
nand U17164 (N_17164,N_13235,N_13735);
xor U17165 (N_17165,N_15499,N_13474);
nand U17166 (N_17166,N_13336,N_15362);
and U17167 (N_17167,N_13419,N_14840);
and U17168 (N_17168,N_14589,N_15153);
or U17169 (N_17169,N_13342,N_13097);
nor U17170 (N_17170,N_14449,N_13857);
and U17171 (N_17171,N_13822,N_15205);
nor U17172 (N_17172,N_14788,N_13560);
nor U17173 (N_17173,N_13351,N_14878);
nand U17174 (N_17174,N_13826,N_15078);
nor U17175 (N_17175,N_14973,N_15079);
and U17176 (N_17176,N_12780,N_13796);
xnor U17177 (N_17177,N_12961,N_14000);
xor U17178 (N_17178,N_13644,N_13227);
nand U17179 (N_17179,N_13676,N_15365);
nor U17180 (N_17180,N_12653,N_14592);
and U17181 (N_17181,N_13790,N_15448);
xor U17182 (N_17182,N_14131,N_14779);
and U17183 (N_17183,N_14033,N_14841);
nand U17184 (N_17184,N_12559,N_15592);
nand U17185 (N_17185,N_13245,N_13756);
nand U17186 (N_17186,N_13997,N_12529);
nor U17187 (N_17187,N_13024,N_14966);
xnor U17188 (N_17188,N_14803,N_12874);
and U17189 (N_17189,N_13087,N_14047);
and U17190 (N_17190,N_14957,N_15363);
xnor U17191 (N_17191,N_13497,N_14404);
or U17192 (N_17192,N_15352,N_15256);
nand U17193 (N_17193,N_13389,N_13459);
and U17194 (N_17194,N_13134,N_14511);
and U17195 (N_17195,N_12549,N_15467);
or U17196 (N_17196,N_14473,N_14833);
and U17197 (N_17197,N_12839,N_13542);
or U17198 (N_17198,N_14759,N_14331);
or U17199 (N_17199,N_13919,N_13336);
nand U17200 (N_17200,N_14320,N_14064);
nand U17201 (N_17201,N_12715,N_14226);
xor U17202 (N_17202,N_14252,N_14894);
and U17203 (N_17203,N_15372,N_14254);
nor U17204 (N_17204,N_13794,N_14232);
or U17205 (N_17205,N_13180,N_15593);
nor U17206 (N_17206,N_15340,N_14815);
xor U17207 (N_17207,N_13624,N_14713);
xnor U17208 (N_17208,N_14010,N_12751);
nand U17209 (N_17209,N_12982,N_12806);
and U17210 (N_17210,N_13170,N_12946);
and U17211 (N_17211,N_13729,N_15589);
nor U17212 (N_17212,N_15457,N_13606);
xor U17213 (N_17213,N_14675,N_13130);
and U17214 (N_17214,N_12926,N_13920);
nand U17215 (N_17215,N_12684,N_13139);
and U17216 (N_17216,N_13208,N_13984);
nor U17217 (N_17217,N_13589,N_12936);
or U17218 (N_17218,N_12936,N_12781);
nand U17219 (N_17219,N_14992,N_13779);
or U17220 (N_17220,N_14599,N_14447);
nand U17221 (N_17221,N_12946,N_13302);
xor U17222 (N_17222,N_13986,N_14008);
or U17223 (N_17223,N_15130,N_12809);
or U17224 (N_17224,N_13379,N_15014);
xor U17225 (N_17225,N_14761,N_14635);
nand U17226 (N_17226,N_14091,N_13659);
nand U17227 (N_17227,N_15391,N_13425);
nor U17228 (N_17228,N_14743,N_13069);
nor U17229 (N_17229,N_15086,N_14004);
nor U17230 (N_17230,N_14331,N_15392);
nand U17231 (N_17231,N_14532,N_13896);
nor U17232 (N_17232,N_13352,N_12549);
nor U17233 (N_17233,N_13348,N_13669);
and U17234 (N_17234,N_13459,N_13363);
xnor U17235 (N_17235,N_15142,N_12952);
nand U17236 (N_17236,N_12750,N_15242);
nand U17237 (N_17237,N_15307,N_14053);
nand U17238 (N_17238,N_15070,N_14796);
xor U17239 (N_17239,N_13408,N_14531);
nor U17240 (N_17240,N_13797,N_13393);
and U17241 (N_17241,N_13811,N_14604);
nor U17242 (N_17242,N_12964,N_15395);
nand U17243 (N_17243,N_13145,N_12665);
nand U17244 (N_17244,N_14173,N_13544);
nand U17245 (N_17245,N_13531,N_14717);
or U17246 (N_17246,N_12706,N_12961);
nand U17247 (N_17247,N_12837,N_15475);
xor U17248 (N_17248,N_12633,N_14506);
and U17249 (N_17249,N_14127,N_12890);
and U17250 (N_17250,N_13590,N_13679);
xor U17251 (N_17251,N_14737,N_13217);
and U17252 (N_17252,N_14965,N_15580);
nand U17253 (N_17253,N_13307,N_13857);
xor U17254 (N_17254,N_15404,N_13060);
xnor U17255 (N_17255,N_14925,N_14215);
xor U17256 (N_17256,N_13438,N_12547);
and U17257 (N_17257,N_14708,N_14348);
nand U17258 (N_17258,N_14124,N_13709);
and U17259 (N_17259,N_14159,N_15206);
or U17260 (N_17260,N_14364,N_13305);
or U17261 (N_17261,N_14858,N_14753);
xor U17262 (N_17262,N_13593,N_13664);
or U17263 (N_17263,N_14087,N_14580);
and U17264 (N_17264,N_15114,N_14712);
nor U17265 (N_17265,N_13324,N_13201);
xnor U17266 (N_17266,N_12751,N_13341);
nand U17267 (N_17267,N_13025,N_13155);
and U17268 (N_17268,N_14631,N_15302);
nor U17269 (N_17269,N_12891,N_13786);
and U17270 (N_17270,N_14910,N_12856);
nand U17271 (N_17271,N_15493,N_14810);
xor U17272 (N_17272,N_13150,N_13152);
and U17273 (N_17273,N_14150,N_12737);
or U17274 (N_17274,N_14667,N_12975);
nor U17275 (N_17275,N_15102,N_14573);
or U17276 (N_17276,N_14707,N_15573);
and U17277 (N_17277,N_13744,N_14282);
or U17278 (N_17278,N_13990,N_12891);
nor U17279 (N_17279,N_12895,N_14068);
or U17280 (N_17280,N_13367,N_13262);
xnor U17281 (N_17281,N_14573,N_14556);
or U17282 (N_17282,N_13771,N_14126);
nand U17283 (N_17283,N_14847,N_12849);
nor U17284 (N_17284,N_14983,N_14539);
or U17285 (N_17285,N_14567,N_13501);
and U17286 (N_17286,N_14546,N_14196);
nand U17287 (N_17287,N_14830,N_13051);
xnor U17288 (N_17288,N_12973,N_15396);
xnor U17289 (N_17289,N_14529,N_14755);
xnor U17290 (N_17290,N_15157,N_14769);
and U17291 (N_17291,N_14645,N_13151);
nand U17292 (N_17292,N_12822,N_13268);
xnor U17293 (N_17293,N_14571,N_13316);
nor U17294 (N_17294,N_15612,N_15525);
and U17295 (N_17295,N_15358,N_15106);
nand U17296 (N_17296,N_13897,N_13249);
nor U17297 (N_17297,N_13446,N_15103);
and U17298 (N_17298,N_14196,N_14755);
xor U17299 (N_17299,N_13288,N_13268);
nand U17300 (N_17300,N_15325,N_15594);
xor U17301 (N_17301,N_12817,N_13455);
or U17302 (N_17302,N_14525,N_14642);
nor U17303 (N_17303,N_14112,N_15227);
xnor U17304 (N_17304,N_15359,N_13634);
or U17305 (N_17305,N_14800,N_15290);
or U17306 (N_17306,N_14556,N_15483);
nor U17307 (N_17307,N_12582,N_14388);
nand U17308 (N_17308,N_12673,N_13244);
nor U17309 (N_17309,N_15538,N_14610);
nor U17310 (N_17310,N_12722,N_12709);
nand U17311 (N_17311,N_14435,N_14322);
nand U17312 (N_17312,N_14959,N_14554);
nand U17313 (N_17313,N_14748,N_15162);
nor U17314 (N_17314,N_15318,N_13723);
or U17315 (N_17315,N_13022,N_14931);
nand U17316 (N_17316,N_13802,N_12832);
nand U17317 (N_17317,N_14797,N_14096);
and U17318 (N_17318,N_13317,N_14020);
or U17319 (N_17319,N_13141,N_12773);
or U17320 (N_17320,N_13862,N_13517);
nor U17321 (N_17321,N_13416,N_15563);
and U17322 (N_17322,N_13339,N_12853);
nor U17323 (N_17323,N_13863,N_13722);
nand U17324 (N_17324,N_13794,N_13044);
nor U17325 (N_17325,N_13358,N_13859);
nor U17326 (N_17326,N_15597,N_15465);
nor U17327 (N_17327,N_13972,N_13762);
xnor U17328 (N_17328,N_13793,N_15376);
nand U17329 (N_17329,N_12524,N_13479);
nor U17330 (N_17330,N_14361,N_12718);
or U17331 (N_17331,N_14529,N_14939);
and U17332 (N_17332,N_13724,N_14144);
or U17333 (N_17333,N_12752,N_13948);
and U17334 (N_17334,N_12793,N_15054);
or U17335 (N_17335,N_12789,N_12685);
or U17336 (N_17336,N_14791,N_14043);
and U17337 (N_17337,N_15165,N_15511);
or U17338 (N_17338,N_13732,N_14576);
and U17339 (N_17339,N_15334,N_14812);
and U17340 (N_17340,N_13518,N_13540);
nand U17341 (N_17341,N_15443,N_14148);
nor U17342 (N_17342,N_15210,N_13821);
nand U17343 (N_17343,N_13560,N_14991);
xnor U17344 (N_17344,N_15128,N_13839);
and U17345 (N_17345,N_12625,N_14701);
or U17346 (N_17346,N_14495,N_12870);
nor U17347 (N_17347,N_15247,N_15535);
or U17348 (N_17348,N_14925,N_15168);
nand U17349 (N_17349,N_14790,N_12742);
and U17350 (N_17350,N_15235,N_12920);
nand U17351 (N_17351,N_12667,N_15346);
xor U17352 (N_17352,N_13451,N_14414);
xnor U17353 (N_17353,N_14131,N_12691);
xnor U17354 (N_17354,N_13459,N_12879);
nor U17355 (N_17355,N_15360,N_14515);
or U17356 (N_17356,N_14761,N_14938);
and U17357 (N_17357,N_13523,N_12978);
or U17358 (N_17358,N_13652,N_13554);
nor U17359 (N_17359,N_14910,N_13546);
or U17360 (N_17360,N_14194,N_12863);
or U17361 (N_17361,N_14122,N_13789);
and U17362 (N_17362,N_13550,N_15120);
nand U17363 (N_17363,N_13390,N_14305);
and U17364 (N_17364,N_13980,N_13114);
and U17365 (N_17365,N_13312,N_12860);
nand U17366 (N_17366,N_14971,N_14218);
xnor U17367 (N_17367,N_13399,N_12916);
nor U17368 (N_17368,N_12716,N_12677);
nor U17369 (N_17369,N_15361,N_13128);
nand U17370 (N_17370,N_12687,N_12788);
nand U17371 (N_17371,N_15576,N_13094);
nand U17372 (N_17372,N_13357,N_13636);
xnor U17373 (N_17373,N_14235,N_14207);
or U17374 (N_17374,N_13068,N_13476);
or U17375 (N_17375,N_13002,N_13028);
nor U17376 (N_17376,N_14626,N_13500);
nor U17377 (N_17377,N_14394,N_13692);
nand U17378 (N_17378,N_12907,N_15525);
nand U17379 (N_17379,N_14446,N_12586);
or U17380 (N_17380,N_13067,N_15055);
nand U17381 (N_17381,N_14257,N_15307);
nor U17382 (N_17382,N_12502,N_12609);
nor U17383 (N_17383,N_15107,N_12668);
nor U17384 (N_17384,N_15396,N_14534);
xor U17385 (N_17385,N_14288,N_13695);
nand U17386 (N_17386,N_12726,N_14545);
xor U17387 (N_17387,N_14036,N_13910);
xnor U17388 (N_17388,N_13115,N_15051);
nand U17389 (N_17389,N_13923,N_13048);
and U17390 (N_17390,N_13808,N_14087);
and U17391 (N_17391,N_13155,N_14741);
xnor U17392 (N_17392,N_15164,N_14687);
and U17393 (N_17393,N_13189,N_13341);
xor U17394 (N_17394,N_12665,N_13127);
nor U17395 (N_17395,N_14193,N_14111);
nand U17396 (N_17396,N_13787,N_12578);
xor U17397 (N_17397,N_13482,N_13014);
nor U17398 (N_17398,N_14846,N_12729);
nand U17399 (N_17399,N_13415,N_14711);
and U17400 (N_17400,N_13649,N_14330);
nor U17401 (N_17401,N_14526,N_15275);
xnor U17402 (N_17402,N_13220,N_14822);
or U17403 (N_17403,N_14832,N_14588);
nor U17404 (N_17404,N_14906,N_13660);
nor U17405 (N_17405,N_13475,N_14803);
nor U17406 (N_17406,N_15158,N_14253);
nand U17407 (N_17407,N_12868,N_12593);
xnor U17408 (N_17408,N_13482,N_13679);
nand U17409 (N_17409,N_12978,N_15473);
nor U17410 (N_17410,N_13713,N_12598);
nor U17411 (N_17411,N_15260,N_14565);
nor U17412 (N_17412,N_15539,N_12573);
nand U17413 (N_17413,N_14587,N_14104);
nor U17414 (N_17414,N_13456,N_14668);
xnor U17415 (N_17415,N_12684,N_12555);
or U17416 (N_17416,N_14795,N_13460);
and U17417 (N_17417,N_13434,N_13446);
xor U17418 (N_17418,N_14863,N_12742);
nor U17419 (N_17419,N_13470,N_14725);
nand U17420 (N_17420,N_13495,N_14535);
or U17421 (N_17421,N_15027,N_13232);
nand U17422 (N_17422,N_14654,N_13004);
and U17423 (N_17423,N_13711,N_15401);
and U17424 (N_17424,N_13222,N_12882);
nand U17425 (N_17425,N_15586,N_15422);
and U17426 (N_17426,N_15464,N_13644);
and U17427 (N_17427,N_13179,N_13974);
nor U17428 (N_17428,N_12856,N_15328);
nor U17429 (N_17429,N_12545,N_15549);
or U17430 (N_17430,N_13777,N_15405);
nor U17431 (N_17431,N_15089,N_15257);
nor U17432 (N_17432,N_13339,N_12808);
nor U17433 (N_17433,N_12953,N_14317);
nand U17434 (N_17434,N_14864,N_13048);
and U17435 (N_17435,N_15504,N_14316);
and U17436 (N_17436,N_12531,N_13518);
nand U17437 (N_17437,N_12850,N_15120);
nand U17438 (N_17438,N_15006,N_15605);
and U17439 (N_17439,N_14920,N_13678);
and U17440 (N_17440,N_15092,N_13962);
or U17441 (N_17441,N_15315,N_14839);
xor U17442 (N_17442,N_13544,N_13253);
xnor U17443 (N_17443,N_14840,N_15169);
nor U17444 (N_17444,N_14401,N_13732);
nand U17445 (N_17445,N_14970,N_14437);
nor U17446 (N_17446,N_14221,N_12613);
and U17447 (N_17447,N_14273,N_15123);
nor U17448 (N_17448,N_13404,N_15166);
or U17449 (N_17449,N_12868,N_14640);
nor U17450 (N_17450,N_14042,N_14528);
xnor U17451 (N_17451,N_15285,N_14365);
nor U17452 (N_17452,N_13687,N_13856);
xor U17453 (N_17453,N_12771,N_13759);
and U17454 (N_17454,N_13005,N_13191);
and U17455 (N_17455,N_13471,N_13574);
and U17456 (N_17456,N_14409,N_12719);
nor U17457 (N_17457,N_13081,N_14157);
and U17458 (N_17458,N_14198,N_12869);
nand U17459 (N_17459,N_14311,N_13171);
or U17460 (N_17460,N_13224,N_14363);
nor U17461 (N_17461,N_14207,N_13236);
and U17462 (N_17462,N_15122,N_12925);
or U17463 (N_17463,N_14283,N_12732);
and U17464 (N_17464,N_15547,N_14197);
nor U17465 (N_17465,N_14867,N_12964);
xnor U17466 (N_17466,N_13537,N_13857);
or U17467 (N_17467,N_14111,N_13789);
nand U17468 (N_17468,N_14272,N_13130);
nor U17469 (N_17469,N_14041,N_14252);
and U17470 (N_17470,N_15615,N_15389);
nor U17471 (N_17471,N_15111,N_15426);
xor U17472 (N_17472,N_14118,N_13040);
or U17473 (N_17473,N_13637,N_14856);
nand U17474 (N_17474,N_14287,N_12934);
or U17475 (N_17475,N_14792,N_12952);
xnor U17476 (N_17476,N_13499,N_14389);
or U17477 (N_17477,N_13668,N_13940);
or U17478 (N_17478,N_12889,N_13355);
nor U17479 (N_17479,N_14130,N_13360);
or U17480 (N_17480,N_13803,N_13066);
nand U17481 (N_17481,N_13191,N_13592);
xnor U17482 (N_17482,N_14691,N_14957);
xnor U17483 (N_17483,N_12776,N_15500);
and U17484 (N_17484,N_15344,N_13713);
and U17485 (N_17485,N_13003,N_12686);
xor U17486 (N_17486,N_14191,N_14235);
xor U17487 (N_17487,N_12763,N_14107);
nand U17488 (N_17488,N_14656,N_13099);
xnor U17489 (N_17489,N_13833,N_12832);
nor U17490 (N_17490,N_13382,N_13505);
or U17491 (N_17491,N_15230,N_13519);
or U17492 (N_17492,N_15019,N_12551);
xor U17493 (N_17493,N_13488,N_15049);
nand U17494 (N_17494,N_15460,N_12995);
nor U17495 (N_17495,N_13919,N_14396);
and U17496 (N_17496,N_13573,N_12577);
nor U17497 (N_17497,N_14246,N_14801);
or U17498 (N_17498,N_14208,N_12790);
nand U17499 (N_17499,N_13988,N_14553);
and U17500 (N_17500,N_14701,N_14862);
xnor U17501 (N_17501,N_12740,N_15214);
and U17502 (N_17502,N_12771,N_12758);
or U17503 (N_17503,N_14407,N_15269);
or U17504 (N_17504,N_13498,N_13565);
nand U17505 (N_17505,N_12810,N_12893);
nand U17506 (N_17506,N_13776,N_14485);
and U17507 (N_17507,N_14192,N_15097);
or U17508 (N_17508,N_12923,N_14214);
or U17509 (N_17509,N_12690,N_12822);
xnor U17510 (N_17510,N_13453,N_14953);
xnor U17511 (N_17511,N_15130,N_13258);
nor U17512 (N_17512,N_13715,N_14803);
xor U17513 (N_17513,N_13573,N_13777);
and U17514 (N_17514,N_14307,N_14395);
and U17515 (N_17515,N_14908,N_13711);
and U17516 (N_17516,N_12934,N_13502);
and U17517 (N_17517,N_13158,N_12898);
or U17518 (N_17518,N_15101,N_14824);
and U17519 (N_17519,N_14615,N_15405);
and U17520 (N_17520,N_14185,N_14620);
nand U17521 (N_17521,N_14666,N_13408);
and U17522 (N_17522,N_13490,N_14348);
xnor U17523 (N_17523,N_12668,N_14336);
or U17524 (N_17524,N_12701,N_12944);
or U17525 (N_17525,N_12990,N_12822);
or U17526 (N_17526,N_14430,N_15240);
and U17527 (N_17527,N_15184,N_14705);
nor U17528 (N_17528,N_13275,N_14838);
nand U17529 (N_17529,N_13160,N_14463);
nor U17530 (N_17530,N_13126,N_14059);
xnor U17531 (N_17531,N_13862,N_15351);
xnor U17532 (N_17532,N_14349,N_14490);
nand U17533 (N_17533,N_14063,N_14449);
xor U17534 (N_17534,N_12743,N_15383);
and U17535 (N_17535,N_14676,N_14485);
and U17536 (N_17536,N_14403,N_13389);
and U17537 (N_17537,N_14044,N_14536);
and U17538 (N_17538,N_12891,N_14157);
and U17539 (N_17539,N_15480,N_14835);
or U17540 (N_17540,N_14088,N_13182);
nand U17541 (N_17541,N_13374,N_13473);
nand U17542 (N_17542,N_15460,N_12545);
nand U17543 (N_17543,N_13955,N_14553);
nor U17544 (N_17544,N_15425,N_13777);
xor U17545 (N_17545,N_12622,N_13005);
nor U17546 (N_17546,N_12633,N_14547);
and U17547 (N_17547,N_14222,N_14659);
or U17548 (N_17548,N_14492,N_14171);
and U17549 (N_17549,N_14273,N_12801);
and U17550 (N_17550,N_15108,N_13053);
xnor U17551 (N_17551,N_15528,N_12963);
and U17552 (N_17552,N_12910,N_13421);
nor U17553 (N_17553,N_13269,N_13783);
or U17554 (N_17554,N_15463,N_13451);
or U17555 (N_17555,N_13011,N_15380);
or U17556 (N_17556,N_14204,N_14170);
xnor U17557 (N_17557,N_12966,N_13248);
nor U17558 (N_17558,N_13218,N_15280);
and U17559 (N_17559,N_12796,N_14642);
nor U17560 (N_17560,N_15220,N_15287);
nand U17561 (N_17561,N_14908,N_14781);
or U17562 (N_17562,N_13198,N_14354);
nor U17563 (N_17563,N_12830,N_12793);
nor U17564 (N_17564,N_15343,N_14218);
and U17565 (N_17565,N_13139,N_15053);
and U17566 (N_17566,N_14779,N_14752);
and U17567 (N_17567,N_13048,N_13200);
nor U17568 (N_17568,N_13144,N_15567);
xor U17569 (N_17569,N_14125,N_13500);
xnor U17570 (N_17570,N_14940,N_14224);
nand U17571 (N_17571,N_15091,N_15039);
xor U17572 (N_17572,N_14832,N_13242);
nand U17573 (N_17573,N_15610,N_13936);
xor U17574 (N_17574,N_12852,N_13700);
or U17575 (N_17575,N_12991,N_14567);
or U17576 (N_17576,N_12869,N_13555);
and U17577 (N_17577,N_14650,N_15217);
or U17578 (N_17578,N_15017,N_13378);
and U17579 (N_17579,N_14542,N_13028);
nand U17580 (N_17580,N_12891,N_14170);
xnor U17581 (N_17581,N_13812,N_12593);
nor U17582 (N_17582,N_14266,N_15269);
xor U17583 (N_17583,N_14912,N_14572);
nor U17584 (N_17584,N_14365,N_12866);
nor U17585 (N_17585,N_15057,N_14621);
xor U17586 (N_17586,N_12548,N_15434);
and U17587 (N_17587,N_14695,N_15328);
or U17588 (N_17588,N_12824,N_15137);
nand U17589 (N_17589,N_13449,N_12805);
and U17590 (N_17590,N_13950,N_15385);
nand U17591 (N_17591,N_14527,N_15360);
xor U17592 (N_17592,N_12590,N_13613);
and U17593 (N_17593,N_12653,N_15122);
or U17594 (N_17594,N_15553,N_14281);
and U17595 (N_17595,N_13202,N_13467);
nand U17596 (N_17596,N_14277,N_15197);
xnor U17597 (N_17597,N_13781,N_13036);
nand U17598 (N_17598,N_15596,N_14631);
nor U17599 (N_17599,N_14390,N_14471);
nor U17600 (N_17600,N_13511,N_13213);
or U17601 (N_17601,N_14055,N_14117);
and U17602 (N_17602,N_14219,N_12825);
nor U17603 (N_17603,N_13697,N_15118);
nor U17604 (N_17604,N_15430,N_14218);
and U17605 (N_17605,N_13735,N_14147);
and U17606 (N_17606,N_14787,N_14296);
xor U17607 (N_17607,N_13217,N_15343);
or U17608 (N_17608,N_14783,N_15281);
xnor U17609 (N_17609,N_14823,N_13865);
nand U17610 (N_17610,N_15593,N_13507);
nand U17611 (N_17611,N_12797,N_13851);
and U17612 (N_17612,N_14643,N_14247);
nand U17613 (N_17613,N_14444,N_14890);
and U17614 (N_17614,N_15580,N_13962);
nand U17615 (N_17615,N_15271,N_15545);
xnor U17616 (N_17616,N_14827,N_15208);
or U17617 (N_17617,N_15349,N_14032);
xor U17618 (N_17618,N_14599,N_12987);
xnor U17619 (N_17619,N_13235,N_14264);
nand U17620 (N_17620,N_13123,N_13020);
nor U17621 (N_17621,N_15094,N_13252);
or U17622 (N_17622,N_14754,N_13681);
xor U17623 (N_17623,N_14420,N_13992);
xor U17624 (N_17624,N_15142,N_14276);
nand U17625 (N_17625,N_13087,N_12707);
or U17626 (N_17626,N_14501,N_12780);
nor U17627 (N_17627,N_15358,N_15318);
nand U17628 (N_17628,N_12943,N_14244);
nand U17629 (N_17629,N_15158,N_15312);
nand U17630 (N_17630,N_13627,N_13140);
nand U17631 (N_17631,N_12927,N_15055);
and U17632 (N_17632,N_13571,N_13970);
and U17633 (N_17633,N_13451,N_13020);
or U17634 (N_17634,N_14008,N_14392);
nor U17635 (N_17635,N_14957,N_13682);
nand U17636 (N_17636,N_14589,N_15559);
nand U17637 (N_17637,N_13471,N_14052);
or U17638 (N_17638,N_14599,N_12892);
xnor U17639 (N_17639,N_14953,N_15351);
xor U17640 (N_17640,N_13631,N_13005);
xnor U17641 (N_17641,N_14146,N_15243);
and U17642 (N_17642,N_15030,N_12871);
xor U17643 (N_17643,N_14767,N_13221);
and U17644 (N_17644,N_13961,N_12627);
or U17645 (N_17645,N_13122,N_13143);
or U17646 (N_17646,N_15369,N_12564);
nand U17647 (N_17647,N_13146,N_14059);
nor U17648 (N_17648,N_12988,N_13446);
or U17649 (N_17649,N_13452,N_15535);
xor U17650 (N_17650,N_13391,N_12758);
nand U17651 (N_17651,N_12612,N_13605);
nor U17652 (N_17652,N_13357,N_14143);
nand U17653 (N_17653,N_13627,N_14679);
or U17654 (N_17654,N_14903,N_14792);
xnor U17655 (N_17655,N_13219,N_13856);
xor U17656 (N_17656,N_13889,N_14002);
nand U17657 (N_17657,N_12884,N_12875);
nor U17658 (N_17658,N_13180,N_13544);
xnor U17659 (N_17659,N_15151,N_14658);
or U17660 (N_17660,N_13015,N_13510);
nor U17661 (N_17661,N_12825,N_13233);
xor U17662 (N_17662,N_13294,N_13880);
nor U17663 (N_17663,N_13220,N_14095);
nand U17664 (N_17664,N_15384,N_12757);
nand U17665 (N_17665,N_14127,N_14013);
xnor U17666 (N_17666,N_15538,N_14633);
nor U17667 (N_17667,N_12849,N_13926);
xnor U17668 (N_17668,N_13789,N_14961);
or U17669 (N_17669,N_14948,N_15564);
nand U17670 (N_17670,N_14702,N_14189);
nor U17671 (N_17671,N_14748,N_14660);
nor U17672 (N_17672,N_14820,N_13494);
nand U17673 (N_17673,N_15602,N_14313);
or U17674 (N_17674,N_14237,N_14736);
nand U17675 (N_17675,N_13179,N_14049);
nand U17676 (N_17676,N_14417,N_13677);
and U17677 (N_17677,N_14908,N_14574);
nor U17678 (N_17678,N_13571,N_15205);
or U17679 (N_17679,N_14818,N_12545);
xnor U17680 (N_17680,N_13203,N_14618);
and U17681 (N_17681,N_14533,N_15315);
and U17682 (N_17682,N_15521,N_14140);
and U17683 (N_17683,N_12735,N_12546);
or U17684 (N_17684,N_14245,N_14191);
or U17685 (N_17685,N_13593,N_14956);
or U17686 (N_17686,N_13438,N_12973);
xor U17687 (N_17687,N_15345,N_13052);
nand U17688 (N_17688,N_15448,N_14350);
or U17689 (N_17689,N_15002,N_13449);
nand U17690 (N_17690,N_12715,N_13190);
nand U17691 (N_17691,N_14748,N_14016);
nor U17692 (N_17692,N_15251,N_13687);
xnor U17693 (N_17693,N_14553,N_13979);
nand U17694 (N_17694,N_15272,N_14071);
and U17695 (N_17695,N_12616,N_15560);
nand U17696 (N_17696,N_15025,N_13366);
and U17697 (N_17697,N_13908,N_14694);
xor U17698 (N_17698,N_13724,N_14024);
and U17699 (N_17699,N_15619,N_15278);
xor U17700 (N_17700,N_12612,N_14268);
nand U17701 (N_17701,N_15464,N_13374);
nand U17702 (N_17702,N_15160,N_13713);
or U17703 (N_17703,N_14666,N_14879);
nor U17704 (N_17704,N_15367,N_13233);
nand U17705 (N_17705,N_13917,N_15334);
nand U17706 (N_17706,N_14764,N_13835);
nand U17707 (N_17707,N_14435,N_12915);
and U17708 (N_17708,N_13554,N_12833);
nor U17709 (N_17709,N_13845,N_14403);
nand U17710 (N_17710,N_13545,N_13386);
xor U17711 (N_17711,N_14182,N_13561);
xor U17712 (N_17712,N_14476,N_14025);
and U17713 (N_17713,N_14350,N_15581);
xnor U17714 (N_17714,N_15098,N_15064);
nand U17715 (N_17715,N_15457,N_12995);
or U17716 (N_17716,N_13238,N_12934);
or U17717 (N_17717,N_15579,N_12927);
xnor U17718 (N_17718,N_14609,N_13350);
xnor U17719 (N_17719,N_14013,N_13266);
or U17720 (N_17720,N_13055,N_14675);
and U17721 (N_17721,N_15136,N_14188);
nor U17722 (N_17722,N_15571,N_15380);
and U17723 (N_17723,N_15616,N_13172);
xnor U17724 (N_17724,N_12988,N_12535);
or U17725 (N_17725,N_13262,N_12786);
nor U17726 (N_17726,N_14363,N_13757);
and U17727 (N_17727,N_15034,N_13477);
xor U17728 (N_17728,N_13522,N_15039);
nor U17729 (N_17729,N_12965,N_14836);
nor U17730 (N_17730,N_13258,N_13063);
xnor U17731 (N_17731,N_13737,N_14157);
and U17732 (N_17732,N_12875,N_15431);
and U17733 (N_17733,N_12857,N_12576);
nand U17734 (N_17734,N_13517,N_14542);
xor U17735 (N_17735,N_13664,N_14080);
and U17736 (N_17736,N_15380,N_15560);
or U17737 (N_17737,N_12798,N_14850);
xor U17738 (N_17738,N_14081,N_15512);
xor U17739 (N_17739,N_13912,N_12933);
xor U17740 (N_17740,N_15194,N_13956);
nor U17741 (N_17741,N_15440,N_13901);
and U17742 (N_17742,N_13836,N_14952);
or U17743 (N_17743,N_15579,N_14767);
nand U17744 (N_17744,N_12749,N_12883);
xnor U17745 (N_17745,N_12583,N_12838);
or U17746 (N_17746,N_14118,N_13297);
or U17747 (N_17747,N_14566,N_13276);
and U17748 (N_17748,N_14365,N_13762);
or U17749 (N_17749,N_13614,N_15268);
xor U17750 (N_17750,N_13151,N_15609);
nor U17751 (N_17751,N_14202,N_15301);
nand U17752 (N_17752,N_14734,N_14580);
nand U17753 (N_17753,N_14388,N_14243);
or U17754 (N_17754,N_14879,N_14800);
nand U17755 (N_17755,N_12701,N_13318);
nor U17756 (N_17756,N_13924,N_13437);
xnor U17757 (N_17757,N_14706,N_12838);
nand U17758 (N_17758,N_14749,N_13170);
or U17759 (N_17759,N_13649,N_15432);
xor U17760 (N_17760,N_13773,N_14177);
or U17761 (N_17761,N_12828,N_15491);
and U17762 (N_17762,N_14953,N_13779);
or U17763 (N_17763,N_13068,N_14948);
nand U17764 (N_17764,N_12776,N_15569);
and U17765 (N_17765,N_12626,N_13554);
xor U17766 (N_17766,N_14397,N_14050);
and U17767 (N_17767,N_13380,N_14992);
and U17768 (N_17768,N_14191,N_15543);
nor U17769 (N_17769,N_13743,N_14109);
or U17770 (N_17770,N_15618,N_13436);
or U17771 (N_17771,N_15289,N_13134);
and U17772 (N_17772,N_15156,N_14688);
and U17773 (N_17773,N_13411,N_15539);
nor U17774 (N_17774,N_14052,N_14014);
xor U17775 (N_17775,N_15616,N_14214);
nor U17776 (N_17776,N_14703,N_12965);
nor U17777 (N_17777,N_14878,N_14760);
nand U17778 (N_17778,N_13909,N_15072);
and U17779 (N_17779,N_14292,N_15612);
or U17780 (N_17780,N_14001,N_13892);
or U17781 (N_17781,N_15057,N_13320);
xnor U17782 (N_17782,N_13439,N_15601);
nand U17783 (N_17783,N_15108,N_12624);
nor U17784 (N_17784,N_14877,N_13019);
or U17785 (N_17785,N_12732,N_13949);
or U17786 (N_17786,N_15372,N_12997);
xor U17787 (N_17787,N_12702,N_14890);
or U17788 (N_17788,N_15154,N_14346);
xor U17789 (N_17789,N_13635,N_14473);
nand U17790 (N_17790,N_14409,N_13751);
nand U17791 (N_17791,N_14911,N_13692);
xnor U17792 (N_17792,N_12671,N_13695);
nand U17793 (N_17793,N_13693,N_13480);
or U17794 (N_17794,N_13865,N_15015);
nor U17795 (N_17795,N_13120,N_14516);
nor U17796 (N_17796,N_13537,N_15362);
xor U17797 (N_17797,N_14940,N_14867);
or U17798 (N_17798,N_13524,N_14425);
and U17799 (N_17799,N_13244,N_14628);
nor U17800 (N_17800,N_15589,N_12818);
nor U17801 (N_17801,N_12800,N_15336);
nor U17802 (N_17802,N_12654,N_13257);
and U17803 (N_17803,N_13129,N_13512);
nand U17804 (N_17804,N_14224,N_14911);
nand U17805 (N_17805,N_14923,N_12754);
nand U17806 (N_17806,N_13605,N_12775);
and U17807 (N_17807,N_12828,N_15309);
or U17808 (N_17808,N_14273,N_15187);
and U17809 (N_17809,N_13568,N_14620);
or U17810 (N_17810,N_13655,N_14119);
nor U17811 (N_17811,N_14237,N_13734);
and U17812 (N_17812,N_14873,N_13048);
or U17813 (N_17813,N_14970,N_13269);
nor U17814 (N_17814,N_14821,N_15364);
or U17815 (N_17815,N_13596,N_13150);
and U17816 (N_17816,N_13833,N_13708);
and U17817 (N_17817,N_15413,N_14742);
or U17818 (N_17818,N_12753,N_15282);
xor U17819 (N_17819,N_13104,N_13599);
or U17820 (N_17820,N_13259,N_13509);
xor U17821 (N_17821,N_13193,N_13934);
nand U17822 (N_17822,N_14070,N_14800);
nor U17823 (N_17823,N_13276,N_14790);
or U17824 (N_17824,N_13042,N_14624);
nor U17825 (N_17825,N_14964,N_12952);
and U17826 (N_17826,N_13458,N_12895);
and U17827 (N_17827,N_15502,N_14335);
nor U17828 (N_17828,N_13444,N_14371);
nor U17829 (N_17829,N_15273,N_15131);
nand U17830 (N_17830,N_12706,N_12584);
and U17831 (N_17831,N_13531,N_15090);
xor U17832 (N_17832,N_12709,N_15190);
and U17833 (N_17833,N_14984,N_13233);
and U17834 (N_17834,N_13810,N_12662);
nand U17835 (N_17835,N_13634,N_12822);
nand U17836 (N_17836,N_13021,N_14809);
and U17837 (N_17837,N_14431,N_15503);
nand U17838 (N_17838,N_14473,N_13107);
and U17839 (N_17839,N_12816,N_15143);
xnor U17840 (N_17840,N_14097,N_13165);
and U17841 (N_17841,N_13459,N_13484);
nand U17842 (N_17842,N_13722,N_15373);
and U17843 (N_17843,N_14102,N_15295);
or U17844 (N_17844,N_13438,N_15271);
or U17845 (N_17845,N_12557,N_13734);
or U17846 (N_17846,N_12706,N_14582);
or U17847 (N_17847,N_13457,N_13525);
and U17848 (N_17848,N_13720,N_12564);
xnor U17849 (N_17849,N_12949,N_13396);
xor U17850 (N_17850,N_12522,N_12578);
and U17851 (N_17851,N_14086,N_14771);
or U17852 (N_17852,N_14328,N_15144);
nor U17853 (N_17853,N_13636,N_12714);
and U17854 (N_17854,N_12981,N_13812);
nor U17855 (N_17855,N_13760,N_13821);
nand U17856 (N_17856,N_13779,N_13055);
and U17857 (N_17857,N_14783,N_12623);
nand U17858 (N_17858,N_15207,N_15172);
xnor U17859 (N_17859,N_13808,N_13848);
nand U17860 (N_17860,N_12788,N_13578);
xor U17861 (N_17861,N_12664,N_15269);
xnor U17862 (N_17862,N_14225,N_14353);
nor U17863 (N_17863,N_13787,N_13642);
xnor U17864 (N_17864,N_12733,N_13173);
or U17865 (N_17865,N_12698,N_13281);
nand U17866 (N_17866,N_13912,N_14249);
nand U17867 (N_17867,N_15130,N_13772);
nor U17868 (N_17868,N_12965,N_14997);
nand U17869 (N_17869,N_14997,N_13996);
or U17870 (N_17870,N_13477,N_13465);
xor U17871 (N_17871,N_12582,N_13420);
and U17872 (N_17872,N_13078,N_14032);
xor U17873 (N_17873,N_12794,N_14311);
and U17874 (N_17874,N_13675,N_13234);
and U17875 (N_17875,N_15272,N_14484);
nand U17876 (N_17876,N_13165,N_15370);
xnor U17877 (N_17877,N_15391,N_13088);
or U17878 (N_17878,N_14745,N_15556);
or U17879 (N_17879,N_14565,N_12781);
nand U17880 (N_17880,N_14859,N_13808);
nor U17881 (N_17881,N_13298,N_15598);
and U17882 (N_17882,N_14430,N_15394);
nand U17883 (N_17883,N_14962,N_14213);
nand U17884 (N_17884,N_14741,N_12961);
nand U17885 (N_17885,N_14779,N_15352);
and U17886 (N_17886,N_14954,N_13204);
or U17887 (N_17887,N_15177,N_12667);
or U17888 (N_17888,N_13560,N_14175);
and U17889 (N_17889,N_13340,N_14601);
and U17890 (N_17890,N_14574,N_14657);
and U17891 (N_17891,N_12786,N_14092);
and U17892 (N_17892,N_13982,N_15520);
nor U17893 (N_17893,N_14937,N_15095);
xor U17894 (N_17894,N_13240,N_12879);
xnor U17895 (N_17895,N_12808,N_14574);
nor U17896 (N_17896,N_14719,N_13236);
nor U17897 (N_17897,N_14403,N_14714);
or U17898 (N_17898,N_13444,N_15082);
nor U17899 (N_17899,N_14953,N_12572);
nor U17900 (N_17900,N_15480,N_14455);
nand U17901 (N_17901,N_14048,N_14581);
or U17902 (N_17902,N_15605,N_12841);
and U17903 (N_17903,N_15118,N_15575);
nand U17904 (N_17904,N_14906,N_12709);
nor U17905 (N_17905,N_12687,N_14123);
nor U17906 (N_17906,N_13892,N_13021);
and U17907 (N_17907,N_14360,N_14326);
nand U17908 (N_17908,N_15067,N_13459);
xor U17909 (N_17909,N_12711,N_13736);
nor U17910 (N_17910,N_12563,N_15370);
nor U17911 (N_17911,N_13432,N_13689);
nand U17912 (N_17912,N_15412,N_14666);
nor U17913 (N_17913,N_13339,N_14687);
nor U17914 (N_17914,N_15513,N_12957);
nand U17915 (N_17915,N_14882,N_15600);
xor U17916 (N_17916,N_12837,N_13753);
nand U17917 (N_17917,N_12759,N_14860);
and U17918 (N_17918,N_13008,N_13560);
xnor U17919 (N_17919,N_14325,N_12860);
nand U17920 (N_17920,N_12567,N_15594);
and U17921 (N_17921,N_14015,N_14979);
and U17922 (N_17922,N_13050,N_12821);
xnor U17923 (N_17923,N_15190,N_12974);
or U17924 (N_17924,N_14274,N_15433);
nand U17925 (N_17925,N_12685,N_13269);
nand U17926 (N_17926,N_13551,N_14017);
nand U17927 (N_17927,N_13927,N_13567);
nand U17928 (N_17928,N_15061,N_13728);
nand U17929 (N_17929,N_15295,N_13089);
nand U17930 (N_17930,N_13279,N_14699);
or U17931 (N_17931,N_14976,N_12515);
nand U17932 (N_17932,N_12750,N_15209);
nor U17933 (N_17933,N_14707,N_14729);
and U17934 (N_17934,N_12826,N_13039);
or U17935 (N_17935,N_12849,N_13718);
or U17936 (N_17936,N_14566,N_15114);
nand U17937 (N_17937,N_12524,N_15362);
and U17938 (N_17938,N_14611,N_12818);
nor U17939 (N_17939,N_15437,N_12543);
xnor U17940 (N_17940,N_14071,N_13661);
and U17941 (N_17941,N_14952,N_14686);
or U17942 (N_17942,N_14682,N_15380);
nand U17943 (N_17943,N_12919,N_14278);
and U17944 (N_17944,N_12837,N_13934);
and U17945 (N_17945,N_13436,N_13036);
nor U17946 (N_17946,N_14117,N_14598);
xnor U17947 (N_17947,N_14911,N_14393);
or U17948 (N_17948,N_14325,N_14137);
nand U17949 (N_17949,N_13333,N_13400);
and U17950 (N_17950,N_15351,N_14940);
and U17951 (N_17951,N_14002,N_14862);
nand U17952 (N_17952,N_12914,N_15531);
nor U17953 (N_17953,N_15109,N_14427);
nand U17954 (N_17954,N_13112,N_15137);
nor U17955 (N_17955,N_14030,N_15540);
nor U17956 (N_17956,N_14185,N_15533);
or U17957 (N_17957,N_15124,N_12999);
nor U17958 (N_17958,N_14493,N_15382);
or U17959 (N_17959,N_13912,N_14984);
and U17960 (N_17960,N_12835,N_14122);
or U17961 (N_17961,N_13305,N_14230);
xor U17962 (N_17962,N_13198,N_13680);
nand U17963 (N_17963,N_14609,N_14763);
xor U17964 (N_17964,N_14123,N_13735);
xor U17965 (N_17965,N_15461,N_15043);
nand U17966 (N_17966,N_14405,N_13680);
or U17967 (N_17967,N_14771,N_15504);
nor U17968 (N_17968,N_14560,N_14013);
xor U17969 (N_17969,N_13364,N_12796);
nand U17970 (N_17970,N_12843,N_13884);
xnor U17971 (N_17971,N_15103,N_12595);
and U17972 (N_17972,N_15107,N_13454);
xnor U17973 (N_17973,N_14371,N_13906);
xor U17974 (N_17974,N_13993,N_14794);
nor U17975 (N_17975,N_14815,N_13070);
nor U17976 (N_17976,N_12879,N_14865);
xnor U17977 (N_17977,N_15467,N_15249);
xnor U17978 (N_17978,N_14785,N_13493);
or U17979 (N_17979,N_14918,N_13073);
and U17980 (N_17980,N_12799,N_12641);
or U17981 (N_17981,N_13314,N_12681);
or U17982 (N_17982,N_14413,N_14212);
xor U17983 (N_17983,N_12960,N_12575);
nor U17984 (N_17984,N_15285,N_14198);
and U17985 (N_17985,N_13099,N_14375);
xor U17986 (N_17986,N_13716,N_13972);
and U17987 (N_17987,N_14055,N_12511);
and U17988 (N_17988,N_12963,N_13817);
and U17989 (N_17989,N_12972,N_13351);
nor U17990 (N_17990,N_13221,N_15192);
and U17991 (N_17991,N_13768,N_14795);
and U17992 (N_17992,N_14679,N_13537);
xnor U17993 (N_17993,N_14052,N_13619);
and U17994 (N_17994,N_15513,N_14708);
xnor U17995 (N_17995,N_13047,N_12645);
or U17996 (N_17996,N_13257,N_14688);
or U17997 (N_17997,N_14263,N_13119);
xor U17998 (N_17998,N_14581,N_13532);
or U17999 (N_17999,N_12830,N_13841);
or U18000 (N_18000,N_12881,N_15263);
and U18001 (N_18001,N_12827,N_14791);
xor U18002 (N_18002,N_12860,N_15187);
or U18003 (N_18003,N_12858,N_12660);
nor U18004 (N_18004,N_14229,N_14585);
xor U18005 (N_18005,N_14769,N_13914);
nor U18006 (N_18006,N_14607,N_12730);
or U18007 (N_18007,N_13316,N_13023);
nand U18008 (N_18008,N_13263,N_12820);
nand U18009 (N_18009,N_15450,N_13570);
nand U18010 (N_18010,N_15241,N_13866);
and U18011 (N_18011,N_14363,N_14381);
or U18012 (N_18012,N_14674,N_15609);
xor U18013 (N_18013,N_13127,N_13096);
nor U18014 (N_18014,N_12953,N_14466);
and U18015 (N_18015,N_12627,N_14646);
nor U18016 (N_18016,N_14919,N_15531);
nand U18017 (N_18017,N_15366,N_13116);
xor U18018 (N_18018,N_13915,N_14675);
xnor U18019 (N_18019,N_15137,N_15139);
and U18020 (N_18020,N_13086,N_12926);
or U18021 (N_18021,N_15315,N_14659);
xor U18022 (N_18022,N_14140,N_14985);
and U18023 (N_18023,N_15218,N_13007);
xnor U18024 (N_18024,N_13998,N_15317);
nor U18025 (N_18025,N_14106,N_12762);
nand U18026 (N_18026,N_14742,N_13689);
nand U18027 (N_18027,N_12943,N_13401);
nand U18028 (N_18028,N_15479,N_15032);
nand U18029 (N_18029,N_15130,N_12912);
nor U18030 (N_18030,N_14636,N_13989);
nor U18031 (N_18031,N_13761,N_13720);
or U18032 (N_18032,N_15096,N_15506);
nand U18033 (N_18033,N_13820,N_14429);
and U18034 (N_18034,N_13903,N_13269);
xnor U18035 (N_18035,N_12623,N_15431);
nor U18036 (N_18036,N_12873,N_13695);
nor U18037 (N_18037,N_12845,N_15586);
nor U18038 (N_18038,N_13191,N_14255);
nor U18039 (N_18039,N_13265,N_14332);
nor U18040 (N_18040,N_14868,N_13278);
or U18041 (N_18041,N_14206,N_12935);
or U18042 (N_18042,N_12931,N_14339);
nor U18043 (N_18043,N_13442,N_13435);
nor U18044 (N_18044,N_13185,N_15375);
xnor U18045 (N_18045,N_15361,N_12713);
or U18046 (N_18046,N_14275,N_14099);
xor U18047 (N_18047,N_14984,N_12549);
or U18048 (N_18048,N_14015,N_14586);
xnor U18049 (N_18049,N_13163,N_14980);
nor U18050 (N_18050,N_13686,N_14116);
nor U18051 (N_18051,N_14592,N_13741);
and U18052 (N_18052,N_12791,N_12667);
xor U18053 (N_18053,N_14409,N_12680);
xor U18054 (N_18054,N_14059,N_13134);
and U18055 (N_18055,N_14462,N_15035);
xor U18056 (N_18056,N_14734,N_14907);
xnor U18057 (N_18057,N_15055,N_14984);
xor U18058 (N_18058,N_14404,N_14041);
and U18059 (N_18059,N_15369,N_14718);
or U18060 (N_18060,N_13327,N_14868);
and U18061 (N_18061,N_13135,N_14412);
and U18062 (N_18062,N_12967,N_13722);
and U18063 (N_18063,N_12626,N_14931);
and U18064 (N_18064,N_14038,N_13600);
and U18065 (N_18065,N_12917,N_13379);
and U18066 (N_18066,N_15231,N_13347);
xor U18067 (N_18067,N_13484,N_12802);
xnor U18068 (N_18068,N_13438,N_15072);
nand U18069 (N_18069,N_13690,N_13747);
and U18070 (N_18070,N_14706,N_14797);
or U18071 (N_18071,N_13673,N_13998);
nand U18072 (N_18072,N_14278,N_14771);
nor U18073 (N_18073,N_15107,N_12592);
xnor U18074 (N_18074,N_15260,N_15090);
and U18075 (N_18075,N_13779,N_13037);
nor U18076 (N_18076,N_14849,N_15025);
or U18077 (N_18077,N_14966,N_13513);
or U18078 (N_18078,N_13155,N_13338);
nor U18079 (N_18079,N_12857,N_15154);
and U18080 (N_18080,N_12693,N_12829);
nor U18081 (N_18081,N_15623,N_14125);
and U18082 (N_18082,N_14635,N_12780);
xnor U18083 (N_18083,N_14099,N_12526);
xnor U18084 (N_18084,N_12895,N_13815);
and U18085 (N_18085,N_14514,N_12867);
nor U18086 (N_18086,N_15576,N_13584);
and U18087 (N_18087,N_12837,N_14599);
nor U18088 (N_18088,N_14761,N_15552);
nand U18089 (N_18089,N_14826,N_14434);
and U18090 (N_18090,N_14449,N_12981);
and U18091 (N_18091,N_14193,N_15493);
nor U18092 (N_18092,N_15406,N_15124);
or U18093 (N_18093,N_14947,N_15355);
xnor U18094 (N_18094,N_14258,N_14189);
or U18095 (N_18095,N_12914,N_14716);
nor U18096 (N_18096,N_13165,N_12730);
or U18097 (N_18097,N_12520,N_13269);
nand U18098 (N_18098,N_14106,N_12562);
xnor U18099 (N_18099,N_13686,N_14937);
and U18100 (N_18100,N_13616,N_13010);
or U18101 (N_18101,N_15148,N_13617);
nand U18102 (N_18102,N_14466,N_13266);
xnor U18103 (N_18103,N_15313,N_13416);
nand U18104 (N_18104,N_13877,N_13097);
and U18105 (N_18105,N_14514,N_14816);
or U18106 (N_18106,N_13856,N_14540);
or U18107 (N_18107,N_14548,N_15102);
nand U18108 (N_18108,N_13444,N_12518);
nand U18109 (N_18109,N_13172,N_14790);
nand U18110 (N_18110,N_14802,N_14758);
nor U18111 (N_18111,N_13778,N_13210);
nand U18112 (N_18112,N_15195,N_14711);
xor U18113 (N_18113,N_13855,N_14254);
nand U18114 (N_18114,N_14363,N_15484);
nand U18115 (N_18115,N_13491,N_14598);
and U18116 (N_18116,N_14303,N_13450);
nand U18117 (N_18117,N_12633,N_13982);
xor U18118 (N_18118,N_15322,N_14866);
nor U18119 (N_18119,N_14529,N_12589);
and U18120 (N_18120,N_12765,N_14853);
xor U18121 (N_18121,N_12576,N_12959);
or U18122 (N_18122,N_12681,N_12978);
and U18123 (N_18123,N_14081,N_14756);
xor U18124 (N_18124,N_12716,N_13564);
and U18125 (N_18125,N_12504,N_13944);
nand U18126 (N_18126,N_15300,N_12829);
and U18127 (N_18127,N_15406,N_14690);
nand U18128 (N_18128,N_14301,N_14601);
nand U18129 (N_18129,N_13163,N_13617);
and U18130 (N_18130,N_15104,N_15204);
nor U18131 (N_18131,N_13231,N_13918);
and U18132 (N_18132,N_12825,N_14444);
or U18133 (N_18133,N_13246,N_15310);
nand U18134 (N_18134,N_13160,N_14024);
nand U18135 (N_18135,N_13672,N_14753);
xor U18136 (N_18136,N_15119,N_13799);
and U18137 (N_18137,N_14518,N_13492);
xnor U18138 (N_18138,N_13367,N_14964);
or U18139 (N_18139,N_13043,N_13244);
and U18140 (N_18140,N_14360,N_15385);
or U18141 (N_18141,N_14228,N_15422);
or U18142 (N_18142,N_13311,N_13244);
nor U18143 (N_18143,N_15282,N_15130);
xor U18144 (N_18144,N_14704,N_13597);
nand U18145 (N_18145,N_12961,N_12786);
xor U18146 (N_18146,N_12658,N_12524);
nor U18147 (N_18147,N_14828,N_13707);
and U18148 (N_18148,N_13724,N_14761);
xor U18149 (N_18149,N_12802,N_14692);
xnor U18150 (N_18150,N_15119,N_12976);
or U18151 (N_18151,N_12939,N_14051);
and U18152 (N_18152,N_14520,N_14291);
and U18153 (N_18153,N_13710,N_12731);
and U18154 (N_18154,N_15073,N_15336);
nor U18155 (N_18155,N_14410,N_13523);
xnor U18156 (N_18156,N_14276,N_14231);
and U18157 (N_18157,N_13951,N_13350);
nand U18158 (N_18158,N_13654,N_13387);
xor U18159 (N_18159,N_13312,N_13976);
nor U18160 (N_18160,N_13801,N_15306);
or U18161 (N_18161,N_14256,N_14883);
and U18162 (N_18162,N_15476,N_15276);
nor U18163 (N_18163,N_12756,N_13787);
or U18164 (N_18164,N_13236,N_13556);
xor U18165 (N_18165,N_14010,N_13453);
xor U18166 (N_18166,N_12883,N_15589);
xnor U18167 (N_18167,N_15164,N_13539);
xnor U18168 (N_18168,N_13424,N_13726);
nand U18169 (N_18169,N_13531,N_15386);
or U18170 (N_18170,N_13812,N_14736);
xnor U18171 (N_18171,N_14980,N_14532);
or U18172 (N_18172,N_13258,N_15530);
xnor U18173 (N_18173,N_13405,N_14935);
nand U18174 (N_18174,N_12512,N_13627);
xnor U18175 (N_18175,N_15310,N_14877);
or U18176 (N_18176,N_14584,N_12576);
xnor U18177 (N_18177,N_13875,N_15498);
nor U18178 (N_18178,N_15047,N_14619);
or U18179 (N_18179,N_14930,N_14269);
xor U18180 (N_18180,N_15180,N_15154);
nor U18181 (N_18181,N_14410,N_13342);
xnor U18182 (N_18182,N_13508,N_13088);
or U18183 (N_18183,N_15546,N_12544);
nand U18184 (N_18184,N_12863,N_12735);
nand U18185 (N_18185,N_13345,N_12933);
xnor U18186 (N_18186,N_13898,N_14267);
nor U18187 (N_18187,N_14955,N_13830);
and U18188 (N_18188,N_13381,N_12509);
nand U18189 (N_18189,N_14618,N_15072);
xor U18190 (N_18190,N_13195,N_14101);
and U18191 (N_18191,N_12775,N_14375);
and U18192 (N_18192,N_14574,N_12926);
and U18193 (N_18193,N_13930,N_14102);
nand U18194 (N_18194,N_14886,N_13867);
or U18195 (N_18195,N_14032,N_15053);
and U18196 (N_18196,N_13764,N_13897);
and U18197 (N_18197,N_13918,N_14081);
xnor U18198 (N_18198,N_13633,N_14559);
and U18199 (N_18199,N_14894,N_14936);
and U18200 (N_18200,N_12661,N_15250);
nor U18201 (N_18201,N_15026,N_13765);
and U18202 (N_18202,N_14837,N_12671);
and U18203 (N_18203,N_13669,N_14261);
xnor U18204 (N_18204,N_15463,N_14574);
and U18205 (N_18205,N_12879,N_13064);
and U18206 (N_18206,N_15415,N_14439);
and U18207 (N_18207,N_14394,N_13528);
nor U18208 (N_18208,N_14980,N_13362);
or U18209 (N_18209,N_14953,N_15317);
xor U18210 (N_18210,N_15139,N_15341);
xor U18211 (N_18211,N_14834,N_14746);
or U18212 (N_18212,N_13321,N_15460);
nand U18213 (N_18213,N_14925,N_13676);
nand U18214 (N_18214,N_14143,N_14049);
nand U18215 (N_18215,N_15142,N_15541);
and U18216 (N_18216,N_12940,N_15413);
and U18217 (N_18217,N_14529,N_13367);
nand U18218 (N_18218,N_14488,N_15215);
xnor U18219 (N_18219,N_12687,N_14589);
or U18220 (N_18220,N_14564,N_12545);
or U18221 (N_18221,N_13279,N_12911);
nand U18222 (N_18222,N_14384,N_14357);
xnor U18223 (N_18223,N_14639,N_15388);
or U18224 (N_18224,N_13663,N_13829);
nor U18225 (N_18225,N_13157,N_13624);
and U18226 (N_18226,N_14079,N_12748);
or U18227 (N_18227,N_13806,N_13363);
and U18228 (N_18228,N_15406,N_13393);
nand U18229 (N_18229,N_13697,N_15224);
nand U18230 (N_18230,N_14842,N_15089);
and U18231 (N_18231,N_13419,N_13590);
nand U18232 (N_18232,N_14370,N_13447);
nor U18233 (N_18233,N_12657,N_14621);
nor U18234 (N_18234,N_12570,N_15358);
or U18235 (N_18235,N_13476,N_14049);
xnor U18236 (N_18236,N_15088,N_13859);
nor U18237 (N_18237,N_14748,N_12650);
nand U18238 (N_18238,N_14447,N_15152);
nand U18239 (N_18239,N_15408,N_13150);
nor U18240 (N_18240,N_14283,N_13575);
xnor U18241 (N_18241,N_14576,N_13977);
and U18242 (N_18242,N_12626,N_13155);
and U18243 (N_18243,N_14197,N_15281);
or U18244 (N_18244,N_14353,N_15540);
or U18245 (N_18245,N_15402,N_12712);
xor U18246 (N_18246,N_13905,N_13993);
nand U18247 (N_18247,N_14241,N_12518);
nand U18248 (N_18248,N_13421,N_14366);
or U18249 (N_18249,N_14606,N_15091);
nor U18250 (N_18250,N_14272,N_12887);
xnor U18251 (N_18251,N_13818,N_14816);
and U18252 (N_18252,N_14128,N_13592);
and U18253 (N_18253,N_13610,N_14773);
or U18254 (N_18254,N_13594,N_13325);
xor U18255 (N_18255,N_15509,N_14537);
nand U18256 (N_18256,N_14446,N_13310);
xnor U18257 (N_18257,N_13608,N_14719);
and U18258 (N_18258,N_13442,N_13839);
xor U18259 (N_18259,N_13385,N_15037);
or U18260 (N_18260,N_12893,N_14791);
nand U18261 (N_18261,N_14342,N_15021);
and U18262 (N_18262,N_15044,N_13916);
xor U18263 (N_18263,N_13158,N_13340);
nor U18264 (N_18264,N_15031,N_15129);
nor U18265 (N_18265,N_13399,N_13558);
xnor U18266 (N_18266,N_15451,N_14966);
xor U18267 (N_18267,N_14473,N_12825);
and U18268 (N_18268,N_13080,N_13367);
and U18269 (N_18269,N_12791,N_14114);
nor U18270 (N_18270,N_13366,N_14770);
nand U18271 (N_18271,N_13873,N_13312);
and U18272 (N_18272,N_15531,N_15368);
nand U18273 (N_18273,N_13547,N_14303);
or U18274 (N_18274,N_15216,N_12947);
nand U18275 (N_18275,N_13327,N_13718);
nor U18276 (N_18276,N_15486,N_13453);
nor U18277 (N_18277,N_12727,N_13698);
or U18278 (N_18278,N_13217,N_12699);
or U18279 (N_18279,N_14331,N_12901);
and U18280 (N_18280,N_14467,N_13538);
nor U18281 (N_18281,N_14546,N_12992);
xnor U18282 (N_18282,N_15598,N_12880);
nand U18283 (N_18283,N_15360,N_13700);
or U18284 (N_18284,N_14259,N_14846);
and U18285 (N_18285,N_13370,N_15011);
nand U18286 (N_18286,N_14046,N_13829);
nand U18287 (N_18287,N_13921,N_14782);
and U18288 (N_18288,N_14717,N_15415);
nand U18289 (N_18289,N_14443,N_14384);
or U18290 (N_18290,N_15160,N_13710);
or U18291 (N_18291,N_12894,N_12983);
nand U18292 (N_18292,N_15013,N_15438);
or U18293 (N_18293,N_15544,N_13733);
xor U18294 (N_18294,N_14073,N_15317);
and U18295 (N_18295,N_13087,N_15251);
or U18296 (N_18296,N_14962,N_14990);
nor U18297 (N_18297,N_13961,N_13375);
or U18298 (N_18298,N_12504,N_12699);
and U18299 (N_18299,N_14034,N_14855);
xnor U18300 (N_18300,N_14443,N_14473);
nand U18301 (N_18301,N_13498,N_13445);
nor U18302 (N_18302,N_13827,N_14764);
and U18303 (N_18303,N_13469,N_12697);
xnor U18304 (N_18304,N_14473,N_14297);
and U18305 (N_18305,N_13564,N_14040);
or U18306 (N_18306,N_13904,N_13850);
nand U18307 (N_18307,N_14385,N_14580);
xor U18308 (N_18308,N_14601,N_13390);
and U18309 (N_18309,N_12934,N_15155);
xnor U18310 (N_18310,N_13241,N_12504);
xor U18311 (N_18311,N_13393,N_13398);
nor U18312 (N_18312,N_15058,N_13067);
or U18313 (N_18313,N_13047,N_15005);
and U18314 (N_18314,N_14165,N_14151);
nand U18315 (N_18315,N_14594,N_13060);
and U18316 (N_18316,N_15010,N_15397);
nor U18317 (N_18317,N_15365,N_13060);
and U18318 (N_18318,N_15001,N_15376);
xnor U18319 (N_18319,N_14286,N_13923);
nor U18320 (N_18320,N_13666,N_12831);
xor U18321 (N_18321,N_13375,N_14301);
nor U18322 (N_18322,N_13489,N_13371);
and U18323 (N_18323,N_14320,N_13500);
and U18324 (N_18324,N_13354,N_14968);
or U18325 (N_18325,N_14293,N_15190);
nand U18326 (N_18326,N_13833,N_12586);
or U18327 (N_18327,N_13710,N_15494);
or U18328 (N_18328,N_12781,N_13559);
nor U18329 (N_18329,N_14777,N_13010);
nand U18330 (N_18330,N_13672,N_13070);
xor U18331 (N_18331,N_13983,N_12739);
and U18332 (N_18332,N_14657,N_15250);
xnor U18333 (N_18333,N_14035,N_13018);
and U18334 (N_18334,N_14929,N_13353);
xor U18335 (N_18335,N_14257,N_15408);
xnor U18336 (N_18336,N_14713,N_13431);
and U18337 (N_18337,N_14781,N_14238);
and U18338 (N_18338,N_12969,N_13362);
or U18339 (N_18339,N_13159,N_14334);
or U18340 (N_18340,N_15095,N_14598);
or U18341 (N_18341,N_12724,N_12946);
nor U18342 (N_18342,N_12563,N_15033);
or U18343 (N_18343,N_15405,N_14811);
or U18344 (N_18344,N_14442,N_14987);
or U18345 (N_18345,N_13537,N_15584);
and U18346 (N_18346,N_14829,N_15150);
nand U18347 (N_18347,N_13696,N_13637);
nand U18348 (N_18348,N_13181,N_13636);
or U18349 (N_18349,N_14174,N_14474);
xnor U18350 (N_18350,N_14938,N_14620);
nand U18351 (N_18351,N_15490,N_15616);
nand U18352 (N_18352,N_14914,N_15564);
or U18353 (N_18353,N_15231,N_13927);
xnor U18354 (N_18354,N_12607,N_12932);
and U18355 (N_18355,N_13943,N_14263);
and U18356 (N_18356,N_12570,N_12830);
or U18357 (N_18357,N_14750,N_15305);
xnor U18358 (N_18358,N_13056,N_15250);
nand U18359 (N_18359,N_14454,N_14775);
nand U18360 (N_18360,N_15512,N_14767);
nor U18361 (N_18361,N_12712,N_15581);
and U18362 (N_18362,N_12954,N_14238);
and U18363 (N_18363,N_13912,N_13970);
xnor U18364 (N_18364,N_14687,N_14641);
and U18365 (N_18365,N_13769,N_13148);
or U18366 (N_18366,N_12800,N_14085);
and U18367 (N_18367,N_14459,N_14771);
or U18368 (N_18368,N_15006,N_13423);
and U18369 (N_18369,N_12626,N_15358);
or U18370 (N_18370,N_12523,N_14633);
xnor U18371 (N_18371,N_15564,N_13044);
nor U18372 (N_18372,N_15563,N_14155);
nor U18373 (N_18373,N_14945,N_12997);
xnor U18374 (N_18374,N_12971,N_14956);
nor U18375 (N_18375,N_13332,N_13409);
and U18376 (N_18376,N_13842,N_13665);
or U18377 (N_18377,N_14189,N_13066);
xnor U18378 (N_18378,N_15400,N_14375);
and U18379 (N_18379,N_13874,N_13510);
or U18380 (N_18380,N_12557,N_14190);
or U18381 (N_18381,N_12512,N_13413);
and U18382 (N_18382,N_15409,N_15025);
nor U18383 (N_18383,N_14451,N_14288);
and U18384 (N_18384,N_15426,N_13964);
nand U18385 (N_18385,N_14557,N_15474);
nor U18386 (N_18386,N_13500,N_13572);
xnor U18387 (N_18387,N_15172,N_13174);
or U18388 (N_18388,N_12941,N_14326);
xor U18389 (N_18389,N_13039,N_13746);
and U18390 (N_18390,N_14213,N_15293);
nor U18391 (N_18391,N_15318,N_14838);
xnor U18392 (N_18392,N_14007,N_12928);
nor U18393 (N_18393,N_12745,N_14154);
and U18394 (N_18394,N_13165,N_12558);
or U18395 (N_18395,N_15532,N_13983);
nand U18396 (N_18396,N_13677,N_13099);
nor U18397 (N_18397,N_14064,N_15198);
xnor U18398 (N_18398,N_13198,N_12963);
and U18399 (N_18399,N_14895,N_15365);
and U18400 (N_18400,N_15272,N_13102);
or U18401 (N_18401,N_13733,N_13099);
and U18402 (N_18402,N_12500,N_13214);
nand U18403 (N_18403,N_14578,N_14412);
nand U18404 (N_18404,N_15412,N_15235);
xnor U18405 (N_18405,N_14681,N_13612);
or U18406 (N_18406,N_12598,N_15586);
and U18407 (N_18407,N_15134,N_13875);
or U18408 (N_18408,N_14566,N_15435);
nand U18409 (N_18409,N_15504,N_15209);
xor U18410 (N_18410,N_14544,N_13103);
or U18411 (N_18411,N_12739,N_12628);
and U18412 (N_18412,N_14413,N_13484);
or U18413 (N_18413,N_13990,N_13274);
xor U18414 (N_18414,N_15601,N_13217);
xnor U18415 (N_18415,N_13994,N_15050);
nor U18416 (N_18416,N_14430,N_14617);
and U18417 (N_18417,N_15487,N_13105);
xor U18418 (N_18418,N_15216,N_15582);
or U18419 (N_18419,N_12883,N_15281);
xnor U18420 (N_18420,N_15554,N_14936);
nor U18421 (N_18421,N_14825,N_14631);
nand U18422 (N_18422,N_12689,N_13080);
xnor U18423 (N_18423,N_15036,N_13932);
nor U18424 (N_18424,N_13796,N_13620);
nor U18425 (N_18425,N_13097,N_14190);
xnor U18426 (N_18426,N_13477,N_14835);
or U18427 (N_18427,N_14527,N_13701);
nor U18428 (N_18428,N_12821,N_13197);
and U18429 (N_18429,N_12650,N_15246);
nand U18430 (N_18430,N_13618,N_14786);
xnor U18431 (N_18431,N_14946,N_12544);
nor U18432 (N_18432,N_15428,N_13925);
nand U18433 (N_18433,N_14391,N_14019);
or U18434 (N_18434,N_14763,N_12541);
nand U18435 (N_18435,N_14524,N_14204);
nor U18436 (N_18436,N_13963,N_13676);
nor U18437 (N_18437,N_13582,N_12627);
and U18438 (N_18438,N_14491,N_15078);
xnor U18439 (N_18439,N_12968,N_13346);
nand U18440 (N_18440,N_12915,N_13777);
nor U18441 (N_18441,N_12717,N_15436);
nor U18442 (N_18442,N_14530,N_12849);
nand U18443 (N_18443,N_14112,N_13089);
nor U18444 (N_18444,N_13642,N_14700);
or U18445 (N_18445,N_13643,N_13851);
and U18446 (N_18446,N_15333,N_14055);
nor U18447 (N_18447,N_13384,N_15495);
nand U18448 (N_18448,N_14806,N_13162);
nor U18449 (N_18449,N_12884,N_14779);
and U18450 (N_18450,N_12525,N_14142);
xnor U18451 (N_18451,N_12678,N_14976);
nand U18452 (N_18452,N_15364,N_12603);
or U18453 (N_18453,N_13164,N_14149);
nand U18454 (N_18454,N_15119,N_13097);
nor U18455 (N_18455,N_13958,N_14383);
and U18456 (N_18456,N_14951,N_14851);
xnor U18457 (N_18457,N_13015,N_15047);
or U18458 (N_18458,N_13543,N_13362);
and U18459 (N_18459,N_15135,N_15417);
or U18460 (N_18460,N_13829,N_14056);
xor U18461 (N_18461,N_14939,N_12686);
and U18462 (N_18462,N_13810,N_13239);
or U18463 (N_18463,N_12719,N_13411);
and U18464 (N_18464,N_12803,N_12558);
nand U18465 (N_18465,N_14932,N_15429);
or U18466 (N_18466,N_13799,N_13543);
nor U18467 (N_18467,N_14510,N_12794);
or U18468 (N_18468,N_13058,N_13640);
and U18469 (N_18469,N_14926,N_14653);
nand U18470 (N_18470,N_12636,N_15033);
nor U18471 (N_18471,N_14451,N_14232);
nand U18472 (N_18472,N_13530,N_13723);
nand U18473 (N_18473,N_13304,N_14621);
or U18474 (N_18474,N_12648,N_14288);
or U18475 (N_18475,N_13395,N_15006);
nor U18476 (N_18476,N_14327,N_14813);
nand U18477 (N_18477,N_14391,N_15592);
nand U18478 (N_18478,N_14616,N_13389);
and U18479 (N_18479,N_15515,N_15363);
nand U18480 (N_18480,N_15014,N_13104);
nor U18481 (N_18481,N_13579,N_13212);
nand U18482 (N_18482,N_13834,N_13002);
nor U18483 (N_18483,N_15352,N_15322);
xnor U18484 (N_18484,N_15073,N_15329);
and U18485 (N_18485,N_15377,N_12651);
nand U18486 (N_18486,N_14558,N_12708);
xor U18487 (N_18487,N_13147,N_13349);
xnor U18488 (N_18488,N_12888,N_13275);
nor U18489 (N_18489,N_15204,N_14617);
or U18490 (N_18490,N_12604,N_12738);
nand U18491 (N_18491,N_13512,N_14411);
xor U18492 (N_18492,N_15227,N_12754);
xor U18493 (N_18493,N_13086,N_13776);
and U18494 (N_18494,N_12513,N_13431);
xor U18495 (N_18495,N_15254,N_12758);
nand U18496 (N_18496,N_15553,N_12615);
nand U18497 (N_18497,N_13382,N_12975);
nor U18498 (N_18498,N_14830,N_13933);
or U18499 (N_18499,N_13342,N_14614);
xor U18500 (N_18500,N_14733,N_13360);
xnor U18501 (N_18501,N_13629,N_13744);
xnor U18502 (N_18502,N_15107,N_15119);
or U18503 (N_18503,N_13701,N_13196);
xnor U18504 (N_18504,N_12569,N_14242);
or U18505 (N_18505,N_14416,N_13447);
nand U18506 (N_18506,N_15076,N_13808);
and U18507 (N_18507,N_14366,N_13324);
nor U18508 (N_18508,N_12645,N_15053);
xnor U18509 (N_18509,N_12633,N_14646);
or U18510 (N_18510,N_15017,N_13572);
or U18511 (N_18511,N_15282,N_14354);
or U18512 (N_18512,N_13399,N_14827);
nand U18513 (N_18513,N_13627,N_13172);
nor U18514 (N_18514,N_14942,N_14957);
xnor U18515 (N_18515,N_15439,N_12939);
or U18516 (N_18516,N_14562,N_14199);
or U18517 (N_18517,N_14950,N_14987);
and U18518 (N_18518,N_12636,N_14286);
nand U18519 (N_18519,N_14770,N_15347);
xnor U18520 (N_18520,N_14908,N_15147);
or U18521 (N_18521,N_12673,N_14318);
xor U18522 (N_18522,N_15385,N_13433);
xnor U18523 (N_18523,N_15527,N_14532);
and U18524 (N_18524,N_12605,N_13068);
nand U18525 (N_18525,N_13424,N_14978);
xor U18526 (N_18526,N_14951,N_13406);
nor U18527 (N_18527,N_15039,N_14631);
nor U18528 (N_18528,N_12993,N_12961);
and U18529 (N_18529,N_13826,N_13113);
and U18530 (N_18530,N_15524,N_13401);
nor U18531 (N_18531,N_12709,N_15009);
nor U18532 (N_18532,N_14579,N_13989);
nand U18533 (N_18533,N_14551,N_14968);
xor U18534 (N_18534,N_13294,N_15497);
nor U18535 (N_18535,N_13939,N_15253);
or U18536 (N_18536,N_12893,N_14067);
nor U18537 (N_18537,N_15207,N_14084);
xor U18538 (N_18538,N_13767,N_13466);
and U18539 (N_18539,N_15119,N_14527);
or U18540 (N_18540,N_14398,N_13598);
or U18541 (N_18541,N_13970,N_13768);
and U18542 (N_18542,N_14618,N_13253);
nand U18543 (N_18543,N_14218,N_14363);
xor U18544 (N_18544,N_12723,N_15373);
xor U18545 (N_18545,N_12796,N_13428);
xnor U18546 (N_18546,N_14036,N_15530);
nand U18547 (N_18547,N_14386,N_15541);
and U18548 (N_18548,N_13470,N_14384);
xor U18549 (N_18549,N_15225,N_15038);
and U18550 (N_18550,N_14894,N_13286);
nand U18551 (N_18551,N_15048,N_14216);
or U18552 (N_18552,N_15148,N_13155);
nand U18553 (N_18553,N_12626,N_14111);
xnor U18554 (N_18554,N_14311,N_14430);
and U18555 (N_18555,N_13866,N_14439);
or U18556 (N_18556,N_12530,N_13419);
nor U18557 (N_18557,N_12788,N_15441);
and U18558 (N_18558,N_15120,N_13892);
xnor U18559 (N_18559,N_13030,N_14063);
xor U18560 (N_18560,N_13253,N_12762);
or U18561 (N_18561,N_13972,N_13940);
nand U18562 (N_18562,N_13843,N_12814);
nor U18563 (N_18563,N_13786,N_13618);
nor U18564 (N_18564,N_14228,N_14627);
nor U18565 (N_18565,N_14290,N_12671);
and U18566 (N_18566,N_13559,N_12641);
and U18567 (N_18567,N_14111,N_13161);
or U18568 (N_18568,N_14997,N_14464);
or U18569 (N_18569,N_14074,N_13192);
and U18570 (N_18570,N_13874,N_12582);
xnor U18571 (N_18571,N_14950,N_12807);
or U18572 (N_18572,N_14791,N_13338);
or U18573 (N_18573,N_13142,N_13631);
xnor U18574 (N_18574,N_12928,N_13367);
nor U18575 (N_18575,N_13811,N_13218);
nor U18576 (N_18576,N_13820,N_13167);
xnor U18577 (N_18577,N_13876,N_12755);
or U18578 (N_18578,N_15412,N_13169);
nor U18579 (N_18579,N_13287,N_13213);
and U18580 (N_18580,N_14527,N_13942);
or U18581 (N_18581,N_15451,N_13764);
xor U18582 (N_18582,N_14563,N_15489);
nand U18583 (N_18583,N_13252,N_15072);
xor U18584 (N_18584,N_15123,N_14322);
xor U18585 (N_18585,N_13929,N_13668);
and U18586 (N_18586,N_13328,N_13029);
and U18587 (N_18587,N_12510,N_14961);
nand U18588 (N_18588,N_13724,N_14926);
xnor U18589 (N_18589,N_13498,N_15557);
xor U18590 (N_18590,N_13019,N_13504);
nor U18591 (N_18591,N_15450,N_14836);
nand U18592 (N_18592,N_13552,N_15547);
nand U18593 (N_18593,N_12584,N_12699);
nor U18594 (N_18594,N_14480,N_15385);
or U18595 (N_18595,N_12771,N_14919);
nand U18596 (N_18596,N_15612,N_12730);
nor U18597 (N_18597,N_13323,N_14886);
nand U18598 (N_18598,N_13095,N_14210);
and U18599 (N_18599,N_13265,N_13814);
nor U18600 (N_18600,N_13916,N_13099);
or U18601 (N_18601,N_13735,N_12618);
xnor U18602 (N_18602,N_14637,N_14525);
or U18603 (N_18603,N_12654,N_13127);
or U18604 (N_18604,N_12786,N_14225);
or U18605 (N_18605,N_12623,N_15073);
xnor U18606 (N_18606,N_14843,N_13800);
and U18607 (N_18607,N_14725,N_12544);
or U18608 (N_18608,N_13940,N_14780);
nand U18609 (N_18609,N_15557,N_15402);
and U18610 (N_18610,N_13323,N_12746);
nand U18611 (N_18611,N_15052,N_14722);
nand U18612 (N_18612,N_15622,N_14220);
or U18613 (N_18613,N_14064,N_14580);
nand U18614 (N_18614,N_13659,N_15358);
nor U18615 (N_18615,N_12831,N_13815);
nor U18616 (N_18616,N_14986,N_15201);
nor U18617 (N_18617,N_15360,N_15206);
xor U18618 (N_18618,N_14017,N_13459);
nor U18619 (N_18619,N_12926,N_14638);
nor U18620 (N_18620,N_13174,N_14369);
nor U18621 (N_18621,N_15459,N_13527);
or U18622 (N_18622,N_14126,N_15393);
and U18623 (N_18623,N_13268,N_12581);
nand U18624 (N_18624,N_13982,N_15068);
or U18625 (N_18625,N_13276,N_15449);
or U18626 (N_18626,N_13839,N_13544);
nand U18627 (N_18627,N_12667,N_14073);
and U18628 (N_18628,N_15257,N_14630);
and U18629 (N_18629,N_13455,N_12751);
nand U18630 (N_18630,N_13410,N_14881);
xnor U18631 (N_18631,N_13453,N_14330);
xnor U18632 (N_18632,N_13928,N_14484);
and U18633 (N_18633,N_14215,N_14780);
xor U18634 (N_18634,N_13372,N_15201);
xor U18635 (N_18635,N_12894,N_15370);
xor U18636 (N_18636,N_14870,N_13989);
nor U18637 (N_18637,N_14478,N_14358);
nand U18638 (N_18638,N_14862,N_13829);
and U18639 (N_18639,N_15499,N_15257);
nand U18640 (N_18640,N_12708,N_14744);
nand U18641 (N_18641,N_12566,N_13902);
nor U18642 (N_18642,N_13523,N_12571);
or U18643 (N_18643,N_15409,N_14126);
and U18644 (N_18644,N_14630,N_12549);
nand U18645 (N_18645,N_13449,N_15530);
and U18646 (N_18646,N_15245,N_13642);
and U18647 (N_18647,N_15301,N_13340);
nand U18648 (N_18648,N_14781,N_12684);
nor U18649 (N_18649,N_15349,N_13590);
nand U18650 (N_18650,N_13498,N_14531);
and U18651 (N_18651,N_12999,N_15532);
and U18652 (N_18652,N_14581,N_14264);
and U18653 (N_18653,N_12752,N_12809);
nor U18654 (N_18654,N_14665,N_13430);
xnor U18655 (N_18655,N_13942,N_13439);
and U18656 (N_18656,N_15600,N_13309);
xor U18657 (N_18657,N_13294,N_15412);
nand U18658 (N_18658,N_15543,N_14359);
xor U18659 (N_18659,N_12712,N_12636);
and U18660 (N_18660,N_15614,N_13181);
or U18661 (N_18661,N_15542,N_13062);
and U18662 (N_18662,N_13395,N_12694);
nand U18663 (N_18663,N_14086,N_14512);
xnor U18664 (N_18664,N_13684,N_15201);
nand U18665 (N_18665,N_13154,N_15099);
or U18666 (N_18666,N_15236,N_13654);
and U18667 (N_18667,N_12720,N_15266);
and U18668 (N_18668,N_13733,N_13138);
nor U18669 (N_18669,N_14517,N_12851);
xnor U18670 (N_18670,N_12539,N_12897);
xor U18671 (N_18671,N_15228,N_13946);
or U18672 (N_18672,N_13790,N_14281);
xnor U18673 (N_18673,N_12998,N_15087);
nand U18674 (N_18674,N_12589,N_13536);
nand U18675 (N_18675,N_14594,N_14683);
nand U18676 (N_18676,N_15068,N_15468);
and U18677 (N_18677,N_15437,N_12694);
or U18678 (N_18678,N_14000,N_13454);
nor U18679 (N_18679,N_12933,N_12853);
nand U18680 (N_18680,N_14556,N_15442);
and U18681 (N_18681,N_14547,N_13083);
and U18682 (N_18682,N_15383,N_15270);
nor U18683 (N_18683,N_12663,N_13267);
and U18684 (N_18684,N_13911,N_13159);
and U18685 (N_18685,N_14736,N_13588);
or U18686 (N_18686,N_12957,N_14856);
or U18687 (N_18687,N_12597,N_12618);
nor U18688 (N_18688,N_14662,N_15290);
nor U18689 (N_18689,N_12690,N_14472);
xor U18690 (N_18690,N_15085,N_12857);
and U18691 (N_18691,N_13568,N_14146);
and U18692 (N_18692,N_14501,N_13286);
xnor U18693 (N_18693,N_14215,N_15595);
or U18694 (N_18694,N_15359,N_13665);
xor U18695 (N_18695,N_15480,N_14184);
xor U18696 (N_18696,N_13931,N_14147);
xnor U18697 (N_18697,N_12913,N_12921);
or U18698 (N_18698,N_14621,N_14265);
xnor U18699 (N_18699,N_14387,N_13643);
xnor U18700 (N_18700,N_14349,N_13655);
nor U18701 (N_18701,N_12557,N_14260);
nand U18702 (N_18702,N_13248,N_15621);
nor U18703 (N_18703,N_13164,N_15419);
xnor U18704 (N_18704,N_15596,N_13346);
or U18705 (N_18705,N_12880,N_14736);
and U18706 (N_18706,N_15133,N_12538);
nand U18707 (N_18707,N_14679,N_13752);
xor U18708 (N_18708,N_12874,N_12928);
nor U18709 (N_18709,N_13517,N_15575);
or U18710 (N_18710,N_13550,N_15099);
nand U18711 (N_18711,N_13163,N_13967);
or U18712 (N_18712,N_13145,N_14161);
or U18713 (N_18713,N_14548,N_14375);
nor U18714 (N_18714,N_12765,N_14911);
xnor U18715 (N_18715,N_13908,N_15308);
nand U18716 (N_18716,N_15485,N_14763);
xnor U18717 (N_18717,N_14733,N_13824);
xnor U18718 (N_18718,N_12997,N_14575);
nor U18719 (N_18719,N_14193,N_13510);
nand U18720 (N_18720,N_12795,N_13857);
and U18721 (N_18721,N_14699,N_14290);
xnor U18722 (N_18722,N_15569,N_15041);
xor U18723 (N_18723,N_15353,N_14330);
xor U18724 (N_18724,N_13219,N_13112);
and U18725 (N_18725,N_14816,N_14799);
or U18726 (N_18726,N_14733,N_13186);
xnor U18727 (N_18727,N_12634,N_13035);
or U18728 (N_18728,N_14200,N_15512);
nand U18729 (N_18729,N_13352,N_13892);
nand U18730 (N_18730,N_14436,N_13733);
xor U18731 (N_18731,N_14030,N_12556);
or U18732 (N_18732,N_14159,N_13932);
or U18733 (N_18733,N_14853,N_12990);
xnor U18734 (N_18734,N_13330,N_15485);
xnor U18735 (N_18735,N_12560,N_15586);
nand U18736 (N_18736,N_13900,N_13705);
or U18737 (N_18737,N_15121,N_15039);
nand U18738 (N_18738,N_13586,N_13538);
xor U18739 (N_18739,N_15241,N_12658);
nor U18740 (N_18740,N_13232,N_14679);
and U18741 (N_18741,N_13808,N_14201);
nand U18742 (N_18742,N_13737,N_15520);
or U18743 (N_18743,N_14662,N_15061);
xnor U18744 (N_18744,N_15041,N_15507);
nand U18745 (N_18745,N_14140,N_15491);
or U18746 (N_18746,N_13169,N_14548);
and U18747 (N_18747,N_13628,N_15544);
or U18748 (N_18748,N_12865,N_15585);
or U18749 (N_18749,N_12755,N_15525);
or U18750 (N_18750,N_15790,N_17346);
or U18751 (N_18751,N_17176,N_15978);
xor U18752 (N_18752,N_17776,N_17304);
xor U18753 (N_18753,N_16067,N_16188);
nand U18754 (N_18754,N_16644,N_18604);
nand U18755 (N_18755,N_18525,N_16918);
and U18756 (N_18756,N_17379,N_16261);
xor U18757 (N_18757,N_18008,N_15796);
and U18758 (N_18758,N_17539,N_16842);
or U18759 (N_18759,N_17545,N_16814);
xor U18760 (N_18760,N_16055,N_17127);
or U18761 (N_18761,N_17954,N_15879);
nor U18762 (N_18762,N_16401,N_16900);
or U18763 (N_18763,N_18541,N_17150);
xnor U18764 (N_18764,N_17745,N_17772);
and U18765 (N_18765,N_18291,N_18017);
nor U18766 (N_18766,N_16184,N_16137);
and U18767 (N_18767,N_18345,N_17731);
xnor U18768 (N_18768,N_17461,N_16048);
nor U18769 (N_18769,N_18386,N_18686);
and U18770 (N_18770,N_18088,N_16684);
or U18771 (N_18771,N_17746,N_17302);
xor U18772 (N_18772,N_17218,N_15820);
and U18773 (N_18773,N_16697,N_16078);
nand U18774 (N_18774,N_18420,N_18747);
and U18775 (N_18775,N_17674,N_16162);
xnor U18776 (N_18776,N_17944,N_16595);
and U18777 (N_18777,N_17178,N_18249);
xor U18778 (N_18778,N_16957,N_17006);
or U18779 (N_18779,N_16764,N_18623);
xor U18780 (N_18780,N_15913,N_17765);
and U18781 (N_18781,N_16369,N_16290);
and U18782 (N_18782,N_16452,N_17956);
or U18783 (N_18783,N_17925,N_17720);
nor U18784 (N_18784,N_17675,N_15749);
and U18785 (N_18785,N_15779,N_18699);
xnor U18786 (N_18786,N_16468,N_16110);
nor U18787 (N_18787,N_16765,N_18262);
xor U18788 (N_18788,N_16723,N_16377);
nand U18789 (N_18789,N_16938,N_17578);
nor U18790 (N_18790,N_18179,N_17982);
nand U18791 (N_18791,N_17484,N_18125);
and U18792 (N_18792,N_16703,N_16260);
nor U18793 (N_18793,N_16691,N_18584);
xnor U18794 (N_18794,N_16618,N_17732);
or U18795 (N_18795,N_17485,N_17316);
xnor U18796 (N_18796,N_18329,N_18535);
or U18797 (N_18797,N_16730,N_15739);
and U18798 (N_18798,N_18046,N_16302);
or U18799 (N_18799,N_18685,N_17777);
xor U18800 (N_18800,N_18078,N_15873);
xnor U18801 (N_18801,N_17350,N_16748);
or U18802 (N_18802,N_16913,N_15658);
nand U18803 (N_18803,N_17195,N_18471);
nand U18804 (N_18804,N_17865,N_15828);
nand U18805 (N_18805,N_17275,N_17128);
and U18806 (N_18806,N_18599,N_17964);
and U18807 (N_18807,N_17285,N_16872);
nand U18808 (N_18808,N_18193,N_17754);
or U18809 (N_18809,N_18229,N_16163);
xnor U18810 (N_18810,N_18530,N_16019);
or U18811 (N_18811,N_18305,N_18028);
nand U18812 (N_18812,N_16892,N_17743);
and U18813 (N_18813,N_15682,N_17473);
nor U18814 (N_18814,N_15912,N_16421);
xnor U18815 (N_18815,N_16641,N_16570);
or U18816 (N_18816,N_16733,N_18620);
and U18817 (N_18817,N_16683,N_18073);
xor U18818 (N_18818,N_17453,N_16330);
xnor U18819 (N_18819,N_18407,N_17175);
nor U18820 (N_18820,N_17198,N_18113);
or U18821 (N_18821,N_17038,N_15831);
nand U18822 (N_18822,N_18692,N_15845);
or U18823 (N_18823,N_17655,N_15667);
nand U18824 (N_18824,N_18368,N_17377);
and U18825 (N_18825,N_17976,N_18103);
nor U18826 (N_18826,N_18168,N_18134);
nor U18827 (N_18827,N_17605,N_16530);
or U18828 (N_18828,N_16996,N_17403);
or U18829 (N_18829,N_16665,N_16130);
and U18830 (N_18830,N_16845,N_17297);
and U18831 (N_18831,N_15850,N_17594);
or U18832 (N_18832,N_16364,N_15743);
and U18833 (N_18833,N_17154,N_18481);
nor U18834 (N_18834,N_17404,N_18352);
xnor U18835 (N_18835,N_15706,N_17309);
or U18836 (N_18836,N_18333,N_18534);
nand U18837 (N_18837,N_16075,N_15650);
nor U18838 (N_18838,N_16890,N_17244);
and U18839 (N_18839,N_18441,N_16399);
nand U18840 (N_18840,N_16552,N_15807);
nor U18841 (N_18841,N_17536,N_16874);
xor U18842 (N_18842,N_17519,N_15769);
and U18843 (N_18843,N_16158,N_17645);
and U18844 (N_18844,N_16967,N_17253);
nand U18845 (N_18845,N_17002,N_18739);
nor U18846 (N_18846,N_18332,N_18156);
xor U18847 (N_18847,N_18694,N_18722);
or U18848 (N_18848,N_16865,N_18278);
or U18849 (N_18849,N_18720,N_17026);
nor U18850 (N_18850,N_17805,N_16266);
nor U18851 (N_18851,N_17163,N_16018);
nand U18852 (N_18852,N_17395,N_17948);
and U18853 (N_18853,N_15712,N_15719);
nand U18854 (N_18854,N_16669,N_16170);
xor U18855 (N_18855,N_17567,N_15761);
nor U18856 (N_18856,N_17803,N_18299);
nand U18857 (N_18857,N_18337,N_17436);
and U18858 (N_18858,N_17882,N_18477);
and U18859 (N_18859,N_16455,N_16870);
xor U18860 (N_18860,N_16803,N_16152);
and U18861 (N_18861,N_16580,N_16529);
nand U18862 (N_18862,N_17718,N_16187);
nor U18863 (N_18863,N_17631,N_17854);
nand U18864 (N_18864,N_15781,N_17557);
xnor U18865 (N_18865,N_17546,N_15922);
nand U18866 (N_18866,N_16389,N_16471);
or U18867 (N_18867,N_18313,N_16275);
or U18868 (N_18868,N_16979,N_18309);
nand U18869 (N_18869,N_17156,N_17458);
nor U18870 (N_18870,N_15695,N_18085);
nand U18871 (N_18871,N_18612,N_17270);
xnor U18872 (N_18872,N_16607,N_18141);
or U18873 (N_18873,N_16658,N_16576);
and U18874 (N_18874,N_17866,N_17110);
or U18875 (N_18875,N_17372,N_17749);
or U18876 (N_18876,N_16951,N_16922);
xor U18877 (N_18877,N_16715,N_17054);
xor U18878 (N_18878,N_16398,N_15698);
or U18879 (N_18879,N_17817,N_16283);
or U18880 (N_18880,N_17587,N_18598);
xor U18881 (N_18881,N_15629,N_16177);
and U18882 (N_18882,N_17843,N_17035);
nand U18883 (N_18883,N_18216,N_17997);
or U18884 (N_18884,N_16749,N_17474);
nand U18885 (N_18885,N_16566,N_17575);
xor U18886 (N_18886,N_17688,N_16511);
and U18887 (N_18887,N_17554,N_17106);
nand U18888 (N_18888,N_15928,N_18413);
xnor U18889 (N_18889,N_15763,N_17367);
nor U18890 (N_18890,N_17602,N_16027);
and U18891 (N_18891,N_16481,N_17452);
and U18892 (N_18892,N_16277,N_15856);
xnor U18893 (N_18893,N_15877,N_16447);
nand U18894 (N_18894,N_16035,N_18116);
xor U18895 (N_18895,N_16439,N_18241);
or U18896 (N_18896,N_18126,N_17623);
nand U18897 (N_18897,N_17989,N_18095);
nor U18898 (N_18898,N_17293,N_17599);
nor U18899 (N_18899,N_16759,N_16961);
or U18900 (N_18900,N_17648,N_18399);
nand U18901 (N_18901,N_16560,N_17827);
and U18902 (N_18902,N_16171,N_16855);
and U18903 (N_18903,N_18220,N_16943);
xnor U18904 (N_18904,N_16994,N_17763);
xnor U18905 (N_18905,N_18167,N_16719);
or U18906 (N_18906,N_16798,N_15801);
nor U18907 (N_18907,N_17335,N_16857);
or U18908 (N_18908,N_16532,N_17024);
nor U18909 (N_18909,N_16516,N_17569);
and U18910 (N_18910,N_18568,N_18545);
nand U18911 (N_18911,N_17226,N_16449);
nand U18912 (N_18912,N_16174,N_18674);
or U18913 (N_18913,N_16651,N_17862);
xor U18914 (N_18914,N_17325,N_17928);
xnor U18915 (N_18915,N_17683,N_17751);
and U18916 (N_18916,N_17052,N_16136);
nand U18917 (N_18917,N_15919,N_17615);
and U18918 (N_18918,N_16375,N_17012);
xnor U18919 (N_18919,N_17931,N_16986);
nand U18920 (N_18920,N_16248,N_17913);
nor U18921 (N_18921,N_18411,N_16013);
or U18922 (N_18922,N_17238,N_17703);
or U18923 (N_18923,N_17523,N_17283);
and U18924 (N_18924,N_16592,N_18234);
xnor U18925 (N_18925,N_18667,N_18079);
and U18926 (N_18926,N_17081,N_15986);
xor U18927 (N_18927,N_18641,N_17585);
and U18928 (N_18928,N_18061,N_18364);
or U18929 (N_18929,N_18222,N_16555);
nand U18930 (N_18930,N_17040,N_18265);
nand U18931 (N_18931,N_16756,N_17492);
nand U18932 (N_18932,N_17728,N_16573);
nand U18933 (N_18933,N_16080,N_15925);
nor U18934 (N_18934,N_15728,N_18043);
nor U18935 (N_18935,N_18310,N_16939);
and U18936 (N_18936,N_15990,N_17894);
nand U18937 (N_18937,N_18202,N_17059);
nand U18938 (N_18938,N_16742,N_18675);
and U18939 (N_18939,N_16475,N_17247);
or U18940 (N_18940,N_16992,N_17103);
or U18941 (N_18941,N_17354,N_16643);
nand U18942 (N_18942,N_18024,N_18198);
and U18943 (N_18943,N_16254,N_16175);
xor U18944 (N_18944,N_16408,N_17830);
or U18945 (N_18945,N_16832,N_15776);
or U18946 (N_18946,N_17626,N_16229);
xor U18947 (N_18947,N_18225,N_17466);
nand U18948 (N_18948,N_16863,N_16244);
and U18949 (N_18949,N_15690,N_17034);
nor U18950 (N_18950,N_16598,N_18392);
or U18951 (N_18951,N_16538,N_16417);
and U18952 (N_18952,N_17885,N_17891);
nand U18953 (N_18953,N_15999,N_17971);
or U18954 (N_18954,N_18414,N_17242);
nor U18955 (N_18955,N_17193,N_17938);
nand U18956 (N_18956,N_15931,N_17442);
nor U18957 (N_18957,N_16826,N_17232);
nor U18958 (N_18958,N_18365,N_17482);
nor U18959 (N_18959,N_18665,N_18361);
or U18960 (N_18960,N_17203,N_15655);
nand U18961 (N_18961,N_18710,N_16639);
nor U18962 (N_18962,N_17700,N_17665);
nor U18963 (N_18963,N_18140,N_17916);
nand U18964 (N_18964,N_17300,N_16797);
and U18965 (N_18965,N_16213,N_16569);
nor U18966 (N_18966,N_15843,N_18741);
or U18967 (N_18967,N_18376,N_17062);
or U18968 (N_18968,N_16030,N_17291);
nand U18969 (N_18969,N_17676,N_16657);
xnor U18970 (N_18970,N_17868,N_16496);
xor U18971 (N_18971,N_18145,N_18176);
xor U18972 (N_18972,N_16628,N_18470);
nor U18973 (N_18973,N_18183,N_15899);
nand U18974 (N_18974,N_17699,N_15969);
xnor U18975 (N_18975,N_17747,N_16732);
nor U18976 (N_18976,N_17206,N_16325);
nor U18977 (N_18977,N_16624,N_17744);
and U18978 (N_18978,N_17561,N_18303);
nor U18979 (N_18979,N_16240,N_17196);
and U18980 (N_18980,N_18090,N_17902);
nor U18981 (N_18981,N_15971,N_18356);
xor U18982 (N_18982,N_16789,N_16501);
or U18983 (N_18983,N_18678,N_16740);
or U18984 (N_18984,N_16751,N_17422);
and U18985 (N_18985,N_16300,N_16739);
nor U18986 (N_18986,N_17651,N_18485);
or U18987 (N_18987,N_16396,N_18069);
and U18988 (N_18988,N_17426,N_18417);
and U18989 (N_18989,N_17121,N_17841);
nand U18990 (N_18990,N_16914,N_15907);
xor U18991 (N_18991,N_18260,N_18574);
and U18992 (N_18992,N_18185,N_18719);
xnor U18993 (N_18993,N_18314,N_17808);
nand U18994 (N_18994,N_15689,N_16824);
or U18995 (N_18995,N_18230,N_17089);
nand U18996 (N_18996,N_16862,N_18732);
nor U18997 (N_18997,N_18170,N_16489);
or U18998 (N_18998,N_18548,N_18657);
xor U18999 (N_18999,N_15939,N_17317);
or U19000 (N_19000,N_18203,N_15837);
nand U19001 (N_19001,N_16966,N_18276);
and U19002 (N_19002,N_17807,N_16426);
and U19003 (N_19003,N_16285,N_17467);
nand U19004 (N_19004,N_15984,N_17953);
and U19005 (N_19005,N_18245,N_15628);
xnor U19006 (N_19006,N_17601,N_16514);
or U19007 (N_19007,N_17368,N_17895);
nor U19008 (N_19008,N_17050,N_18362);
or U19009 (N_19009,N_17500,N_16921);
and U19010 (N_19010,N_17955,N_17071);
and U19011 (N_19011,N_17709,N_17382);
nor U19012 (N_19012,N_17217,N_16061);
nand U19013 (N_19013,N_18507,N_17952);
or U19014 (N_19014,N_16104,N_17767);
and U19015 (N_19015,N_16004,N_18591);
xnor U19016 (N_19016,N_16263,N_17820);
and U19017 (N_19017,N_16761,N_16512);
xor U19018 (N_19018,N_17396,N_17962);
or U19019 (N_19019,N_18503,N_15740);
and U19020 (N_19020,N_16689,N_17305);
xor U19021 (N_19021,N_18331,N_18552);
nand U19022 (N_19022,N_16526,N_16534);
or U19023 (N_19023,N_16677,N_18377);
nor U19024 (N_19024,N_16333,N_17656);
nand U19025 (N_19025,N_17251,N_17506);
nand U19026 (N_19026,N_17102,N_17907);
xnor U19027 (N_19027,N_17632,N_16473);
and U19028 (N_19028,N_16249,N_15847);
nor U19029 (N_19029,N_17398,N_18250);
and U19030 (N_19030,N_16477,N_18740);
nor U19031 (N_19031,N_17153,N_17834);
nor U19032 (N_19032,N_17490,N_18082);
xor U19033 (N_19033,N_18379,N_18738);
and U19034 (N_19034,N_18419,N_17996);
xor U19035 (N_19035,N_17873,N_16806);
and U19036 (N_19036,N_16387,N_16718);
nand U19037 (N_19037,N_15640,N_17311);
xnor U19038 (N_19038,N_17824,N_16919);
xnor U19039 (N_19039,N_16692,N_17282);
and U19040 (N_19040,N_16392,N_17710);
xnor U19041 (N_19041,N_16594,N_18606);
and U19042 (N_19042,N_16069,N_17503);
or U19043 (N_19043,N_17423,N_16975);
nand U19044 (N_19044,N_17137,N_17529);
or U19045 (N_19045,N_16391,N_15849);
and U19046 (N_19046,N_17541,N_17255);
xor U19047 (N_19047,N_17220,N_17294);
or U19048 (N_19048,N_16429,N_18318);
nor U19049 (N_19049,N_15888,N_18427);
and U19050 (N_19050,N_18253,N_18453);
nor U19051 (N_19051,N_18089,N_16344);
nand U19052 (N_19052,N_17845,N_16791);
or U19053 (N_19053,N_18464,N_18542);
nand U19054 (N_19054,N_16313,N_16207);
nor U19055 (N_19055,N_16154,N_18067);
xnor U19056 (N_19056,N_16005,N_18695);
xnor U19057 (N_19057,N_18280,N_15691);
xor U19058 (N_19058,N_16197,N_16853);
xor U19059 (N_19059,N_17850,N_16156);
and U19060 (N_19060,N_18371,N_16070);
nand U19061 (N_19061,N_18474,N_18281);
or U19062 (N_19062,N_17399,N_17618);
nand U19063 (N_19063,N_15935,N_18594);
and U19064 (N_19064,N_16107,N_17671);
and U19065 (N_19065,N_17409,N_17055);
and U19066 (N_19066,N_16120,N_17421);
nor U19067 (N_19067,N_16746,N_18160);
and U19068 (N_19068,N_17373,N_17307);
or U19069 (N_19069,N_16507,N_16049);
nand U19070 (N_19070,N_16402,N_16625);
and U19071 (N_19071,N_16852,N_16884);
xnor U19072 (N_19072,N_17721,N_18610);
or U19073 (N_19073,N_18522,N_16525);
nor U19074 (N_19074,N_17786,N_17277);
xor U19075 (N_19075,N_18486,N_16517);
or U19076 (N_19076,N_17796,N_17353);
xnor U19077 (N_19077,N_17172,N_16972);
and U19078 (N_19078,N_16485,N_17652);
and U19079 (N_19079,N_16617,N_18264);
nand U19080 (N_19080,N_17021,N_16584);
nor U19081 (N_19081,N_17117,N_16672);
nor U19082 (N_19082,N_17160,N_17550);
nor U19083 (N_19083,N_18235,N_18504);
xor U19084 (N_19084,N_17123,N_17861);
or U19085 (N_19085,N_15741,N_18120);
xor U19086 (N_19086,N_17933,N_16953);
and U19087 (N_19087,N_16458,N_18581);
nand U19088 (N_19088,N_15916,N_18493);
nand U19089 (N_19089,N_16166,N_17240);
and U19090 (N_19090,N_16499,N_16026);
nand U19091 (N_19091,N_17104,N_16822);
xor U19092 (N_19092,N_16747,N_15881);
xor U19093 (N_19093,N_18544,N_16542);
or U19094 (N_19094,N_18308,N_15909);
or U19095 (N_19095,N_16668,N_17464);
xnor U19096 (N_19096,N_17846,N_16502);
or U19097 (N_19097,N_16021,N_18445);
and U19098 (N_19098,N_16666,N_15675);
xnor U19099 (N_19099,N_16982,N_16472);
nor U19100 (N_19100,N_16415,N_17857);
nor U19101 (N_19101,N_15930,N_17290);
nor U19102 (N_19102,N_17066,N_18153);
and U19103 (N_19103,N_16101,N_16142);
xor U19104 (N_19104,N_17990,N_15768);
or U19105 (N_19105,N_17011,N_18239);
xnor U19106 (N_19106,N_17375,N_16370);
nand U19107 (N_19107,N_16381,N_15645);
and U19108 (N_19108,N_15630,N_17152);
xnor U19109 (N_19109,N_16423,N_17782);
and U19110 (N_19110,N_17004,N_18143);
nor U19111 (N_19111,N_16696,N_17323);
and U19112 (N_19112,N_17741,N_17249);
and U19113 (N_19113,N_17730,N_17598);
nor U19114 (N_19114,N_18723,N_17096);
nor U19115 (N_19115,N_15898,N_17540);
nor U19116 (N_19116,N_18139,N_18395);
nor U19117 (N_19117,N_15934,N_15653);
xor U19118 (N_19118,N_15734,N_17388);
and U19119 (N_19119,N_15832,N_15764);
nand U19120 (N_19120,N_17723,N_15681);
or U19121 (N_19121,N_17416,N_15733);
nand U19122 (N_19122,N_17331,N_18144);
nand U19123 (N_19123,N_18290,N_16947);
nor U19124 (N_19124,N_17658,N_17892);
nand U19125 (N_19125,N_17559,N_16636);
nand U19126 (N_19126,N_16902,N_16880);
and U19127 (N_19127,N_18721,N_15964);
or U19128 (N_19128,N_18633,N_16394);
and U19129 (N_19129,N_18171,N_17690);
and U19130 (N_19130,N_16016,N_18208);
xor U19131 (N_19131,N_16574,N_16821);
nor U19132 (N_19132,N_17061,N_16937);
and U19133 (N_19133,N_16486,N_15785);
nand U19134 (N_19134,N_18194,N_17789);
nand U19135 (N_19135,N_16647,N_16340);
xnor U19136 (N_19136,N_18547,N_18573);
xnor U19137 (N_19137,N_16988,N_18506);
or U19138 (N_19138,N_18055,N_15885);
xor U19139 (N_19139,N_18593,N_17852);
and U19140 (N_19140,N_17164,N_18304);
nor U19141 (N_19141,N_17480,N_16233);
nand U19142 (N_19142,N_17194,N_16589);
or U19143 (N_19143,N_16906,N_16056);
nor U19144 (N_19144,N_17397,N_17687);
xor U19145 (N_19145,N_18688,N_16653);
nand U19146 (N_19146,N_17448,N_16359);
nand U19147 (N_19147,N_17667,N_17909);
nand U19148 (N_19148,N_18439,N_17994);
or U19149 (N_19149,N_16823,N_15694);
nand U19150 (N_19150,N_17241,N_16114);
nand U19151 (N_19151,N_18524,N_16817);
nor U19152 (N_19152,N_16442,N_18161);
nor U19153 (N_19153,N_17447,N_18714);
nor U19154 (N_19154,N_17814,N_18000);
nand U19155 (N_19155,N_17552,N_17572);
nand U19156 (N_19156,N_17494,N_18131);
and U19157 (N_19157,N_18020,N_18023);
or U19158 (N_19158,N_17433,N_18048);
nor U19159 (N_19159,N_18472,N_17424);
nand U19160 (N_19160,N_18068,N_16384);
or U19161 (N_19161,N_18187,N_18513);
and U19162 (N_19162,N_17308,N_18444);
or U19163 (N_19163,N_18270,N_17950);
or U19164 (N_19164,N_16637,N_17941);
or U19165 (N_19165,N_17093,N_18554);
xnor U19166 (N_19166,N_18261,N_17243);
or U19167 (N_19167,N_16716,N_18076);
and U19168 (N_19168,N_16737,N_16802);
nand U19169 (N_19169,N_18580,N_15692);
nand U19170 (N_19170,N_18698,N_17312);
and U19171 (N_19171,N_17125,N_18360);
and U19172 (N_19172,N_16282,N_17187);
and U19173 (N_19173,N_18502,N_15824);
xor U19174 (N_19174,N_16204,N_15862);
nor U19175 (N_19175,N_16571,N_17622);
or U19176 (N_19176,N_15905,N_16024);
nand U19177 (N_19177,N_15810,N_18070);
and U19178 (N_19178,N_17060,N_17517);
nand U19179 (N_19179,N_17074,N_17274);
or U19180 (N_19180,N_16433,N_16453);
nor U19181 (N_19181,N_18433,N_16276);
nand U19182 (N_19182,N_17223,N_17836);
or U19183 (N_19183,N_18372,N_16050);
nor U19184 (N_19184,N_17009,N_16941);
nand U19185 (N_19185,N_17704,N_16729);
nand U19186 (N_19186,N_17879,N_17965);
nand U19187 (N_19187,N_16117,N_15738);
nor U19188 (N_19188,N_17405,N_18045);
or U19189 (N_19189,N_17670,N_17239);
nor U19190 (N_19190,N_17625,N_16338);
nor U19191 (N_19191,N_16998,N_15880);
and U19192 (N_19192,N_17215,N_17580);
nor U19193 (N_19193,N_16882,N_16172);
nor U19194 (N_19194,N_17046,N_16456);
nand U19195 (N_19195,N_16416,N_18124);
nand U19196 (N_19196,N_17105,N_15980);
nor U19197 (N_19197,N_16124,N_15730);
or U19198 (N_19198,N_18560,N_17742);
and U19199 (N_19199,N_16971,N_16168);
nor U19200 (N_19200,N_16693,N_16504);
nor U19201 (N_19201,N_17619,N_18326);
and U19202 (N_19202,N_16378,N_18159);
nand U19203 (N_19203,N_17787,N_16958);
xor U19204 (N_19204,N_16459,N_16128);
nor U19205 (N_19205,N_17949,N_15863);
nand U19206 (N_19206,N_18190,N_18680);
nand U19207 (N_19207,N_17413,N_18663);
and U19208 (N_19208,N_16631,N_18632);
and U19209 (N_19209,N_16133,N_18035);
nor U19210 (N_19210,N_17514,N_17600);
or U19211 (N_19211,N_17930,N_15715);
nor U19212 (N_19212,N_18147,N_17161);
and U19213 (N_19213,N_17037,N_18520);
or U19214 (N_19214,N_18370,N_18283);
nand U19215 (N_19215,N_16084,N_17917);
nor U19216 (N_19216,N_15709,N_18173);
or U19217 (N_19217,N_18182,N_16605);
or U19218 (N_19218,N_17927,N_16609);
nor U19219 (N_19219,N_17092,N_16058);
or U19220 (N_19220,N_16878,N_18683);
nand U19221 (N_19221,N_17534,N_16790);
nand U19222 (N_19222,N_16879,N_16769);
nor U19223 (N_19223,N_18162,N_18514);
or U19224 (N_19224,N_17008,N_16328);
xor U19225 (N_19225,N_16224,N_17993);
nand U19226 (N_19226,N_17593,N_15783);
or U19227 (N_19227,N_16036,N_17007);
nor U19228 (N_19228,N_16936,N_17822);
xnor U19229 (N_19229,N_17985,N_16616);
or U19230 (N_19230,N_15747,N_15816);
nor U19231 (N_19231,N_17190,N_17015);
nand U19232 (N_19232,N_17488,N_15883);
xnor U19233 (N_19233,N_18592,N_17165);
xor U19234 (N_19234,N_16661,N_18224);
and U19235 (N_19235,N_17087,N_17493);
and U19236 (N_19236,N_18529,N_15826);
or U19237 (N_19237,N_17418,N_15817);
xnor U19238 (N_19238,N_17498,N_16850);
or U19239 (N_19239,N_16564,N_16536);
xnor U19240 (N_19240,N_18661,N_16519);
xor U19241 (N_19241,N_17348,N_17736);
nand U19242 (N_19242,N_17823,N_18049);
or U19243 (N_19243,N_18666,N_18018);
nand U19244 (N_19244,N_15631,N_15742);
nand U19245 (N_19245,N_18518,N_16169);
or U19246 (N_19246,N_17935,N_16220);
and U19247 (N_19247,N_17961,N_15647);
nor U19248 (N_19248,N_16498,N_17288);
nand U19249 (N_19249,N_17281,N_18717);
nand U19250 (N_19250,N_17570,N_18232);
and U19251 (N_19251,N_17511,N_18174);
xnor U19252 (N_19252,N_16917,N_16029);
xor U19253 (N_19253,N_17677,N_16373);
and U19254 (N_19254,N_16216,N_16102);
nand U19255 (N_19255,N_18437,N_17264);
nor U19256 (N_19256,N_16811,N_17968);
or U19257 (N_19257,N_15657,N_18032);
or U19258 (N_19258,N_16704,N_18645);
or U19259 (N_19259,N_16222,N_16281);
or U19260 (N_19260,N_16911,N_18551);
nand U19261 (N_19261,N_18373,N_16854);
xnor U19262 (N_19262,N_18629,N_16363);
nor U19263 (N_19263,N_16227,N_17100);
xor U19264 (N_19264,N_16757,N_15882);
xnor U19265 (N_19265,N_17155,N_18509);
nand U19266 (N_19266,N_17644,N_15937);
nand U19267 (N_19267,N_16970,N_18307);
or U19268 (N_19268,N_16296,N_15659);
nand U19269 (N_19269,N_18354,N_17722);
or U19270 (N_19270,N_18521,N_15987);
or U19271 (N_19271,N_15721,N_15656);
nor U19272 (N_19272,N_18027,N_18064);
or U19273 (N_19273,N_18696,N_18091);
nand U19274 (N_19274,N_17044,N_18127);
and U19275 (N_19275,N_17973,N_18549);
or U19276 (N_19276,N_16183,N_17998);
or U19277 (N_19277,N_16242,N_17696);
or U19278 (N_19278,N_18536,N_15977);
or U19279 (N_19279,N_18204,N_16223);
nand U19280 (N_19280,N_18094,N_18083);
and U19281 (N_19281,N_17179,N_17435);
or U19282 (N_19282,N_16195,N_16563);
nand U19283 (N_19283,N_17412,N_16527);
nor U19284 (N_19284,N_18642,N_18065);
xor U19285 (N_19285,N_16259,N_18300);
xor U19286 (N_19286,N_18404,N_17717);
xnor U19287 (N_19287,N_18567,N_16727);
and U19288 (N_19288,N_16482,N_17266);
or U19289 (N_19289,N_18480,N_16366);
nand U19290 (N_19290,N_18650,N_18748);
or U19291 (N_19291,N_16268,N_17438);
or U19292 (N_19292,N_17337,N_16308);
nor U19293 (N_19293,N_18537,N_18442);
nor U19294 (N_19294,N_17637,N_18213);
nor U19295 (N_19295,N_17064,N_15693);
or U19296 (N_19296,N_17278,N_16648);
nor U19297 (N_19297,N_16767,N_15662);
nand U19298 (N_19298,N_18689,N_16780);
or U19299 (N_19299,N_18077,N_18109);
xor U19300 (N_19300,N_17298,N_16464);
nand U19301 (N_19301,N_17849,N_18031);
nor U19302 (N_19302,N_15685,N_15735);
and U19303 (N_19303,N_18684,N_16776);
nor U19304 (N_19304,N_16303,N_17538);
or U19305 (N_19305,N_16888,N_17781);
xor U19306 (N_19306,N_16834,N_16664);
nand U19307 (N_19307,N_17785,N_16141);
or U19308 (N_19308,N_17505,N_16923);
nand U19309 (N_19309,N_16934,N_16773);
or U19310 (N_19310,N_18558,N_18041);
and U19311 (N_19311,N_15771,N_17326);
and U19312 (N_19312,N_16243,N_17900);
or U19313 (N_19313,N_17793,N_17136);
nand U19314 (N_19314,N_17496,N_16813);
and U19315 (N_19315,N_17522,N_17333);
xnor U19316 (N_19316,N_17926,N_17975);
nor U19317 (N_19317,N_16755,N_17792);
and U19318 (N_19318,N_17666,N_16997);
or U19319 (N_19319,N_16079,N_17662);
and U19320 (N_19320,N_17812,N_17945);
or U19321 (N_19321,N_17947,N_17649);
or U19322 (N_19322,N_16535,N_18679);
and U19323 (N_19323,N_18426,N_16210);
nor U19324 (N_19324,N_15963,N_16688);
or U19325 (N_19325,N_15962,N_16006);
or U19326 (N_19326,N_17932,N_16403);
and U19327 (N_19327,N_18543,N_16710);
xor U19328 (N_19328,N_15664,N_15637);
xor U19329 (N_19329,N_18409,N_18637);
xor U19330 (N_19330,N_17692,N_16062);
or U19331 (N_19331,N_15994,N_18112);
nor U19332 (N_19332,N_16521,N_17359);
xor U19333 (N_19333,N_18293,N_15988);
and U19334 (N_19334,N_18500,N_18708);
and U19335 (N_19335,N_17088,N_16280);
nand U19336 (N_19336,N_17431,N_16219);
nand U19337 (N_19337,N_17289,N_18335);
xor U19338 (N_19338,N_16008,N_17564);
and U19339 (N_19339,N_15891,N_16901);
nor U19340 (N_19340,N_18093,N_17831);
xor U19341 (N_19341,N_15901,N_17755);
and U19342 (N_19342,N_16599,N_17299);
or U19343 (N_19343,N_15711,N_18431);
or U19344 (N_19344,N_16237,N_15677);
nand U19345 (N_19345,N_17313,N_17725);
nor U19346 (N_19346,N_18106,N_16371);
nor U19347 (N_19347,N_15857,N_16272);
nand U19348 (N_19348,N_18033,N_17988);
nor U19349 (N_19349,N_16082,N_16662);
or U19350 (N_19350,N_16097,N_16738);
xnor U19351 (N_19351,N_15992,N_17981);
nor U19352 (N_19352,N_17851,N_15720);
and U19353 (N_19353,N_15802,N_15947);
xnor U19354 (N_19354,N_18646,N_16645);
and U19355 (N_19355,N_16553,N_16505);
or U19356 (N_19356,N_18231,N_18624);
xor U19357 (N_19357,N_17679,N_16708);
nand U19358 (N_19358,N_17358,N_17528);
xnor U19359 (N_19359,N_15940,N_15893);
xnor U19360 (N_19360,N_16575,N_18374);
xnor U19361 (N_19361,N_17250,N_16491);
or U19362 (N_19362,N_18517,N_18080);
nand U19363 (N_19363,N_17795,N_17076);
xor U19364 (N_19364,N_15757,N_18512);
nor U19365 (N_19365,N_17957,N_17939);
nor U19366 (N_19366,N_16129,N_18669);
xor U19367 (N_19367,N_17257,N_17260);
nand U19368 (N_19368,N_15704,N_16985);
nor U19369 (N_19369,N_15746,N_17635);
nand U19370 (N_19370,N_17364,N_18589);
or U19371 (N_19371,N_17750,N_16293);
or U19372 (N_19372,N_17295,N_15737);
and U19373 (N_19373,N_18658,N_16218);
xor U19374 (N_19374,N_16987,N_18617);
nand U19375 (N_19375,N_18746,N_18728);
xnor U19376 (N_19376,N_16072,N_15663);
xor U19377 (N_19377,N_16270,N_16225);
and U19378 (N_19378,N_16588,N_16581);
nor U19379 (N_19379,N_18288,N_17036);
or U19380 (N_19380,N_15997,N_18330);
nor U19381 (N_19381,N_17049,N_17376);
or U19382 (N_19382,N_17177,N_18351);
xnor U19383 (N_19383,N_17157,N_16428);
nand U19384 (N_19384,N_16777,N_17181);
and U19385 (N_19385,N_18030,N_18550);
xnor U19386 (N_19386,N_16579,N_18191);
xor U19387 (N_19387,N_17880,N_17272);
or U19388 (N_19388,N_18359,N_16619);
nor U19389 (N_19389,N_18217,N_18454);
nand U19390 (N_19390,N_18559,N_17604);
and U19391 (N_19391,N_16954,N_16724);
nor U19392 (N_19392,N_16274,N_16745);
nor U19393 (N_19393,N_17606,N_16386);
xor U19394 (N_19394,N_16071,N_18478);
nand U19395 (N_19395,N_17429,N_15811);
nand U19396 (N_19396,N_15639,N_18210);
nand U19397 (N_19397,N_18460,N_16074);
nand U19398 (N_19398,N_17018,N_16413);
nor U19399 (N_19399,N_15967,N_16446);
and U19400 (N_19400,N_16681,N_17122);
and U19401 (N_19401,N_18393,N_16151);
xor U19402 (N_19402,N_18448,N_16318);
xnor U19403 (N_19403,N_18366,N_16908);
xnor U19404 (N_19404,N_17419,N_17086);
nor U19405 (N_19405,N_18556,N_16964);
nor U19406 (N_19406,N_17205,N_17908);
nor U19407 (N_19407,N_15989,N_16469);
or U19408 (N_19408,N_16076,N_16356);
xnor U19409 (N_19409,N_16596,N_16652);
xnor U19410 (N_19410,N_16457,N_16467);
nor U19411 (N_19411,N_17224,N_16810);
nand U19412 (N_19412,N_17057,N_16762);
xor U19413 (N_19413,N_17871,N_16940);
and U19414 (N_19414,N_17689,N_15732);
nor U19415 (N_19415,N_18286,N_18575);
and U19416 (N_19416,N_16991,N_17292);
or U19417 (N_19417,N_16753,N_18451);
nand U19418 (N_19418,N_16040,N_17329);
nand U19419 (N_19419,N_16623,N_17799);
nand U19420 (N_19420,N_15726,N_16314);
or U19421 (N_19421,N_17596,N_16606);
xnor U19422 (N_19422,N_17821,N_16087);
or U19423 (N_19423,N_18489,N_18175);
nor U19424 (N_19424,N_17607,N_18107);
and U19425 (N_19425,N_18292,N_17355);
nor U19426 (N_19426,N_16420,N_18284);
nor U19427 (N_19427,N_17958,N_18749);
nor U19428 (N_19428,N_16509,N_15762);
nor U19429 (N_19429,N_17000,N_18651);
xnor U19430 (N_19430,N_17904,N_18342);
or U19431 (N_19431,N_16676,N_17586);
nand U19432 (N_19432,N_18060,N_15825);
nand U19433 (N_19433,N_17963,N_15970);
nor U19434 (N_19434,N_15791,N_17231);
nand U19435 (N_19435,N_16840,N_17548);
nor U19436 (N_19436,N_16770,N_17462);
and U19437 (N_19437,N_18189,N_17469);
nand U19438 (N_19438,N_17780,N_16812);
or U19439 (N_19439,N_15927,N_17245);
xor U19440 (N_19440,N_17487,N_17112);
nor U19441 (N_19441,N_18713,N_18609);
nor U19442 (N_19442,N_17972,N_16194);
nor U19443 (N_19443,N_17825,N_17562);
nor U19444 (N_19444,N_17597,N_16500);
nor U19445 (N_19445,N_16685,N_17174);
nand U19446 (N_19446,N_18122,N_18271);
nor U19447 (N_19447,N_17135,N_16608);
and U19448 (N_19448,N_15686,N_16109);
and U19449 (N_19449,N_16436,N_18226);
nand U19450 (N_19450,N_16173,N_16465);
nor U19451 (N_19451,N_17207,N_18476);
nor U19452 (N_19452,N_18233,N_18214);
nor U19453 (N_19453,N_15646,N_17186);
nor U19454 (N_19454,N_17695,N_16835);
and U19455 (N_19455,N_16531,N_16711);
and U19456 (N_19456,N_15627,N_18618);
xnor U19457 (N_19457,N_17811,N_18062);
nor U19458 (N_19458,N_16434,N_15854);
and U19459 (N_19459,N_17627,N_16157);
or U19460 (N_19460,N_17073,N_15789);
nand U19461 (N_19461,N_17284,N_18257);
xor U19462 (N_19462,N_16032,N_15958);
nor U19463 (N_19463,N_15788,N_16602);
nor U19464 (N_19464,N_17028,N_17508);
nand U19465 (N_19465,N_17872,N_16887);
nor U19466 (N_19466,N_16950,N_18627);
and U19467 (N_19467,N_16337,N_16134);
and U19468 (N_19468,N_18533,N_18129);
nand U19469 (N_19469,N_16786,N_17848);
xor U19470 (N_19470,N_15979,N_17013);
and U19471 (N_19471,N_16952,N_15775);
nor U19472 (N_19472,N_17609,N_18608);
nor U19473 (N_19473,N_16963,N_16066);
and U19474 (N_19474,N_15915,N_16883);
or U19475 (N_19475,N_16445,N_17919);
or U19476 (N_19476,N_16347,N_17146);
and U19477 (N_19477,N_17440,N_15727);
or U19478 (N_19478,N_18677,N_18058);
nand U19479 (N_19479,N_17478,N_16912);
xor U19480 (N_19480,N_18341,N_16698);
nor U19481 (N_19481,N_17078,N_16319);
nor U19482 (N_19482,N_17672,N_15836);
xor U19483 (N_19483,N_18724,N_16354);
nand U19484 (N_19484,N_17896,N_17167);
xnor U19485 (N_19485,N_18155,N_18311);
or U19486 (N_19486,N_18390,N_18440);
nand U19487 (N_19487,N_17370,N_16875);
or U19488 (N_19488,N_18295,N_16965);
nor U19489 (N_19489,N_15773,N_17204);
nand U19490 (N_19490,N_15892,N_18488);
xnor U19491 (N_19491,N_18243,N_16962);
or U19492 (N_19492,N_16041,N_17212);
or U19493 (N_19493,N_17608,N_15670);
or U19494 (N_19494,N_16787,N_18421);
xnor U19495 (N_19495,N_16886,N_16920);
and U19496 (N_19496,N_17338,N_18597);
nand U19497 (N_19497,N_17434,N_18227);
and U19498 (N_19498,N_18511,N_16694);
xnor U19499 (N_19499,N_16678,N_15814);
or U19500 (N_19500,N_16192,N_16196);
nand U19501 (N_19501,N_17636,N_17769);
xor U19502 (N_19502,N_18242,N_17149);
or U19503 (N_19503,N_15945,N_18571);
nor U19504 (N_19504,N_16077,N_18003);
or U19505 (N_19505,N_17653,N_17783);
or U19506 (N_19506,N_16148,N_16198);
xor U19507 (N_19507,N_18151,N_17171);
nor U19508 (N_19508,N_17216,N_18343);
or U19509 (N_19509,N_17027,N_18044);
nand U19510 (N_19510,N_15765,N_18118);
nor U19511 (N_19511,N_17685,N_15813);
nor U19512 (N_19512,N_16524,N_18561);
nand U19513 (N_19513,N_16208,N_17320);
xor U19514 (N_19514,N_16493,N_17535);
or U19515 (N_19515,N_18670,N_16804);
nor U19516 (N_19516,N_15815,N_18654);
nand U19517 (N_19517,N_16860,N_16794);
or U19518 (N_19518,N_18375,N_17643);
or U19519 (N_19519,N_18693,N_15684);
xor U19520 (N_19520,N_15902,N_16284);
nor U19521 (N_19521,N_17048,N_18682);
or U19522 (N_19522,N_18465,N_18398);
xor U19523 (N_19523,N_18466,N_18705);
nor U19524 (N_19524,N_16989,N_15809);
nand U19525 (N_19525,N_16217,N_16744);
nor U19526 (N_19526,N_17124,N_15860);
and U19527 (N_19527,N_16712,N_16916);
nand U19528 (N_19528,N_16831,N_17715);
xnor U19529 (N_19529,N_18499,N_17225);
nand U19530 (N_19530,N_17937,N_17099);
xor U19531 (N_19531,N_17483,N_18207);
xnor U19532 (N_19532,N_16721,N_17719);
or U19533 (N_19533,N_15672,N_15792);
nand U19534 (N_19534,N_16924,N_18218);
or U19535 (N_19535,N_18306,N_16153);
nand U19536 (N_19536,N_15699,N_18539);
and U19537 (N_19537,N_17842,N_16868);
xor U19538 (N_19538,N_18338,N_16815);
nand U19539 (N_19539,N_18647,N_17791);
nand U19540 (N_19540,N_15777,N_17591);
or U19541 (N_19541,N_17457,N_16135);
nor U19542 (N_19542,N_15806,N_16830);
or U19543 (N_19543,N_16633,N_17713);
or U19544 (N_19544,N_15722,N_18557);
nor U19545 (N_19545,N_18690,N_16792);
nor U19546 (N_19546,N_17801,N_17708);
xnor U19547 (N_19547,N_16339,N_17518);
xnor U19548 (N_19548,N_18132,N_17693);
and U19549 (N_19549,N_16051,N_16065);
or U19550 (N_19550,N_17735,N_18117);
or U19551 (N_19551,N_18643,N_18635);
and U19552 (N_19552,N_16081,N_16903);
and U19553 (N_19553,N_16587,N_17802);
nand U19554 (N_19554,N_16001,N_17261);
or U19555 (N_19555,N_18206,N_17761);
nor U19556 (N_19556,N_17051,N_16660);
nand U19557 (N_19557,N_17612,N_16113);
or U19558 (N_19558,N_16709,N_16028);
or U19559 (N_19559,N_18267,N_15961);
nand U19560 (N_19560,N_17169,N_16871);
xnor U19561 (N_19561,N_18215,N_17533);
xnor U19562 (N_19562,N_16766,N_16546);
or U19563 (N_19563,N_16788,N_17058);
and U19564 (N_19564,N_16278,N_16342);
nand U19565 (N_19565,N_16298,N_18546);
and U19566 (N_19566,N_18586,N_16981);
and U19567 (N_19567,N_16893,N_17633);
nand U19568 (N_19568,N_18001,N_18712);
nand U19569 (N_19569,N_15835,N_16310);
xnor U19570 (N_19570,N_18378,N_15636);
and U19571 (N_19571,N_16973,N_15900);
and U19572 (N_19572,N_18729,N_18515);
nand U19573 (N_19573,N_18154,N_16206);
and U19574 (N_19574,N_16935,N_16349);
nand U19575 (N_19575,N_15723,N_16848);
xor U19576 (N_19576,N_17840,N_16116);
xnor U19577 (N_19577,N_17610,N_16382);
xnor U19578 (N_19578,N_16007,N_16583);
nand U19579 (N_19579,N_16063,N_15756);
and U19580 (N_19580,N_17042,N_17884);
or U19581 (N_19581,N_16425,N_16627);
nor U19582 (N_19582,N_16343,N_17443);
nand U19583 (N_19583,N_16215,N_17869);
or U19584 (N_19584,N_17694,N_16269);
nand U19585 (N_19585,N_16232,N_17911);
nor U19586 (N_19586,N_15869,N_18621);
or U19587 (N_19587,N_16760,N_18328);
or U19588 (N_19588,N_18051,N_17211);
and U19589 (N_19589,N_16422,N_17098);
nor U19590 (N_19590,N_17402,N_18744);
and U19591 (N_19591,N_17085,N_16544);
nor U19592 (N_19592,N_17682,N_16397);
xor U19593 (N_19593,N_17729,N_18201);
or U19594 (N_19594,N_17481,N_16212);
xnor U19595 (N_19595,N_16483,N_16199);
nor U19596 (N_19596,N_17887,N_17660);
nand U19597 (N_19597,N_17680,N_16699);
nor U19598 (N_19598,N_15804,N_17737);
and U19599 (N_19599,N_18479,N_16106);
nand U19600 (N_19600,N_17966,N_16155);
nand U19601 (N_19601,N_17940,N_16758);
nor U19602 (N_19602,N_18492,N_16138);
or U19603 (N_19603,N_17657,N_17959);
nand U19604 (N_19604,N_18047,N_16725);
nand U19605 (N_19605,N_18272,N_17936);
and U19606 (N_19606,N_16054,N_18172);
xnor U19607 (N_19607,N_16348,N_16889);
xnor U19608 (N_19608,N_16376,N_18010);
nor U19609 (N_19609,N_17544,N_15688);
nor U19610 (N_19610,N_18491,N_18668);
or U19611 (N_19611,N_16031,N_17525);
xnor U19612 (N_19612,N_17979,N_16185);
and U19613 (N_19613,N_15871,N_16849);
nor U19614 (N_19614,N_18579,N_15795);
or U19615 (N_19615,N_15866,N_16289);
xnor U19616 (N_19616,N_15941,N_17507);
nand U19617 (N_19617,N_18057,N_16039);
nand U19618 (N_19618,N_18184,N_16640);
and U19619 (N_19619,N_18071,N_15904);
xor U19620 (N_19620,N_16086,N_17045);
and U19621 (N_19621,N_17810,N_16122);
xnor U19622 (N_19622,N_17033,N_15952);
and U19623 (N_19623,N_16508,N_18148);
xor U19624 (N_19624,N_17923,N_16412);
nand U19625 (N_19625,N_15911,N_17858);
xnor U19626 (N_19626,N_17332,N_17389);
or U19627 (N_19627,N_16059,N_16012);
xor U19628 (N_19628,N_18128,N_17445);
or U19629 (N_19629,N_18301,N_15957);
or U19630 (N_19630,N_17118,N_16334);
nor U19631 (N_19631,N_17444,N_18369);
nand U19632 (N_19632,N_15736,N_18367);
or U19633 (N_19633,N_16480,N_16118);
nor U19634 (N_19634,N_18634,N_16165);
xnor U19635 (N_19635,N_17143,N_18394);
and U19636 (N_19636,N_15830,N_17890);
or U19637 (N_19637,N_16235,N_17532);
and U19638 (N_19638,N_16713,N_17477);
or U19639 (N_19639,N_16929,N_17394);
nor U19640 (N_19640,N_18468,N_16722);
or U19641 (N_19641,N_16182,N_17509);
and U19642 (N_19642,N_17855,N_18246);
and U19643 (N_19643,N_15886,N_15926);
nand U19644 (N_19644,N_15839,N_17120);
xnor U19645 (N_19645,N_17091,N_15751);
nand U19646 (N_19646,N_16825,N_16424);
and U19647 (N_19647,N_18495,N_18195);
xnor U19648 (N_19648,N_18736,N_16667);
nand U19649 (N_19649,N_16547,N_18498);
xnor U19650 (N_19650,N_17408,N_18578);
or U19651 (N_19651,N_17142,N_17878);
nand U19652 (N_19652,N_15661,N_15651);
or U19653 (N_19653,N_18673,N_16324);
and U19654 (N_19654,N_18277,N_17571);
or U19655 (N_19655,N_16611,N_16956);
nand U19656 (N_19656,N_18285,N_18432);
or U19657 (N_19657,N_18279,N_17771);
nand U19658 (N_19658,N_16461,N_17459);
nand U19659 (N_19659,N_16479,N_16360);
and U19660 (N_19660,N_17800,N_16968);
nand U19661 (N_19661,N_18007,N_17809);
nor U19662 (N_19662,N_18209,N_16497);
and U19663 (N_19663,N_18348,N_16726);
xnor U19664 (N_19664,N_18403,N_18562);
or U19665 (N_19665,N_16649,N_18396);
nand U19666 (N_19666,N_16771,N_15669);
or U19667 (N_19667,N_16663,N_17425);
xnor U19668 (N_19668,N_16085,N_16638);
nor U19669 (N_19669,N_16818,N_15942);
and U19670 (N_19670,N_18588,N_16323);
nand U19671 (N_19671,N_15634,N_17838);
or U19672 (N_19672,N_17835,N_16351);
and U19673 (N_19673,N_16690,N_15705);
and U19674 (N_19674,N_18240,N_16864);
xor U19675 (N_19675,N_16897,N_15652);
xor U19676 (N_19676,N_16558,N_16221);
and U19677 (N_19677,N_15760,N_17067);
xnor U19678 (N_19678,N_18505,N_17016);
or U19679 (N_19679,N_17479,N_18607);
or U19680 (N_19680,N_17410,N_15724);
or U19681 (N_19681,N_18602,N_18186);
nor U19682 (N_19682,N_17213,N_15641);
xnor U19683 (N_19683,N_15910,N_16980);
and U19684 (N_19684,N_15955,N_16119);
nor U19685 (N_19685,N_16291,N_18631);
xor U19686 (N_19686,N_18052,N_16948);
xnor U19687 (N_19687,N_16253,N_16586);
or U19688 (N_19688,N_18251,N_16236);
nor U19689 (N_19689,N_18648,N_16095);
and U19690 (N_19690,N_17563,N_17390);
or U19691 (N_19691,N_15772,N_16393);
and U19692 (N_19692,N_15972,N_18735);
xnor U19693 (N_19693,N_16800,N_16488);
or U19694 (N_19694,N_16494,N_18269);
and U19695 (N_19695,N_18672,N_18576);
xor U19696 (N_19696,N_17202,N_17365);
or U19697 (N_19697,N_16925,N_18259);
xnor U19698 (N_19698,N_16045,N_17188);
xnor U19699 (N_19699,N_16717,N_17141);
nor U19700 (N_19700,N_16352,N_18111);
nor U19701 (N_19701,N_17726,N_16686);
xor U19702 (N_19702,N_18026,N_17856);
and U19703 (N_19703,N_17621,N_18563);
nor U19704 (N_19704,N_18037,N_18424);
nor U19705 (N_19705,N_16930,N_18258);
xnor U19706 (N_19706,N_15635,N_17951);
and U19707 (N_19707,N_16513,N_16774);
nor U19708 (N_19708,N_18228,N_15654);
nand U19709 (N_19709,N_18715,N_17228);
nor U19710 (N_19710,N_16350,N_17759);
nor U19711 (N_19711,N_17180,N_16140);
xnor U19712 (N_19712,N_17942,N_17263);
xor U19713 (N_19713,N_16549,N_16368);
nor U19714 (N_19714,N_17788,N_17072);
and U19715 (N_19715,N_17774,N_18266);
nor U19716 (N_19716,N_16557,N_15846);
nand U19717 (N_19717,N_16752,N_16201);
and U19718 (N_19718,N_17144,N_18555);
nor U19719 (N_19719,N_18572,N_17491);
or U19720 (N_19720,N_18566,N_17197);
nor U19721 (N_19721,N_16160,N_17502);
nor U19722 (N_19722,N_17558,N_17097);
nor U19723 (N_19723,N_16894,N_15867);
nor U19724 (N_19724,N_18254,N_18430);
nand U19725 (N_19725,N_18164,N_15903);
xnor U19726 (N_19726,N_18435,N_18423);
or U19727 (N_19727,N_16910,N_17455);
nor U19728 (N_19728,N_18274,N_16038);
nand U19729 (N_19729,N_15758,N_17991);
xor U19730 (N_19730,N_18349,N_17929);
and U19731 (N_19731,N_16895,N_16271);
nor U19732 (N_19732,N_17960,N_18709);
xor U19733 (N_19733,N_15951,N_15803);
xor U19734 (N_19734,N_18158,N_17757);
and U19735 (N_19735,N_17537,N_16112);
or U19736 (N_19736,N_17430,N_18034);
nor U19737 (N_19737,N_17336,N_17616);
and U19738 (N_19738,N_17271,N_17381);
or U19739 (N_19739,N_17330,N_17020);
nand U19740 (N_19740,N_17259,N_16675);
nand U19741 (N_19741,N_17287,N_16768);
and U19742 (N_19742,N_16642,N_17001);
xnor U19743 (N_19743,N_15833,N_18063);
xor U19744 (N_19744,N_15680,N_17918);
xnor U19745 (N_19745,N_16150,N_17512);
nor U19746 (N_19746,N_18463,N_17668);
and U19747 (N_19747,N_18697,N_17642);
nand U19748 (N_19748,N_18346,N_16307);
or U19749 (N_19749,N_16448,N_16105);
or U19750 (N_19750,N_15718,N_18339);
or U19751 (N_19751,N_16837,N_17770);
or U19752 (N_19752,N_16353,N_18711);
or U19753 (N_19753,N_15993,N_16341);
nor U19754 (N_19754,N_16431,N_17303);
or U19755 (N_19755,N_17138,N_16179);
or U19756 (N_19756,N_15897,N_17738);
nor U19757 (N_19757,N_15770,N_17387);
nand U19758 (N_19758,N_15717,N_18494);
and U19759 (N_19759,N_17234,N_16808);
nor U19760 (N_19760,N_17875,N_17516);
and U19761 (N_19761,N_15818,N_16898);
nor U19762 (N_19762,N_17520,N_18622);
xor U19763 (N_19763,N_15920,N_18287);
xnor U19764 (N_19764,N_18181,N_16949);
and U19765 (N_19765,N_18081,N_15889);
nand U19766 (N_19766,N_15687,N_16946);
xor U19767 (N_19767,N_15676,N_15921);
nor U19768 (N_19768,N_15975,N_18483);
and U19769 (N_19769,N_16267,N_16851);
nor U19770 (N_19770,N_16861,N_17075);
nand U19771 (N_19771,N_18084,N_17663);
or U19772 (N_19772,N_17867,N_17090);
xnor U19773 (N_19773,N_17460,N_18092);
xnor U19774 (N_19774,N_17543,N_17129);
xnor U19775 (N_19775,N_17724,N_17832);
or U19776 (N_19776,N_16873,N_17132);
nor U19777 (N_19777,N_16042,N_15981);
and U19778 (N_19778,N_18221,N_18100);
nor U19779 (N_19779,N_16329,N_16309);
and U19780 (N_19780,N_17063,N_16255);
nor U19781 (N_19781,N_17590,N_16577);
nand U19782 (N_19782,N_15714,N_17229);
nor U19783 (N_19783,N_16380,N_16046);
nor U19784 (N_19784,N_15950,N_15982);
and U19785 (N_19785,N_18211,N_18611);
xnor U19786 (N_19786,N_17101,N_17417);
nor U19787 (N_19787,N_16533,N_16190);
nand U19788 (N_19788,N_17921,N_17210);
or U19789 (N_19789,N_16743,N_17620);
and U19790 (N_19790,N_17977,N_17499);
and U19791 (N_19791,N_17369,N_18687);
and U19792 (N_19792,N_18166,N_15956);
xnor U19793 (N_19793,N_17315,N_17248);
and U19794 (N_19794,N_18523,N_18700);
nor U19795 (N_19795,N_16073,N_16928);
nor U19796 (N_19796,N_17356,N_16090);
nor U19797 (N_19797,N_18726,N_17910);
xor U19798 (N_19798,N_18317,N_17393);
and U19799 (N_19799,N_16346,N_16695);
nor U19800 (N_19800,N_18383,N_18180);
xnor U19801 (N_19801,N_16905,N_18294);
and U19802 (N_19802,N_18577,N_18703);
xor U19803 (N_19803,N_16931,N_16867);
nand U19804 (N_19804,N_15823,N_16955);
and U19805 (N_19805,N_16728,N_17352);
nand U19806 (N_19806,N_18484,N_18691);
xor U19807 (N_19807,N_15778,N_16793);
or U19808 (N_19808,N_18163,N_15626);
nand U19809 (N_19809,N_17005,N_16014);
nand U19810 (N_19810,N_18659,N_17542);
nor U19811 (N_19811,N_17401,N_17797);
nand U19812 (N_19812,N_18192,N_17844);
and U19813 (N_19813,N_17111,N_17386);
nand U19814 (N_19814,N_18664,N_17056);
and U19815 (N_19815,N_17158,N_18086);
and U19816 (N_19816,N_15753,N_15974);
nor U19817 (N_19817,N_16582,N_17130);
xor U19818 (N_19818,N_17860,N_18098);
nand U19819 (N_19819,N_17760,N_17347);
nor U19820 (N_19820,N_15991,N_18408);
and U19821 (N_19821,N_17714,N_16211);
or U19822 (N_19822,N_16143,N_18461);
xnor U19823 (N_19823,N_16520,N_15797);
nor U19824 (N_19824,N_16543,N_15787);
and U19825 (N_19825,N_18150,N_17454);
nand U19826 (N_19826,N_16052,N_17641);
nand U19827 (N_19827,N_16750,N_18157);
or U19828 (N_19828,N_18734,N_17327);
xor U19829 (N_19829,N_15924,N_16023);
nand U19830 (N_19830,N_17611,N_17276);
or U19831 (N_19831,N_18625,N_18443);
nor U19832 (N_19832,N_16454,N_16418);
xnor U19833 (N_19833,N_16630,N_15890);
or U19834 (N_19834,N_16357,N_16043);
and U19835 (N_19835,N_17116,N_17697);
nor U19836 (N_19836,N_17818,N_17565);
nor U19837 (N_19837,N_17140,N_16178);
nand U19838 (N_19838,N_17199,N_18105);
and U19839 (N_19839,N_18531,N_17659);
and U19840 (N_19840,N_18733,N_18097);
xor U19841 (N_19841,N_17147,N_18019);
nand U19842 (N_19842,N_16515,N_15996);
nor U19843 (N_19843,N_17384,N_16654);
or U19844 (N_19844,N_15933,N_17131);
xnor U19845 (N_19845,N_16622,N_15759);
nor U19846 (N_19846,N_15852,N_16044);
nand U19847 (N_19847,N_16355,N_16407);
or U19848 (N_19848,N_17083,N_18325);
and U19849 (N_19849,N_17031,N_16365);
nor U19850 (N_19850,N_16969,N_18605);
xor U19851 (N_19851,N_16037,N_18066);
nor U19852 (N_19852,N_18350,N_16484);
nand U19853 (N_19853,N_18197,N_15966);
and U19854 (N_19854,N_18363,N_17230);
nand U19855 (N_19855,N_16650,N_18450);
xnor U19856 (N_19856,N_15766,N_17883);
nor U19857 (N_19857,N_17613,N_17624);
xor U19858 (N_19858,N_18015,N_18133);
nand U19859 (N_19859,N_18320,N_16839);
xnor U19860 (N_19860,N_15906,N_18570);
or U19861 (N_19861,N_16999,N_17145);
or U19862 (N_19862,N_17705,N_15870);
nand U19863 (N_19863,N_16462,N_15851);
and U19864 (N_19864,N_17560,N_16876);
and U19865 (N_19865,N_16635,N_17108);
or U19866 (N_19866,N_17984,N_16121);
and U19867 (N_19867,N_16646,N_18731);
and U19868 (N_19868,N_18636,N_16336);
xor U19869 (N_19869,N_16593,N_16993);
or U19870 (N_19870,N_18273,N_17039);
and U19871 (N_19871,N_18660,N_16367);
and U19872 (N_19872,N_17383,N_18745);
nor U19873 (N_19873,N_18497,N_17702);
or U19874 (N_19874,N_15745,N_15774);
nand U19875 (N_19875,N_17227,N_17740);
nand U19876 (N_19876,N_18038,N_17069);
nor U19877 (N_19877,N_18616,N_16149);
or U19878 (N_19878,N_17265,N_15671);
or U19879 (N_19879,N_18615,N_18487);
nand U19880 (N_19880,N_15665,N_16615);
nand U19881 (N_19881,N_16312,N_18727);
nor U19882 (N_19882,N_17139,N_16836);
nor U19883 (N_19883,N_16613,N_15983);
nand U19884 (N_19884,N_17133,N_18405);
and U19885 (N_19885,N_15679,N_16320);
and U19886 (N_19886,N_18653,N_18002);
and U19887 (N_19887,N_17113,N_15976);
nand U19888 (N_19888,N_18640,N_18036);
or U19889 (N_19889,N_15954,N_16292);
nor U19890 (N_19890,N_17686,N_18401);
or U19891 (N_19891,N_18029,N_16470);
and U19892 (N_19892,N_18152,N_15793);
nor U19893 (N_19893,N_18334,N_17734);
or U19894 (N_19894,N_16933,N_15729);
nor U19895 (N_19895,N_18114,N_17080);
xor U19896 (N_19896,N_16438,N_16257);
or U19897 (N_19897,N_16385,N_16159);
and U19898 (N_19898,N_16540,N_16537);
nand U19899 (N_19899,N_18255,N_16904);
xor U19900 (N_19900,N_18236,N_17170);
and U19901 (N_19901,N_17515,N_16772);
nand U19902 (N_19902,N_15896,N_15948);
xor U19903 (N_19903,N_16186,N_17077);
nand U19904 (N_19904,N_16809,N_16301);
or U19905 (N_19905,N_18353,N_17681);
xor U19906 (N_19906,N_16995,N_16551);
xor U19907 (N_19907,N_16843,N_15878);
or U19908 (N_19908,N_18324,N_17468);
and U19909 (N_19909,N_15713,N_16288);
and U19910 (N_19910,N_15895,N_16311);
nor U19911 (N_19911,N_16614,N_16671);
nor U19912 (N_19912,N_18247,N_16827);
xor U19913 (N_19913,N_16265,N_15995);
nor U19914 (N_19914,N_17378,N_17839);
and U19915 (N_19915,N_17829,N_18730);
and U19916 (N_19916,N_18169,N_17924);
xor U19917 (N_19917,N_18585,N_18638);
xor U19918 (N_19918,N_16167,N_16404);
or U19919 (N_19919,N_17109,N_16626);
and U19920 (N_19920,N_17269,N_16094);
xnor U19921 (N_19921,N_17420,N_17441);
or U19922 (N_19922,N_18115,N_17470);
and U19923 (N_19923,N_17901,N_18418);
xnor U19924 (N_19924,N_16612,N_17634);
nand U19925 (N_19925,N_17362,N_17943);
or U19926 (N_19926,N_15973,N_17214);
xor U19927 (N_19927,N_17023,N_17551);
xnor U19928 (N_19928,N_18296,N_16492);
xor U19929 (N_19929,N_16295,N_17256);
and U19930 (N_19930,N_17254,N_18244);
or U19931 (N_19931,N_15959,N_18108);
xor U19932 (N_19932,N_17010,N_16083);
nor U19933 (N_19933,N_15805,N_17349);
and U19934 (N_19934,N_16214,N_16799);
xor U19935 (N_19935,N_16807,N_17166);
nor U19936 (N_19936,N_17859,N_17614);
and U19937 (N_19937,N_17200,N_17897);
nor U19938 (N_19938,N_18671,N_17914);
or U19939 (N_19939,N_17775,N_16409);
xnor U19940 (N_19940,N_16561,N_18737);
nor U19941 (N_19941,N_17748,N_16603);
nand U19942 (N_19942,N_15944,N_17584);
or U19943 (N_19943,N_18455,N_17764);
nor U19944 (N_19944,N_16466,N_16707);
or U19945 (N_19945,N_18681,N_18121);
nor U19946 (N_19946,N_16565,N_17819);
or U19947 (N_19947,N_16432,N_18382);
nand U19948 (N_19948,N_16245,N_16379);
or U19949 (N_19949,N_16841,N_16601);
and U19950 (N_19950,N_18538,N_17476);
nor U19951 (N_19951,N_16701,N_15923);
xor U19952 (N_19952,N_17603,N_15918);
xnor U19953 (N_19953,N_17568,N_17664);
or U19954 (N_19954,N_17222,N_17669);
xor U19955 (N_19955,N_15936,N_16541);
or U19956 (N_19956,N_17986,N_18256);
nor U19957 (N_19957,N_17784,N_18385);
or U19958 (N_19958,N_18614,N_16262);
xor U19959 (N_19959,N_17650,N_15819);
xnor U19960 (N_19960,N_16600,N_18381);
xnor U19961 (N_19961,N_18416,N_17531);
or U19962 (N_19962,N_15701,N_17070);
nor U19963 (N_19963,N_18527,N_18054);
nand U19964 (N_19964,N_16942,N_15894);
xor U19965 (N_19965,N_17339,N_16754);
or U19966 (N_19966,N_16406,N_17314);
nor U19967 (N_19967,N_16400,N_16287);
nand U19968 (N_19968,N_18268,N_18014);
or U19969 (N_19969,N_17162,N_16620);
xnor U19970 (N_19970,N_18701,N_18676);
or U19971 (N_19971,N_15748,N_16111);
xor U19972 (N_19972,N_17766,N_16092);
nor U19973 (N_19973,N_18021,N_17237);
or U19974 (N_19974,N_17360,N_17524);
or U19975 (N_19975,N_15840,N_16057);
xor U19976 (N_19976,N_18196,N_16011);
xor U19977 (N_19977,N_17853,N_18013);
or U19978 (N_19978,N_16856,N_15660);
nor U19979 (N_19979,N_17555,N_17446);
and U19980 (N_19980,N_18704,N_16017);
and U19981 (N_19981,N_15841,N_15844);
xor U19982 (N_19982,N_15754,N_17758);
or U19983 (N_19983,N_17450,N_16345);
and U19984 (N_19984,N_16145,N_18074);
nor U19985 (N_19985,N_18387,N_17920);
nand U19986 (N_19986,N_17273,N_16705);
and U19987 (N_19987,N_16317,N_17987);
and U19988 (N_19988,N_17967,N_15872);
or U19989 (N_19989,N_16702,N_18200);
nand U19990 (N_19990,N_17922,N_15949);
and U19991 (N_19991,N_16256,N_16306);
or U19992 (N_19992,N_16476,N_17798);
xor U19993 (N_19993,N_17837,N_17877);
and U19994 (N_19994,N_16775,N_17579);
and U19995 (N_19995,N_18263,N_18312);
xnor U19996 (N_19996,N_18528,N_18469);
nor U19997 (N_19997,N_16778,N_15861);
and U19998 (N_19998,N_17510,N_16714);
nor U19999 (N_19999,N_16068,N_18237);
or U20000 (N_20000,N_17790,N_16125);
and U20001 (N_20001,N_16316,N_18662);
nor U20002 (N_20002,N_15710,N_17246);
nand U20003 (N_20003,N_15946,N_17361);
and U20004 (N_20004,N_17526,N_17497);
or U20005 (N_20005,N_18397,N_15868);
nor U20006 (N_20006,N_17504,N_17773);
or U20007 (N_20007,N_17495,N_16896);
and U20008 (N_20008,N_16828,N_16437);
nand U20009 (N_20009,N_17475,N_18649);
or U20010 (N_20010,N_18628,N_17209);
nor U20011 (N_20011,N_18050,N_15838);
or U20012 (N_20012,N_17646,N_17391);
and U20013 (N_20013,N_15858,N_16463);
nor U20014 (N_20014,N_16374,N_17794);
xor U20015 (N_20015,N_17280,N_17233);
nor U20016 (N_20016,N_17547,N_18059);
or U20017 (N_20017,N_17374,N_16891);
xnor U20018 (N_20018,N_18319,N_16487);
nand U20019 (N_20019,N_17654,N_17863);
and U20020 (N_20020,N_16247,N_18582);
or U20021 (N_20021,N_15876,N_16474);
xor U20022 (N_20022,N_16230,N_17678);
xnor U20023 (N_20023,N_15678,N_16983);
nor U20024 (N_20024,N_17995,N_16585);
xor U20025 (N_20025,N_16139,N_15696);
or U20026 (N_20026,N_17640,N_16321);
nor U20027 (N_20027,N_16927,N_17582);
and U20028 (N_20028,N_16020,N_17870);
nand U20029 (N_20029,N_15965,N_18742);
and U20030 (N_20030,N_16189,N_15666);
nand U20031 (N_20031,N_16191,N_18510);
nor U20032 (N_20032,N_17753,N_17082);
nor U20033 (N_20033,N_18149,N_17898);
nand U20034 (N_20034,N_18446,N_18323);
xnor U20035 (N_20035,N_18075,N_17201);
and U20036 (N_20036,N_17406,N_16674);
xnor U20037 (N_20037,N_17449,N_16528);
nor U20038 (N_20038,N_16361,N_15855);
nor U20039 (N_20039,N_15784,N_17826);
xor U20040 (N_20040,N_17159,N_18042);
and U20041 (N_20041,N_16670,N_18553);
nor U20042 (N_20042,N_18564,N_17486);
nor U20043 (N_20043,N_16621,N_16960);
nand U20044 (N_20044,N_15887,N_17301);
or U20045 (N_20045,N_17328,N_16405);
and U20046 (N_20046,N_16246,N_17258);
nand U20047 (N_20047,N_18655,N_15642);
or U20048 (N_20048,N_18336,N_18212);
or U20049 (N_20049,N_15842,N_15648);
and U20050 (N_20050,N_16819,N_17079);
xor U20051 (N_20051,N_16976,N_16932);
xor U20052 (N_20052,N_17022,N_17712);
nor U20053 (N_20053,N_18434,N_15829);
and U20054 (N_20054,N_17756,N_18347);
or U20055 (N_20055,N_17041,N_16286);
or U20056 (N_20056,N_18449,N_18457);
xor U20057 (N_20057,N_18583,N_18590);
nor U20058 (N_20058,N_16984,N_16591);
and U20059 (N_20059,N_15755,N_16326);
nor U20060 (N_20060,N_16805,N_16205);
or U20061 (N_20061,N_17969,N_18652);
xor U20062 (N_20062,N_15865,N_16844);
and U20063 (N_20063,N_18447,N_18473);
xnor U20064 (N_20064,N_15914,N_15716);
nand U20065 (N_20065,N_16411,N_17252);
nor U20066 (N_20066,N_15884,N_17881);
nand U20067 (N_20067,N_15649,N_16273);
and U20068 (N_20068,N_17673,N_17134);
and U20069 (N_20069,N_17437,N_18322);
xor U20070 (N_20070,N_16562,N_17182);
and U20071 (N_20071,N_17813,N_18119);
nor U20072 (N_20072,N_18508,N_16209);
and U20073 (N_20073,N_17029,N_16590);
nand U20074 (N_20074,N_17340,N_16099);
and U20075 (N_20075,N_17456,N_18199);
nor U20076 (N_20076,N_16829,N_17815);
or U20077 (N_20077,N_17711,N_16203);
nand U20078 (N_20078,N_18600,N_18429);
nand U20079 (N_20079,N_18400,N_17889);
nor U20080 (N_20080,N_18138,N_17189);
or U20081 (N_20081,N_18458,N_16518);
nand U20082 (N_20082,N_16064,N_15953);
xor U20083 (N_20083,N_15985,N_16410);
or U20084 (N_20084,N_15798,N_18391);
nand U20085 (N_20085,N_17581,N_17888);
xnor U20086 (N_20086,N_18165,N_18595);
and U20087 (N_20087,N_18039,N_16655);
and U20088 (N_20088,N_17341,N_18188);
nand U20089 (N_20089,N_16846,N_18716);
nand U20090 (N_20090,N_16147,N_17471);
xor U20091 (N_20091,N_15932,N_15697);
or U20092 (N_20092,N_16847,N_17629);
nor U20093 (N_20093,N_18501,N_17392);
xnor U20094 (N_20094,N_18025,N_18223);
nor U20095 (N_20095,N_16550,N_16523);
xor U20096 (N_20096,N_16231,N_16781);
or U20097 (N_20097,N_18297,N_16000);
or U20098 (N_20098,N_17906,N_17999);
or U20099 (N_20099,N_15725,N_18601);
or U20100 (N_20100,N_15875,N_16015);
or U20101 (N_20101,N_17344,N_17915);
nand U20102 (N_20102,N_17053,N_15744);
xnor U20103 (N_20103,N_16763,N_17065);
nand U20104 (N_20104,N_16132,N_18565);
or U20105 (N_20105,N_16430,N_16682);
or U20106 (N_20106,N_17733,N_18406);
xnor U20107 (N_20107,N_16796,N_17983);
nor U20108 (N_20108,N_15960,N_18707);
or U20109 (N_20109,N_18462,N_16327);
or U20110 (N_20110,N_16907,N_16238);
nand U20111 (N_20111,N_18009,N_16881);
nor U20112 (N_20112,N_15731,N_16944);
xor U20113 (N_20113,N_17970,N_16877);
or U20114 (N_20114,N_16414,N_18136);
xor U20115 (N_20115,N_18072,N_18644);
nand U20116 (N_20116,N_17974,N_16435);
or U20117 (N_20117,N_17638,N_15800);
nand U20118 (N_20118,N_15767,N_16795);
or U20119 (N_20119,N_16335,N_16009);
nor U20120 (N_20120,N_18436,N_16003);
xnor U20121 (N_20121,N_18540,N_16033);
nor U20122 (N_20122,N_17530,N_18384);
or U20123 (N_20123,N_15643,N_17806);
and U20124 (N_20124,N_16034,N_18402);
nand U20125 (N_20125,N_18016,N_15702);
nand U20126 (N_20126,N_18205,N_17701);
or U20127 (N_20127,N_18011,N_18490);
xor U20128 (N_20128,N_16974,N_18706);
xor U20129 (N_20129,N_17583,N_18056);
and U20130 (N_20130,N_17980,N_18282);
xnor U20131 (N_20131,N_15874,N_16096);
and U20132 (N_20132,N_17716,N_17573);
nor U20133 (N_20133,N_16388,N_16315);
or U20134 (N_20134,N_18316,N_17343);
or U20135 (N_20135,N_16332,N_18302);
xor U20136 (N_20136,N_18142,N_15834);
nand U20137 (N_20137,N_17191,N_16091);
nand U20138 (N_20138,N_16816,N_15782);
and U20139 (N_20139,N_16959,N_17876);
nand U20140 (N_20140,N_16990,N_18467);
nand U20141 (N_20141,N_17899,N_15908);
nand U20142 (N_20142,N_15707,N_18613);
nand U20143 (N_20143,N_17465,N_16556);
xor U20144 (N_20144,N_16784,N_16060);
or U20145 (N_20145,N_15938,N_17345);
nand U20146 (N_20146,N_15998,N_18459);
nor U20147 (N_20147,N_16548,N_16144);
xor U20148 (N_20148,N_17168,N_16833);
or U20149 (N_20149,N_16176,N_15625);
nand U20150 (N_20150,N_16554,N_16299);
nand U20151 (N_20151,N_17833,N_16331);
nand U20152 (N_20152,N_17768,N_18238);
xnor U20153 (N_20153,N_18137,N_17380);
or U20154 (N_20154,N_17439,N_16239);
xor U20155 (N_20155,N_16801,N_16098);
nand U20156 (N_20156,N_15638,N_15632);
or U20157 (N_20157,N_18248,N_17886);
nand U20158 (N_20158,N_16522,N_17208);
nand U20159 (N_20159,N_16539,N_17752);
xnor U20160 (N_20160,N_16252,N_18516);
xnor U20161 (N_20161,N_16088,N_17003);
nor U20162 (N_20162,N_17489,N_16604);
or U20163 (N_20163,N_15821,N_17221);
nor U20164 (N_20164,N_15929,N_16279);
or U20165 (N_20165,N_16656,N_17400);
or U20166 (N_20166,N_15822,N_18104);
nand U20167 (N_20167,N_17992,N_15864);
nand U20168 (N_20168,N_16115,N_16297);
nand U20169 (N_20169,N_17279,N_17183);
nor U20170 (N_20170,N_17030,N_18438);
nand U20171 (N_20171,N_15673,N_17236);
and U20172 (N_20172,N_17566,N_18219);
xor U20173 (N_20173,N_17779,N_18526);
and U20174 (N_20174,N_16322,N_18519);
nand U20175 (N_20175,N_17934,N_16444);
nand U20176 (N_20176,N_16025,N_18639);
nor U20177 (N_20177,N_17357,N_18452);
or U20178 (N_20178,N_17647,N_18702);
nor U20179 (N_20179,N_18040,N_17778);
or U20180 (N_20180,N_17366,N_18327);
or U20181 (N_20181,N_17319,N_16372);
and U20182 (N_20182,N_16250,N_17727);
or U20183 (N_20183,N_16451,N_18340);
and U20184 (N_20184,N_17235,N_16202);
and U20185 (N_20185,N_17978,N_16241);
and U20186 (N_20186,N_16578,N_16193);
xor U20187 (N_20187,N_17342,N_17706);
and U20188 (N_20188,N_16687,N_18130);
nand U20189 (N_20189,N_17639,N_16181);
nor U20190 (N_20190,N_17816,N_16785);
xnor U20191 (N_20191,N_17864,N_18656);
nand U20192 (N_20192,N_18718,N_17427);
nand U20193 (N_20193,N_17595,N_16510);
or U20194 (N_20194,N_17014,N_16610);
nand U20195 (N_20195,N_16629,N_16779);
and U20196 (N_20196,N_17321,N_15848);
and U20197 (N_20197,N_18569,N_15780);
xnor U20198 (N_20198,N_18099,N_16450);
nand U20199 (N_20199,N_16680,N_18135);
nand U20200 (N_20200,N_17322,N_16915);
or U20201 (N_20201,N_16164,N_15808);
nand U20202 (N_20202,N_17262,N_18475);
nor U20203 (N_20203,N_17428,N_16503);
nand U20204 (N_20204,N_17556,N_16632);
nand U20205 (N_20205,N_17019,N_18004);
or U20206 (N_20206,N_15968,N_18389);
xnor U20207 (N_20207,N_16866,N_16234);
or U20208 (N_20208,N_18456,N_17847);
nand U20209 (N_20209,N_16859,N_16659);
nor U20210 (N_20210,N_15750,N_18743);
xnor U20211 (N_20211,N_16100,N_17296);
xor U20212 (N_20212,N_18357,N_17513);
nand U20213 (N_20213,N_15799,N_16978);
xor U20214 (N_20214,N_18110,N_17173);
or U20215 (N_20215,N_17119,N_17691);
nor U20216 (N_20216,N_16126,N_17126);
and U20217 (N_20217,N_17912,N_18087);
and U20218 (N_20218,N_18355,N_18596);
nand U20219 (N_20219,N_18315,N_17334);
and U20220 (N_20220,N_17617,N_15633);
or U20221 (N_20221,N_17148,N_17828);
or U20222 (N_20222,N_17411,N_16103);
nor U20223 (N_20223,N_17432,N_16720);
nor U20224 (N_20224,N_16783,N_16545);
nand U20225 (N_20225,N_16679,N_16782);
and U20226 (N_20226,N_16264,N_17363);
nor U20227 (N_20227,N_18626,N_16820);
nand U20228 (N_20228,N_16127,N_16838);
xor U20229 (N_20229,N_18102,N_16885);
or U20230 (N_20230,N_17521,N_16443);
or U20231 (N_20231,N_17527,N_18177);
xor U20232 (N_20232,N_16572,N_18006);
and U20233 (N_20233,N_17094,N_16945);
or U20234 (N_20234,N_17903,N_16258);
xor U20235 (N_20235,N_16460,N_17574);
or U20236 (N_20236,N_18012,N_18496);
nand U20237 (N_20237,N_16858,N_18146);
xor U20238 (N_20238,N_17306,N_18252);
xnor U20239 (N_20239,N_17318,N_16228);
or U20240 (N_20240,N_16123,N_17267);
or U20241 (N_20241,N_17661,N_15794);
nand U20242 (N_20242,N_17151,N_18630);
or U20243 (N_20243,N_17804,N_18022);
nor U20244 (N_20244,N_16567,N_17414);
and U20245 (N_20245,N_17047,N_17192);
nand U20246 (N_20246,N_16131,N_16899);
or U20247 (N_20247,N_16053,N_15668);
xnor U20248 (N_20248,N_16441,N_16478);
or U20249 (N_20249,N_17684,N_16089);
nor U20250 (N_20250,N_17762,N_16047);
or U20251 (N_20251,N_16419,N_18298);
xnor U20252 (N_20252,N_16226,N_15644);
nor U20253 (N_20253,N_17589,N_17592);
nand U20254 (N_20254,N_18101,N_18344);
nor U20255 (N_20255,N_17068,N_17310);
xor U20256 (N_20256,N_18005,N_17219);
and U20257 (N_20257,N_18289,N_16700);
or U20258 (N_20258,N_18725,N_18482);
nand U20259 (N_20259,N_15812,N_17107);
or U20260 (N_20260,N_15786,N_16251);
nand U20261 (N_20261,N_17371,N_17463);
and U20262 (N_20262,N_18532,N_17905);
nor U20263 (N_20263,N_15674,N_15859);
xnor U20264 (N_20264,N_16002,N_17451);
and U20265 (N_20265,N_17025,N_18380);
nor U20266 (N_20266,N_17268,N_15703);
or U20267 (N_20267,N_16977,N_18178);
nor U20268 (N_20268,N_16180,N_17415);
or U20269 (N_20269,N_17577,N_17946);
or U20270 (N_20270,N_16440,N_17707);
nor U20271 (N_20271,N_16597,N_18428);
xor U20272 (N_20272,N_16909,N_16304);
or U20273 (N_20273,N_16358,N_15708);
and U20274 (N_20274,N_17874,N_16383);
xor U20275 (N_20275,N_17017,N_17472);
and U20276 (N_20276,N_18358,N_17184);
and U20277 (N_20277,N_18619,N_18096);
or U20278 (N_20278,N_16093,N_18422);
nor U20279 (N_20279,N_16161,N_17553);
and U20280 (N_20280,N_16305,N_16506);
xnor U20281 (N_20281,N_17286,N_16741);
and U20282 (N_20282,N_16634,N_15683);
xnor U20283 (N_20283,N_16731,N_18603);
nor U20284 (N_20284,N_15752,N_17698);
xor U20285 (N_20285,N_16559,N_17084);
and U20286 (N_20286,N_17115,N_16362);
or U20287 (N_20287,N_17628,N_16706);
nand U20288 (N_20288,N_17032,N_16490);
nand U20289 (N_20289,N_16200,N_16735);
or U20290 (N_20290,N_17588,N_17385);
nand U20291 (N_20291,N_16869,N_17324);
and U20292 (N_20292,N_18123,N_17501);
or U20293 (N_20293,N_18410,N_18388);
and U20294 (N_20294,N_15700,N_15853);
xnor U20295 (N_20295,N_17407,N_18275);
and U20296 (N_20296,N_16390,N_18425);
nand U20297 (N_20297,N_18412,N_16734);
xnor U20298 (N_20298,N_17351,N_16108);
or U20299 (N_20299,N_17893,N_15827);
or U20300 (N_20300,N_16736,N_16395);
or U20301 (N_20301,N_16146,N_15943);
nand U20302 (N_20302,N_15917,N_18053);
xnor U20303 (N_20303,N_17095,N_17630);
or U20304 (N_20304,N_17549,N_16010);
xor U20305 (N_20305,N_16294,N_16673);
nor U20306 (N_20306,N_17043,N_17576);
nand U20307 (N_20307,N_17114,N_16568);
nor U20308 (N_20308,N_16427,N_16926);
or U20309 (N_20309,N_17739,N_16022);
and U20310 (N_20310,N_18321,N_16495);
and U20311 (N_20311,N_18587,N_18415);
or U20312 (N_20312,N_17185,N_16823);
and U20313 (N_20313,N_15824,N_16893);
or U20314 (N_20314,N_16613,N_16061);
nand U20315 (N_20315,N_16049,N_17033);
nand U20316 (N_20316,N_18583,N_16490);
and U20317 (N_20317,N_17457,N_17352);
xor U20318 (N_20318,N_17838,N_18406);
nor U20319 (N_20319,N_18673,N_15697);
xnor U20320 (N_20320,N_18262,N_16343);
or U20321 (N_20321,N_17084,N_15974);
and U20322 (N_20322,N_18062,N_18354);
xnor U20323 (N_20323,N_17825,N_18644);
xor U20324 (N_20324,N_18006,N_15882);
and U20325 (N_20325,N_17570,N_17765);
and U20326 (N_20326,N_16901,N_17271);
nand U20327 (N_20327,N_17263,N_16726);
xnor U20328 (N_20328,N_17838,N_17835);
and U20329 (N_20329,N_17216,N_18614);
xor U20330 (N_20330,N_17942,N_17286);
nand U20331 (N_20331,N_17470,N_16266);
xnor U20332 (N_20332,N_16284,N_16018);
xnor U20333 (N_20333,N_16161,N_17098);
and U20334 (N_20334,N_17864,N_16824);
nand U20335 (N_20335,N_16620,N_18244);
xor U20336 (N_20336,N_16095,N_15663);
nand U20337 (N_20337,N_16668,N_17339);
nand U20338 (N_20338,N_18527,N_18183);
and U20339 (N_20339,N_16671,N_17949);
nor U20340 (N_20340,N_17246,N_15699);
or U20341 (N_20341,N_17458,N_18575);
and U20342 (N_20342,N_17042,N_17576);
and U20343 (N_20343,N_18194,N_17871);
xor U20344 (N_20344,N_16668,N_17059);
nor U20345 (N_20345,N_16192,N_17614);
and U20346 (N_20346,N_17131,N_16180);
nor U20347 (N_20347,N_17026,N_17851);
nor U20348 (N_20348,N_18461,N_18638);
or U20349 (N_20349,N_17619,N_15818);
and U20350 (N_20350,N_17427,N_18081);
nor U20351 (N_20351,N_18731,N_16540);
nor U20352 (N_20352,N_15952,N_18625);
and U20353 (N_20353,N_18098,N_16146);
xnor U20354 (N_20354,N_17565,N_17118);
nand U20355 (N_20355,N_17539,N_17253);
nand U20356 (N_20356,N_15962,N_18150);
and U20357 (N_20357,N_18306,N_17676);
and U20358 (N_20358,N_17766,N_17213);
and U20359 (N_20359,N_18033,N_18309);
and U20360 (N_20360,N_17049,N_18657);
or U20361 (N_20361,N_16053,N_15645);
or U20362 (N_20362,N_16815,N_16510);
and U20363 (N_20363,N_17198,N_16891);
or U20364 (N_20364,N_18012,N_18255);
and U20365 (N_20365,N_16415,N_15814);
or U20366 (N_20366,N_16193,N_15664);
or U20367 (N_20367,N_16289,N_16933);
nor U20368 (N_20368,N_18027,N_17459);
and U20369 (N_20369,N_16363,N_17443);
nand U20370 (N_20370,N_16005,N_18745);
and U20371 (N_20371,N_18007,N_18363);
xnor U20372 (N_20372,N_18048,N_15945);
and U20373 (N_20373,N_16265,N_17495);
nor U20374 (N_20374,N_16417,N_17545);
nand U20375 (N_20375,N_18629,N_16215);
nor U20376 (N_20376,N_17366,N_17310);
or U20377 (N_20377,N_16195,N_15710);
nor U20378 (N_20378,N_18078,N_18146);
nor U20379 (N_20379,N_17173,N_18079);
nand U20380 (N_20380,N_16271,N_17328);
and U20381 (N_20381,N_18565,N_17019);
xnor U20382 (N_20382,N_16407,N_18121);
nand U20383 (N_20383,N_15763,N_18156);
xnor U20384 (N_20384,N_17668,N_16739);
and U20385 (N_20385,N_17676,N_17818);
xor U20386 (N_20386,N_17566,N_18021);
or U20387 (N_20387,N_18245,N_17026);
and U20388 (N_20388,N_15806,N_16138);
nor U20389 (N_20389,N_18632,N_17596);
xnor U20390 (N_20390,N_17465,N_16514);
nand U20391 (N_20391,N_16072,N_16014);
nor U20392 (N_20392,N_18688,N_16151);
and U20393 (N_20393,N_16696,N_18383);
and U20394 (N_20394,N_16553,N_18059);
xnor U20395 (N_20395,N_18204,N_16793);
nand U20396 (N_20396,N_16448,N_18588);
nand U20397 (N_20397,N_18370,N_17632);
or U20398 (N_20398,N_18486,N_18187);
or U20399 (N_20399,N_17723,N_15685);
nor U20400 (N_20400,N_16916,N_18492);
and U20401 (N_20401,N_15763,N_16908);
nand U20402 (N_20402,N_18644,N_15952);
xnor U20403 (N_20403,N_17068,N_16259);
or U20404 (N_20404,N_18588,N_18066);
xor U20405 (N_20405,N_16268,N_16869);
xor U20406 (N_20406,N_18658,N_16585);
and U20407 (N_20407,N_18170,N_18490);
nor U20408 (N_20408,N_17816,N_18161);
and U20409 (N_20409,N_18383,N_18081);
nor U20410 (N_20410,N_17381,N_17320);
nor U20411 (N_20411,N_17298,N_18313);
nor U20412 (N_20412,N_17020,N_15673);
or U20413 (N_20413,N_18248,N_18240);
xnor U20414 (N_20414,N_16092,N_17658);
or U20415 (N_20415,N_18142,N_15818);
nand U20416 (N_20416,N_16891,N_18637);
and U20417 (N_20417,N_16422,N_17057);
xor U20418 (N_20418,N_16677,N_16744);
nor U20419 (N_20419,N_16075,N_17592);
nor U20420 (N_20420,N_18556,N_17846);
nand U20421 (N_20421,N_18560,N_18181);
or U20422 (N_20422,N_16398,N_17874);
and U20423 (N_20423,N_16848,N_16816);
nor U20424 (N_20424,N_17375,N_16138);
xnor U20425 (N_20425,N_17414,N_18558);
and U20426 (N_20426,N_16063,N_17430);
xor U20427 (N_20427,N_18608,N_17962);
nand U20428 (N_20428,N_15745,N_17276);
or U20429 (N_20429,N_16267,N_17165);
xor U20430 (N_20430,N_18495,N_17227);
or U20431 (N_20431,N_17272,N_15959);
xnor U20432 (N_20432,N_15849,N_15939);
or U20433 (N_20433,N_16048,N_17178);
or U20434 (N_20434,N_16322,N_18113);
and U20435 (N_20435,N_16913,N_18062);
or U20436 (N_20436,N_17745,N_17458);
nand U20437 (N_20437,N_18116,N_16194);
and U20438 (N_20438,N_16402,N_18713);
or U20439 (N_20439,N_18090,N_18652);
or U20440 (N_20440,N_17510,N_17170);
or U20441 (N_20441,N_17983,N_15801);
or U20442 (N_20442,N_17298,N_17939);
nor U20443 (N_20443,N_17535,N_16380);
nand U20444 (N_20444,N_18075,N_18237);
xnor U20445 (N_20445,N_18540,N_18067);
nor U20446 (N_20446,N_16211,N_17407);
xnor U20447 (N_20447,N_16013,N_17014);
nand U20448 (N_20448,N_18348,N_18026);
and U20449 (N_20449,N_17367,N_16100);
xnor U20450 (N_20450,N_17749,N_18293);
or U20451 (N_20451,N_18026,N_18519);
or U20452 (N_20452,N_15771,N_18233);
xnor U20453 (N_20453,N_16121,N_16270);
nor U20454 (N_20454,N_18020,N_15661);
xnor U20455 (N_20455,N_16799,N_15829);
or U20456 (N_20456,N_18608,N_17947);
xnor U20457 (N_20457,N_17614,N_17791);
and U20458 (N_20458,N_16171,N_16449);
nor U20459 (N_20459,N_17468,N_17172);
xor U20460 (N_20460,N_16414,N_18174);
nand U20461 (N_20461,N_16508,N_16646);
and U20462 (N_20462,N_18605,N_18746);
nand U20463 (N_20463,N_16236,N_18722);
nand U20464 (N_20464,N_16363,N_16389);
xor U20465 (N_20465,N_18560,N_16187);
nand U20466 (N_20466,N_15702,N_17031);
or U20467 (N_20467,N_17020,N_18154);
nor U20468 (N_20468,N_16513,N_17144);
and U20469 (N_20469,N_17895,N_15854);
or U20470 (N_20470,N_15852,N_17819);
nor U20471 (N_20471,N_17075,N_16040);
or U20472 (N_20472,N_17709,N_16684);
xnor U20473 (N_20473,N_18357,N_18499);
nand U20474 (N_20474,N_17614,N_17900);
or U20475 (N_20475,N_17069,N_15979);
nor U20476 (N_20476,N_16831,N_16826);
xor U20477 (N_20477,N_17686,N_18195);
and U20478 (N_20478,N_16903,N_18375);
nand U20479 (N_20479,N_17294,N_16503);
and U20480 (N_20480,N_16091,N_15994);
nand U20481 (N_20481,N_16407,N_16206);
nor U20482 (N_20482,N_17748,N_18353);
nor U20483 (N_20483,N_18182,N_18685);
nand U20484 (N_20484,N_17268,N_16079);
nand U20485 (N_20485,N_16430,N_15907);
nand U20486 (N_20486,N_17672,N_16667);
xor U20487 (N_20487,N_16171,N_18194);
xor U20488 (N_20488,N_17695,N_16109);
or U20489 (N_20489,N_17187,N_18689);
nand U20490 (N_20490,N_18657,N_16959);
or U20491 (N_20491,N_16887,N_18558);
nand U20492 (N_20492,N_18229,N_16020);
nand U20493 (N_20493,N_16045,N_18269);
or U20494 (N_20494,N_16388,N_16953);
xnor U20495 (N_20495,N_18246,N_18053);
or U20496 (N_20496,N_18385,N_17460);
and U20497 (N_20497,N_17576,N_18703);
xnor U20498 (N_20498,N_16767,N_17945);
nand U20499 (N_20499,N_16426,N_16288);
nand U20500 (N_20500,N_15953,N_15795);
and U20501 (N_20501,N_17919,N_16369);
and U20502 (N_20502,N_15978,N_18445);
and U20503 (N_20503,N_16044,N_16917);
or U20504 (N_20504,N_17071,N_16010);
and U20505 (N_20505,N_17089,N_17721);
xor U20506 (N_20506,N_18145,N_17430);
nand U20507 (N_20507,N_15896,N_18740);
xor U20508 (N_20508,N_15831,N_17985);
and U20509 (N_20509,N_16466,N_18399);
and U20510 (N_20510,N_16189,N_15716);
or U20511 (N_20511,N_16853,N_18112);
xor U20512 (N_20512,N_18727,N_16680);
or U20513 (N_20513,N_17769,N_16753);
xnor U20514 (N_20514,N_18709,N_17162);
or U20515 (N_20515,N_18453,N_17801);
or U20516 (N_20516,N_17755,N_15688);
and U20517 (N_20517,N_16274,N_17754);
or U20518 (N_20518,N_18117,N_18430);
or U20519 (N_20519,N_15879,N_16268);
or U20520 (N_20520,N_16563,N_18136);
or U20521 (N_20521,N_18493,N_16059);
nor U20522 (N_20522,N_17315,N_15747);
xor U20523 (N_20523,N_18631,N_17030);
or U20524 (N_20524,N_18131,N_16747);
nand U20525 (N_20525,N_15790,N_16831);
nand U20526 (N_20526,N_18604,N_17295);
or U20527 (N_20527,N_15956,N_15874);
xnor U20528 (N_20528,N_17257,N_15695);
xor U20529 (N_20529,N_17970,N_17128);
or U20530 (N_20530,N_18244,N_18057);
xnor U20531 (N_20531,N_17112,N_17753);
xnor U20532 (N_20532,N_16816,N_15950);
xnor U20533 (N_20533,N_16926,N_17477);
xor U20534 (N_20534,N_15998,N_18239);
nor U20535 (N_20535,N_17982,N_16879);
xnor U20536 (N_20536,N_16688,N_16896);
and U20537 (N_20537,N_18489,N_18633);
and U20538 (N_20538,N_17169,N_18365);
xnor U20539 (N_20539,N_16344,N_16626);
xnor U20540 (N_20540,N_17457,N_16882);
nor U20541 (N_20541,N_16524,N_17477);
xnor U20542 (N_20542,N_17224,N_16288);
nand U20543 (N_20543,N_18669,N_18121);
xor U20544 (N_20544,N_18548,N_18679);
xnor U20545 (N_20545,N_17978,N_17003);
nand U20546 (N_20546,N_18027,N_18510);
nor U20547 (N_20547,N_16872,N_18081);
nand U20548 (N_20548,N_18112,N_15848);
nor U20549 (N_20549,N_17856,N_16761);
nor U20550 (N_20550,N_16413,N_16840);
and U20551 (N_20551,N_18026,N_16247);
and U20552 (N_20552,N_17260,N_15998);
and U20553 (N_20553,N_18595,N_16278);
nand U20554 (N_20554,N_16582,N_16739);
and U20555 (N_20555,N_18666,N_17547);
nor U20556 (N_20556,N_15768,N_15707);
or U20557 (N_20557,N_16022,N_17302);
or U20558 (N_20558,N_16463,N_17070);
nand U20559 (N_20559,N_18161,N_18424);
nand U20560 (N_20560,N_17374,N_17417);
xor U20561 (N_20561,N_16388,N_15825);
nor U20562 (N_20562,N_16401,N_15751);
nor U20563 (N_20563,N_18378,N_16105);
nand U20564 (N_20564,N_16392,N_16066);
and U20565 (N_20565,N_18314,N_15917);
or U20566 (N_20566,N_18159,N_17812);
xor U20567 (N_20567,N_16494,N_17171);
nor U20568 (N_20568,N_17673,N_16586);
and U20569 (N_20569,N_16950,N_17532);
nand U20570 (N_20570,N_17631,N_18296);
nand U20571 (N_20571,N_17228,N_16778);
xnor U20572 (N_20572,N_18619,N_17120);
and U20573 (N_20573,N_18174,N_16887);
or U20574 (N_20574,N_15831,N_18721);
nand U20575 (N_20575,N_16200,N_15976);
and U20576 (N_20576,N_16228,N_17840);
nor U20577 (N_20577,N_16178,N_16250);
nand U20578 (N_20578,N_18425,N_17157);
xnor U20579 (N_20579,N_18574,N_16799);
or U20580 (N_20580,N_15662,N_16790);
xnor U20581 (N_20581,N_18616,N_18462);
xor U20582 (N_20582,N_17592,N_17631);
nor U20583 (N_20583,N_17780,N_15945);
xnor U20584 (N_20584,N_15954,N_17220);
and U20585 (N_20585,N_18663,N_16414);
or U20586 (N_20586,N_17168,N_16931);
nor U20587 (N_20587,N_15893,N_17912);
or U20588 (N_20588,N_15698,N_16320);
xor U20589 (N_20589,N_17258,N_17934);
nand U20590 (N_20590,N_18495,N_16040);
and U20591 (N_20591,N_18125,N_16239);
nand U20592 (N_20592,N_16442,N_18351);
nor U20593 (N_20593,N_17401,N_16251);
or U20594 (N_20594,N_18060,N_18702);
and U20595 (N_20595,N_16465,N_17341);
nor U20596 (N_20596,N_17543,N_17128);
or U20597 (N_20597,N_16615,N_18549);
xnor U20598 (N_20598,N_18059,N_16998);
nor U20599 (N_20599,N_15687,N_16409);
nor U20600 (N_20600,N_16492,N_18621);
nand U20601 (N_20601,N_17830,N_18446);
xnor U20602 (N_20602,N_18146,N_18618);
nor U20603 (N_20603,N_16769,N_18231);
and U20604 (N_20604,N_17550,N_16422);
nor U20605 (N_20605,N_18608,N_16069);
nand U20606 (N_20606,N_17818,N_18385);
xor U20607 (N_20607,N_16680,N_17367);
or U20608 (N_20608,N_16781,N_18310);
nor U20609 (N_20609,N_15797,N_16130);
xor U20610 (N_20610,N_16465,N_17881);
and U20611 (N_20611,N_17999,N_16231);
nand U20612 (N_20612,N_17303,N_16561);
nand U20613 (N_20613,N_17562,N_17886);
or U20614 (N_20614,N_16638,N_16556);
nand U20615 (N_20615,N_16930,N_18449);
xnor U20616 (N_20616,N_17947,N_18012);
nor U20617 (N_20617,N_16027,N_18709);
nand U20618 (N_20618,N_17448,N_15986);
or U20619 (N_20619,N_16242,N_16934);
nand U20620 (N_20620,N_16298,N_17984);
or U20621 (N_20621,N_17288,N_17760);
xor U20622 (N_20622,N_17321,N_16151);
xor U20623 (N_20623,N_15864,N_18141);
and U20624 (N_20624,N_17624,N_16879);
xor U20625 (N_20625,N_18452,N_18272);
xor U20626 (N_20626,N_17874,N_18262);
nand U20627 (N_20627,N_15968,N_16127);
and U20628 (N_20628,N_17010,N_18258);
or U20629 (N_20629,N_18745,N_18540);
xnor U20630 (N_20630,N_17922,N_18330);
xor U20631 (N_20631,N_16712,N_15866);
nor U20632 (N_20632,N_18125,N_16898);
nand U20633 (N_20633,N_18713,N_16388);
xor U20634 (N_20634,N_15882,N_16215);
and U20635 (N_20635,N_16298,N_17770);
xnor U20636 (N_20636,N_18661,N_16573);
nor U20637 (N_20637,N_18497,N_15676);
and U20638 (N_20638,N_17179,N_18458);
and U20639 (N_20639,N_18412,N_15787);
nor U20640 (N_20640,N_17908,N_17186);
xnor U20641 (N_20641,N_17847,N_18434);
nand U20642 (N_20642,N_18007,N_16379);
xor U20643 (N_20643,N_18325,N_17359);
nor U20644 (N_20644,N_18133,N_18626);
or U20645 (N_20645,N_15805,N_17987);
and U20646 (N_20646,N_16182,N_17481);
xnor U20647 (N_20647,N_18522,N_17646);
nor U20648 (N_20648,N_17884,N_17771);
nor U20649 (N_20649,N_18327,N_18408);
or U20650 (N_20650,N_18108,N_17661);
or U20651 (N_20651,N_17309,N_18638);
xor U20652 (N_20652,N_18051,N_18053);
nor U20653 (N_20653,N_18550,N_16022);
or U20654 (N_20654,N_15941,N_16266);
nand U20655 (N_20655,N_16051,N_15721);
nor U20656 (N_20656,N_17830,N_17368);
nand U20657 (N_20657,N_18001,N_18162);
nand U20658 (N_20658,N_15844,N_18361);
xnor U20659 (N_20659,N_17476,N_18587);
and U20660 (N_20660,N_17082,N_16090);
xor U20661 (N_20661,N_16698,N_18433);
or U20662 (N_20662,N_18251,N_16800);
and U20663 (N_20663,N_17062,N_16398);
and U20664 (N_20664,N_16854,N_18721);
nor U20665 (N_20665,N_15843,N_18604);
xor U20666 (N_20666,N_16757,N_17522);
or U20667 (N_20667,N_17891,N_18574);
or U20668 (N_20668,N_18736,N_17278);
or U20669 (N_20669,N_15849,N_15671);
and U20670 (N_20670,N_17988,N_16312);
xor U20671 (N_20671,N_16080,N_17192);
nand U20672 (N_20672,N_15803,N_18325);
nor U20673 (N_20673,N_15659,N_16765);
xor U20674 (N_20674,N_18519,N_17683);
xor U20675 (N_20675,N_17648,N_16233);
or U20676 (N_20676,N_17130,N_18352);
or U20677 (N_20677,N_16489,N_16810);
nand U20678 (N_20678,N_17858,N_18530);
nand U20679 (N_20679,N_16164,N_16938);
nand U20680 (N_20680,N_16700,N_17651);
xnor U20681 (N_20681,N_17914,N_16610);
or U20682 (N_20682,N_17820,N_17210);
nor U20683 (N_20683,N_18549,N_17457);
nand U20684 (N_20684,N_16789,N_16195);
xor U20685 (N_20685,N_17792,N_16248);
or U20686 (N_20686,N_17395,N_16277);
nand U20687 (N_20687,N_16002,N_17082);
and U20688 (N_20688,N_16775,N_18268);
nand U20689 (N_20689,N_15733,N_16647);
or U20690 (N_20690,N_15720,N_18733);
or U20691 (N_20691,N_16799,N_15774);
xor U20692 (N_20692,N_17712,N_15874);
nor U20693 (N_20693,N_18731,N_16788);
nand U20694 (N_20694,N_18117,N_18507);
xor U20695 (N_20695,N_15960,N_17565);
nand U20696 (N_20696,N_16039,N_17148);
nor U20697 (N_20697,N_18473,N_17901);
nor U20698 (N_20698,N_18734,N_16936);
xnor U20699 (N_20699,N_15941,N_16430);
or U20700 (N_20700,N_16904,N_17433);
or U20701 (N_20701,N_17094,N_15828);
and U20702 (N_20702,N_17131,N_17933);
or U20703 (N_20703,N_16977,N_18697);
and U20704 (N_20704,N_18094,N_17003);
or U20705 (N_20705,N_16690,N_16095);
nand U20706 (N_20706,N_18212,N_15876);
or U20707 (N_20707,N_17203,N_17101);
and U20708 (N_20708,N_17792,N_17394);
or U20709 (N_20709,N_18429,N_18099);
and U20710 (N_20710,N_16365,N_16130);
and U20711 (N_20711,N_16469,N_18676);
nand U20712 (N_20712,N_18457,N_16667);
nor U20713 (N_20713,N_17557,N_15913);
nand U20714 (N_20714,N_18743,N_15968);
nand U20715 (N_20715,N_17959,N_16510);
xnor U20716 (N_20716,N_16818,N_16406);
or U20717 (N_20717,N_17463,N_17633);
and U20718 (N_20718,N_16685,N_17633);
xnor U20719 (N_20719,N_17734,N_15661);
nor U20720 (N_20720,N_17041,N_16107);
nand U20721 (N_20721,N_18208,N_16114);
nor U20722 (N_20722,N_18119,N_16896);
and U20723 (N_20723,N_16871,N_18542);
nand U20724 (N_20724,N_16155,N_16097);
and U20725 (N_20725,N_16083,N_18650);
nand U20726 (N_20726,N_18456,N_15799);
or U20727 (N_20727,N_16090,N_16911);
nor U20728 (N_20728,N_18283,N_18173);
nand U20729 (N_20729,N_16251,N_15794);
nand U20730 (N_20730,N_17390,N_16670);
and U20731 (N_20731,N_17121,N_18660);
and U20732 (N_20732,N_16584,N_16412);
nor U20733 (N_20733,N_17608,N_17473);
nor U20734 (N_20734,N_15689,N_18685);
xor U20735 (N_20735,N_16256,N_18052);
or U20736 (N_20736,N_16118,N_17716);
nor U20737 (N_20737,N_17395,N_18486);
and U20738 (N_20738,N_16611,N_18347);
nand U20739 (N_20739,N_16311,N_16969);
or U20740 (N_20740,N_16696,N_16169);
and U20741 (N_20741,N_16921,N_17029);
nand U20742 (N_20742,N_18706,N_18598);
xor U20743 (N_20743,N_15817,N_17733);
xnor U20744 (N_20744,N_17832,N_18113);
nor U20745 (N_20745,N_17061,N_16456);
or U20746 (N_20746,N_17694,N_18380);
nor U20747 (N_20747,N_16060,N_16017);
nand U20748 (N_20748,N_15847,N_18113);
nand U20749 (N_20749,N_18469,N_17698);
xnor U20750 (N_20750,N_17973,N_16039);
nor U20751 (N_20751,N_16885,N_18586);
nor U20752 (N_20752,N_17853,N_18094);
or U20753 (N_20753,N_16444,N_18199);
xor U20754 (N_20754,N_18034,N_15935);
or U20755 (N_20755,N_18435,N_17677);
or U20756 (N_20756,N_15972,N_17690);
and U20757 (N_20757,N_17582,N_17060);
nand U20758 (N_20758,N_17531,N_15689);
nand U20759 (N_20759,N_18688,N_16294);
xnor U20760 (N_20760,N_15995,N_18172);
and U20761 (N_20761,N_17200,N_16695);
or U20762 (N_20762,N_16231,N_16232);
nand U20763 (N_20763,N_18648,N_16070);
and U20764 (N_20764,N_17130,N_16305);
xnor U20765 (N_20765,N_16484,N_18699);
nor U20766 (N_20766,N_17766,N_16245);
nor U20767 (N_20767,N_18321,N_17605);
nand U20768 (N_20768,N_18338,N_18400);
and U20769 (N_20769,N_16984,N_16987);
or U20770 (N_20770,N_16997,N_16823);
nor U20771 (N_20771,N_17221,N_17700);
or U20772 (N_20772,N_17784,N_17102);
and U20773 (N_20773,N_15772,N_17813);
or U20774 (N_20774,N_17249,N_16652);
nand U20775 (N_20775,N_17216,N_15998);
xor U20776 (N_20776,N_16461,N_17093);
xor U20777 (N_20777,N_16835,N_16089);
nor U20778 (N_20778,N_17062,N_18685);
xor U20779 (N_20779,N_17589,N_16643);
nor U20780 (N_20780,N_16503,N_16906);
nand U20781 (N_20781,N_18028,N_18247);
nor U20782 (N_20782,N_16981,N_16770);
xor U20783 (N_20783,N_16510,N_16117);
and U20784 (N_20784,N_17484,N_17666);
or U20785 (N_20785,N_16504,N_17819);
nor U20786 (N_20786,N_17849,N_17016);
nand U20787 (N_20787,N_15714,N_16424);
nand U20788 (N_20788,N_16307,N_18128);
nand U20789 (N_20789,N_17173,N_16714);
nand U20790 (N_20790,N_16822,N_17146);
or U20791 (N_20791,N_16125,N_18527);
and U20792 (N_20792,N_16912,N_18593);
xor U20793 (N_20793,N_18074,N_17552);
xor U20794 (N_20794,N_15930,N_18307);
xor U20795 (N_20795,N_17049,N_16823);
nor U20796 (N_20796,N_16227,N_17607);
nor U20797 (N_20797,N_16227,N_17725);
or U20798 (N_20798,N_15649,N_18514);
nand U20799 (N_20799,N_17815,N_18238);
and U20800 (N_20800,N_17944,N_17251);
nand U20801 (N_20801,N_16234,N_18369);
and U20802 (N_20802,N_16538,N_17909);
and U20803 (N_20803,N_16941,N_17386);
or U20804 (N_20804,N_16624,N_17052);
nor U20805 (N_20805,N_15706,N_18034);
nor U20806 (N_20806,N_16797,N_17816);
nor U20807 (N_20807,N_17830,N_17182);
and U20808 (N_20808,N_18668,N_15908);
and U20809 (N_20809,N_17326,N_15851);
and U20810 (N_20810,N_16571,N_18624);
xnor U20811 (N_20811,N_16913,N_16958);
and U20812 (N_20812,N_17743,N_16816);
and U20813 (N_20813,N_18401,N_16077);
and U20814 (N_20814,N_17821,N_18616);
nand U20815 (N_20815,N_16213,N_16449);
nand U20816 (N_20816,N_16958,N_18280);
nand U20817 (N_20817,N_18278,N_16844);
xnor U20818 (N_20818,N_16091,N_15847);
or U20819 (N_20819,N_15879,N_16719);
nand U20820 (N_20820,N_15937,N_16280);
or U20821 (N_20821,N_18191,N_17098);
nor U20822 (N_20822,N_16970,N_17571);
or U20823 (N_20823,N_16060,N_18154);
and U20824 (N_20824,N_17804,N_17596);
or U20825 (N_20825,N_17546,N_16656);
and U20826 (N_20826,N_17008,N_16884);
nand U20827 (N_20827,N_16128,N_16586);
nor U20828 (N_20828,N_16604,N_18127);
and U20829 (N_20829,N_17172,N_17259);
nand U20830 (N_20830,N_16204,N_18373);
xor U20831 (N_20831,N_17713,N_16810);
and U20832 (N_20832,N_17957,N_16373);
and U20833 (N_20833,N_15795,N_16201);
and U20834 (N_20834,N_18428,N_17487);
xor U20835 (N_20835,N_18444,N_16434);
nand U20836 (N_20836,N_16395,N_15652);
and U20837 (N_20837,N_16339,N_18313);
and U20838 (N_20838,N_17457,N_18460);
and U20839 (N_20839,N_15973,N_16557);
or U20840 (N_20840,N_18531,N_17770);
or U20841 (N_20841,N_17843,N_18464);
and U20842 (N_20842,N_17886,N_17742);
nor U20843 (N_20843,N_16538,N_18454);
nand U20844 (N_20844,N_18676,N_17769);
nand U20845 (N_20845,N_17680,N_17251);
xnor U20846 (N_20846,N_18274,N_15821);
xor U20847 (N_20847,N_16470,N_18290);
nor U20848 (N_20848,N_16753,N_18373);
and U20849 (N_20849,N_16453,N_15674);
nand U20850 (N_20850,N_18075,N_16006);
nor U20851 (N_20851,N_17536,N_15649);
xor U20852 (N_20852,N_17985,N_17751);
nor U20853 (N_20853,N_18431,N_17772);
xnor U20854 (N_20854,N_15631,N_18215);
xnor U20855 (N_20855,N_18320,N_18602);
and U20856 (N_20856,N_17819,N_17837);
or U20857 (N_20857,N_16383,N_16049);
and U20858 (N_20858,N_16170,N_18625);
xor U20859 (N_20859,N_16604,N_17847);
nand U20860 (N_20860,N_16705,N_15798);
nor U20861 (N_20861,N_16918,N_16142);
nor U20862 (N_20862,N_17256,N_16260);
xor U20863 (N_20863,N_17843,N_16480);
or U20864 (N_20864,N_16932,N_17424);
nor U20865 (N_20865,N_18729,N_17675);
nor U20866 (N_20866,N_18143,N_17188);
nand U20867 (N_20867,N_15870,N_18217);
xnor U20868 (N_20868,N_17869,N_18140);
and U20869 (N_20869,N_16054,N_18098);
and U20870 (N_20870,N_17553,N_18484);
nor U20871 (N_20871,N_17793,N_17838);
and U20872 (N_20872,N_16006,N_16957);
and U20873 (N_20873,N_16657,N_16695);
and U20874 (N_20874,N_16359,N_17197);
or U20875 (N_20875,N_17507,N_15827);
nor U20876 (N_20876,N_16613,N_18046);
nand U20877 (N_20877,N_17693,N_16777);
nor U20878 (N_20878,N_15804,N_16915);
nand U20879 (N_20879,N_15792,N_17169);
xnor U20880 (N_20880,N_17354,N_16661);
nor U20881 (N_20881,N_15784,N_17161);
xnor U20882 (N_20882,N_17275,N_16442);
or U20883 (N_20883,N_18692,N_17082);
nand U20884 (N_20884,N_17699,N_17578);
nand U20885 (N_20885,N_18318,N_17485);
nor U20886 (N_20886,N_16349,N_18188);
xnor U20887 (N_20887,N_17303,N_16964);
nand U20888 (N_20888,N_18721,N_17172);
nand U20889 (N_20889,N_15766,N_16519);
nor U20890 (N_20890,N_18685,N_16715);
or U20891 (N_20891,N_17825,N_17735);
xnor U20892 (N_20892,N_17812,N_17453);
nor U20893 (N_20893,N_17666,N_15907);
nand U20894 (N_20894,N_18005,N_15689);
or U20895 (N_20895,N_16542,N_16084);
nor U20896 (N_20896,N_17502,N_18491);
or U20897 (N_20897,N_18162,N_17118);
xor U20898 (N_20898,N_16741,N_17538);
nand U20899 (N_20899,N_15796,N_17070);
or U20900 (N_20900,N_16829,N_15940);
xor U20901 (N_20901,N_17264,N_15823);
xor U20902 (N_20902,N_16299,N_17800);
or U20903 (N_20903,N_15730,N_15739);
and U20904 (N_20904,N_17995,N_16477);
xor U20905 (N_20905,N_16908,N_18521);
or U20906 (N_20906,N_17861,N_18231);
nand U20907 (N_20907,N_17687,N_17816);
xnor U20908 (N_20908,N_17354,N_17601);
nand U20909 (N_20909,N_17407,N_18091);
or U20910 (N_20910,N_16333,N_17212);
nand U20911 (N_20911,N_17541,N_17077);
or U20912 (N_20912,N_18316,N_16491);
nand U20913 (N_20913,N_16745,N_17675);
or U20914 (N_20914,N_16785,N_16589);
and U20915 (N_20915,N_17527,N_16802);
or U20916 (N_20916,N_16535,N_16104);
xnor U20917 (N_20917,N_17520,N_15855);
or U20918 (N_20918,N_16929,N_16703);
nor U20919 (N_20919,N_17161,N_18417);
and U20920 (N_20920,N_17540,N_17213);
or U20921 (N_20921,N_15779,N_17100);
or U20922 (N_20922,N_16168,N_18709);
xor U20923 (N_20923,N_17418,N_16075);
xor U20924 (N_20924,N_16177,N_17899);
or U20925 (N_20925,N_18375,N_18369);
nand U20926 (N_20926,N_18618,N_16601);
or U20927 (N_20927,N_18351,N_16450);
and U20928 (N_20928,N_18243,N_17793);
nor U20929 (N_20929,N_18628,N_17315);
nor U20930 (N_20930,N_17935,N_16979);
or U20931 (N_20931,N_16125,N_17654);
nor U20932 (N_20932,N_18564,N_17221);
nor U20933 (N_20933,N_17432,N_17774);
nor U20934 (N_20934,N_17183,N_17135);
nand U20935 (N_20935,N_18506,N_16516);
nor U20936 (N_20936,N_16937,N_18655);
xnor U20937 (N_20937,N_15892,N_18720);
nand U20938 (N_20938,N_18360,N_16743);
nor U20939 (N_20939,N_17004,N_17334);
and U20940 (N_20940,N_18245,N_16373);
and U20941 (N_20941,N_16848,N_17303);
or U20942 (N_20942,N_17808,N_17496);
xor U20943 (N_20943,N_17676,N_17873);
and U20944 (N_20944,N_16800,N_16917);
and U20945 (N_20945,N_17334,N_17396);
xnor U20946 (N_20946,N_18492,N_15896);
or U20947 (N_20947,N_17426,N_15854);
and U20948 (N_20948,N_17092,N_18017);
or U20949 (N_20949,N_18077,N_15763);
nand U20950 (N_20950,N_16605,N_17401);
nor U20951 (N_20951,N_16596,N_18719);
or U20952 (N_20952,N_18138,N_18619);
xor U20953 (N_20953,N_16964,N_17328);
nand U20954 (N_20954,N_17627,N_16831);
and U20955 (N_20955,N_16398,N_17676);
or U20956 (N_20956,N_15703,N_16185);
and U20957 (N_20957,N_16273,N_17459);
or U20958 (N_20958,N_15935,N_17743);
nor U20959 (N_20959,N_18105,N_17470);
xor U20960 (N_20960,N_16299,N_16954);
and U20961 (N_20961,N_15801,N_18577);
and U20962 (N_20962,N_16739,N_17656);
and U20963 (N_20963,N_17489,N_17200);
and U20964 (N_20964,N_16122,N_15825);
nor U20965 (N_20965,N_17618,N_17643);
nor U20966 (N_20966,N_15860,N_16707);
xnor U20967 (N_20967,N_16817,N_17565);
or U20968 (N_20968,N_18376,N_16665);
xor U20969 (N_20969,N_15830,N_18498);
nand U20970 (N_20970,N_17049,N_17859);
xor U20971 (N_20971,N_16865,N_17395);
xor U20972 (N_20972,N_16185,N_16028);
nor U20973 (N_20973,N_16062,N_16533);
nand U20974 (N_20974,N_17944,N_16143);
or U20975 (N_20975,N_15769,N_16719);
nor U20976 (N_20976,N_18334,N_18210);
and U20977 (N_20977,N_16384,N_18152);
and U20978 (N_20978,N_17716,N_16231);
nor U20979 (N_20979,N_18098,N_17857);
and U20980 (N_20980,N_15824,N_15671);
xnor U20981 (N_20981,N_16883,N_16685);
or U20982 (N_20982,N_15896,N_15734);
xnor U20983 (N_20983,N_18660,N_17827);
nor U20984 (N_20984,N_17508,N_17636);
nor U20985 (N_20985,N_18603,N_16885);
nand U20986 (N_20986,N_17932,N_15752);
xnor U20987 (N_20987,N_15716,N_17539);
nand U20988 (N_20988,N_16925,N_17110);
and U20989 (N_20989,N_15702,N_18060);
nor U20990 (N_20990,N_16512,N_15666);
and U20991 (N_20991,N_17241,N_18711);
xnor U20992 (N_20992,N_18388,N_17709);
or U20993 (N_20993,N_16465,N_16771);
and U20994 (N_20994,N_16498,N_16372);
xnor U20995 (N_20995,N_15765,N_17990);
nor U20996 (N_20996,N_15669,N_17110);
or U20997 (N_20997,N_16342,N_17436);
or U20998 (N_20998,N_17354,N_15639);
or U20999 (N_20999,N_15983,N_15711);
nor U21000 (N_21000,N_18337,N_17121);
xor U21001 (N_21001,N_16184,N_17075);
and U21002 (N_21002,N_17370,N_17424);
xor U21003 (N_21003,N_18637,N_16053);
nor U21004 (N_21004,N_15806,N_16434);
nor U21005 (N_21005,N_17260,N_18575);
nor U21006 (N_21006,N_15887,N_16670);
nor U21007 (N_21007,N_17076,N_18595);
nand U21008 (N_21008,N_15702,N_17578);
or U21009 (N_21009,N_16686,N_18575);
nor U21010 (N_21010,N_16602,N_17170);
xor U21011 (N_21011,N_17045,N_17420);
or U21012 (N_21012,N_15835,N_16419);
nand U21013 (N_21013,N_17819,N_15813);
nand U21014 (N_21014,N_18743,N_16755);
xnor U21015 (N_21015,N_18686,N_17181);
nor U21016 (N_21016,N_18295,N_17984);
or U21017 (N_21017,N_16199,N_18543);
nor U21018 (N_21018,N_16235,N_18446);
and U21019 (N_21019,N_17069,N_15688);
nand U21020 (N_21020,N_17848,N_18255);
nand U21021 (N_21021,N_15635,N_18562);
nand U21022 (N_21022,N_16985,N_18625);
nor U21023 (N_21023,N_17970,N_18260);
or U21024 (N_21024,N_18065,N_15906);
xor U21025 (N_21025,N_17585,N_16448);
nand U21026 (N_21026,N_18427,N_17428);
nor U21027 (N_21027,N_17368,N_16816);
or U21028 (N_21028,N_17359,N_15829);
nand U21029 (N_21029,N_16437,N_18602);
xnor U21030 (N_21030,N_18443,N_15893);
nor U21031 (N_21031,N_18142,N_16835);
xor U21032 (N_21032,N_16830,N_17914);
xor U21033 (N_21033,N_16902,N_18175);
nand U21034 (N_21034,N_16809,N_17081);
or U21035 (N_21035,N_17145,N_17366);
nor U21036 (N_21036,N_18192,N_16722);
nor U21037 (N_21037,N_17445,N_16017);
xnor U21038 (N_21038,N_16916,N_16998);
nand U21039 (N_21039,N_15686,N_17088);
or U21040 (N_21040,N_16541,N_17881);
or U21041 (N_21041,N_18725,N_16362);
nand U21042 (N_21042,N_16740,N_16376);
nand U21043 (N_21043,N_17088,N_16803);
or U21044 (N_21044,N_16270,N_17481);
and U21045 (N_21045,N_17368,N_16328);
and U21046 (N_21046,N_17115,N_16466);
nor U21047 (N_21047,N_16329,N_15942);
or U21048 (N_21048,N_18149,N_16570);
or U21049 (N_21049,N_18114,N_18329);
xnor U21050 (N_21050,N_18496,N_17040);
nor U21051 (N_21051,N_17005,N_17589);
xor U21052 (N_21052,N_17938,N_17777);
and U21053 (N_21053,N_18661,N_17142);
nor U21054 (N_21054,N_16219,N_17603);
nor U21055 (N_21055,N_16678,N_18720);
and U21056 (N_21056,N_18046,N_15779);
nor U21057 (N_21057,N_18506,N_18619);
xnor U21058 (N_21058,N_17130,N_17374);
nand U21059 (N_21059,N_18335,N_16281);
xnor U21060 (N_21060,N_17142,N_16782);
xnor U21061 (N_21061,N_16333,N_16521);
and U21062 (N_21062,N_18704,N_18178);
nand U21063 (N_21063,N_17198,N_16290);
nand U21064 (N_21064,N_17628,N_16341);
xnor U21065 (N_21065,N_16115,N_18177);
nor U21066 (N_21066,N_17043,N_17693);
or U21067 (N_21067,N_17429,N_15891);
or U21068 (N_21068,N_18289,N_18089);
or U21069 (N_21069,N_17516,N_18303);
nor U21070 (N_21070,N_16220,N_16566);
nor U21071 (N_21071,N_16473,N_16594);
nand U21072 (N_21072,N_17411,N_17443);
nand U21073 (N_21073,N_16813,N_17765);
and U21074 (N_21074,N_18265,N_18295);
or U21075 (N_21075,N_17530,N_16466);
xnor U21076 (N_21076,N_16845,N_18414);
xnor U21077 (N_21077,N_16031,N_18335);
and U21078 (N_21078,N_16294,N_17354);
or U21079 (N_21079,N_17439,N_18224);
nand U21080 (N_21080,N_16802,N_16298);
nor U21081 (N_21081,N_16459,N_16900);
nor U21082 (N_21082,N_15942,N_18008);
or U21083 (N_21083,N_16846,N_17626);
or U21084 (N_21084,N_16052,N_15776);
xnor U21085 (N_21085,N_16008,N_16744);
nand U21086 (N_21086,N_15751,N_17894);
nand U21087 (N_21087,N_15760,N_18284);
nand U21088 (N_21088,N_18105,N_17234);
or U21089 (N_21089,N_18681,N_18565);
and U21090 (N_21090,N_17258,N_17873);
and U21091 (N_21091,N_18015,N_15967);
nand U21092 (N_21092,N_17984,N_17474);
nand U21093 (N_21093,N_17425,N_17621);
nor U21094 (N_21094,N_16123,N_16298);
nor U21095 (N_21095,N_17712,N_15684);
or U21096 (N_21096,N_16704,N_16788);
xor U21097 (N_21097,N_17198,N_17691);
nor U21098 (N_21098,N_17851,N_17422);
nand U21099 (N_21099,N_18351,N_17988);
nor U21100 (N_21100,N_18306,N_17345);
nand U21101 (N_21101,N_17915,N_18669);
nor U21102 (N_21102,N_16251,N_16784);
nand U21103 (N_21103,N_15723,N_17476);
xnor U21104 (N_21104,N_17000,N_17303);
xnor U21105 (N_21105,N_17547,N_18489);
xor U21106 (N_21106,N_17714,N_17756);
nor U21107 (N_21107,N_17826,N_15850);
xnor U21108 (N_21108,N_17941,N_15887);
xnor U21109 (N_21109,N_17576,N_17766);
nand U21110 (N_21110,N_16408,N_18194);
nor U21111 (N_21111,N_16478,N_18595);
xnor U21112 (N_21112,N_17461,N_16108);
nor U21113 (N_21113,N_18144,N_17506);
and U21114 (N_21114,N_15689,N_15773);
nand U21115 (N_21115,N_16316,N_18369);
xnor U21116 (N_21116,N_17050,N_17377);
and U21117 (N_21117,N_18467,N_17594);
nand U21118 (N_21118,N_17753,N_16110);
and U21119 (N_21119,N_15786,N_18419);
xor U21120 (N_21120,N_16148,N_16043);
or U21121 (N_21121,N_16931,N_16443);
or U21122 (N_21122,N_17113,N_15917);
or U21123 (N_21123,N_16331,N_17912);
nand U21124 (N_21124,N_17627,N_17542);
or U21125 (N_21125,N_17158,N_16861);
and U21126 (N_21126,N_16679,N_15759);
or U21127 (N_21127,N_16347,N_16776);
or U21128 (N_21128,N_17991,N_16446);
nand U21129 (N_21129,N_17975,N_18568);
or U21130 (N_21130,N_16359,N_17180);
xnor U21131 (N_21131,N_17403,N_15791);
or U21132 (N_21132,N_17673,N_17385);
nand U21133 (N_21133,N_17119,N_17512);
and U21134 (N_21134,N_18642,N_16617);
nor U21135 (N_21135,N_17210,N_17514);
and U21136 (N_21136,N_18485,N_17844);
nand U21137 (N_21137,N_17479,N_15785);
nor U21138 (N_21138,N_17916,N_18462);
and U21139 (N_21139,N_16797,N_17613);
xor U21140 (N_21140,N_18311,N_16775);
and U21141 (N_21141,N_18578,N_16232);
nor U21142 (N_21142,N_17772,N_15627);
and U21143 (N_21143,N_17317,N_18115);
nor U21144 (N_21144,N_16222,N_17984);
or U21145 (N_21145,N_16277,N_18277);
or U21146 (N_21146,N_18533,N_17941);
and U21147 (N_21147,N_17961,N_17807);
nor U21148 (N_21148,N_16304,N_18117);
nor U21149 (N_21149,N_15815,N_17937);
and U21150 (N_21150,N_15827,N_15937);
or U21151 (N_21151,N_17961,N_18566);
or U21152 (N_21152,N_17102,N_17971);
nor U21153 (N_21153,N_16731,N_16730);
nor U21154 (N_21154,N_16768,N_18425);
nand U21155 (N_21155,N_16598,N_16664);
or U21156 (N_21156,N_17150,N_18462);
nor U21157 (N_21157,N_17981,N_15663);
nor U21158 (N_21158,N_18218,N_17967);
nand U21159 (N_21159,N_17531,N_15777);
or U21160 (N_21160,N_16717,N_15980);
nand U21161 (N_21161,N_17011,N_15649);
nand U21162 (N_21162,N_18466,N_17199);
nand U21163 (N_21163,N_16817,N_15785);
nand U21164 (N_21164,N_16466,N_16412);
nand U21165 (N_21165,N_16094,N_16061);
and U21166 (N_21166,N_16997,N_18412);
nor U21167 (N_21167,N_18335,N_17347);
nor U21168 (N_21168,N_16930,N_18450);
and U21169 (N_21169,N_16660,N_16382);
and U21170 (N_21170,N_17689,N_16068);
or U21171 (N_21171,N_18217,N_18385);
xnor U21172 (N_21172,N_17916,N_16558);
nor U21173 (N_21173,N_18520,N_16310);
nor U21174 (N_21174,N_18442,N_17406);
nor U21175 (N_21175,N_15716,N_18040);
xor U21176 (N_21176,N_17091,N_17627);
or U21177 (N_21177,N_17172,N_18379);
xor U21178 (N_21178,N_15937,N_17679);
and U21179 (N_21179,N_18206,N_15941);
xor U21180 (N_21180,N_16600,N_18632);
xor U21181 (N_21181,N_16357,N_15967);
xnor U21182 (N_21182,N_16002,N_17510);
or U21183 (N_21183,N_18535,N_16425);
and U21184 (N_21184,N_18547,N_16247);
or U21185 (N_21185,N_18385,N_17682);
and U21186 (N_21186,N_16128,N_16782);
nand U21187 (N_21187,N_17923,N_18158);
and U21188 (N_21188,N_17248,N_15726);
and U21189 (N_21189,N_18069,N_16974);
xor U21190 (N_21190,N_16410,N_17875);
or U21191 (N_21191,N_15952,N_16613);
nand U21192 (N_21192,N_17076,N_18567);
and U21193 (N_21193,N_16888,N_16380);
and U21194 (N_21194,N_17627,N_18328);
nand U21195 (N_21195,N_15897,N_17610);
nor U21196 (N_21196,N_16319,N_18413);
nor U21197 (N_21197,N_17576,N_16058);
nor U21198 (N_21198,N_18541,N_18443);
or U21199 (N_21199,N_18322,N_18116);
and U21200 (N_21200,N_17413,N_16147);
nor U21201 (N_21201,N_16883,N_16899);
xor U21202 (N_21202,N_18475,N_17835);
nand U21203 (N_21203,N_17660,N_18103);
or U21204 (N_21204,N_17011,N_15868);
or U21205 (N_21205,N_15643,N_16626);
xnor U21206 (N_21206,N_16438,N_16590);
or U21207 (N_21207,N_15859,N_16010);
nand U21208 (N_21208,N_17845,N_16169);
xnor U21209 (N_21209,N_16256,N_16737);
nor U21210 (N_21210,N_15908,N_15962);
xor U21211 (N_21211,N_16292,N_15655);
nor U21212 (N_21212,N_17456,N_16964);
and U21213 (N_21213,N_16227,N_17927);
xnor U21214 (N_21214,N_18689,N_16319);
xnor U21215 (N_21215,N_17666,N_17124);
and U21216 (N_21216,N_17380,N_17443);
nand U21217 (N_21217,N_18262,N_17220);
xor U21218 (N_21218,N_17405,N_15919);
nand U21219 (N_21219,N_17729,N_17547);
or U21220 (N_21220,N_17852,N_16865);
or U21221 (N_21221,N_17390,N_16707);
nand U21222 (N_21222,N_17976,N_17755);
nor U21223 (N_21223,N_17764,N_17441);
nor U21224 (N_21224,N_18275,N_16750);
nand U21225 (N_21225,N_15633,N_15913);
nand U21226 (N_21226,N_18745,N_17270);
or U21227 (N_21227,N_17056,N_16533);
xnor U21228 (N_21228,N_18617,N_18111);
or U21229 (N_21229,N_16363,N_17280);
and U21230 (N_21230,N_16924,N_17405);
nand U21231 (N_21231,N_16118,N_16132);
nor U21232 (N_21232,N_17109,N_16879);
or U21233 (N_21233,N_16322,N_18698);
nand U21234 (N_21234,N_18486,N_15999);
and U21235 (N_21235,N_17960,N_16390);
or U21236 (N_21236,N_18272,N_17385);
or U21237 (N_21237,N_15706,N_18548);
or U21238 (N_21238,N_15754,N_16767);
xor U21239 (N_21239,N_16721,N_15963);
nand U21240 (N_21240,N_18528,N_17796);
and U21241 (N_21241,N_16193,N_15716);
nand U21242 (N_21242,N_16208,N_17036);
xor U21243 (N_21243,N_15761,N_16836);
or U21244 (N_21244,N_17583,N_16654);
nor U21245 (N_21245,N_15749,N_16015);
nand U21246 (N_21246,N_15710,N_16416);
nor U21247 (N_21247,N_17398,N_18081);
xor U21248 (N_21248,N_18289,N_18585);
nand U21249 (N_21249,N_15655,N_16520);
or U21250 (N_21250,N_17178,N_18115);
and U21251 (N_21251,N_16348,N_17644);
nor U21252 (N_21252,N_18166,N_16614);
nor U21253 (N_21253,N_16898,N_18178);
nand U21254 (N_21254,N_17315,N_16231);
nor U21255 (N_21255,N_16660,N_16612);
or U21256 (N_21256,N_18234,N_18244);
nand U21257 (N_21257,N_15822,N_17796);
or U21258 (N_21258,N_16121,N_16147);
xor U21259 (N_21259,N_16007,N_17724);
nor U21260 (N_21260,N_16734,N_18547);
nor U21261 (N_21261,N_16797,N_16735);
xnor U21262 (N_21262,N_17654,N_15963);
xor U21263 (N_21263,N_16905,N_18501);
nand U21264 (N_21264,N_16066,N_16440);
or U21265 (N_21265,N_15835,N_16166);
or U21266 (N_21266,N_17396,N_15655);
nand U21267 (N_21267,N_16671,N_16808);
or U21268 (N_21268,N_17153,N_18288);
nand U21269 (N_21269,N_16969,N_17762);
nor U21270 (N_21270,N_17159,N_17573);
or U21271 (N_21271,N_16880,N_18566);
nor U21272 (N_21272,N_16736,N_18107);
nor U21273 (N_21273,N_17638,N_16005);
nand U21274 (N_21274,N_17907,N_18469);
or U21275 (N_21275,N_16507,N_15785);
and U21276 (N_21276,N_16525,N_17353);
nand U21277 (N_21277,N_18603,N_17235);
and U21278 (N_21278,N_18660,N_16645);
and U21279 (N_21279,N_16259,N_16677);
and U21280 (N_21280,N_18386,N_17846);
or U21281 (N_21281,N_16333,N_18740);
or U21282 (N_21282,N_18384,N_17747);
nor U21283 (N_21283,N_16167,N_18492);
and U21284 (N_21284,N_17412,N_18021);
and U21285 (N_21285,N_18332,N_17637);
and U21286 (N_21286,N_17619,N_16078);
or U21287 (N_21287,N_15974,N_17930);
nor U21288 (N_21288,N_16591,N_18670);
or U21289 (N_21289,N_15729,N_16121);
and U21290 (N_21290,N_17081,N_18401);
xnor U21291 (N_21291,N_17554,N_18065);
nor U21292 (N_21292,N_18700,N_18648);
or U21293 (N_21293,N_16225,N_17577);
nor U21294 (N_21294,N_17184,N_17655);
and U21295 (N_21295,N_17036,N_16850);
nand U21296 (N_21296,N_17575,N_17145);
nand U21297 (N_21297,N_16892,N_17775);
xnor U21298 (N_21298,N_16468,N_18518);
xnor U21299 (N_21299,N_16574,N_17787);
or U21300 (N_21300,N_16159,N_16947);
and U21301 (N_21301,N_16221,N_15630);
or U21302 (N_21302,N_17659,N_16395);
and U21303 (N_21303,N_17397,N_17376);
or U21304 (N_21304,N_17894,N_15783);
xnor U21305 (N_21305,N_16585,N_17532);
xnor U21306 (N_21306,N_16500,N_18596);
xor U21307 (N_21307,N_15881,N_18561);
or U21308 (N_21308,N_15627,N_16270);
nor U21309 (N_21309,N_15729,N_16125);
or U21310 (N_21310,N_17971,N_16177);
xor U21311 (N_21311,N_18089,N_17303);
or U21312 (N_21312,N_16315,N_17314);
xnor U21313 (N_21313,N_18606,N_17383);
or U21314 (N_21314,N_17371,N_16045);
or U21315 (N_21315,N_16914,N_17493);
and U21316 (N_21316,N_16956,N_16358);
or U21317 (N_21317,N_16202,N_17120);
and U21318 (N_21318,N_18372,N_15941);
or U21319 (N_21319,N_16148,N_16487);
nor U21320 (N_21320,N_17446,N_16883);
or U21321 (N_21321,N_16248,N_17744);
xnor U21322 (N_21322,N_16135,N_18236);
and U21323 (N_21323,N_18628,N_17517);
or U21324 (N_21324,N_18558,N_17254);
and U21325 (N_21325,N_15973,N_16769);
nand U21326 (N_21326,N_18642,N_16257);
nand U21327 (N_21327,N_16369,N_16045);
xor U21328 (N_21328,N_16815,N_16561);
xor U21329 (N_21329,N_17559,N_18024);
xor U21330 (N_21330,N_17808,N_16171);
nand U21331 (N_21331,N_17892,N_17487);
or U21332 (N_21332,N_17512,N_16174);
xnor U21333 (N_21333,N_15873,N_16110);
xnor U21334 (N_21334,N_16003,N_17358);
nor U21335 (N_21335,N_17167,N_17487);
xnor U21336 (N_21336,N_17837,N_16619);
nand U21337 (N_21337,N_16885,N_16866);
or U21338 (N_21338,N_17419,N_16045);
or U21339 (N_21339,N_17668,N_16195);
or U21340 (N_21340,N_16723,N_17326);
and U21341 (N_21341,N_15739,N_16282);
nor U21342 (N_21342,N_16497,N_16176);
nand U21343 (N_21343,N_16220,N_17940);
or U21344 (N_21344,N_16205,N_16091);
nor U21345 (N_21345,N_17500,N_15817);
nand U21346 (N_21346,N_17936,N_16376);
xor U21347 (N_21347,N_18277,N_18630);
xnor U21348 (N_21348,N_17743,N_15782);
and U21349 (N_21349,N_18162,N_17029);
nand U21350 (N_21350,N_16803,N_17717);
and U21351 (N_21351,N_18407,N_17527);
xor U21352 (N_21352,N_16767,N_17729);
and U21353 (N_21353,N_17140,N_16991);
xor U21354 (N_21354,N_17426,N_17491);
and U21355 (N_21355,N_15849,N_16565);
or U21356 (N_21356,N_15668,N_17924);
nand U21357 (N_21357,N_18364,N_17584);
or U21358 (N_21358,N_15826,N_17246);
nor U21359 (N_21359,N_18556,N_16022);
nand U21360 (N_21360,N_16250,N_15696);
xor U21361 (N_21361,N_17785,N_16675);
nand U21362 (N_21362,N_17581,N_17655);
or U21363 (N_21363,N_17913,N_17231);
and U21364 (N_21364,N_17579,N_16590);
and U21365 (N_21365,N_16540,N_16114);
xor U21366 (N_21366,N_16852,N_17659);
or U21367 (N_21367,N_16592,N_16298);
nand U21368 (N_21368,N_18183,N_15777);
and U21369 (N_21369,N_17994,N_15802);
xnor U21370 (N_21370,N_18687,N_17283);
and U21371 (N_21371,N_15787,N_16049);
nor U21372 (N_21372,N_17210,N_18025);
nand U21373 (N_21373,N_17087,N_16402);
nor U21374 (N_21374,N_15918,N_17201);
nand U21375 (N_21375,N_17270,N_16181);
nand U21376 (N_21376,N_17779,N_17583);
nor U21377 (N_21377,N_17397,N_16309);
and U21378 (N_21378,N_18578,N_17552);
or U21379 (N_21379,N_16648,N_16225);
xnor U21380 (N_21380,N_18643,N_18320);
and U21381 (N_21381,N_16665,N_16147);
or U21382 (N_21382,N_16623,N_17551);
or U21383 (N_21383,N_17714,N_17675);
nor U21384 (N_21384,N_16238,N_18049);
nor U21385 (N_21385,N_15766,N_17625);
nand U21386 (N_21386,N_16985,N_16674);
nand U21387 (N_21387,N_16282,N_16832);
and U21388 (N_21388,N_17510,N_17631);
nand U21389 (N_21389,N_16307,N_16318);
nor U21390 (N_21390,N_16372,N_17889);
xor U21391 (N_21391,N_17569,N_18674);
nor U21392 (N_21392,N_17081,N_16055);
or U21393 (N_21393,N_17750,N_16379);
xnor U21394 (N_21394,N_15827,N_17495);
xnor U21395 (N_21395,N_17711,N_18577);
and U21396 (N_21396,N_18305,N_17138);
nand U21397 (N_21397,N_16886,N_16139);
and U21398 (N_21398,N_17749,N_17614);
and U21399 (N_21399,N_15839,N_17550);
and U21400 (N_21400,N_16300,N_17150);
or U21401 (N_21401,N_16490,N_16295);
or U21402 (N_21402,N_18583,N_16422);
or U21403 (N_21403,N_18356,N_16590);
xor U21404 (N_21404,N_18012,N_17288);
nor U21405 (N_21405,N_17096,N_16995);
or U21406 (N_21406,N_18259,N_17133);
and U21407 (N_21407,N_18702,N_17277);
or U21408 (N_21408,N_16743,N_18246);
or U21409 (N_21409,N_17761,N_18631);
nand U21410 (N_21410,N_17519,N_18139);
and U21411 (N_21411,N_16890,N_18266);
xor U21412 (N_21412,N_18059,N_16198);
nor U21413 (N_21413,N_16710,N_17922);
nand U21414 (N_21414,N_18497,N_17374);
nand U21415 (N_21415,N_17361,N_17079);
xnor U21416 (N_21416,N_16758,N_17555);
xor U21417 (N_21417,N_16161,N_17159);
and U21418 (N_21418,N_16821,N_18252);
xnor U21419 (N_21419,N_16460,N_16351);
or U21420 (N_21420,N_16826,N_16519);
nand U21421 (N_21421,N_17331,N_16716);
nor U21422 (N_21422,N_15922,N_15677);
xor U21423 (N_21423,N_18115,N_16914);
and U21424 (N_21424,N_15789,N_18661);
and U21425 (N_21425,N_16761,N_18210);
or U21426 (N_21426,N_18654,N_16188);
nand U21427 (N_21427,N_16951,N_15783);
and U21428 (N_21428,N_16367,N_17648);
nand U21429 (N_21429,N_17683,N_17895);
nand U21430 (N_21430,N_16107,N_18261);
nand U21431 (N_21431,N_18718,N_15766);
nor U21432 (N_21432,N_16840,N_15724);
or U21433 (N_21433,N_15914,N_15976);
or U21434 (N_21434,N_17380,N_17066);
and U21435 (N_21435,N_18398,N_17905);
nor U21436 (N_21436,N_17168,N_17740);
nor U21437 (N_21437,N_17234,N_17239);
xor U21438 (N_21438,N_18438,N_17790);
nand U21439 (N_21439,N_17561,N_16533);
nor U21440 (N_21440,N_17989,N_17919);
or U21441 (N_21441,N_17991,N_18090);
nor U21442 (N_21442,N_15712,N_16084);
and U21443 (N_21443,N_15873,N_16298);
nor U21444 (N_21444,N_16137,N_15628);
and U21445 (N_21445,N_17312,N_15723);
or U21446 (N_21446,N_17322,N_15811);
and U21447 (N_21447,N_16974,N_16030);
nor U21448 (N_21448,N_16322,N_17501);
and U21449 (N_21449,N_16783,N_16234);
and U21450 (N_21450,N_18033,N_17795);
nand U21451 (N_21451,N_16991,N_16824);
or U21452 (N_21452,N_16905,N_16147);
xor U21453 (N_21453,N_17960,N_16768);
nand U21454 (N_21454,N_18164,N_16717);
nand U21455 (N_21455,N_16354,N_18617);
nand U21456 (N_21456,N_18744,N_15812);
xor U21457 (N_21457,N_17706,N_16146);
nor U21458 (N_21458,N_15826,N_16982);
and U21459 (N_21459,N_18368,N_18518);
nand U21460 (N_21460,N_16664,N_15953);
nand U21461 (N_21461,N_18249,N_18583);
or U21462 (N_21462,N_16907,N_17421);
nand U21463 (N_21463,N_17256,N_16218);
nor U21464 (N_21464,N_17380,N_18032);
and U21465 (N_21465,N_16985,N_18058);
and U21466 (N_21466,N_16617,N_16375);
or U21467 (N_21467,N_16253,N_17834);
xor U21468 (N_21468,N_16358,N_16451);
nor U21469 (N_21469,N_16725,N_17406);
or U21470 (N_21470,N_18279,N_17364);
nand U21471 (N_21471,N_18248,N_16938);
or U21472 (N_21472,N_18490,N_15790);
xor U21473 (N_21473,N_15651,N_15860);
nor U21474 (N_21474,N_18340,N_15682);
or U21475 (N_21475,N_15825,N_16730);
and U21476 (N_21476,N_17105,N_15819);
nor U21477 (N_21477,N_16446,N_16925);
nand U21478 (N_21478,N_18493,N_16911);
nand U21479 (N_21479,N_17234,N_15955);
or U21480 (N_21480,N_15970,N_17337);
xor U21481 (N_21481,N_16928,N_16140);
nand U21482 (N_21482,N_17422,N_17137);
and U21483 (N_21483,N_18152,N_18733);
and U21484 (N_21484,N_18217,N_18617);
nand U21485 (N_21485,N_18736,N_16848);
nand U21486 (N_21486,N_16133,N_15860);
nand U21487 (N_21487,N_17926,N_18645);
xnor U21488 (N_21488,N_17149,N_18054);
nor U21489 (N_21489,N_18446,N_17301);
nor U21490 (N_21490,N_16726,N_17663);
nand U21491 (N_21491,N_18728,N_16849);
nand U21492 (N_21492,N_17928,N_18375);
nand U21493 (N_21493,N_16585,N_16164);
nor U21494 (N_21494,N_17748,N_15930);
nand U21495 (N_21495,N_16502,N_18675);
nand U21496 (N_21496,N_15759,N_18158);
nand U21497 (N_21497,N_17321,N_17224);
nand U21498 (N_21498,N_17788,N_18178);
and U21499 (N_21499,N_16642,N_17265);
nand U21500 (N_21500,N_16665,N_16383);
or U21501 (N_21501,N_16340,N_16949);
or U21502 (N_21502,N_18480,N_18749);
and U21503 (N_21503,N_16962,N_15926);
or U21504 (N_21504,N_16905,N_16037);
and U21505 (N_21505,N_17664,N_17767);
and U21506 (N_21506,N_18695,N_17586);
nand U21507 (N_21507,N_17150,N_16920);
xnor U21508 (N_21508,N_17194,N_16453);
or U21509 (N_21509,N_16534,N_16412);
nand U21510 (N_21510,N_16149,N_17002);
and U21511 (N_21511,N_16096,N_18168);
nor U21512 (N_21512,N_16035,N_16641);
nor U21513 (N_21513,N_18608,N_18597);
or U21514 (N_21514,N_18533,N_18475);
xor U21515 (N_21515,N_17349,N_17914);
xnor U21516 (N_21516,N_16076,N_15770);
and U21517 (N_21517,N_15818,N_18037);
and U21518 (N_21518,N_16989,N_15905);
nor U21519 (N_21519,N_18490,N_17186);
and U21520 (N_21520,N_16747,N_16694);
nor U21521 (N_21521,N_16973,N_15856);
nor U21522 (N_21522,N_15943,N_17270);
nand U21523 (N_21523,N_18084,N_17620);
xor U21524 (N_21524,N_16936,N_18440);
nand U21525 (N_21525,N_16792,N_15955);
xnor U21526 (N_21526,N_16863,N_17676);
nand U21527 (N_21527,N_15961,N_16554);
and U21528 (N_21528,N_18526,N_18471);
nor U21529 (N_21529,N_16752,N_17646);
or U21530 (N_21530,N_16403,N_17459);
or U21531 (N_21531,N_17966,N_17586);
nand U21532 (N_21532,N_16286,N_17856);
nand U21533 (N_21533,N_18370,N_16832);
or U21534 (N_21534,N_17637,N_17690);
or U21535 (N_21535,N_18227,N_16206);
nor U21536 (N_21536,N_18219,N_16655);
or U21537 (N_21537,N_17427,N_17929);
and U21538 (N_21538,N_16182,N_18674);
xnor U21539 (N_21539,N_16040,N_17596);
nand U21540 (N_21540,N_15669,N_17182);
nand U21541 (N_21541,N_18276,N_18569);
nand U21542 (N_21542,N_18502,N_18624);
nand U21543 (N_21543,N_16359,N_15958);
xor U21544 (N_21544,N_18140,N_16600);
nor U21545 (N_21545,N_16585,N_15841);
nor U21546 (N_21546,N_17130,N_18627);
and U21547 (N_21547,N_18644,N_18457);
nor U21548 (N_21548,N_16211,N_18553);
and U21549 (N_21549,N_16733,N_16375);
nand U21550 (N_21550,N_16228,N_17276);
or U21551 (N_21551,N_16927,N_17719);
nor U21552 (N_21552,N_18256,N_17910);
or U21553 (N_21553,N_18580,N_16236);
xor U21554 (N_21554,N_16218,N_18143);
nor U21555 (N_21555,N_17525,N_16892);
nor U21556 (N_21556,N_17794,N_18704);
or U21557 (N_21557,N_18663,N_15899);
nand U21558 (N_21558,N_18449,N_16485);
and U21559 (N_21559,N_17544,N_17234);
or U21560 (N_21560,N_17004,N_18199);
xor U21561 (N_21561,N_16257,N_16162);
nor U21562 (N_21562,N_17537,N_16668);
xnor U21563 (N_21563,N_16077,N_17170);
xnor U21564 (N_21564,N_16019,N_17165);
xor U21565 (N_21565,N_18711,N_16609);
or U21566 (N_21566,N_16558,N_18405);
nor U21567 (N_21567,N_16129,N_18259);
or U21568 (N_21568,N_18189,N_17552);
xnor U21569 (N_21569,N_18314,N_16733);
or U21570 (N_21570,N_16615,N_15831);
xnor U21571 (N_21571,N_16089,N_17960);
nand U21572 (N_21572,N_17599,N_16061);
or U21573 (N_21573,N_15656,N_17094);
nor U21574 (N_21574,N_15687,N_15804);
nor U21575 (N_21575,N_16244,N_15972);
and U21576 (N_21576,N_17058,N_16986);
nand U21577 (N_21577,N_18113,N_15848);
or U21578 (N_21578,N_15913,N_16134);
or U21579 (N_21579,N_15905,N_18689);
or U21580 (N_21580,N_15977,N_18318);
nor U21581 (N_21581,N_18575,N_17576);
and U21582 (N_21582,N_16720,N_18152);
nand U21583 (N_21583,N_18188,N_17728);
nor U21584 (N_21584,N_18412,N_18350);
xor U21585 (N_21585,N_17453,N_16951);
nand U21586 (N_21586,N_18073,N_16047);
xor U21587 (N_21587,N_17051,N_18747);
or U21588 (N_21588,N_18447,N_18673);
and U21589 (N_21589,N_16569,N_16697);
nand U21590 (N_21590,N_16073,N_16313);
xor U21591 (N_21591,N_15847,N_16198);
xnor U21592 (N_21592,N_16452,N_16724);
and U21593 (N_21593,N_16038,N_18458);
and U21594 (N_21594,N_16186,N_16130);
or U21595 (N_21595,N_17741,N_15905);
or U21596 (N_21596,N_18712,N_16273);
nor U21597 (N_21597,N_18214,N_16750);
xnor U21598 (N_21598,N_18246,N_16778);
nor U21599 (N_21599,N_17959,N_16432);
nor U21600 (N_21600,N_15853,N_17183);
or U21601 (N_21601,N_18047,N_18522);
nor U21602 (N_21602,N_18292,N_16946);
nand U21603 (N_21603,N_17521,N_17073);
nor U21604 (N_21604,N_17619,N_16725);
and U21605 (N_21605,N_17166,N_15916);
xor U21606 (N_21606,N_16694,N_18053);
nand U21607 (N_21607,N_16854,N_17598);
nand U21608 (N_21608,N_16830,N_18074);
nor U21609 (N_21609,N_17525,N_15803);
nor U21610 (N_21610,N_18677,N_16787);
nor U21611 (N_21611,N_16907,N_15662);
nand U21612 (N_21612,N_16915,N_17592);
nand U21613 (N_21613,N_18653,N_15784);
or U21614 (N_21614,N_17819,N_18510);
or U21615 (N_21615,N_15639,N_17741);
nand U21616 (N_21616,N_16421,N_16656);
xor U21617 (N_21617,N_17856,N_16375);
or U21618 (N_21618,N_17274,N_17651);
and U21619 (N_21619,N_16055,N_16522);
xnor U21620 (N_21620,N_18253,N_17241);
nand U21621 (N_21621,N_16060,N_17249);
and U21622 (N_21622,N_15962,N_16829);
nor U21623 (N_21623,N_18063,N_16409);
and U21624 (N_21624,N_16089,N_16179);
or U21625 (N_21625,N_16932,N_15749);
xnor U21626 (N_21626,N_16722,N_18554);
nand U21627 (N_21627,N_18037,N_17571);
and U21628 (N_21628,N_16604,N_17522);
or U21629 (N_21629,N_18501,N_15879);
or U21630 (N_21630,N_16590,N_18328);
nand U21631 (N_21631,N_18009,N_16434);
and U21632 (N_21632,N_18681,N_17536);
nor U21633 (N_21633,N_17393,N_16789);
nor U21634 (N_21634,N_15890,N_16705);
or U21635 (N_21635,N_15904,N_17737);
nor U21636 (N_21636,N_15752,N_17012);
or U21637 (N_21637,N_15655,N_16437);
nand U21638 (N_21638,N_17233,N_17174);
or U21639 (N_21639,N_18288,N_18622);
or U21640 (N_21640,N_17264,N_16096);
nor U21641 (N_21641,N_17925,N_17608);
xor U21642 (N_21642,N_16628,N_18158);
nand U21643 (N_21643,N_15796,N_17396);
and U21644 (N_21644,N_15750,N_16643);
nor U21645 (N_21645,N_15860,N_17226);
nor U21646 (N_21646,N_16732,N_17117);
nand U21647 (N_21647,N_16499,N_16218);
nor U21648 (N_21648,N_16420,N_16796);
nand U21649 (N_21649,N_17081,N_15683);
or U21650 (N_21650,N_17861,N_15699);
or U21651 (N_21651,N_16387,N_17190);
and U21652 (N_21652,N_18118,N_16281);
or U21653 (N_21653,N_15867,N_18583);
xnor U21654 (N_21654,N_17132,N_16372);
and U21655 (N_21655,N_17098,N_17692);
and U21656 (N_21656,N_18601,N_18224);
and U21657 (N_21657,N_18126,N_17920);
and U21658 (N_21658,N_16155,N_17096);
nor U21659 (N_21659,N_17790,N_16002);
or U21660 (N_21660,N_18049,N_18074);
nor U21661 (N_21661,N_16498,N_16548);
or U21662 (N_21662,N_15834,N_16790);
nor U21663 (N_21663,N_17167,N_18222);
nand U21664 (N_21664,N_16534,N_17153);
nor U21665 (N_21665,N_17591,N_16504);
or U21666 (N_21666,N_16224,N_18033);
nand U21667 (N_21667,N_17913,N_16406);
xnor U21668 (N_21668,N_16928,N_18364);
or U21669 (N_21669,N_15755,N_18709);
or U21670 (N_21670,N_17216,N_17510);
or U21671 (N_21671,N_17346,N_16305);
and U21672 (N_21672,N_17592,N_18332);
nand U21673 (N_21673,N_17798,N_18163);
or U21674 (N_21674,N_18680,N_17849);
nor U21675 (N_21675,N_16948,N_18692);
xnor U21676 (N_21676,N_16463,N_17880);
and U21677 (N_21677,N_18200,N_17045);
or U21678 (N_21678,N_16423,N_17701);
or U21679 (N_21679,N_17279,N_17018);
and U21680 (N_21680,N_17247,N_17430);
and U21681 (N_21681,N_15655,N_15825);
nor U21682 (N_21682,N_16195,N_17969);
xor U21683 (N_21683,N_18197,N_18579);
xnor U21684 (N_21684,N_17731,N_15729);
nand U21685 (N_21685,N_17191,N_17521);
nand U21686 (N_21686,N_16442,N_17441);
or U21687 (N_21687,N_16762,N_18001);
nand U21688 (N_21688,N_17631,N_18625);
xnor U21689 (N_21689,N_15953,N_17069);
and U21690 (N_21690,N_17408,N_15634);
nor U21691 (N_21691,N_18645,N_16076);
or U21692 (N_21692,N_16590,N_17359);
xor U21693 (N_21693,N_17116,N_17844);
or U21694 (N_21694,N_17134,N_16578);
and U21695 (N_21695,N_16188,N_18325);
nor U21696 (N_21696,N_16972,N_18453);
nor U21697 (N_21697,N_16585,N_17238);
nand U21698 (N_21698,N_17469,N_17905);
nor U21699 (N_21699,N_18407,N_17259);
xor U21700 (N_21700,N_17950,N_15990);
nand U21701 (N_21701,N_15752,N_18260);
nand U21702 (N_21702,N_16785,N_16648);
nor U21703 (N_21703,N_17310,N_17468);
nor U21704 (N_21704,N_17426,N_16144);
nor U21705 (N_21705,N_15834,N_18623);
or U21706 (N_21706,N_18203,N_18649);
or U21707 (N_21707,N_17028,N_17104);
and U21708 (N_21708,N_17457,N_17172);
and U21709 (N_21709,N_17843,N_18609);
nand U21710 (N_21710,N_15918,N_17154);
nand U21711 (N_21711,N_17763,N_15858);
xor U21712 (N_21712,N_18297,N_18351);
xor U21713 (N_21713,N_16871,N_17529);
xnor U21714 (N_21714,N_17988,N_17249);
nor U21715 (N_21715,N_16163,N_17511);
nand U21716 (N_21716,N_18264,N_17795);
nor U21717 (N_21717,N_18423,N_16499);
nand U21718 (N_21718,N_17177,N_16822);
or U21719 (N_21719,N_17172,N_17102);
nor U21720 (N_21720,N_15715,N_15903);
or U21721 (N_21721,N_17206,N_17527);
and U21722 (N_21722,N_16544,N_17282);
or U21723 (N_21723,N_16316,N_16095);
or U21724 (N_21724,N_16651,N_17130);
xor U21725 (N_21725,N_17000,N_16972);
or U21726 (N_21726,N_17494,N_18354);
nor U21727 (N_21727,N_16551,N_18479);
xnor U21728 (N_21728,N_17915,N_15750);
xnor U21729 (N_21729,N_17610,N_17793);
nand U21730 (N_21730,N_16694,N_16285);
nor U21731 (N_21731,N_16390,N_15769);
nor U21732 (N_21732,N_16291,N_17953);
xnor U21733 (N_21733,N_18315,N_18047);
xor U21734 (N_21734,N_15812,N_17007);
or U21735 (N_21735,N_16136,N_15853);
nand U21736 (N_21736,N_17897,N_17356);
or U21737 (N_21737,N_16893,N_18037);
nor U21738 (N_21738,N_15688,N_18608);
nor U21739 (N_21739,N_17387,N_18193);
nor U21740 (N_21740,N_17260,N_17743);
xor U21741 (N_21741,N_17929,N_16604);
and U21742 (N_21742,N_17366,N_17760);
and U21743 (N_21743,N_17304,N_16839);
and U21744 (N_21744,N_18478,N_18296);
nor U21745 (N_21745,N_18181,N_17713);
or U21746 (N_21746,N_16893,N_17154);
nand U21747 (N_21747,N_17471,N_15936);
nand U21748 (N_21748,N_16527,N_16541);
and U21749 (N_21749,N_16306,N_16188);
nor U21750 (N_21750,N_15634,N_18065);
nand U21751 (N_21751,N_17192,N_17013);
and U21752 (N_21752,N_17362,N_17850);
nor U21753 (N_21753,N_17309,N_17650);
or U21754 (N_21754,N_17501,N_18138);
nand U21755 (N_21755,N_16878,N_18524);
nand U21756 (N_21756,N_17467,N_16908);
xor U21757 (N_21757,N_17212,N_15970);
nor U21758 (N_21758,N_15941,N_16001);
xnor U21759 (N_21759,N_17640,N_15925);
and U21760 (N_21760,N_17140,N_17874);
or U21761 (N_21761,N_18044,N_16800);
xor U21762 (N_21762,N_16322,N_18240);
nor U21763 (N_21763,N_18454,N_18536);
nor U21764 (N_21764,N_18206,N_16488);
and U21765 (N_21765,N_15701,N_16500);
nor U21766 (N_21766,N_16073,N_16796);
or U21767 (N_21767,N_17212,N_17881);
xor U21768 (N_21768,N_18036,N_16455);
nor U21769 (N_21769,N_16967,N_17751);
or U21770 (N_21770,N_15889,N_18304);
xor U21771 (N_21771,N_15965,N_16793);
nor U21772 (N_21772,N_18610,N_16325);
or U21773 (N_21773,N_16594,N_17519);
xnor U21774 (N_21774,N_17704,N_16396);
nor U21775 (N_21775,N_17910,N_17988);
nor U21776 (N_21776,N_16395,N_15814);
or U21777 (N_21777,N_18290,N_17210);
nor U21778 (N_21778,N_18708,N_17711);
and U21779 (N_21779,N_17175,N_15985);
xnor U21780 (N_21780,N_18650,N_17445);
nand U21781 (N_21781,N_17992,N_16638);
nor U21782 (N_21782,N_17878,N_15726);
xor U21783 (N_21783,N_16105,N_16708);
or U21784 (N_21784,N_17958,N_15823);
nand U21785 (N_21785,N_16483,N_17591);
nor U21786 (N_21786,N_16072,N_18260);
nand U21787 (N_21787,N_18636,N_18141);
nor U21788 (N_21788,N_16180,N_16684);
and U21789 (N_21789,N_16196,N_17506);
and U21790 (N_21790,N_17369,N_16662);
nand U21791 (N_21791,N_17728,N_15859);
nand U21792 (N_21792,N_15923,N_18007);
or U21793 (N_21793,N_15923,N_17279);
nand U21794 (N_21794,N_15862,N_17706);
or U21795 (N_21795,N_17194,N_16394);
nor U21796 (N_21796,N_16124,N_16357);
nor U21797 (N_21797,N_17684,N_16594);
nand U21798 (N_21798,N_17338,N_18306);
nand U21799 (N_21799,N_18356,N_17982);
xnor U21800 (N_21800,N_15981,N_17567);
and U21801 (N_21801,N_18261,N_17418);
xnor U21802 (N_21802,N_15666,N_15805);
xnor U21803 (N_21803,N_17011,N_18123);
nor U21804 (N_21804,N_18214,N_17422);
nor U21805 (N_21805,N_17768,N_16665);
nand U21806 (N_21806,N_18722,N_16519);
or U21807 (N_21807,N_17533,N_16374);
or U21808 (N_21808,N_18690,N_15736);
nand U21809 (N_21809,N_17713,N_17111);
and U21810 (N_21810,N_16853,N_17525);
and U21811 (N_21811,N_17694,N_18006);
nor U21812 (N_21812,N_15790,N_17285);
and U21813 (N_21813,N_18639,N_18102);
xnor U21814 (N_21814,N_16511,N_16968);
nor U21815 (N_21815,N_17350,N_17627);
xor U21816 (N_21816,N_17717,N_16266);
nand U21817 (N_21817,N_16428,N_16991);
xor U21818 (N_21818,N_17843,N_16789);
or U21819 (N_21819,N_16406,N_16580);
nor U21820 (N_21820,N_16794,N_15791);
and U21821 (N_21821,N_18533,N_18333);
nor U21822 (N_21822,N_15786,N_16984);
nor U21823 (N_21823,N_18426,N_16456);
xnor U21824 (N_21824,N_17181,N_17856);
and U21825 (N_21825,N_18600,N_16778);
and U21826 (N_21826,N_17276,N_16129);
xnor U21827 (N_21827,N_16852,N_18671);
or U21828 (N_21828,N_15962,N_16182);
nor U21829 (N_21829,N_15761,N_17954);
xor U21830 (N_21830,N_16730,N_15843);
xnor U21831 (N_21831,N_15912,N_17589);
nor U21832 (N_21832,N_17597,N_15793);
nor U21833 (N_21833,N_17725,N_15672);
and U21834 (N_21834,N_17748,N_15737);
or U21835 (N_21835,N_16363,N_15806);
or U21836 (N_21836,N_16084,N_15749);
xnor U21837 (N_21837,N_17663,N_17920);
nor U21838 (N_21838,N_16577,N_18600);
or U21839 (N_21839,N_16808,N_18664);
nor U21840 (N_21840,N_16507,N_17138);
nor U21841 (N_21841,N_18402,N_16480);
and U21842 (N_21842,N_18389,N_18655);
and U21843 (N_21843,N_17911,N_16254);
or U21844 (N_21844,N_17718,N_17209);
xor U21845 (N_21845,N_18179,N_17615);
xor U21846 (N_21846,N_16394,N_17516);
nor U21847 (N_21847,N_17396,N_15848);
or U21848 (N_21848,N_17481,N_16816);
and U21849 (N_21849,N_16210,N_16901);
or U21850 (N_21850,N_16584,N_16873);
and U21851 (N_21851,N_18531,N_17146);
nand U21852 (N_21852,N_17638,N_18380);
and U21853 (N_21853,N_15662,N_18194);
nor U21854 (N_21854,N_18644,N_15839);
nand U21855 (N_21855,N_15659,N_15673);
nand U21856 (N_21856,N_18680,N_15967);
or U21857 (N_21857,N_17596,N_18390);
xor U21858 (N_21858,N_16336,N_18337);
or U21859 (N_21859,N_17417,N_18639);
and U21860 (N_21860,N_16259,N_18359);
xnor U21861 (N_21861,N_17231,N_15964);
xor U21862 (N_21862,N_16564,N_18566);
nor U21863 (N_21863,N_17798,N_16566);
or U21864 (N_21864,N_16311,N_16482);
and U21865 (N_21865,N_15664,N_16415);
nor U21866 (N_21866,N_15767,N_16607);
nor U21867 (N_21867,N_16459,N_18687);
xnor U21868 (N_21868,N_16081,N_15881);
xnor U21869 (N_21869,N_17313,N_17635);
or U21870 (N_21870,N_15864,N_15629);
nor U21871 (N_21871,N_18124,N_15934);
xnor U21872 (N_21872,N_16122,N_17534);
and U21873 (N_21873,N_18709,N_16920);
nor U21874 (N_21874,N_17278,N_17731);
and U21875 (N_21875,N_20975,N_21047);
xor U21876 (N_21876,N_21435,N_20042);
and U21877 (N_21877,N_20798,N_20791);
and U21878 (N_21878,N_20530,N_18957);
nor U21879 (N_21879,N_19389,N_18963);
and U21880 (N_21880,N_19543,N_21443);
or U21881 (N_21881,N_20177,N_21065);
and U21882 (N_21882,N_20965,N_20990);
and U21883 (N_21883,N_20859,N_19070);
nor U21884 (N_21884,N_21067,N_19210);
nand U21885 (N_21885,N_19889,N_19770);
nor U21886 (N_21886,N_21105,N_20300);
xor U21887 (N_21887,N_19186,N_19209);
nand U21888 (N_21888,N_20688,N_20149);
nor U21889 (N_21889,N_20991,N_21217);
xor U21890 (N_21890,N_19379,N_20871);
and U21891 (N_21891,N_21606,N_19040);
nor U21892 (N_21892,N_20396,N_20727);
xor U21893 (N_21893,N_20045,N_20813);
xor U21894 (N_21894,N_21235,N_19973);
xor U21895 (N_21895,N_20610,N_20782);
nor U21896 (N_21896,N_20778,N_20661);
and U21897 (N_21897,N_19666,N_21275);
and U21898 (N_21898,N_20186,N_21501);
and U21899 (N_21899,N_19659,N_21244);
xor U21900 (N_21900,N_19034,N_20378);
nor U21901 (N_21901,N_21118,N_18765);
and U21902 (N_21902,N_19514,N_19180);
nor U21903 (N_21903,N_21327,N_20844);
nor U21904 (N_21904,N_19317,N_18916);
nand U21905 (N_21905,N_21376,N_20191);
nand U21906 (N_21906,N_20482,N_19565);
or U21907 (N_21907,N_20505,N_19432);
nand U21908 (N_21908,N_21325,N_20170);
nor U21909 (N_21909,N_20678,N_20897);
nand U21910 (N_21910,N_19971,N_19160);
xor U21911 (N_21911,N_19304,N_21765);
xnor U21912 (N_21912,N_20298,N_19545);
xor U21913 (N_21913,N_18782,N_19581);
or U21914 (N_21914,N_20315,N_19610);
or U21915 (N_21915,N_21767,N_21056);
and U21916 (N_21916,N_18810,N_20028);
nand U21917 (N_21917,N_20265,N_19936);
nand U21918 (N_21918,N_20091,N_18880);
or U21919 (N_21919,N_20421,N_21704);
xnor U21920 (N_21920,N_21324,N_21441);
or U21921 (N_21921,N_20805,N_21861);
nand U21922 (N_21922,N_19353,N_19567);
nor U21923 (N_21923,N_20003,N_20051);
nand U21924 (N_21924,N_21811,N_18942);
or U21925 (N_21925,N_20526,N_20107);
or U21926 (N_21926,N_19957,N_21461);
nand U21927 (N_21927,N_21845,N_19910);
nand U21928 (N_21928,N_20738,N_19743);
or U21929 (N_21929,N_19934,N_19916);
and U21930 (N_21930,N_18973,N_21731);
nor U21931 (N_21931,N_21402,N_21781);
nand U21932 (N_21932,N_19645,N_21107);
and U21933 (N_21933,N_19885,N_20679);
or U21934 (N_21934,N_19541,N_20979);
nor U21935 (N_21935,N_20751,N_20692);
or U21936 (N_21936,N_20046,N_20318);
and U21937 (N_21937,N_19284,N_20153);
and U21938 (N_21938,N_20174,N_20572);
and U21939 (N_21939,N_21361,N_19720);
nor U21940 (N_21940,N_19462,N_19446);
or U21941 (N_21941,N_21028,N_20409);
and U21942 (N_21942,N_20986,N_21026);
and U21943 (N_21943,N_18900,N_19516);
nand U21944 (N_21944,N_20030,N_19879);
xor U21945 (N_21945,N_21084,N_21592);
xnor U21946 (N_21946,N_19112,N_20527);
or U21947 (N_21947,N_20748,N_21014);
or U21948 (N_21948,N_20529,N_19238);
or U21949 (N_21949,N_21387,N_18998);
nand U21950 (N_21950,N_20617,N_19901);
xnor U21951 (N_21951,N_19853,N_19595);
nand U21952 (N_21952,N_19786,N_20079);
and U21953 (N_21953,N_20918,N_21718);
and U21954 (N_21954,N_19488,N_18848);
nor U21955 (N_21955,N_20896,N_20402);
xnor U21956 (N_21956,N_21011,N_21155);
and U21957 (N_21957,N_19893,N_20311);
nand U21958 (N_21958,N_21591,N_21309);
nand U21959 (N_21959,N_21379,N_18953);
nor U21960 (N_21960,N_19725,N_19792);
xnor U21961 (N_21961,N_19810,N_20476);
nor U21962 (N_21962,N_20664,N_21572);
xnor U21963 (N_21963,N_21810,N_20207);
nand U21964 (N_21964,N_21775,N_20250);
and U21965 (N_21965,N_19240,N_20743);
xor U21966 (N_21966,N_20014,N_19998);
and U21967 (N_21967,N_20539,N_21405);
nor U21968 (N_21968,N_19865,N_18834);
or U21969 (N_21969,N_21157,N_21142);
xnor U21970 (N_21970,N_21460,N_19115);
and U21971 (N_21971,N_20627,N_19182);
xnor U21972 (N_21972,N_19144,N_19781);
nand U21973 (N_21973,N_21007,N_20256);
xor U21974 (N_21974,N_21131,N_20070);
xnor U21975 (N_21975,N_21308,N_18873);
nand U21976 (N_21976,N_20123,N_18752);
or U21977 (N_21977,N_20460,N_20078);
and U21978 (N_21978,N_19146,N_20632);
nand U21979 (N_21979,N_19760,N_19278);
xnor U21980 (N_21980,N_19806,N_20506);
xnor U21981 (N_21981,N_19883,N_18972);
nand U21982 (N_21982,N_19305,N_21147);
nor U21983 (N_21983,N_19871,N_19218);
and U21984 (N_21984,N_20510,N_20034);
or U21985 (N_21985,N_19797,N_20371);
nor U21986 (N_21986,N_21380,N_19308);
and U21987 (N_21987,N_21796,N_19033);
nand U21988 (N_21988,N_20455,N_20905);
and U21989 (N_21989,N_21478,N_20596);
and U21990 (N_21990,N_18828,N_21676);
or U21991 (N_21991,N_19417,N_21373);
xor U21992 (N_21992,N_19007,N_21040);
and U21993 (N_21993,N_19440,N_20874);
xnor U21994 (N_21994,N_21366,N_18960);
or U21995 (N_21995,N_20124,N_19126);
nor U21996 (N_21996,N_20445,N_19461);
nand U21997 (N_21997,N_19912,N_19987);
xnor U21998 (N_21998,N_20837,N_19326);
or U21999 (N_21999,N_20521,N_20876);
nor U22000 (N_22000,N_21108,N_18915);
xnor U22001 (N_22001,N_18909,N_21162);
nand U22002 (N_22002,N_21567,N_21522);
nand U22003 (N_22003,N_20493,N_21024);
xnor U22004 (N_22004,N_19949,N_18894);
or U22005 (N_22005,N_19964,N_19966);
nor U22006 (N_22006,N_21078,N_19074);
nand U22007 (N_22007,N_18977,N_21643);
xor U22008 (N_22008,N_19108,N_19418);
nor U22009 (N_22009,N_20220,N_19481);
or U22010 (N_22010,N_21849,N_20291);
xor U22011 (N_22011,N_19489,N_20397);
xnor U22012 (N_22012,N_21653,N_21214);
or U22013 (N_22013,N_20806,N_20308);
xnor U22014 (N_22014,N_21289,N_20940);
xor U22015 (N_22015,N_19832,N_20607);
nand U22016 (N_22016,N_21495,N_18844);
or U22017 (N_22017,N_19153,N_19260);
and U22018 (N_22018,N_20763,N_18927);
nor U22019 (N_22019,N_20525,N_21374);
nand U22020 (N_22020,N_21805,N_19321);
nor U22021 (N_22021,N_21648,N_18947);
nor U22022 (N_22022,N_20077,N_19377);
nor U22023 (N_22023,N_21426,N_20713);
and U22024 (N_22024,N_18776,N_20148);
nor U22025 (N_22025,N_21196,N_20417);
nor U22026 (N_22026,N_20152,N_19731);
or U22027 (N_22027,N_20249,N_19371);
xor U22028 (N_22028,N_20057,N_19570);
and U22029 (N_22029,N_19322,N_20788);
xor U22030 (N_22030,N_21552,N_18911);
and U22031 (N_22031,N_19614,N_19709);
nand U22032 (N_22032,N_18903,N_18962);
xor U22033 (N_22033,N_19038,N_19136);
or U22034 (N_22034,N_19911,N_19137);
xor U22035 (N_22035,N_19161,N_20932);
xor U22036 (N_22036,N_20559,N_20089);
nor U22037 (N_22037,N_21473,N_20669);
nand U22038 (N_22038,N_21663,N_20629);
or U22039 (N_22039,N_19081,N_19085);
xnor U22040 (N_22040,N_18847,N_21021);
or U22041 (N_22041,N_20056,N_20228);
nand U22042 (N_22042,N_19564,N_21139);
nand U22043 (N_22043,N_20229,N_19517);
and U22044 (N_22044,N_19424,N_21239);
nand U22045 (N_22045,N_21492,N_21513);
nand U22046 (N_22046,N_20992,N_19644);
nand U22047 (N_22047,N_20670,N_20446);
or U22048 (N_22048,N_20840,N_19704);
xnor U22049 (N_22049,N_19458,N_19044);
and U22050 (N_22050,N_21317,N_21785);
nor U22051 (N_22051,N_21408,N_21415);
xor U22052 (N_22052,N_21077,N_20216);
xnor U22053 (N_22053,N_18816,N_21560);
nand U22054 (N_22054,N_19140,N_20535);
and U22055 (N_22055,N_20296,N_19403);
or U22056 (N_22056,N_19301,N_18943);
xnor U22057 (N_22057,N_19199,N_20496);
nand U22058 (N_22058,N_20821,N_19896);
or U22059 (N_22059,N_18805,N_20923);
nand U22060 (N_22060,N_20930,N_21311);
nor U22061 (N_22061,N_20646,N_18822);
xor U22062 (N_22062,N_19362,N_19863);
or U22063 (N_22063,N_19422,N_18845);
or U22064 (N_22064,N_19054,N_20066);
xnor U22065 (N_22065,N_21550,N_19356);
and U22066 (N_22066,N_20978,N_20400);
xor U22067 (N_22067,N_19174,N_21207);
xor U22068 (N_22068,N_20049,N_19525);
xor U22069 (N_22069,N_20954,N_19550);
or U22070 (N_22070,N_19017,N_19110);
nand U22071 (N_22071,N_19549,N_19454);
or U22072 (N_22072,N_19537,N_18898);
xnor U22073 (N_22073,N_19601,N_20106);
xnor U22074 (N_22074,N_19120,N_20803);
nor U22075 (N_22075,N_18882,N_21458);
xor U22076 (N_22076,N_18974,N_21534);
nor U22077 (N_22077,N_20804,N_21568);
and U22078 (N_22078,N_19181,N_20414);
and U22079 (N_22079,N_19124,N_20094);
nor U22080 (N_22080,N_19821,N_20882);
nand U22081 (N_22081,N_18854,N_20656);
xnor U22082 (N_22082,N_20531,N_20942);
nor U22083 (N_22083,N_21123,N_20736);
nand U22084 (N_22084,N_18952,N_19306);
nor U22085 (N_22085,N_21870,N_20739);
and U22086 (N_22086,N_21679,N_20586);
xnor U22087 (N_22087,N_19960,N_19862);
nand U22088 (N_22088,N_20474,N_21628);
and U22089 (N_22089,N_20029,N_21271);
or U22090 (N_22090,N_19176,N_18946);
xor U22091 (N_22091,N_21755,N_21843);
xnor U22092 (N_22092,N_19974,N_19900);
nand U22093 (N_22093,N_20000,N_21520);
nand U22094 (N_22094,N_21614,N_19063);
and U22095 (N_22095,N_19560,N_21430);
nor U22096 (N_22096,N_20305,N_19012);
or U22097 (N_22097,N_18867,N_19193);
nand U22098 (N_22098,N_21396,N_20420);
or U22099 (N_22099,N_19930,N_21146);
xor U22100 (N_22100,N_21215,N_19309);
nand U22101 (N_22101,N_19069,N_21283);
nor U22102 (N_22102,N_20558,N_19277);
xor U22103 (N_22103,N_21697,N_21708);
nor U22104 (N_22104,N_20784,N_21322);
and U22105 (N_22105,N_21867,N_19706);
nand U22106 (N_22106,N_20587,N_18928);
xor U22107 (N_22107,N_20828,N_21585);
nor U22108 (N_22108,N_19090,N_19848);
nor U22109 (N_22109,N_21316,N_21536);
nor U22110 (N_22110,N_19303,N_20582);
nor U22111 (N_22111,N_19808,N_19060);
xor U22112 (N_22112,N_20197,N_21348);
or U22113 (N_22113,N_19285,N_18931);
nor U22114 (N_22114,N_20624,N_18986);
xor U22115 (N_22115,N_21093,N_18933);
xor U22116 (N_22116,N_18887,N_19803);
xor U22117 (N_22117,N_21281,N_21677);
or U22118 (N_22118,N_19433,N_18951);
nor U22119 (N_22119,N_19932,N_20480);
nand U22120 (N_22120,N_21245,N_19876);
xnor U22121 (N_22121,N_18879,N_21280);
nor U22122 (N_22122,N_19700,N_21449);
xnor U22123 (N_22123,N_20618,N_20353);
nand U22124 (N_22124,N_21641,N_21795);
and U22125 (N_22125,N_20548,N_20479);
or U22126 (N_22126,N_20184,N_19057);
nand U22127 (N_22127,N_20257,N_19102);
nor U22128 (N_22128,N_19449,N_19342);
and U22129 (N_22129,N_21241,N_21259);
or U22130 (N_22130,N_21313,N_20035);
or U22131 (N_22131,N_21599,N_20113);
xor U22132 (N_22132,N_19854,N_21303);
nand U22133 (N_22133,N_21206,N_19336);
or U22134 (N_22134,N_19639,N_20753);
nand U22135 (N_22135,N_20040,N_21032);
nor U22136 (N_22136,N_20895,N_19401);
or U22137 (N_22137,N_19859,N_20227);
nand U22138 (N_22138,N_19620,N_21012);
nor U22139 (N_22139,N_19021,N_20438);
nor U22140 (N_22140,N_19948,N_20909);
nand U22141 (N_22141,N_19684,N_21295);
nor U22142 (N_22142,N_21638,N_21821);
nand U22143 (N_22143,N_21530,N_19767);
nand U22144 (N_22144,N_18890,N_19100);
or U22145 (N_22145,N_19697,N_20551);
and U22146 (N_22146,N_20450,N_20999);
nor U22147 (N_22147,N_20765,N_19997);
nor U22148 (N_22148,N_21595,N_21545);
and U22149 (N_22149,N_19339,N_21858);
nor U22150 (N_22150,N_19654,N_18792);
xor U22151 (N_22151,N_21645,N_21230);
xnor U22152 (N_22152,N_19650,N_18839);
nor U22153 (N_22153,N_21386,N_18888);
nand U22154 (N_22154,N_20533,N_19105);
or U22155 (N_22155,N_21326,N_19250);
nor U22156 (N_22156,N_19927,N_20443);
nand U22157 (N_22157,N_20393,N_19472);
xor U22158 (N_22158,N_21001,N_19191);
and U22159 (N_22159,N_19492,N_19029);
and U22160 (N_22160,N_20498,N_18851);
or U22161 (N_22161,N_20372,N_20958);
nand U22162 (N_22162,N_21496,N_21231);
nor U22163 (N_22163,N_20473,N_19275);
and U22164 (N_22164,N_20890,N_21787);
nand U22165 (N_22165,N_19925,N_19217);
or U22166 (N_22166,N_20033,N_18785);
or U22167 (N_22167,N_21400,N_20797);
xnor U22168 (N_22168,N_19080,N_21276);
xor U22169 (N_22169,N_21434,N_20201);
or U22170 (N_22170,N_21487,N_20866);
and U22171 (N_22171,N_21174,N_18862);
and U22172 (N_22172,N_19690,N_19861);
or U22173 (N_22173,N_21356,N_20108);
xnor U22174 (N_22174,N_19372,N_21068);
nand U22175 (N_22175,N_19696,N_19387);
nand U22176 (N_22176,N_19826,N_18773);
and U22177 (N_22177,N_20910,N_21031);
nand U22178 (N_22178,N_21249,N_20854);
and U22179 (N_22179,N_21516,N_20781);
nand U22180 (N_22180,N_20831,N_19055);
xnor U22181 (N_22181,N_21654,N_20764);
nor U22182 (N_22182,N_20603,N_19754);
and U22183 (N_22183,N_20605,N_19621);
xor U22184 (N_22184,N_19018,N_19635);
nand U22185 (N_22185,N_19167,N_19702);
and U22186 (N_22186,N_20973,N_19116);
nor U22187 (N_22187,N_19122,N_20219);
nand U22188 (N_22188,N_20137,N_19224);
and U22189 (N_22189,N_20246,N_20967);
or U22190 (N_22190,N_20024,N_19628);
xnor U22191 (N_22191,N_21442,N_21529);
xnor U22192 (N_22192,N_19678,N_18902);
nor U22193 (N_22193,N_18863,N_21871);
nor U22194 (N_22194,N_21110,N_20281);
xnor U22195 (N_22195,N_19302,N_21204);
nor U22196 (N_22196,N_19508,N_20584);
or U22197 (N_22197,N_19269,N_20855);
xor U22198 (N_22198,N_21699,N_21847);
nand U22199 (N_22199,N_18945,N_20331);
nor U22200 (N_22200,N_20136,N_19198);
or U22201 (N_22201,N_19824,N_20109);
xor U22202 (N_22202,N_21144,N_20016);
and U22203 (N_22203,N_20364,N_18774);
and U22204 (N_22204,N_20815,N_20340);
and U22205 (N_22205,N_20581,N_19358);
or U22206 (N_22206,N_21687,N_21286);
and U22207 (N_22207,N_21830,N_20841);
and U22208 (N_22208,N_19231,N_21824);
xnor U22209 (N_22209,N_19364,N_19248);
nand U22210 (N_22210,N_21265,N_19970);
or U22211 (N_22211,N_18840,N_20208);
nor U22212 (N_22212,N_21344,N_19216);
and U22213 (N_22213,N_19359,N_18788);
or U22214 (N_22214,N_21800,N_18905);
nand U22215 (N_22215,N_21055,N_21323);
nor U22216 (N_22216,N_20122,N_19068);
and U22217 (N_22217,N_19800,N_20367);
nor U22218 (N_22218,N_18874,N_21476);
and U22219 (N_22219,N_21855,N_19898);
or U22220 (N_22220,N_19150,N_19577);
or U22221 (N_22221,N_18913,N_19815);
nand U22222 (N_22222,N_19145,N_20933);
xnor U22223 (N_22223,N_19933,N_18907);
nand U22224 (N_22224,N_21127,N_20687);
nand U22225 (N_22225,N_20159,N_21119);
xnor U22226 (N_22226,N_19207,N_19943);
and U22227 (N_22227,N_18976,N_18783);
or U22228 (N_22228,N_21583,N_19171);
nand U22229 (N_22229,N_21034,N_20299);
nor U22230 (N_22230,N_20647,N_20620);
nand U22231 (N_22231,N_21571,N_19147);
or U22232 (N_22232,N_21189,N_19773);
nor U22233 (N_22233,N_21691,N_20156);
nor U22234 (N_22234,N_19544,N_20466);
xor U22235 (N_22235,N_20488,N_20719);
nor U22236 (N_22236,N_21412,N_19744);
or U22237 (N_22237,N_20520,N_21822);
nor U22238 (N_22238,N_20503,N_20494);
and U22239 (N_22239,N_19811,N_19954);
or U22240 (N_22240,N_20935,N_20931);
nand U22241 (N_22241,N_20566,N_19453);
nor U22242 (N_22242,N_20255,N_20358);
and U22243 (N_22243,N_19431,N_19683);
nand U22244 (N_22244,N_20245,N_21723);
and U22245 (N_22245,N_19009,N_21357);
xor U22246 (N_22246,N_19399,N_19427);
nand U22247 (N_22247,N_19232,N_21616);
xor U22248 (N_22248,N_19204,N_19434);
nand U22249 (N_22249,N_21334,N_21193);
nand U22250 (N_22250,N_20852,N_20274);
and U22251 (N_22251,N_19348,N_20823);
nor U22252 (N_22252,N_20084,N_20131);
nor U22253 (N_22253,N_21355,N_21705);
nand U22254 (N_22254,N_20872,N_18922);
xnor U22255 (N_22255,N_19681,N_21082);
xnor U22256 (N_22256,N_19527,N_18884);
and U22257 (N_22257,N_20723,N_18883);
or U22258 (N_22258,N_19676,N_21419);
xor U22259 (N_22259,N_19822,N_19737);
nand U22260 (N_22260,N_18889,N_20115);
or U22261 (N_22261,N_19783,N_21675);
nor U22262 (N_22262,N_21427,N_20427);
nand U22263 (N_22263,N_20222,N_21042);
nor U22264 (N_22264,N_19178,N_19503);
nand U22265 (N_22265,N_19627,N_21741);
nor U22266 (N_22266,N_20063,N_19314);
xnor U22267 (N_22267,N_20168,N_21126);
nand U22268 (N_22268,N_19734,N_20811);
xor U22269 (N_22269,N_20059,N_21825);
and U22270 (N_22270,N_21840,N_20707);
and U22271 (N_22271,N_20114,N_19523);
nor U22272 (N_22272,N_21485,N_21254);
nor U22273 (N_22273,N_19318,N_20902);
and U22274 (N_22274,N_20983,N_21300);
and U22275 (N_22275,N_20894,N_19469);
nor U22276 (N_22276,N_20018,N_20199);
or U22277 (N_22277,N_19867,N_20720);
nor U22278 (N_22278,N_20356,N_19498);
nand U22279 (N_22279,N_20212,N_19035);
nor U22280 (N_22280,N_20619,N_19518);
and U22281 (N_22281,N_20477,N_19740);
and U22282 (N_22282,N_21857,N_19226);
xor U22283 (N_22283,N_18823,N_19311);
nor U22284 (N_22284,N_19125,N_21816);
nor U22285 (N_22285,N_21175,N_19874);
xnor U22286 (N_22286,N_19222,N_19886);
or U22287 (N_22287,N_21158,N_21820);
or U22288 (N_22288,N_19575,N_21062);
nor U22289 (N_22289,N_19988,N_21694);
or U22290 (N_22290,N_21505,N_20075);
and U22291 (N_22291,N_21526,N_19675);
nor U22292 (N_22292,N_21216,N_21610);
xnor U22293 (N_22293,N_20908,N_19816);
nor U22294 (N_22294,N_20175,N_18793);
or U22295 (N_22295,N_19955,N_21632);
nand U22296 (N_22296,N_18861,N_19631);
xnor U22297 (N_22297,N_20297,N_19649);
nand U22298 (N_22298,N_19297,N_21532);
nand U22299 (N_22299,N_21198,N_20458);
xnor U22300 (N_22300,N_20283,N_20074);
xor U22301 (N_22301,N_20667,N_19784);
xor U22302 (N_22302,N_20634,N_20638);
nor U22303 (N_22303,N_20337,N_21002);
nor U22304 (N_22304,N_20190,N_21392);
xor U22305 (N_22305,N_18864,N_20915);
nand U22306 (N_22306,N_20759,N_19374);
nand U22307 (N_22307,N_20594,N_20453);
nor U22308 (N_22308,N_21088,N_19945);
or U22309 (N_22309,N_19633,N_20573);
and U22310 (N_22310,N_20547,N_21575);
nand U22311 (N_22311,N_19761,N_20792);
xor U22312 (N_22312,N_19989,N_19239);
xnor U22313 (N_22313,N_18771,N_19764);
xor U22314 (N_22314,N_18770,N_20317);
nand U22315 (N_22315,N_20247,N_21185);
and U22316 (N_22316,N_21834,N_20047);
or U22317 (N_22317,N_21659,N_21517);
and U22318 (N_22318,N_19465,N_21145);
nand U22319 (N_22319,N_19726,N_20376);
nand U22320 (N_22320,N_20399,N_20972);
nand U22321 (N_22321,N_20889,N_19027);
xnor U22322 (N_22322,N_20912,N_20981);
xnor U22323 (N_22323,N_19512,N_19736);
nor U22324 (N_22324,N_21804,N_20668);
or U22325 (N_22325,N_20685,N_19258);
nor U22326 (N_22326,N_20770,N_21424);
nor U22327 (N_22327,N_18997,N_20484);
nor U22328 (N_22328,N_18969,N_19665);
or U22329 (N_22329,N_20746,N_21510);
nor U22330 (N_22330,N_19707,N_19190);
nand U22331 (N_22331,N_20943,N_20509);
xnor U22332 (N_22332,N_19682,N_20927);
and U22333 (N_22333,N_20637,N_20171);
and U22334 (N_22334,N_20887,N_21046);
xor U22335 (N_22335,N_21406,N_20883);
nand U22336 (N_22336,N_18767,N_21543);
nor U22337 (N_22337,N_20072,N_19864);
or U22338 (N_22338,N_20644,N_21578);
nor U22339 (N_22339,N_20740,N_18875);
nor U22340 (N_22340,N_20665,N_20717);
xor U22341 (N_22341,N_21394,N_21171);
or U22342 (N_22342,N_20266,N_20657);
and U22343 (N_22343,N_20666,N_19128);
nand U22344 (N_22344,N_19331,N_21742);
or U22345 (N_22345,N_20556,N_19748);
nor U22346 (N_22346,N_21627,N_19630);
or U22347 (N_22347,N_21365,N_19907);
and U22348 (N_22348,N_20608,N_19172);
or U22349 (N_22349,N_20756,N_21714);
xnor U22350 (N_22350,N_19780,N_19014);
nor U22351 (N_22351,N_19251,N_21090);
and U22352 (N_22352,N_21160,N_19652);
or U22353 (N_22353,N_18996,N_20676);
nor U22354 (N_22354,N_20833,N_21038);
or U22355 (N_22355,N_20893,N_21268);
nand U22356 (N_22356,N_19230,N_19598);
or U22357 (N_22357,N_21393,N_21403);
nor U22358 (N_22358,N_19114,N_19478);
or U22359 (N_22359,N_21459,N_20497);
nand U22360 (N_22360,N_20236,N_20185);
and U22361 (N_22361,N_21306,N_19552);
nor U22362 (N_22362,N_20082,N_19051);
nor U22363 (N_22363,N_20877,N_19490);
nor U22364 (N_22364,N_19011,N_20585);
nand U22365 (N_22365,N_19670,N_20456);
nand U22366 (N_22366,N_20195,N_19892);
and U22367 (N_22367,N_19227,N_20442);
nand U22368 (N_22368,N_21263,N_20758);
or U22369 (N_22369,N_20861,N_19276);
or U22370 (N_22370,N_20544,N_21416);
xnor U22371 (N_22371,N_19839,N_19390);
or U22372 (N_22372,N_21688,N_19903);
or U22373 (N_22373,N_21321,N_21115);
or U22374 (N_22374,N_21190,N_21363);
nor U22375 (N_22375,N_20528,N_21582);
or U22376 (N_22376,N_20574,N_19264);
nand U22377 (N_22377,N_20277,N_19976);
or U22378 (N_22378,N_21130,N_20892);
nand U22379 (N_22379,N_19255,N_21183);
and U22380 (N_22380,N_20832,N_21869);
nand U22381 (N_22381,N_18784,N_19759);
xnor U22382 (N_22382,N_19653,N_19118);
and U22383 (N_22383,N_21342,N_21735);
or U22384 (N_22384,N_21260,N_21229);
nor U22385 (N_22385,N_21170,N_20917);
and U22386 (N_22386,N_21512,N_19531);
and U22387 (N_22387,N_19438,N_20926);
nand U22388 (N_22388,N_19695,N_21669);
or U22389 (N_22389,N_20853,N_19787);
or U22390 (N_22390,N_20110,N_20052);
and U22391 (N_22391,N_19320,N_21188);
nand U22392 (N_22392,N_21161,N_19777);
xnor U22393 (N_22393,N_20313,N_20188);
or U22394 (N_22394,N_19920,N_21091);
or U22395 (N_22395,N_20278,N_21726);
and U22396 (N_22396,N_21750,N_21634);
or U22397 (N_22397,N_20776,N_21644);
and U22398 (N_22398,N_21745,N_21018);
and U22399 (N_22399,N_21338,N_21555);
and U22400 (N_22400,N_18981,N_18849);
and U22401 (N_22401,N_20752,N_21725);
or U22402 (N_22402,N_20880,N_21646);
nor U22403 (N_22403,N_18855,N_19495);
nor U22404 (N_22404,N_19506,N_20773);
xor U22405 (N_22405,N_20939,N_21747);
nand U22406 (N_22406,N_18830,N_19154);
nand U22407 (N_22407,N_19804,N_21409);
xor U22408 (N_22408,N_20677,N_21828);
xor U22409 (N_22409,N_19299,N_19429);
and U22410 (N_22410,N_20189,N_19166);
nor U22411 (N_22411,N_21404,N_19919);
xor U22412 (N_22412,N_21036,N_19395);
nand U22413 (N_22413,N_21457,N_20426);
and U22414 (N_22414,N_19421,N_19106);
and U22415 (N_22415,N_20839,N_19435);
nor U22416 (N_22416,N_19600,N_19235);
xor U22417 (N_22417,N_21279,N_21116);
or U22418 (N_22418,N_21594,N_19753);
or U22419 (N_22419,N_21794,N_19420);
nand U22420 (N_22420,N_19705,N_19662);
and U22421 (N_22421,N_20215,N_20293);
and U22422 (N_22422,N_19613,N_21255);
or U22423 (N_22423,N_20243,N_20478);
and U22424 (N_22424,N_19163,N_19423);
or U22425 (N_22425,N_20911,N_19894);
xor U22426 (N_22426,N_20459,N_19938);
or U22427 (N_22427,N_20700,N_19292);
xnor U22428 (N_22428,N_20641,N_21807);
nand U22429 (N_22429,N_21191,N_21452);
or U22430 (N_22430,N_19629,N_20718);
and U22431 (N_22431,N_19830,N_21769);
nand U22432 (N_22432,N_18781,N_18842);
xnor U22433 (N_22433,N_20702,N_20938);
nand U22434 (N_22434,N_21464,N_19170);
nand U22435 (N_22435,N_21003,N_20963);
nor U22436 (N_22436,N_20119,N_19738);
or U22437 (N_22437,N_20095,N_20541);
nor U22438 (N_22438,N_20203,N_21851);
and U22439 (N_22439,N_21589,N_21749);
nor U22440 (N_22440,N_19319,N_19836);
nand U22441 (N_22441,N_18935,N_20651);
nor U22442 (N_22442,N_19827,N_19749);
xnor U22443 (N_22443,N_19158,N_18841);
xor U22444 (N_22444,N_21390,N_19094);
nor U22445 (N_22445,N_21226,N_21238);
nand U22446 (N_22446,N_21506,N_21744);
nand U22447 (N_22447,N_21753,N_20069);
or U22448 (N_22448,N_21444,N_18868);
nor U22449 (N_22449,N_20373,N_18899);
xnor U22450 (N_22450,N_18800,N_19796);
nand U22451 (N_22451,N_21192,N_19298);
or U22452 (N_22452,N_19468,N_21823);
nand U22453 (N_22453,N_19052,N_19286);
nand U22454 (N_22454,N_21391,N_20611);
or U22455 (N_22455,N_20578,N_19623);
and U22456 (N_22456,N_20303,N_21069);
nand U22457 (N_22457,N_19316,N_20816);
nor U22458 (N_22458,N_20636,N_20012);
or U22459 (N_22459,N_20253,N_19323);
and U22460 (N_22460,N_18757,N_21278);
nand U22461 (N_22461,N_21719,N_19817);
xnor U22462 (N_22462,N_20642,N_19741);
nand U22463 (N_22463,N_21015,N_20829);
nor U22464 (N_22464,N_20725,N_19099);
or U22465 (N_22465,N_19135,N_21509);
nor U22466 (N_22466,N_21853,N_19263);
nor U22467 (N_22467,N_18756,N_18989);
xor U22468 (N_22468,N_21601,N_19370);
and U22469 (N_22469,N_20783,N_20457);
nand U22470 (N_22470,N_21773,N_20928);
and U22471 (N_22471,N_20058,N_20920);
xor U22472 (N_22472,N_21339,N_21329);
or U22473 (N_22473,N_20270,N_20276);
and U22474 (N_22474,N_20922,N_19015);
xnor U22475 (N_22475,N_21681,N_20157);
nor U22476 (N_22476,N_20698,N_19315);
xor U22477 (N_22477,N_20098,N_21647);
nand U22478 (N_22478,N_19984,N_21331);
or U22479 (N_22479,N_20731,N_19189);
xnor U22480 (N_22480,N_20937,N_21554);
or U22481 (N_22481,N_19041,N_19719);
and U22482 (N_22482,N_20583,N_20126);
or U22483 (N_22483,N_20511,N_21657);
nor U22484 (N_22484,N_21163,N_19165);
xnor U22485 (N_22485,N_19742,N_21598);
nand U22486 (N_22486,N_20538,N_20512);
nor U22487 (N_22487,N_21482,N_21087);
nand U22488 (N_22488,N_21528,N_18866);
xor U22489 (N_22489,N_18937,N_21557);
and U22490 (N_22490,N_19294,N_20690);
nor U22491 (N_22491,N_21730,N_21236);
or U22492 (N_22492,N_20779,N_19244);
xnor U22493 (N_22493,N_19716,N_20310);
nor U22494 (N_22494,N_21490,N_21101);
and U22495 (N_22495,N_20501,N_19795);
nor U22496 (N_22496,N_21122,N_20716);
nor U22497 (N_22497,N_20294,N_21564);
xor U22498 (N_22498,N_20234,N_20172);
nor U22499 (N_22499,N_20434,N_19194);
and U22500 (N_22500,N_20160,N_20086);
and U22501 (N_22501,N_19888,N_21692);
xor U22502 (N_22502,N_19849,N_21410);
nand U22503 (N_22503,N_19829,N_20169);
and U22504 (N_22504,N_20344,N_19333);
and U22505 (N_22505,N_20683,N_19123);
nand U22506 (N_22506,N_19929,N_20848);
nor U22507 (N_22507,N_21341,N_20817);
or U22508 (N_22508,N_20118,N_21418);
and U22509 (N_22509,N_19405,N_21227);
xor U22510 (N_22510,N_19604,N_20004);
nand U22511 (N_22511,N_21508,N_18966);
xor U22512 (N_22512,N_18865,N_19177);
and U22513 (N_22513,N_18819,N_20360);
nand U22514 (N_22514,N_18790,N_18924);
xor U22515 (N_22515,N_19247,N_20843);
or U22516 (N_22516,N_19113,N_20514);
or U22517 (N_22517,N_18769,N_21079);
xnor U22518 (N_22518,N_19307,N_19612);
or U22519 (N_22519,N_21706,N_20490);
nor U22520 (N_22520,N_20518,N_21129);
or U22521 (N_22521,N_21786,N_21631);
xnor U22522 (N_22522,N_19024,N_21609);
nor U22523 (N_22523,N_20810,N_18808);
or U22524 (N_22524,N_18768,N_20742);
and U22525 (N_22525,N_18797,N_18970);
and U22526 (N_22526,N_20674,N_19407);
and U22527 (N_22527,N_21337,N_19259);
nor U22528 (N_22528,N_21792,N_19437);
nand U22529 (N_22529,N_19533,N_20794);
and U22530 (N_22530,N_19775,N_20363);
nor U22531 (N_22531,N_20885,N_21104);
nand U22532 (N_22532,N_20320,N_18815);
nor U22533 (N_22533,N_20771,N_18925);
nand U22534 (N_22534,N_20708,N_21044);
or U22535 (N_22535,N_18881,N_20565);
and U22536 (N_22536,N_20575,N_19608);
nor U22537 (N_22537,N_21738,N_21121);
xor U22538 (N_22538,N_19799,N_20862);
and U22539 (N_22539,N_20158,N_19048);
or U22540 (N_22540,N_21698,N_20231);
and U22541 (N_22541,N_20233,N_20134);
or U22542 (N_22542,N_20093,N_19562);
or U22543 (N_22543,N_19188,N_21025);
nor U22544 (N_22544,N_19026,N_19831);
nor U22545 (N_22545,N_20863,N_20648);
xor U22546 (N_22546,N_18971,N_21071);
or U22547 (N_22547,N_19755,N_18763);
xor U22548 (N_22548,N_21030,N_20609);
nand U22549 (N_22549,N_21383,N_21081);
xnor U22550 (N_22550,N_20374,N_20235);
or U22551 (N_22551,N_21397,N_20869);
nor U22552 (N_22552,N_21600,N_20284);
xor U22553 (N_22553,N_19522,N_20261);
or U22554 (N_22554,N_21291,N_19366);
nand U22555 (N_22555,N_21752,N_20254);
nand U22556 (N_22556,N_19819,N_18878);
xnor U22557 (N_22557,N_19617,N_21095);
nor U22558 (N_22558,N_20873,N_21751);
nor U22559 (N_22559,N_20264,N_20849);
and U22560 (N_22560,N_20330,N_19393);
or U22561 (N_22561,N_19891,N_19246);
xnor U22562 (N_22562,N_20431,N_19658);
xnor U22563 (N_22563,N_18950,N_20166);
nor U22564 (N_22564,N_19774,N_19291);
or U22565 (N_22565,N_18965,N_18772);
nor U22566 (N_22566,N_20329,N_20422);
or U22567 (N_22567,N_21045,N_20306);
and U22568 (N_22568,N_19037,N_20335);
or U22569 (N_22569,N_20562,N_20085);
xnor U22570 (N_22570,N_21448,N_19837);
and U22571 (N_22571,N_19445,N_21862);
nand U22572 (N_22572,N_20673,N_21848);
or U22573 (N_22573,N_20697,N_19935);
xor U22574 (N_22574,N_20011,N_19219);
or U22575 (N_22575,N_19312,N_20424);
xor U22576 (N_22576,N_19396,N_21551);
or U22577 (N_22577,N_20998,N_21491);
nand U22578 (N_22578,N_19368,N_19557);
nor U22579 (N_22579,N_20796,N_19426);
nor U22580 (N_22580,N_20662,N_21721);
xor U22581 (N_22581,N_21051,N_21479);
and U22582 (N_22582,N_18939,N_19584);
xor U22583 (N_22583,N_18985,N_21340);
and U22584 (N_22584,N_19484,N_21558);
and U22585 (N_22585,N_20023,N_20639);
xnor U22586 (N_22586,N_21399,N_19553);
and U22587 (N_22587,N_20508,N_21009);
and U22588 (N_22588,N_20630,N_18838);
xor U22589 (N_22589,N_20947,N_21436);
or U22590 (N_22590,N_19568,N_21273);
nand U22591 (N_22591,N_20454,N_20615);
nand U22592 (N_22592,N_21136,N_20121);
xor U22593 (N_22593,N_21250,N_19959);
and U22594 (N_22594,N_19963,N_19625);
or U22595 (N_22595,N_20513,N_19618);
xnor U22596 (N_22596,N_21760,N_21282);
nand U22597 (N_22597,N_19391,N_19020);
nor U22598 (N_22598,N_20307,N_18779);
nor U22599 (N_22599,N_19729,N_19882);
nor U22600 (N_22600,N_21177,N_18967);
xor U22601 (N_22601,N_21728,N_21378);
and U22602 (N_22602,N_19386,N_20621);
nand U22603 (N_22603,N_19556,N_21468);
nor U22604 (N_22604,N_21307,N_21076);
nor U22605 (N_22605,N_20950,N_21208);
nor U22606 (N_22606,N_21748,N_20301);
and U22607 (N_22607,N_20903,N_21700);
and U22608 (N_22608,N_19511,N_19179);
xnor U22609 (N_22609,N_18803,N_19646);
nand U22610 (N_22610,N_21237,N_20543);
nand U22611 (N_22611,N_20139,N_19637);
nand U22612 (N_22612,N_19300,N_19467);
xor U22613 (N_22613,N_21580,N_20415);
nand U22614 (N_22614,N_21854,N_21054);
or U22615 (N_22615,N_20799,N_20081);
or U22616 (N_22616,N_19352,N_19609);
or U22617 (N_22617,N_18814,N_21381);
and U22618 (N_22618,N_18801,N_21305);
nand U22619 (N_22619,N_18835,N_21080);
nand U22620 (N_22620,N_20757,N_21336);
nand U22621 (N_22621,N_19413,N_18777);
or U22622 (N_22622,N_21852,N_18857);
nand U22623 (N_22623,N_18958,N_20271);
nand U22624 (N_22624,N_19921,N_21422);
and U22625 (N_22625,N_20316,N_21799);
and U22626 (N_22626,N_21006,N_20428);
or U22627 (N_22627,N_18917,N_19715);
nand U22628 (N_22628,N_19605,N_21106);
nor U22629 (N_22629,N_20080,N_20127);
or U22630 (N_22630,N_21111,N_19109);
xnor U22631 (N_22631,N_19569,N_19103);
nand U22632 (N_22632,N_19520,N_19691);
or U22633 (N_22633,N_21246,N_19708);
nor U22634 (N_22634,N_18751,N_19036);
and U22635 (N_22635,N_21613,N_21125);
nor U22636 (N_22636,N_20336,N_18791);
or U22637 (N_22637,N_21690,N_21302);
xor U22638 (N_22638,N_19159,N_20907);
xor U22639 (N_22639,N_20223,N_20167);
or U22640 (N_22640,N_20067,N_19636);
nand U22641 (N_22641,N_21368,N_21388);
or U22642 (N_22642,N_20631,N_21294);
nand U22643 (N_22643,N_21117,N_20825);
and U22644 (N_22644,N_18833,N_19926);
and U22645 (N_22645,N_18908,N_21395);
xnor U22646 (N_22646,N_19077,N_21073);
xor U22647 (N_22647,N_21270,N_19130);
and U22648 (N_22648,N_20971,N_19460);
xor U22649 (N_22649,N_21224,N_21109);
and U22650 (N_22650,N_21156,N_19451);
nor U22651 (N_22651,N_20968,N_19476);
and U22652 (N_22652,N_19555,N_20633);
nor U22653 (N_22653,N_19793,N_20392);
xor U22654 (N_22654,N_21484,N_20043);
nor U22655 (N_22655,N_20013,N_20452);
and U22656 (N_22656,N_21685,N_18780);
xnor U22657 (N_22657,N_21213,N_20130);
nor U22658 (N_22658,N_20292,N_20359);
and U22659 (N_22659,N_19439,N_19043);
or U22660 (N_22660,N_20919,N_21205);
nand U22661 (N_22661,N_21169,N_20333);
nand U22662 (N_22662,N_21736,N_21603);
nor U22663 (N_22663,N_20824,N_19046);
nand U22664 (N_22664,N_20597,N_20423);
or U22665 (N_22665,N_21242,N_21353);
xor U22666 (N_22666,N_21319,N_21343);
or U22667 (N_22667,N_19977,N_20600);
and U22668 (N_22668,N_19908,N_20934);
and U22669 (N_22669,N_20242,N_20224);
xnor U22670 (N_22670,N_19647,N_20437);
xnor U22671 (N_22671,N_19918,N_19599);
or U22672 (N_22672,N_20285,N_20412);
or U22673 (N_22673,N_21298,N_19360);
nand U22674 (N_22674,N_19969,N_20182);
or U22675 (N_22675,N_21466,N_20354);
nor U22676 (N_22676,N_19638,N_18877);
nand U22677 (N_22677,N_20394,N_19718);
xnor U22678 (N_22678,N_19546,N_21314);
nor U22679 (N_22679,N_20323,N_21168);
nand U22680 (N_22680,N_20659,N_20588);
nor U22681 (N_22681,N_20592,N_21085);
nor U22682 (N_22682,N_19016,N_20341);
xnor U22683 (N_22683,N_19010,N_21838);
nand U22684 (N_22684,N_21665,N_19699);
and U22685 (N_22685,N_18829,N_18895);
or U22686 (N_22686,N_21086,N_21411);
or U22687 (N_22687,N_20712,N_20645);
and U22688 (N_22688,N_21777,N_21842);
or U22689 (N_22689,N_19626,N_21179);
nor U22690 (N_22690,N_19878,N_21740);
xnor U22691 (N_22691,N_19162,N_20789);
and U22692 (N_22692,N_20790,N_20087);
xnor U22693 (N_22693,N_21808,N_20516);
nor U22694 (N_22694,N_19812,N_21702);
xor U22695 (N_22695,N_19534,N_20290);
and U22696 (N_22696,N_21288,N_19008);
nor U22697 (N_22697,N_19473,N_19845);
xor U22698 (N_22698,N_20068,N_19843);
and U22699 (N_22699,N_19142,N_19872);
nor U22700 (N_22700,N_20785,N_20312);
nand U22701 (N_22701,N_21836,N_20944);
or U22702 (N_22702,N_21172,N_19347);
or U22703 (N_22703,N_21022,N_18778);
xnor U22704 (N_22704,N_19538,N_20660);
or U22705 (N_22705,N_21841,N_20461);
nand U22706 (N_22706,N_19980,N_19999);
and U22707 (N_22707,N_18994,N_19535);
and U22708 (N_22708,N_20626,N_18999);
nor U22709 (N_22709,N_19589,N_19841);
xnor U22710 (N_22710,N_20860,N_19672);
xor U22711 (N_22711,N_20288,N_20211);
and U22712 (N_22712,N_19985,N_21352);
and U22713 (N_22713,N_20178,N_19986);
nand U22714 (N_22714,N_19290,N_20613);
nand U22715 (N_22715,N_19361,N_19596);
and U22716 (N_22716,N_20929,N_20280);
or U22717 (N_22717,N_20612,N_20322);
xor U22718 (N_22718,N_20411,N_19494);
nor U22719 (N_22719,N_20576,N_21000);
xor U22720 (N_22720,N_19346,N_20769);
and U22721 (N_22721,N_21253,N_19404);
or U22722 (N_22722,N_20002,N_18896);
and U22723 (N_22723,N_21099,N_19640);
and U22724 (N_22724,N_21630,N_19131);
nand U22725 (N_22725,N_20348,N_19698);
nor U22726 (N_22726,N_21037,N_21489);
nand U22727 (N_22727,N_21262,N_21414);
xor U22728 (N_22728,N_20730,N_19592);
or U22729 (N_22729,N_20961,N_18940);
nor U22730 (N_22730,N_19521,N_19530);
and U22731 (N_22731,N_21425,N_18991);
or U22732 (N_22732,N_19384,N_21774);
and U22733 (N_22733,N_19078,N_19809);
and U22734 (N_22734,N_20240,N_21619);
and U22735 (N_22735,N_18827,N_21264);
or U22736 (N_22736,N_19591,N_18753);
xnor U22737 (N_22737,N_21292,N_19559);
nor U22738 (N_22738,N_19664,N_21839);
xnor U22739 (N_22739,N_21758,N_21837);
and U22740 (N_22740,N_19200,N_20206);
xor U22741 (N_22741,N_18910,N_20868);
and U22742 (N_22742,N_21097,N_18954);
nand U22743 (N_22743,N_21385,N_21017);
xnor U22744 (N_22744,N_21519,N_19689);
nor U22745 (N_22745,N_21483,N_18956);
or U22746 (N_22746,N_18870,N_20545);
xor U22747 (N_22747,N_20226,N_21371);
and U22748 (N_22748,N_21650,N_18938);
xor U22749 (N_22749,N_20696,N_19961);
xnor U22750 (N_22750,N_21061,N_21666);
nor U22751 (N_22751,N_21581,N_20568);
nand U22752 (N_22752,N_21538,N_20154);
xnor U22753 (N_22753,N_19397,N_20187);
nand U22754 (N_22754,N_21100,N_20366);
xor U22755 (N_22755,N_19444,N_21201);
nand U22756 (N_22756,N_21548,N_20135);
and U22757 (N_22757,N_18802,N_20365);
and U22758 (N_22758,N_19857,N_19703);
or U22759 (N_22759,N_20279,N_20304);
nor U22760 (N_22760,N_20384,N_21209);
or U22761 (N_22761,N_19031,N_20324);
nor U22762 (N_22762,N_21511,N_20515);
xnor U22763 (N_22763,N_19624,N_21671);
or U22764 (N_22764,N_19456,N_20904);
nand U22765 (N_22765,N_21114,N_19542);
and U22766 (N_22766,N_20689,N_20553);
nand U22767 (N_22767,N_20827,N_19728);
xnor U22768 (N_22768,N_21074,N_19881);
or U22769 (N_22769,N_21771,N_21713);
nor U22770 (N_22770,N_19768,N_20925);
nor U22771 (N_22771,N_21480,N_21624);
and U22772 (N_22772,N_20111,N_21809);
nor U22773 (N_22773,N_20092,N_19148);
or U22774 (N_22774,N_20675,N_21102);
xor U22775 (N_22775,N_21565,N_20745);
xnor U22776 (N_22776,N_19474,N_21092);
nand U22777 (N_22777,N_20655,N_18821);
or U22778 (N_22778,N_18995,N_20984);
xor U22779 (N_22779,N_21301,N_19953);
nand U22780 (N_22780,N_21033,N_20694);
nor U22781 (N_22781,N_19287,N_20263);
and U22782 (N_22782,N_19897,N_20686);
or U22783 (N_22783,N_19073,N_20977);
nand U22784 (N_22784,N_20561,N_21563);
or U22785 (N_22785,N_19087,N_21202);
nor U22786 (N_22786,N_21128,N_19677);
nor U22787 (N_22787,N_18795,N_19905);
or U22788 (N_22788,N_21539,N_19479);
xnor U22789 (N_22789,N_20218,N_19151);
nand U22790 (N_22790,N_19443,N_21020);
xnor U22791 (N_22791,N_20181,N_20941);
xor U22792 (N_22792,N_20801,N_21788);
and U22793 (N_22793,N_19692,N_21178);
xor U22794 (N_22794,N_19203,N_21717);
and U22795 (N_22795,N_19419,N_21098);
or U22796 (N_22796,N_19818,N_21330);
or U22797 (N_22797,N_19402,N_20146);
or U22798 (N_22798,N_20388,N_20774);
or U22799 (N_22799,N_19895,N_19772);
and U22800 (N_22800,N_19724,N_20814);
nand U22801 (N_22801,N_19983,N_19282);
nor U22802 (N_22802,N_21525,N_19940);
xor U22803 (N_22803,N_19752,N_18876);
and U22804 (N_22804,N_20132,N_19788);
xnor U22805 (N_22805,N_21072,N_19338);
nand U22806 (N_22806,N_18886,N_20955);
nor U22807 (N_22807,N_20948,N_21445);
or U22808 (N_22808,N_19751,N_19201);
and U22809 (N_22809,N_18919,N_21312);
nand U22810 (N_22810,N_18897,N_21518);
or U22811 (N_22811,N_19807,N_20251);
nor U22812 (N_22812,N_21818,N_21428);
or U22813 (N_22813,N_18980,N_21332);
and U22814 (N_22814,N_21438,N_21507);
nand U22815 (N_22815,N_21746,N_21269);
xnor U22816 (N_22816,N_19002,N_20328);
or U22817 (N_22817,N_21463,N_20591);
nand U22818 (N_22818,N_19851,N_20194);
xnor U22819 (N_22819,N_19762,N_19972);
xnor U22820 (N_22820,N_21149,N_20120);
xnor U22821 (N_22821,N_21166,N_21739);
or U22822 (N_22822,N_21566,N_21683);
or U22823 (N_22823,N_19663,N_21500);
nor U22824 (N_22824,N_19962,N_20053);
xor U22825 (N_22825,N_19597,N_21743);
nand U22826 (N_22826,N_19642,N_18796);
nor U22827 (N_22827,N_19447,N_19713);
xor U22828 (N_22828,N_21070,N_20867);
xor U22829 (N_22829,N_19228,N_21347);
nor U22830 (N_22830,N_19979,N_19272);
or U22831 (N_22831,N_21864,N_19295);
nor U22832 (N_22832,N_19245,N_21359);
xnor U22833 (N_22833,N_21335,N_19981);
nand U22834 (N_22834,N_20142,N_20386);
or U22835 (N_22835,N_19607,N_19132);
nand U22836 (N_22836,N_21608,N_21194);
xnor U22837 (N_22837,N_20165,N_20440);
nand U22838 (N_22838,N_20008,N_21058);
nor U22839 (N_22839,N_19526,N_20993);
and U22840 (N_22840,N_20786,N_21661);
xnor U22841 (N_22841,N_19212,N_21623);
nor U22842 (N_22842,N_21048,N_19651);
xor U22843 (N_22843,N_20936,N_19571);
or U22844 (N_22844,N_20321,N_21184);
xnor U22845 (N_22845,N_21553,N_20486);
and U22846 (N_22846,N_20946,N_19602);
xnor U22847 (N_22847,N_20767,N_20432);
xnor U22848 (N_22848,N_20032,N_19648);
nor U22849 (N_22849,N_21531,N_20916);
or U22850 (N_22850,N_21083,N_21693);
xnor U22851 (N_22851,N_19169,N_20425);
and U22852 (N_22852,N_20048,N_21783);
nor U22853 (N_22853,N_21605,N_19262);
nand U22854 (N_22854,N_20875,N_19332);
and U22855 (N_22855,N_20462,N_19674);
nor U22856 (N_22856,N_19367,N_19868);
xor U22857 (N_22857,N_19271,N_21225);
and U22858 (N_22858,N_19958,N_21574);
nand U22859 (N_22859,N_18871,N_19028);
or U22860 (N_22860,N_21540,N_20534);
nor U22861 (N_22861,N_19802,N_20248);
xnor U22862 (N_22862,N_20325,N_20262);
nor U22863 (N_22863,N_19220,N_21499);
nand U22864 (N_22864,N_19330,N_19582);
or U22865 (N_22865,N_19611,N_20104);
xor U22866 (N_22866,N_20398,N_19714);
and U22867 (N_22867,N_19168,N_19840);
nor U22868 (N_22868,N_19991,N_20144);
or U22869 (N_22869,N_19441,N_20327);
nor U22870 (N_22870,N_21113,N_19873);
nand U22871 (N_22871,N_19902,N_20834);
xor U22872 (N_22872,N_19414,N_19039);
or U22873 (N_22873,N_19117,N_20744);
nand U22874 (N_22874,N_19950,N_20995);
or U22875 (N_22875,N_19615,N_20387);
xor U22876 (N_22876,N_19071,N_18786);
nand U22877 (N_22877,N_21733,N_19504);
and U22878 (N_22878,N_20065,N_20750);
or U22879 (N_22879,N_19914,N_19785);
xnor U22880 (N_22880,N_19324,N_19477);
nor U22881 (N_22881,N_20957,N_19471);
nor U22882 (N_22882,N_20198,N_20851);
xnor U22883 (N_22883,N_21027,N_21135);
or U22884 (N_22884,N_21132,N_21577);
or U22885 (N_22885,N_19416,N_18826);
xor U22886 (N_22886,N_19756,N_19411);
nor U22887 (N_22887,N_21502,N_19668);
xor U22888 (N_22888,N_21763,N_18858);
or U22889 (N_22889,N_21389,N_18941);
nor U22890 (N_22890,N_18920,N_20272);
nand U22891 (N_22891,N_21005,N_20780);
nand U22892 (N_22892,N_21433,N_19273);
nand U22893 (N_22893,N_20039,N_21137);
nand U22894 (N_22894,N_20038,N_19365);
or U22895 (N_22895,N_19732,N_21546);
xnor U22896 (N_22896,N_20357,N_19133);
xor U22897 (N_22897,N_21846,N_20524);
xnor U22898 (N_22898,N_18914,N_20590);
nand U22899 (N_22899,N_19825,N_19050);
or U22900 (N_22900,N_21815,N_21835);
nand U22901 (N_22901,N_21266,N_20010);
nor U22902 (N_22902,N_21096,N_21770);
xnor U22903 (N_22903,N_21454,N_20475);
nor U22904 (N_22904,N_20962,N_21284);
and U22905 (N_22905,N_21524,N_20970);
xor U22906 (N_22906,N_19157,N_21290);
xnor U22907 (N_22907,N_19013,N_19152);
xor U22908 (N_22908,N_20150,N_18850);
nor U22909 (N_22909,N_19847,N_19206);
xor U22910 (N_22910,N_20103,N_21148);
nor U22911 (N_22911,N_19084,N_21456);
nor U22912 (N_22912,N_21440,N_19345);
or U22913 (N_22913,N_21640,N_21696);
xor U22914 (N_22914,N_20116,N_20309);
and U22915 (N_22915,N_18820,N_19129);
or U22916 (N_22916,N_21813,N_19329);
or U22917 (N_22917,N_19656,N_20579);
nor U22918 (N_22918,N_21827,N_21789);
nor U22919 (N_22919,N_20463,N_21488);
and U22920 (N_22920,N_21200,N_20577);
xor U22921 (N_22921,N_19139,N_20362);
nor U22922 (N_22922,N_20268,N_18859);
nor U22923 (N_22923,N_18831,N_20595);
nand U22924 (N_22924,N_21233,N_19335);
or U22925 (N_22925,N_20062,N_19003);
and U22926 (N_22926,N_20623,N_20275);
and U22927 (N_22927,N_19093,N_19887);
xnor U22928 (N_22928,N_20681,N_20989);
or U22929 (N_22929,N_19745,N_19813);
and U22930 (N_22930,N_19641,N_19448);
xnor U22931 (N_22931,N_20960,N_20467);
xnor U22932 (N_22932,N_20706,N_20326);
or U22933 (N_22933,N_19501,N_20210);
nor U22934 (N_22934,N_20076,N_18949);
and U22935 (N_22935,N_19234,N_21779);
and U22936 (N_22936,N_19042,N_19539);
nand U22937 (N_22937,N_21515,N_20649);
or U22938 (N_22938,N_19834,N_19464);
xnor U22939 (N_22939,N_21868,N_19846);
and U22940 (N_22940,N_20495,N_21094);
or U22941 (N_22941,N_19266,N_19350);
nor U22942 (N_22942,N_20945,N_21256);
nand U22943 (N_22943,N_20129,N_19580);
xor U22944 (N_22944,N_19325,N_21527);
nor U22945 (N_22945,N_19047,N_19835);
xnor U22946 (N_22946,N_21737,N_20532);
nand U22947 (N_22947,N_20886,N_20856);
nand U22948 (N_22948,N_19254,N_20350);
nor U22949 (N_22949,N_20395,N_21349);
and U22950 (N_22950,N_20601,N_20870);
xnor U22951 (N_22951,N_20857,N_21151);
nor U22952 (N_22952,N_20163,N_20349);
nand U22953 (N_22953,N_20361,N_21655);
xnor U22954 (N_22954,N_20747,N_21803);
xnor U22955 (N_22955,N_20369,N_18904);
nor U22956 (N_22956,N_18934,N_20985);
nand U22957 (N_22957,N_20635,N_21455);
or U22958 (N_22958,N_19213,N_21642);
nor U22959 (N_22959,N_21481,N_20258);
and U22960 (N_22960,N_19735,N_19996);
or U22961 (N_22961,N_19066,N_19064);
nor U22962 (N_22962,N_20680,N_20845);
nand U22963 (N_22963,N_21382,N_21874);
and U22964 (N_22964,N_20151,N_18982);
nor U22965 (N_22965,N_21791,N_19382);
or U22966 (N_22966,N_21367,N_19951);
xor U22967 (N_22967,N_20006,N_21429);
nand U22968 (N_22968,N_20906,N_19942);
and U22969 (N_22969,N_20711,N_21680);
xor U22970 (N_22970,N_21013,N_20221);
nor U22971 (N_22971,N_21477,N_20138);
nand U22972 (N_22972,N_20145,N_18798);
or U22973 (N_22973,N_18811,N_20732);
and U22974 (N_22974,N_18860,N_20385);
xor U22975 (N_22975,N_20709,N_21503);
xnor U22976 (N_22976,N_20465,N_20762);
nor U22977 (N_22977,N_18926,N_19510);
or U22978 (N_22978,N_21649,N_20289);
xnor U22979 (N_22979,N_19410,N_19237);
and U22980 (N_22980,N_21844,N_20729);
and U22981 (N_22981,N_20822,N_21686);
xor U22982 (N_22982,N_19355,N_20976);
nand U22983 (N_22983,N_19875,N_18968);
nand U22984 (N_22984,N_21212,N_19723);
nand U22985 (N_22985,N_18837,N_20760);
nor U22986 (N_22986,N_21611,N_20865);
and U22987 (N_22987,N_21521,N_21210);
xnor U22988 (N_22988,N_19844,N_21384);
or U22989 (N_22989,N_20083,N_21569);
nand U22990 (N_22990,N_20777,N_20179);
xnor U22991 (N_22991,N_20836,N_21039);
nand U22992 (N_22992,N_20557,N_19884);
or U22993 (N_22993,N_20710,N_20616);
nand U22994 (N_22994,N_21570,N_19801);
nor U22995 (N_22995,N_21588,N_20622);
and U22996 (N_22996,N_19328,N_18984);
and U22997 (N_22997,N_21439,N_19083);
nor U22998 (N_22998,N_19711,N_19519);
xnor U22999 (N_22999,N_20703,N_18993);
and U23000 (N_23000,N_18918,N_19965);
nor U23001 (N_23001,N_18983,N_20517);
or U23002 (N_23002,N_20567,N_19643);
and U23003 (N_23003,N_21590,N_19376);
nand U23004 (N_23004,N_20071,N_18944);
xor U23005 (N_23005,N_20370,N_20105);
nand U23006 (N_23006,N_21547,N_18955);
nor U23007 (N_23007,N_19457,N_20850);
nand U23008 (N_23008,N_19730,N_20734);
nand U23009 (N_23009,N_20772,N_19616);
and U23010 (N_23010,N_20055,N_20847);
xnor U23011 (N_23011,N_20812,N_20022);
nand U23012 (N_23012,N_20128,N_21446);
nor U23013 (N_23013,N_19667,N_19576);
nor U23014 (N_23014,N_21817,N_19850);
or U23015 (N_23015,N_21049,N_19375);
or U23016 (N_23016,N_21333,N_21801);
xor U23017 (N_23017,N_19354,N_21066);
or U23018 (N_23018,N_19288,N_19019);
xnor U23019 (N_23019,N_21450,N_18755);
and U23020 (N_23020,N_20025,N_20682);
or U23021 (N_23021,N_18799,N_21859);
xor U23022 (N_23022,N_21401,N_19579);
and U23023 (N_23023,N_19022,N_19994);
and U23024 (N_23024,N_21471,N_19586);
xor U23025 (N_23025,N_19127,N_21872);
nor U23026 (N_23026,N_20980,N_19572);
nor U23027 (N_23027,N_19233,N_20749);
xnor U23028 (N_23028,N_19412,N_19185);
and U23029 (N_23029,N_19249,N_19805);
or U23030 (N_23030,N_20728,N_19045);
and U23031 (N_23031,N_20754,N_19253);
xnor U23032 (N_23032,N_20408,N_20901);
nor U23033 (N_23033,N_19655,N_19814);
nor U23034 (N_23034,N_19134,N_19101);
nor U23035 (N_23035,N_19392,N_19782);
nor U23036 (N_23036,N_19502,N_19195);
and U23037 (N_23037,N_20064,N_20099);
nand U23038 (N_23038,N_19686,N_19092);
xnor U23039 (N_23039,N_21533,N_20410);
nand U23040 (N_23040,N_21833,N_21267);
xnor U23041 (N_23041,N_20802,N_19588);
nor U23042 (N_23042,N_20761,N_21625);
xnor U23043 (N_23043,N_20418,N_21793);
and U23044 (N_23044,N_21651,N_19497);
xnor U23045 (N_23045,N_21228,N_20663);
xor U23046 (N_23046,N_21222,N_20343);
and U23047 (N_23047,N_21797,N_20560);
and U23048 (N_23048,N_19904,N_20390);
or U23049 (N_23049,N_19794,N_21220);
and U23050 (N_23050,N_21431,N_21474);
nor U23051 (N_23051,N_21299,N_19241);
nor U23052 (N_23052,N_19442,N_21004);
or U23053 (N_23053,N_19594,N_19121);
or U23054 (N_23054,N_19917,N_20205);
or U23055 (N_23055,N_19408,N_20554);
nor U23056 (N_23056,N_19223,N_19899);
nand U23057 (N_23057,N_21369,N_19944);
xnor U23058 (N_23058,N_20956,N_20988);
and U23059 (N_23059,N_19947,N_21218);
nand U23060 (N_23060,N_21597,N_21234);
xnor U23061 (N_23061,N_19791,N_18921);
nand U23062 (N_23062,N_18760,N_18809);
or U23063 (N_23063,N_21364,N_19739);
nand U23064 (N_23064,N_20031,N_19913);
nor U23065 (N_23065,N_20451,N_19475);
and U23066 (N_23066,N_19776,N_19225);
nand U23067 (N_23067,N_21063,N_19138);
and U23068 (N_23068,N_21617,N_19349);
or U23069 (N_23069,N_19095,N_18832);
nor U23070 (N_23070,N_21724,N_21711);
and U23071 (N_23071,N_21346,N_20342);
nand U23072 (N_23072,N_19982,N_19937);
nor U23073 (N_23073,N_18978,N_18754);
nor U23074 (N_23074,N_19067,N_21626);
and U23075 (N_23075,N_21715,N_19006);
xnor U23076 (N_23076,N_19141,N_19156);
xor U23077 (N_23077,N_19975,N_20898);
or U23078 (N_23078,N_19205,N_21586);
nand U23079 (N_23079,N_20141,N_20652);
xnor U23080 (N_23080,N_19482,N_21602);
or U23081 (N_23081,N_21154,N_21089);
nor U23082 (N_23082,N_19771,N_21010);
nand U23083 (N_23083,N_21140,N_21727);
xnor U23084 (N_23084,N_20914,N_20606);
nor U23085 (N_23085,N_21420,N_21658);
xnor U23086 (N_23086,N_21832,N_18990);
xnor U23087 (N_23087,N_18759,N_19758);
xor U23088 (N_23088,N_20604,N_19378);
nor U23089 (N_23089,N_21050,N_20355);
nor U23090 (N_23090,N_19915,N_19340);
nand U23091 (N_23091,N_19603,N_21498);
nand U23092 (N_23092,N_19558,N_19634);
xor U23093 (N_23093,N_21850,N_21451);
nand U23094 (N_23094,N_19343,N_21257);
nand U23095 (N_23095,N_19727,N_20964);
nand U23096 (N_23096,N_20564,N_20900);
nor U23097 (N_23097,N_20383,N_21633);
or U23098 (N_23098,N_18813,N_18885);
and U23099 (N_23099,N_21287,N_21729);
nor U23100 (N_23100,N_19529,N_18959);
nand U23101 (N_23101,N_20269,N_19310);
nor U23102 (N_23102,N_20204,N_20037);
nor U23103 (N_23103,N_19547,N_19712);
and U23104 (N_23104,N_19866,N_19660);
or U23105 (N_23105,N_20117,N_21716);
nor U23106 (N_23106,N_20143,N_19363);
nor U23107 (N_23107,N_19214,N_20112);
xor U23108 (N_23108,N_20017,N_20913);
nor U23109 (N_23109,N_21695,N_19561);
xor U23110 (N_23110,N_19992,N_20193);
or U23111 (N_23111,N_21243,N_19030);
nor U23112 (N_23112,N_20351,N_21757);
nor U23113 (N_23113,N_21075,N_20826);
nor U23114 (N_23114,N_20161,N_20835);
xnor U23115 (N_23115,N_21453,N_19243);
xor U23116 (N_23116,N_19296,N_19267);
nor U23117 (N_23117,N_21596,N_20088);
and U23118 (N_23118,N_20001,N_20147);
nor U23119 (N_23119,N_20183,N_21612);
and U23120 (N_23120,N_20949,N_19470);
nand U23121 (N_23121,N_20640,N_18932);
xnor U23122 (N_23122,N_20125,N_21494);
nor U23123 (N_23123,N_19415,N_20273);
nand U23124 (N_23124,N_21195,N_20209);
xor U23125 (N_23125,N_19000,N_20721);
nor U23126 (N_23126,N_20726,N_18789);
or U23127 (N_23127,N_20830,N_21621);
or U23128 (N_23128,N_18992,N_20020);
nor U23129 (N_23129,N_21826,N_20430);
nand U23130 (N_23130,N_21710,N_21023);
nand U23131 (N_23131,N_20230,N_19593);
and U23132 (N_23132,N_20819,N_20555);
and U23133 (N_23133,N_21762,N_20519);
nor U23134 (N_23134,N_21667,N_21689);
and U23135 (N_23135,N_19483,N_19383);
xnor U23136 (N_23136,N_19528,N_19183);
or U23137 (N_23137,N_19380,N_21462);
xnor U23138 (N_23138,N_21432,N_19946);
nor U23139 (N_23139,N_20196,N_21133);
nand U23140 (N_23140,N_20625,N_21622);
xnor U23141 (N_23141,N_19928,N_19532);
xnor U23142 (N_23142,N_19750,N_21629);
or U23143 (N_23143,N_21035,N_19833);
and U23144 (N_23144,N_20969,N_21377);
nor U23145 (N_23145,N_21829,N_20287);
or U23146 (N_23146,N_21052,N_21593);
and U23147 (N_23147,N_20403,N_20470);
nor U23148 (N_23148,N_19828,N_19001);
nor U23149 (N_23149,N_19722,N_20406);
nand U23150 (N_23150,N_21607,N_21223);
or U23151 (N_23151,N_20502,N_19524);
and U23152 (N_23152,N_20489,N_19798);
and U23153 (N_23153,N_19398,N_20244);
xnor U23154 (N_23154,N_21537,N_19877);
nand U23155 (N_23155,N_21164,N_20339);
or U23156 (N_23156,N_20021,N_19091);
nand U23157 (N_23157,N_20953,N_20295);
xnor U23158 (N_23158,N_21856,N_19990);
nor U23159 (N_23159,N_20202,N_20007);
xnor U23160 (N_23160,N_20569,N_20589);
nor U23161 (N_23161,N_20162,N_20101);
xnor U23162 (N_23162,N_19710,N_21143);
or U23163 (N_23163,N_21819,N_20691);
nand U23164 (N_23164,N_20684,N_20176);
nand U23165 (N_23165,N_21375,N_20737);
nor U23166 (N_23166,N_21351,N_20252);
and U23167 (N_23167,N_19733,N_21514);
and U23168 (N_23168,N_19995,N_20793);
nor U23169 (N_23169,N_19256,N_19554);
or U23170 (N_23170,N_19184,N_18750);
or U23171 (N_23171,N_20192,N_19164);
and U23172 (N_23172,N_21544,N_20061);
nand U23173 (N_23173,N_19274,N_21165);
and U23174 (N_23174,N_18818,N_19583);
or U23175 (N_23175,N_20416,N_19388);
or U23176 (N_23176,N_19585,N_18891);
nor U23177 (N_23177,N_19406,N_20391);
nand U23178 (N_23178,N_20027,N_18964);
xor U23179 (N_23179,N_20173,N_21272);
xnor U23180 (N_23180,N_19563,N_20500);
and U23181 (N_23181,N_21447,N_18987);
nand U23182 (N_23182,N_21814,N_20879);
nor U23183 (N_23183,N_21318,N_21701);
or U23184 (N_23184,N_19890,N_19265);
and U23185 (N_23185,N_19823,N_20401);
nor U23186 (N_23186,N_19119,N_21790);
and U23187 (N_23187,N_19507,N_21768);
nor U23188 (N_23188,N_21360,N_20602);
nand U23189 (N_23189,N_19062,N_18758);
xor U23190 (N_23190,N_19334,N_19515);
or U23191 (N_23191,N_18893,N_18824);
and U23192 (N_23192,N_19540,N_19931);
nor U23193 (N_23193,N_21167,N_19880);
nor U23194 (N_23194,N_21523,N_21467);
or U23195 (N_23195,N_18852,N_19192);
nand U23196 (N_23196,N_20714,N_19869);
nand U23197 (N_23197,N_19053,N_21766);
nor U23198 (N_23198,N_21057,N_20334);
and U23199 (N_23199,N_20491,N_20468);
and U23200 (N_23200,N_20987,N_19500);
nor U23201 (N_23201,N_21873,N_19566);
nor U23202 (N_23202,N_19870,N_21019);
nand U23203 (N_23203,N_19671,N_20580);
xnor U23204 (N_23204,N_19491,N_19757);
nand U23205 (N_23205,N_19924,N_20671);
xor U23206 (N_23206,N_20404,N_20036);
and U23207 (N_23207,N_20507,N_20380);
and U23208 (N_23208,N_19341,N_21865);
xnor U23209 (N_23209,N_19313,N_20073);
and U23210 (N_23210,N_20469,N_19509);
and U23211 (N_23211,N_19606,N_21756);
nand U23212 (N_23212,N_20054,N_21636);
or U23213 (N_23213,N_21472,N_21759);
nand U23214 (N_23214,N_19385,N_19175);
nor U23215 (N_23215,N_19149,N_21297);
or U23216 (N_23216,N_18988,N_19747);
and U23217 (N_23217,N_21274,N_19236);
or U23218 (N_23218,N_21437,N_21652);
and U23219 (N_23219,N_21285,N_18787);
nor U23220 (N_23220,N_21587,N_19280);
xnor U23221 (N_23221,N_21060,N_20650);
xnor U23222 (N_23222,N_19661,N_19058);
nand U23223 (N_23223,N_21712,N_21635);
nor U23224 (N_23224,N_21053,N_21656);
nand U23225 (N_23225,N_19436,N_21678);
and U23226 (N_23226,N_18906,N_19075);
or U23227 (N_23227,N_21542,N_19221);
nand U23228 (N_23228,N_19852,N_18869);
and U23229 (N_23229,N_19025,N_19551);
nor U23230 (N_23230,N_21187,N_20722);
nor U23231 (N_23231,N_19082,N_19430);
xor U23232 (N_23232,N_19369,N_20599);
xor U23233 (N_23233,N_20050,N_19486);
xnor U23234 (N_23234,N_19978,N_20375);
and U23235 (N_23235,N_19065,N_19856);
xnor U23236 (N_23236,N_20413,N_19790);
or U23237 (N_23237,N_19769,N_20200);
or U23238 (N_23238,N_20809,N_19694);
nand U23239 (N_23239,N_19941,N_19701);
nand U23240 (N_23240,N_19721,N_20492);
xor U23241 (N_23241,N_18892,N_19685);
or U23242 (N_23242,N_21660,N_20439);
or U23243 (N_23243,N_20155,N_20499);
xnor U23244 (N_23244,N_19906,N_21732);
or U23245 (N_23245,N_21579,N_19283);
nand U23246 (N_23246,N_20180,N_20487);
nand U23247 (N_23247,N_21573,N_19587);
xor U23248 (N_23248,N_20433,N_20314);
nand U23249 (N_23249,N_21398,N_19452);
and U23250 (N_23250,N_20654,N_20540);
nand U23251 (N_23251,N_20858,N_19293);
or U23252 (N_23252,N_19032,N_21637);
xor U23253 (N_23253,N_21240,N_19211);
or U23254 (N_23254,N_21421,N_21423);
nor U23255 (N_23255,N_21584,N_20379);
nand U23256 (N_23256,N_19261,N_20571);
xnor U23257 (N_23257,N_20653,N_20695);
or U23258 (N_23258,N_21008,N_20693);
xnor U23259 (N_23259,N_20214,N_19242);
or U23260 (N_23260,N_21304,N_19187);
nor U23261 (N_23261,N_20239,N_20041);
or U23262 (N_23262,N_19215,N_21620);
and U23263 (N_23263,N_20241,N_21831);
and U23264 (N_23264,N_21684,N_20319);
or U23265 (N_23265,N_21776,N_19505);
nor U23266 (N_23266,N_19088,N_21802);
xnor U23267 (N_23267,N_18975,N_21221);
nor U23268 (N_23268,N_20213,N_20924);
xor U23269 (N_23269,N_19023,N_19107);
nand U23270 (N_23270,N_20921,N_21120);
and U23271 (N_23271,N_21258,N_21138);
or U23272 (N_23272,N_20140,N_19463);
nand U23273 (N_23273,N_21134,N_19717);
nand U23274 (N_23274,N_21251,N_19956);
nand U23275 (N_23275,N_20755,N_21203);
and U23276 (N_23276,N_20481,N_18936);
or U23277 (N_23277,N_20429,N_21772);
nor U23278 (N_23278,N_19281,N_18923);
or U23279 (N_23279,N_20550,N_20225);
nand U23280 (N_23280,N_20009,N_18807);
nand U23281 (N_23281,N_21152,N_19669);
nor U23282 (N_23282,N_21576,N_21780);
and U23283 (N_23283,N_21664,N_20996);
and U23284 (N_23284,N_20435,N_19279);
nand U23285 (N_23285,N_20838,N_20537);
xnor U23286 (N_23286,N_19746,N_21219);
or U23287 (N_23287,N_20741,N_20808);
and U23288 (N_23288,N_21764,N_21504);
and U23289 (N_23289,N_21559,N_18806);
xor U23290 (N_23290,N_19289,N_20436);
nand U23291 (N_23291,N_21673,N_20570);
xnor U23292 (N_23292,N_21798,N_20133);
nor U23293 (N_23293,N_21535,N_18856);
xnor U23294 (N_23294,N_21541,N_21417);
and U23295 (N_23295,N_20026,N_20552);
and U23296 (N_23296,N_20448,N_20523);
nand U23297 (N_23297,N_21674,N_20382);
or U23298 (N_23298,N_20951,N_19257);
xnor U23299 (N_23299,N_19196,N_18930);
or U23300 (N_23300,N_19373,N_21486);
xor U23301 (N_23301,N_18912,N_21720);
nor U23302 (N_23302,N_19485,N_21812);
xnor U23303 (N_23303,N_21778,N_21493);
or U23304 (N_23304,N_19789,N_20332);
and U23305 (N_23305,N_21124,N_19049);
or U23306 (N_23306,N_20019,N_20347);
xor U23307 (N_23307,N_19104,N_20878);
xnor U23308 (N_23308,N_19173,N_19680);
xor U23309 (N_23309,N_20614,N_19657);
or U23310 (N_23310,N_19459,N_19425);
nor U23311 (N_23311,N_19344,N_21016);
xnor U23312 (N_23312,N_19059,N_21784);
and U23313 (N_23313,N_21709,N_18775);
xnor U23314 (N_23314,N_20444,N_21497);
xor U23315 (N_23315,N_19098,N_21296);
xor U23316 (N_23316,N_19056,N_19337);
nand U23317 (N_23317,N_19493,N_20542);
or U23318 (N_23318,N_21703,N_20522);
xnor U23319 (N_23319,N_21354,N_18961);
nand U23320 (N_23320,N_19993,N_21199);
nor U23321 (N_23321,N_18812,N_18764);
and U23322 (N_23322,N_21782,N_21662);
nand U23323 (N_23323,N_19496,N_20768);
nand U23324 (N_23324,N_21310,N_19673);
nand U23325 (N_23325,N_19357,N_21211);
or U23326 (N_23326,N_20842,N_19548);
xnor U23327 (N_23327,N_21315,N_20164);
xor U23328 (N_23328,N_21722,N_21604);
or U23329 (N_23329,N_18825,N_20888);
nor U23330 (N_23330,N_20472,N_20441);
and U23331 (N_23331,N_19466,N_19381);
or U23332 (N_23332,N_19143,N_19409);
and U23333 (N_23333,N_19086,N_19450);
or U23334 (N_23334,N_21345,N_19922);
and U23335 (N_23335,N_20044,N_19952);
nand U23336 (N_23336,N_20217,N_18794);
nor U23337 (N_23337,N_21232,N_18817);
nand U23338 (N_23338,N_19096,N_20100);
xor U23339 (N_23339,N_19089,N_19688);
and U23340 (N_23340,N_20899,N_20346);
nor U23341 (N_23341,N_20864,N_20820);
xnor U23342 (N_23342,N_20546,N_20345);
or U23343 (N_23343,N_21247,N_19765);
or U23344 (N_23344,N_19622,N_20593);
or U23345 (N_23345,N_19855,N_18762);
xnor U23346 (N_23346,N_20377,N_21043);
nand U23347 (N_23347,N_18846,N_20966);
or U23348 (N_23348,N_19632,N_20302);
nor U23349 (N_23349,N_21358,N_21806);
nor U23350 (N_23350,N_19004,N_21754);
or U23351 (N_23351,N_19072,N_20800);
and U23352 (N_23352,N_21180,N_21465);
and U23353 (N_23353,N_20563,N_20005);
nand U23354 (N_23354,N_19573,N_21668);
nand U23355 (N_23355,N_20715,N_19763);
or U23356 (N_23356,N_20536,N_20097);
or U23357 (N_23357,N_19351,N_19923);
xnor U23358 (N_23358,N_21556,N_20884);
and U23359 (N_23359,N_20598,N_20982);
nand U23360 (N_23360,N_20705,N_21186);
nor U23361 (N_23361,N_20419,N_20286);
or U23362 (N_23362,N_20658,N_20471);
xor U23363 (N_23363,N_21370,N_21112);
nor U23364 (N_23364,N_18872,N_20282);
nand U23365 (N_23365,N_20549,N_20389);
nand U23366 (N_23366,N_19909,N_21761);
or U23367 (N_23367,N_21320,N_20704);
nor U23368 (N_23368,N_19939,N_19766);
or U23369 (N_23369,N_21328,N_21618);
xnor U23370 (N_23370,N_21176,N_20260);
nand U23371 (N_23371,N_20959,N_21029);
or U23372 (N_23372,N_19536,N_21469);
xor U23373 (N_23373,N_20775,N_21182);
nor U23374 (N_23374,N_19229,N_21475);
and U23375 (N_23375,N_19619,N_21159);
nor U23376 (N_23376,N_19687,N_21197);
nor U23377 (N_23377,N_19590,N_21059);
and U23378 (N_23378,N_21615,N_20485);
or U23379 (N_23379,N_19860,N_19208);
nand U23380 (N_23380,N_19779,N_21672);
or U23381 (N_23381,N_18804,N_21153);
or U23382 (N_23382,N_21863,N_21470);
nor U23383 (N_23383,N_21413,N_21734);
or U23384 (N_23384,N_21261,N_21181);
xor U23385 (N_23385,N_20643,N_20405);
or U23386 (N_23386,N_20238,N_21064);
xnor U23387 (N_23387,N_20891,N_19858);
or U23388 (N_23388,N_18948,N_21682);
nor U23389 (N_23389,N_18761,N_19197);
nand U23390 (N_23390,N_19079,N_20338);
or U23391 (N_23391,N_18766,N_20259);
or U23392 (N_23392,N_20483,N_20952);
xor U23393 (N_23393,N_19693,N_20733);
nand U23394 (N_23394,N_18853,N_20447);
or U23395 (N_23395,N_21103,N_20974);
or U23396 (N_23396,N_21866,N_21350);
nor U23397 (N_23397,N_21860,N_20096);
or U23398 (N_23398,N_19487,N_19005);
nand U23399 (N_23399,N_20724,N_20628);
nor U23400 (N_23400,N_20701,N_18901);
xor U23401 (N_23401,N_19428,N_20368);
xnor U23402 (N_23402,N_20504,N_20102);
nor U23403 (N_23403,N_21561,N_21150);
nor U23404 (N_23404,N_19820,N_19838);
nor U23405 (N_23405,N_21549,N_19578);
and U23406 (N_23406,N_18929,N_21362);
or U23407 (N_23407,N_20237,N_20997);
and U23408 (N_23408,N_20735,N_21372);
nand U23409 (N_23409,N_20464,N_21562);
and U23410 (N_23410,N_21670,N_21293);
nand U23411 (N_23411,N_19270,N_20699);
or U23412 (N_23412,N_20994,N_20449);
and U23413 (N_23413,N_19155,N_19842);
and U23414 (N_23414,N_21407,N_20381);
nand U23415 (N_23415,N_19252,N_19967);
or U23416 (N_23416,N_19778,N_20267);
and U23417 (N_23417,N_20407,N_20787);
xor U23418 (N_23418,N_21041,N_21248);
and U23419 (N_23419,N_19394,N_19202);
and U23420 (N_23420,N_20881,N_21707);
and U23421 (N_23421,N_19574,N_19400);
nand U23422 (N_23422,N_19327,N_21252);
or U23423 (N_23423,N_20818,N_19268);
nor U23424 (N_23424,N_19513,N_19968);
and U23425 (N_23425,N_20015,N_18836);
nand U23426 (N_23426,N_18979,N_19480);
nor U23427 (N_23427,N_20352,N_20232);
xor U23428 (N_23428,N_21277,N_20795);
xnor U23429 (N_23429,N_20846,N_21639);
nand U23430 (N_23430,N_19679,N_19076);
nand U23431 (N_23431,N_20060,N_21141);
and U23432 (N_23432,N_20090,N_19097);
or U23433 (N_23433,N_19061,N_20766);
nor U23434 (N_23434,N_19499,N_20807);
or U23435 (N_23435,N_19111,N_18843);
or U23436 (N_23436,N_20672,N_19455);
nor U23437 (N_23437,N_21173,N_21018);
nor U23438 (N_23438,N_20409,N_19271);
and U23439 (N_23439,N_20426,N_18798);
and U23440 (N_23440,N_20976,N_19153);
xor U23441 (N_23441,N_20951,N_19760);
nand U23442 (N_23442,N_20020,N_19188);
or U23443 (N_23443,N_21210,N_21658);
nor U23444 (N_23444,N_18934,N_19870);
and U23445 (N_23445,N_20704,N_19396);
xor U23446 (N_23446,N_19062,N_20827);
or U23447 (N_23447,N_20643,N_20116);
or U23448 (N_23448,N_19761,N_19713);
or U23449 (N_23449,N_20627,N_20194);
nand U23450 (N_23450,N_20033,N_19074);
and U23451 (N_23451,N_20028,N_20636);
or U23452 (N_23452,N_20450,N_21370);
nor U23453 (N_23453,N_21853,N_20994);
nor U23454 (N_23454,N_19708,N_18757);
and U23455 (N_23455,N_18912,N_20515);
nand U23456 (N_23456,N_20489,N_21566);
xor U23457 (N_23457,N_18796,N_21609);
and U23458 (N_23458,N_21861,N_20700);
and U23459 (N_23459,N_20518,N_19114);
or U23460 (N_23460,N_21754,N_20994);
xnor U23461 (N_23461,N_19190,N_18886);
or U23462 (N_23462,N_20741,N_20677);
nor U23463 (N_23463,N_20191,N_20995);
xnor U23464 (N_23464,N_18974,N_19887);
nand U23465 (N_23465,N_21788,N_19068);
or U23466 (N_23466,N_21233,N_19240);
or U23467 (N_23467,N_19781,N_21573);
or U23468 (N_23468,N_21632,N_20829);
and U23469 (N_23469,N_19756,N_19113);
nand U23470 (N_23470,N_20048,N_21194);
xor U23471 (N_23471,N_18886,N_21317);
nor U23472 (N_23472,N_20058,N_19068);
nor U23473 (N_23473,N_21348,N_19938);
xor U23474 (N_23474,N_19758,N_19465);
xnor U23475 (N_23475,N_20785,N_18822);
nand U23476 (N_23476,N_19602,N_20418);
nor U23477 (N_23477,N_20347,N_20200);
or U23478 (N_23478,N_19474,N_19335);
xnor U23479 (N_23479,N_20457,N_19123);
xor U23480 (N_23480,N_19827,N_20494);
xnor U23481 (N_23481,N_20310,N_19844);
xor U23482 (N_23482,N_21546,N_20245);
and U23483 (N_23483,N_21250,N_21848);
or U23484 (N_23484,N_21842,N_20507);
and U23485 (N_23485,N_19529,N_21214);
or U23486 (N_23486,N_20131,N_19650);
nand U23487 (N_23487,N_21190,N_21803);
xnor U23488 (N_23488,N_20588,N_20255);
or U23489 (N_23489,N_21688,N_20070);
or U23490 (N_23490,N_20627,N_21163);
xnor U23491 (N_23491,N_19621,N_20856);
or U23492 (N_23492,N_19676,N_21597);
xor U23493 (N_23493,N_21069,N_19377);
nor U23494 (N_23494,N_20973,N_21240);
and U23495 (N_23495,N_21597,N_21748);
or U23496 (N_23496,N_20436,N_20708);
and U23497 (N_23497,N_19987,N_19523);
nand U23498 (N_23498,N_19159,N_19251);
xnor U23499 (N_23499,N_21585,N_19851);
xnor U23500 (N_23500,N_20875,N_19475);
or U23501 (N_23501,N_21240,N_20450);
nor U23502 (N_23502,N_20032,N_20786);
xor U23503 (N_23503,N_21693,N_19350);
and U23504 (N_23504,N_19719,N_19589);
and U23505 (N_23505,N_21358,N_20296);
nor U23506 (N_23506,N_19598,N_18850);
nand U23507 (N_23507,N_21441,N_21715);
and U23508 (N_23508,N_20032,N_19761);
nor U23509 (N_23509,N_19868,N_18997);
nor U23510 (N_23510,N_18988,N_19267);
nand U23511 (N_23511,N_20718,N_20843);
or U23512 (N_23512,N_21132,N_21474);
and U23513 (N_23513,N_20752,N_21126);
or U23514 (N_23514,N_19931,N_18830);
and U23515 (N_23515,N_19877,N_20009);
and U23516 (N_23516,N_21708,N_21784);
or U23517 (N_23517,N_20413,N_21458);
xnor U23518 (N_23518,N_18867,N_21376);
or U23519 (N_23519,N_21086,N_21705);
nand U23520 (N_23520,N_20503,N_21333);
nor U23521 (N_23521,N_21264,N_19894);
and U23522 (N_23522,N_19513,N_20723);
xnor U23523 (N_23523,N_21588,N_20616);
nor U23524 (N_23524,N_19812,N_20385);
nand U23525 (N_23525,N_19121,N_21551);
xnor U23526 (N_23526,N_20420,N_19583);
nor U23527 (N_23527,N_19201,N_20800);
nor U23528 (N_23528,N_21558,N_20845);
nor U23529 (N_23529,N_21677,N_21857);
or U23530 (N_23530,N_20255,N_18970);
nor U23531 (N_23531,N_20487,N_21140);
and U23532 (N_23532,N_21091,N_20186);
and U23533 (N_23533,N_19045,N_21606);
and U23534 (N_23534,N_19880,N_20387);
and U23535 (N_23535,N_21213,N_20758);
or U23536 (N_23536,N_20410,N_21455);
nand U23537 (N_23537,N_19369,N_19186);
nand U23538 (N_23538,N_20029,N_20364);
or U23539 (N_23539,N_21322,N_19951);
nor U23540 (N_23540,N_19047,N_19304);
nand U23541 (N_23541,N_21434,N_20297);
nand U23542 (N_23542,N_20469,N_21476);
xnor U23543 (N_23543,N_19954,N_20509);
and U23544 (N_23544,N_20037,N_18847);
xnor U23545 (N_23545,N_21247,N_21824);
or U23546 (N_23546,N_21748,N_20743);
or U23547 (N_23547,N_19715,N_21178);
nor U23548 (N_23548,N_21324,N_19308);
xor U23549 (N_23549,N_21084,N_20756);
xnor U23550 (N_23550,N_20887,N_19326);
and U23551 (N_23551,N_19660,N_21859);
nor U23552 (N_23552,N_21737,N_18842);
xnor U23553 (N_23553,N_21172,N_21728);
nor U23554 (N_23554,N_19988,N_20944);
xor U23555 (N_23555,N_21737,N_21387);
or U23556 (N_23556,N_19139,N_19203);
nand U23557 (N_23557,N_21378,N_21229);
xor U23558 (N_23558,N_21530,N_21669);
nand U23559 (N_23559,N_21328,N_21622);
nor U23560 (N_23560,N_19607,N_21705);
xnor U23561 (N_23561,N_19395,N_21187);
xor U23562 (N_23562,N_18998,N_21282);
and U23563 (N_23563,N_21626,N_21063);
xnor U23564 (N_23564,N_20116,N_21247);
and U23565 (N_23565,N_20976,N_21801);
nor U23566 (N_23566,N_19567,N_19784);
or U23567 (N_23567,N_19476,N_18992);
nor U23568 (N_23568,N_19699,N_19070);
xor U23569 (N_23569,N_20993,N_19403);
xnor U23570 (N_23570,N_21863,N_20607);
or U23571 (N_23571,N_20865,N_19716);
nand U23572 (N_23572,N_21028,N_21783);
nand U23573 (N_23573,N_18822,N_19938);
nor U23574 (N_23574,N_19035,N_20676);
xor U23575 (N_23575,N_19629,N_20877);
or U23576 (N_23576,N_19545,N_20744);
nor U23577 (N_23577,N_21169,N_19054);
xnor U23578 (N_23578,N_19177,N_21101);
and U23579 (N_23579,N_20010,N_19889);
xnor U23580 (N_23580,N_19640,N_21280);
nor U23581 (N_23581,N_18960,N_21116);
or U23582 (N_23582,N_19628,N_21157);
and U23583 (N_23583,N_20561,N_19395);
xnor U23584 (N_23584,N_21335,N_21525);
nand U23585 (N_23585,N_19977,N_19016);
and U23586 (N_23586,N_21787,N_20152);
nor U23587 (N_23587,N_21186,N_18916);
xnor U23588 (N_23588,N_20205,N_19684);
nand U23589 (N_23589,N_21201,N_18941);
nor U23590 (N_23590,N_19566,N_21207);
and U23591 (N_23591,N_21573,N_21719);
xor U23592 (N_23592,N_20727,N_19014);
or U23593 (N_23593,N_20734,N_19136);
xor U23594 (N_23594,N_20950,N_20495);
nor U23595 (N_23595,N_19358,N_18865);
and U23596 (N_23596,N_20446,N_19815);
nand U23597 (N_23597,N_19116,N_21811);
and U23598 (N_23598,N_21436,N_19836);
xor U23599 (N_23599,N_21132,N_19884);
nand U23600 (N_23600,N_21673,N_19110);
xnor U23601 (N_23601,N_19767,N_19937);
and U23602 (N_23602,N_19649,N_19929);
xnor U23603 (N_23603,N_19111,N_21209);
or U23604 (N_23604,N_21616,N_19971);
or U23605 (N_23605,N_19120,N_20809);
nor U23606 (N_23606,N_21577,N_19680);
and U23607 (N_23607,N_18816,N_20223);
nor U23608 (N_23608,N_20155,N_20321);
and U23609 (N_23609,N_20759,N_19958);
or U23610 (N_23610,N_20405,N_20930);
nand U23611 (N_23611,N_19888,N_21688);
nand U23612 (N_23612,N_21813,N_21844);
nor U23613 (N_23613,N_21631,N_19688);
nor U23614 (N_23614,N_20472,N_21500);
and U23615 (N_23615,N_21462,N_20404);
and U23616 (N_23616,N_21086,N_20509);
or U23617 (N_23617,N_19251,N_20897);
xor U23618 (N_23618,N_20655,N_20557);
and U23619 (N_23619,N_19251,N_19538);
or U23620 (N_23620,N_19804,N_19757);
xor U23621 (N_23621,N_20236,N_19745);
nor U23622 (N_23622,N_20281,N_19277);
or U23623 (N_23623,N_19252,N_20188);
and U23624 (N_23624,N_21256,N_20232);
or U23625 (N_23625,N_19460,N_18951);
nor U23626 (N_23626,N_20054,N_18882);
or U23627 (N_23627,N_20501,N_21816);
and U23628 (N_23628,N_19114,N_19495);
or U23629 (N_23629,N_20667,N_20936);
nand U23630 (N_23630,N_21183,N_21262);
nand U23631 (N_23631,N_19666,N_19612);
nand U23632 (N_23632,N_19686,N_21674);
nand U23633 (N_23633,N_19992,N_19063);
nor U23634 (N_23634,N_21460,N_20847);
xnor U23635 (N_23635,N_19768,N_20502);
nor U23636 (N_23636,N_21552,N_19896);
or U23637 (N_23637,N_21215,N_19230);
xnor U23638 (N_23638,N_21383,N_18948);
nor U23639 (N_23639,N_21713,N_19648);
and U23640 (N_23640,N_19583,N_19919);
and U23641 (N_23641,N_20337,N_18768);
and U23642 (N_23642,N_20558,N_20133);
nand U23643 (N_23643,N_21432,N_20018);
nand U23644 (N_23644,N_19125,N_21804);
xnor U23645 (N_23645,N_21114,N_19594);
xor U23646 (N_23646,N_20248,N_21142);
xor U23647 (N_23647,N_19168,N_19553);
nand U23648 (N_23648,N_20150,N_19234);
nand U23649 (N_23649,N_19866,N_20214);
or U23650 (N_23650,N_21728,N_20666);
nand U23651 (N_23651,N_19090,N_20709);
or U23652 (N_23652,N_19710,N_20473);
or U23653 (N_23653,N_18755,N_19191);
and U23654 (N_23654,N_20682,N_19898);
xor U23655 (N_23655,N_19282,N_21067);
nor U23656 (N_23656,N_21847,N_19093);
and U23657 (N_23657,N_19487,N_20797);
or U23658 (N_23658,N_20226,N_19653);
and U23659 (N_23659,N_19068,N_20505);
xnor U23660 (N_23660,N_20553,N_21829);
nor U23661 (N_23661,N_19641,N_19689);
nor U23662 (N_23662,N_18843,N_21213);
or U23663 (N_23663,N_21021,N_20492);
xor U23664 (N_23664,N_20230,N_21416);
xor U23665 (N_23665,N_20002,N_20351);
and U23666 (N_23666,N_19359,N_21667);
or U23667 (N_23667,N_19880,N_19743);
and U23668 (N_23668,N_20882,N_19372);
nor U23669 (N_23669,N_19618,N_19859);
nor U23670 (N_23670,N_20756,N_18834);
nand U23671 (N_23671,N_21242,N_21428);
xnor U23672 (N_23672,N_19776,N_19974);
or U23673 (N_23673,N_21797,N_20352);
and U23674 (N_23674,N_21779,N_19648);
or U23675 (N_23675,N_21823,N_19649);
nor U23676 (N_23676,N_19494,N_20284);
nand U23677 (N_23677,N_19931,N_21102);
xnor U23678 (N_23678,N_20587,N_20980);
xnor U23679 (N_23679,N_20453,N_21575);
nor U23680 (N_23680,N_19023,N_21407);
and U23681 (N_23681,N_21640,N_20204);
xor U23682 (N_23682,N_19280,N_21855);
nand U23683 (N_23683,N_21337,N_20296);
nand U23684 (N_23684,N_19482,N_20900);
nor U23685 (N_23685,N_18788,N_21795);
and U23686 (N_23686,N_19529,N_21095);
nor U23687 (N_23687,N_21130,N_19278);
nand U23688 (N_23688,N_20010,N_19968);
nor U23689 (N_23689,N_20254,N_19400);
nand U23690 (N_23690,N_20938,N_20582);
and U23691 (N_23691,N_21506,N_21036);
nor U23692 (N_23692,N_20085,N_20779);
nand U23693 (N_23693,N_20448,N_19024);
or U23694 (N_23694,N_19029,N_20576);
nor U23695 (N_23695,N_21409,N_20898);
xnor U23696 (N_23696,N_19822,N_20467);
nand U23697 (N_23697,N_18758,N_19282);
nor U23698 (N_23698,N_20781,N_20050);
and U23699 (N_23699,N_20400,N_19876);
xor U23700 (N_23700,N_21403,N_21394);
nor U23701 (N_23701,N_19785,N_20433);
and U23702 (N_23702,N_20151,N_19136);
nor U23703 (N_23703,N_20447,N_21372);
and U23704 (N_23704,N_21066,N_20872);
and U23705 (N_23705,N_21871,N_18966);
nor U23706 (N_23706,N_21223,N_18980);
nand U23707 (N_23707,N_20628,N_21374);
nand U23708 (N_23708,N_21574,N_20254);
and U23709 (N_23709,N_18800,N_20259);
xor U23710 (N_23710,N_20873,N_20253);
and U23711 (N_23711,N_19829,N_20122);
nor U23712 (N_23712,N_20945,N_20229);
and U23713 (N_23713,N_19518,N_20918);
xnor U23714 (N_23714,N_19855,N_21193);
xnor U23715 (N_23715,N_20256,N_21249);
nor U23716 (N_23716,N_20285,N_19870);
or U23717 (N_23717,N_19608,N_21434);
xor U23718 (N_23718,N_21301,N_19113);
and U23719 (N_23719,N_21672,N_21599);
or U23720 (N_23720,N_19842,N_20964);
or U23721 (N_23721,N_19628,N_19163);
nand U23722 (N_23722,N_21479,N_21387);
nand U23723 (N_23723,N_19337,N_20902);
and U23724 (N_23724,N_21583,N_19997);
or U23725 (N_23725,N_21747,N_20661);
nand U23726 (N_23726,N_21243,N_20501);
and U23727 (N_23727,N_21220,N_21034);
nor U23728 (N_23728,N_19214,N_21145);
nand U23729 (N_23729,N_21132,N_21054);
or U23730 (N_23730,N_19421,N_21499);
nand U23731 (N_23731,N_19677,N_20010);
or U23732 (N_23732,N_21707,N_21435);
xor U23733 (N_23733,N_21321,N_19105);
or U23734 (N_23734,N_20247,N_20684);
or U23735 (N_23735,N_19830,N_19027);
or U23736 (N_23736,N_19679,N_19999);
xor U23737 (N_23737,N_20279,N_19898);
or U23738 (N_23738,N_20060,N_19171);
xor U23739 (N_23739,N_21352,N_21501);
xnor U23740 (N_23740,N_19035,N_19622);
nor U23741 (N_23741,N_19467,N_20400);
and U23742 (N_23742,N_19213,N_19337);
xnor U23743 (N_23743,N_20736,N_21293);
nand U23744 (N_23744,N_21549,N_20617);
and U23745 (N_23745,N_20977,N_21300);
nor U23746 (N_23746,N_20062,N_20442);
xnor U23747 (N_23747,N_21477,N_19924);
nand U23748 (N_23748,N_21356,N_21697);
or U23749 (N_23749,N_20611,N_18935);
nand U23750 (N_23750,N_21312,N_20541);
nor U23751 (N_23751,N_20604,N_19458);
xor U23752 (N_23752,N_19038,N_21159);
or U23753 (N_23753,N_21512,N_20548);
or U23754 (N_23754,N_20204,N_20687);
nand U23755 (N_23755,N_21413,N_21084);
xor U23756 (N_23756,N_21711,N_20411);
or U23757 (N_23757,N_20350,N_19334);
nand U23758 (N_23758,N_21799,N_19576);
nand U23759 (N_23759,N_19897,N_19268);
xor U23760 (N_23760,N_20691,N_21830);
or U23761 (N_23761,N_21275,N_20679);
xnor U23762 (N_23762,N_20117,N_19733);
nand U23763 (N_23763,N_21334,N_20714);
xor U23764 (N_23764,N_20812,N_19987);
nor U23765 (N_23765,N_19250,N_20164);
xor U23766 (N_23766,N_18807,N_20642);
nor U23767 (N_23767,N_20570,N_18987);
and U23768 (N_23768,N_18838,N_19933);
nand U23769 (N_23769,N_18781,N_21608);
nor U23770 (N_23770,N_19111,N_20592);
xor U23771 (N_23771,N_19037,N_21357);
xor U23772 (N_23772,N_21024,N_21865);
and U23773 (N_23773,N_20729,N_18781);
nor U23774 (N_23774,N_19483,N_19132);
nand U23775 (N_23775,N_19084,N_20161);
or U23776 (N_23776,N_19045,N_19201);
and U23777 (N_23777,N_20423,N_20384);
and U23778 (N_23778,N_20554,N_19454);
xnor U23779 (N_23779,N_20952,N_21031);
nor U23780 (N_23780,N_19001,N_19666);
nand U23781 (N_23781,N_19156,N_20285);
xor U23782 (N_23782,N_19113,N_19626);
and U23783 (N_23783,N_19019,N_18907);
xor U23784 (N_23784,N_20193,N_19240);
nor U23785 (N_23785,N_20886,N_19902);
xnor U23786 (N_23786,N_19925,N_21464);
nand U23787 (N_23787,N_21639,N_20992);
nor U23788 (N_23788,N_19875,N_20368);
nand U23789 (N_23789,N_20256,N_21071);
and U23790 (N_23790,N_20161,N_19241);
nand U23791 (N_23791,N_19167,N_20196);
xor U23792 (N_23792,N_21673,N_19746);
xnor U23793 (N_23793,N_20099,N_19297);
xnor U23794 (N_23794,N_21320,N_19017);
or U23795 (N_23795,N_18924,N_18821);
xnor U23796 (N_23796,N_18877,N_19466);
and U23797 (N_23797,N_20065,N_20159);
or U23798 (N_23798,N_19922,N_19652);
xnor U23799 (N_23799,N_20990,N_20093);
nor U23800 (N_23800,N_20139,N_19209);
nand U23801 (N_23801,N_20161,N_19703);
xnor U23802 (N_23802,N_20514,N_19384);
xor U23803 (N_23803,N_20917,N_20364);
nor U23804 (N_23804,N_20650,N_19387);
and U23805 (N_23805,N_21315,N_21416);
and U23806 (N_23806,N_19436,N_20626);
xor U23807 (N_23807,N_21264,N_21338);
or U23808 (N_23808,N_20214,N_20850);
xor U23809 (N_23809,N_21499,N_20093);
or U23810 (N_23810,N_21050,N_21859);
and U23811 (N_23811,N_19664,N_21748);
or U23812 (N_23812,N_18935,N_21508);
xnor U23813 (N_23813,N_20904,N_21061);
nor U23814 (N_23814,N_19884,N_19792);
and U23815 (N_23815,N_21555,N_19320);
nor U23816 (N_23816,N_19515,N_20044);
xor U23817 (N_23817,N_18954,N_20410);
nor U23818 (N_23818,N_21283,N_18956);
xor U23819 (N_23819,N_19844,N_20828);
and U23820 (N_23820,N_21171,N_21679);
xor U23821 (N_23821,N_21598,N_21421);
nand U23822 (N_23822,N_21837,N_19809);
nor U23823 (N_23823,N_19435,N_18828);
nand U23824 (N_23824,N_18819,N_21373);
nand U23825 (N_23825,N_19062,N_19961);
nand U23826 (N_23826,N_21145,N_20615);
and U23827 (N_23827,N_21837,N_21750);
nand U23828 (N_23828,N_20658,N_19372);
nor U23829 (N_23829,N_19960,N_19750);
nand U23830 (N_23830,N_21057,N_19989);
nand U23831 (N_23831,N_18936,N_20343);
nor U23832 (N_23832,N_21217,N_19541);
or U23833 (N_23833,N_19469,N_19824);
nand U23834 (N_23834,N_18779,N_20348);
xnor U23835 (N_23835,N_19970,N_18811);
and U23836 (N_23836,N_21141,N_19622);
or U23837 (N_23837,N_19717,N_21638);
and U23838 (N_23838,N_20486,N_19328);
xnor U23839 (N_23839,N_21739,N_20874);
nand U23840 (N_23840,N_19450,N_21470);
xnor U23841 (N_23841,N_21707,N_20547);
or U23842 (N_23842,N_20883,N_20214);
or U23843 (N_23843,N_20294,N_20897);
nor U23844 (N_23844,N_21610,N_21067);
nand U23845 (N_23845,N_21121,N_19360);
xnor U23846 (N_23846,N_20370,N_21790);
nor U23847 (N_23847,N_21751,N_21181);
or U23848 (N_23848,N_21731,N_19556);
nand U23849 (N_23849,N_19765,N_18802);
or U23850 (N_23850,N_20089,N_18916);
nand U23851 (N_23851,N_19163,N_19882);
nand U23852 (N_23852,N_21088,N_21395);
and U23853 (N_23853,N_20781,N_20740);
xnor U23854 (N_23854,N_20436,N_20176);
nor U23855 (N_23855,N_18796,N_19300);
xnor U23856 (N_23856,N_19506,N_19568);
and U23857 (N_23857,N_21400,N_20099);
nor U23858 (N_23858,N_20011,N_20673);
nor U23859 (N_23859,N_20759,N_20444);
nand U23860 (N_23860,N_20569,N_20730);
and U23861 (N_23861,N_20023,N_19028);
xnor U23862 (N_23862,N_19022,N_20243);
xor U23863 (N_23863,N_19221,N_20757);
nand U23864 (N_23864,N_18809,N_20296);
nor U23865 (N_23865,N_21064,N_19382);
xnor U23866 (N_23866,N_18894,N_21249);
nand U23867 (N_23867,N_19749,N_20234);
or U23868 (N_23868,N_20616,N_18776);
and U23869 (N_23869,N_20071,N_19592);
and U23870 (N_23870,N_21034,N_20751);
or U23871 (N_23871,N_20756,N_19240);
or U23872 (N_23872,N_20929,N_19574);
nand U23873 (N_23873,N_20643,N_21701);
xnor U23874 (N_23874,N_21484,N_20186);
or U23875 (N_23875,N_21441,N_20886);
nand U23876 (N_23876,N_20355,N_21659);
and U23877 (N_23877,N_20195,N_20941);
nor U23878 (N_23878,N_19521,N_19783);
and U23879 (N_23879,N_19783,N_19437);
nand U23880 (N_23880,N_19978,N_19365);
and U23881 (N_23881,N_21738,N_19391);
xnor U23882 (N_23882,N_20780,N_18962);
nor U23883 (N_23883,N_20583,N_21418);
xor U23884 (N_23884,N_20949,N_19720);
or U23885 (N_23885,N_20392,N_19272);
and U23886 (N_23886,N_21855,N_19486);
and U23887 (N_23887,N_20356,N_20520);
or U23888 (N_23888,N_20205,N_20464);
nor U23889 (N_23889,N_20870,N_20383);
and U23890 (N_23890,N_19579,N_19359);
nand U23891 (N_23891,N_21638,N_20341);
and U23892 (N_23892,N_20361,N_21846);
or U23893 (N_23893,N_20432,N_19394);
or U23894 (N_23894,N_18774,N_20211);
nor U23895 (N_23895,N_21585,N_20813);
or U23896 (N_23896,N_20131,N_19794);
nand U23897 (N_23897,N_19325,N_20256);
nor U23898 (N_23898,N_21096,N_21099);
xnor U23899 (N_23899,N_21364,N_21731);
and U23900 (N_23900,N_19947,N_19477);
nand U23901 (N_23901,N_21867,N_21155);
nor U23902 (N_23902,N_20391,N_18798);
nor U23903 (N_23903,N_21641,N_19848);
and U23904 (N_23904,N_19150,N_19934);
and U23905 (N_23905,N_20399,N_21726);
xnor U23906 (N_23906,N_21152,N_21055);
xnor U23907 (N_23907,N_20420,N_20472);
or U23908 (N_23908,N_20920,N_19999);
nor U23909 (N_23909,N_21068,N_19243);
and U23910 (N_23910,N_18996,N_20646);
nand U23911 (N_23911,N_20801,N_21132);
nor U23912 (N_23912,N_21003,N_18952);
nand U23913 (N_23913,N_20016,N_20376);
nor U23914 (N_23914,N_19223,N_20058);
nor U23915 (N_23915,N_20777,N_20114);
or U23916 (N_23916,N_19191,N_20283);
nand U23917 (N_23917,N_19906,N_19594);
xor U23918 (N_23918,N_20086,N_21152);
nand U23919 (N_23919,N_19437,N_19723);
nand U23920 (N_23920,N_20798,N_21751);
nor U23921 (N_23921,N_20064,N_21480);
and U23922 (N_23922,N_21250,N_19746);
xor U23923 (N_23923,N_20201,N_20542);
or U23924 (N_23924,N_21623,N_20277);
nand U23925 (N_23925,N_20037,N_21693);
xor U23926 (N_23926,N_21094,N_21323);
nand U23927 (N_23927,N_19302,N_19373);
or U23928 (N_23928,N_21761,N_19520);
xnor U23929 (N_23929,N_20869,N_20525);
nand U23930 (N_23930,N_18800,N_21009);
or U23931 (N_23931,N_21350,N_18982);
nand U23932 (N_23932,N_20131,N_19182);
or U23933 (N_23933,N_19272,N_20946);
xor U23934 (N_23934,N_19655,N_20118);
or U23935 (N_23935,N_21871,N_20969);
nor U23936 (N_23936,N_19194,N_20199);
xor U23937 (N_23937,N_19534,N_20950);
or U23938 (N_23938,N_21150,N_19415);
nand U23939 (N_23939,N_20645,N_21005);
xnor U23940 (N_23940,N_19416,N_21327);
nor U23941 (N_23941,N_20019,N_19661);
nor U23942 (N_23942,N_18836,N_19513);
nor U23943 (N_23943,N_19991,N_20461);
or U23944 (N_23944,N_19679,N_20907);
xnor U23945 (N_23945,N_19228,N_19316);
nor U23946 (N_23946,N_21584,N_21546);
nand U23947 (N_23947,N_19195,N_19105);
xnor U23948 (N_23948,N_19164,N_19759);
xor U23949 (N_23949,N_19548,N_18839);
xor U23950 (N_23950,N_19813,N_18760);
nor U23951 (N_23951,N_20513,N_20406);
nor U23952 (N_23952,N_19461,N_21645);
nor U23953 (N_23953,N_21555,N_19541);
xnor U23954 (N_23954,N_20956,N_21718);
and U23955 (N_23955,N_20869,N_21681);
nor U23956 (N_23956,N_21648,N_19353);
or U23957 (N_23957,N_19147,N_19840);
nand U23958 (N_23958,N_19977,N_19441);
nand U23959 (N_23959,N_19378,N_20270);
or U23960 (N_23960,N_21570,N_19063);
nand U23961 (N_23961,N_21324,N_18901);
or U23962 (N_23962,N_20487,N_20818);
nor U23963 (N_23963,N_21614,N_18823);
xnor U23964 (N_23964,N_21298,N_20961);
nand U23965 (N_23965,N_21122,N_20465);
nor U23966 (N_23966,N_20995,N_19043);
xor U23967 (N_23967,N_19700,N_20402);
xor U23968 (N_23968,N_18958,N_21134);
nand U23969 (N_23969,N_20192,N_19424);
nand U23970 (N_23970,N_18981,N_21309);
and U23971 (N_23971,N_19214,N_21704);
or U23972 (N_23972,N_20454,N_20585);
and U23973 (N_23973,N_19759,N_18890);
or U23974 (N_23974,N_21149,N_18904);
and U23975 (N_23975,N_21467,N_20734);
and U23976 (N_23976,N_21830,N_21600);
nor U23977 (N_23977,N_21601,N_19900);
and U23978 (N_23978,N_19674,N_20950);
nand U23979 (N_23979,N_20947,N_19788);
xnor U23980 (N_23980,N_20210,N_21091);
xor U23981 (N_23981,N_20961,N_21399);
xnor U23982 (N_23982,N_19172,N_19194);
nor U23983 (N_23983,N_20101,N_19197);
or U23984 (N_23984,N_21335,N_20648);
xor U23985 (N_23985,N_19014,N_21012);
and U23986 (N_23986,N_21098,N_20650);
nor U23987 (N_23987,N_19170,N_19175);
nor U23988 (N_23988,N_19661,N_21000);
nor U23989 (N_23989,N_21237,N_19352);
nand U23990 (N_23990,N_19263,N_19848);
or U23991 (N_23991,N_18988,N_19261);
and U23992 (N_23992,N_19394,N_19688);
xor U23993 (N_23993,N_20862,N_19817);
or U23994 (N_23994,N_20038,N_18997);
nand U23995 (N_23995,N_20651,N_20052);
nor U23996 (N_23996,N_21297,N_21036);
and U23997 (N_23997,N_20391,N_21370);
nand U23998 (N_23998,N_21440,N_21451);
or U23999 (N_23999,N_20233,N_20717);
or U24000 (N_24000,N_19530,N_21423);
and U24001 (N_24001,N_20691,N_20056);
and U24002 (N_24002,N_19353,N_19588);
nor U24003 (N_24003,N_21253,N_20129);
nand U24004 (N_24004,N_21193,N_21013);
nand U24005 (N_24005,N_20596,N_19120);
or U24006 (N_24006,N_19791,N_21186);
xor U24007 (N_24007,N_19265,N_18931);
nor U24008 (N_24008,N_19937,N_20261);
and U24009 (N_24009,N_20875,N_20037);
nand U24010 (N_24010,N_20441,N_19530);
nor U24011 (N_24011,N_19039,N_18769);
nor U24012 (N_24012,N_21787,N_20329);
or U24013 (N_24013,N_18841,N_21675);
nor U24014 (N_24014,N_21489,N_19296);
or U24015 (N_24015,N_20321,N_21035);
nand U24016 (N_24016,N_18970,N_20420);
or U24017 (N_24017,N_19859,N_18773);
nand U24018 (N_24018,N_21239,N_18920);
nor U24019 (N_24019,N_20608,N_21197);
nand U24020 (N_24020,N_19820,N_21497);
nand U24021 (N_24021,N_21513,N_19738);
nor U24022 (N_24022,N_21603,N_19946);
nand U24023 (N_24023,N_21163,N_19275);
xnor U24024 (N_24024,N_19263,N_21109);
nand U24025 (N_24025,N_18865,N_20052);
and U24026 (N_24026,N_21674,N_21503);
xor U24027 (N_24027,N_20980,N_21266);
or U24028 (N_24028,N_19379,N_21284);
nor U24029 (N_24029,N_21080,N_18971);
nor U24030 (N_24030,N_20648,N_19478);
or U24031 (N_24031,N_19794,N_19741);
nor U24032 (N_24032,N_20886,N_21571);
nor U24033 (N_24033,N_21613,N_20978);
or U24034 (N_24034,N_20229,N_20643);
nor U24035 (N_24035,N_19294,N_19729);
nor U24036 (N_24036,N_21116,N_19170);
xor U24037 (N_24037,N_19316,N_20125);
xnor U24038 (N_24038,N_20151,N_21258);
nor U24039 (N_24039,N_19488,N_21870);
nor U24040 (N_24040,N_18943,N_20489);
and U24041 (N_24041,N_21094,N_20001);
xor U24042 (N_24042,N_19009,N_20788);
nor U24043 (N_24043,N_21357,N_19757);
nand U24044 (N_24044,N_18876,N_18804);
xnor U24045 (N_24045,N_20127,N_21863);
or U24046 (N_24046,N_21771,N_21783);
or U24047 (N_24047,N_19239,N_19442);
nand U24048 (N_24048,N_21398,N_20401);
or U24049 (N_24049,N_21519,N_20667);
xor U24050 (N_24050,N_20646,N_20138);
nand U24051 (N_24051,N_19146,N_19115);
xnor U24052 (N_24052,N_19715,N_21036);
xor U24053 (N_24053,N_19420,N_19170);
nand U24054 (N_24054,N_21732,N_21607);
nand U24055 (N_24055,N_19862,N_20278);
or U24056 (N_24056,N_20181,N_20744);
nor U24057 (N_24057,N_20214,N_19114);
xnor U24058 (N_24058,N_19859,N_21030);
or U24059 (N_24059,N_20192,N_21439);
and U24060 (N_24060,N_20681,N_18866);
nand U24061 (N_24061,N_20254,N_20982);
and U24062 (N_24062,N_21122,N_20578);
nor U24063 (N_24063,N_18938,N_20530);
and U24064 (N_24064,N_19743,N_19065);
or U24065 (N_24065,N_20596,N_19842);
nor U24066 (N_24066,N_20292,N_19264);
xor U24067 (N_24067,N_19459,N_21771);
xnor U24068 (N_24068,N_20341,N_20034);
xnor U24069 (N_24069,N_19780,N_21181);
and U24070 (N_24070,N_19765,N_19511);
xor U24071 (N_24071,N_21759,N_21058);
nor U24072 (N_24072,N_19072,N_20853);
nor U24073 (N_24073,N_20698,N_20017);
xnor U24074 (N_24074,N_21707,N_19564);
or U24075 (N_24075,N_21118,N_18816);
or U24076 (N_24076,N_21546,N_19840);
nor U24077 (N_24077,N_21534,N_21549);
and U24078 (N_24078,N_19730,N_19789);
or U24079 (N_24079,N_21274,N_20027);
nand U24080 (N_24080,N_18926,N_19053);
xnor U24081 (N_24081,N_20194,N_20922);
nor U24082 (N_24082,N_20386,N_19962);
nand U24083 (N_24083,N_20840,N_21274);
nand U24084 (N_24084,N_21162,N_20536);
xnor U24085 (N_24085,N_18955,N_20808);
nor U24086 (N_24086,N_19132,N_19911);
nor U24087 (N_24087,N_20410,N_19030);
or U24088 (N_24088,N_18843,N_19440);
xor U24089 (N_24089,N_20763,N_21824);
or U24090 (N_24090,N_20056,N_19260);
and U24091 (N_24091,N_19174,N_19035);
xnor U24092 (N_24092,N_19182,N_21514);
xnor U24093 (N_24093,N_21171,N_20826);
nand U24094 (N_24094,N_20053,N_21312);
xnor U24095 (N_24095,N_21428,N_20747);
nand U24096 (N_24096,N_21616,N_19453);
nor U24097 (N_24097,N_19942,N_21191);
and U24098 (N_24098,N_21495,N_20284);
nor U24099 (N_24099,N_19169,N_20951);
or U24100 (N_24100,N_20263,N_19095);
nand U24101 (N_24101,N_21339,N_20424);
or U24102 (N_24102,N_21183,N_18815);
nand U24103 (N_24103,N_21087,N_21520);
and U24104 (N_24104,N_21495,N_21167);
xor U24105 (N_24105,N_20352,N_20774);
nand U24106 (N_24106,N_20854,N_21695);
nor U24107 (N_24107,N_21874,N_19587);
or U24108 (N_24108,N_20902,N_20304);
nor U24109 (N_24109,N_21146,N_20003);
and U24110 (N_24110,N_20167,N_21461);
and U24111 (N_24111,N_18865,N_20215);
nand U24112 (N_24112,N_20028,N_21313);
or U24113 (N_24113,N_21704,N_20077);
xor U24114 (N_24114,N_21730,N_21251);
xnor U24115 (N_24115,N_20390,N_19379);
and U24116 (N_24116,N_21398,N_20990);
and U24117 (N_24117,N_18891,N_19929);
nor U24118 (N_24118,N_19437,N_18956);
xor U24119 (N_24119,N_19000,N_19206);
or U24120 (N_24120,N_19741,N_20780);
xnor U24121 (N_24121,N_18841,N_19534);
nand U24122 (N_24122,N_19768,N_21195);
or U24123 (N_24123,N_19950,N_21236);
and U24124 (N_24124,N_20947,N_19825);
nor U24125 (N_24125,N_19100,N_21232);
xor U24126 (N_24126,N_19851,N_20923);
and U24127 (N_24127,N_21518,N_20106);
nand U24128 (N_24128,N_20347,N_21418);
nand U24129 (N_24129,N_19177,N_19557);
nor U24130 (N_24130,N_20326,N_19931);
or U24131 (N_24131,N_20653,N_18943);
xor U24132 (N_24132,N_19238,N_18784);
nor U24133 (N_24133,N_19301,N_21682);
nand U24134 (N_24134,N_20532,N_19640);
or U24135 (N_24135,N_20283,N_21559);
and U24136 (N_24136,N_20577,N_20114);
or U24137 (N_24137,N_20873,N_20303);
nand U24138 (N_24138,N_21275,N_21313);
nand U24139 (N_24139,N_19833,N_21621);
and U24140 (N_24140,N_19069,N_21012);
nand U24141 (N_24141,N_19238,N_19103);
and U24142 (N_24142,N_21358,N_21573);
xor U24143 (N_24143,N_19163,N_21511);
nand U24144 (N_24144,N_18974,N_20911);
xor U24145 (N_24145,N_20414,N_21123);
nor U24146 (N_24146,N_21099,N_19455);
and U24147 (N_24147,N_19874,N_19793);
nor U24148 (N_24148,N_21511,N_20894);
and U24149 (N_24149,N_19480,N_19893);
nand U24150 (N_24150,N_19319,N_20329);
nand U24151 (N_24151,N_21559,N_20791);
and U24152 (N_24152,N_20247,N_19374);
and U24153 (N_24153,N_18789,N_20038);
nand U24154 (N_24154,N_20564,N_20166);
nor U24155 (N_24155,N_19726,N_20359);
nand U24156 (N_24156,N_21326,N_21366);
nor U24157 (N_24157,N_20289,N_20632);
or U24158 (N_24158,N_21441,N_18846);
nand U24159 (N_24159,N_19481,N_21278);
and U24160 (N_24160,N_20814,N_19144);
xor U24161 (N_24161,N_18786,N_20585);
nor U24162 (N_24162,N_19854,N_19894);
or U24163 (N_24163,N_19377,N_21640);
and U24164 (N_24164,N_19757,N_20976);
and U24165 (N_24165,N_19027,N_21531);
and U24166 (N_24166,N_19732,N_21177);
nor U24167 (N_24167,N_20011,N_19393);
nand U24168 (N_24168,N_21764,N_20105);
nor U24169 (N_24169,N_19866,N_20752);
nor U24170 (N_24170,N_18857,N_19649);
and U24171 (N_24171,N_19296,N_18962);
nor U24172 (N_24172,N_19464,N_19604);
or U24173 (N_24173,N_21822,N_19969);
nand U24174 (N_24174,N_19909,N_20519);
xnor U24175 (N_24175,N_21534,N_20927);
or U24176 (N_24176,N_21680,N_19775);
nand U24177 (N_24177,N_21662,N_21074);
or U24178 (N_24178,N_20743,N_18886);
xor U24179 (N_24179,N_21078,N_19175);
xnor U24180 (N_24180,N_19118,N_19981);
and U24181 (N_24181,N_19970,N_21002);
nor U24182 (N_24182,N_19983,N_20048);
nor U24183 (N_24183,N_20293,N_18965);
xnor U24184 (N_24184,N_21199,N_19911);
xor U24185 (N_24185,N_19742,N_19059);
and U24186 (N_24186,N_21789,N_18762);
xor U24187 (N_24187,N_18824,N_18806);
or U24188 (N_24188,N_20195,N_20196);
and U24189 (N_24189,N_21288,N_19366);
or U24190 (N_24190,N_19324,N_19121);
or U24191 (N_24191,N_21415,N_21640);
or U24192 (N_24192,N_19383,N_18865);
nor U24193 (N_24193,N_19109,N_20116);
nand U24194 (N_24194,N_20848,N_18910);
xor U24195 (N_24195,N_19860,N_20337);
nand U24196 (N_24196,N_18975,N_21515);
nor U24197 (N_24197,N_21870,N_21787);
nor U24198 (N_24198,N_21530,N_21058);
or U24199 (N_24199,N_21292,N_20666);
xnor U24200 (N_24200,N_20388,N_19814);
and U24201 (N_24201,N_20080,N_19332);
nor U24202 (N_24202,N_21173,N_21181);
and U24203 (N_24203,N_20941,N_19630);
or U24204 (N_24204,N_20811,N_20853);
and U24205 (N_24205,N_21571,N_18907);
and U24206 (N_24206,N_21143,N_20172);
xor U24207 (N_24207,N_19150,N_20987);
nand U24208 (N_24208,N_21353,N_19293);
xnor U24209 (N_24209,N_19562,N_19435);
and U24210 (N_24210,N_20802,N_20121);
nor U24211 (N_24211,N_19053,N_21572);
or U24212 (N_24212,N_20289,N_19691);
nand U24213 (N_24213,N_21623,N_21370);
xnor U24214 (N_24214,N_19583,N_19236);
and U24215 (N_24215,N_21342,N_19517);
nand U24216 (N_24216,N_19969,N_19471);
xor U24217 (N_24217,N_21535,N_21456);
xnor U24218 (N_24218,N_20223,N_19099);
nand U24219 (N_24219,N_21804,N_19096);
and U24220 (N_24220,N_19795,N_20207);
and U24221 (N_24221,N_19887,N_20792);
and U24222 (N_24222,N_19210,N_19553);
and U24223 (N_24223,N_19073,N_21113);
and U24224 (N_24224,N_19961,N_21157);
nor U24225 (N_24225,N_18751,N_18860);
xnor U24226 (N_24226,N_21605,N_20707);
xor U24227 (N_24227,N_20352,N_19979);
and U24228 (N_24228,N_21065,N_21350);
nand U24229 (N_24229,N_21664,N_21804);
nor U24230 (N_24230,N_19559,N_21122);
xor U24231 (N_24231,N_19058,N_18798);
nor U24232 (N_24232,N_20455,N_20506);
nor U24233 (N_24233,N_21536,N_19278);
nand U24234 (N_24234,N_19355,N_20927);
nor U24235 (N_24235,N_21592,N_21668);
or U24236 (N_24236,N_19343,N_20786);
xor U24237 (N_24237,N_20853,N_20007);
or U24238 (N_24238,N_21840,N_20283);
xnor U24239 (N_24239,N_19083,N_19075);
xor U24240 (N_24240,N_20121,N_21572);
and U24241 (N_24241,N_20116,N_20399);
nand U24242 (N_24242,N_21616,N_20355);
or U24243 (N_24243,N_21708,N_20843);
and U24244 (N_24244,N_18780,N_21108);
xor U24245 (N_24245,N_19780,N_20899);
xnor U24246 (N_24246,N_21182,N_21793);
nand U24247 (N_24247,N_18750,N_19242);
nor U24248 (N_24248,N_21105,N_21066);
and U24249 (N_24249,N_21107,N_19375);
or U24250 (N_24250,N_21736,N_21096);
nand U24251 (N_24251,N_18998,N_21272);
xnor U24252 (N_24252,N_19187,N_21112);
xnor U24253 (N_24253,N_21248,N_19670);
xor U24254 (N_24254,N_20613,N_20383);
nand U24255 (N_24255,N_20995,N_19574);
and U24256 (N_24256,N_19675,N_20574);
nor U24257 (N_24257,N_20703,N_18756);
nand U24258 (N_24258,N_20438,N_19114);
nand U24259 (N_24259,N_19456,N_19193);
xnor U24260 (N_24260,N_20199,N_20071);
and U24261 (N_24261,N_20657,N_19429);
nor U24262 (N_24262,N_21115,N_21098);
nor U24263 (N_24263,N_20168,N_20527);
and U24264 (N_24264,N_21480,N_21491);
xor U24265 (N_24265,N_21574,N_21671);
nand U24266 (N_24266,N_20212,N_20166);
xor U24267 (N_24267,N_19645,N_19963);
xnor U24268 (N_24268,N_21621,N_21854);
xor U24269 (N_24269,N_21146,N_21031);
nand U24270 (N_24270,N_20128,N_20200);
nor U24271 (N_24271,N_21058,N_18816);
and U24272 (N_24272,N_19681,N_20607);
or U24273 (N_24273,N_21869,N_20638);
and U24274 (N_24274,N_21063,N_21089);
and U24275 (N_24275,N_21695,N_19720);
nor U24276 (N_24276,N_19278,N_19370);
or U24277 (N_24277,N_18849,N_18844);
and U24278 (N_24278,N_18888,N_21189);
and U24279 (N_24279,N_21809,N_19701);
and U24280 (N_24280,N_20364,N_20795);
nand U24281 (N_24281,N_20514,N_20278);
nor U24282 (N_24282,N_19772,N_18883);
nand U24283 (N_24283,N_19569,N_21359);
xor U24284 (N_24284,N_19760,N_20659);
nand U24285 (N_24285,N_21464,N_19319);
or U24286 (N_24286,N_18946,N_20693);
and U24287 (N_24287,N_21226,N_19193);
nor U24288 (N_24288,N_18845,N_20141);
and U24289 (N_24289,N_21455,N_18924);
or U24290 (N_24290,N_21696,N_19269);
nor U24291 (N_24291,N_21619,N_19231);
or U24292 (N_24292,N_19620,N_19446);
and U24293 (N_24293,N_19049,N_20281);
nand U24294 (N_24294,N_20473,N_21687);
or U24295 (N_24295,N_20691,N_19762);
nand U24296 (N_24296,N_21857,N_20473);
nor U24297 (N_24297,N_19224,N_21791);
nand U24298 (N_24298,N_21698,N_20316);
nand U24299 (N_24299,N_18974,N_21602);
and U24300 (N_24300,N_20007,N_20880);
and U24301 (N_24301,N_18810,N_19617);
nand U24302 (N_24302,N_21088,N_19889);
nand U24303 (N_24303,N_21703,N_21414);
nor U24304 (N_24304,N_20334,N_20077);
xor U24305 (N_24305,N_20709,N_18842);
xor U24306 (N_24306,N_21874,N_20067);
xnor U24307 (N_24307,N_18785,N_21226);
nand U24308 (N_24308,N_18936,N_19787);
and U24309 (N_24309,N_19535,N_21838);
nor U24310 (N_24310,N_19449,N_21592);
xnor U24311 (N_24311,N_20160,N_20185);
nand U24312 (N_24312,N_19945,N_20509);
nand U24313 (N_24313,N_21517,N_20470);
and U24314 (N_24314,N_19821,N_20489);
or U24315 (N_24315,N_19970,N_21420);
nor U24316 (N_24316,N_21043,N_19020);
xnor U24317 (N_24317,N_21770,N_20972);
nor U24318 (N_24318,N_21476,N_19186);
nor U24319 (N_24319,N_21338,N_20258);
nor U24320 (N_24320,N_21277,N_21683);
or U24321 (N_24321,N_21833,N_20363);
and U24322 (N_24322,N_20633,N_20752);
nand U24323 (N_24323,N_20831,N_20030);
nand U24324 (N_24324,N_19741,N_21199);
and U24325 (N_24325,N_19095,N_21814);
nor U24326 (N_24326,N_20352,N_20413);
or U24327 (N_24327,N_20400,N_19360);
xor U24328 (N_24328,N_20282,N_21492);
or U24329 (N_24329,N_19749,N_20382);
nand U24330 (N_24330,N_18958,N_19090);
xnor U24331 (N_24331,N_20848,N_20454);
nor U24332 (N_24332,N_19967,N_19178);
xor U24333 (N_24333,N_18982,N_20927);
xor U24334 (N_24334,N_20575,N_20393);
nand U24335 (N_24335,N_19608,N_20510);
nand U24336 (N_24336,N_21644,N_20152);
and U24337 (N_24337,N_21276,N_19210);
nor U24338 (N_24338,N_21029,N_19406);
xnor U24339 (N_24339,N_21001,N_19373);
or U24340 (N_24340,N_21276,N_19815);
xor U24341 (N_24341,N_19210,N_20539);
xor U24342 (N_24342,N_20277,N_20060);
nand U24343 (N_24343,N_20236,N_20099);
or U24344 (N_24344,N_21338,N_19215);
and U24345 (N_24345,N_20151,N_18948);
xnor U24346 (N_24346,N_18827,N_21640);
nor U24347 (N_24347,N_19897,N_19659);
nor U24348 (N_24348,N_21864,N_21700);
nand U24349 (N_24349,N_21023,N_19748);
and U24350 (N_24350,N_19879,N_21034);
nand U24351 (N_24351,N_21716,N_21667);
and U24352 (N_24352,N_21509,N_20570);
nand U24353 (N_24353,N_20390,N_20327);
nor U24354 (N_24354,N_19216,N_20625);
xnor U24355 (N_24355,N_20444,N_19883);
or U24356 (N_24356,N_20923,N_20111);
nand U24357 (N_24357,N_18772,N_21739);
xor U24358 (N_24358,N_19026,N_20481);
xnor U24359 (N_24359,N_19657,N_21130);
and U24360 (N_24360,N_20667,N_21298);
nor U24361 (N_24361,N_19243,N_21749);
and U24362 (N_24362,N_21211,N_19903);
nand U24363 (N_24363,N_20251,N_18957);
or U24364 (N_24364,N_19765,N_21338);
or U24365 (N_24365,N_21224,N_21341);
xor U24366 (N_24366,N_20862,N_20205);
nand U24367 (N_24367,N_21759,N_20990);
and U24368 (N_24368,N_21519,N_20530);
xor U24369 (N_24369,N_20198,N_20370);
nor U24370 (N_24370,N_19531,N_20282);
nand U24371 (N_24371,N_21487,N_20195);
xor U24372 (N_24372,N_19677,N_21874);
and U24373 (N_24373,N_19396,N_21386);
xor U24374 (N_24374,N_19015,N_20136);
or U24375 (N_24375,N_20993,N_20507);
nand U24376 (N_24376,N_20526,N_21095);
xor U24377 (N_24377,N_19472,N_20616);
or U24378 (N_24378,N_19660,N_19160);
nor U24379 (N_24379,N_21398,N_21799);
or U24380 (N_24380,N_20090,N_18963);
and U24381 (N_24381,N_19561,N_19858);
or U24382 (N_24382,N_21842,N_21308);
and U24383 (N_24383,N_20696,N_19792);
nand U24384 (N_24384,N_21138,N_20704);
or U24385 (N_24385,N_19369,N_21489);
and U24386 (N_24386,N_20792,N_21028);
nand U24387 (N_24387,N_19259,N_21192);
nor U24388 (N_24388,N_20732,N_21118);
xnor U24389 (N_24389,N_21749,N_21420);
nand U24390 (N_24390,N_20804,N_18909);
and U24391 (N_24391,N_21610,N_21144);
or U24392 (N_24392,N_20872,N_20397);
nor U24393 (N_24393,N_21665,N_18758);
or U24394 (N_24394,N_19225,N_20671);
and U24395 (N_24395,N_20340,N_19912);
xnor U24396 (N_24396,N_19653,N_20098);
nor U24397 (N_24397,N_19813,N_21660);
or U24398 (N_24398,N_20126,N_21209);
nand U24399 (N_24399,N_18757,N_19802);
nor U24400 (N_24400,N_20133,N_18857);
and U24401 (N_24401,N_20794,N_20242);
and U24402 (N_24402,N_20950,N_21244);
nand U24403 (N_24403,N_19788,N_20201);
xor U24404 (N_24404,N_20562,N_18923);
xor U24405 (N_24405,N_19317,N_19104);
nand U24406 (N_24406,N_20614,N_20203);
and U24407 (N_24407,N_19093,N_19968);
nor U24408 (N_24408,N_20358,N_18920);
nor U24409 (N_24409,N_20455,N_21623);
nand U24410 (N_24410,N_18975,N_20784);
nand U24411 (N_24411,N_21184,N_19257);
or U24412 (N_24412,N_21702,N_21219);
nor U24413 (N_24413,N_20513,N_21857);
nor U24414 (N_24414,N_21151,N_21844);
nand U24415 (N_24415,N_19233,N_21479);
xor U24416 (N_24416,N_21153,N_19517);
and U24417 (N_24417,N_19351,N_18825);
and U24418 (N_24418,N_19503,N_19451);
xnor U24419 (N_24419,N_21052,N_18760);
nor U24420 (N_24420,N_19810,N_21716);
nor U24421 (N_24421,N_18932,N_20239);
nor U24422 (N_24422,N_20239,N_21197);
nand U24423 (N_24423,N_18949,N_21212);
nor U24424 (N_24424,N_19315,N_20113);
or U24425 (N_24425,N_20701,N_19095);
or U24426 (N_24426,N_19931,N_20570);
and U24427 (N_24427,N_21675,N_20087);
and U24428 (N_24428,N_19237,N_18764);
xor U24429 (N_24429,N_20806,N_20587);
xor U24430 (N_24430,N_21092,N_21409);
or U24431 (N_24431,N_19869,N_20102);
or U24432 (N_24432,N_20610,N_21627);
nor U24433 (N_24433,N_20744,N_21350);
or U24434 (N_24434,N_20178,N_19523);
or U24435 (N_24435,N_20959,N_20463);
and U24436 (N_24436,N_20177,N_21134);
nand U24437 (N_24437,N_20392,N_21837);
nand U24438 (N_24438,N_20574,N_20604);
xor U24439 (N_24439,N_21426,N_20054);
xor U24440 (N_24440,N_21749,N_19893);
and U24441 (N_24441,N_21476,N_21621);
xor U24442 (N_24442,N_21225,N_20784);
xnor U24443 (N_24443,N_21383,N_19104);
xor U24444 (N_24444,N_20739,N_21283);
nor U24445 (N_24445,N_19818,N_19503);
xnor U24446 (N_24446,N_20328,N_20380);
xnor U24447 (N_24447,N_21583,N_20475);
and U24448 (N_24448,N_21274,N_20359);
nand U24449 (N_24449,N_20593,N_20083);
nand U24450 (N_24450,N_18954,N_21853);
or U24451 (N_24451,N_20295,N_18763);
or U24452 (N_24452,N_19115,N_19712);
nor U24453 (N_24453,N_21083,N_19438);
nor U24454 (N_24454,N_20423,N_20781);
or U24455 (N_24455,N_20326,N_20937);
or U24456 (N_24456,N_18840,N_21194);
xnor U24457 (N_24457,N_19300,N_20773);
or U24458 (N_24458,N_19517,N_21706);
or U24459 (N_24459,N_20994,N_19906);
and U24460 (N_24460,N_20434,N_19281);
nor U24461 (N_24461,N_19658,N_20754);
nor U24462 (N_24462,N_20632,N_19122);
or U24463 (N_24463,N_21643,N_21244);
xor U24464 (N_24464,N_21335,N_21377);
xnor U24465 (N_24465,N_19154,N_21694);
nor U24466 (N_24466,N_20263,N_19890);
nand U24467 (N_24467,N_20919,N_21087);
nor U24468 (N_24468,N_19357,N_20437);
xor U24469 (N_24469,N_19633,N_20711);
or U24470 (N_24470,N_21808,N_18930);
and U24471 (N_24471,N_19757,N_18947);
or U24472 (N_24472,N_21467,N_21171);
and U24473 (N_24473,N_18859,N_19721);
nand U24474 (N_24474,N_20231,N_21805);
nand U24475 (N_24475,N_19209,N_20785);
or U24476 (N_24476,N_20698,N_19900);
nor U24477 (N_24477,N_19163,N_19094);
nor U24478 (N_24478,N_19965,N_20273);
xnor U24479 (N_24479,N_20011,N_19579);
and U24480 (N_24480,N_19320,N_19080);
and U24481 (N_24481,N_21096,N_21217);
and U24482 (N_24482,N_19002,N_21357);
xor U24483 (N_24483,N_19537,N_20893);
xnor U24484 (N_24484,N_20727,N_20512);
or U24485 (N_24485,N_20277,N_20638);
nand U24486 (N_24486,N_21071,N_19088);
or U24487 (N_24487,N_19524,N_20993);
nand U24488 (N_24488,N_19050,N_21688);
xor U24489 (N_24489,N_21488,N_20645);
xor U24490 (N_24490,N_20160,N_21227);
nand U24491 (N_24491,N_19779,N_18832);
nor U24492 (N_24492,N_19464,N_21705);
nand U24493 (N_24493,N_19551,N_21350);
nand U24494 (N_24494,N_21873,N_20622);
nand U24495 (N_24495,N_20081,N_21012);
nand U24496 (N_24496,N_19366,N_19015);
nor U24497 (N_24497,N_21816,N_19379);
and U24498 (N_24498,N_19789,N_21403);
xnor U24499 (N_24499,N_19895,N_19378);
xnor U24500 (N_24500,N_21124,N_19651);
or U24501 (N_24501,N_21572,N_20167);
xnor U24502 (N_24502,N_21706,N_21554);
and U24503 (N_24503,N_19294,N_19470);
xor U24504 (N_24504,N_19192,N_19620);
and U24505 (N_24505,N_20939,N_20878);
nand U24506 (N_24506,N_21263,N_21713);
xnor U24507 (N_24507,N_21646,N_20389);
nor U24508 (N_24508,N_20617,N_20271);
nand U24509 (N_24509,N_20148,N_20342);
and U24510 (N_24510,N_21803,N_20598);
or U24511 (N_24511,N_21836,N_19056);
or U24512 (N_24512,N_20035,N_21450);
nor U24513 (N_24513,N_21513,N_19372);
nor U24514 (N_24514,N_21306,N_21057);
nand U24515 (N_24515,N_21076,N_20774);
or U24516 (N_24516,N_21828,N_20619);
or U24517 (N_24517,N_19944,N_20366);
xnor U24518 (N_24518,N_20718,N_20204);
and U24519 (N_24519,N_21853,N_21639);
xnor U24520 (N_24520,N_19799,N_19562);
nand U24521 (N_24521,N_20524,N_19401);
and U24522 (N_24522,N_20826,N_19425);
xor U24523 (N_24523,N_19614,N_18759);
nor U24524 (N_24524,N_20516,N_18804);
xor U24525 (N_24525,N_20014,N_21253);
nor U24526 (N_24526,N_18982,N_21109);
nor U24527 (N_24527,N_19433,N_21656);
nand U24528 (N_24528,N_19435,N_21099);
nor U24529 (N_24529,N_19940,N_19991);
nor U24530 (N_24530,N_20182,N_19507);
or U24531 (N_24531,N_20387,N_20449);
nand U24532 (N_24532,N_18992,N_20206);
and U24533 (N_24533,N_19836,N_18784);
nand U24534 (N_24534,N_21848,N_20602);
xnor U24535 (N_24535,N_19343,N_19414);
and U24536 (N_24536,N_21022,N_19374);
or U24537 (N_24537,N_20853,N_20270);
nand U24538 (N_24538,N_18889,N_19757);
xor U24539 (N_24539,N_20190,N_19769);
nor U24540 (N_24540,N_19182,N_19792);
and U24541 (N_24541,N_18752,N_21871);
or U24542 (N_24542,N_19985,N_19639);
or U24543 (N_24543,N_20123,N_19047);
and U24544 (N_24544,N_20596,N_19845);
nor U24545 (N_24545,N_19595,N_20683);
and U24546 (N_24546,N_19802,N_18786);
nor U24547 (N_24547,N_21775,N_21794);
nor U24548 (N_24548,N_18784,N_20700);
nand U24549 (N_24549,N_20382,N_21683);
xor U24550 (N_24550,N_19841,N_19534);
nor U24551 (N_24551,N_18849,N_18902);
nand U24552 (N_24552,N_19102,N_19552);
or U24553 (N_24553,N_21229,N_21667);
nand U24554 (N_24554,N_21213,N_18965);
or U24555 (N_24555,N_20213,N_19130);
and U24556 (N_24556,N_20411,N_20939);
nor U24557 (N_24557,N_19105,N_19540);
nor U24558 (N_24558,N_21228,N_20561);
nor U24559 (N_24559,N_19720,N_19150);
nor U24560 (N_24560,N_21444,N_20748);
or U24561 (N_24561,N_19993,N_20826);
or U24562 (N_24562,N_19086,N_19718);
nor U24563 (N_24563,N_21782,N_21637);
and U24564 (N_24564,N_18764,N_19703);
or U24565 (N_24565,N_19134,N_20033);
or U24566 (N_24566,N_19536,N_19638);
nor U24567 (N_24567,N_21855,N_19006);
xor U24568 (N_24568,N_18923,N_18875);
or U24569 (N_24569,N_19154,N_18782);
nor U24570 (N_24570,N_19253,N_21668);
nand U24571 (N_24571,N_18758,N_20903);
and U24572 (N_24572,N_21760,N_20858);
or U24573 (N_24573,N_19271,N_18796);
nor U24574 (N_24574,N_21057,N_20958);
xnor U24575 (N_24575,N_18914,N_21873);
nand U24576 (N_24576,N_21777,N_19830);
nor U24577 (N_24577,N_20043,N_19219);
and U24578 (N_24578,N_21081,N_20251);
nand U24579 (N_24579,N_19232,N_20693);
nor U24580 (N_24580,N_19421,N_18849);
or U24581 (N_24581,N_21116,N_21664);
nand U24582 (N_24582,N_21221,N_21641);
xnor U24583 (N_24583,N_19746,N_20263);
or U24584 (N_24584,N_21652,N_21816);
or U24585 (N_24585,N_21837,N_19946);
nand U24586 (N_24586,N_19231,N_20690);
nor U24587 (N_24587,N_21407,N_19007);
or U24588 (N_24588,N_20659,N_20063);
nor U24589 (N_24589,N_20094,N_20522);
nand U24590 (N_24590,N_19770,N_18991);
and U24591 (N_24591,N_20230,N_21550);
or U24592 (N_24592,N_20254,N_21223);
or U24593 (N_24593,N_19316,N_19682);
nor U24594 (N_24594,N_21107,N_19181);
or U24595 (N_24595,N_19046,N_19699);
nor U24596 (N_24596,N_19228,N_20067);
and U24597 (N_24597,N_21641,N_19381);
nand U24598 (N_24598,N_19848,N_21426);
and U24599 (N_24599,N_19862,N_21458);
nand U24600 (N_24600,N_20230,N_18956);
nor U24601 (N_24601,N_19238,N_21581);
and U24602 (N_24602,N_20396,N_19751);
nand U24603 (N_24603,N_21147,N_19416);
xnor U24604 (N_24604,N_18881,N_19234);
nor U24605 (N_24605,N_18878,N_21812);
and U24606 (N_24606,N_20472,N_21502);
nor U24607 (N_24607,N_20956,N_18900);
xnor U24608 (N_24608,N_21730,N_21088);
xnor U24609 (N_24609,N_18807,N_19479);
nand U24610 (N_24610,N_19981,N_19931);
xnor U24611 (N_24611,N_18818,N_20462);
xor U24612 (N_24612,N_20900,N_19674);
nand U24613 (N_24613,N_21667,N_18978);
xnor U24614 (N_24614,N_19804,N_21845);
and U24615 (N_24615,N_20580,N_18850);
nand U24616 (N_24616,N_20821,N_19997);
xor U24617 (N_24617,N_21160,N_21534);
and U24618 (N_24618,N_19522,N_19367);
nand U24619 (N_24619,N_18858,N_18947);
nor U24620 (N_24620,N_21503,N_19956);
or U24621 (N_24621,N_19162,N_20012);
nand U24622 (N_24622,N_20514,N_19412);
or U24623 (N_24623,N_19896,N_20937);
nand U24624 (N_24624,N_19498,N_19364);
xnor U24625 (N_24625,N_20979,N_19576);
xor U24626 (N_24626,N_20543,N_20430);
xor U24627 (N_24627,N_19130,N_20061);
and U24628 (N_24628,N_20907,N_20505);
xnor U24629 (N_24629,N_20545,N_20746);
or U24630 (N_24630,N_21423,N_19424);
xnor U24631 (N_24631,N_21013,N_20183);
xnor U24632 (N_24632,N_18893,N_19091);
and U24633 (N_24633,N_21871,N_20810);
and U24634 (N_24634,N_21369,N_21855);
nand U24635 (N_24635,N_20343,N_19369);
xor U24636 (N_24636,N_20923,N_19426);
nand U24637 (N_24637,N_19679,N_19801);
xnor U24638 (N_24638,N_20257,N_21419);
xnor U24639 (N_24639,N_19180,N_21843);
or U24640 (N_24640,N_20990,N_19244);
nor U24641 (N_24641,N_19171,N_20278);
and U24642 (N_24642,N_20455,N_19681);
nor U24643 (N_24643,N_20296,N_20689);
xnor U24644 (N_24644,N_19283,N_21350);
nor U24645 (N_24645,N_18786,N_20819);
xor U24646 (N_24646,N_19413,N_19460);
xnor U24647 (N_24647,N_21813,N_21023);
nand U24648 (N_24648,N_20957,N_20351);
xnor U24649 (N_24649,N_20800,N_18988);
and U24650 (N_24650,N_21213,N_19956);
or U24651 (N_24651,N_21138,N_21612);
xnor U24652 (N_24652,N_20221,N_19884);
and U24653 (N_24653,N_20740,N_19544);
or U24654 (N_24654,N_19732,N_19106);
xor U24655 (N_24655,N_21399,N_20574);
xnor U24656 (N_24656,N_20015,N_21150);
nand U24657 (N_24657,N_18856,N_21275);
nor U24658 (N_24658,N_19035,N_19079);
nand U24659 (N_24659,N_18914,N_19002);
xnor U24660 (N_24660,N_21257,N_21391);
nor U24661 (N_24661,N_19272,N_19936);
or U24662 (N_24662,N_19340,N_20996);
and U24663 (N_24663,N_19007,N_19175);
xor U24664 (N_24664,N_19283,N_21624);
or U24665 (N_24665,N_19666,N_21210);
and U24666 (N_24666,N_21734,N_20407);
and U24667 (N_24667,N_19112,N_19026);
or U24668 (N_24668,N_21207,N_20313);
nor U24669 (N_24669,N_19717,N_21067);
xnor U24670 (N_24670,N_20714,N_20882);
and U24671 (N_24671,N_18850,N_19946);
or U24672 (N_24672,N_21435,N_21576);
or U24673 (N_24673,N_21132,N_20761);
and U24674 (N_24674,N_18933,N_21820);
nor U24675 (N_24675,N_19106,N_21658);
nor U24676 (N_24676,N_20337,N_19002);
xnor U24677 (N_24677,N_21414,N_20251);
and U24678 (N_24678,N_19790,N_21245);
nand U24679 (N_24679,N_21129,N_21791);
or U24680 (N_24680,N_20308,N_19934);
and U24681 (N_24681,N_21433,N_19226);
or U24682 (N_24682,N_18927,N_20732);
nor U24683 (N_24683,N_20389,N_20197);
nand U24684 (N_24684,N_21816,N_21503);
xnor U24685 (N_24685,N_18865,N_20561);
nor U24686 (N_24686,N_21291,N_19570);
nand U24687 (N_24687,N_19306,N_20111);
or U24688 (N_24688,N_18986,N_19525);
nor U24689 (N_24689,N_19752,N_19468);
or U24690 (N_24690,N_19764,N_19696);
xor U24691 (N_24691,N_18823,N_20557);
nor U24692 (N_24692,N_20054,N_18927);
nand U24693 (N_24693,N_19041,N_19515);
xor U24694 (N_24694,N_20774,N_20351);
nor U24695 (N_24695,N_20593,N_18928);
and U24696 (N_24696,N_21408,N_20913);
nand U24697 (N_24697,N_21561,N_19194);
or U24698 (N_24698,N_19395,N_20635);
nor U24699 (N_24699,N_19234,N_21388);
or U24700 (N_24700,N_21122,N_19092);
and U24701 (N_24701,N_20536,N_19563);
nor U24702 (N_24702,N_19437,N_20327);
nand U24703 (N_24703,N_20775,N_20494);
or U24704 (N_24704,N_20997,N_19975);
or U24705 (N_24705,N_19814,N_21832);
xor U24706 (N_24706,N_19585,N_19561);
xor U24707 (N_24707,N_19718,N_21762);
or U24708 (N_24708,N_19600,N_18910);
nand U24709 (N_24709,N_19053,N_21631);
nor U24710 (N_24710,N_21556,N_18770);
nor U24711 (N_24711,N_19490,N_21801);
nor U24712 (N_24712,N_19051,N_19204);
or U24713 (N_24713,N_19738,N_20531);
nor U24714 (N_24714,N_20036,N_20714);
and U24715 (N_24715,N_20109,N_20007);
and U24716 (N_24716,N_20900,N_21386);
or U24717 (N_24717,N_20386,N_19533);
and U24718 (N_24718,N_21500,N_19279);
xor U24719 (N_24719,N_18906,N_19717);
xor U24720 (N_24720,N_19097,N_21710);
or U24721 (N_24721,N_19583,N_18842);
xnor U24722 (N_24722,N_20786,N_21655);
or U24723 (N_24723,N_19422,N_21128);
nor U24724 (N_24724,N_21306,N_19265);
nor U24725 (N_24725,N_20841,N_21244);
nor U24726 (N_24726,N_20409,N_20941);
nand U24727 (N_24727,N_20058,N_18765);
and U24728 (N_24728,N_19210,N_21142);
and U24729 (N_24729,N_20408,N_18864);
or U24730 (N_24730,N_18979,N_21234);
and U24731 (N_24731,N_21263,N_20971);
or U24732 (N_24732,N_20942,N_20229);
nor U24733 (N_24733,N_19095,N_19628);
nand U24734 (N_24734,N_19649,N_21495);
xnor U24735 (N_24735,N_19104,N_19927);
or U24736 (N_24736,N_21568,N_20204);
and U24737 (N_24737,N_19655,N_19288);
xor U24738 (N_24738,N_20024,N_20348);
nor U24739 (N_24739,N_20650,N_19492);
and U24740 (N_24740,N_21193,N_21801);
and U24741 (N_24741,N_21090,N_19536);
nor U24742 (N_24742,N_21117,N_20336);
or U24743 (N_24743,N_20046,N_19153);
and U24744 (N_24744,N_20962,N_19749);
and U24745 (N_24745,N_21257,N_19039);
nor U24746 (N_24746,N_20606,N_20394);
nor U24747 (N_24747,N_19754,N_20033);
or U24748 (N_24748,N_21726,N_20248);
xnor U24749 (N_24749,N_20397,N_19603);
and U24750 (N_24750,N_19757,N_18852);
nor U24751 (N_24751,N_18985,N_20305);
nand U24752 (N_24752,N_20628,N_21685);
xor U24753 (N_24753,N_21576,N_18931);
and U24754 (N_24754,N_21381,N_20249);
nand U24755 (N_24755,N_18752,N_20031);
or U24756 (N_24756,N_21184,N_20089);
xor U24757 (N_24757,N_18946,N_21580);
nand U24758 (N_24758,N_19359,N_20817);
or U24759 (N_24759,N_20146,N_19591);
and U24760 (N_24760,N_19736,N_21507);
or U24761 (N_24761,N_20163,N_21388);
nor U24762 (N_24762,N_20638,N_20002);
nor U24763 (N_24763,N_21290,N_20861);
xnor U24764 (N_24764,N_19519,N_19754);
xor U24765 (N_24765,N_20187,N_19083);
nand U24766 (N_24766,N_21611,N_19989);
xnor U24767 (N_24767,N_21785,N_19473);
nor U24768 (N_24768,N_21636,N_19563);
and U24769 (N_24769,N_19987,N_21019);
or U24770 (N_24770,N_20990,N_21429);
nand U24771 (N_24771,N_21367,N_19769);
and U24772 (N_24772,N_21267,N_21573);
nand U24773 (N_24773,N_19991,N_20333);
xnor U24774 (N_24774,N_21528,N_19360);
nand U24775 (N_24775,N_21032,N_20726);
nor U24776 (N_24776,N_20599,N_20947);
nor U24777 (N_24777,N_19842,N_21738);
nor U24778 (N_24778,N_20577,N_20005);
nand U24779 (N_24779,N_21022,N_20417);
nand U24780 (N_24780,N_21151,N_21508);
nand U24781 (N_24781,N_21536,N_21273);
or U24782 (N_24782,N_21859,N_21207);
nand U24783 (N_24783,N_21392,N_19408);
nor U24784 (N_24784,N_19855,N_19010);
and U24785 (N_24785,N_20204,N_20660);
nand U24786 (N_24786,N_19875,N_19196);
or U24787 (N_24787,N_21576,N_21535);
or U24788 (N_24788,N_18832,N_20963);
and U24789 (N_24789,N_19039,N_21260);
nand U24790 (N_24790,N_19501,N_20461);
xnor U24791 (N_24791,N_20075,N_20891);
xor U24792 (N_24792,N_21345,N_19471);
nand U24793 (N_24793,N_19491,N_21453);
nand U24794 (N_24794,N_20174,N_20981);
and U24795 (N_24795,N_20213,N_19070);
or U24796 (N_24796,N_20529,N_20812);
nand U24797 (N_24797,N_20282,N_21813);
xor U24798 (N_24798,N_18965,N_21594);
or U24799 (N_24799,N_20323,N_21367);
and U24800 (N_24800,N_20035,N_18758);
nor U24801 (N_24801,N_19501,N_18789);
nand U24802 (N_24802,N_19790,N_20661);
xor U24803 (N_24803,N_21763,N_18831);
or U24804 (N_24804,N_21855,N_21227);
or U24805 (N_24805,N_21109,N_20736);
or U24806 (N_24806,N_18889,N_18972);
nor U24807 (N_24807,N_21606,N_20772);
nor U24808 (N_24808,N_19658,N_18823);
xor U24809 (N_24809,N_18995,N_19802);
or U24810 (N_24810,N_19596,N_21726);
nand U24811 (N_24811,N_20968,N_20977);
nor U24812 (N_24812,N_21382,N_19463);
xor U24813 (N_24813,N_21725,N_20947);
or U24814 (N_24814,N_19097,N_19148);
nor U24815 (N_24815,N_19714,N_19030);
nor U24816 (N_24816,N_19247,N_19821);
and U24817 (N_24817,N_20067,N_20415);
or U24818 (N_24818,N_18781,N_20247);
nor U24819 (N_24819,N_19180,N_21468);
xor U24820 (N_24820,N_21390,N_19016);
xnor U24821 (N_24821,N_19342,N_19320);
and U24822 (N_24822,N_20777,N_19882);
nand U24823 (N_24823,N_18909,N_19784);
xor U24824 (N_24824,N_19904,N_21002);
nand U24825 (N_24825,N_20198,N_20616);
nor U24826 (N_24826,N_20915,N_19731);
or U24827 (N_24827,N_18957,N_21216);
nor U24828 (N_24828,N_19627,N_19886);
xor U24829 (N_24829,N_20398,N_21028);
and U24830 (N_24830,N_21271,N_21165);
nand U24831 (N_24831,N_20641,N_20891);
nand U24832 (N_24832,N_20281,N_20584);
or U24833 (N_24833,N_19232,N_19687);
nand U24834 (N_24834,N_19466,N_21719);
xnor U24835 (N_24835,N_20864,N_19951);
nand U24836 (N_24836,N_20014,N_21222);
xor U24837 (N_24837,N_19316,N_19289);
and U24838 (N_24838,N_19404,N_19548);
nand U24839 (N_24839,N_20806,N_20931);
nand U24840 (N_24840,N_20322,N_18976);
nand U24841 (N_24841,N_18769,N_21472);
nor U24842 (N_24842,N_21706,N_18960);
or U24843 (N_24843,N_21508,N_19769);
or U24844 (N_24844,N_19084,N_19812);
nand U24845 (N_24845,N_20737,N_19133);
nor U24846 (N_24846,N_19672,N_21779);
or U24847 (N_24847,N_21730,N_19900);
and U24848 (N_24848,N_21676,N_21422);
xor U24849 (N_24849,N_21090,N_21317);
or U24850 (N_24850,N_20898,N_21815);
xnor U24851 (N_24851,N_19484,N_20629);
xor U24852 (N_24852,N_18869,N_21327);
nand U24853 (N_24853,N_21450,N_19156);
xnor U24854 (N_24854,N_19684,N_18986);
and U24855 (N_24855,N_20622,N_18896);
xnor U24856 (N_24856,N_20270,N_21215);
nand U24857 (N_24857,N_19418,N_19958);
nand U24858 (N_24858,N_21830,N_18937);
xnor U24859 (N_24859,N_21541,N_20953);
nand U24860 (N_24860,N_19841,N_20876);
or U24861 (N_24861,N_18969,N_19252);
nand U24862 (N_24862,N_19217,N_21724);
or U24863 (N_24863,N_18968,N_21809);
nand U24864 (N_24864,N_19163,N_20826);
and U24865 (N_24865,N_20882,N_18951);
xor U24866 (N_24866,N_19887,N_20822);
and U24867 (N_24867,N_21118,N_19871);
nor U24868 (N_24868,N_21342,N_20119);
or U24869 (N_24869,N_20902,N_19574);
nor U24870 (N_24870,N_20488,N_20268);
nor U24871 (N_24871,N_20510,N_20001);
and U24872 (N_24872,N_19908,N_19818);
and U24873 (N_24873,N_20637,N_19044);
or U24874 (N_24874,N_20138,N_21313);
nand U24875 (N_24875,N_19474,N_19097);
nand U24876 (N_24876,N_20497,N_20944);
and U24877 (N_24877,N_19518,N_19152);
and U24878 (N_24878,N_20766,N_20220);
nand U24879 (N_24879,N_21311,N_19283);
nor U24880 (N_24880,N_20362,N_19702);
xor U24881 (N_24881,N_20725,N_21585);
or U24882 (N_24882,N_19952,N_19135);
or U24883 (N_24883,N_20141,N_21400);
xor U24884 (N_24884,N_19026,N_19881);
xor U24885 (N_24885,N_19441,N_19561);
nor U24886 (N_24886,N_20566,N_19769);
nor U24887 (N_24887,N_20892,N_19559);
xnor U24888 (N_24888,N_18944,N_20231);
and U24889 (N_24889,N_19186,N_21711);
xor U24890 (N_24890,N_21549,N_21222);
or U24891 (N_24891,N_19647,N_18880);
xnor U24892 (N_24892,N_20924,N_19352);
xor U24893 (N_24893,N_19126,N_21651);
and U24894 (N_24894,N_19401,N_19603);
nand U24895 (N_24895,N_20384,N_20975);
or U24896 (N_24896,N_19747,N_19365);
or U24897 (N_24897,N_18972,N_19910);
and U24898 (N_24898,N_19409,N_20846);
nor U24899 (N_24899,N_20479,N_21703);
nor U24900 (N_24900,N_20735,N_20432);
and U24901 (N_24901,N_19509,N_18782);
or U24902 (N_24902,N_21836,N_18844);
xor U24903 (N_24903,N_19057,N_20591);
nor U24904 (N_24904,N_20127,N_20716);
and U24905 (N_24905,N_19129,N_20902);
nand U24906 (N_24906,N_20760,N_20478);
and U24907 (N_24907,N_20438,N_21720);
xnor U24908 (N_24908,N_20173,N_21468);
xor U24909 (N_24909,N_19376,N_21487);
nor U24910 (N_24910,N_21166,N_21390);
or U24911 (N_24911,N_20256,N_19584);
nor U24912 (N_24912,N_20460,N_19908);
or U24913 (N_24913,N_18948,N_19036);
nand U24914 (N_24914,N_20443,N_21269);
and U24915 (N_24915,N_18974,N_19408);
xor U24916 (N_24916,N_19059,N_20879);
xnor U24917 (N_24917,N_20376,N_21810);
or U24918 (N_24918,N_19030,N_20136);
or U24919 (N_24919,N_21504,N_18883);
nor U24920 (N_24920,N_19761,N_20413);
and U24921 (N_24921,N_18869,N_19986);
or U24922 (N_24922,N_20529,N_21492);
nor U24923 (N_24923,N_19463,N_21468);
nor U24924 (N_24924,N_19261,N_19672);
xnor U24925 (N_24925,N_20690,N_20327);
nor U24926 (N_24926,N_21799,N_19052);
nand U24927 (N_24927,N_19082,N_21544);
or U24928 (N_24928,N_19402,N_19540);
or U24929 (N_24929,N_19336,N_19120);
or U24930 (N_24930,N_20943,N_21379);
nor U24931 (N_24931,N_19002,N_19115);
and U24932 (N_24932,N_20254,N_21142);
xnor U24933 (N_24933,N_19198,N_19745);
or U24934 (N_24934,N_20520,N_18753);
nand U24935 (N_24935,N_19327,N_21721);
nand U24936 (N_24936,N_20236,N_19553);
xor U24937 (N_24937,N_21083,N_20722);
or U24938 (N_24938,N_20003,N_18961);
xor U24939 (N_24939,N_20862,N_20397);
nand U24940 (N_24940,N_20456,N_20503);
nor U24941 (N_24941,N_21616,N_19331);
nor U24942 (N_24942,N_20390,N_20020);
nor U24943 (N_24943,N_20850,N_20877);
xor U24944 (N_24944,N_20642,N_19187);
or U24945 (N_24945,N_21775,N_21800);
xor U24946 (N_24946,N_20532,N_21707);
or U24947 (N_24947,N_21481,N_21491);
or U24948 (N_24948,N_19948,N_19037);
xor U24949 (N_24949,N_19022,N_18911);
xnor U24950 (N_24950,N_21458,N_21577);
xor U24951 (N_24951,N_21309,N_18761);
nand U24952 (N_24952,N_20767,N_18900);
and U24953 (N_24953,N_19154,N_18899);
nor U24954 (N_24954,N_20210,N_18911);
and U24955 (N_24955,N_19134,N_20002);
xor U24956 (N_24956,N_21163,N_21185);
and U24957 (N_24957,N_19176,N_18963);
nand U24958 (N_24958,N_19660,N_19358);
xor U24959 (N_24959,N_18966,N_18942);
nor U24960 (N_24960,N_20760,N_20357);
xnor U24961 (N_24961,N_20752,N_19266);
nand U24962 (N_24962,N_20872,N_20800);
and U24963 (N_24963,N_21170,N_19431);
nor U24964 (N_24964,N_20199,N_20647);
and U24965 (N_24965,N_20040,N_21414);
xnor U24966 (N_24966,N_21410,N_20634);
nor U24967 (N_24967,N_20199,N_19410);
xnor U24968 (N_24968,N_21076,N_21772);
and U24969 (N_24969,N_20644,N_21134);
nand U24970 (N_24970,N_19318,N_20242);
or U24971 (N_24971,N_21707,N_21590);
xor U24972 (N_24972,N_21380,N_18937);
and U24973 (N_24973,N_19185,N_21517);
or U24974 (N_24974,N_19142,N_20524);
nor U24975 (N_24975,N_20504,N_20292);
nand U24976 (N_24976,N_20742,N_20285);
nand U24977 (N_24977,N_20239,N_21746);
or U24978 (N_24978,N_19430,N_21206);
or U24979 (N_24979,N_19947,N_20207);
xor U24980 (N_24980,N_21392,N_20255);
nand U24981 (N_24981,N_20134,N_20109);
xnor U24982 (N_24982,N_19193,N_19924);
nand U24983 (N_24983,N_20453,N_18800);
nor U24984 (N_24984,N_21474,N_19840);
nand U24985 (N_24985,N_21299,N_19042);
nor U24986 (N_24986,N_20019,N_21679);
xor U24987 (N_24987,N_20389,N_18788);
nand U24988 (N_24988,N_20046,N_21041);
nand U24989 (N_24989,N_21398,N_21401);
nor U24990 (N_24990,N_20810,N_19687);
nor U24991 (N_24991,N_18871,N_21254);
or U24992 (N_24992,N_19922,N_20456);
or U24993 (N_24993,N_19499,N_21689);
and U24994 (N_24994,N_18999,N_21754);
or U24995 (N_24995,N_19402,N_20195);
or U24996 (N_24996,N_19575,N_20229);
or U24997 (N_24997,N_20263,N_20382);
and U24998 (N_24998,N_21430,N_19803);
or U24999 (N_24999,N_19376,N_19050);
nand UO_0 (O_0,N_22932,N_22892);
nor UO_1 (O_1,N_22549,N_22482);
or UO_2 (O_2,N_24956,N_23365);
xnor UO_3 (O_3,N_23484,N_24700);
and UO_4 (O_4,N_22885,N_21899);
or UO_5 (O_5,N_24094,N_24801);
or UO_6 (O_6,N_24422,N_24464);
and UO_7 (O_7,N_23627,N_24066);
and UO_8 (O_8,N_24593,N_23065);
nor UO_9 (O_9,N_23548,N_22598);
xor UO_10 (O_10,N_24634,N_24431);
nor UO_11 (O_11,N_23987,N_24779);
nand UO_12 (O_12,N_22069,N_24039);
xor UO_13 (O_13,N_22292,N_21905);
nand UO_14 (O_14,N_23039,N_23165);
nand UO_15 (O_15,N_22622,N_23741);
xor UO_16 (O_16,N_24460,N_24982);
xnor UO_17 (O_17,N_23344,N_24459);
nand UO_18 (O_18,N_24358,N_22277);
or UO_19 (O_19,N_23535,N_24374);
nand UO_20 (O_20,N_24591,N_22075);
nor UO_21 (O_21,N_24028,N_22456);
nand UO_22 (O_22,N_24698,N_22116);
and UO_23 (O_23,N_22923,N_22788);
xor UO_24 (O_24,N_22125,N_24230);
or UO_25 (O_25,N_21991,N_24708);
xnor UO_26 (O_26,N_22301,N_24138);
nor UO_27 (O_27,N_24117,N_23498);
and UO_28 (O_28,N_24636,N_24868);
or UO_29 (O_29,N_23454,N_24471);
or UO_30 (O_30,N_22603,N_22385);
or UO_31 (O_31,N_24174,N_23709);
or UO_32 (O_32,N_24862,N_24935);
xnor UO_33 (O_33,N_24263,N_23087);
or UO_34 (O_34,N_22959,N_24482);
nand UO_35 (O_35,N_22178,N_22046);
nor UO_36 (O_36,N_24725,N_22585);
nor UO_37 (O_37,N_23685,N_23421);
nor UO_38 (O_38,N_23300,N_23049);
nand UO_39 (O_39,N_23791,N_24297);
nor UO_40 (O_40,N_23128,N_21901);
or UO_41 (O_41,N_24666,N_24999);
xnor UO_42 (O_42,N_24254,N_21975);
or UO_43 (O_43,N_22085,N_22538);
nor UO_44 (O_44,N_23567,N_22865);
nand UO_45 (O_45,N_24293,N_23771);
nand UO_46 (O_46,N_22105,N_22400);
and UO_47 (O_47,N_24723,N_24490);
or UO_48 (O_48,N_24947,N_23358);
xnor UO_49 (O_49,N_23982,N_24484);
and UO_50 (O_50,N_24560,N_24571);
and UO_51 (O_51,N_22479,N_24467);
nand UO_52 (O_52,N_23700,N_24913);
nand UO_53 (O_53,N_24200,N_24001);
xor UO_54 (O_54,N_21990,N_24056);
or UO_55 (O_55,N_24266,N_22605);
nor UO_56 (O_56,N_22147,N_22316);
xor UO_57 (O_57,N_23657,N_24368);
xnor UO_58 (O_58,N_23983,N_22853);
and UO_59 (O_59,N_24645,N_23582);
xnor UO_60 (O_60,N_23889,N_23642);
or UO_61 (O_61,N_23540,N_22615);
nand UO_62 (O_62,N_22650,N_21880);
nand UO_63 (O_63,N_22851,N_23763);
xnor UO_64 (O_64,N_23171,N_22429);
nor UO_65 (O_65,N_24992,N_22079);
nand UO_66 (O_66,N_22729,N_22383);
xnor UO_67 (O_67,N_24295,N_24895);
or UO_68 (O_68,N_24470,N_24410);
or UO_69 (O_69,N_23179,N_24069);
or UO_70 (O_70,N_24510,N_21922);
and UO_71 (O_71,N_22869,N_23356);
nor UO_72 (O_72,N_22396,N_24438);
and UO_73 (O_73,N_24364,N_23021);
nand UO_74 (O_74,N_24535,N_23005);
nor UO_75 (O_75,N_23729,N_23139);
nor UO_76 (O_76,N_23821,N_22483);
and UO_77 (O_77,N_24648,N_24633);
and UO_78 (O_78,N_23203,N_23321);
nand UO_79 (O_79,N_24531,N_22874);
or UO_80 (O_80,N_22269,N_22347);
nand UO_81 (O_81,N_24301,N_23743);
and UO_82 (O_82,N_22665,N_22058);
xor UO_83 (O_83,N_24639,N_22290);
xnor UO_84 (O_84,N_23731,N_23011);
and UO_85 (O_85,N_24567,N_24215);
or UO_86 (O_86,N_23302,N_24188);
nand UO_87 (O_87,N_21893,N_22230);
or UO_88 (O_88,N_22312,N_22578);
and UO_89 (O_89,N_24447,N_24048);
or UO_90 (O_90,N_23490,N_24541);
xor UO_91 (O_91,N_23591,N_24413);
nor UO_92 (O_92,N_24125,N_23470);
nand UO_93 (O_93,N_24092,N_23032);
xnor UO_94 (O_94,N_24345,N_23249);
nor UO_95 (O_95,N_23904,N_23148);
or UO_96 (O_96,N_22397,N_24803);
xor UO_97 (O_97,N_24772,N_22379);
nand UO_98 (O_98,N_22274,N_24565);
nor UO_99 (O_99,N_22144,N_21981);
or UO_100 (O_100,N_22083,N_24338);
nand UO_101 (O_101,N_23383,N_24225);
nor UO_102 (O_102,N_23501,N_24930);
nor UO_103 (O_103,N_24155,N_22670);
nor UO_104 (O_104,N_24549,N_23696);
and UO_105 (O_105,N_22203,N_22737);
and UO_106 (O_106,N_23975,N_24176);
and UO_107 (O_107,N_23584,N_22451);
nor UO_108 (O_108,N_23668,N_24060);
or UO_109 (O_109,N_21908,N_22242);
nand UO_110 (O_110,N_23955,N_22883);
nand UO_111 (O_111,N_22082,N_24475);
or UO_112 (O_112,N_22110,N_22593);
or UO_113 (O_113,N_22698,N_23341);
and UO_114 (O_114,N_22754,N_24850);
or UO_115 (O_115,N_22661,N_24332);
xnor UO_116 (O_116,N_23984,N_22284);
nor UO_117 (O_117,N_24024,N_23655);
and UO_118 (O_118,N_22489,N_24390);
xor UO_119 (O_119,N_22070,N_21997);
nor UO_120 (O_120,N_24748,N_23089);
nor UO_121 (O_121,N_22461,N_22188);
nor UO_122 (O_122,N_24169,N_22699);
xor UO_123 (O_123,N_22162,N_23328);
and UO_124 (O_124,N_22283,N_24903);
nor UO_125 (O_125,N_24749,N_23835);
and UO_126 (O_126,N_23558,N_23331);
nand UO_127 (O_127,N_23831,N_22955);
xnor UO_128 (O_128,N_23518,N_24908);
xnor UO_129 (O_129,N_24319,N_21993);
and UO_130 (O_130,N_22835,N_24971);
or UO_131 (O_131,N_22246,N_24557);
xor UO_132 (O_132,N_22989,N_22264);
and UO_133 (O_133,N_24082,N_22010);
nor UO_134 (O_134,N_24519,N_23440);
nand UO_135 (O_135,N_24622,N_22167);
nor UO_136 (O_136,N_22543,N_22308);
nor UO_137 (O_137,N_24409,N_24106);
nor UO_138 (O_138,N_24950,N_23527);
nor UO_139 (O_139,N_24329,N_22368);
nand UO_140 (O_140,N_24785,N_23986);
xnor UO_141 (O_141,N_24341,N_24035);
and UO_142 (O_142,N_22163,N_23172);
nand UO_143 (O_143,N_24281,N_24185);
and UO_144 (O_144,N_24796,N_23464);
xnor UO_145 (O_145,N_24685,N_23661);
and UO_146 (O_146,N_23739,N_22993);
or UO_147 (O_147,N_23303,N_24370);
nand UO_148 (O_148,N_24916,N_23911);
xor UO_149 (O_149,N_23543,N_22651);
nor UO_150 (O_150,N_21967,N_22027);
xnor UO_151 (O_151,N_23592,N_23812);
xnor UO_152 (O_152,N_23929,N_22848);
or UO_153 (O_153,N_23631,N_23375);
nand UO_154 (O_154,N_24737,N_24610);
nor UO_155 (O_155,N_24638,N_22200);
nand UO_156 (O_156,N_22618,N_24898);
xnor UO_157 (O_157,N_24624,N_23413);
or UO_158 (O_158,N_24896,N_24975);
nand UO_159 (O_159,N_22221,N_21930);
nand UO_160 (O_160,N_22755,N_23467);
nor UO_161 (O_161,N_23168,N_22182);
or UO_162 (O_162,N_24960,N_24403);
nand UO_163 (O_163,N_22502,N_24811);
nand UO_164 (O_164,N_24775,N_23836);
xor UO_165 (O_165,N_22903,N_23541);
nand UO_166 (O_166,N_22638,N_23735);
nand UO_167 (O_167,N_23227,N_23636);
nand UO_168 (O_168,N_24515,N_23216);
nor UO_169 (O_169,N_22157,N_21881);
or UO_170 (O_170,N_24984,N_22793);
xor UO_171 (O_171,N_22506,N_22223);
or UO_172 (O_172,N_23914,N_22683);
xnor UO_173 (O_173,N_22297,N_24857);
nand UO_174 (O_174,N_22669,N_22621);
or UO_175 (O_175,N_22662,N_22189);
or UO_176 (O_176,N_24837,N_24500);
xnor UO_177 (O_177,N_24030,N_22612);
or UO_178 (O_178,N_24335,N_21875);
nor UO_179 (O_179,N_24049,N_23422);
nand UO_180 (O_180,N_22779,N_21999);
xnor UO_181 (O_181,N_22627,N_23083);
nand UO_182 (O_182,N_23802,N_21951);
nand UO_183 (O_183,N_23629,N_22518);
xnor UO_184 (O_184,N_23967,N_24559);
xor UO_185 (O_185,N_23207,N_23517);
xor UO_186 (O_186,N_24613,N_22298);
nand UO_187 (O_187,N_23095,N_24325);
nor UO_188 (O_188,N_23145,N_23441);
nor UO_189 (O_189,N_24417,N_21982);
and UO_190 (O_190,N_23732,N_23676);
nand UO_191 (O_191,N_22108,N_24197);
nand UO_192 (O_192,N_23869,N_24781);
and UO_193 (O_193,N_23251,N_24569);
nand UO_194 (O_194,N_23519,N_22407);
nor UO_195 (O_195,N_22623,N_22315);
nor UO_196 (O_196,N_23725,N_22090);
xnor UO_197 (O_197,N_24420,N_21896);
nand UO_198 (O_198,N_22440,N_23728);
nor UO_199 (O_199,N_24934,N_24282);
and UO_200 (O_200,N_23730,N_21961);
nor UO_201 (O_201,N_24443,N_24695);
nand UO_202 (O_202,N_22752,N_23574);
nor UO_203 (O_203,N_24177,N_23839);
nand UO_204 (O_204,N_24555,N_23220);
and UO_205 (O_205,N_24219,N_22911);
nand UO_206 (O_206,N_24929,N_23794);
nand UO_207 (O_207,N_22417,N_22735);
xor UO_208 (O_208,N_22318,N_24681);
nor UO_209 (O_209,N_22330,N_23536);
or UO_210 (O_210,N_22153,N_24642);
or UO_211 (O_211,N_24096,N_23160);
or UO_212 (O_212,N_22926,N_24608);
or UO_213 (O_213,N_22691,N_24159);
nand UO_214 (O_214,N_21962,N_23840);
and UO_215 (O_215,N_22837,N_24717);
and UO_216 (O_216,N_22654,N_24970);
xor UO_217 (O_217,N_23183,N_23691);
xnor UO_218 (O_218,N_23516,N_24157);
nor UO_219 (O_219,N_24814,N_24211);
xnor UO_220 (O_220,N_23443,N_21944);
nand UO_221 (O_221,N_23803,N_22380);
and UO_222 (O_222,N_24561,N_22204);
or UO_223 (O_223,N_23617,N_22427);
xor UO_224 (O_224,N_21892,N_22310);
xor UO_225 (O_225,N_22378,N_22453);
and UO_226 (O_226,N_24827,N_23876);
nand UO_227 (O_227,N_24037,N_22697);
xor UO_228 (O_228,N_22876,N_24804);
nor UO_229 (O_229,N_22834,N_24978);
xnor UO_230 (O_230,N_24365,N_22859);
or UO_231 (O_231,N_23182,N_23782);
and UO_232 (O_232,N_24290,N_24339);
nand UO_233 (O_233,N_22843,N_23446);
xor UO_234 (O_234,N_24799,N_21978);
nand UO_235 (O_235,N_22106,N_21952);
nor UO_236 (O_236,N_22820,N_24308);
xnor UO_237 (O_237,N_24248,N_22325);
and UO_238 (O_238,N_21945,N_22646);
nand UO_239 (O_239,N_23043,N_23656);
nand UO_240 (O_240,N_23336,N_24356);
nand UO_241 (O_241,N_22761,N_22015);
or UO_242 (O_242,N_22857,N_24946);
or UO_243 (O_243,N_22282,N_24378);
xnor UO_244 (O_244,N_23618,N_22233);
or UO_245 (O_245,N_24952,N_24141);
and UO_246 (O_246,N_22476,N_22012);
xnor UO_247 (O_247,N_22252,N_22652);
or UO_248 (O_248,N_23176,N_24881);
xnor UO_249 (O_249,N_22139,N_22565);
nor UO_250 (O_250,N_24637,N_22135);
nor UO_251 (O_251,N_23395,N_24711);
xnor UO_252 (O_252,N_23632,N_22057);
xnor UO_253 (O_253,N_23202,N_24939);
or UO_254 (O_254,N_21938,N_23265);
nand UO_255 (O_255,N_22171,N_22887);
nor UO_256 (O_256,N_24554,N_23092);
xnor UO_257 (O_257,N_24179,N_23100);
nor UO_258 (O_258,N_22966,N_22248);
nand UO_259 (O_259,N_24265,N_23744);
xnor UO_260 (O_260,N_24053,N_23916);
xor UO_261 (O_261,N_23275,N_24388);
xor UO_262 (O_262,N_24525,N_22634);
nand UO_263 (O_263,N_24387,N_24943);
nand UO_264 (O_264,N_23684,N_23430);
and UO_265 (O_265,N_23279,N_24103);
or UO_266 (O_266,N_23166,N_23210);
nor UO_267 (O_267,N_22151,N_23890);
or UO_268 (O_268,N_23236,N_21947);
xor UO_269 (O_269,N_21927,N_23273);
xor UO_270 (O_270,N_23532,N_22713);
and UO_271 (O_271,N_21992,N_23660);
or UO_272 (O_272,N_21941,N_23297);
xor UO_273 (O_273,N_24016,N_24757);
or UO_274 (O_274,N_22224,N_22327);
nand UO_275 (O_275,N_22013,N_23118);
xor UO_276 (O_276,N_22401,N_24307);
xnor UO_277 (O_277,N_23854,N_23779);
and UO_278 (O_278,N_24000,N_21932);
or UO_279 (O_279,N_22706,N_24474);
nor UO_280 (O_280,N_22728,N_24210);
xor UO_281 (O_281,N_23801,N_23019);
or UO_282 (O_282,N_23526,N_22405);
and UO_283 (O_283,N_24823,N_22500);
or UO_284 (O_284,N_23809,N_24260);
or UO_285 (O_285,N_23943,N_23439);
xnor UO_286 (O_286,N_23956,N_23020);
or UO_287 (O_287,N_22542,N_23740);
nor UO_288 (O_288,N_23958,N_23834);
and UO_289 (O_289,N_22433,N_24243);
nand UO_290 (O_290,N_22709,N_23832);
or UO_291 (O_291,N_23828,N_22474);
and UO_292 (O_292,N_24574,N_24678);
nand UO_293 (O_293,N_24062,N_22954);
nor UO_294 (O_294,N_22152,N_24366);
or UO_295 (O_295,N_22969,N_21907);
nand UO_296 (O_296,N_24452,N_22562);
and UO_297 (O_297,N_24523,N_24668);
nor UO_298 (O_298,N_22340,N_24171);
xor UO_299 (O_299,N_22191,N_23286);
xnor UO_300 (O_300,N_22700,N_23376);
nand UO_301 (O_301,N_22055,N_23368);
nand UO_302 (O_302,N_23351,N_21943);
xor UO_303 (O_303,N_24380,N_22617);
or UO_304 (O_304,N_24831,N_22839);
nand UO_305 (O_305,N_24318,N_22444);
and UO_306 (O_306,N_23350,N_22939);
or UO_307 (O_307,N_23615,N_24488);
nor UO_308 (O_308,N_24227,N_24437);
or UO_309 (O_309,N_24126,N_22904);
or UO_310 (O_310,N_22810,N_24166);
xor UO_311 (O_311,N_22580,N_23616);
and UO_312 (O_312,N_22552,N_23865);
nor UO_313 (O_313,N_24257,N_22856);
nand UO_314 (O_314,N_22637,N_23170);
nor UO_315 (O_315,N_22514,N_24679);
and UO_316 (O_316,N_24396,N_23481);
or UO_317 (O_317,N_23968,N_24373);
xnor UO_318 (O_318,N_24832,N_23770);
xor UO_319 (O_319,N_24118,N_24235);
nor UO_320 (O_320,N_23082,N_23733);
or UO_321 (O_321,N_22493,N_22148);
nand UO_322 (O_322,N_23322,N_23537);
xor UO_323 (O_323,N_24888,N_22100);
or UO_324 (O_324,N_21903,N_22997);
nor UO_325 (O_325,N_24596,N_22778);
xor UO_326 (O_326,N_24316,N_22335);
nor UO_327 (O_327,N_22767,N_22443);
nor UO_328 (O_328,N_24451,N_22421);
nor UO_329 (O_329,N_24556,N_24239);
or UO_330 (O_330,N_24033,N_23442);
nand UO_331 (O_331,N_23923,N_23436);
and UO_332 (O_332,N_22909,N_23724);
nor UO_333 (O_333,N_21895,N_24922);
and UO_334 (O_334,N_23169,N_24280);
xor UO_335 (O_335,N_23387,N_24528);
nand UO_336 (O_336,N_22832,N_22109);
nand UO_337 (O_337,N_23643,N_24603);
and UO_338 (O_338,N_23564,N_23306);
nor UO_339 (O_339,N_24466,N_22648);
nor UO_340 (O_340,N_23283,N_22631);
and UO_341 (O_341,N_22068,N_23244);
and UO_342 (O_342,N_23380,N_23962);
xor UO_343 (O_343,N_24289,N_21897);
and UO_344 (O_344,N_23121,N_24505);
nand UO_345 (O_345,N_23680,N_23980);
nand UO_346 (O_346,N_23882,N_23897);
or UO_347 (O_347,N_22094,N_22672);
and UO_348 (O_348,N_24404,N_23280);
nand UO_349 (O_349,N_24847,N_22146);
and UO_350 (O_350,N_24963,N_22115);
nor UO_351 (O_351,N_24167,N_22293);
and UO_352 (O_352,N_22497,N_23091);
nor UO_353 (O_353,N_23901,N_22168);
or UO_354 (O_354,N_22470,N_24566);
or UO_355 (O_355,N_22642,N_24444);
and UO_356 (O_356,N_21894,N_24958);
nand UO_357 (O_357,N_22219,N_22731);
nor UO_358 (O_358,N_23263,N_24981);
or UO_359 (O_359,N_23742,N_22093);
nand UO_360 (O_360,N_23458,N_24376);
or UO_361 (O_361,N_24303,N_22468);
nand UO_362 (O_362,N_24479,N_22430);
xor UO_363 (O_363,N_24629,N_23424);
xnor UO_364 (O_364,N_24813,N_24778);
and UO_365 (O_365,N_23381,N_23237);
nor UO_366 (O_366,N_24285,N_23648);
nor UO_367 (O_367,N_22925,N_22428);
xnor UO_368 (O_368,N_24109,N_23152);
or UO_369 (O_369,N_24544,N_24650);
and UO_370 (O_370,N_23282,N_24462);
nand UO_371 (O_371,N_23206,N_24936);
or UO_372 (O_372,N_23683,N_22101);
and UO_373 (O_373,N_23056,N_24029);
nand UO_374 (O_374,N_23063,N_23900);
nor UO_375 (O_375,N_22686,N_23106);
nand UO_376 (O_376,N_24229,N_22555);
nand UO_377 (O_377,N_24580,N_23124);
nand UO_378 (O_378,N_24392,N_23465);
nand UO_379 (O_379,N_22088,N_24760);
nand UO_380 (O_380,N_23159,N_22893);
and UO_381 (O_381,N_23068,N_24761);
nor UO_382 (O_382,N_23193,N_23504);
nand UO_383 (O_383,N_23506,N_22673);
nand UO_384 (O_384,N_21876,N_21911);
nand UO_385 (O_385,N_23402,N_23959);
xnor UO_386 (O_386,N_22991,N_23090);
nor UO_387 (O_387,N_24866,N_24925);
or UO_388 (O_388,N_23186,N_24383);
and UO_389 (O_389,N_23213,N_23130);
nor UO_390 (O_390,N_22038,N_23158);
nand UO_391 (O_391,N_23222,N_24040);
nand UO_392 (O_392,N_23167,N_22568);
or UO_393 (O_393,N_24083,N_23602);
nor UO_394 (O_394,N_23879,N_23639);
nor UO_395 (O_395,N_24721,N_22557);
nand UO_396 (O_396,N_24587,N_22990);
xor UO_397 (O_397,N_23462,N_23468);
nor UO_398 (O_398,N_22948,N_22712);
xnor UO_399 (O_399,N_22968,N_24601);
nor UO_400 (O_400,N_23954,N_22973);
or UO_401 (O_401,N_23188,N_22566);
and UO_402 (O_402,N_22358,N_22207);
nand UO_403 (O_403,N_24730,N_22376);
and UO_404 (O_404,N_24232,N_22987);
nand UO_405 (O_405,N_24027,N_24321);
nand UO_406 (O_406,N_22575,N_22439);
or UO_407 (O_407,N_23241,N_22112);
xor UO_408 (O_408,N_22394,N_22352);
nand UO_409 (O_409,N_23852,N_23099);
and UO_410 (O_410,N_22745,N_24792);
or UO_411 (O_411,N_23486,N_23933);
nor UO_412 (O_412,N_24630,N_23940);
xor UO_413 (O_413,N_23154,N_22520);
xor UO_414 (O_414,N_23664,N_22722);
and UO_415 (O_415,N_24269,N_24607);
and UO_416 (O_416,N_22127,N_23748);
nor UO_417 (O_417,N_23931,N_23960);
nor UO_418 (O_418,N_22913,N_21965);
and UO_419 (O_419,N_23530,N_23494);
or UO_420 (O_420,N_24480,N_22229);
or UO_421 (O_421,N_22256,N_22052);
nor UO_422 (O_422,N_23925,N_22632);
nand UO_423 (O_423,N_23784,N_23194);
or UO_424 (O_424,N_22854,N_22464);
nand UO_425 (O_425,N_22759,N_23059);
or UO_426 (O_426,N_22087,N_24191);
xnor UO_427 (O_427,N_21998,N_24842);
and UO_428 (O_428,N_24296,N_22604);
and UO_429 (O_429,N_23457,N_24416);
nand UO_430 (O_430,N_22322,N_24445);
or UO_431 (O_431,N_22721,N_24546);
or UO_432 (O_432,N_22080,N_24495);
xnor UO_433 (O_433,N_22936,N_23822);
or UO_434 (O_434,N_23508,N_23399);
nand UO_435 (O_435,N_24399,N_23572);
nor UO_436 (O_436,N_24920,N_22158);
nand UO_437 (O_437,N_23335,N_24507);
or UO_438 (O_438,N_22225,N_23776);
and UO_439 (O_439,N_23229,N_23147);
and UO_440 (O_440,N_23247,N_22216);
or UO_441 (O_441,N_23654,N_23524);
or UO_442 (O_442,N_24520,N_22956);
xor UO_443 (O_443,N_22689,N_23102);
or UO_444 (O_444,N_22360,N_23198);
or UO_445 (O_445,N_23476,N_24770);
nor UO_446 (O_446,N_23703,N_23444);
nand UO_447 (O_447,N_24806,N_24110);
or UO_448 (O_448,N_22704,N_24870);
nor UO_449 (O_449,N_23001,N_23348);
nor UO_450 (O_450,N_23971,N_23094);
or UO_451 (O_451,N_23093,N_24855);
and UO_452 (O_452,N_22197,N_23769);
xor UO_453 (O_453,N_24738,N_22947);
nor UO_454 (O_454,N_22845,N_24463);
xnor UO_455 (O_455,N_22600,N_24043);
and UO_456 (O_456,N_24545,N_24133);
xnor UO_457 (O_457,N_23233,N_22595);
nand UO_458 (O_458,N_22798,N_22446);
and UO_459 (O_459,N_24222,N_22475);
xor UO_460 (O_460,N_23425,N_24627);
nor UO_461 (O_461,N_23266,N_21954);
and UO_462 (O_462,N_22594,N_22355);
and UO_463 (O_463,N_23401,N_22445);
or UO_464 (O_464,N_22361,N_21900);
and UO_465 (O_465,N_22384,N_22748);
nand UO_466 (O_466,N_22041,N_23204);
nor UO_467 (O_467,N_23354,N_24497);
nand UO_468 (O_468,N_24506,N_23562);
or UO_469 (O_469,N_23717,N_22777);
or UO_470 (O_470,N_21889,N_22763);
or UO_471 (O_471,N_23410,N_21995);
nand UO_472 (O_472,N_22460,N_23754);
nor UO_473 (O_473,N_24893,N_24237);
xor UO_474 (O_474,N_22424,N_23581);
or UO_475 (O_475,N_22756,N_23420);
nand UO_476 (O_476,N_22681,N_23529);
or UO_477 (O_477,N_24489,N_22694);
xnor UO_478 (O_478,N_22334,N_21935);
and UO_479 (O_479,N_21996,N_22916);
nand UO_480 (O_480,N_22227,N_23891);
or UO_481 (O_481,N_22020,N_24384);
or UO_482 (O_482,N_23333,N_24744);
xor UO_483 (O_483,N_24747,N_22527);
or UO_484 (O_484,N_22138,N_24931);
nor UO_485 (O_485,N_23972,N_22123);
nor UO_486 (O_486,N_22348,N_22420);
nand UO_487 (O_487,N_22550,N_23327);
nand UO_488 (O_488,N_23910,N_23042);
xor UO_489 (O_489,N_24894,N_24707);
xor UO_490 (O_490,N_23793,N_23755);
or UO_491 (O_491,N_24588,N_24874);
or UO_492 (O_492,N_23449,N_24287);
nand UO_493 (O_493,N_24100,N_22061);
and UO_494 (O_494,N_24713,N_23583);
or UO_495 (O_495,N_22862,N_24647);
or UO_496 (O_496,N_23539,N_22448);
nor UO_497 (O_497,N_22553,N_24820);
nor UO_498 (O_498,N_24203,N_23597);
xnor UO_499 (O_499,N_24848,N_24741);
nor UO_500 (O_500,N_24421,N_24104);
or UO_501 (O_501,N_23843,N_23577);
xor UO_502 (O_502,N_23080,N_23277);
nor UO_503 (O_503,N_24492,N_24932);
nand UO_504 (O_504,N_22036,N_24328);
or UO_505 (O_505,N_21949,N_24268);
nor UO_506 (O_506,N_24472,N_23845);
nor UO_507 (O_507,N_23447,N_22332);
nand UO_508 (O_508,N_24754,N_23290);
and UO_509 (O_509,N_21878,N_24824);
or UO_510 (O_510,N_22881,N_23573);
nor UO_511 (O_511,N_22114,N_22343);
nor UO_512 (O_512,N_22695,N_22986);
or UO_513 (O_513,N_23463,N_22899);
nand UO_514 (O_514,N_22096,N_23699);
and UO_515 (O_515,N_24865,N_24822);
nor UO_516 (O_516,N_23177,N_24284);
nand UO_517 (O_517,N_22739,N_23261);
nor UO_518 (O_518,N_22273,N_23364);
or UO_519 (O_519,N_22608,N_24455);
or UO_520 (O_520,N_24899,N_23565);
xor UO_521 (O_521,N_23818,N_23837);
and UO_522 (O_522,N_24724,N_23930);
nor UO_523 (O_523,N_22510,N_22812);
or UO_524 (O_524,N_24693,N_22048);
nor UO_525 (O_525,N_22970,N_23781);
and UO_526 (O_526,N_24797,N_24209);
and UO_527 (O_527,N_24871,N_22150);
xor UO_528 (O_528,N_24651,N_22403);
nand UO_529 (O_529,N_24733,N_23509);
or UO_530 (O_530,N_23600,N_24694);
or UO_531 (O_531,N_22303,N_23939);
xor UO_532 (O_532,N_23480,N_23448);
nand UO_533 (O_533,N_23450,N_23132);
and UO_534 (O_534,N_23620,N_22888);
nor UO_535 (O_535,N_22091,N_23292);
nand UO_536 (O_536,N_22732,N_24632);
nor UO_537 (O_537,N_23775,N_23459);
nand UO_538 (O_538,N_24954,N_24270);
nor UO_539 (O_539,N_24620,N_24068);
and UO_540 (O_540,N_22607,N_21888);
nand UO_541 (O_541,N_24305,N_24578);
nor UO_542 (O_542,N_23310,N_23515);
or UO_543 (O_543,N_23619,N_21933);
nor UO_544 (O_544,N_22131,N_21939);
or UO_545 (O_545,N_22588,N_23815);
or UO_546 (O_546,N_21980,N_24706);
nor UO_547 (O_547,N_22996,N_24299);
or UO_548 (O_548,N_22641,N_24671);
or UO_549 (O_549,N_22441,N_22934);
nor UO_550 (O_550,N_24148,N_24010);
and UO_551 (O_551,N_24701,N_23569);
nor UO_552 (O_552,N_24113,N_24055);
and UO_553 (O_553,N_24461,N_23624);
or UO_554 (O_554,N_23675,N_23579);
or UO_555 (O_555,N_24716,N_24509);
nor UO_556 (O_556,N_22677,N_22611);
nor UO_557 (O_557,N_21877,N_22043);
and UO_558 (O_558,N_23318,N_22583);
nor UO_559 (O_559,N_23920,N_22202);
nor UO_560 (O_560,N_22363,N_23008);
xor UO_561 (O_561,N_24306,N_24019);
nand UO_562 (O_562,N_24604,N_22306);
xnor UO_563 (O_563,N_23197,N_22323);
xor UO_564 (O_564,N_24252,N_24663);
nand UO_565 (O_565,N_23884,N_23824);
and UO_566 (O_566,N_22126,N_22772);
and UO_567 (O_567,N_22077,N_24496);
and UO_568 (O_568,N_24655,N_22165);
xor UO_569 (O_569,N_22907,N_22491);
nand UO_570 (O_570,N_23223,N_23074);
or UO_571 (O_571,N_23587,N_23066);
or UO_572 (O_572,N_23038,N_24729);
and UO_573 (O_573,N_24542,N_23892);
xor UO_574 (O_574,N_23362,N_24928);
xor UO_575 (O_575,N_22032,N_22978);
or UO_576 (O_576,N_24526,N_23786);
xor UO_577 (O_577,N_23034,N_24802);
xor UO_578 (O_578,N_22828,N_22567);
xnor UO_579 (O_579,N_23998,N_23231);
nor UO_580 (O_580,N_22140,N_21918);
or UO_581 (O_581,N_24057,N_24786);
or UO_582 (O_582,N_24712,N_23386);
and UO_583 (O_583,N_24530,N_22179);
and UO_584 (O_584,N_24324,N_24734);
xnor UO_585 (O_585,N_23308,N_22056);
xor UO_586 (O_586,N_21984,N_22251);
or UO_587 (O_587,N_24833,N_23808);
nor UO_588 (O_588,N_23963,N_22922);
nor UO_589 (O_589,N_24377,N_23403);
and UO_590 (O_590,N_22792,N_23307);
nand UO_591 (O_591,N_23885,N_24382);
or UO_592 (O_592,N_22485,N_23418);
and UO_593 (O_593,N_23859,N_24527);
or UO_594 (O_594,N_23894,N_23941);
or UO_595 (O_595,N_23334,N_24063);
nor UO_596 (O_596,N_23667,N_24830);
nand UO_597 (O_597,N_22022,N_22940);
and UO_598 (O_598,N_23215,N_24736);
or UO_599 (O_599,N_24501,N_23557);
xor UO_600 (O_600,N_23004,N_22558);
or UO_601 (O_601,N_23614,N_23738);
xor UO_602 (O_602,N_21925,N_22784);
and UO_603 (O_603,N_21885,N_22659);
xnor UO_604 (O_604,N_24614,N_24783);
nor UO_605 (O_605,N_21985,N_24087);
xnor UO_606 (O_606,N_24398,N_24327);
nor UO_607 (O_607,N_22213,N_23598);
xnor UO_608 (O_608,N_23133,N_22432);
and UO_609 (O_609,N_24766,N_22742);
nor UO_610 (O_610,N_24623,N_22133);
and UO_611 (O_611,N_22003,N_24592);
or UO_612 (O_612,N_23257,N_23497);
and UO_613 (O_613,N_24071,N_24320);
and UO_614 (O_614,N_24143,N_22898);
or UO_615 (O_615,N_23295,N_24142);
and UO_616 (O_616,N_24054,N_24626);
nand UO_617 (O_617,N_22173,N_22279);
or UO_618 (O_618,N_23713,N_24579);
xnor UO_619 (O_619,N_23605,N_23291);
nor UO_620 (O_620,N_21983,N_23604);
nor UO_621 (O_621,N_24375,N_22818);
nand UO_622 (O_622,N_23585,N_22176);
nor UO_623 (O_623,N_22212,N_22750);
nor UO_624 (O_624,N_23363,N_24955);
nand UO_625 (O_625,N_22826,N_23305);
and UO_626 (O_626,N_24397,N_24017);
and UO_627 (O_627,N_23922,N_22042);
or UO_628 (O_628,N_23281,N_22597);
and UO_629 (O_629,N_24890,N_23847);
nand UO_630 (O_630,N_23329,N_21914);
nand UO_631 (O_631,N_24199,N_23814);
nor UO_632 (O_632,N_22582,N_21942);
xnor UO_633 (O_633,N_24718,N_24805);
nor UO_634 (O_634,N_24393,N_23666);
and UO_635 (O_635,N_24773,N_22534);
nand UO_636 (O_636,N_23314,N_22829);
or UO_637 (O_637,N_24121,N_22855);
xnor UO_638 (O_638,N_23199,N_22289);
and UO_639 (O_639,N_24491,N_22124);
nor UO_640 (O_640,N_24826,N_22645);
nand UO_641 (O_641,N_22504,N_22917);
or UO_642 (O_642,N_22620,N_22438);
xor UO_643 (O_643,N_23571,N_24139);
nor UO_644 (O_644,N_24080,N_22921);
xnor UO_645 (O_645,N_21879,N_22769);
or UO_646 (O_646,N_23949,N_22258);
or UO_647 (O_647,N_22018,N_24816);
nor UO_648 (O_648,N_24617,N_22785);
xnor UO_649 (O_649,N_22389,N_22074);
nand UO_650 (O_650,N_23390,N_24228);
nor UO_651 (O_651,N_23027,N_23479);
and UO_652 (O_652,N_22508,N_24849);
nor UO_653 (O_653,N_24149,N_22831);
or UO_654 (O_654,N_22338,N_24156);
xor UO_655 (O_655,N_24953,N_24808);
nand UO_656 (O_656,N_24605,N_24189);
nand UO_657 (O_657,N_23745,N_23347);
or UO_658 (O_658,N_22195,N_24988);
nor UO_659 (O_659,N_22198,N_24787);
xor UO_660 (O_660,N_24611,N_24344);
and UO_661 (O_661,N_24957,N_23451);
nor UO_662 (O_662,N_23379,N_24547);
or UO_663 (O_663,N_24310,N_24722);
xnor UO_664 (O_664,N_24261,N_23064);
xor UO_665 (O_665,N_23270,N_22095);
or UO_666 (O_666,N_23819,N_24059);
nand UO_667 (O_667,N_22353,N_22145);
xor UO_668 (O_668,N_22764,N_24234);
xor UO_669 (O_669,N_21973,N_23811);
and UO_670 (O_670,N_24046,N_21921);
and UO_671 (O_671,N_23687,N_24715);
nor UO_672 (O_672,N_23412,N_22507);
nor UO_673 (O_673,N_24845,N_23478);
and UO_674 (O_674,N_22309,N_24765);
and UO_675 (O_675,N_23560,N_23895);
nand UO_676 (O_676,N_22743,N_23205);
or UO_677 (O_677,N_22367,N_23150);
and UO_678 (O_678,N_22858,N_24690);
or UO_679 (O_679,N_22344,N_24841);
nand UO_680 (O_680,N_23325,N_23003);
or UO_681 (O_681,N_23966,N_22897);
xnor UO_682 (O_682,N_23077,N_23874);
xor UO_683 (O_683,N_22039,N_23239);
or UO_684 (O_684,N_21920,N_24764);
and UO_685 (O_685,N_24991,N_23499);
nor UO_686 (O_686,N_23384,N_22571);
nand UO_687 (O_687,N_23969,N_22243);
nor UO_688 (O_688,N_22701,N_24277);
nand UO_689 (O_689,N_24271,N_22800);
xor UO_690 (O_690,N_23455,N_22406);
and UO_691 (O_691,N_23903,N_22076);
nand UO_692 (O_692,N_23252,N_24919);
nand UO_693 (O_693,N_24672,N_21956);
nand UO_694 (O_694,N_22636,N_23477);
or UO_695 (O_695,N_23672,N_22035);
nor UO_696 (O_696,N_23164,N_24331);
nand UO_697 (O_697,N_22537,N_22257);
xnor UO_698 (O_698,N_22501,N_22512);
nor UO_699 (O_699,N_24658,N_24440);
xnor UO_700 (O_700,N_24099,N_23758);
xnor UO_701 (O_701,N_22245,N_24732);
xnor UO_702 (O_702,N_24311,N_22418);
and UO_703 (O_703,N_22574,N_24442);
nor UO_704 (O_704,N_23682,N_24021);
xor UO_705 (O_705,N_24120,N_23103);
or UO_706 (O_706,N_23848,N_22516);
nor UO_707 (O_707,N_22640,N_21955);
or UO_708 (O_708,N_23271,N_24381);
and UO_709 (O_709,N_23419,N_24134);
nand UO_710 (O_710,N_24883,N_23311);
and UO_711 (O_711,N_22238,N_23235);
nor UO_712 (O_712,N_23951,N_23370);
nor UO_713 (O_713,N_22214,N_22628);
and UO_714 (O_714,N_22121,N_22169);
or UO_715 (O_715,N_24145,N_24192);
and UO_716 (O_716,N_22692,N_24818);
or UO_717 (O_717,N_23195,N_24949);
nand UO_718 (O_718,N_24294,N_24322);
or UO_719 (O_719,N_22668,N_24670);
or UO_720 (O_720,N_22410,N_23670);
nor UO_721 (O_721,N_23645,N_22643);
and UO_722 (O_722,N_22024,N_23071);
nand UO_723 (O_723,N_22590,N_22045);
and UO_724 (O_724,N_24077,N_23330);
or UO_725 (O_725,N_22547,N_24573);
and UO_726 (O_726,N_22736,N_22840);
xor UO_727 (O_727,N_21994,N_22649);
nor UO_728 (O_728,N_23997,N_24217);
xnor UO_729 (O_729,N_23023,N_24244);
or UO_730 (O_730,N_23714,N_23640);
and UO_731 (O_731,N_24807,N_24882);
nor UO_732 (O_732,N_24979,N_23533);
nor UO_733 (O_733,N_23267,N_24423);
xor UO_734 (O_734,N_23495,N_24635);
and UO_735 (O_735,N_24485,N_23817);
or UO_736 (O_736,N_24709,N_22375);
xor UO_737 (O_737,N_22920,N_22525);
and UO_738 (O_738,N_22321,N_22192);
nand UO_739 (O_739,N_23936,N_22159);
nor UO_740 (O_740,N_22240,N_24927);
and UO_741 (O_741,N_24326,N_24869);
nand UO_742 (O_742,N_23414,N_23146);
nor UO_743 (O_743,N_24575,N_23841);
xor UO_744 (O_744,N_24313,N_22016);
nor UO_745 (O_745,N_23012,N_24386);
or UO_746 (O_746,N_22795,N_24540);
nor UO_747 (O_747,N_24061,N_21916);
and UO_748 (O_748,N_23471,N_24272);
xor UO_749 (O_749,N_24763,N_22259);
nand UO_750 (O_750,N_21923,N_24524);
nor UO_751 (O_751,N_23323,N_22073);
xnor UO_752 (O_752,N_23340,N_23992);
nor UO_753 (O_753,N_23461,N_22369);
nand UO_754 (O_754,N_24187,N_23887);
xnor UO_755 (O_755,N_23805,N_23912);
nand UO_756 (O_756,N_22805,N_24619);
xnor UO_757 (O_757,N_22236,N_23635);
xnor UO_758 (O_758,N_23137,N_23423);
nand UO_759 (O_759,N_22398,N_22962);
xor UO_760 (O_760,N_23453,N_23899);
nand UO_761 (O_761,N_23542,N_22462);
or UO_762 (O_762,N_23861,N_23787);
nor UO_763 (O_763,N_24669,N_24255);
nor UO_764 (O_764,N_23795,N_24330);
or UO_765 (O_765,N_23711,N_24691);
nand UO_766 (O_766,N_23599,N_24508);
nand UO_767 (O_767,N_23698,N_22031);
nor UO_768 (O_768,N_24965,N_22878);
and UO_769 (O_769,N_23907,N_22773);
or UO_770 (O_770,N_22072,N_22569);
or UO_771 (O_771,N_24817,N_22879);
or UO_772 (O_772,N_23438,N_22675);
and UO_773 (O_773,N_22164,N_23877);
or UO_774 (O_774,N_23970,N_23678);
nand UO_775 (O_775,N_22724,N_23262);
or UO_776 (O_776,N_24846,N_21958);
xnor UO_777 (O_777,N_22584,N_23829);
nor UO_778 (O_778,N_23719,N_22783);
nor UO_779 (O_779,N_23031,N_23086);
or UO_780 (O_780,N_24130,N_23369);
and UO_781 (O_781,N_22050,N_23760);
or UO_782 (O_782,N_22941,N_21909);
nand UO_783 (O_783,N_24070,N_24279);
or UO_784 (O_784,N_24684,N_23114);
and UO_785 (O_785,N_24606,N_22809);
nand UO_786 (O_786,N_23488,N_23646);
or UO_787 (O_787,N_24628,N_23669);
and UO_788 (O_788,N_24940,N_23878);
xor UO_789 (O_789,N_23482,N_22875);
xnor UO_790 (O_790,N_22572,N_22299);
nor UO_791 (O_791,N_22753,N_22924);
xnor UO_792 (O_792,N_24728,N_22599);
xnor UO_793 (O_793,N_22237,N_23312);
and UO_794 (O_794,N_22836,N_22806);
nand UO_795 (O_795,N_23218,N_24562);
nor UO_796 (O_796,N_22864,N_23069);
nand UO_797 (O_797,N_22725,N_22281);
or UO_798 (O_798,N_22149,N_23595);
xnor UO_799 (O_799,N_22247,N_23294);
and UO_800 (O_800,N_24058,N_23394);
and UO_801 (O_801,N_23208,N_24091);
xnor UO_802 (O_802,N_23790,N_24727);
or UO_803 (O_803,N_24116,N_22868);
or UO_804 (O_804,N_22919,N_22452);
and UO_805 (O_805,N_22331,N_23830);
and UO_806 (O_806,N_23919,N_24045);
nor UO_807 (O_807,N_23674,N_22827);
or UO_808 (O_808,N_22768,N_22313);
nor UO_809 (O_809,N_24221,N_24878);
nor UO_810 (O_810,N_24346,N_24714);
xor UO_811 (O_811,N_23634,N_22546);
and UO_812 (O_812,N_23060,N_22730);
nor UO_813 (O_813,N_24664,N_22944);
or UO_814 (O_814,N_24915,N_24184);
xor UO_815 (O_815,N_23751,N_22180);
nand UO_816 (O_816,N_22426,N_23772);
nand UO_817 (O_817,N_24917,N_23695);
nand UO_818 (O_818,N_24275,N_23580);
xor UO_819 (O_819,N_23965,N_22847);
or UO_820 (O_820,N_22625,N_23374);
nand UO_821 (O_821,N_22296,N_23298);
xor UO_822 (O_822,N_23337,N_24660);
nor UO_823 (O_823,N_24078,N_24692);
nand UO_824 (O_824,N_23606,N_23378);
or UO_825 (O_825,N_23913,N_23456);
xnor UO_826 (O_826,N_22791,N_22602);
nor UO_827 (O_827,N_23136,N_23588);
nor UO_828 (O_828,N_24864,N_22177);
xor UO_829 (O_829,N_22496,N_24625);
and UO_830 (O_830,N_23993,N_24705);
nand UO_831 (O_831,N_22766,N_24406);
and UO_832 (O_832,N_22317,N_23129);
nand UO_833 (O_833,N_23245,N_22120);
or UO_834 (O_834,N_21887,N_24202);
nand UO_835 (O_835,N_23545,N_22624);
or UO_836 (O_836,N_23985,N_24434);
xnor UO_837 (O_837,N_22591,N_22596);
nor UO_838 (O_838,N_24697,N_22842);
nor UO_839 (O_839,N_23994,N_22263);
nand UO_840 (O_840,N_22435,N_24923);
xnor UO_841 (O_841,N_22678,N_24673);
nor UO_842 (O_842,N_22589,N_24590);
nand UO_843 (O_843,N_23734,N_23762);
and UO_844 (O_844,N_24997,N_23946);
xor UO_845 (O_845,N_22183,N_22170);
and UO_846 (O_846,N_22351,N_23045);
or UO_847 (O_847,N_22824,N_22660);
nor UO_848 (O_848,N_23144,N_23044);
nor UO_849 (O_849,N_23917,N_22218);
or UO_850 (O_850,N_24755,N_24767);
or UO_851 (O_851,N_23964,N_23209);
nor UO_852 (O_852,N_23029,N_24859);
nor UO_853 (O_853,N_21946,N_24007);
nand UO_854 (O_854,N_22789,N_22155);
xnor UO_855 (O_855,N_22821,N_23076);
and UO_856 (O_856,N_22688,N_22184);
nor UO_857 (O_857,N_23342,N_22690);
nor UO_858 (O_858,N_22528,N_23594);
and UO_859 (O_859,N_22117,N_23823);
xor UO_860 (O_860,N_22872,N_22026);
xnor UO_861 (O_861,N_22674,N_24987);
and UO_862 (O_862,N_23293,N_23881);
nand UO_863 (O_863,N_24369,N_23033);
xnor UO_864 (O_864,N_22387,N_23816);
xnor UO_865 (O_865,N_24880,N_23737);
and UO_866 (O_866,N_24676,N_24385);
and UO_867 (O_867,N_24933,N_23007);
and UO_868 (O_868,N_22253,N_22981);
nor UO_869 (O_869,N_22174,N_22365);
nand UO_870 (O_870,N_21979,N_22577);
nand UO_871 (O_871,N_21886,N_22972);
xor UO_872 (O_872,N_24493,N_23372);
xnor UO_873 (O_873,N_24851,N_24577);
xor UO_874 (O_874,N_22244,N_23367);
xor UO_875 (O_875,N_22463,N_22413);
xor UO_876 (O_876,N_24348,N_22029);
or UO_877 (O_877,N_23633,N_22328);
or UO_878 (O_878,N_22033,N_23221);
and UO_879 (O_879,N_24689,N_23827);
and UO_880 (O_880,N_23407,N_23162);
nand UO_881 (O_881,N_23934,N_22733);
and UO_882 (O_882,N_24581,N_22097);
nor UO_883 (O_883,N_24128,N_24115);
or UO_884 (O_884,N_21950,N_22586);
xnor UO_885 (O_885,N_23650,N_24433);
or UO_886 (O_886,N_24517,N_23035);
or UO_887 (O_887,N_23570,N_22040);
nand UO_888 (O_888,N_24391,N_23534);
or UO_889 (O_889,N_22492,N_21974);
nor UO_890 (O_890,N_22945,N_23768);
nand UO_891 (O_891,N_23452,N_24250);
or UO_892 (O_892,N_22007,N_24583);
nand UO_893 (O_893,N_23320,N_24008);
nor UO_894 (O_894,N_24503,N_24173);
nand UO_895 (O_895,N_22776,N_22006);
or UO_896 (O_896,N_24810,N_24834);
or UO_897 (O_897,N_22710,N_23016);
and UO_898 (O_898,N_23609,N_22610);
or UO_899 (O_899,N_24262,N_24704);
nor UO_900 (O_900,N_24951,N_23345);
nand UO_901 (O_901,N_22034,N_23433);
nand UO_902 (O_902,N_22098,N_22132);
or UO_903 (O_903,N_24563,N_24178);
nor UO_904 (O_904,N_22350,N_22908);
or UO_905 (O_905,N_23142,N_21924);
nor UO_906 (O_906,N_24214,N_24012);
or UO_907 (O_907,N_23196,N_24002);
and UO_908 (O_908,N_24990,N_22342);
xnor UO_909 (O_909,N_23697,N_24966);
nor UO_910 (O_910,N_22209,N_23692);
nor UO_911 (O_911,N_22630,N_22799);
nor UO_912 (O_912,N_23797,N_23608);
xnor UO_913 (O_913,N_23511,N_23988);
nor UO_914 (O_914,N_22494,N_23041);
nor UO_915 (O_915,N_22044,N_23224);
or UO_916 (O_916,N_24815,N_22532);
xor UO_917 (O_917,N_24050,N_23686);
xnor UO_918 (O_918,N_24891,N_24224);
and UO_919 (O_919,N_24347,N_23906);
nand UO_920 (O_920,N_24825,N_22053);
nor UO_921 (O_921,N_24323,N_24948);
nand UO_922 (O_922,N_23996,N_24205);
and UO_923 (O_923,N_24075,N_24513);
and UO_924 (O_924,N_23647,N_22942);
nand UO_925 (O_925,N_24640,N_22544);
nor UO_926 (O_926,N_23405,N_24137);
nor UO_927 (O_927,N_23067,N_23621);
and UO_928 (O_928,N_22220,N_24361);
and UO_929 (O_929,N_24877,N_22285);
xnor UO_930 (O_930,N_22128,N_22633);
nand UO_931 (O_931,N_21917,N_24876);
xnor UO_932 (O_932,N_22503,N_22684);
nand UO_933 (O_933,N_22187,N_23551);
nor UO_934 (O_934,N_22559,N_24745);
and UO_935 (O_935,N_24353,N_22314);
nor UO_936 (O_936,N_23690,N_23799);
or UO_937 (O_937,N_24032,N_23234);
nand UO_938 (O_938,N_22844,N_24844);
and UO_939 (O_939,N_23935,N_24789);
nand UO_940 (O_940,N_22134,N_24750);
nor UO_941 (O_941,N_24389,N_23974);
nand UO_942 (O_942,N_22472,N_22521);
or UO_943 (O_943,N_22037,N_24759);
nand UO_944 (O_944,N_23947,N_22957);
and UO_945 (O_945,N_24430,N_22129);
xnor UO_946 (O_946,N_23382,N_23550);
xor UO_947 (O_947,N_22931,N_24912);
or UO_948 (O_948,N_22122,N_22781);
nor UO_949 (O_949,N_24206,N_24314);
or UO_950 (O_950,N_23396,N_22235);
nor UO_951 (O_951,N_23316,N_22971);
or UO_952 (O_952,N_21977,N_22272);
nor UO_953 (O_953,N_23278,N_23662);
or UO_954 (O_954,N_24616,N_23902);
xnor UO_955 (O_955,N_24131,N_22531);
nor UO_956 (O_956,N_22092,N_24426);
nand UO_957 (O_957,N_23360,N_23641);
xnor UO_958 (O_958,N_24753,N_24534);
or UO_959 (O_959,N_23025,N_22196);
nand UO_960 (O_960,N_23757,N_23568);
nor UO_961 (O_961,N_23849,N_22536);
xnor UO_962 (O_962,N_24022,N_24967);
or UO_963 (O_963,N_24703,N_23437);
or UO_964 (O_964,N_23723,N_23120);
and UO_965 (O_965,N_23649,N_23792);
and UO_966 (O_966,N_22601,N_23028);
xnor UO_967 (O_967,N_22288,N_24873);
and UO_968 (O_968,N_22530,N_22081);
or UO_969 (O_969,N_24959,N_24516);
nand UO_970 (O_970,N_22391,N_24972);
nand UO_971 (O_971,N_24656,N_23110);
or UO_972 (O_972,N_24351,N_24400);
nand UO_973 (O_973,N_24158,N_24476);
and UO_974 (O_974,N_24446,N_23301);
xor UO_975 (O_975,N_24095,N_24473);
or UO_976 (O_976,N_23746,N_22786);
and UO_977 (O_977,N_23937,N_24904);
nand UO_978 (O_978,N_22466,N_23324);
or UO_979 (O_979,N_22228,N_24667);
or UO_980 (O_980,N_24253,N_22241);
nor UO_981 (O_981,N_23932,N_24182);
nor UO_982 (O_982,N_23549,N_22930);
xnor UO_983 (O_983,N_22873,N_22490);
nor UO_984 (O_984,N_23050,N_22703);
and UO_985 (O_985,N_23109,N_22587);
xor UO_986 (O_986,N_23628,N_24558);
or UO_987 (O_987,N_22811,N_24146);
xor UO_988 (O_988,N_22980,N_23346);
xor UO_989 (O_989,N_22425,N_21884);
or UO_990 (O_990,N_23926,N_24198);
or UO_991 (O_991,N_22307,N_24769);
or UO_992 (O_992,N_22671,N_22199);
nor UO_993 (O_993,N_24233,N_23860);
and UO_994 (O_994,N_23397,N_24315);
or UO_995 (O_995,N_24828,N_22780);
xnor UO_996 (O_996,N_22563,N_23623);
or UO_997 (O_997,N_24276,N_23510);
nand UO_998 (O_998,N_22261,N_24696);
and UO_999 (O_999,N_23752,N_22062);
or UO_1000 (O_1000,N_22967,N_23864);
and UO_1001 (O_1001,N_23976,N_23434);
nor UO_1002 (O_1002,N_23555,N_24892);
xnor UO_1003 (O_1003,N_23915,N_22647);
and UO_1004 (O_1004,N_22816,N_24494);
nand UO_1005 (O_1005,N_22556,N_23727);
nor UO_1006 (O_1006,N_23174,N_22723);
nand UO_1007 (O_1007,N_22653,N_24312);
or UO_1008 (O_1008,N_23072,N_24107);
and UO_1009 (O_1009,N_22336,N_24273);
xnor UO_1010 (O_1010,N_22071,N_23192);
nand UO_1011 (O_1011,N_23006,N_23406);
and UO_1012 (O_1012,N_22513,N_22477);
nor UO_1013 (O_1013,N_22963,N_21989);
and UO_1014 (O_1014,N_24976,N_22382);
or UO_1015 (O_1015,N_22030,N_22841);
nor UO_1016 (O_1016,N_23153,N_24469);
and UO_1017 (O_1017,N_22679,N_23804);
xor UO_1018 (O_1018,N_24020,N_22442);
xor UO_1019 (O_1019,N_23546,N_24968);
xor UO_1020 (O_1020,N_22409,N_22107);
xnor UO_1021 (O_1021,N_24751,N_24532);
or UO_1022 (O_1022,N_24570,N_22629);
nand UO_1023 (O_1023,N_22877,N_23472);
xor UO_1024 (O_1024,N_23313,N_23688);
nor UO_1025 (O_1025,N_24595,N_23055);
xor UO_1026 (O_1026,N_23105,N_22481);
or UO_1027 (O_1027,N_24111,N_23671);
nor UO_1028 (O_1028,N_23088,N_22938);
nand UO_1029 (O_1029,N_22867,N_24242);
or UO_1030 (O_1030,N_24044,N_22850);
nand UO_1031 (O_1031,N_24538,N_24465);
nand UO_1032 (O_1032,N_22863,N_24969);
nor UO_1033 (O_1033,N_24897,N_22912);
nand UO_1034 (O_1034,N_22005,N_23825);
or UO_1035 (O_1035,N_22457,N_22366);
or UO_1036 (O_1036,N_23689,N_24247);
and UO_1037 (O_1037,N_24419,N_21891);
nand UO_1038 (O_1038,N_23255,N_23953);
and UO_1039 (O_1039,N_23774,N_24129);
nor UO_1040 (O_1040,N_23134,N_22469);
nor UO_1041 (O_1041,N_23058,N_23866);
nor UO_1042 (O_1042,N_24291,N_24119);
and UO_1043 (O_1043,N_23979,N_24112);
xnor UO_1044 (O_1044,N_22415,N_24288);
and UO_1045 (O_1045,N_22801,N_23973);
nand UO_1046 (O_1046,N_22300,N_23749);
and UO_1047 (O_1047,N_23037,N_24791);
xor UO_1048 (O_1048,N_24181,N_24914);
nand UO_1049 (O_1049,N_23015,N_24144);
and UO_1050 (O_1050,N_23214,N_22802);
nor UO_1051 (O_1051,N_24011,N_21976);
nand UO_1052 (O_1052,N_22813,N_22541);
xor UO_1053 (O_1053,N_23556,N_22374);
nor UO_1054 (O_1054,N_22254,N_22419);
xor UO_1055 (O_1055,N_22262,N_24836);
and UO_1056 (O_1056,N_21883,N_22664);
or UO_1057 (O_1057,N_23264,N_23590);
xnor UO_1058 (O_1058,N_23211,N_23905);
nor UO_1059 (O_1059,N_24401,N_22803);
nand UO_1060 (O_1060,N_22614,N_22656);
xnor UO_1061 (O_1061,N_22302,N_22141);
and UO_1062 (O_1062,N_24025,N_22175);
or UO_1063 (O_1063,N_22084,N_22143);
nor UO_1064 (O_1064,N_23528,N_24101);
xor UO_1065 (O_1065,N_21926,N_22935);
nor UO_1066 (O_1066,N_22866,N_24425);
nor UO_1067 (O_1067,N_24165,N_23726);
nor UO_1068 (O_1068,N_22119,N_24408);
nor UO_1069 (O_1069,N_22716,N_22267);
or UO_1070 (O_1070,N_24889,N_23415);
or UO_1071 (O_1071,N_23736,N_24884);
and UO_1072 (O_1072,N_23856,N_23844);
xor UO_1073 (O_1073,N_22918,N_22746);
or UO_1074 (O_1074,N_23990,N_23013);
and UO_1075 (O_1075,N_23187,N_24342);
nand UO_1076 (O_1076,N_24572,N_22232);
or UO_1077 (O_1077,N_24264,N_23126);
and UO_1078 (O_1078,N_22422,N_22319);
nor UO_1079 (O_1079,N_21936,N_22393);
xnor UO_1080 (O_1080,N_22609,N_22390);
and UO_1081 (O_1081,N_24031,N_24909);
nand UO_1082 (O_1082,N_23761,N_22270);
and UO_1083 (O_1083,N_23141,N_23212);
xor UO_1084 (O_1084,N_22009,N_23131);
nor UO_1085 (O_1085,N_24352,N_22161);
or UO_1086 (O_1086,N_22255,N_24609);
or UO_1087 (O_1087,N_22995,N_22359);
nand UO_1088 (O_1088,N_23693,N_22581);
nand UO_1089 (O_1089,N_22201,N_23589);
and UO_1090 (O_1090,N_22749,N_22311);
or UO_1091 (O_1091,N_24201,N_24355);
and UO_1092 (O_1092,N_22994,N_23638);
nor UO_1093 (O_1093,N_23612,N_22860);
nand UO_1094 (O_1094,N_24394,N_22324);
xor UO_1095 (O_1095,N_23896,N_23432);
and UO_1096 (O_1096,N_22346,N_24521);
xor UO_1097 (O_1097,N_24140,N_23151);
nand UO_1098 (O_1098,N_22111,N_23416);
nand UO_1099 (O_1099,N_22822,N_22751);
or UO_1100 (O_1100,N_23140,N_23022);
or UO_1101 (O_1101,N_23081,N_24858);
nand UO_1102 (O_1102,N_23681,N_24589);
nand UO_1103 (O_1103,N_24241,N_24097);
nor UO_1104 (O_1104,N_22222,N_23858);
and UO_1105 (O_1105,N_24402,N_24405);
nand UO_1106 (O_1106,N_22362,N_22915);
xnor UO_1107 (O_1107,N_22304,N_24108);
or UO_1108 (O_1108,N_24776,N_23226);
nor UO_1109 (O_1109,N_24756,N_22089);
or UO_1110 (O_1110,N_22714,N_23503);
nor UO_1111 (O_1111,N_23652,N_23554);
nor UO_1112 (O_1112,N_21972,N_22974);
nand UO_1113 (O_1113,N_23123,N_23052);
nand UO_1114 (O_1114,N_23596,N_23232);
or UO_1115 (O_1115,N_24190,N_24081);
nor UO_1116 (O_1116,N_22771,N_23181);
or UO_1117 (O_1117,N_23813,N_22329);
and UO_1118 (O_1118,N_24812,N_22548);
xnor UO_1119 (O_1119,N_22437,N_23888);
and UO_1120 (O_1120,N_22280,N_23009);
nor UO_1121 (O_1121,N_24362,N_22370);
nand UO_1122 (O_1122,N_22431,N_24584);
nor UO_1123 (O_1123,N_22998,N_24731);
nor UO_1124 (O_1124,N_23122,N_24942);
or UO_1125 (O_1125,N_24548,N_23927);
xnor UO_1126 (O_1126,N_24962,N_23626);
nor UO_1127 (O_1127,N_22804,N_24151);
xnor UO_1128 (O_1128,N_24172,N_22626);
and UO_1129 (O_1129,N_23276,N_22765);
nand UO_1130 (O_1130,N_22774,N_22983);
or UO_1131 (O_1131,N_23576,N_24514);
nand UO_1132 (O_1132,N_22579,N_23961);
or UO_1133 (O_1133,N_22949,N_24800);
xnor UO_1134 (O_1134,N_22054,N_21959);
xor UO_1135 (O_1135,N_23873,N_22488);
nand UO_1136 (O_1136,N_22592,N_24994);
nand UO_1137 (O_1137,N_22411,N_24887);
nand UO_1138 (O_1138,N_24599,N_24675);
and UO_1139 (O_1139,N_24843,N_23637);
nor UO_1140 (O_1140,N_24902,N_23785);
or UO_1141 (O_1141,N_24003,N_22193);
xor UO_1142 (O_1142,N_23796,N_22696);
nand UO_1143 (O_1143,N_24586,N_24457);
or UO_1144 (O_1144,N_24918,N_22961);
nand UO_1145 (O_1145,N_22889,N_24441);
or UO_1146 (O_1146,N_24788,N_22208);
nand UO_1147 (O_1147,N_23073,N_23780);
xnor UO_1148 (O_1148,N_22682,N_24996);
nand UO_1149 (O_1149,N_23010,N_24743);
nand UO_1150 (O_1150,N_22511,N_23217);
nand UO_1151 (O_1151,N_24079,N_23789);
or UO_1152 (O_1152,N_24085,N_22937);
and UO_1153 (O_1153,N_22345,N_24259);
nand UO_1154 (O_1154,N_23863,N_22519);
nor UO_1155 (O_1155,N_22928,N_22357);
nand UO_1156 (O_1156,N_24758,N_23319);
xor UO_1157 (O_1157,N_24477,N_23720);
nor UO_1158 (O_1158,N_22113,N_24795);
or UO_1159 (O_1159,N_24298,N_23062);
nand UO_1160 (O_1160,N_22099,N_23750);
or UO_1161 (O_1161,N_23538,N_21929);
and UO_1162 (O_1162,N_22814,N_22408);
xnor UO_1163 (O_1163,N_23883,N_22616);
or UO_1164 (O_1164,N_22976,N_22613);
nor UO_1165 (O_1165,N_23898,N_22059);
and UO_1166 (O_1166,N_23259,N_23002);
or UO_1167 (O_1167,N_22927,N_22535);
nand UO_1168 (O_1168,N_23101,N_24995);
xnor UO_1169 (O_1169,N_22894,N_23445);
nand UO_1170 (O_1170,N_22902,N_23428);
or UO_1171 (O_1171,N_23474,N_24659);
xor UO_1172 (O_1172,N_24518,N_24090);
nand UO_1173 (O_1173,N_24852,N_22953);
nand UO_1174 (O_1174,N_24486,N_24161);
nand UO_1175 (O_1175,N_23357,N_22830);
xnor UO_1176 (O_1176,N_24653,N_22726);
nor UO_1177 (O_1177,N_22066,N_22870);
nand UO_1178 (O_1178,N_23523,N_23173);
nand UO_1179 (O_1179,N_23607,N_22658);
and UO_1180 (O_1180,N_23500,N_23553);
nand UO_1181 (O_1181,N_22717,N_22635);
xor UO_1182 (O_1182,N_24193,N_22666);
or UO_1183 (O_1183,N_24359,N_24009);
or UO_1184 (O_1184,N_22136,N_23677);
nand UO_1185 (O_1185,N_23185,N_22137);
or UO_1186 (O_1186,N_22564,N_24600);
nand UO_1187 (O_1187,N_23127,N_24015);
xnor UO_1188 (O_1188,N_22522,N_24317);
nand UO_1189 (O_1189,N_23520,N_21971);
or UO_1190 (O_1190,N_23559,N_21966);
and UO_1191 (O_1191,N_23928,N_23868);
or UO_1192 (O_1192,N_22551,N_22423);
xor UO_1193 (O_1193,N_24334,N_24553);
xnor UO_1194 (O_1194,N_24218,N_23078);
nor UO_1195 (O_1195,N_24710,N_22740);
or UO_1196 (O_1196,N_23502,N_24006);
or UO_1197 (O_1197,N_24537,N_22693);
nand UO_1198 (O_1198,N_24938,N_23810);
or UO_1199 (O_1199,N_23918,N_23981);
or UO_1200 (O_1200,N_22891,N_22294);
or UO_1201 (O_1201,N_23189,N_22060);
or UO_1202 (O_1202,N_22741,N_23332);
nand UO_1203 (O_1203,N_23644,N_24989);
xor UO_1204 (O_1204,N_24005,N_22979);
xor UO_1205 (O_1205,N_22454,N_23250);
xnor UO_1206 (O_1206,N_24371,N_23460);
and UO_1207 (O_1207,N_23807,N_24762);
nor UO_1208 (O_1208,N_24771,N_24336);
and UO_1209 (O_1209,N_24478,N_22655);
xor UO_1210 (O_1210,N_22975,N_22487);
and UO_1211 (O_1211,N_22561,N_23366);
nor UO_1212 (O_1212,N_24631,N_24941);
xor UO_1213 (O_1213,N_24512,N_24292);
or UO_1214 (O_1214,N_22402,N_24867);
nor UO_1215 (O_1215,N_22166,N_23846);
and UO_1216 (O_1216,N_24739,N_24089);
nor UO_1217 (O_1217,N_23427,N_23288);
nand UO_1218 (O_1218,N_21960,N_22349);
xnor UO_1219 (O_1219,N_24152,N_22364);
xor UO_1220 (O_1220,N_22950,N_23544);
xor UO_1221 (O_1221,N_22011,N_24212);
nor UO_1222 (O_1222,N_22757,N_23798);
and UO_1223 (O_1223,N_24164,N_23201);
xnor UO_1224 (O_1224,N_24226,N_23701);
nand UO_1225 (O_1225,N_24418,N_22985);
nand UO_1226 (O_1226,N_24088,N_23184);
and UO_1227 (O_1227,N_22190,N_24945);
xnor UO_1228 (O_1228,N_23191,N_23716);
or UO_1229 (O_1229,N_24983,N_22064);
nor UO_1230 (O_1230,N_24041,N_24170);
xnor UO_1231 (O_1231,N_24379,N_23575);
nand UO_1232 (O_1232,N_22484,N_22871);
nor UO_1233 (O_1233,N_23175,N_22825);
xor UO_1234 (O_1234,N_24350,N_24042);
nor UO_1235 (O_1235,N_23258,N_23806);
or UO_1236 (O_1236,N_24674,N_23908);
nor UO_1237 (O_1237,N_24036,N_24964);
nand UO_1238 (O_1238,N_23287,N_23219);
nor UO_1239 (O_1239,N_23361,N_24699);
nand UO_1240 (O_1240,N_23240,N_23857);
nor UO_1241 (O_1241,N_22952,N_24782);
nand UO_1242 (O_1242,N_24429,N_23853);
nand UO_1243 (O_1243,N_22320,N_22639);
and UO_1244 (O_1244,N_22333,N_23256);
xnor UO_1245 (O_1245,N_23285,N_24594);
xnor UO_1246 (O_1246,N_22782,N_23135);
and UO_1247 (O_1247,N_24564,N_23269);
nor UO_1248 (O_1248,N_22880,N_24539);
or UO_1249 (O_1249,N_24498,N_22205);
xnor UO_1250 (O_1250,N_22882,N_22102);
or UO_1251 (O_1251,N_23057,N_24886);
nand UO_1252 (O_1252,N_24682,N_23492);
and UO_1253 (O_1253,N_24456,N_24768);
or UO_1254 (O_1254,N_22014,N_24481);
nor UO_1255 (O_1255,N_21969,N_24123);
or UO_1256 (O_1256,N_24977,N_23978);
nor UO_1257 (O_1257,N_22392,N_23409);
nor UO_1258 (O_1258,N_23163,N_24504);
nor UO_1259 (O_1259,N_23948,N_24340);
nand UO_1260 (O_1260,N_22371,N_23851);
nand UO_1261 (O_1261,N_23253,N_23143);
nor UO_1262 (O_1262,N_23704,N_23521);
and UO_1263 (O_1263,N_23673,N_24618);
or UO_1264 (O_1264,N_22051,N_24124);
and UO_1265 (O_1265,N_23070,N_24924);
nor UO_1266 (O_1266,N_22958,N_23909);
and UO_1267 (O_1267,N_23024,N_24986);
nand UO_1268 (O_1268,N_22929,N_22895);
or UO_1269 (O_1269,N_22539,N_23466);
nor UO_1270 (O_1270,N_24283,N_22797);
and UO_1271 (O_1271,N_22760,N_23315);
or UO_1272 (O_1272,N_24661,N_23872);
xnor UO_1273 (O_1273,N_22480,N_22770);
or UO_1274 (O_1274,N_24026,N_22554);
xnor UO_1275 (O_1275,N_24160,N_23352);
nor UO_1276 (O_1276,N_23400,N_22265);
xor UO_1277 (O_1277,N_22271,N_22744);
nor UO_1278 (O_1278,N_22708,N_22458);
xnor UO_1279 (O_1279,N_22478,N_22373);
nand UO_1280 (O_1280,N_22896,N_22808);
nor UO_1281 (O_1281,N_22906,N_22796);
xor UO_1282 (O_1282,N_24944,N_22545);
nand UO_1283 (O_1283,N_22217,N_22275);
or UO_1284 (O_1284,N_24856,N_21988);
xor UO_1285 (O_1285,N_24240,N_22738);
xor UO_1286 (O_1286,N_21913,N_24993);
nand UO_1287 (O_1287,N_23242,N_22404);
nand UO_1288 (O_1288,N_23097,N_24652);
nor UO_1289 (O_1289,N_23601,N_24487);
nor UO_1290 (O_1290,N_24168,N_24216);
nand UO_1291 (O_1291,N_24127,N_23886);
nand UO_1292 (O_1292,N_22447,N_24220);
xnor UO_1293 (O_1293,N_21963,N_24499);
or UO_1294 (O_1294,N_23408,N_22194);
xnor UO_1295 (O_1295,N_24612,N_23777);
nand UO_1296 (O_1296,N_23766,N_22023);
and UO_1297 (O_1297,N_23149,N_22910);
xnor UO_1298 (O_1298,N_22386,N_23921);
xnor UO_1299 (O_1299,N_23469,N_22946);
nor UO_1300 (O_1300,N_22529,N_21953);
or UO_1301 (O_1301,N_23339,N_24395);
xnor UO_1302 (O_1302,N_24790,N_23417);
or UO_1303 (O_1303,N_22762,N_23343);
or UO_1304 (O_1304,N_24543,N_22000);
xor UO_1305 (O_1305,N_24576,N_24654);
nand UO_1306 (O_1306,N_22372,N_24135);
or UO_1307 (O_1307,N_24853,N_24207);
xnor UO_1308 (O_1308,N_23663,N_24136);
and UO_1309 (O_1309,N_23513,N_24901);
and UO_1310 (O_1310,N_24363,N_23079);
nand UO_1311 (O_1311,N_22295,N_23708);
nand UO_1312 (O_1312,N_23820,N_24657);
or UO_1313 (O_1313,N_23659,N_22416);
or UO_1314 (O_1314,N_22606,N_24582);
and UO_1315 (O_1315,N_22523,N_24921);
xnor UO_1316 (O_1316,N_24256,N_24649);
or UO_1317 (O_1317,N_24067,N_24449);
and UO_1318 (O_1318,N_24450,N_22434);
and UO_1319 (O_1319,N_24662,N_24536);
and UO_1320 (O_1320,N_22185,N_23991);
and UO_1321 (O_1321,N_22450,N_22861);
xnor UO_1322 (O_1322,N_22819,N_24163);
nand UO_1323 (O_1323,N_23871,N_23359);
nand UO_1324 (O_1324,N_22815,N_22250);
or UO_1325 (O_1325,N_24439,N_24780);
or UO_1326 (O_1326,N_24646,N_24047);
and UO_1327 (O_1327,N_23429,N_24854);
and UO_1328 (O_1328,N_23112,N_22160);
nor UO_1329 (O_1329,N_23800,N_24819);
nand UO_1330 (O_1330,N_24267,N_24407);
or UO_1331 (O_1331,N_23783,N_22573);
xor UO_1332 (O_1332,N_23952,N_22852);
xnor UO_1333 (O_1333,N_23238,N_23505);
nor UO_1334 (O_1334,N_24213,N_24236);
nor UO_1335 (O_1335,N_24074,N_23392);
xor UO_1336 (O_1336,N_22680,N_24551);
nand UO_1337 (O_1337,N_24175,N_21964);
and UO_1338 (O_1338,N_22715,N_24302);
nor UO_1339 (O_1339,N_24084,N_23487);
xnor UO_1340 (O_1340,N_23706,N_23272);
and UO_1341 (O_1341,N_23243,N_24102);
or UO_1342 (O_1342,N_24098,N_22377);
or UO_1343 (O_1343,N_23349,N_24726);
nor UO_1344 (O_1344,N_23371,N_21902);
or UO_1345 (O_1345,N_21928,N_24702);
xnor UO_1346 (O_1346,N_23155,N_24742);
and UO_1347 (O_1347,N_22291,N_23875);
xor UO_1348 (O_1348,N_24186,N_22002);
or UO_1349 (O_1349,N_22211,N_24643);
nand UO_1350 (O_1350,N_22960,N_23630);
xor UO_1351 (O_1351,N_22172,N_23000);
or UO_1352 (O_1352,N_24838,N_23040);
and UO_1353 (O_1353,N_22215,N_22455);
nand UO_1354 (O_1354,N_24286,N_23679);
xor UO_1355 (O_1355,N_21882,N_22459);
or UO_1356 (O_1356,N_24483,N_24415);
xor UO_1357 (O_1357,N_23893,N_23061);
or UO_1358 (O_1358,N_24875,N_23507);
and UO_1359 (O_1359,N_24051,N_24746);
and UO_1360 (O_1360,N_23426,N_22231);
nor UO_1361 (O_1361,N_24349,N_23338);
and UO_1362 (O_1362,N_24093,N_22505);
and UO_1363 (O_1363,N_24677,N_23119);
xnor UO_1364 (O_1364,N_24998,N_23944);
or UO_1365 (O_1365,N_24424,N_22838);
nand UO_1366 (O_1366,N_22619,N_22495);
and UO_1367 (O_1367,N_23563,N_23788);
nor UO_1368 (O_1368,N_24821,N_23833);
xor UO_1369 (O_1369,N_22707,N_24052);
xnor UO_1370 (O_1370,N_24343,N_23036);
nor UO_1371 (O_1371,N_24196,N_24720);
nor UO_1372 (O_1372,N_23304,N_21915);
and UO_1373 (O_1373,N_24644,N_23054);
nor UO_1374 (O_1374,N_22846,N_22644);
nor UO_1375 (O_1375,N_23707,N_22266);
and UO_1376 (O_1376,N_23522,N_24568);
xor UO_1377 (O_1377,N_24428,N_24980);
nor UO_1378 (O_1378,N_24246,N_24304);
xnor UO_1379 (O_1379,N_24829,N_23098);
xnor UO_1380 (O_1380,N_23248,N_23722);
xnor UO_1381 (O_1381,N_24973,N_22268);
nand UO_1382 (O_1382,N_23880,N_24435);
nand UO_1383 (O_1383,N_22992,N_23850);
or UO_1384 (O_1384,N_24300,N_24238);
and UO_1385 (O_1385,N_23096,N_24245);
nand UO_1386 (O_1386,N_21898,N_23046);
or UO_1387 (O_1387,N_23870,N_24794);
nor UO_1388 (O_1388,N_24018,N_22399);
or UO_1389 (O_1389,N_23942,N_23613);
or UO_1390 (O_1390,N_22078,N_24122);
xor UO_1391 (O_1391,N_23157,N_22977);
xnor UO_1392 (O_1392,N_23694,N_24777);
nand UO_1393 (O_1393,N_23653,N_24337);
xnor UO_1394 (O_1394,N_22326,N_24014);
nor UO_1395 (O_1395,N_23491,N_21890);
or UO_1396 (O_1396,N_22471,N_24900);
nand UO_1397 (O_1397,N_23658,N_24585);
and UO_1398 (O_1398,N_24154,N_22156);
and UO_1399 (O_1399,N_22103,N_24194);
nand UO_1400 (O_1400,N_22999,N_23048);
nor UO_1401 (O_1401,N_24879,N_22118);
nor UO_1402 (O_1402,N_23496,N_22526);
or UO_1403 (O_1403,N_24907,N_24740);
or UO_1404 (O_1404,N_24453,N_24458);
and UO_1405 (O_1405,N_22206,N_21906);
or UO_1406 (O_1406,N_23284,N_21910);
and UO_1407 (O_1407,N_23778,N_23353);
xnor UO_1408 (O_1408,N_23610,N_22001);
nand UO_1409 (O_1409,N_23026,N_22540);
xnor UO_1410 (O_1410,N_22965,N_24511);
nand UO_1411 (O_1411,N_22395,N_23924);
or UO_1412 (O_1412,N_24038,N_22354);
nand UO_1413 (O_1413,N_24180,N_23651);
xor UO_1414 (O_1414,N_22711,N_23593);
nor UO_1415 (O_1415,N_23999,N_21912);
or UO_1416 (O_1416,N_24839,N_22775);
and UO_1417 (O_1417,N_24258,N_21948);
xnor UO_1418 (O_1418,N_24468,N_22287);
xor UO_1419 (O_1419,N_21919,N_23950);
or UO_1420 (O_1420,N_24114,N_24357);
nor UO_1421 (O_1421,N_22790,N_24251);
nand UO_1422 (O_1422,N_22900,N_23075);
xnor UO_1423 (O_1423,N_22509,N_22028);
and UO_1424 (O_1424,N_24034,N_22337);
nand UO_1425 (O_1425,N_22249,N_22154);
xnor UO_1426 (O_1426,N_24597,N_23289);
nor UO_1427 (O_1427,N_23299,N_23989);
nor UO_1428 (O_1428,N_24926,N_23355);
and UO_1429 (O_1429,N_24150,N_24023);
xnor UO_1430 (O_1430,N_22570,N_24147);
xnor UO_1431 (O_1431,N_24911,N_22982);
nor UO_1432 (O_1432,N_23561,N_23622);
or UO_1433 (O_1433,N_23705,N_23268);
or UO_1434 (O_1434,N_24360,N_22286);
nor UO_1435 (O_1435,N_24231,N_21940);
nor UO_1436 (O_1436,N_21934,N_23747);
nand UO_1437 (O_1437,N_22988,N_23867);
nand UO_1438 (O_1438,N_23108,N_24086);
or UO_1439 (O_1439,N_22339,N_23514);
or UO_1440 (O_1440,N_24985,N_23200);
nor UO_1441 (O_1441,N_22086,N_22833);
and UO_1442 (O_1442,N_24208,N_22933);
and UO_1443 (O_1443,N_23718,N_22657);
xor UO_1444 (O_1444,N_23053,N_24004);
or UO_1445 (O_1445,N_23125,N_22718);
nor UO_1446 (O_1446,N_23178,N_24072);
nand UO_1447 (O_1447,N_23190,N_24105);
and UO_1448 (O_1448,N_24552,N_22747);
nor UO_1449 (O_1449,N_24153,N_24885);
nor UO_1450 (O_1450,N_22705,N_23230);
or UO_1451 (O_1451,N_23773,N_23047);
or UO_1452 (O_1452,N_23309,N_24719);
and UO_1453 (O_1453,N_24427,N_24448);
nor UO_1454 (O_1454,N_23111,N_23104);
xnor UO_1455 (O_1455,N_22524,N_24961);
or UO_1456 (O_1456,N_24412,N_22727);
or UO_1457 (O_1457,N_23017,N_23489);
nor UO_1458 (O_1458,N_22498,N_23391);
nor UO_1459 (O_1459,N_23113,N_23435);
or UO_1460 (O_1460,N_22142,N_24436);
xor UO_1461 (O_1461,N_24522,N_24502);
or UO_1462 (O_1462,N_23586,N_22905);
xor UO_1463 (O_1463,N_23767,N_22734);
or UO_1464 (O_1464,N_23473,N_23838);
xnor UO_1465 (O_1465,N_23115,N_23702);
and UO_1466 (O_1466,N_22239,N_24937);
or UO_1467 (O_1467,N_24204,N_22807);
nor UO_1468 (O_1468,N_24065,N_24798);
and UO_1469 (O_1469,N_22663,N_23710);
nand UO_1470 (O_1470,N_24861,N_22886);
nand UO_1471 (O_1471,N_21904,N_23117);
and UO_1472 (O_1472,N_24687,N_24076);
nand UO_1473 (O_1473,N_23014,N_22004);
and UO_1474 (O_1474,N_22065,N_23138);
and UO_1475 (O_1475,N_24183,N_22305);
or UO_1476 (O_1476,N_24872,N_23246);
or UO_1477 (O_1477,N_23116,N_22414);
and UO_1478 (O_1478,N_23957,N_24860);
and UO_1479 (O_1479,N_24309,N_21968);
nor UO_1480 (O_1480,N_24372,N_24835);
nor UO_1481 (O_1481,N_22890,N_23552);
xor UO_1482 (O_1482,N_22499,N_22063);
xnor UO_1483 (O_1483,N_22794,N_22260);
xor UO_1484 (O_1484,N_23393,N_22210);
nand UO_1485 (O_1485,N_22884,N_24735);
xnor UO_1486 (O_1486,N_24974,N_24367);
xnor UO_1487 (O_1487,N_23611,N_24683);
and UO_1488 (O_1488,N_22517,N_22412);
nor UO_1489 (O_1489,N_24274,N_24223);
or UO_1490 (O_1490,N_22234,N_23377);
nand UO_1491 (O_1491,N_23531,N_21986);
xnor UO_1492 (O_1492,N_22049,N_23254);
and UO_1493 (O_1493,N_22130,N_22984);
nand UO_1494 (O_1494,N_24665,N_23030);
nand UO_1495 (O_1495,N_23296,N_22486);
xnor UO_1496 (O_1496,N_21987,N_23493);
or UO_1497 (O_1497,N_23051,N_24784);
xor UO_1498 (O_1498,N_24411,N_24863);
and UO_1499 (O_1499,N_22104,N_24529);
nor UO_1500 (O_1500,N_23842,N_23475);
or UO_1501 (O_1501,N_23018,N_23180);
nand UO_1502 (O_1502,N_22467,N_24641);
nand UO_1503 (O_1503,N_24774,N_23411);
and UO_1504 (O_1504,N_22047,N_22067);
or UO_1505 (O_1505,N_23753,N_23389);
nand UO_1506 (O_1506,N_23274,N_24793);
and UO_1507 (O_1507,N_21970,N_23485);
xor UO_1508 (O_1508,N_22533,N_24249);
and UO_1509 (O_1509,N_23715,N_23228);
or UO_1510 (O_1510,N_22823,N_24680);
nand UO_1511 (O_1511,N_22226,N_22719);
nor UO_1512 (O_1512,N_23665,N_23862);
nor UO_1513 (O_1513,N_23764,N_22576);
and UO_1514 (O_1514,N_23388,N_24432);
nor UO_1515 (O_1515,N_24906,N_22449);
nand UO_1516 (O_1516,N_22017,N_22278);
and UO_1517 (O_1517,N_22914,N_23759);
nor UO_1518 (O_1518,N_22951,N_23161);
xnor UO_1519 (O_1519,N_22341,N_22181);
and UO_1520 (O_1520,N_24598,N_22436);
nor UO_1521 (O_1521,N_23756,N_22515);
and UO_1522 (O_1522,N_23826,N_23156);
and UO_1523 (O_1523,N_23317,N_23398);
or UO_1524 (O_1524,N_23085,N_23260);
or UO_1525 (O_1525,N_24195,N_23603);
nand UO_1526 (O_1526,N_24414,N_21931);
and UO_1527 (O_1527,N_22685,N_24621);
nand UO_1528 (O_1528,N_23326,N_24073);
xnor UO_1529 (O_1529,N_24533,N_24910);
nand UO_1530 (O_1530,N_23404,N_22849);
xor UO_1531 (O_1531,N_23765,N_23483);
nand UO_1532 (O_1532,N_22276,N_24686);
xnor UO_1533 (O_1533,N_23855,N_23385);
and UO_1534 (O_1534,N_24278,N_22021);
and UO_1535 (O_1535,N_23977,N_22676);
nor UO_1536 (O_1536,N_23578,N_23525);
nand UO_1537 (O_1537,N_22186,N_24132);
nand UO_1538 (O_1538,N_23107,N_24064);
xnor UO_1539 (O_1539,N_24454,N_23721);
and UO_1540 (O_1540,N_22964,N_24809);
and UO_1541 (O_1541,N_24162,N_23995);
xor UO_1542 (O_1542,N_22465,N_24013);
or UO_1543 (O_1543,N_22473,N_22356);
and UO_1544 (O_1544,N_22702,N_22720);
nor UO_1545 (O_1545,N_21957,N_23512);
xor UO_1546 (O_1546,N_23373,N_21937);
nand UO_1547 (O_1547,N_23938,N_24602);
or UO_1548 (O_1548,N_22901,N_22019);
and UO_1549 (O_1549,N_22560,N_24615);
nor UO_1550 (O_1550,N_22381,N_23084);
and UO_1551 (O_1551,N_24840,N_23225);
nor UO_1552 (O_1552,N_23547,N_24752);
xnor UO_1553 (O_1553,N_22388,N_22817);
nor UO_1554 (O_1554,N_23625,N_22008);
or UO_1555 (O_1555,N_23566,N_24905);
or UO_1556 (O_1556,N_22943,N_23431);
or UO_1557 (O_1557,N_22787,N_23712);
xnor UO_1558 (O_1558,N_24688,N_24333);
and UO_1559 (O_1559,N_22667,N_22758);
xor UO_1560 (O_1560,N_23945,N_22025);
xor UO_1561 (O_1561,N_24550,N_22687);
nor UO_1562 (O_1562,N_24354,N_24920);
or UO_1563 (O_1563,N_22679,N_23658);
xnor UO_1564 (O_1564,N_24759,N_24668);
and UO_1565 (O_1565,N_24261,N_23372);
and UO_1566 (O_1566,N_23745,N_23859);
and UO_1567 (O_1567,N_22295,N_24143);
nor UO_1568 (O_1568,N_24479,N_22953);
or UO_1569 (O_1569,N_22857,N_23783);
or UO_1570 (O_1570,N_23206,N_24708);
nor UO_1571 (O_1571,N_23690,N_24641);
nor UO_1572 (O_1572,N_24029,N_21981);
nor UO_1573 (O_1573,N_22646,N_24731);
nor UO_1574 (O_1574,N_24103,N_22308);
xnor UO_1575 (O_1575,N_23919,N_22965);
or UO_1576 (O_1576,N_21946,N_22593);
and UO_1577 (O_1577,N_22071,N_22976);
or UO_1578 (O_1578,N_23111,N_23138);
and UO_1579 (O_1579,N_22225,N_24285);
or UO_1580 (O_1580,N_24813,N_24912);
nor UO_1581 (O_1581,N_24933,N_23871);
nor UO_1582 (O_1582,N_22346,N_23243);
nor UO_1583 (O_1583,N_23075,N_24083);
nand UO_1584 (O_1584,N_24681,N_23215);
or UO_1585 (O_1585,N_22553,N_24504);
xnor UO_1586 (O_1586,N_23626,N_22356);
nand UO_1587 (O_1587,N_23912,N_22427);
or UO_1588 (O_1588,N_21976,N_24061);
xor UO_1589 (O_1589,N_22944,N_24444);
nor UO_1590 (O_1590,N_22989,N_22457);
nor UO_1591 (O_1591,N_23148,N_23650);
or UO_1592 (O_1592,N_24121,N_21895);
and UO_1593 (O_1593,N_22680,N_22171);
xnor UO_1594 (O_1594,N_24409,N_24236);
or UO_1595 (O_1595,N_23200,N_24609);
nor UO_1596 (O_1596,N_24347,N_22314);
or UO_1597 (O_1597,N_21983,N_24965);
nand UO_1598 (O_1598,N_21904,N_23425);
nand UO_1599 (O_1599,N_24424,N_23952);
nor UO_1600 (O_1600,N_24763,N_21923);
or UO_1601 (O_1601,N_24230,N_24183);
or UO_1602 (O_1602,N_22437,N_23634);
or UO_1603 (O_1603,N_23015,N_23445);
or UO_1604 (O_1604,N_22178,N_22402);
nor UO_1605 (O_1605,N_24822,N_22567);
nor UO_1606 (O_1606,N_24265,N_23889);
xor UO_1607 (O_1607,N_24999,N_23220);
nand UO_1608 (O_1608,N_23523,N_24649);
or UO_1609 (O_1609,N_22062,N_22971);
nor UO_1610 (O_1610,N_23960,N_23613);
xnor UO_1611 (O_1611,N_23421,N_24843);
xnor UO_1612 (O_1612,N_22167,N_22528);
nor UO_1613 (O_1613,N_23992,N_22336);
nor UO_1614 (O_1614,N_24996,N_24243);
or UO_1615 (O_1615,N_24184,N_23477);
nand UO_1616 (O_1616,N_24191,N_23073);
and UO_1617 (O_1617,N_23786,N_23305);
nand UO_1618 (O_1618,N_24722,N_23299);
and UO_1619 (O_1619,N_23742,N_21939);
and UO_1620 (O_1620,N_23166,N_21935);
nor UO_1621 (O_1621,N_24645,N_24914);
or UO_1622 (O_1622,N_24172,N_22976);
nor UO_1623 (O_1623,N_23122,N_24453);
and UO_1624 (O_1624,N_23900,N_23868);
or UO_1625 (O_1625,N_22414,N_22973);
or UO_1626 (O_1626,N_22577,N_23022);
and UO_1627 (O_1627,N_24914,N_22637);
nor UO_1628 (O_1628,N_22963,N_24592);
nor UO_1629 (O_1629,N_24962,N_23689);
or UO_1630 (O_1630,N_24234,N_22363);
xor UO_1631 (O_1631,N_22425,N_22462);
and UO_1632 (O_1632,N_23178,N_23385);
xnor UO_1633 (O_1633,N_23099,N_24181);
and UO_1634 (O_1634,N_22301,N_24729);
nand UO_1635 (O_1635,N_22585,N_24722);
or UO_1636 (O_1636,N_24514,N_24408);
xnor UO_1637 (O_1637,N_24846,N_22147);
and UO_1638 (O_1638,N_24845,N_22651);
and UO_1639 (O_1639,N_23228,N_24722);
nand UO_1640 (O_1640,N_22030,N_22647);
and UO_1641 (O_1641,N_24359,N_22127);
nor UO_1642 (O_1642,N_22257,N_24458);
nor UO_1643 (O_1643,N_23768,N_23090);
and UO_1644 (O_1644,N_22886,N_24521);
nor UO_1645 (O_1645,N_22540,N_21877);
and UO_1646 (O_1646,N_23950,N_24014);
xor UO_1647 (O_1647,N_24798,N_24535);
and UO_1648 (O_1648,N_23290,N_24048);
nor UO_1649 (O_1649,N_24126,N_23450);
and UO_1650 (O_1650,N_24340,N_22944);
or UO_1651 (O_1651,N_23319,N_22355);
and UO_1652 (O_1652,N_24597,N_22384);
or UO_1653 (O_1653,N_24679,N_22630);
or UO_1654 (O_1654,N_24011,N_24143);
xor UO_1655 (O_1655,N_23488,N_23174);
or UO_1656 (O_1656,N_24537,N_23716);
nor UO_1657 (O_1657,N_23671,N_24823);
nand UO_1658 (O_1658,N_24496,N_24445);
nand UO_1659 (O_1659,N_23466,N_24239);
nand UO_1660 (O_1660,N_23930,N_24428);
xor UO_1661 (O_1661,N_24664,N_24346);
xnor UO_1662 (O_1662,N_24483,N_24249);
nor UO_1663 (O_1663,N_24726,N_24660);
and UO_1664 (O_1664,N_24390,N_23082);
and UO_1665 (O_1665,N_22754,N_24288);
and UO_1666 (O_1666,N_23815,N_23144);
nor UO_1667 (O_1667,N_23678,N_22519);
xor UO_1668 (O_1668,N_22388,N_22386);
xnor UO_1669 (O_1669,N_24442,N_23992);
or UO_1670 (O_1670,N_23070,N_22886);
and UO_1671 (O_1671,N_23713,N_23386);
or UO_1672 (O_1672,N_24279,N_23962);
xor UO_1673 (O_1673,N_23864,N_24743);
nand UO_1674 (O_1674,N_24830,N_22346);
nor UO_1675 (O_1675,N_21989,N_21953);
nor UO_1676 (O_1676,N_23485,N_23926);
nand UO_1677 (O_1677,N_22256,N_22515);
nor UO_1678 (O_1678,N_23442,N_22230);
nand UO_1679 (O_1679,N_22975,N_23730);
and UO_1680 (O_1680,N_22787,N_24964);
and UO_1681 (O_1681,N_22386,N_22366);
or UO_1682 (O_1682,N_23111,N_22095);
nor UO_1683 (O_1683,N_24537,N_23995);
nor UO_1684 (O_1684,N_24776,N_23840);
nand UO_1685 (O_1685,N_22859,N_24831);
nand UO_1686 (O_1686,N_22467,N_22047);
nand UO_1687 (O_1687,N_22445,N_24568);
xor UO_1688 (O_1688,N_24332,N_24940);
or UO_1689 (O_1689,N_22104,N_23554);
or UO_1690 (O_1690,N_23913,N_23143);
or UO_1691 (O_1691,N_22944,N_21911);
and UO_1692 (O_1692,N_22139,N_23386);
nand UO_1693 (O_1693,N_24700,N_22783);
nand UO_1694 (O_1694,N_22811,N_21977);
xnor UO_1695 (O_1695,N_24988,N_22537);
or UO_1696 (O_1696,N_24167,N_21901);
nand UO_1697 (O_1697,N_23860,N_24856);
nor UO_1698 (O_1698,N_24732,N_24893);
nand UO_1699 (O_1699,N_22427,N_22233);
or UO_1700 (O_1700,N_22182,N_21881);
xor UO_1701 (O_1701,N_23788,N_24681);
nor UO_1702 (O_1702,N_23526,N_24848);
or UO_1703 (O_1703,N_22040,N_24244);
nor UO_1704 (O_1704,N_22893,N_22669);
nand UO_1705 (O_1705,N_23245,N_24874);
xnor UO_1706 (O_1706,N_22291,N_22202);
or UO_1707 (O_1707,N_22025,N_22318);
or UO_1708 (O_1708,N_22651,N_22103);
and UO_1709 (O_1709,N_23908,N_23851);
xor UO_1710 (O_1710,N_23432,N_22525);
or UO_1711 (O_1711,N_23996,N_22402);
nor UO_1712 (O_1712,N_24255,N_22545);
nor UO_1713 (O_1713,N_22869,N_22270);
and UO_1714 (O_1714,N_22873,N_21935);
and UO_1715 (O_1715,N_22918,N_23089);
or UO_1716 (O_1716,N_22965,N_23096);
xor UO_1717 (O_1717,N_24235,N_24633);
nor UO_1718 (O_1718,N_23680,N_24741);
xnor UO_1719 (O_1719,N_23197,N_23946);
nand UO_1720 (O_1720,N_21973,N_21961);
nor UO_1721 (O_1721,N_24490,N_24530);
nor UO_1722 (O_1722,N_24837,N_23081);
and UO_1723 (O_1723,N_23327,N_23810);
xor UO_1724 (O_1724,N_23375,N_24155);
xor UO_1725 (O_1725,N_23592,N_22750);
or UO_1726 (O_1726,N_21909,N_22764);
xor UO_1727 (O_1727,N_22773,N_24152);
or UO_1728 (O_1728,N_23856,N_22816);
and UO_1729 (O_1729,N_23745,N_22758);
and UO_1730 (O_1730,N_22991,N_23399);
and UO_1731 (O_1731,N_24549,N_24495);
nor UO_1732 (O_1732,N_24913,N_24982);
xnor UO_1733 (O_1733,N_23328,N_21927);
nand UO_1734 (O_1734,N_24283,N_22289);
or UO_1735 (O_1735,N_24351,N_21878);
and UO_1736 (O_1736,N_22041,N_24276);
and UO_1737 (O_1737,N_23835,N_22766);
xor UO_1738 (O_1738,N_23695,N_22327);
and UO_1739 (O_1739,N_23411,N_24581);
xnor UO_1740 (O_1740,N_24017,N_24155);
or UO_1741 (O_1741,N_22843,N_23343);
nor UO_1742 (O_1742,N_24327,N_24027);
xor UO_1743 (O_1743,N_22705,N_23122);
xnor UO_1744 (O_1744,N_23256,N_22490);
xor UO_1745 (O_1745,N_23018,N_22626);
xor UO_1746 (O_1746,N_24522,N_22633);
and UO_1747 (O_1747,N_23315,N_22080);
xnor UO_1748 (O_1748,N_24206,N_22307);
or UO_1749 (O_1749,N_24732,N_23445);
xnor UO_1750 (O_1750,N_23543,N_24435);
xor UO_1751 (O_1751,N_24187,N_22765);
and UO_1752 (O_1752,N_23570,N_24054);
nand UO_1753 (O_1753,N_24668,N_24928);
and UO_1754 (O_1754,N_23156,N_23779);
or UO_1755 (O_1755,N_23541,N_22647);
nand UO_1756 (O_1756,N_23005,N_23265);
or UO_1757 (O_1757,N_22346,N_22895);
and UO_1758 (O_1758,N_24891,N_24096);
nand UO_1759 (O_1759,N_23536,N_24234);
nor UO_1760 (O_1760,N_23490,N_23589);
nor UO_1761 (O_1761,N_23283,N_23036);
and UO_1762 (O_1762,N_22731,N_23240);
or UO_1763 (O_1763,N_24299,N_24301);
nor UO_1764 (O_1764,N_24736,N_22981);
or UO_1765 (O_1765,N_23949,N_23762);
nand UO_1766 (O_1766,N_24132,N_23812);
nor UO_1767 (O_1767,N_22475,N_22495);
xor UO_1768 (O_1768,N_24270,N_21980);
or UO_1769 (O_1769,N_22444,N_21889);
nand UO_1770 (O_1770,N_23586,N_23213);
or UO_1771 (O_1771,N_24014,N_24633);
xor UO_1772 (O_1772,N_24132,N_24136);
and UO_1773 (O_1773,N_23301,N_22559);
xor UO_1774 (O_1774,N_24635,N_24036);
or UO_1775 (O_1775,N_22609,N_22926);
nand UO_1776 (O_1776,N_23693,N_23352);
and UO_1777 (O_1777,N_24883,N_22980);
xor UO_1778 (O_1778,N_22009,N_22276);
or UO_1779 (O_1779,N_23619,N_23456);
nor UO_1780 (O_1780,N_23211,N_22142);
nand UO_1781 (O_1781,N_21976,N_23778);
nor UO_1782 (O_1782,N_21981,N_22527);
nor UO_1783 (O_1783,N_22563,N_22598);
nor UO_1784 (O_1784,N_24007,N_23087);
nand UO_1785 (O_1785,N_22749,N_23172);
xor UO_1786 (O_1786,N_22164,N_22789);
xnor UO_1787 (O_1787,N_23967,N_24051);
and UO_1788 (O_1788,N_23172,N_23460);
xor UO_1789 (O_1789,N_24781,N_23594);
xor UO_1790 (O_1790,N_22250,N_24426);
nand UO_1791 (O_1791,N_22911,N_23150);
xor UO_1792 (O_1792,N_23612,N_24609);
xnor UO_1793 (O_1793,N_22747,N_23491);
nand UO_1794 (O_1794,N_24629,N_22364);
nand UO_1795 (O_1795,N_22866,N_23917);
and UO_1796 (O_1796,N_23532,N_23815);
or UO_1797 (O_1797,N_24241,N_23185);
or UO_1798 (O_1798,N_22866,N_22891);
nor UO_1799 (O_1799,N_22304,N_23839);
nand UO_1800 (O_1800,N_22163,N_22269);
nor UO_1801 (O_1801,N_21929,N_24396);
and UO_1802 (O_1802,N_23734,N_22029);
nand UO_1803 (O_1803,N_22874,N_24263);
or UO_1804 (O_1804,N_23059,N_23736);
and UO_1805 (O_1805,N_22831,N_22124);
or UO_1806 (O_1806,N_22729,N_23625);
nand UO_1807 (O_1807,N_23385,N_22145);
and UO_1808 (O_1808,N_23637,N_23721);
or UO_1809 (O_1809,N_23343,N_23549);
or UO_1810 (O_1810,N_24509,N_22045);
nand UO_1811 (O_1811,N_22269,N_23140);
xnor UO_1812 (O_1812,N_23566,N_23857);
xnor UO_1813 (O_1813,N_23682,N_23121);
nor UO_1814 (O_1814,N_24082,N_24013);
and UO_1815 (O_1815,N_22393,N_23270);
nand UO_1816 (O_1816,N_24850,N_22679);
nor UO_1817 (O_1817,N_23196,N_23272);
or UO_1818 (O_1818,N_22958,N_22944);
and UO_1819 (O_1819,N_22940,N_23182);
or UO_1820 (O_1820,N_23146,N_24705);
xnor UO_1821 (O_1821,N_22795,N_23239);
or UO_1822 (O_1822,N_24446,N_24361);
nor UO_1823 (O_1823,N_22092,N_24811);
nand UO_1824 (O_1824,N_23308,N_21937);
xor UO_1825 (O_1825,N_24538,N_23124);
xor UO_1826 (O_1826,N_24265,N_24090);
xor UO_1827 (O_1827,N_23421,N_24309);
or UO_1828 (O_1828,N_23216,N_23647);
or UO_1829 (O_1829,N_22819,N_23849);
or UO_1830 (O_1830,N_23020,N_22601);
and UO_1831 (O_1831,N_23543,N_22567);
nand UO_1832 (O_1832,N_22498,N_24906);
or UO_1833 (O_1833,N_22070,N_24701);
nand UO_1834 (O_1834,N_22822,N_24422);
or UO_1835 (O_1835,N_24316,N_24416);
and UO_1836 (O_1836,N_24581,N_24459);
nor UO_1837 (O_1837,N_22830,N_24842);
or UO_1838 (O_1838,N_24677,N_24126);
nor UO_1839 (O_1839,N_24713,N_23836);
or UO_1840 (O_1840,N_24840,N_24657);
or UO_1841 (O_1841,N_22056,N_24860);
nor UO_1842 (O_1842,N_24286,N_23329);
xor UO_1843 (O_1843,N_24049,N_22203);
or UO_1844 (O_1844,N_22667,N_24207);
nor UO_1845 (O_1845,N_24197,N_22995);
nand UO_1846 (O_1846,N_24343,N_24462);
nor UO_1847 (O_1847,N_24032,N_24095);
or UO_1848 (O_1848,N_24775,N_23796);
nor UO_1849 (O_1849,N_23326,N_24440);
xor UO_1850 (O_1850,N_23767,N_24419);
nand UO_1851 (O_1851,N_21893,N_23749);
nand UO_1852 (O_1852,N_24497,N_22127);
nand UO_1853 (O_1853,N_23416,N_24063);
nor UO_1854 (O_1854,N_23498,N_23112);
xor UO_1855 (O_1855,N_22896,N_22002);
nand UO_1856 (O_1856,N_23356,N_23429);
or UO_1857 (O_1857,N_24920,N_23407);
nand UO_1858 (O_1858,N_22288,N_23864);
nor UO_1859 (O_1859,N_23421,N_22929);
nor UO_1860 (O_1860,N_23806,N_22505);
xnor UO_1861 (O_1861,N_22981,N_24526);
nor UO_1862 (O_1862,N_24217,N_22317);
xnor UO_1863 (O_1863,N_24012,N_22210);
or UO_1864 (O_1864,N_23472,N_21978);
or UO_1865 (O_1865,N_23211,N_23273);
or UO_1866 (O_1866,N_22336,N_23475);
and UO_1867 (O_1867,N_23646,N_24896);
nand UO_1868 (O_1868,N_22824,N_23884);
and UO_1869 (O_1869,N_22327,N_23426);
or UO_1870 (O_1870,N_24548,N_24113);
or UO_1871 (O_1871,N_22084,N_22502);
or UO_1872 (O_1872,N_23326,N_23767);
xor UO_1873 (O_1873,N_22282,N_23812);
and UO_1874 (O_1874,N_23566,N_24586);
and UO_1875 (O_1875,N_22465,N_23265);
and UO_1876 (O_1876,N_22262,N_24860);
nor UO_1877 (O_1877,N_23250,N_24427);
or UO_1878 (O_1878,N_24522,N_24982);
nor UO_1879 (O_1879,N_24709,N_22529);
and UO_1880 (O_1880,N_22388,N_23084);
xor UO_1881 (O_1881,N_23170,N_24943);
or UO_1882 (O_1882,N_23077,N_22567);
and UO_1883 (O_1883,N_24426,N_23927);
and UO_1884 (O_1884,N_23653,N_23254);
and UO_1885 (O_1885,N_24441,N_23833);
and UO_1886 (O_1886,N_22947,N_22560);
nand UO_1887 (O_1887,N_24481,N_24595);
xnor UO_1888 (O_1888,N_21907,N_24164);
or UO_1889 (O_1889,N_24250,N_24942);
xnor UO_1890 (O_1890,N_24503,N_23962);
or UO_1891 (O_1891,N_22896,N_22822);
or UO_1892 (O_1892,N_23855,N_22658);
nor UO_1893 (O_1893,N_21904,N_22694);
nand UO_1894 (O_1894,N_23854,N_24152);
nor UO_1895 (O_1895,N_21999,N_23813);
and UO_1896 (O_1896,N_24110,N_23320);
nor UO_1897 (O_1897,N_22453,N_23903);
nand UO_1898 (O_1898,N_22947,N_22897);
nand UO_1899 (O_1899,N_23365,N_23022);
nand UO_1900 (O_1900,N_21977,N_24864);
xor UO_1901 (O_1901,N_24457,N_24311);
or UO_1902 (O_1902,N_24345,N_23844);
or UO_1903 (O_1903,N_23092,N_23679);
nor UO_1904 (O_1904,N_24775,N_24715);
nor UO_1905 (O_1905,N_23690,N_22975);
xor UO_1906 (O_1906,N_22903,N_23205);
and UO_1907 (O_1907,N_23393,N_23707);
xnor UO_1908 (O_1908,N_23365,N_23731);
xor UO_1909 (O_1909,N_23438,N_24077);
or UO_1910 (O_1910,N_24615,N_24605);
nand UO_1911 (O_1911,N_24895,N_21986);
nand UO_1912 (O_1912,N_23289,N_23701);
xor UO_1913 (O_1913,N_23273,N_24952);
nand UO_1914 (O_1914,N_22693,N_24816);
or UO_1915 (O_1915,N_24631,N_24547);
nor UO_1916 (O_1916,N_23005,N_22354);
and UO_1917 (O_1917,N_23169,N_21968);
xor UO_1918 (O_1918,N_23765,N_23535);
xor UO_1919 (O_1919,N_24411,N_22764);
or UO_1920 (O_1920,N_24731,N_24989);
nor UO_1921 (O_1921,N_22565,N_23165);
and UO_1922 (O_1922,N_24381,N_23030);
xor UO_1923 (O_1923,N_22354,N_23749);
or UO_1924 (O_1924,N_23255,N_24848);
or UO_1925 (O_1925,N_24894,N_24150);
xnor UO_1926 (O_1926,N_24906,N_23434);
and UO_1927 (O_1927,N_23371,N_22202);
or UO_1928 (O_1928,N_23144,N_22357);
nand UO_1929 (O_1929,N_23742,N_24691);
xor UO_1930 (O_1930,N_24950,N_24567);
xnor UO_1931 (O_1931,N_23321,N_24084);
and UO_1932 (O_1932,N_23228,N_24481);
xnor UO_1933 (O_1933,N_23796,N_23803);
xor UO_1934 (O_1934,N_22737,N_24508);
nor UO_1935 (O_1935,N_22036,N_24208);
xnor UO_1936 (O_1936,N_24043,N_22909);
nand UO_1937 (O_1937,N_23017,N_24234);
nor UO_1938 (O_1938,N_23274,N_23701);
and UO_1939 (O_1939,N_23117,N_22664);
nor UO_1940 (O_1940,N_24208,N_23567);
nor UO_1941 (O_1941,N_23103,N_24288);
xor UO_1942 (O_1942,N_22344,N_24900);
or UO_1943 (O_1943,N_24483,N_23033);
and UO_1944 (O_1944,N_22228,N_22996);
nor UO_1945 (O_1945,N_22006,N_23458);
or UO_1946 (O_1946,N_23446,N_22913);
or UO_1947 (O_1947,N_22192,N_23908);
xor UO_1948 (O_1948,N_23306,N_24466);
or UO_1949 (O_1949,N_24145,N_24896);
or UO_1950 (O_1950,N_24560,N_24237);
or UO_1951 (O_1951,N_23061,N_24887);
or UO_1952 (O_1952,N_24613,N_24047);
or UO_1953 (O_1953,N_23737,N_23380);
and UO_1954 (O_1954,N_23807,N_23046);
nor UO_1955 (O_1955,N_24180,N_24354);
nor UO_1956 (O_1956,N_22582,N_22908);
nor UO_1957 (O_1957,N_23168,N_21999);
nand UO_1958 (O_1958,N_23886,N_22272);
and UO_1959 (O_1959,N_24312,N_24867);
or UO_1960 (O_1960,N_23602,N_24928);
xnor UO_1961 (O_1961,N_23885,N_24078);
nor UO_1962 (O_1962,N_22357,N_23824);
nor UO_1963 (O_1963,N_22754,N_24888);
or UO_1964 (O_1964,N_21952,N_23879);
or UO_1965 (O_1965,N_23715,N_21876);
nand UO_1966 (O_1966,N_22488,N_23998);
or UO_1967 (O_1967,N_24456,N_24700);
or UO_1968 (O_1968,N_23459,N_22190);
or UO_1969 (O_1969,N_23301,N_22843);
nor UO_1970 (O_1970,N_24089,N_22617);
xnor UO_1971 (O_1971,N_24033,N_22242);
nand UO_1972 (O_1972,N_23107,N_23738);
nand UO_1973 (O_1973,N_22650,N_24511);
or UO_1974 (O_1974,N_22825,N_22261);
xor UO_1975 (O_1975,N_23298,N_24568);
and UO_1976 (O_1976,N_22930,N_23440);
and UO_1977 (O_1977,N_22499,N_24405);
xor UO_1978 (O_1978,N_23311,N_22096);
xor UO_1979 (O_1979,N_23449,N_22738);
nand UO_1980 (O_1980,N_22411,N_24907);
xnor UO_1981 (O_1981,N_23013,N_22365);
nand UO_1982 (O_1982,N_24505,N_23866);
nand UO_1983 (O_1983,N_23180,N_22360);
nand UO_1984 (O_1984,N_24515,N_24165);
xor UO_1985 (O_1985,N_24565,N_23187);
and UO_1986 (O_1986,N_21892,N_22177);
nand UO_1987 (O_1987,N_23079,N_23928);
xnor UO_1988 (O_1988,N_24009,N_23249);
or UO_1989 (O_1989,N_23891,N_23577);
or UO_1990 (O_1990,N_22669,N_22310);
nand UO_1991 (O_1991,N_24842,N_23571);
xnor UO_1992 (O_1992,N_23129,N_21970);
nand UO_1993 (O_1993,N_24150,N_23704);
xor UO_1994 (O_1994,N_24806,N_23497);
or UO_1995 (O_1995,N_21909,N_24359);
xnor UO_1996 (O_1996,N_23197,N_23918);
or UO_1997 (O_1997,N_22334,N_22282);
nor UO_1998 (O_1998,N_24731,N_23533);
or UO_1999 (O_1999,N_23518,N_23004);
and UO_2000 (O_2000,N_23622,N_24525);
xor UO_2001 (O_2001,N_23962,N_23252);
and UO_2002 (O_2002,N_24691,N_23678);
or UO_2003 (O_2003,N_24887,N_22181);
nand UO_2004 (O_2004,N_24761,N_22165);
or UO_2005 (O_2005,N_22411,N_22320);
nor UO_2006 (O_2006,N_24883,N_24570);
nand UO_2007 (O_2007,N_23757,N_22302);
nand UO_2008 (O_2008,N_24914,N_23332);
xor UO_2009 (O_2009,N_23308,N_24099);
and UO_2010 (O_2010,N_24379,N_23928);
nor UO_2011 (O_2011,N_24618,N_22375);
or UO_2012 (O_2012,N_23400,N_23731);
xor UO_2013 (O_2013,N_23712,N_23089);
or UO_2014 (O_2014,N_24684,N_24381);
nand UO_2015 (O_2015,N_22930,N_24834);
or UO_2016 (O_2016,N_22254,N_22065);
and UO_2017 (O_2017,N_23317,N_23893);
or UO_2018 (O_2018,N_24823,N_23030);
xor UO_2019 (O_2019,N_24674,N_22846);
and UO_2020 (O_2020,N_24720,N_23446);
nor UO_2021 (O_2021,N_22857,N_22732);
or UO_2022 (O_2022,N_24178,N_23760);
or UO_2023 (O_2023,N_23921,N_23350);
nand UO_2024 (O_2024,N_24503,N_23227);
or UO_2025 (O_2025,N_22469,N_22495);
and UO_2026 (O_2026,N_22540,N_24165);
or UO_2027 (O_2027,N_24207,N_24111);
or UO_2028 (O_2028,N_23908,N_21999);
and UO_2029 (O_2029,N_24362,N_24980);
or UO_2030 (O_2030,N_23836,N_24083);
or UO_2031 (O_2031,N_23475,N_24719);
xnor UO_2032 (O_2032,N_22775,N_23071);
nand UO_2033 (O_2033,N_24829,N_23369);
nand UO_2034 (O_2034,N_23691,N_24560);
and UO_2035 (O_2035,N_23368,N_24205);
nand UO_2036 (O_2036,N_22179,N_24914);
nand UO_2037 (O_2037,N_23824,N_23592);
xor UO_2038 (O_2038,N_23022,N_22831);
or UO_2039 (O_2039,N_24216,N_22173);
and UO_2040 (O_2040,N_22138,N_23785);
xor UO_2041 (O_2041,N_24024,N_21965);
nor UO_2042 (O_2042,N_22176,N_24927);
or UO_2043 (O_2043,N_23875,N_22626);
and UO_2044 (O_2044,N_23511,N_24655);
nand UO_2045 (O_2045,N_22226,N_24104);
or UO_2046 (O_2046,N_23797,N_23964);
nand UO_2047 (O_2047,N_22208,N_22895);
nor UO_2048 (O_2048,N_22237,N_22396);
or UO_2049 (O_2049,N_24580,N_24001);
xnor UO_2050 (O_2050,N_24077,N_23714);
or UO_2051 (O_2051,N_22538,N_22467);
and UO_2052 (O_2052,N_23758,N_22309);
xnor UO_2053 (O_2053,N_22694,N_24312);
nand UO_2054 (O_2054,N_22719,N_23861);
nand UO_2055 (O_2055,N_21951,N_23084);
or UO_2056 (O_2056,N_22184,N_23605);
nor UO_2057 (O_2057,N_23473,N_24115);
and UO_2058 (O_2058,N_22377,N_22536);
nand UO_2059 (O_2059,N_22588,N_22647);
xor UO_2060 (O_2060,N_23087,N_23003);
nor UO_2061 (O_2061,N_22054,N_23352);
nand UO_2062 (O_2062,N_22779,N_22818);
nand UO_2063 (O_2063,N_24725,N_24964);
nand UO_2064 (O_2064,N_21978,N_22955);
or UO_2065 (O_2065,N_23358,N_24549);
nand UO_2066 (O_2066,N_23346,N_24605);
and UO_2067 (O_2067,N_22649,N_23671);
and UO_2068 (O_2068,N_24676,N_22371);
or UO_2069 (O_2069,N_24259,N_22006);
nor UO_2070 (O_2070,N_22451,N_24592);
nand UO_2071 (O_2071,N_23730,N_23118);
or UO_2072 (O_2072,N_24747,N_23930);
and UO_2073 (O_2073,N_22001,N_24212);
and UO_2074 (O_2074,N_23948,N_22287);
xor UO_2075 (O_2075,N_23818,N_23026);
and UO_2076 (O_2076,N_24791,N_23862);
nor UO_2077 (O_2077,N_22158,N_23825);
or UO_2078 (O_2078,N_23310,N_24331);
and UO_2079 (O_2079,N_24047,N_22996);
or UO_2080 (O_2080,N_22398,N_24520);
nor UO_2081 (O_2081,N_24678,N_22148);
nor UO_2082 (O_2082,N_24833,N_24719);
nor UO_2083 (O_2083,N_23481,N_24400);
nand UO_2084 (O_2084,N_24376,N_23611);
nor UO_2085 (O_2085,N_23181,N_24732);
xor UO_2086 (O_2086,N_23959,N_23628);
or UO_2087 (O_2087,N_23461,N_21878);
nand UO_2088 (O_2088,N_22278,N_22911);
nor UO_2089 (O_2089,N_22969,N_23668);
and UO_2090 (O_2090,N_22990,N_22044);
nand UO_2091 (O_2091,N_23634,N_23317);
nand UO_2092 (O_2092,N_22709,N_22288);
nand UO_2093 (O_2093,N_23957,N_23060);
nor UO_2094 (O_2094,N_24134,N_22668);
nand UO_2095 (O_2095,N_22178,N_23509);
xnor UO_2096 (O_2096,N_21938,N_24992);
and UO_2097 (O_2097,N_22533,N_22528);
or UO_2098 (O_2098,N_21943,N_22656);
nand UO_2099 (O_2099,N_23807,N_23951);
or UO_2100 (O_2100,N_21978,N_24207);
and UO_2101 (O_2101,N_24327,N_22646);
xnor UO_2102 (O_2102,N_22271,N_22819);
nor UO_2103 (O_2103,N_23941,N_24149);
nor UO_2104 (O_2104,N_23666,N_23352);
nor UO_2105 (O_2105,N_23378,N_24474);
and UO_2106 (O_2106,N_24209,N_22631);
or UO_2107 (O_2107,N_23863,N_23496);
nor UO_2108 (O_2108,N_24410,N_23713);
and UO_2109 (O_2109,N_24137,N_23535);
nor UO_2110 (O_2110,N_23838,N_23494);
and UO_2111 (O_2111,N_21889,N_23492);
and UO_2112 (O_2112,N_23971,N_24625);
xor UO_2113 (O_2113,N_23667,N_24114);
and UO_2114 (O_2114,N_22704,N_22524);
xor UO_2115 (O_2115,N_24320,N_21924);
xnor UO_2116 (O_2116,N_22487,N_22536);
nand UO_2117 (O_2117,N_24807,N_22558);
nor UO_2118 (O_2118,N_24205,N_24804);
or UO_2119 (O_2119,N_23615,N_23396);
and UO_2120 (O_2120,N_24579,N_24306);
nand UO_2121 (O_2121,N_23972,N_23343);
xnor UO_2122 (O_2122,N_23903,N_21997);
and UO_2123 (O_2123,N_22558,N_24327);
nor UO_2124 (O_2124,N_24181,N_23545);
nor UO_2125 (O_2125,N_23399,N_24715);
xor UO_2126 (O_2126,N_24906,N_24106);
nand UO_2127 (O_2127,N_23516,N_22659);
nand UO_2128 (O_2128,N_22932,N_24425);
or UO_2129 (O_2129,N_22911,N_22401);
or UO_2130 (O_2130,N_23750,N_23528);
xor UO_2131 (O_2131,N_24999,N_23700);
xor UO_2132 (O_2132,N_22025,N_23621);
or UO_2133 (O_2133,N_23090,N_23806);
nor UO_2134 (O_2134,N_22180,N_24894);
nand UO_2135 (O_2135,N_23871,N_23473);
and UO_2136 (O_2136,N_24009,N_22360);
or UO_2137 (O_2137,N_24155,N_22784);
nand UO_2138 (O_2138,N_24081,N_24895);
xnor UO_2139 (O_2139,N_22123,N_23909);
nor UO_2140 (O_2140,N_22694,N_23645);
or UO_2141 (O_2141,N_22373,N_24471);
nand UO_2142 (O_2142,N_24349,N_24371);
xnor UO_2143 (O_2143,N_24570,N_21983);
nor UO_2144 (O_2144,N_23435,N_21963);
nor UO_2145 (O_2145,N_23158,N_24658);
or UO_2146 (O_2146,N_24512,N_22872);
nand UO_2147 (O_2147,N_23425,N_22396);
or UO_2148 (O_2148,N_24640,N_23878);
xnor UO_2149 (O_2149,N_24007,N_22657);
or UO_2150 (O_2150,N_23624,N_24512);
or UO_2151 (O_2151,N_21950,N_22406);
and UO_2152 (O_2152,N_24645,N_22970);
xnor UO_2153 (O_2153,N_23934,N_22500);
and UO_2154 (O_2154,N_24612,N_23385);
nand UO_2155 (O_2155,N_23027,N_22290);
and UO_2156 (O_2156,N_24218,N_23090);
nand UO_2157 (O_2157,N_24508,N_22932);
nand UO_2158 (O_2158,N_24087,N_23682);
nor UO_2159 (O_2159,N_22218,N_24920);
nand UO_2160 (O_2160,N_22442,N_24048);
nand UO_2161 (O_2161,N_23166,N_23407);
nor UO_2162 (O_2162,N_22461,N_22239);
or UO_2163 (O_2163,N_24405,N_23889);
and UO_2164 (O_2164,N_24609,N_22432);
or UO_2165 (O_2165,N_23078,N_22763);
nand UO_2166 (O_2166,N_24171,N_21951);
xnor UO_2167 (O_2167,N_22446,N_24337);
nand UO_2168 (O_2168,N_22867,N_23127);
or UO_2169 (O_2169,N_24943,N_22966);
xnor UO_2170 (O_2170,N_22611,N_22154);
and UO_2171 (O_2171,N_23551,N_23994);
and UO_2172 (O_2172,N_24936,N_22088);
and UO_2173 (O_2173,N_23405,N_22690);
or UO_2174 (O_2174,N_23406,N_24672);
and UO_2175 (O_2175,N_24495,N_23421);
nor UO_2176 (O_2176,N_23087,N_23227);
or UO_2177 (O_2177,N_22343,N_23251);
and UO_2178 (O_2178,N_24818,N_23022);
xnor UO_2179 (O_2179,N_24939,N_23669);
or UO_2180 (O_2180,N_24854,N_22458);
nor UO_2181 (O_2181,N_24776,N_24841);
nor UO_2182 (O_2182,N_24859,N_23929);
or UO_2183 (O_2183,N_24182,N_22138);
nor UO_2184 (O_2184,N_23584,N_24887);
and UO_2185 (O_2185,N_22124,N_22712);
and UO_2186 (O_2186,N_22660,N_23524);
or UO_2187 (O_2187,N_24850,N_24158);
xnor UO_2188 (O_2188,N_22737,N_23945);
nand UO_2189 (O_2189,N_22603,N_23042);
nor UO_2190 (O_2190,N_24825,N_22092);
or UO_2191 (O_2191,N_23595,N_23574);
xor UO_2192 (O_2192,N_23989,N_22391);
nand UO_2193 (O_2193,N_22489,N_24329);
nor UO_2194 (O_2194,N_22301,N_24015);
nand UO_2195 (O_2195,N_21949,N_23058);
nand UO_2196 (O_2196,N_22114,N_23538);
nor UO_2197 (O_2197,N_22971,N_23785);
nand UO_2198 (O_2198,N_23765,N_22534);
xor UO_2199 (O_2199,N_23803,N_23013);
and UO_2200 (O_2200,N_24904,N_24333);
nor UO_2201 (O_2201,N_23301,N_24363);
and UO_2202 (O_2202,N_24008,N_23917);
nand UO_2203 (O_2203,N_24589,N_22509);
nand UO_2204 (O_2204,N_23407,N_22847);
nor UO_2205 (O_2205,N_24692,N_22304);
xor UO_2206 (O_2206,N_22770,N_22250);
nor UO_2207 (O_2207,N_22675,N_24683);
nand UO_2208 (O_2208,N_22375,N_24815);
nor UO_2209 (O_2209,N_24361,N_24482);
nor UO_2210 (O_2210,N_22936,N_22444);
xnor UO_2211 (O_2211,N_24685,N_21973);
and UO_2212 (O_2212,N_23795,N_22576);
nor UO_2213 (O_2213,N_23963,N_23366);
nand UO_2214 (O_2214,N_22165,N_24156);
and UO_2215 (O_2215,N_22505,N_23213);
xor UO_2216 (O_2216,N_22881,N_23554);
and UO_2217 (O_2217,N_23360,N_22927);
and UO_2218 (O_2218,N_24434,N_22586);
nand UO_2219 (O_2219,N_23556,N_22242);
and UO_2220 (O_2220,N_24425,N_23452);
nand UO_2221 (O_2221,N_24854,N_22053);
or UO_2222 (O_2222,N_22804,N_23522);
nand UO_2223 (O_2223,N_24240,N_24667);
nor UO_2224 (O_2224,N_23461,N_24844);
nor UO_2225 (O_2225,N_21946,N_24935);
and UO_2226 (O_2226,N_23998,N_23132);
nand UO_2227 (O_2227,N_23637,N_24685);
or UO_2228 (O_2228,N_22663,N_24214);
nor UO_2229 (O_2229,N_22789,N_23708);
nor UO_2230 (O_2230,N_22349,N_24124);
nor UO_2231 (O_2231,N_22305,N_22260);
or UO_2232 (O_2232,N_24356,N_23539);
xor UO_2233 (O_2233,N_24439,N_24700);
or UO_2234 (O_2234,N_24388,N_24597);
and UO_2235 (O_2235,N_24492,N_23921);
and UO_2236 (O_2236,N_22799,N_23648);
xnor UO_2237 (O_2237,N_23918,N_23209);
nor UO_2238 (O_2238,N_23938,N_23920);
xor UO_2239 (O_2239,N_22434,N_22296);
and UO_2240 (O_2240,N_22784,N_23011);
nand UO_2241 (O_2241,N_22932,N_23425);
nor UO_2242 (O_2242,N_24390,N_22820);
nor UO_2243 (O_2243,N_24769,N_22961);
or UO_2244 (O_2244,N_23471,N_22189);
or UO_2245 (O_2245,N_23939,N_22596);
or UO_2246 (O_2246,N_24385,N_24219);
or UO_2247 (O_2247,N_23196,N_21906);
and UO_2248 (O_2248,N_22138,N_23661);
xor UO_2249 (O_2249,N_22030,N_23998);
nand UO_2250 (O_2250,N_22125,N_24837);
xnor UO_2251 (O_2251,N_24277,N_23349);
xnor UO_2252 (O_2252,N_22565,N_21999);
or UO_2253 (O_2253,N_24947,N_22481);
nand UO_2254 (O_2254,N_23700,N_23316);
xor UO_2255 (O_2255,N_22618,N_23828);
and UO_2256 (O_2256,N_23250,N_23879);
nand UO_2257 (O_2257,N_23130,N_22966);
and UO_2258 (O_2258,N_22546,N_22805);
xnor UO_2259 (O_2259,N_23358,N_22476);
nor UO_2260 (O_2260,N_23266,N_22867);
or UO_2261 (O_2261,N_24331,N_22427);
or UO_2262 (O_2262,N_23169,N_22093);
and UO_2263 (O_2263,N_24623,N_21959);
and UO_2264 (O_2264,N_23441,N_22450);
nand UO_2265 (O_2265,N_24977,N_24119);
xnor UO_2266 (O_2266,N_24143,N_23409);
or UO_2267 (O_2267,N_23104,N_23059);
or UO_2268 (O_2268,N_24230,N_23113);
and UO_2269 (O_2269,N_24324,N_23536);
and UO_2270 (O_2270,N_23815,N_21988);
nand UO_2271 (O_2271,N_23093,N_23502);
nand UO_2272 (O_2272,N_24097,N_22686);
or UO_2273 (O_2273,N_22388,N_23664);
or UO_2274 (O_2274,N_24733,N_22024);
and UO_2275 (O_2275,N_23756,N_24017);
and UO_2276 (O_2276,N_24990,N_24517);
and UO_2277 (O_2277,N_23070,N_23002);
and UO_2278 (O_2278,N_23258,N_23842);
and UO_2279 (O_2279,N_21993,N_23707);
or UO_2280 (O_2280,N_24326,N_22343);
xnor UO_2281 (O_2281,N_22770,N_24533);
xor UO_2282 (O_2282,N_22114,N_23837);
xnor UO_2283 (O_2283,N_22232,N_24553);
nand UO_2284 (O_2284,N_22526,N_22745);
or UO_2285 (O_2285,N_24651,N_24814);
nand UO_2286 (O_2286,N_23713,N_23641);
or UO_2287 (O_2287,N_23461,N_23210);
nand UO_2288 (O_2288,N_23530,N_23579);
xnor UO_2289 (O_2289,N_22641,N_22243);
nand UO_2290 (O_2290,N_24790,N_22750);
and UO_2291 (O_2291,N_24462,N_23536);
nand UO_2292 (O_2292,N_22493,N_23025);
nor UO_2293 (O_2293,N_24133,N_24950);
nor UO_2294 (O_2294,N_23369,N_21957);
nor UO_2295 (O_2295,N_22639,N_24044);
nor UO_2296 (O_2296,N_23130,N_23533);
nand UO_2297 (O_2297,N_22473,N_22067);
or UO_2298 (O_2298,N_22935,N_22182);
xnor UO_2299 (O_2299,N_23047,N_23217);
nor UO_2300 (O_2300,N_24921,N_24531);
and UO_2301 (O_2301,N_23661,N_23754);
or UO_2302 (O_2302,N_23333,N_23791);
nor UO_2303 (O_2303,N_23148,N_24884);
nand UO_2304 (O_2304,N_22239,N_23848);
nand UO_2305 (O_2305,N_22959,N_24581);
or UO_2306 (O_2306,N_24024,N_24820);
or UO_2307 (O_2307,N_23740,N_23656);
xor UO_2308 (O_2308,N_24002,N_23445);
xor UO_2309 (O_2309,N_23719,N_23503);
nand UO_2310 (O_2310,N_24785,N_24352);
and UO_2311 (O_2311,N_24650,N_23407);
or UO_2312 (O_2312,N_24305,N_22877);
nor UO_2313 (O_2313,N_23001,N_23582);
or UO_2314 (O_2314,N_22340,N_24296);
and UO_2315 (O_2315,N_22352,N_22097);
xnor UO_2316 (O_2316,N_24626,N_23844);
nor UO_2317 (O_2317,N_24457,N_22417);
xor UO_2318 (O_2318,N_24930,N_24358);
nor UO_2319 (O_2319,N_24555,N_24065);
or UO_2320 (O_2320,N_22050,N_24698);
or UO_2321 (O_2321,N_22946,N_23539);
and UO_2322 (O_2322,N_22540,N_22346);
xnor UO_2323 (O_2323,N_24382,N_24283);
or UO_2324 (O_2324,N_24401,N_22754);
or UO_2325 (O_2325,N_24416,N_24812);
nor UO_2326 (O_2326,N_23067,N_23432);
and UO_2327 (O_2327,N_24601,N_22207);
nor UO_2328 (O_2328,N_23157,N_24288);
nor UO_2329 (O_2329,N_22526,N_23423);
nand UO_2330 (O_2330,N_23953,N_23516);
nand UO_2331 (O_2331,N_24743,N_22255);
nand UO_2332 (O_2332,N_22346,N_23276);
xnor UO_2333 (O_2333,N_23380,N_22326);
nor UO_2334 (O_2334,N_23323,N_24749);
nor UO_2335 (O_2335,N_24915,N_24129);
nand UO_2336 (O_2336,N_23341,N_23943);
or UO_2337 (O_2337,N_24020,N_23068);
and UO_2338 (O_2338,N_22565,N_23356);
nor UO_2339 (O_2339,N_22709,N_23192);
xnor UO_2340 (O_2340,N_24080,N_23881);
nand UO_2341 (O_2341,N_23751,N_22535);
or UO_2342 (O_2342,N_22227,N_24800);
nand UO_2343 (O_2343,N_24043,N_23285);
or UO_2344 (O_2344,N_24726,N_22184);
and UO_2345 (O_2345,N_24934,N_24528);
or UO_2346 (O_2346,N_24092,N_22719);
xor UO_2347 (O_2347,N_21902,N_23034);
nand UO_2348 (O_2348,N_23405,N_22417);
nand UO_2349 (O_2349,N_22162,N_23905);
nand UO_2350 (O_2350,N_22783,N_24633);
nor UO_2351 (O_2351,N_22400,N_22092);
nor UO_2352 (O_2352,N_23284,N_24584);
nand UO_2353 (O_2353,N_22222,N_23138);
or UO_2354 (O_2354,N_21942,N_23196);
or UO_2355 (O_2355,N_24658,N_24923);
or UO_2356 (O_2356,N_23476,N_24963);
or UO_2357 (O_2357,N_22768,N_23577);
and UO_2358 (O_2358,N_23240,N_22268);
nand UO_2359 (O_2359,N_24238,N_24162);
xnor UO_2360 (O_2360,N_21931,N_22499);
nand UO_2361 (O_2361,N_22161,N_21992);
or UO_2362 (O_2362,N_22451,N_22737);
and UO_2363 (O_2363,N_23892,N_24820);
xnor UO_2364 (O_2364,N_23771,N_24307);
nor UO_2365 (O_2365,N_22362,N_23585);
or UO_2366 (O_2366,N_23337,N_22084);
nor UO_2367 (O_2367,N_24212,N_23733);
or UO_2368 (O_2368,N_24178,N_24992);
or UO_2369 (O_2369,N_23768,N_23554);
nor UO_2370 (O_2370,N_24623,N_23221);
nand UO_2371 (O_2371,N_23860,N_23331);
or UO_2372 (O_2372,N_22649,N_24519);
or UO_2373 (O_2373,N_23441,N_24295);
nor UO_2374 (O_2374,N_23739,N_22986);
nand UO_2375 (O_2375,N_23028,N_22061);
nand UO_2376 (O_2376,N_22481,N_23450);
xnor UO_2377 (O_2377,N_24092,N_23064);
nor UO_2378 (O_2378,N_22936,N_24276);
and UO_2379 (O_2379,N_24473,N_24703);
nor UO_2380 (O_2380,N_23215,N_24483);
nand UO_2381 (O_2381,N_24134,N_23711);
nor UO_2382 (O_2382,N_22627,N_23185);
nand UO_2383 (O_2383,N_22679,N_24400);
nor UO_2384 (O_2384,N_21969,N_24756);
xnor UO_2385 (O_2385,N_22624,N_21926);
or UO_2386 (O_2386,N_22479,N_24951);
nor UO_2387 (O_2387,N_24723,N_24312);
nand UO_2388 (O_2388,N_23610,N_24524);
nor UO_2389 (O_2389,N_22765,N_22266);
nor UO_2390 (O_2390,N_23677,N_23896);
or UO_2391 (O_2391,N_23785,N_23498);
nand UO_2392 (O_2392,N_24140,N_24855);
nand UO_2393 (O_2393,N_23717,N_23998);
nand UO_2394 (O_2394,N_22975,N_23937);
xnor UO_2395 (O_2395,N_24233,N_23696);
xnor UO_2396 (O_2396,N_23975,N_22354);
xnor UO_2397 (O_2397,N_24745,N_24179);
nand UO_2398 (O_2398,N_24981,N_23769);
nand UO_2399 (O_2399,N_24737,N_23749);
nor UO_2400 (O_2400,N_23221,N_24794);
xnor UO_2401 (O_2401,N_23911,N_23447);
nand UO_2402 (O_2402,N_23803,N_22596);
nor UO_2403 (O_2403,N_24823,N_22608);
nor UO_2404 (O_2404,N_24321,N_24853);
or UO_2405 (O_2405,N_21969,N_24902);
nor UO_2406 (O_2406,N_23359,N_22669);
or UO_2407 (O_2407,N_24319,N_24932);
and UO_2408 (O_2408,N_23186,N_23808);
or UO_2409 (O_2409,N_22975,N_22183);
nor UO_2410 (O_2410,N_23769,N_23085);
xor UO_2411 (O_2411,N_23580,N_22798);
xor UO_2412 (O_2412,N_24911,N_22338);
and UO_2413 (O_2413,N_24205,N_23579);
xor UO_2414 (O_2414,N_24276,N_24383);
xor UO_2415 (O_2415,N_22556,N_23531);
and UO_2416 (O_2416,N_23629,N_23538);
xnor UO_2417 (O_2417,N_24632,N_21923);
nor UO_2418 (O_2418,N_21995,N_22257);
xor UO_2419 (O_2419,N_23704,N_23406);
and UO_2420 (O_2420,N_23942,N_21935);
nand UO_2421 (O_2421,N_24957,N_22426);
nor UO_2422 (O_2422,N_22926,N_22819);
and UO_2423 (O_2423,N_24635,N_24823);
nor UO_2424 (O_2424,N_22997,N_22542);
and UO_2425 (O_2425,N_22925,N_23861);
nand UO_2426 (O_2426,N_24583,N_23008);
or UO_2427 (O_2427,N_24842,N_23138);
and UO_2428 (O_2428,N_22438,N_23285);
nand UO_2429 (O_2429,N_24312,N_24779);
nor UO_2430 (O_2430,N_24664,N_24166);
or UO_2431 (O_2431,N_24608,N_24110);
and UO_2432 (O_2432,N_22713,N_23966);
nor UO_2433 (O_2433,N_23584,N_22607);
nor UO_2434 (O_2434,N_23898,N_24170);
and UO_2435 (O_2435,N_22110,N_23211);
and UO_2436 (O_2436,N_24950,N_22412);
or UO_2437 (O_2437,N_24409,N_22474);
and UO_2438 (O_2438,N_23557,N_22017);
nor UO_2439 (O_2439,N_21936,N_23857);
nand UO_2440 (O_2440,N_22319,N_23139);
and UO_2441 (O_2441,N_24996,N_24357);
and UO_2442 (O_2442,N_22674,N_23523);
and UO_2443 (O_2443,N_23292,N_23623);
or UO_2444 (O_2444,N_22336,N_23574);
nand UO_2445 (O_2445,N_24168,N_22646);
and UO_2446 (O_2446,N_22790,N_22769);
nand UO_2447 (O_2447,N_23304,N_22966);
or UO_2448 (O_2448,N_23960,N_23049);
nor UO_2449 (O_2449,N_22607,N_22144);
xor UO_2450 (O_2450,N_23249,N_24780);
xor UO_2451 (O_2451,N_23146,N_22844);
or UO_2452 (O_2452,N_23364,N_23593);
nor UO_2453 (O_2453,N_24594,N_22660);
nor UO_2454 (O_2454,N_23939,N_23878);
xor UO_2455 (O_2455,N_24657,N_24554);
and UO_2456 (O_2456,N_23761,N_22460);
and UO_2457 (O_2457,N_22900,N_22544);
nor UO_2458 (O_2458,N_24437,N_24702);
and UO_2459 (O_2459,N_23320,N_22536);
or UO_2460 (O_2460,N_23216,N_22672);
and UO_2461 (O_2461,N_23611,N_24160);
nor UO_2462 (O_2462,N_22434,N_22332);
or UO_2463 (O_2463,N_24848,N_23606);
nor UO_2464 (O_2464,N_22121,N_23144);
nand UO_2465 (O_2465,N_23170,N_23238);
nor UO_2466 (O_2466,N_22931,N_23762);
nand UO_2467 (O_2467,N_24429,N_24092);
or UO_2468 (O_2468,N_24767,N_24630);
nand UO_2469 (O_2469,N_22252,N_22452);
or UO_2470 (O_2470,N_24972,N_21988);
nand UO_2471 (O_2471,N_22789,N_23417);
nand UO_2472 (O_2472,N_22703,N_23519);
and UO_2473 (O_2473,N_24708,N_24709);
nor UO_2474 (O_2474,N_23873,N_22968);
nor UO_2475 (O_2475,N_23192,N_22349);
xor UO_2476 (O_2476,N_24209,N_24700);
nand UO_2477 (O_2477,N_24703,N_22453);
and UO_2478 (O_2478,N_22039,N_24264);
nand UO_2479 (O_2479,N_23160,N_22357);
xor UO_2480 (O_2480,N_24107,N_24555);
xnor UO_2481 (O_2481,N_22950,N_22568);
or UO_2482 (O_2482,N_22911,N_24583);
nand UO_2483 (O_2483,N_23513,N_22463);
and UO_2484 (O_2484,N_22632,N_24173);
or UO_2485 (O_2485,N_23287,N_23349);
nor UO_2486 (O_2486,N_23219,N_24334);
nand UO_2487 (O_2487,N_24472,N_23900);
or UO_2488 (O_2488,N_23765,N_23738);
and UO_2489 (O_2489,N_24294,N_23910);
and UO_2490 (O_2490,N_22488,N_24091);
xnor UO_2491 (O_2491,N_22451,N_22903);
and UO_2492 (O_2492,N_24115,N_22976);
and UO_2493 (O_2493,N_23768,N_23395);
or UO_2494 (O_2494,N_24529,N_24649);
nor UO_2495 (O_2495,N_22267,N_23083);
or UO_2496 (O_2496,N_24596,N_24774);
xor UO_2497 (O_2497,N_22480,N_23282);
nand UO_2498 (O_2498,N_24891,N_22847);
nor UO_2499 (O_2499,N_24261,N_22599);
or UO_2500 (O_2500,N_24829,N_22280);
or UO_2501 (O_2501,N_24444,N_21993);
xor UO_2502 (O_2502,N_24631,N_22362);
nor UO_2503 (O_2503,N_22784,N_23266);
nor UO_2504 (O_2504,N_23494,N_22169);
xor UO_2505 (O_2505,N_23192,N_22271);
and UO_2506 (O_2506,N_23825,N_23191);
nand UO_2507 (O_2507,N_24655,N_23764);
nor UO_2508 (O_2508,N_23415,N_22496);
nor UO_2509 (O_2509,N_22155,N_24363);
nor UO_2510 (O_2510,N_24839,N_23362);
or UO_2511 (O_2511,N_22310,N_24054);
xnor UO_2512 (O_2512,N_23427,N_21879);
and UO_2513 (O_2513,N_22258,N_21884);
and UO_2514 (O_2514,N_22798,N_23006);
nand UO_2515 (O_2515,N_23293,N_22488);
and UO_2516 (O_2516,N_22820,N_22700);
nor UO_2517 (O_2517,N_24140,N_24388);
or UO_2518 (O_2518,N_22994,N_23083);
nand UO_2519 (O_2519,N_23490,N_23259);
nand UO_2520 (O_2520,N_23780,N_24248);
nor UO_2521 (O_2521,N_22658,N_22846);
nor UO_2522 (O_2522,N_22540,N_23001);
or UO_2523 (O_2523,N_23093,N_23647);
nand UO_2524 (O_2524,N_22115,N_24501);
xnor UO_2525 (O_2525,N_23007,N_22428);
and UO_2526 (O_2526,N_24084,N_24638);
xor UO_2527 (O_2527,N_24606,N_23151);
nand UO_2528 (O_2528,N_23298,N_24481);
and UO_2529 (O_2529,N_22414,N_23933);
or UO_2530 (O_2530,N_23308,N_22684);
or UO_2531 (O_2531,N_24893,N_22061);
nor UO_2532 (O_2532,N_23580,N_23043);
nor UO_2533 (O_2533,N_23468,N_22356);
nor UO_2534 (O_2534,N_22651,N_22135);
or UO_2535 (O_2535,N_24711,N_24673);
and UO_2536 (O_2536,N_22635,N_23635);
and UO_2537 (O_2537,N_23734,N_23957);
nor UO_2538 (O_2538,N_24171,N_24637);
nor UO_2539 (O_2539,N_24057,N_22785);
xnor UO_2540 (O_2540,N_24470,N_22022);
nor UO_2541 (O_2541,N_22958,N_22050);
nand UO_2542 (O_2542,N_23123,N_22284);
xnor UO_2543 (O_2543,N_23137,N_24329);
xor UO_2544 (O_2544,N_24688,N_24644);
xnor UO_2545 (O_2545,N_24796,N_24351);
and UO_2546 (O_2546,N_24487,N_23519);
nand UO_2547 (O_2547,N_22630,N_22712);
or UO_2548 (O_2548,N_23097,N_22143);
and UO_2549 (O_2549,N_24605,N_23687);
nor UO_2550 (O_2550,N_22186,N_22206);
xnor UO_2551 (O_2551,N_24741,N_24767);
nor UO_2552 (O_2552,N_24378,N_22482);
nor UO_2553 (O_2553,N_22969,N_22789);
nor UO_2554 (O_2554,N_22595,N_24497);
nand UO_2555 (O_2555,N_22911,N_23627);
nor UO_2556 (O_2556,N_23982,N_24795);
xor UO_2557 (O_2557,N_22079,N_24278);
xor UO_2558 (O_2558,N_24267,N_22995);
and UO_2559 (O_2559,N_22958,N_23303);
xnor UO_2560 (O_2560,N_24628,N_22327);
nor UO_2561 (O_2561,N_22479,N_24658);
nand UO_2562 (O_2562,N_22882,N_24137);
or UO_2563 (O_2563,N_21900,N_23862);
or UO_2564 (O_2564,N_24037,N_22254);
xnor UO_2565 (O_2565,N_24590,N_23729);
or UO_2566 (O_2566,N_22561,N_24555);
and UO_2567 (O_2567,N_23786,N_24037);
nand UO_2568 (O_2568,N_23039,N_23714);
or UO_2569 (O_2569,N_24598,N_24510);
xor UO_2570 (O_2570,N_22735,N_23231);
nand UO_2571 (O_2571,N_23781,N_23723);
nor UO_2572 (O_2572,N_22212,N_24447);
xor UO_2573 (O_2573,N_23124,N_24338);
nor UO_2574 (O_2574,N_23181,N_23681);
xnor UO_2575 (O_2575,N_23457,N_23503);
xor UO_2576 (O_2576,N_23182,N_22762);
xor UO_2577 (O_2577,N_23364,N_23767);
and UO_2578 (O_2578,N_24952,N_23534);
nor UO_2579 (O_2579,N_23438,N_23174);
xor UO_2580 (O_2580,N_23604,N_24055);
nor UO_2581 (O_2581,N_24685,N_24308);
and UO_2582 (O_2582,N_22315,N_24597);
xor UO_2583 (O_2583,N_24748,N_24605);
and UO_2584 (O_2584,N_23426,N_22252);
or UO_2585 (O_2585,N_24783,N_22100);
or UO_2586 (O_2586,N_21908,N_23906);
or UO_2587 (O_2587,N_24431,N_23324);
or UO_2588 (O_2588,N_23497,N_24056);
xor UO_2589 (O_2589,N_22602,N_24978);
nor UO_2590 (O_2590,N_22221,N_22334);
or UO_2591 (O_2591,N_23637,N_24830);
nand UO_2592 (O_2592,N_22934,N_23321);
or UO_2593 (O_2593,N_24863,N_22398);
and UO_2594 (O_2594,N_23434,N_23539);
or UO_2595 (O_2595,N_22815,N_23504);
xnor UO_2596 (O_2596,N_22487,N_23657);
nor UO_2597 (O_2597,N_24308,N_23300);
xor UO_2598 (O_2598,N_21883,N_24362);
xor UO_2599 (O_2599,N_24427,N_23085);
nor UO_2600 (O_2600,N_23358,N_22446);
nand UO_2601 (O_2601,N_24002,N_22684);
nor UO_2602 (O_2602,N_24951,N_24476);
and UO_2603 (O_2603,N_23769,N_22050);
nand UO_2604 (O_2604,N_24613,N_22436);
and UO_2605 (O_2605,N_22099,N_24108);
xor UO_2606 (O_2606,N_24439,N_23794);
nor UO_2607 (O_2607,N_22879,N_23019);
and UO_2608 (O_2608,N_23787,N_24836);
nand UO_2609 (O_2609,N_23945,N_22508);
or UO_2610 (O_2610,N_24251,N_24140);
xor UO_2611 (O_2611,N_22250,N_24924);
xnor UO_2612 (O_2612,N_23467,N_22365);
xor UO_2613 (O_2613,N_24162,N_24065);
or UO_2614 (O_2614,N_24882,N_23336);
nand UO_2615 (O_2615,N_24166,N_22395);
or UO_2616 (O_2616,N_23634,N_22877);
xnor UO_2617 (O_2617,N_21893,N_23477);
nand UO_2618 (O_2618,N_23452,N_22974);
xor UO_2619 (O_2619,N_24220,N_22535);
xor UO_2620 (O_2620,N_22922,N_23422);
xnor UO_2621 (O_2621,N_24128,N_22213);
xor UO_2622 (O_2622,N_23764,N_24811);
or UO_2623 (O_2623,N_23128,N_23222);
and UO_2624 (O_2624,N_23918,N_22669);
nand UO_2625 (O_2625,N_24395,N_24630);
nor UO_2626 (O_2626,N_22717,N_24884);
or UO_2627 (O_2627,N_23950,N_23594);
nor UO_2628 (O_2628,N_23930,N_23464);
xor UO_2629 (O_2629,N_23648,N_23668);
nor UO_2630 (O_2630,N_24803,N_23771);
or UO_2631 (O_2631,N_24991,N_23257);
and UO_2632 (O_2632,N_24576,N_22255);
and UO_2633 (O_2633,N_23409,N_22841);
nand UO_2634 (O_2634,N_22877,N_22197);
nor UO_2635 (O_2635,N_24288,N_23953);
nand UO_2636 (O_2636,N_23196,N_24281);
nor UO_2637 (O_2637,N_22644,N_23588);
and UO_2638 (O_2638,N_23987,N_23767);
or UO_2639 (O_2639,N_22354,N_22827);
nor UO_2640 (O_2640,N_23323,N_23923);
nor UO_2641 (O_2641,N_22448,N_22436);
nor UO_2642 (O_2642,N_23446,N_24294);
nand UO_2643 (O_2643,N_23930,N_22124);
or UO_2644 (O_2644,N_21909,N_24858);
nor UO_2645 (O_2645,N_24054,N_24391);
nor UO_2646 (O_2646,N_24897,N_23279);
xnor UO_2647 (O_2647,N_22133,N_24038);
and UO_2648 (O_2648,N_24927,N_24756);
xnor UO_2649 (O_2649,N_23493,N_22104);
xor UO_2650 (O_2650,N_23035,N_23132);
xnor UO_2651 (O_2651,N_22638,N_23179);
nor UO_2652 (O_2652,N_24914,N_23448);
or UO_2653 (O_2653,N_22412,N_23734);
xnor UO_2654 (O_2654,N_22202,N_24892);
and UO_2655 (O_2655,N_24302,N_22401);
or UO_2656 (O_2656,N_21893,N_24907);
nor UO_2657 (O_2657,N_24109,N_24398);
and UO_2658 (O_2658,N_23779,N_23231);
nor UO_2659 (O_2659,N_24047,N_22378);
and UO_2660 (O_2660,N_22875,N_23267);
xor UO_2661 (O_2661,N_22687,N_22213);
xor UO_2662 (O_2662,N_22678,N_23761);
xor UO_2663 (O_2663,N_23890,N_23524);
nor UO_2664 (O_2664,N_22782,N_22937);
or UO_2665 (O_2665,N_24259,N_24015);
nand UO_2666 (O_2666,N_22367,N_21932);
nand UO_2667 (O_2667,N_22102,N_22692);
nand UO_2668 (O_2668,N_24277,N_23531);
xor UO_2669 (O_2669,N_21920,N_22645);
and UO_2670 (O_2670,N_22559,N_23228);
nand UO_2671 (O_2671,N_24489,N_23557);
nor UO_2672 (O_2672,N_22328,N_24409);
nand UO_2673 (O_2673,N_22019,N_24960);
or UO_2674 (O_2674,N_24899,N_22626);
or UO_2675 (O_2675,N_21929,N_22359);
xnor UO_2676 (O_2676,N_21962,N_23327);
nand UO_2677 (O_2677,N_24122,N_23322);
or UO_2678 (O_2678,N_24647,N_23060);
nor UO_2679 (O_2679,N_23446,N_21981);
nand UO_2680 (O_2680,N_22080,N_23519);
nor UO_2681 (O_2681,N_23998,N_24592);
xnor UO_2682 (O_2682,N_22724,N_21988);
xor UO_2683 (O_2683,N_22786,N_22865);
xor UO_2684 (O_2684,N_23802,N_23175);
nor UO_2685 (O_2685,N_24783,N_24653);
or UO_2686 (O_2686,N_22363,N_24644);
or UO_2687 (O_2687,N_23245,N_23666);
nor UO_2688 (O_2688,N_24051,N_22075);
nor UO_2689 (O_2689,N_23947,N_24464);
nand UO_2690 (O_2690,N_23792,N_24111);
or UO_2691 (O_2691,N_24949,N_23922);
and UO_2692 (O_2692,N_24798,N_24914);
or UO_2693 (O_2693,N_22678,N_24442);
nor UO_2694 (O_2694,N_22034,N_24195);
and UO_2695 (O_2695,N_24053,N_24022);
and UO_2696 (O_2696,N_22262,N_23831);
and UO_2697 (O_2697,N_22910,N_21931);
nand UO_2698 (O_2698,N_22626,N_22181);
nand UO_2699 (O_2699,N_23501,N_22073);
nor UO_2700 (O_2700,N_22211,N_22070);
or UO_2701 (O_2701,N_23252,N_24685);
and UO_2702 (O_2702,N_22122,N_23159);
nand UO_2703 (O_2703,N_23326,N_24998);
xnor UO_2704 (O_2704,N_23005,N_22232);
xor UO_2705 (O_2705,N_22058,N_23455);
nor UO_2706 (O_2706,N_24891,N_23604);
nand UO_2707 (O_2707,N_23713,N_22991);
nand UO_2708 (O_2708,N_24061,N_22640);
xor UO_2709 (O_2709,N_24307,N_24847);
xor UO_2710 (O_2710,N_24895,N_24046);
or UO_2711 (O_2711,N_22150,N_21999);
xnor UO_2712 (O_2712,N_23464,N_23196);
nand UO_2713 (O_2713,N_22924,N_24744);
and UO_2714 (O_2714,N_22180,N_23090);
nand UO_2715 (O_2715,N_24672,N_23643);
or UO_2716 (O_2716,N_23441,N_24439);
or UO_2717 (O_2717,N_24414,N_23271);
nor UO_2718 (O_2718,N_23905,N_24662);
nand UO_2719 (O_2719,N_24137,N_22105);
nor UO_2720 (O_2720,N_23898,N_24898);
and UO_2721 (O_2721,N_22367,N_23619);
nand UO_2722 (O_2722,N_24263,N_24175);
nor UO_2723 (O_2723,N_23772,N_24313);
and UO_2724 (O_2724,N_24093,N_22901);
nor UO_2725 (O_2725,N_23254,N_23634);
and UO_2726 (O_2726,N_23575,N_22208);
nor UO_2727 (O_2727,N_24197,N_24291);
nand UO_2728 (O_2728,N_23519,N_23569);
and UO_2729 (O_2729,N_21882,N_24053);
nand UO_2730 (O_2730,N_23194,N_22836);
nand UO_2731 (O_2731,N_22530,N_22102);
and UO_2732 (O_2732,N_22784,N_22398);
nor UO_2733 (O_2733,N_23255,N_22718);
nor UO_2734 (O_2734,N_22749,N_24978);
and UO_2735 (O_2735,N_23946,N_22547);
nand UO_2736 (O_2736,N_23977,N_22160);
xor UO_2737 (O_2737,N_22759,N_24163);
nand UO_2738 (O_2738,N_24002,N_22510);
and UO_2739 (O_2739,N_22141,N_23040);
and UO_2740 (O_2740,N_24521,N_22553);
nand UO_2741 (O_2741,N_24112,N_22254);
or UO_2742 (O_2742,N_22917,N_24979);
or UO_2743 (O_2743,N_24809,N_22738);
nor UO_2744 (O_2744,N_24888,N_22551);
and UO_2745 (O_2745,N_24389,N_22256);
xnor UO_2746 (O_2746,N_22547,N_23326);
and UO_2747 (O_2747,N_24955,N_23111);
nor UO_2748 (O_2748,N_24877,N_24250);
nand UO_2749 (O_2749,N_23461,N_23388);
nand UO_2750 (O_2750,N_24081,N_24178);
nor UO_2751 (O_2751,N_24170,N_24341);
nor UO_2752 (O_2752,N_23051,N_22476);
xnor UO_2753 (O_2753,N_23004,N_21931);
nand UO_2754 (O_2754,N_22468,N_23190);
or UO_2755 (O_2755,N_22443,N_24605);
or UO_2756 (O_2756,N_22305,N_22164);
and UO_2757 (O_2757,N_23220,N_22775);
nand UO_2758 (O_2758,N_22740,N_22236);
nor UO_2759 (O_2759,N_24294,N_24331);
and UO_2760 (O_2760,N_23462,N_24049);
xnor UO_2761 (O_2761,N_23167,N_23698);
xor UO_2762 (O_2762,N_22331,N_24103);
nand UO_2763 (O_2763,N_24959,N_22335);
or UO_2764 (O_2764,N_24624,N_23811);
or UO_2765 (O_2765,N_24407,N_23602);
or UO_2766 (O_2766,N_22772,N_22723);
xnor UO_2767 (O_2767,N_22706,N_24233);
nor UO_2768 (O_2768,N_22536,N_23487);
nand UO_2769 (O_2769,N_24135,N_22588);
and UO_2770 (O_2770,N_23179,N_22677);
or UO_2771 (O_2771,N_23598,N_22025);
nand UO_2772 (O_2772,N_24283,N_23924);
and UO_2773 (O_2773,N_22762,N_24102);
nand UO_2774 (O_2774,N_24655,N_23087);
and UO_2775 (O_2775,N_24238,N_23217);
nor UO_2776 (O_2776,N_23140,N_23260);
nor UO_2777 (O_2777,N_23477,N_24247);
nor UO_2778 (O_2778,N_21927,N_22064);
nor UO_2779 (O_2779,N_22879,N_24720);
nor UO_2780 (O_2780,N_24866,N_22154);
xnor UO_2781 (O_2781,N_22173,N_21955);
nand UO_2782 (O_2782,N_22878,N_22449);
and UO_2783 (O_2783,N_23051,N_23744);
and UO_2784 (O_2784,N_23631,N_23687);
or UO_2785 (O_2785,N_23500,N_22474);
and UO_2786 (O_2786,N_22040,N_24863);
xnor UO_2787 (O_2787,N_24098,N_23974);
nand UO_2788 (O_2788,N_24444,N_24602);
xor UO_2789 (O_2789,N_22358,N_23279);
nor UO_2790 (O_2790,N_23651,N_22506);
nand UO_2791 (O_2791,N_22825,N_23738);
nand UO_2792 (O_2792,N_22909,N_22657);
and UO_2793 (O_2793,N_23794,N_24152);
and UO_2794 (O_2794,N_24313,N_22208);
and UO_2795 (O_2795,N_24628,N_23701);
nand UO_2796 (O_2796,N_23300,N_22399);
nand UO_2797 (O_2797,N_23361,N_24190);
nand UO_2798 (O_2798,N_22238,N_22493);
nor UO_2799 (O_2799,N_22216,N_24807);
nand UO_2800 (O_2800,N_22313,N_24860);
nand UO_2801 (O_2801,N_24653,N_21904);
or UO_2802 (O_2802,N_22989,N_23306);
and UO_2803 (O_2803,N_23470,N_22910);
nand UO_2804 (O_2804,N_23366,N_23309);
nand UO_2805 (O_2805,N_23474,N_23852);
and UO_2806 (O_2806,N_23372,N_23463);
and UO_2807 (O_2807,N_22142,N_24871);
nand UO_2808 (O_2808,N_22433,N_24270);
nand UO_2809 (O_2809,N_22022,N_22517);
or UO_2810 (O_2810,N_23397,N_22172);
and UO_2811 (O_2811,N_22658,N_23780);
and UO_2812 (O_2812,N_24150,N_22360);
nor UO_2813 (O_2813,N_23031,N_23760);
nand UO_2814 (O_2814,N_24336,N_23092);
and UO_2815 (O_2815,N_22410,N_22739);
and UO_2816 (O_2816,N_22643,N_22268);
and UO_2817 (O_2817,N_24563,N_24874);
nor UO_2818 (O_2818,N_22445,N_23174);
or UO_2819 (O_2819,N_22979,N_22187);
nand UO_2820 (O_2820,N_22356,N_22867);
or UO_2821 (O_2821,N_22351,N_23123);
or UO_2822 (O_2822,N_24637,N_24362);
or UO_2823 (O_2823,N_23229,N_24179);
xnor UO_2824 (O_2824,N_23680,N_22903);
nor UO_2825 (O_2825,N_22426,N_23338);
or UO_2826 (O_2826,N_23356,N_23381);
nor UO_2827 (O_2827,N_24937,N_22783);
nand UO_2828 (O_2828,N_22764,N_23278);
or UO_2829 (O_2829,N_23619,N_23051);
nor UO_2830 (O_2830,N_24306,N_23649);
and UO_2831 (O_2831,N_21963,N_23367);
xnor UO_2832 (O_2832,N_24044,N_24908);
or UO_2833 (O_2833,N_23113,N_22392);
nor UO_2834 (O_2834,N_22559,N_24209);
nand UO_2835 (O_2835,N_23668,N_23808);
or UO_2836 (O_2836,N_22297,N_21989);
or UO_2837 (O_2837,N_22116,N_24086);
xor UO_2838 (O_2838,N_23719,N_22802);
xor UO_2839 (O_2839,N_23708,N_23980);
xnor UO_2840 (O_2840,N_23028,N_22101);
nand UO_2841 (O_2841,N_24224,N_23573);
nor UO_2842 (O_2842,N_23171,N_24531);
and UO_2843 (O_2843,N_22061,N_23832);
and UO_2844 (O_2844,N_22568,N_22248);
nor UO_2845 (O_2845,N_22690,N_23474);
nor UO_2846 (O_2846,N_22080,N_22331);
nor UO_2847 (O_2847,N_24730,N_21964);
and UO_2848 (O_2848,N_24426,N_23920);
and UO_2849 (O_2849,N_24290,N_24964);
or UO_2850 (O_2850,N_22036,N_23542);
xor UO_2851 (O_2851,N_22814,N_22341);
nand UO_2852 (O_2852,N_24276,N_22352);
and UO_2853 (O_2853,N_24772,N_24684);
nand UO_2854 (O_2854,N_24607,N_22479);
and UO_2855 (O_2855,N_23147,N_22840);
xnor UO_2856 (O_2856,N_22832,N_22662);
or UO_2857 (O_2857,N_23087,N_23620);
nor UO_2858 (O_2858,N_23696,N_23042);
nor UO_2859 (O_2859,N_21933,N_23808);
or UO_2860 (O_2860,N_24442,N_24589);
or UO_2861 (O_2861,N_24400,N_22232);
and UO_2862 (O_2862,N_22017,N_24247);
nor UO_2863 (O_2863,N_22982,N_24335);
and UO_2864 (O_2864,N_24228,N_22244);
or UO_2865 (O_2865,N_23853,N_22475);
nor UO_2866 (O_2866,N_22699,N_23796);
and UO_2867 (O_2867,N_24880,N_23842);
or UO_2868 (O_2868,N_23606,N_22991);
and UO_2869 (O_2869,N_24336,N_22410);
nor UO_2870 (O_2870,N_24991,N_22636);
and UO_2871 (O_2871,N_24104,N_24321);
xnor UO_2872 (O_2872,N_24198,N_22481);
and UO_2873 (O_2873,N_24901,N_23836);
and UO_2874 (O_2874,N_24228,N_22499);
nor UO_2875 (O_2875,N_22174,N_23549);
and UO_2876 (O_2876,N_23546,N_22482);
xnor UO_2877 (O_2877,N_23750,N_24425);
xnor UO_2878 (O_2878,N_22212,N_21977);
nor UO_2879 (O_2879,N_22723,N_23988);
xnor UO_2880 (O_2880,N_24961,N_22917);
or UO_2881 (O_2881,N_24860,N_23352);
and UO_2882 (O_2882,N_22433,N_23108);
or UO_2883 (O_2883,N_22871,N_24131);
and UO_2884 (O_2884,N_22525,N_23262);
xor UO_2885 (O_2885,N_24201,N_22313);
nor UO_2886 (O_2886,N_24537,N_23153);
or UO_2887 (O_2887,N_22663,N_23905);
or UO_2888 (O_2888,N_23110,N_24138);
or UO_2889 (O_2889,N_24767,N_24212);
and UO_2890 (O_2890,N_22025,N_24935);
nand UO_2891 (O_2891,N_24938,N_22999);
and UO_2892 (O_2892,N_24654,N_22738);
or UO_2893 (O_2893,N_23986,N_22781);
xor UO_2894 (O_2894,N_24829,N_24299);
or UO_2895 (O_2895,N_23371,N_24652);
nand UO_2896 (O_2896,N_23063,N_24748);
xnor UO_2897 (O_2897,N_22514,N_22073);
nor UO_2898 (O_2898,N_23464,N_22870);
nor UO_2899 (O_2899,N_23534,N_23780);
xor UO_2900 (O_2900,N_21975,N_22268);
xor UO_2901 (O_2901,N_23729,N_22476);
or UO_2902 (O_2902,N_23142,N_24543);
nor UO_2903 (O_2903,N_22444,N_24078);
nor UO_2904 (O_2904,N_22356,N_24699);
nor UO_2905 (O_2905,N_24761,N_21942);
and UO_2906 (O_2906,N_24626,N_23965);
and UO_2907 (O_2907,N_23561,N_23019);
or UO_2908 (O_2908,N_22113,N_23835);
xor UO_2909 (O_2909,N_23847,N_22750);
and UO_2910 (O_2910,N_24437,N_23852);
and UO_2911 (O_2911,N_22026,N_24054);
nor UO_2912 (O_2912,N_23572,N_24441);
xor UO_2913 (O_2913,N_24815,N_22759);
and UO_2914 (O_2914,N_22228,N_22064);
nor UO_2915 (O_2915,N_23890,N_24261);
xor UO_2916 (O_2916,N_23619,N_24586);
nor UO_2917 (O_2917,N_24363,N_21920);
nand UO_2918 (O_2918,N_24549,N_22883);
nand UO_2919 (O_2919,N_24371,N_22863);
nor UO_2920 (O_2920,N_22084,N_24207);
or UO_2921 (O_2921,N_22004,N_23567);
and UO_2922 (O_2922,N_24175,N_24638);
and UO_2923 (O_2923,N_22237,N_22167);
nor UO_2924 (O_2924,N_23601,N_23173);
xnor UO_2925 (O_2925,N_24738,N_22614);
xnor UO_2926 (O_2926,N_22871,N_24274);
and UO_2927 (O_2927,N_23538,N_24588);
nor UO_2928 (O_2928,N_23004,N_24410);
xor UO_2929 (O_2929,N_23277,N_24197);
nand UO_2930 (O_2930,N_23811,N_22399);
nand UO_2931 (O_2931,N_23761,N_22966);
nand UO_2932 (O_2932,N_24342,N_22762);
nor UO_2933 (O_2933,N_22953,N_23549);
nand UO_2934 (O_2934,N_24548,N_23785);
or UO_2935 (O_2935,N_24791,N_22510);
or UO_2936 (O_2936,N_22235,N_22578);
xor UO_2937 (O_2937,N_24187,N_24233);
or UO_2938 (O_2938,N_24442,N_23445);
and UO_2939 (O_2939,N_22348,N_24242);
xnor UO_2940 (O_2940,N_22646,N_24485);
and UO_2941 (O_2941,N_22076,N_24580);
nand UO_2942 (O_2942,N_24081,N_23460);
nor UO_2943 (O_2943,N_23041,N_21996);
xnor UO_2944 (O_2944,N_22560,N_22321);
nand UO_2945 (O_2945,N_24628,N_24678);
xnor UO_2946 (O_2946,N_24818,N_23283);
or UO_2947 (O_2947,N_22905,N_22553);
and UO_2948 (O_2948,N_24587,N_22571);
or UO_2949 (O_2949,N_21990,N_22186);
and UO_2950 (O_2950,N_22630,N_23518);
nand UO_2951 (O_2951,N_23841,N_24470);
or UO_2952 (O_2952,N_22137,N_22081);
or UO_2953 (O_2953,N_24262,N_24476);
and UO_2954 (O_2954,N_24835,N_22992);
nand UO_2955 (O_2955,N_24567,N_24578);
nand UO_2956 (O_2956,N_23012,N_22858);
nor UO_2957 (O_2957,N_22392,N_24921);
nor UO_2958 (O_2958,N_23491,N_24843);
and UO_2959 (O_2959,N_22710,N_23909);
xnor UO_2960 (O_2960,N_24308,N_24276);
or UO_2961 (O_2961,N_23246,N_22676);
nor UO_2962 (O_2962,N_24401,N_22433);
xnor UO_2963 (O_2963,N_23075,N_23815);
and UO_2964 (O_2964,N_22210,N_23267);
xor UO_2965 (O_2965,N_23115,N_22101);
nand UO_2966 (O_2966,N_24895,N_22097);
or UO_2967 (O_2967,N_22098,N_23570);
nand UO_2968 (O_2968,N_23608,N_24639);
and UO_2969 (O_2969,N_23878,N_22789);
and UO_2970 (O_2970,N_22788,N_24827);
nand UO_2971 (O_2971,N_22307,N_24797);
and UO_2972 (O_2972,N_24616,N_23721);
nand UO_2973 (O_2973,N_23733,N_23012);
nor UO_2974 (O_2974,N_24092,N_22328);
nand UO_2975 (O_2975,N_24510,N_22410);
nand UO_2976 (O_2976,N_23282,N_23334);
and UO_2977 (O_2977,N_23563,N_22149);
xor UO_2978 (O_2978,N_24182,N_24822);
nor UO_2979 (O_2979,N_24592,N_22880);
nand UO_2980 (O_2980,N_24816,N_23990);
xnor UO_2981 (O_2981,N_23050,N_24436);
nor UO_2982 (O_2982,N_23180,N_23193);
xor UO_2983 (O_2983,N_23817,N_23152);
nand UO_2984 (O_2984,N_24184,N_24216);
nor UO_2985 (O_2985,N_22343,N_24842);
nor UO_2986 (O_2986,N_24874,N_23663);
nand UO_2987 (O_2987,N_23585,N_23744);
nand UO_2988 (O_2988,N_23022,N_23670);
nand UO_2989 (O_2989,N_24804,N_22836);
and UO_2990 (O_2990,N_22636,N_24816);
nand UO_2991 (O_2991,N_22687,N_24820);
nand UO_2992 (O_2992,N_24311,N_22438);
and UO_2993 (O_2993,N_22984,N_22098);
xnor UO_2994 (O_2994,N_23860,N_22229);
xnor UO_2995 (O_2995,N_24626,N_24479);
xor UO_2996 (O_2996,N_22702,N_21972);
and UO_2997 (O_2997,N_24050,N_24940);
nor UO_2998 (O_2998,N_23790,N_24255);
xnor UO_2999 (O_2999,N_23274,N_22798);
endmodule