module basic_500_3000_500_4_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_209,In_15);
and U1 (N_1,In_422,In_49);
nor U2 (N_2,In_172,In_173);
nor U3 (N_3,In_52,In_461);
nor U4 (N_4,In_152,In_392);
xnor U5 (N_5,In_463,In_363);
and U6 (N_6,In_319,In_382);
nor U7 (N_7,In_322,In_101);
nand U8 (N_8,In_34,In_132);
xor U9 (N_9,In_161,In_185);
nand U10 (N_10,In_198,In_378);
nand U11 (N_11,In_199,In_139);
nor U12 (N_12,In_43,In_408);
nor U13 (N_13,In_64,In_343);
and U14 (N_14,In_246,In_241);
nand U15 (N_15,In_379,In_292);
or U16 (N_16,In_487,In_76);
nor U17 (N_17,In_341,In_149);
nor U18 (N_18,In_486,In_11);
and U19 (N_19,In_81,In_360);
nor U20 (N_20,In_270,In_208);
or U21 (N_21,In_446,In_3);
and U22 (N_22,In_476,In_53);
or U23 (N_23,In_239,In_140);
nor U24 (N_24,In_311,In_125);
or U25 (N_25,In_218,In_248);
nor U26 (N_26,In_485,In_36);
nand U27 (N_27,In_260,In_89);
and U28 (N_28,In_389,In_69);
xor U29 (N_29,In_250,In_370);
and U30 (N_30,In_308,In_60);
nor U31 (N_31,In_236,In_37);
nor U32 (N_32,In_57,In_414);
nor U33 (N_33,In_336,In_74);
xnor U34 (N_34,In_405,In_478);
or U35 (N_35,In_168,In_334);
nand U36 (N_36,In_399,In_26);
and U37 (N_37,In_268,In_313);
nor U38 (N_38,In_397,In_95);
or U39 (N_39,In_471,In_421);
or U40 (N_40,In_212,In_238);
and U41 (N_41,In_456,In_479);
nand U42 (N_42,In_99,In_348);
and U43 (N_43,In_20,In_96);
nand U44 (N_44,In_327,In_70);
nand U45 (N_45,In_430,In_449);
xor U46 (N_46,In_32,In_438);
and U47 (N_47,In_123,In_155);
nand U48 (N_48,In_483,In_41);
and U49 (N_49,In_184,In_50);
or U50 (N_50,In_420,In_51);
or U51 (N_51,In_317,In_42);
and U52 (N_52,In_63,In_273);
xnor U53 (N_53,In_200,In_91);
nand U54 (N_54,In_44,In_359);
and U55 (N_55,In_277,In_169);
or U56 (N_56,In_281,In_332);
nor U57 (N_57,In_264,In_75);
nand U58 (N_58,In_371,In_349);
nand U59 (N_59,In_289,In_230);
and U60 (N_60,In_47,In_165);
and U61 (N_61,In_119,In_297);
nand U62 (N_62,In_423,In_80);
or U63 (N_63,In_345,In_90);
and U64 (N_64,In_367,In_195);
or U65 (N_65,In_354,In_416);
nor U66 (N_66,In_104,In_434);
nand U67 (N_67,In_303,In_194);
nand U68 (N_68,In_204,In_127);
xnor U69 (N_69,In_78,In_72);
nand U70 (N_70,In_192,In_495);
nor U71 (N_71,In_451,In_13);
nand U72 (N_72,In_112,In_162);
nand U73 (N_73,In_84,In_150);
xnor U74 (N_74,In_35,In_58);
nand U75 (N_75,In_376,In_138);
nor U76 (N_76,In_267,In_439);
nor U77 (N_77,In_288,In_33);
and U78 (N_78,In_103,In_386);
nor U79 (N_79,In_462,In_419);
nor U80 (N_80,In_175,In_144);
nor U81 (N_81,In_488,In_489);
nand U82 (N_82,In_337,In_22);
or U83 (N_83,In_201,In_255);
nand U84 (N_84,In_153,In_46);
or U85 (N_85,In_251,In_458);
nor U86 (N_86,In_79,In_178);
xor U87 (N_87,In_290,In_100);
or U88 (N_88,In_117,In_65);
nor U89 (N_89,In_98,In_235);
or U90 (N_90,In_432,In_299);
or U91 (N_91,In_364,In_325);
nor U92 (N_92,In_443,In_448);
and U93 (N_93,In_480,In_259);
nand U94 (N_94,In_221,In_324);
xnor U95 (N_95,In_4,In_492);
xor U96 (N_96,In_445,In_122);
or U97 (N_97,In_205,In_7);
nand U98 (N_98,In_460,In_442);
xnor U99 (N_99,In_14,In_30);
nand U100 (N_100,In_331,In_272);
nor U101 (N_101,In_197,In_309);
or U102 (N_102,In_186,In_436);
and U103 (N_103,In_231,In_494);
nand U104 (N_104,In_312,In_431);
nor U105 (N_105,In_293,In_223);
and U106 (N_106,In_130,In_244);
xor U107 (N_107,In_181,In_473);
and U108 (N_108,In_249,In_437);
nand U109 (N_109,In_291,In_224);
and U110 (N_110,In_187,In_394);
nor U111 (N_111,In_202,In_409);
and U112 (N_112,In_284,In_48);
nor U113 (N_113,In_428,In_373);
or U114 (N_114,In_131,In_377);
nand U115 (N_115,In_111,In_450);
or U116 (N_116,In_306,In_86);
or U117 (N_117,In_316,In_315);
nand U118 (N_118,In_128,In_83);
nor U119 (N_119,In_31,In_177);
or U120 (N_120,In_118,In_280);
nand U121 (N_121,In_94,In_18);
and U122 (N_122,In_163,In_158);
and U123 (N_123,In_116,In_245);
or U124 (N_124,In_134,In_302);
and U125 (N_125,In_258,In_365);
nor U126 (N_126,In_114,In_242);
xnor U127 (N_127,In_38,In_253);
or U128 (N_128,In_469,In_464);
nor U129 (N_129,In_427,In_351);
xnor U130 (N_130,In_368,In_411);
nor U131 (N_131,In_429,In_228);
or U132 (N_132,In_180,In_148);
xor U133 (N_133,In_383,In_93);
and U134 (N_134,In_453,In_137);
and U135 (N_135,In_55,In_404);
and U136 (N_136,In_124,In_358);
nor U137 (N_137,In_179,In_109);
nand U138 (N_138,In_157,In_225);
or U139 (N_139,In_490,In_240);
or U140 (N_140,In_452,In_335);
nor U141 (N_141,In_474,In_301);
xor U142 (N_142,In_286,In_222);
nor U143 (N_143,In_207,In_323);
and U144 (N_144,In_418,In_285);
nor U145 (N_145,In_384,In_88);
or U146 (N_146,In_328,In_66);
nor U147 (N_147,In_484,In_415);
or U148 (N_148,In_355,In_441);
nor U149 (N_149,In_82,In_107);
or U150 (N_150,In_497,In_435);
and U151 (N_151,In_45,In_220);
nor U152 (N_152,In_388,In_143);
nor U153 (N_153,In_5,In_499);
nor U154 (N_154,In_444,In_135);
nor U155 (N_155,In_307,In_191);
nor U156 (N_156,In_387,In_196);
and U157 (N_157,In_10,In_347);
and U158 (N_158,In_25,In_237);
nor U159 (N_159,In_403,In_183);
or U160 (N_160,In_40,In_390);
and U161 (N_161,In_396,In_385);
or U162 (N_162,In_320,In_372);
nand U163 (N_163,In_330,In_424);
nand U164 (N_164,In_275,In_375);
nand U165 (N_165,In_344,In_468);
nor U166 (N_166,In_190,In_481);
nor U167 (N_167,In_188,In_8);
nand U168 (N_168,In_263,In_407);
and U169 (N_169,In_401,In_97);
or U170 (N_170,In_357,In_85);
nor U171 (N_171,In_12,In_59);
xnor U172 (N_172,In_219,In_276);
nand U173 (N_173,In_433,In_466);
and U174 (N_174,In_229,In_23);
and U175 (N_175,In_174,In_269);
or U176 (N_176,In_211,In_110);
nor U177 (N_177,In_266,In_457);
or U178 (N_178,In_472,In_213);
and U179 (N_179,In_170,In_247);
and U180 (N_180,In_234,In_321);
nand U181 (N_181,In_356,In_374);
xor U182 (N_182,In_77,In_0);
nor U183 (N_183,In_115,In_120);
nor U184 (N_184,In_206,In_164);
nand U185 (N_185,In_381,In_151);
xnor U186 (N_186,In_28,In_252);
or U187 (N_187,In_304,In_6);
or U188 (N_188,In_27,In_283);
nor U189 (N_189,In_278,In_193);
and U190 (N_190,In_413,In_274);
nor U191 (N_191,In_146,In_166);
or U192 (N_192,In_257,In_340);
nand U193 (N_193,In_68,In_243);
or U194 (N_194,In_366,In_393);
nor U195 (N_195,In_24,In_102);
or U196 (N_196,In_296,In_133);
nor U197 (N_197,In_454,In_333);
nand U198 (N_198,In_369,In_310);
nor U199 (N_199,In_136,In_400);
or U200 (N_200,In_71,In_261);
nand U201 (N_201,In_217,In_156);
nand U202 (N_202,In_493,In_346);
and U203 (N_203,In_145,In_106);
or U204 (N_204,In_159,In_17);
or U205 (N_205,In_477,In_459);
nor U206 (N_206,In_147,In_210);
and U207 (N_207,In_214,In_314);
and U208 (N_208,In_121,In_326);
or U209 (N_209,In_342,In_167);
nor U210 (N_210,In_440,In_226);
xor U211 (N_211,In_318,In_1);
or U212 (N_212,In_279,In_227);
or U213 (N_213,In_380,In_67);
nand U214 (N_214,In_294,In_447);
xnor U215 (N_215,In_29,In_298);
xor U216 (N_216,In_295,In_129);
nand U217 (N_217,In_154,In_412);
or U218 (N_218,In_498,In_87);
nor U219 (N_219,In_491,In_426);
nor U220 (N_220,In_105,In_391);
nand U221 (N_221,In_467,In_287);
and U222 (N_222,In_352,In_425);
or U223 (N_223,In_54,In_455);
xnor U224 (N_224,In_282,In_475);
and U225 (N_225,In_402,In_338);
and U226 (N_226,In_271,In_176);
and U227 (N_227,In_262,In_203);
or U228 (N_228,In_410,In_216);
nand U229 (N_229,In_108,In_350);
and U230 (N_230,In_92,In_256);
nand U231 (N_231,In_39,In_61);
nand U232 (N_232,In_2,In_182);
nand U233 (N_233,In_215,In_171);
and U234 (N_234,In_329,In_482);
nand U235 (N_235,In_265,In_62);
nand U236 (N_236,In_160,In_395);
nand U237 (N_237,In_470,In_465);
nand U238 (N_238,In_19,In_232);
nand U239 (N_239,In_361,In_141);
nand U240 (N_240,In_73,In_56);
or U241 (N_241,In_353,In_496);
nand U242 (N_242,In_9,In_233);
nand U243 (N_243,In_339,In_113);
nand U244 (N_244,In_417,In_406);
xor U245 (N_245,In_21,In_305);
or U246 (N_246,In_16,In_362);
and U247 (N_247,In_254,In_189);
nor U248 (N_248,In_142,In_398);
or U249 (N_249,In_126,In_300);
or U250 (N_250,In_133,In_370);
and U251 (N_251,In_439,In_477);
and U252 (N_252,In_369,In_496);
or U253 (N_253,In_400,In_397);
and U254 (N_254,In_460,In_261);
nor U255 (N_255,In_191,In_417);
nand U256 (N_256,In_386,In_367);
nand U257 (N_257,In_100,In_451);
or U258 (N_258,In_23,In_436);
or U259 (N_259,In_205,In_489);
nand U260 (N_260,In_488,In_372);
nor U261 (N_261,In_174,In_5);
nor U262 (N_262,In_427,In_118);
nand U263 (N_263,In_291,In_266);
nor U264 (N_264,In_122,In_80);
nand U265 (N_265,In_483,In_99);
nand U266 (N_266,In_381,In_338);
nand U267 (N_267,In_330,In_188);
nor U268 (N_268,In_273,In_285);
nand U269 (N_269,In_271,In_143);
nand U270 (N_270,In_420,In_260);
nor U271 (N_271,In_337,In_73);
nor U272 (N_272,In_72,In_343);
nor U273 (N_273,In_55,In_400);
and U274 (N_274,In_197,In_269);
or U275 (N_275,In_62,In_130);
nor U276 (N_276,In_3,In_284);
nand U277 (N_277,In_295,In_451);
nand U278 (N_278,In_184,In_286);
or U279 (N_279,In_263,In_350);
nand U280 (N_280,In_163,In_396);
and U281 (N_281,In_459,In_82);
xor U282 (N_282,In_369,In_243);
and U283 (N_283,In_258,In_230);
nand U284 (N_284,In_242,In_174);
or U285 (N_285,In_337,In_423);
xnor U286 (N_286,In_253,In_167);
or U287 (N_287,In_245,In_58);
xnor U288 (N_288,In_55,In_281);
nand U289 (N_289,In_60,In_351);
nor U290 (N_290,In_497,In_248);
and U291 (N_291,In_336,In_383);
or U292 (N_292,In_289,In_258);
and U293 (N_293,In_341,In_190);
or U294 (N_294,In_338,In_245);
and U295 (N_295,In_401,In_211);
nor U296 (N_296,In_237,In_198);
nor U297 (N_297,In_470,In_322);
nor U298 (N_298,In_424,In_53);
nand U299 (N_299,In_310,In_215);
nand U300 (N_300,In_453,In_12);
or U301 (N_301,In_418,In_150);
nand U302 (N_302,In_76,In_368);
or U303 (N_303,In_467,In_455);
or U304 (N_304,In_305,In_285);
nand U305 (N_305,In_459,In_284);
nand U306 (N_306,In_220,In_75);
and U307 (N_307,In_122,In_187);
nand U308 (N_308,In_89,In_437);
or U309 (N_309,In_35,In_33);
or U310 (N_310,In_224,In_441);
nor U311 (N_311,In_92,In_374);
and U312 (N_312,In_92,In_186);
nand U313 (N_313,In_2,In_267);
nor U314 (N_314,In_96,In_53);
or U315 (N_315,In_284,In_392);
and U316 (N_316,In_309,In_482);
and U317 (N_317,In_351,In_285);
and U318 (N_318,In_174,In_442);
and U319 (N_319,In_497,In_43);
and U320 (N_320,In_332,In_203);
nand U321 (N_321,In_439,In_142);
or U322 (N_322,In_472,In_228);
or U323 (N_323,In_481,In_361);
or U324 (N_324,In_357,In_360);
and U325 (N_325,In_10,In_284);
or U326 (N_326,In_17,In_115);
nor U327 (N_327,In_376,In_322);
nand U328 (N_328,In_296,In_466);
nor U329 (N_329,In_255,In_261);
or U330 (N_330,In_363,In_190);
nand U331 (N_331,In_134,In_200);
nor U332 (N_332,In_491,In_131);
or U333 (N_333,In_165,In_424);
xnor U334 (N_334,In_165,In_7);
nand U335 (N_335,In_0,In_407);
or U336 (N_336,In_480,In_240);
nand U337 (N_337,In_470,In_223);
nor U338 (N_338,In_260,In_1);
nor U339 (N_339,In_437,In_28);
nand U340 (N_340,In_427,In_131);
nand U341 (N_341,In_399,In_417);
and U342 (N_342,In_196,In_156);
nor U343 (N_343,In_60,In_299);
nor U344 (N_344,In_25,In_272);
nor U345 (N_345,In_312,In_494);
xnor U346 (N_346,In_282,In_113);
or U347 (N_347,In_248,In_32);
nand U348 (N_348,In_247,In_104);
nand U349 (N_349,In_85,In_441);
and U350 (N_350,In_263,In_141);
and U351 (N_351,In_478,In_368);
nand U352 (N_352,In_218,In_40);
nor U353 (N_353,In_424,In_266);
nand U354 (N_354,In_352,In_486);
xnor U355 (N_355,In_38,In_7);
or U356 (N_356,In_148,In_321);
nor U357 (N_357,In_27,In_433);
xnor U358 (N_358,In_349,In_68);
nand U359 (N_359,In_493,In_273);
or U360 (N_360,In_228,In_102);
xnor U361 (N_361,In_150,In_169);
nand U362 (N_362,In_359,In_126);
and U363 (N_363,In_231,In_471);
nor U364 (N_364,In_88,In_142);
nand U365 (N_365,In_49,In_456);
and U366 (N_366,In_312,In_438);
or U367 (N_367,In_242,In_289);
nand U368 (N_368,In_319,In_26);
nand U369 (N_369,In_478,In_262);
or U370 (N_370,In_48,In_0);
or U371 (N_371,In_433,In_490);
and U372 (N_372,In_154,In_39);
nand U373 (N_373,In_115,In_108);
or U374 (N_374,In_202,In_317);
xnor U375 (N_375,In_146,In_49);
nand U376 (N_376,In_407,In_259);
or U377 (N_377,In_107,In_455);
and U378 (N_378,In_199,In_266);
nor U379 (N_379,In_269,In_326);
and U380 (N_380,In_19,In_57);
or U381 (N_381,In_368,In_173);
and U382 (N_382,In_75,In_198);
or U383 (N_383,In_138,In_401);
or U384 (N_384,In_303,In_249);
nor U385 (N_385,In_381,In_303);
and U386 (N_386,In_395,In_396);
nor U387 (N_387,In_308,In_343);
nor U388 (N_388,In_399,In_44);
or U389 (N_389,In_255,In_360);
or U390 (N_390,In_115,In_237);
nand U391 (N_391,In_202,In_437);
nand U392 (N_392,In_468,In_12);
and U393 (N_393,In_83,In_350);
or U394 (N_394,In_254,In_182);
and U395 (N_395,In_296,In_303);
and U396 (N_396,In_98,In_358);
and U397 (N_397,In_348,In_241);
nand U398 (N_398,In_217,In_153);
nor U399 (N_399,In_346,In_108);
and U400 (N_400,In_383,In_13);
and U401 (N_401,In_130,In_52);
nor U402 (N_402,In_40,In_33);
nor U403 (N_403,In_275,In_399);
and U404 (N_404,In_305,In_41);
nand U405 (N_405,In_398,In_242);
nand U406 (N_406,In_138,In_374);
nand U407 (N_407,In_133,In_190);
nand U408 (N_408,In_376,In_157);
xnor U409 (N_409,In_232,In_115);
or U410 (N_410,In_284,In_486);
nand U411 (N_411,In_264,In_308);
nand U412 (N_412,In_385,In_479);
nor U413 (N_413,In_187,In_407);
nor U414 (N_414,In_151,In_299);
nor U415 (N_415,In_379,In_83);
nand U416 (N_416,In_306,In_10);
xor U417 (N_417,In_281,In_6);
and U418 (N_418,In_188,In_94);
and U419 (N_419,In_440,In_350);
xor U420 (N_420,In_318,In_109);
nand U421 (N_421,In_160,In_28);
or U422 (N_422,In_412,In_48);
or U423 (N_423,In_450,In_43);
or U424 (N_424,In_120,In_57);
nor U425 (N_425,In_70,In_393);
or U426 (N_426,In_305,In_325);
or U427 (N_427,In_300,In_252);
nand U428 (N_428,In_170,In_418);
nand U429 (N_429,In_261,In_128);
or U430 (N_430,In_75,In_458);
or U431 (N_431,In_328,In_413);
nand U432 (N_432,In_422,In_399);
nor U433 (N_433,In_343,In_212);
nor U434 (N_434,In_477,In_318);
or U435 (N_435,In_117,In_403);
xor U436 (N_436,In_350,In_140);
nor U437 (N_437,In_240,In_62);
or U438 (N_438,In_288,In_274);
or U439 (N_439,In_58,In_386);
nor U440 (N_440,In_347,In_375);
and U441 (N_441,In_157,In_419);
nor U442 (N_442,In_199,In_287);
nor U443 (N_443,In_89,In_36);
or U444 (N_444,In_461,In_358);
or U445 (N_445,In_464,In_106);
nor U446 (N_446,In_360,In_34);
and U447 (N_447,In_334,In_485);
xor U448 (N_448,In_261,In_33);
and U449 (N_449,In_116,In_499);
or U450 (N_450,In_413,In_279);
and U451 (N_451,In_314,In_41);
nor U452 (N_452,In_18,In_480);
nor U453 (N_453,In_360,In_359);
or U454 (N_454,In_303,In_443);
nand U455 (N_455,In_151,In_472);
xor U456 (N_456,In_262,In_277);
nor U457 (N_457,In_223,In_302);
nor U458 (N_458,In_178,In_252);
xnor U459 (N_459,In_141,In_103);
xor U460 (N_460,In_74,In_443);
or U461 (N_461,In_473,In_371);
nor U462 (N_462,In_56,In_283);
or U463 (N_463,In_442,In_437);
and U464 (N_464,In_118,In_367);
nand U465 (N_465,In_86,In_311);
xnor U466 (N_466,In_50,In_61);
nand U467 (N_467,In_345,In_116);
nand U468 (N_468,In_369,In_297);
nand U469 (N_469,In_386,In_473);
or U470 (N_470,In_347,In_346);
nor U471 (N_471,In_395,In_280);
nor U472 (N_472,In_431,In_427);
nand U473 (N_473,In_251,In_102);
or U474 (N_474,In_46,In_266);
nand U475 (N_475,In_121,In_88);
nor U476 (N_476,In_160,In_430);
nor U477 (N_477,In_419,In_41);
nor U478 (N_478,In_200,In_431);
or U479 (N_479,In_41,In_467);
and U480 (N_480,In_386,In_9);
or U481 (N_481,In_156,In_209);
and U482 (N_482,In_429,In_207);
or U483 (N_483,In_409,In_437);
and U484 (N_484,In_13,In_323);
nand U485 (N_485,In_354,In_25);
xor U486 (N_486,In_401,In_81);
nand U487 (N_487,In_51,In_153);
nand U488 (N_488,In_134,In_252);
nor U489 (N_489,In_1,In_46);
nand U490 (N_490,In_257,In_291);
and U491 (N_491,In_65,In_475);
or U492 (N_492,In_485,In_450);
nand U493 (N_493,In_451,In_290);
or U494 (N_494,In_445,In_461);
or U495 (N_495,In_475,In_404);
or U496 (N_496,In_382,In_463);
nand U497 (N_497,In_370,In_354);
or U498 (N_498,In_213,In_424);
and U499 (N_499,In_490,In_337);
xor U500 (N_500,In_231,In_312);
nand U501 (N_501,In_271,In_210);
nor U502 (N_502,In_479,In_131);
nand U503 (N_503,In_106,In_318);
nor U504 (N_504,In_370,In_429);
or U505 (N_505,In_387,In_206);
or U506 (N_506,In_384,In_484);
nand U507 (N_507,In_345,In_94);
or U508 (N_508,In_85,In_173);
and U509 (N_509,In_294,In_390);
nand U510 (N_510,In_303,In_441);
xor U511 (N_511,In_60,In_74);
and U512 (N_512,In_73,In_96);
xor U513 (N_513,In_368,In_396);
or U514 (N_514,In_444,In_299);
and U515 (N_515,In_215,In_427);
or U516 (N_516,In_453,In_215);
xnor U517 (N_517,In_118,In_423);
nand U518 (N_518,In_34,In_472);
xnor U519 (N_519,In_366,In_412);
or U520 (N_520,In_123,In_19);
nor U521 (N_521,In_336,In_339);
and U522 (N_522,In_40,In_9);
or U523 (N_523,In_142,In_462);
nor U524 (N_524,In_399,In_413);
nor U525 (N_525,In_455,In_328);
nand U526 (N_526,In_421,In_25);
and U527 (N_527,In_114,In_137);
and U528 (N_528,In_327,In_306);
and U529 (N_529,In_312,In_262);
nor U530 (N_530,In_378,In_267);
xnor U531 (N_531,In_328,In_166);
and U532 (N_532,In_216,In_163);
nand U533 (N_533,In_151,In_337);
or U534 (N_534,In_88,In_87);
nand U535 (N_535,In_497,In_131);
or U536 (N_536,In_495,In_356);
nand U537 (N_537,In_284,In_6);
or U538 (N_538,In_297,In_128);
or U539 (N_539,In_231,In_497);
or U540 (N_540,In_429,In_321);
and U541 (N_541,In_167,In_144);
nand U542 (N_542,In_115,In_399);
or U543 (N_543,In_13,In_181);
nand U544 (N_544,In_169,In_74);
and U545 (N_545,In_302,In_264);
nor U546 (N_546,In_219,In_249);
or U547 (N_547,In_337,In_217);
or U548 (N_548,In_208,In_148);
nand U549 (N_549,In_325,In_359);
or U550 (N_550,In_52,In_440);
and U551 (N_551,In_407,In_309);
nand U552 (N_552,In_278,In_9);
or U553 (N_553,In_190,In_462);
or U554 (N_554,In_422,In_245);
nand U555 (N_555,In_156,In_72);
and U556 (N_556,In_404,In_340);
xnor U557 (N_557,In_115,In_220);
nor U558 (N_558,In_73,In_23);
and U559 (N_559,In_39,In_29);
or U560 (N_560,In_114,In_99);
or U561 (N_561,In_256,In_186);
and U562 (N_562,In_407,In_236);
and U563 (N_563,In_444,In_131);
xor U564 (N_564,In_223,In_67);
nor U565 (N_565,In_92,In_2);
or U566 (N_566,In_426,In_210);
or U567 (N_567,In_308,In_440);
nor U568 (N_568,In_257,In_69);
nand U569 (N_569,In_138,In_173);
nor U570 (N_570,In_360,In_468);
or U571 (N_571,In_483,In_201);
xor U572 (N_572,In_106,In_349);
or U573 (N_573,In_17,In_74);
or U574 (N_574,In_129,In_87);
or U575 (N_575,In_187,In_320);
xor U576 (N_576,In_84,In_56);
xor U577 (N_577,In_251,In_343);
and U578 (N_578,In_40,In_238);
nand U579 (N_579,In_158,In_442);
nor U580 (N_580,In_399,In_304);
nand U581 (N_581,In_293,In_463);
xor U582 (N_582,In_471,In_455);
and U583 (N_583,In_261,In_73);
nand U584 (N_584,In_209,In_241);
nor U585 (N_585,In_110,In_224);
xnor U586 (N_586,In_281,In_435);
nand U587 (N_587,In_178,In_379);
or U588 (N_588,In_63,In_451);
xnor U589 (N_589,In_295,In_434);
or U590 (N_590,In_250,In_244);
or U591 (N_591,In_406,In_303);
and U592 (N_592,In_322,In_417);
and U593 (N_593,In_74,In_197);
or U594 (N_594,In_199,In_369);
nand U595 (N_595,In_109,In_471);
nand U596 (N_596,In_196,In_286);
and U597 (N_597,In_196,In_408);
nand U598 (N_598,In_120,In_482);
xor U599 (N_599,In_430,In_313);
or U600 (N_600,In_257,In_212);
nor U601 (N_601,In_64,In_101);
or U602 (N_602,In_161,In_427);
and U603 (N_603,In_214,In_443);
or U604 (N_604,In_15,In_189);
nor U605 (N_605,In_470,In_320);
xor U606 (N_606,In_26,In_463);
nand U607 (N_607,In_139,In_100);
or U608 (N_608,In_464,In_483);
or U609 (N_609,In_494,In_340);
nand U610 (N_610,In_70,In_493);
nand U611 (N_611,In_15,In_208);
xnor U612 (N_612,In_126,In_187);
xnor U613 (N_613,In_330,In_477);
xnor U614 (N_614,In_177,In_15);
and U615 (N_615,In_50,In_323);
and U616 (N_616,In_212,In_353);
or U617 (N_617,In_86,In_324);
or U618 (N_618,In_312,In_17);
nor U619 (N_619,In_377,In_151);
nand U620 (N_620,In_157,In_463);
nand U621 (N_621,In_194,In_180);
and U622 (N_622,In_443,In_273);
or U623 (N_623,In_109,In_273);
nand U624 (N_624,In_148,In_289);
or U625 (N_625,In_467,In_150);
nand U626 (N_626,In_464,In_465);
nand U627 (N_627,In_378,In_269);
nand U628 (N_628,In_348,In_134);
and U629 (N_629,In_61,In_334);
or U630 (N_630,In_95,In_10);
nand U631 (N_631,In_309,In_347);
xnor U632 (N_632,In_469,In_150);
nand U633 (N_633,In_58,In_145);
nor U634 (N_634,In_200,In_48);
and U635 (N_635,In_195,In_322);
nor U636 (N_636,In_395,In_99);
nand U637 (N_637,In_72,In_454);
nor U638 (N_638,In_83,In_365);
nor U639 (N_639,In_161,In_289);
nor U640 (N_640,In_252,In_448);
nand U641 (N_641,In_483,In_159);
nor U642 (N_642,In_347,In_340);
nor U643 (N_643,In_40,In_269);
xnor U644 (N_644,In_304,In_366);
nor U645 (N_645,In_413,In_113);
or U646 (N_646,In_269,In_359);
xnor U647 (N_647,In_287,In_81);
nor U648 (N_648,In_476,In_334);
or U649 (N_649,In_302,In_452);
nor U650 (N_650,In_147,In_243);
or U651 (N_651,In_227,In_356);
or U652 (N_652,In_497,In_426);
nand U653 (N_653,In_346,In_232);
nor U654 (N_654,In_257,In_379);
nand U655 (N_655,In_495,In_75);
and U656 (N_656,In_273,In_247);
nand U657 (N_657,In_338,In_44);
nand U658 (N_658,In_367,In_168);
nor U659 (N_659,In_72,In_410);
nand U660 (N_660,In_374,In_56);
or U661 (N_661,In_229,In_383);
or U662 (N_662,In_157,In_49);
and U663 (N_663,In_191,In_185);
nand U664 (N_664,In_111,In_278);
nand U665 (N_665,In_384,In_319);
xor U666 (N_666,In_494,In_388);
nor U667 (N_667,In_352,In_434);
or U668 (N_668,In_278,In_196);
nand U669 (N_669,In_312,In_273);
nand U670 (N_670,In_18,In_299);
nand U671 (N_671,In_298,In_294);
nand U672 (N_672,In_255,In_368);
nand U673 (N_673,In_102,In_388);
nand U674 (N_674,In_359,In_419);
xor U675 (N_675,In_147,In_230);
nor U676 (N_676,In_138,In_474);
or U677 (N_677,In_426,In_278);
or U678 (N_678,In_168,In_233);
nor U679 (N_679,In_163,In_49);
nand U680 (N_680,In_36,In_29);
nor U681 (N_681,In_459,In_180);
or U682 (N_682,In_435,In_230);
nand U683 (N_683,In_73,In_64);
or U684 (N_684,In_183,In_400);
or U685 (N_685,In_135,In_314);
or U686 (N_686,In_358,In_378);
or U687 (N_687,In_370,In_28);
nor U688 (N_688,In_401,In_0);
xnor U689 (N_689,In_42,In_86);
and U690 (N_690,In_478,In_49);
nor U691 (N_691,In_299,In_277);
or U692 (N_692,In_487,In_180);
nor U693 (N_693,In_131,In_222);
nand U694 (N_694,In_231,In_280);
nor U695 (N_695,In_5,In_468);
nor U696 (N_696,In_215,In_363);
nand U697 (N_697,In_494,In_361);
nand U698 (N_698,In_138,In_154);
or U699 (N_699,In_404,In_318);
xor U700 (N_700,In_328,In_243);
nand U701 (N_701,In_353,In_21);
or U702 (N_702,In_478,In_222);
nand U703 (N_703,In_417,In_112);
nor U704 (N_704,In_101,In_263);
xnor U705 (N_705,In_55,In_204);
or U706 (N_706,In_100,In_69);
nand U707 (N_707,In_39,In_63);
or U708 (N_708,In_6,In_111);
and U709 (N_709,In_210,In_127);
or U710 (N_710,In_339,In_22);
and U711 (N_711,In_274,In_94);
and U712 (N_712,In_416,In_95);
and U713 (N_713,In_59,In_109);
xnor U714 (N_714,In_117,In_52);
nor U715 (N_715,In_491,In_19);
and U716 (N_716,In_371,In_14);
or U717 (N_717,In_221,In_348);
nor U718 (N_718,In_498,In_436);
or U719 (N_719,In_418,In_100);
and U720 (N_720,In_103,In_499);
xor U721 (N_721,In_462,In_491);
nor U722 (N_722,In_341,In_136);
and U723 (N_723,In_72,In_427);
xnor U724 (N_724,In_166,In_397);
nand U725 (N_725,In_89,In_359);
and U726 (N_726,In_375,In_407);
xnor U727 (N_727,In_310,In_150);
nor U728 (N_728,In_83,In_419);
nor U729 (N_729,In_380,In_360);
or U730 (N_730,In_475,In_178);
nor U731 (N_731,In_434,In_330);
nor U732 (N_732,In_169,In_119);
nand U733 (N_733,In_129,In_314);
nand U734 (N_734,In_210,In_32);
nor U735 (N_735,In_400,In_148);
xor U736 (N_736,In_428,In_113);
nor U737 (N_737,In_309,In_334);
nand U738 (N_738,In_389,In_208);
nand U739 (N_739,In_306,In_419);
nor U740 (N_740,In_159,In_16);
or U741 (N_741,In_248,In_46);
nand U742 (N_742,In_341,In_221);
or U743 (N_743,In_170,In_19);
nand U744 (N_744,In_56,In_59);
nor U745 (N_745,In_136,In_106);
nor U746 (N_746,In_380,In_258);
nor U747 (N_747,In_306,In_356);
nor U748 (N_748,In_21,In_445);
nor U749 (N_749,In_419,In_295);
nand U750 (N_750,N_239,N_739);
nand U751 (N_751,N_546,N_63);
or U752 (N_752,N_200,N_749);
and U753 (N_753,N_424,N_324);
and U754 (N_754,N_641,N_561);
xor U755 (N_755,N_307,N_464);
nor U756 (N_756,N_402,N_562);
and U757 (N_757,N_625,N_181);
and U758 (N_758,N_488,N_446);
nand U759 (N_759,N_355,N_80);
nor U760 (N_760,N_320,N_408);
and U761 (N_761,N_353,N_194);
nor U762 (N_762,N_204,N_333);
and U763 (N_763,N_77,N_621);
nor U764 (N_764,N_727,N_737);
nor U765 (N_765,N_125,N_132);
and U766 (N_766,N_622,N_152);
nor U767 (N_767,N_157,N_213);
nand U768 (N_768,N_315,N_723);
and U769 (N_769,N_410,N_443);
xor U770 (N_770,N_109,N_235);
and U771 (N_771,N_187,N_26);
or U772 (N_772,N_559,N_260);
and U773 (N_773,N_107,N_663);
nand U774 (N_774,N_516,N_694);
nand U775 (N_775,N_198,N_159);
nand U776 (N_776,N_558,N_237);
or U777 (N_777,N_726,N_470);
nor U778 (N_778,N_454,N_334);
and U779 (N_779,N_648,N_614);
nor U780 (N_780,N_69,N_169);
nand U781 (N_781,N_602,N_719);
nor U782 (N_782,N_613,N_623);
or U783 (N_783,N_746,N_242);
and U784 (N_784,N_684,N_712);
nand U785 (N_785,N_441,N_345);
nor U786 (N_786,N_612,N_91);
nor U787 (N_787,N_369,N_645);
nor U788 (N_788,N_246,N_168);
or U789 (N_789,N_372,N_394);
nor U790 (N_790,N_23,N_225);
nor U791 (N_791,N_455,N_421);
or U792 (N_792,N_92,N_154);
nand U793 (N_793,N_126,N_31);
or U794 (N_794,N_747,N_177);
and U795 (N_795,N_388,N_227);
nor U796 (N_796,N_566,N_2);
and U797 (N_797,N_106,N_456);
nor U798 (N_798,N_180,N_356);
nand U799 (N_799,N_238,N_396);
and U800 (N_800,N_316,N_644);
nor U801 (N_801,N_722,N_318);
nand U802 (N_802,N_428,N_450);
nor U803 (N_803,N_277,N_474);
nand U804 (N_804,N_555,N_729);
or U805 (N_805,N_725,N_743);
nor U806 (N_806,N_32,N_76);
and U807 (N_807,N_733,N_53);
and U808 (N_808,N_512,N_607);
and U809 (N_809,N_64,N_635);
and U810 (N_810,N_147,N_111);
and U811 (N_811,N_68,N_496);
nand U812 (N_812,N_659,N_609);
and U813 (N_813,N_281,N_49);
or U814 (N_814,N_241,N_292);
and U815 (N_815,N_630,N_331);
nor U816 (N_816,N_585,N_425);
nor U817 (N_817,N_432,N_37);
and U818 (N_818,N_138,N_223);
and U819 (N_819,N_230,N_485);
nor U820 (N_820,N_8,N_461);
and U821 (N_821,N_536,N_270);
nor U822 (N_822,N_339,N_375);
xnor U823 (N_823,N_205,N_721);
and U824 (N_824,N_472,N_411);
nor U825 (N_825,N_224,N_453);
and U826 (N_826,N_104,N_211);
xnor U827 (N_827,N_604,N_321);
xor U828 (N_828,N_526,N_95);
nor U829 (N_829,N_337,N_459);
nand U830 (N_830,N_24,N_386);
nand U831 (N_831,N_403,N_278);
or U832 (N_832,N_423,N_574);
or U833 (N_833,N_709,N_549);
and U834 (N_834,N_553,N_710);
xnor U835 (N_835,N_415,N_473);
and U836 (N_836,N_702,N_244);
and U837 (N_837,N_48,N_185);
nand U838 (N_838,N_38,N_460);
nand U839 (N_839,N_540,N_681);
nand U840 (N_840,N_196,N_370);
nor U841 (N_841,N_151,N_517);
nor U842 (N_842,N_303,N_228);
nand U843 (N_843,N_218,N_184);
nand U844 (N_844,N_366,N_434);
or U845 (N_845,N_258,N_207);
or U846 (N_846,N_667,N_462);
or U847 (N_847,N_16,N_301);
nand U848 (N_848,N_458,N_673);
nand U849 (N_849,N_598,N_266);
xnor U850 (N_850,N_240,N_543);
and U851 (N_851,N_576,N_6);
or U852 (N_852,N_210,N_679);
nor U853 (N_853,N_409,N_275);
and U854 (N_854,N_309,N_18);
and U855 (N_855,N_678,N_121);
and U856 (N_856,N_43,N_490);
nor U857 (N_857,N_178,N_219);
or U858 (N_858,N_20,N_584);
nand U859 (N_859,N_166,N_542);
or U860 (N_860,N_478,N_52);
and U861 (N_861,N_59,N_267);
nand U862 (N_862,N_253,N_539);
and U863 (N_863,N_108,N_65);
and U864 (N_864,N_465,N_597);
nor U865 (N_865,N_362,N_509);
xor U866 (N_866,N_715,N_101);
nor U867 (N_867,N_530,N_136);
nand U868 (N_868,N_271,N_697);
nor U869 (N_869,N_544,N_689);
xnor U870 (N_870,N_497,N_98);
or U871 (N_871,N_222,N_717);
nor U872 (N_872,N_294,N_669);
nor U873 (N_873,N_305,N_256);
and U874 (N_874,N_564,N_554);
nand U875 (N_875,N_380,N_418);
nor U876 (N_876,N_62,N_664);
or U877 (N_877,N_385,N_4);
and U878 (N_878,N_550,N_588);
and U879 (N_879,N_164,N_534);
or U880 (N_880,N_170,N_519);
nor U881 (N_881,N_489,N_1);
nor U882 (N_882,N_39,N_600);
nand U883 (N_883,N_487,N_520);
nand U884 (N_884,N_482,N_329);
and U885 (N_885,N_420,N_274);
and U886 (N_886,N_313,N_736);
xnor U887 (N_887,N_261,N_680);
and U888 (N_888,N_273,N_378);
and U889 (N_889,N_720,N_67);
and U890 (N_890,N_647,N_595);
or U891 (N_891,N_58,N_259);
nand U892 (N_892,N_131,N_11);
nand U893 (N_893,N_572,N_269);
or U894 (N_894,N_35,N_404);
xor U895 (N_895,N_79,N_144);
or U896 (N_896,N_262,N_744);
nor U897 (N_897,N_188,N_633);
nor U898 (N_898,N_658,N_714);
xor U899 (N_899,N_646,N_636);
and U900 (N_900,N_118,N_703);
and U901 (N_901,N_72,N_155);
nand U902 (N_902,N_525,N_97);
or U903 (N_903,N_9,N_367);
nor U904 (N_904,N_21,N_78);
or U905 (N_905,N_300,N_390);
or U906 (N_906,N_165,N_405);
or U907 (N_907,N_389,N_344);
or U908 (N_908,N_156,N_413);
nand U909 (N_909,N_143,N_114);
nor U910 (N_910,N_548,N_399);
nor U911 (N_911,N_55,N_685);
or U912 (N_912,N_439,N_501);
nand U913 (N_913,N_603,N_384);
and U914 (N_914,N_234,N_51);
nand U915 (N_915,N_245,N_491);
or U916 (N_916,N_740,N_400);
and U917 (N_917,N_336,N_704);
nor U918 (N_918,N_247,N_427);
nand U919 (N_919,N_284,N_732);
nor U920 (N_920,N_265,N_93);
xor U921 (N_921,N_236,N_445);
and U922 (N_922,N_606,N_148);
xor U923 (N_923,N_383,N_652);
and U924 (N_924,N_128,N_656);
or U925 (N_925,N_671,N_422);
nand U926 (N_926,N_291,N_351);
and U927 (N_927,N_494,N_713);
xnor U928 (N_928,N_221,N_691);
nor U929 (N_929,N_575,N_568);
or U930 (N_930,N_706,N_172);
and U931 (N_931,N_475,N_708);
nand U932 (N_932,N_286,N_401);
or U933 (N_933,N_60,N_632);
or U934 (N_934,N_346,N_480);
and U935 (N_935,N_521,N_85);
nor U936 (N_936,N_73,N_96);
and U937 (N_937,N_532,N_731);
nand U938 (N_938,N_343,N_142);
nand U939 (N_939,N_297,N_387);
nor U940 (N_940,N_229,N_317);
and U941 (N_941,N_134,N_734);
or U942 (N_942,N_430,N_88);
nand U943 (N_943,N_451,N_586);
nand U944 (N_944,N_3,N_583);
nor U945 (N_945,N_493,N_699);
xnor U946 (N_946,N_611,N_416);
nor U947 (N_947,N_533,N_233);
or U948 (N_948,N_538,N_392);
nand U949 (N_949,N_208,N_202);
and U950 (N_950,N_440,N_735);
or U951 (N_951,N_677,N_406);
and U952 (N_952,N_249,N_359);
or U953 (N_953,N_327,N_655);
nand U954 (N_954,N_250,N_203);
or U955 (N_955,N_314,N_711);
or U956 (N_956,N_90,N_117);
and U957 (N_957,N_570,N_41);
and U958 (N_958,N_70,N_209);
or U959 (N_959,N_304,N_195);
and U960 (N_960,N_302,N_263);
nand U961 (N_961,N_13,N_57);
and U962 (N_962,N_513,N_199);
nand U963 (N_963,N_189,N_571);
nor U964 (N_964,N_44,N_212);
and U965 (N_965,N_14,N_174);
or U966 (N_966,N_190,N_433);
nor U967 (N_967,N_634,N_639);
nor U968 (N_968,N_398,N_582);
nor U969 (N_969,N_115,N_283);
and U970 (N_970,N_29,N_150);
or U971 (N_971,N_105,N_173);
nand U972 (N_972,N_466,N_193);
and U973 (N_973,N_25,N_524);
and U974 (N_974,N_183,N_395);
nand U975 (N_975,N_567,N_591);
and U976 (N_976,N_643,N_163);
and U977 (N_977,N_692,N_285);
nand U978 (N_978,N_654,N_569);
and U979 (N_979,N_676,N_0);
nor U980 (N_980,N_499,N_357);
and U981 (N_981,N_328,N_46);
or U982 (N_982,N_330,N_508);
nand U983 (N_983,N_87,N_522);
or U984 (N_984,N_463,N_672);
and U985 (N_985,N_518,N_123);
nor U986 (N_986,N_514,N_27);
xor U987 (N_987,N_146,N_354);
and U988 (N_988,N_730,N_310);
nor U989 (N_989,N_662,N_596);
or U990 (N_990,N_745,N_10);
or U991 (N_991,N_171,N_231);
or U992 (N_992,N_61,N_541);
xor U993 (N_993,N_500,N_119);
and U994 (N_994,N_577,N_718);
nand U995 (N_995,N_335,N_348);
xor U996 (N_996,N_688,N_360);
nor U997 (N_997,N_197,N_486);
or U998 (N_998,N_535,N_693);
nand U999 (N_999,N_338,N_153);
or U1000 (N_1000,N_298,N_374);
and U1001 (N_1001,N_299,N_528);
and U1002 (N_1002,N_593,N_99);
or U1003 (N_1003,N_272,N_627);
and U1004 (N_1004,N_220,N_120);
or U1005 (N_1005,N_54,N_340);
xnor U1006 (N_1006,N_137,N_74);
nor U1007 (N_1007,N_376,N_616);
nand U1008 (N_1008,N_363,N_206);
nand U1009 (N_1009,N_650,N_510);
or U1010 (N_1010,N_377,N_293);
and U1011 (N_1011,N_7,N_707);
nor U1012 (N_1012,N_129,N_638);
nor U1013 (N_1013,N_551,N_352);
xor U1014 (N_1014,N_332,N_12);
xor U1015 (N_1015,N_716,N_34);
nor U1016 (N_1016,N_545,N_17);
xor U1017 (N_1017,N_179,N_506);
xnor U1018 (N_1018,N_748,N_28);
or U1019 (N_1019,N_523,N_449);
or U1020 (N_1020,N_81,N_349);
or U1021 (N_1021,N_620,N_290);
or U1022 (N_1022,N_563,N_527);
nand U1023 (N_1023,N_36,N_492);
nor U1024 (N_1024,N_268,N_471);
and U1025 (N_1025,N_116,N_102);
or U1026 (N_1026,N_557,N_665);
and U1027 (N_1027,N_511,N_670);
or U1028 (N_1028,N_33,N_419);
xnor U1029 (N_1029,N_560,N_45);
nand U1030 (N_1030,N_312,N_214);
nand U1031 (N_1031,N_40,N_592);
or U1032 (N_1032,N_503,N_295);
nand U1033 (N_1033,N_252,N_201);
xnor U1034 (N_1034,N_47,N_502);
and U1035 (N_1035,N_217,N_15);
nand U1036 (N_1036,N_112,N_140);
nor U1037 (N_1037,N_637,N_690);
xnor U1038 (N_1038,N_468,N_407);
nor U1039 (N_1039,N_83,N_135);
and U1040 (N_1040,N_615,N_279);
nand U1041 (N_1041,N_580,N_323);
and U1042 (N_1042,N_365,N_495);
xnor U1043 (N_1043,N_599,N_608);
xnor U1044 (N_1044,N_589,N_556);
and U1045 (N_1045,N_447,N_226);
nor U1046 (N_1046,N_182,N_122);
nor U1047 (N_1047,N_617,N_476);
and U1048 (N_1048,N_5,N_139);
or U1049 (N_1049,N_86,N_547);
nand U1050 (N_1050,N_373,N_287);
and U1051 (N_1051,N_381,N_186);
or U1052 (N_1052,N_368,N_113);
nor U1053 (N_1053,N_103,N_660);
nand U1054 (N_1054,N_705,N_431);
nand U1055 (N_1055,N_695,N_435);
and U1056 (N_1056,N_624,N_393);
and U1057 (N_1057,N_71,N_243);
and U1058 (N_1058,N_232,N_700);
or U1059 (N_1059,N_573,N_361);
or U1060 (N_1060,N_133,N_601);
or U1061 (N_1061,N_657,N_498);
nor U1062 (N_1062,N_412,N_444);
nand U1063 (N_1063,N_724,N_537);
nand U1064 (N_1064,N_683,N_110);
or U1065 (N_1065,N_30,N_149);
or U1066 (N_1066,N_326,N_280);
xnor U1067 (N_1067,N_429,N_145);
nor U1068 (N_1068,N_127,N_22);
and U1069 (N_1069,N_618,N_176);
nand U1070 (N_1070,N_565,N_649);
and U1071 (N_1071,N_100,N_282);
nor U1072 (N_1072,N_619,N_426);
nor U1073 (N_1073,N_319,N_590);
and U1074 (N_1074,N_162,N_610);
and U1075 (N_1075,N_322,N_668);
or U1076 (N_1076,N_391,N_653);
xor U1077 (N_1077,N_579,N_50);
xnor U1078 (N_1078,N_289,N_255);
nor U1079 (N_1079,N_436,N_481);
or U1080 (N_1080,N_75,N_191);
nor U1081 (N_1081,N_483,N_728);
nand U1082 (N_1082,N_379,N_417);
and U1083 (N_1083,N_437,N_306);
xnor U1084 (N_1084,N_741,N_587);
nand U1085 (N_1085,N_452,N_342);
or U1086 (N_1086,N_371,N_124);
nand U1087 (N_1087,N_66,N_504);
or U1088 (N_1088,N_257,N_311);
nand U1089 (N_1089,N_640,N_251);
nor U1090 (N_1090,N_505,N_161);
nor U1091 (N_1091,N_442,N_56);
nor U1092 (N_1092,N_581,N_84);
and U1093 (N_1093,N_254,N_469);
or U1094 (N_1094,N_82,N_160);
nor U1095 (N_1095,N_605,N_288);
and U1096 (N_1096,N_642,N_529);
or U1097 (N_1097,N_479,N_738);
and U1098 (N_1098,N_594,N_515);
nor U1099 (N_1099,N_19,N_675);
nand U1100 (N_1100,N_552,N_467);
or U1101 (N_1101,N_698,N_631);
and U1102 (N_1102,N_477,N_175);
nand U1103 (N_1103,N_158,N_696);
and U1104 (N_1104,N_629,N_325);
nor U1105 (N_1105,N_661,N_42);
and U1106 (N_1106,N_674,N_742);
and U1107 (N_1107,N_484,N_457);
and U1108 (N_1108,N_686,N_666);
and U1109 (N_1109,N_626,N_130);
or U1110 (N_1110,N_531,N_264);
nand U1111 (N_1111,N_215,N_341);
nand U1112 (N_1112,N_701,N_578);
or U1113 (N_1113,N_382,N_651);
and U1114 (N_1114,N_397,N_358);
and U1115 (N_1115,N_507,N_216);
or U1116 (N_1116,N_347,N_94);
nor U1117 (N_1117,N_414,N_438);
nand U1118 (N_1118,N_350,N_364);
and U1119 (N_1119,N_628,N_141);
and U1120 (N_1120,N_276,N_89);
nor U1121 (N_1121,N_192,N_682);
nand U1122 (N_1122,N_448,N_296);
or U1123 (N_1123,N_308,N_248);
nor U1124 (N_1124,N_167,N_687);
or U1125 (N_1125,N_577,N_15);
or U1126 (N_1126,N_363,N_717);
nor U1127 (N_1127,N_388,N_549);
or U1128 (N_1128,N_40,N_185);
and U1129 (N_1129,N_669,N_319);
or U1130 (N_1130,N_365,N_509);
nand U1131 (N_1131,N_654,N_596);
and U1132 (N_1132,N_557,N_498);
nand U1133 (N_1133,N_29,N_312);
nor U1134 (N_1134,N_649,N_615);
nand U1135 (N_1135,N_380,N_54);
or U1136 (N_1136,N_256,N_166);
nor U1137 (N_1137,N_609,N_8);
and U1138 (N_1138,N_38,N_574);
and U1139 (N_1139,N_530,N_347);
nor U1140 (N_1140,N_269,N_221);
or U1141 (N_1141,N_44,N_268);
nand U1142 (N_1142,N_456,N_690);
or U1143 (N_1143,N_220,N_575);
nor U1144 (N_1144,N_478,N_40);
nor U1145 (N_1145,N_639,N_168);
or U1146 (N_1146,N_338,N_160);
nor U1147 (N_1147,N_547,N_347);
nor U1148 (N_1148,N_187,N_252);
nor U1149 (N_1149,N_422,N_555);
and U1150 (N_1150,N_602,N_491);
nand U1151 (N_1151,N_138,N_117);
xor U1152 (N_1152,N_304,N_572);
or U1153 (N_1153,N_96,N_55);
and U1154 (N_1154,N_746,N_302);
xnor U1155 (N_1155,N_296,N_398);
and U1156 (N_1156,N_270,N_703);
xor U1157 (N_1157,N_261,N_6);
or U1158 (N_1158,N_151,N_622);
nand U1159 (N_1159,N_523,N_252);
nor U1160 (N_1160,N_631,N_357);
and U1161 (N_1161,N_721,N_197);
and U1162 (N_1162,N_45,N_526);
and U1163 (N_1163,N_114,N_129);
nand U1164 (N_1164,N_107,N_305);
and U1165 (N_1165,N_372,N_534);
or U1166 (N_1166,N_401,N_180);
and U1167 (N_1167,N_617,N_411);
nor U1168 (N_1168,N_211,N_298);
xor U1169 (N_1169,N_246,N_71);
nor U1170 (N_1170,N_655,N_437);
nor U1171 (N_1171,N_633,N_359);
or U1172 (N_1172,N_369,N_235);
and U1173 (N_1173,N_638,N_473);
nand U1174 (N_1174,N_226,N_507);
or U1175 (N_1175,N_103,N_176);
or U1176 (N_1176,N_514,N_637);
nand U1177 (N_1177,N_572,N_147);
xor U1178 (N_1178,N_155,N_678);
or U1179 (N_1179,N_578,N_452);
xor U1180 (N_1180,N_109,N_496);
nand U1181 (N_1181,N_214,N_672);
or U1182 (N_1182,N_578,N_405);
nor U1183 (N_1183,N_265,N_722);
nor U1184 (N_1184,N_419,N_321);
or U1185 (N_1185,N_84,N_173);
nor U1186 (N_1186,N_434,N_744);
nand U1187 (N_1187,N_487,N_442);
nor U1188 (N_1188,N_431,N_742);
nand U1189 (N_1189,N_27,N_227);
nand U1190 (N_1190,N_578,N_333);
xnor U1191 (N_1191,N_551,N_233);
nor U1192 (N_1192,N_299,N_135);
nor U1193 (N_1193,N_611,N_738);
or U1194 (N_1194,N_544,N_314);
and U1195 (N_1195,N_663,N_722);
or U1196 (N_1196,N_169,N_201);
or U1197 (N_1197,N_682,N_439);
and U1198 (N_1198,N_87,N_663);
nor U1199 (N_1199,N_222,N_662);
nor U1200 (N_1200,N_508,N_701);
and U1201 (N_1201,N_304,N_446);
and U1202 (N_1202,N_604,N_397);
nor U1203 (N_1203,N_596,N_1);
nand U1204 (N_1204,N_587,N_418);
nand U1205 (N_1205,N_220,N_646);
and U1206 (N_1206,N_69,N_495);
and U1207 (N_1207,N_254,N_436);
nand U1208 (N_1208,N_607,N_596);
nand U1209 (N_1209,N_503,N_489);
or U1210 (N_1210,N_80,N_571);
nor U1211 (N_1211,N_568,N_71);
xor U1212 (N_1212,N_708,N_346);
nand U1213 (N_1213,N_250,N_129);
nor U1214 (N_1214,N_55,N_291);
and U1215 (N_1215,N_685,N_345);
or U1216 (N_1216,N_227,N_324);
nor U1217 (N_1217,N_576,N_207);
or U1218 (N_1218,N_185,N_487);
and U1219 (N_1219,N_403,N_308);
and U1220 (N_1220,N_376,N_421);
nor U1221 (N_1221,N_460,N_458);
or U1222 (N_1222,N_353,N_125);
nor U1223 (N_1223,N_696,N_206);
nor U1224 (N_1224,N_350,N_430);
or U1225 (N_1225,N_336,N_438);
nand U1226 (N_1226,N_744,N_392);
nand U1227 (N_1227,N_468,N_202);
and U1228 (N_1228,N_264,N_341);
and U1229 (N_1229,N_347,N_656);
nor U1230 (N_1230,N_61,N_625);
nand U1231 (N_1231,N_621,N_726);
nor U1232 (N_1232,N_677,N_293);
or U1233 (N_1233,N_328,N_540);
or U1234 (N_1234,N_118,N_463);
and U1235 (N_1235,N_130,N_542);
nor U1236 (N_1236,N_12,N_492);
xor U1237 (N_1237,N_79,N_53);
nand U1238 (N_1238,N_214,N_399);
nor U1239 (N_1239,N_174,N_87);
or U1240 (N_1240,N_360,N_404);
nand U1241 (N_1241,N_393,N_203);
and U1242 (N_1242,N_111,N_145);
nand U1243 (N_1243,N_587,N_511);
and U1244 (N_1244,N_36,N_13);
nand U1245 (N_1245,N_493,N_468);
nand U1246 (N_1246,N_93,N_14);
nor U1247 (N_1247,N_56,N_429);
nor U1248 (N_1248,N_506,N_586);
xnor U1249 (N_1249,N_675,N_129);
nand U1250 (N_1250,N_124,N_683);
nor U1251 (N_1251,N_175,N_59);
or U1252 (N_1252,N_509,N_288);
or U1253 (N_1253,N_349,N_691);
or U1254 (N_1254,N_336,N_300);
nand U1255 (N_1255,N_124,N_553);
and U1256 (N_1256,N_243,N_162);
and U1257 (N_1257,N_18,N_82);
nand U1258 (N_1258,N_396,N_260);
nor U1259 (N_1259,N_367,N_662);
xor U1260 (N_1260,N_657,N_33);
xnor U1261 (N_1261,N_169,N_612);
nor U1262 (N_1262,N_728,N_143);
and U1263 (N_1263,N_627,N_225);
nor U1264 (N_1264,N_86,N_368);
and U1265 (N_1265,N_304,N_164);
nand U1266 (N_1266,N_694,N_486);
nor U1267 (N_1267,N_171,N_304);
nor U1268 (N_1268,N_613,N_285);
nor U1269 (N_1269,N_125,N_292);
nand U1270 (N_1270,N_251,N_346);
xnor U1271 (N_1271,N_553,N_222);
or U1272 (N_1272,N_490,N_276);
nor U1273 (N_1273,N_259,N_352);
nor U1274 (N_1274,N_384,N_356);
and U1275 (N_1275,N_292,N_383);
nor U1276 (N_1276,N_365,N_670);
xor U1277 (N_1277,N_88,N_365);
xnor U1278 (N_1278,N_242,N_309);
xor U1279 (N_1279,N_30,N_169);
and U1280 (N_1280,N_266,N_710);
nand U1281 (N_1281,N_188,N_51);
nand U1282 (N_1282,N_506,N_633);
nand U1283 (N_1283,N_694,N_749);
or U1284 (N_1284,N_239,N_300);
nand U1285 (N_1285,N_216,N_109);
nand U1286 (N_1286,N_201,N_577);
nand U1287 (N_1287,N_80,N_25);
nand U1288 (N_1288,N_533,N_328);
and U1289 (N_1289,N_695,N_339);
and U1290 (N_1290,N_480,N_377);
or U1291 (N_1291,N_550,N_168);
and U1292 (N_1292,N_55,N_707);
nor U1293 (N_1293,N_219,N_547);
and U1294 (N_1294,N_183,N_542);
or U1295 (N_1295,N_265,N_502);
or U1296 (N_1296,N_673,N_507);
or U1297 (N_1297,N_439,N_228);
or U1298 (N_1298,N_686,N_282);
nand U1299 (N_1299,N_53,N_674);
or U1300 (N_1300,N_400,N_143);
and U1301 (N_1301,N_300,N_653);
xnor U1302 (N_1302,N_2,N_61);
nor U1303 (N_1303,N_675,N_497);
nand U1304 (N_1304,N_202,N_102);
or U1305 (N_1305,N_269,N_261);
or U1306 (N_1306,N_143,N_636);
or U1307 (N_1307,N_659,N_437);
nand U1308 (N_1308,N_670,N_27);
and U1309 (N_1309,N_684,N_82);
nor U1310 (N_1310,N_432,N_527);
nor U1311 (N_1311,N_3,N_377);
or U1312 (N_1312,N_615,N_546);
nand U1313 (N_1313,N_650,N_379);
and U1314 (N_1314,N_213,N_715);
and U1315 (N_1315,N_652,N_78);
nand U1316 (N_1316,N_130,N_77);
and U1317 (N_1317,N_104,N_516);
nor U1318 (N_1318,N_103,N_88);
nor U1319 (N_1319,N_463,N_181);
or U1320 (N_1320,N_447,N_342);
nand U1321 (N_1321,N_738,N_580);
nor U1322 (N_1322,N_474,N_431);
nor U1323 (N_1323,N_400,N_725);
or U1324 (N_1324,N_151,N_503);
nor U1325 (N_1325,N_227,N_176);
nor U1326 (N_1326,N_320,N_504);
and U1327 (N_1327,N_282,N_675);
and U1328 (N_1328,N_128,N_209);
nand U1329 (N_1329,N_629,N_712);
or U1330 (N_1330,N_9,N_78);
nor U1331 (N_1331,N_86,N_4);
and U1332 (N_1332,N_489,N_559);
and U1333 (N_1333,N_261,N_591);
nor U1334 (N_1334,N_525,N_328);
nand U1335 (N_1335,N_221,N_472);
and U1336 (N_1336,N_642,N_113);
and U1337 (N_1337,N_365,N_352);
or U1338 (N_1338,N_98,N_486);
nand U1339 (N_1339,N_67,N_217);
nand U1340 (N_1340,N_183,N_386);
nor U1341 (N_1341,N_648,N_189);
nand U1342 (N_1342,N_436,N_483);
and U1343 (N_1343,N_534,N_689);
xor U1344 (N_1344,N_484,N_297);
nor U1345 (N_1345,N_228,N_643);
or U1346 (N_1346,N_623,N_212);
nor U1347 (N_1347,N_557,N_409);
nor U1348 (N_1348,N_131,N_432);
or U1349 (N_1349,N_587,N_739);
nor U1350 (N_1350,N_320,N_18);
nand U1351 (N_1351,N_144,N_531);
nand U1352 (N_1352,N_329,N_458);
or U1353 (N_1353,N_324,N_635);
and U1354 (N_1354,N_415,N_112);
nand U1355 (N_1355,N_545,N_638);
nand U1356 (N_1356,N_334,N_184);
nor U1357 (N_1357,N_734,N_695);
nand U1358 (N_1358,N_361,N_649);
and U1359 (N_1359,N_147,N_235);
nand U1360 (N_1360,N_10,N_564);
nor U1361 (N_1361,N_2,N_273);
or U1362 (N_1362,N_213,N_266);
nand U1363 (N_1363,N_356,N_558);
and U1364 (N_1364,N_403,N_670);
nor U1365 (N_1365,N_85,N_100);
nor U1366 (N_1366,N_579,N_695);
or U1367 (N_1367,N_144,N_243);
or U1368 (N_1368,N_497,N_94);
and U1369 (N_1369,N_706,N_713);
and U1370 (N_1370,N_514,N_365);
nor U1371 (N_1371,N_476,N_551);
xnor U1372 (N_1372,N_221,N_478);
nor U1373 (N_1373,N_1,N_657);
nor U1374 (N_1374,N_450,N_469);
and U1375 (N_1375,N_505,N_62);
nor U1376 (N_1376,N_731,N_517);
or U1377 (N_1377,N_281,N_312);
xor U1378 (N_1378,N_744,N_736);
or U1379 (N_1379,N_60,N_474);
nor U1380 (N_1380,N_733,N_311);
nand U1381 (N_1381,N_479,N_643);
or U1382 (N_1382,N_19,N_717);
nand U1383 (N_1383,N_145,N_647);
or U1384 (N_1384,N_186,N_69);
and U1385 (N_1385,N_428,N_35);
nor U1386 (N_1386,N_275,N_242);
nand U1387 (N_1387,N_75,N_744);
nand U1388 (N_1388,N_185,N_329);
nor U1389 (N_1389,N_138,N_408);
or U1390 (N_1390,N_433,N_186);
and U1391 (N_1391,N_248,N_732);
or U1392 (N_1392,N_692,N_364);
or U1393 (N_1393,N_250,N_704);
and U1394 (N_1394,N_82,N_422);
and U1395 (N_1395,N_95,N_743);
xnor U1396 (N_1396,N_185,N_227);
nor U1397 (N_1397,N_192,N_745);
and U1398 (N_1398,N_474,N_119);
nand U1399 (N_1399,N_207,N_186);
nand U1400 (N_1400,N_100,N_103);
or U1401 (N_1401,N_487,N_144);
nor U1402 (N_1402,N_570,N_676);
nor U1403 (N_1403,N_75,N_422);
xor U1404 (N_1404,N_641,N_484);
nand U1405 (N_1405,N_262,N_25);
xor U1406 (N_1406,N_491,N_439);
and U1407 (N_1407,N_152,N_730);
or U1408 (N_1408,N_580,N_644);
xor U1409 (N_1409,N_490,N_247);
nor U1410 (N_1410,N_7,N_737);
nor U1411 (N_1411,N_565,N_709);
nor U1412 (N_1412,N_169,N_659);
or U1413 (N_1413,N_589,N_572);
nor U1414 (N_1414,N_69,N_113);
or U1415 (N_1415,N_326,N_425);
nand U1416 (N_1416,N_571,N_402);
and U1417 (N_1417,N_242,N_262);
or U1418 (N_1418,N_486,N_645);
and U1419 (N_1419,N_677,N_617);
or U1420 (N_1420,N_97,N_625);
or U1421 (N_1421,N_457,N_332);
or U1422 (N_1422,N_145,N_7);
xnor U1423 (N_1423,N_63,N_379);
xnor U1424 (N_1424,N_321,N_491);
or U1425 (N_1425,N_579,N_88);
nor U1426 (N_1426,N_303,N_95);
and U1427 (N_1427,N_594,N_724);
nor U1428 (N_1428,N_491,N_512);
nor U1429 (N_1429,N_171,N_386);
and U1430 (N_1430,N_337,N_95);
and U1431 (N_1431,N_511,N_442);
and U1432 (N_1432,N_517,N_670);
or U1433 (N_1433,N_198,N_729);
nor U1434 (N_1434,N_651,N_371);
and U1435 (N_1435,N_279,N_716);
or U1436 (N_1436,N_745,N_128);
or U1437 (N_1437,N_42,N_439);
nand U1438 (N_1438,N_374,N_182);
xor U1439 (N_1439,N_80,N_168);
or U1440 (N_1440,N_224,N_519);
nor U1441 (N_1441,N_313,N_504);
nor U1442 (N_1442,N_328,N_595);
or U1443 (N_1443,N_157,N_627);
and U1444 (N_1444,N_702,N_706);
nor U1445 (N_1445,N_445,N_226);
and U1446 (N_1446,N_530,N_689);
or U1447 (N_1447,N_62,N_522);
and U1448 (N_1448,N_724,N_173);
nand U1449 (N_1449,N_199,N_663);
or U1450 (N_1450,N_444,N_382);
xnor U1451 (N_1451,N_489,N_78);
nor U1452 (N_1452,N_375,N_371);
or U1453 (N_1453,N_690,N_312);
or U1454 (N_1454,N_355,N_9);
xor U1455 (N_1455,N_12,N_514);
and U1456 (N_1456,N_566,N_462);
xnor U1457 (N_1457,N_172,N_222);
or U1458 (N_1458,N_685,N_301);
nand U1459 (N_1459,N_230,N_461);
nand U1460 (N_1460,N_368,N_4);
nor U1461 (N_1461,N_686,N_320);
or U1462 (N_1462,N_166,N_26);
and U1463 (N_1463,N_485,N_568);
or U1464 (N_1464,N_446,N_558);
or U1465 (N_1465,N_468,N_470);
xnor U1466 (N_1466,N_320,N_388);
nand U1467 (N_1467,N_159,N_707);
nand U1468 (N_1468,N_607,N_259);
xnor U1469 (N_1469,N_491,N_523);
and U1470 (N_1470,N_55,N_604);
nand U1471 (N_1471,N_191,N_71);
nand U1472 (N_1472,N_575,N_29);
nor U1473 (N_1473,N_404,N_474);
nand U1474 (N_1474,N_315,N_583);
nor U1475 (N_1475,N_291,N_136);
and U1476 (N_1476,N_3,N_101);
xnor U1477 (N_1477,N_656,N_12);
and U1478 (N_1478,N_133,N_115);
xnor U1479 (N_1479,N_241,N_101);
nand U1480 (N_1480,N_740,N_244);
and U1481 (N_1481,N_2,N_684);
nor U1482 (N_1482,N_538,N_465);
nand U1483 (N_1483,N_620,N_570);
or U1484 (N_1484,N_77,N_513);
or U1485 (N_1485,N_393,N_652);
nand U1486 (N_1486,N_178,N_259);
nor U1487 (N_1487,N_583,N_338);
nor U1488 (N_1488,N_154,N_49);
nor U1489 (N_1489,N_629,N_521);
and U1490 (N_1490,N_256,N_410);
and U1491 (N_1491,N_583,N_179);
or U1492 (N_1492,N_576,N_629);
xnor U1493 (N_1493,N_592,N_676);
xnor U1494 (N_1494,N_73,N_565);
nor U1495 (N_1495,N_727,N_746);
nand U1496 (N_1496,N_159,N_264);
or U1497 (N_1497,N_519,N_152);
or U1498 (N_1498,N_390,N_144);
and U1499 (N_1499,N_103,N_269);
nor U1500 (N_1500,N_1312,N_1322);
nand U1501 (N_1501,N_1232,N_911);
xnor U1502 (N_1502,N_962,N_1198);
nand U1503 (N_1503,N_1490,N_1214);
nor U1504 (N_1504,N_1274,N_906);
xor U1505 (N_1505,N_1083,N_1047);
or U1506 (N_1506,N_1174,N_811);
xor U1507 (N_1507,N_916,N_819);
nand U1508 (N_1508,N_780,N_814);
and U1509 (N_1509,N_1295,N_781);
nor U1510 (N_1510,N_1375,N_1045);
nand U1511 (N_1511,N_1488,N_798);
nand U1512 (N_1512,N_800,N_1075);
xnor U1513 (N_1513,N_1300,N_1194);
or U1514 (N_1514,N_1122,N_1081);
or U1515 (N_1515,N_1285,N_1230);
nor U1516 (N_1516,N_1210,N_1357);
nor U1517 (N_1517,N_970,N_754);
and U1518 (N_1518,N_961,N_1186);
nand U1519 (N_1519,N_776,N_1197);
nand U1520 (N_1520,N_824,N_1044);
nor U1521 (N_1521,N_1138,N_834);
or U1522 (N_1522,N_1199,N_1413);
nor U1523 (N_1523,N_1036,N_950);
and U1524 (N_1524,N_1024,N_1076);
or U1525 (N_1525,N_989,N_1241);
nor U1526 (N_1526,N_991,N_1067);
nor U1527 (N_1527,N_1016,N_851);
nand U1528 (N_1528,N_974,N_979);
nand U1529 (N_1529,N_1273,N_1127);
and U1530 (N_1530,N_1203,N_1020);
or U1531 (N_1531,N_1021,N_1008);
and U1532 (N_1532,N_1330,N_1046);
nand U1533 (N_1533,N_964,N_809);
nand U1534 (N_1534,N_1443,N_765);
or U1535 (N_1535,N_1053,N_1360);
or U1536 (N_1536,N_1004,N_1124);
nor U1537 (N_1537,N_817,N_1377);
and U1538 (N_1538,N_1037,N_1325);
nor U1539 (N_1539,N_1347,N_827);
nand U1540 (N_1540,N_758,N_1227);
nand U1541 (N_1541,N_909,N_905);
and U1542 (N_1542,N_874,N_1183);
and U1543 (N_1543,N_1048,N_772);
nor U1544 (N_1544,N_1050,N_857);
and U1545 (N_1545,N_930,N_1001);
and U1546 (N_1546,N_1104,N_1324);
and U1547 (N_1547,N_1305,N_1267);
or U1548 (N_1548,N_893,N_1465);
or U1549 (N_1549,N_1249,N_1028);
nor U1550 (N_1550,N_802,N_1421);
nand U1551 (N_1551,N_869,N_1329);
and U1552 (N_1552,N_1384,N_820);
xor U1553 (N_1553,N_1304,N_1137);
xor U1554 (N_1554,N_1407,N_790);
and U1555 (N_1555,N_1337,N_1040);
nand U1556 (N_1556,N_779,N_1383);
and U1557 (N_1557,N_1074,N_1463);
xnor U1558 (N_1558,N_1298,N_993);
nor U1559 (N_1559,N_1181,N_915);
or U1560 (N_1560,N_1299,N_1378);
nand U1561 (N_1561,N_902,N_1121);
or U1562 (N_1562,N_1073,N_990);
nand U1563 (N_1563,N_1253,N_789);
nor U1564 (N_1564,N_870,N_888);
nor U1565 (N_1565,N_1255,N_968);
nor U1566 (N_1566,N_1148,N_813);
nor U1567 (N_1567,N_1234,N_1182);
nor U1568 (N_1568,N_1428,N_969);
or U1569 (N_1569,N_978,N_1229);
xnor U1570 (N_1570,N_1101,N_1376);
and U1571 (N_1571,N_1495,N_1043);
and U1572 (N_1572,N_1344,N_1158);
nor U1573 (N_1573,N_882,N_1132);
and U1574 (N_1574,N_1240,N_1339);
and U1575 (N_1575,N_951,N_1291);
or U1576 (N_1576,N_821,N_1417);
and U1577 (N_1577,N_823,N_997);
and U1578 (N_1578,N_895,N_1464);
or U1579 (N_1579,N_1152,N_887);
nor U1580 (N_1580,N_988,N_1320);
nor U1581 (N_1581,N_1477,N_822);
and U1582 (N_1582,N_1366,N_1187);
nor U1583 (N_1583,N_1473,N_1301);
and U1584 (N_1584,N_904,N_762);
or U1585 (N_1585,N_1368,N_1331);
or U1586 (N_1586,N_799,N_1139);
xor U1587 (N_1587,N_1089,N_1434);
and U1588 (N_1588,N_897,N_883);
and U1589 (N_1589,N_879,N_833);
nand U1590 (N_1590,N_1052,N_1367);
or U1591 (N_1591,N_1475,N_770);
nand U1592 (N_1592,N_1491,N_1061);
nor U1593 (N_1593,N_1119,N_1007);
or U1594 (N_1594,N_1173,N_1235);
or U1595 (N_1595,N_1115,N_1480);
nor U1596 (N_1596,N_1242,N_1420);
nor U1597 (N_1597,N_898,N_1486);
nor U1598 (N_1598,N_995,N_808);
and U1599 (N_1599,N_1015,N_1387);
nor U1600 (N_1600,N_865,N_1270);
nand U1601 (N_1601,N_1146,N_1144);
or U1602 (N_1602,N_1401,N_1030);
xnor U1603 (N_1603,N_1391,N_1211);
or U1604 (N_1604,N_1003,N_1216);
or U1605 (N_1605,N_1063,N_1245);
or U1606 (N_1606,N_1114,N_1078);
or U1607 (N_1607,N_1314,N_977);
xor U1608 (N_1608,N_848,N_1151);
or U1609 (N_1609,N_1123,N_1389);
nand U1610 (N_1610,N_1429,N_949);
nor U1611 (N_1611,N_839,N_1056);
nor U1612 (N_1612,N_1257,N_1208);
and U1613 (N_1613,N_1260,N_1147);
nand U1614 (N_1614,N_1411,N_998);
and U1615 (N_1615,N_1239,N_1039);
xnor U1616 (N_1616,N_1354,N_1497);
nor U1617 (N_1617,N_1275,N_1281);
and U1618 (N_1618,N_1102,N_1470);
nand U1619 (N_1619,N_1057,N_1458);
or U1620 (N_1620,N_1358,N_1080);
and U1621 (N_1621,N_1447,N_1394);
and U1622 (N_1622,N_1129,N_788);
and U1623 (N_1623,N_816,N_1088);
nor U1624 (N_1624,N_1436,N_1205);
nand U1625 (N_1625,N_1409,N_1361);
or U1626 (N_1626,N_1496,N_1499);
nand U1627 (N_1627,N_1019,N_1091);
and U1628 (N_1628,N_875,N_1489);
nand U1629 (N_1629,N_1029,N_1031);
or U1630 (N_1630,N_1193,N_1476);
nand U1631 (N_1631,N_914,N_838);
or U1632 (N_1632,N_1113,N_981);
nor U1633 (N_1633,N_1290,N_1396);
nor U1634 (N_1634,N_1334,N_1397);
nand U1635 (N_1635,N_885,N_1335);
nand U1636 (N_1636,N_1392,N_761);
or U1637 (N_1637,N_1192,N_1390);
or U1638 (N_1638,N_1185,N_1303);
and U1639 (N_1639,N_1467,N_957);
and U1640 (N_1640,N_1224,N_1209);
or U1641 (N_1641,N_972,N_766);
or U1642 (N_1642,N_1365,N_1177);
nand U1643 (N_1643,N_1051,N_1092);
and U1644 (N_1644,N_1005,N_1084);
or U1645 (N_1645,N_1131,N_987);
nor U1646 (N_1646,N_1439,N_1018);
nor U1647 (N_1647,N_1450,N_1317);
xnor U1648 (N_1648,N_1425,N_803);
or U1649 (N_1649,N_944,N_1445);
or U1650 (N_1650,N_1179,N_878);
or U1651 (N_1651,N_965,N_891);
and U1652 (N_1652,N_900,N_1220);
and U1653 (N_1653,N_830,N_931);
nand U1654 (N_1654,N_928,N_1374);
nand U1655 (N_1655,N_1195,N_919);
nand U1656 (N_1656,N_1072,N_1379);
nor U1657 (N_1657,N_1117,N_984);
nand U1658 (N_1658,N_877,N_941);
and U1659 (N_1659,N_880,N_1481);
or U1660 (N_1660,N_1041,N_1180);
nor U1661 (N_1661,N_831,N_756);
nand U1662 (N_1662,N_1012,N_1427);
nand U1663 (N_1663,N_976,N_1103);
xor U1664 (N_1664,N_1049,N_1318);
nand U1665 (N_1665,N_1090,N_1125);
or U1666 (N_1666,N_908,N_1297);
nor U1667 (N_1667,N_1424,N_948);
or U1668 (N_1668,N_1011,N_926);
nand U1669 (N_1669,N_1190,N_1065);
nor U1670 (N_1670,N_1448,N_1444);
or U1671 (N_1671,N_1009,N_892);
nand U1672 (N_1672,N_1286,N_959);
nand U1673 (N_1673,N_1404,N_782);
or U1674 (N_1674,N_1271,N_1359);
and U1675 (N_1675,N_1157,N_940);
nor U1676 (N_1676,N_773,N_1408);
or U1677 (N_1677,N_918,N_845);
nand U1678 (N_1678,N_1418,N_1191);
and U1679 (N_1679,N_1308,N_797);
nor U1680 (N_1680,N_1196,N_1026);
nand U1681 (N_1681,N_1256,N_881);
nand U1682 (N_1682,N_1340,N_1386);
nor U1683 (N_1683,N_980,N_1328);
nand U1684 (N_1684,N_942,N_826);
or U1685 (N_1685,N_912,N_1415);
and U1686 (N_1686,N_1142,N_1086);
nand U1687 (N_1687,N_1228,N_1485);
nand U1688 (N_1688,N_971,N_1141);
nor U1689 (N_1689,N_1410,N_764);
nand U1690 (N_1690,N_994,N_1161);
and U1691 (N_1691,N_1393,N_1321);
nand U1692 (N_1692,N_1178,N_999);
nand U1693 (N_1693,N_1494,N_1149);
nand U1694 (N_1694,N_955,N_1289);
and U1695 (N_1695,N_837,N_1350);
or U1696 (N_1696,N_1433,N_1204);
xor U1697 (N_1697,N_1460,N_769);
and U1698 (N_1698,N_1027,N_794);
or U1699 (N_1699,N_890,N_958);
or U1700 (N_1700,N_953,N_1006);
or U1701 (N_1701,N_1380,N_927);
nand U1702 (N_1702,N_1369,N_1284);
nor U1703 (N_1703,N_1206,N_894);
nor U1704 (N_1704,N_1262,N_1356);
or U1705 (N_1705,N_866,N_768);
nand U1706 (N_1706,N_872,N_1170);
nor U1707 (N_1707,N_1277,N_1058);
xor U1708 (N_1708,N_1258,N_983);
nor U1709 (N_1709,N_1017,N_1306);
and U1710 (N_1710,N_1416,N_1250);
and U1711 (N_1711,N_1176,N_1248);
or U1712 (N_1712,N_1098,N_812);
nand U1713 (N_1713,N_1422,N_1215);
and U1714 (N_1714,N_1272,N_1400);
nand U1715 (N_1715,N_804,N_884);
or U1716 (N_1716,N_1484,N_985);
and U1717 (N_1717,N_1287,N_1154);
or U1718 (N_1718,N_1219,N_956);
nor U1719 (N_1719,N_1032,N_1233);
and U1720 (N_1720,N_771,N_1134);
or U1721 (N_1721,N_1120,N_1440);
nor U1722 (N_1722,N_1370,N_1077);
nand U1723 (N_1723,N_1323,N_1034);
and U1724 (N_1724,N_1382,N_1022);
nand U1725 (N_1725,N_876,N_1002);
nor U1726 (N_1726,N_1035,N_775);
or U1727 (N_1727,N_1294,N_1355);
nand U1728 (N_1728,N_1150,N_1118);
and U1729 (N_1729,N_1493,N_842);
nor U1730 (N_1730,N_1373,N_1189);
xor U1731 (N_1731,N_1169,N_1498);
nor U1732 (N_1732,N_925,N_1345);
and U1733 (N_1733,N_1457,N_1363);
nand U1734 (N_1734,N_1435,N_1217);
nor U1735 (N_1735,N_867,N_1326);
and U1736 (N_1736,N_1282,N_1218);
xor U1737 (N_1737,N_896,N_1405);
xnor U1738 (N_1738,N_832,N_920);
nor U1739 (N_1739,N_1292,N_1487);
nor U1740 (N_1740,N_1419,N_1430);
and U1741 (N_1741,N_1060,N_858);
nand U1742 (N_1742,N_1130,N_982);
or U1743 (N_1743,N_852,N_1159);
or U1744 (N_1744,N_860,N_1456);
nor U1745 (N_1745,N_784,N_873);
nand U1746 (N_1746,N_1237,N_1296);
nand U1747 (N_1747,N_992,N_1455);
xor U1748 (N_1748,N_1059,N_1279);
or U1749 (N_1749,N_778,N_954);
or U1750 (N_1750,N_932,N_1168);
and U1751 (N_1751,N_1371,N_1341);
or U1752 (N_1752,N_1243,N_1381);
nor U1753 (N_1753,N_1462,N_924);
or U1754 (N_1754,N_1038,N_1100);
and U1755 (N_1755,N_1268,N_1140);
xor U1756 (N_1756,N_1343,N_1247);
nand U1757 (N_1757,N_1165,N_1094);
nand U1758 (N_1758,N_937,N_815);
or U1759 (N_1759,N_1223,N_1171);
or U1760 (N_1760,N_1441,N_1108);
and U1761 (N_1761,N_1128,N_783);
nand U1762 (N_1762,N_1269,N_1010);
and U1763 (N_1763,N_1202,N_934);
and U1764 (N_1764,N_1085,N_829);
nor U1765 (N_1765,N_921,N_793);
nor U1766 (N_1766,N_975,N_1244);
nor U1767 (N_1767,N_1238,N_1111);
and U1768 (N_1768,N_1055,N_1096);
or U1769 (N_1769,N_946,N_855);
nor U1770 (N_1770,N_913,N_1251);
or U1771 (N_1771,N_1327,N_1483);
or U1772 (N_1772,N_1352,N_1333);
and U1773 (N_1773,N_1164,N_1307);
xor U1774 (N_1774,N_1266,N_952);
nor U1775 (N_1775,N_923,N_1042);
nor U1776 (N_1776,N_1226,N_796);
nand U1777 (N_1777,N_1126,N_807);
or U1778 (N_1778,N_818,N_1188);
and U1779 (N_1779,N_973,N_1212);
and U1780 (N_1780,N_901,N_1222);
nor U1781 (N_1781,N_1469,N_1231);
nand U1782 (N_1782,N_1395,N_777);
or U1783 (N_1783,N_1288,N_922);
xor U1784 (N_1784,N_1116,N_1310);
nor U1785 (N_1785,N_806,N_933);
and U1786 (N_1786,N_1110,N_1175);
nor U1787 (N_1787,N_1263,N_1014);
xor U1788 (N_1788,N_1254,N_1309);
or U1789 (N_1789,N_1025,N_1319);
nor U1790 (N_1790,N_836,N_1013);
nand U1791 (N_1791,N_889,N_1133);
nand U1792 (N_1792,N_1478,N_825);
nand U1793 (N_1793,N_755,N_1466);
nor U1794 (N_1794,N_1402,N_1451);
or U1795 (N_1795,N_840,N_1023);
and U1796 (N_1796,N_1162,N_843);
and U1797 (N_1797,N_963,N_1482);
nand U1798 (N_1798,N_1414,N_903);
nor U1799 (N_1799,N_1143,N_1364);
and U1800 (N_1800,N_945,N_1155);
and U1801 (N_1801,N_753,N_1338);
nor U1802 (N_1802,N_862,N_871);
nor U1803 (N_1803,N_960,N_1105);
xor U1804 (N_1804,N_785,N_966);
nand U1805 (N_1805,N_1474,N_1246);
nor U1806 (N_1806,N_1106,N_1446);
nand U1807 (N_1807,N_1093,N_750);
or U1808 (N_1808,N_864,N_841);
and U1809 (N_1809,N_1087,N_1145);
and U1810 (N_1810,N_1225,N_1252);
and U1811 (N_1811,N_917,N_1062);
nand U1812 (N_1812,N_850,N_1095);
nand U1813 (N_1813,N_1453,N_774);
or U1814 (N_1814,N_835,N_1201);
or U1815 (N_1815,N_1000,N_935);
nor U1816 (N_1816,N_1097,N_786);
nand U1817 (N_1817,N_1468,N_1261);
nor U1818 (N_1818,N_1264,N_757);
or U1819 (N_1819,N_1135,N_996);
nor U1820 (N_1820,N_763,N_1069);
nor U1821 (N_1821,N_801,N_854);
and U1822 (N_1822,N_1068,N_1348);
nand U1823 (N_1823,N_943,N_1492);
nor U1824 (N_1824,N_856,N_886);
or U1825 (N_1825,N_1311,N_1442);
nor U1826 (N_1826,N_1362,N_1200);
nor U1827 (N_1827,N_1398,N_1109);
xor U1828 (N_1828,N_1280,N_1064);
and U1829 (N_1829,N_1412,N_1346);
nor U1830 (N_1830,N_849,N_1342);
and U1831 (N_1831,N_1156,N_1066);
nand U1832 (N_1832,N_1316,N_1426);
nor U1833 (N_1833,N_859,N_1107);
nor U1834 (N_1834,N_1461,N_1112);
nand U1835 (N_1835,N_929,N_1167);
nor U1836 (N_1836,N_1136,N_1406);
nand U1837 (N_1837,N_1479,N_1313);
nor U1838 (N_1838,N_1431,N_1166);
nor U1839 (N_1839,N_1184,N_844);
and U1840 (N_1840,N_1351,N_939);
nor U1841 (N_1841,N_1372,N_1471);
nand U1842 (N_1842,N_1454,N_947);
nor U1843 (N_1843,N_1349,N_1071);
nor U1844 (N_1844,N_907,N_1259);
and U1845 (N_1845,N_1336,N_1437);
and U1846 (N_1846,N_967,N_910);
nor U1847 (N_1847,N_847,N_1213);
xor U1848 (N_1848,N_1079,N_792);
nor U1849 (N_1849,N_1054,N_759);
nand U1850 (N_1850,N_1423,N_760);
nor U1851 (N_1851,N_1438,N_1449);
and U1852 (N_1852,N_938,N_986);
or U1853 (N_1853,N_805,N_861);
and U1854 (N_1854,N_1385,N_795);
and U1855 (N_1855,N_868,N_1082);
xnor U1856 (N_1856,N_1315,N_1070);
or U1857 (N_1857,N_1432,N_828);
nor U1858 (N_1858,N_1302,N_1163);
nor U1859 (N_1859,N_1403,N_1399);
nand U1860 (N_1860,N_1207,N_1278);
and U1861 (N_1861,N_752,N_810);
nand U1862 (N_1862,N_846,N_787);
xor U1863 (N_1863,N_899,N_791);
and U1864 (N_1864,N_853,N_751);
nor U1865 (N_1865,N_767,N_1353);
nand U1866 (N_1866,N_1276,N_1265);
nand U1867 (N_1867,N_1236,N_1153);
and U1868 (N_1868,N_1388,N_1283);
xor U1869 (N_1869,N_1033,N_936);
or U1870 (N_1870,N_1459,N_1172);
or U1871 (N_1871,N_1472,N_863);
nand U1872 (N_1872,N_1099,N_1293);
nor U1873 (N_1873,N_1332,N_1160);
nand U1874 (N_1874,N_1221,N_1452);
and U1875 (N_1875,N_1064,N_1068);
nand U1876 (N_1876,N_1080,N_970);
nor U1877 (N_1877,N_1406,N_1427);
and U1878 (N_1878,N_1095,N_982);
or U1879 (N_1879,N_809,N_977);
or U1880 (N_1880,N_910,N_882);
nor U1881 (N_1881,N_783,N_1103);
nor U1882 (N_1882,N_1225,N_1016);
or U1883 (N_1883,N_1012,N_1157);
or U1884 (N_1884,N_1407,N_782);
nand U1885 (N_1885,N_1363,N_883);
and U1886 (N_1886,N_896,N_1349);
nand U1887 (N_1887,N_1012,N_990);
xnor U1888 (N_1888,N_1080,N_1277);
xor U1889 (N_1889,N_817,N_847);
nand U1890 (N_1890,N_1181,N_1150);
nor U1891 (N_1891,N_1478,N_1279);
and U1892 (N_1892,N_973,N_1150);
or U1893 (N_1893,N_1213,N_1333);
and U1894 (N_1894,N_1059,N_1283);
nand U1895 (N_1895,N_976,N_1379);
xnor U1896 (N_1896,N_829,N_1215);
nand U1897 (N_1897,N_865,N_1038);
xnor U1898 (N_1898,N_1293,N_751);
nand U1899 (N_1899,N_1119,N_778);
nor U1900 (N_1900,N_1054,N_834);
or U1901 (N_1901,N_1340,N_1280);
xor U1902 (N_1902,N_796,N_977);
nand U1903 (N_1903,N_1393,N_1007);
nor U1904 (N_1904,N_964,N_1174);
or U1905 (N_1905,N_1310,N_935);
or U1906 (N_1906,N_1313,N_938);
and U1907 (N_1907,N_1145,N_864);
nand U1908 (N_1908,N_809,N_833);
nand U1909 (N_1909,N_1428,N_771);
and U1910 (N_1910,N_1343,N_1324);
and U1911 (N_1911,N_1365,N_1060);
or U1912 (N_1912,N_956,N_1371);
and U1913 (N_1913,N_1377,N_1042);
nand U1914 (N_1914,N_1392,N_1180);
or U1915 (N_1915,N_1164,N_1038);
xnor U1916 (N_1916,N_1290,N_1027);
nor U1917 (N_1917,N_899,N_867);
nand U1918 (N_1918,N_858,N_1422);
nand U1919 (N_1919,N_1318,N_774);
nor U1920 (N_1920,N_984,N_933);
xor U1921 (N_1921,N_975,N_1443);
nor U1922 (N_1922,N_881,N_1319);
and U1923 (N_1923,N_1045,N_1140);
xnor U1924 (N_1924,N_1419,N_1315);
and U1925 (N_1925,N_799,N_1153);
nand U1926 (N_1926,N_1471,N_1311);
or U1927 (N_1927,N_897,N_875);
or U1928 (N_1928,N_1013,N_862);
and U1929 (N_1929,N_1471,N_799);
and U1930 (N_1930,N_1476,N_979);
nor U1931 (N_1931,N_1115,N_1330);
and U1932 (N_1932,N_1157,N_1098);
or U1933 (N_1933,N_1459,N_824);
nand U1934 (N_1934,N_934,N_1386);
and U1935 (N_1935,N_1347,N_1249);
and U1936 (N_1936,N_1185,N_1238);
or U1937 (N_1937,N_1370,N_1414);
nand U1938 (N_1938,N_1191,N_778);
or U1939 (N_1939,N_1006,N_920);
nand U1940 (N_1940,N_813,N_840);
and U1941 (N_1941,N_1355,N_1166);
or U1942 (N_1942,N_772,N_1084);
and U1943 (N_1943,N_1078,N_852);
nor U1944 (N_1944,N_1076,N_844);
nand U1945 (N_1945,N_1221,N_1033);
nand U1946 (N_1946,N_1393,N_1289);
nand U1947 (N_1947,N_883,N_1285);
and U1948 (N_1948,N_1070,N_1422);
or U1949 (N_1949,N_1007,N_1082);
or U1950 (N_1950,N_1356,N_1232);
nand U1951 (N_1951,N_1169,N_997);
nor U1952 (N_1952,N_1071,N_1422);
nand U1953 (N_1953,N_1172,N_914);
and U1954 (N_1954,N_867,N_1201);
or U1955 (N_1955,N_1460,N_857);
nor U1956 (N_1956,N_896,N_1062);
nand U1957 (N_1957,N_1058,N_1103);
and U1958 (N_1958,N_775,N_1066);
and U1959 (N_1959,N_1182,N_1165);
or U1960 (N_1960,N_1090,N_856);
and U1961 (N_1961,N_1425,N_1253);
and U1962 (N_1962,N_878,N_770);
nand U1963 (N_1963,N_1005,N_1213);
nand U1964 (N_1964,N_1469,N_1240);
xor U1965 (N_1965,N_1357,N_1111);
nand U1966 (N_1966,N_913,N_925);
nor U1967 (N_1967,N_900,N_912);
and U1968 (N_1968,N_902,N_1342);
or U1969 (N_1969,N_786,N_921);
nand U1970 (N_1970,N_1469,N_969);
and U1971 (N_1971,N_1094,N_1308);
xor U1972 (N_1972,N_1315,N_1371);
or U1973 (N_1973,N_1492,N_801);
xnor U1974 (N_1974,N_784,N_1106);
nor U1975 (N_1975,N_1041,N_997);
and U1976 (N_1976,N_1481,N_1314);
or U1977 (N_1977,N_960,N_1028);
nor U1978 (N_1978,N_1191,N_824);
or U1979 (N_1979,N_1041,N_1285);
or U1980 (N_1980,N_840,N_965);
nand U1981 (N_1981,N_1340,N_1293);
nand U1982 (N_1982,N_1134,N_1010);
or U1983 (N_1983,N_829,N_834);
nor U1984 (N_1984,N_762,N_824);
nor U1985 (N_1985,N_1277,N_1415);
nor U1986 (N_1986,N_1421,N_1059);
or U1987 (N_1987,N_1244,N_1153);
nor U1988 (N_1988,N_1374,N_1406);
and U1989 (N_1989,N_1387,N_998);
or U1990 (N_1990,N_958,N_1373);
or U1991 (N_1991,N_860,N_1350);
nand U1992 (N_1992,N_1160,N_1461);
or U1993 (N_1993,N_1286,N_898);
nor U1994 (N_1994,N_967,N_1290);
or U1995 (N_1995,N_1191,N_1412);
xor U1996 (N_1996,N_1366,N_1355);
xor U1997 (N_1997,N_914,N_1480);
or U1998 (N_1998,N_888,N_1302);
nand U1999 (N_1999,N_1342,N_914);
or U2000 (N_2000,N_1302,N_1406);
nand U2001 (N_2001,N_788,N_1148);
and U2002 (N_2002,N_1382,N_923);
nand U2003 (N_2003,N_810,N_1213);
nor U2004 (N_2004,N_1289,N_1491);
and U2005 (N_2005,N_838,N_1485);
nor U2006 (N_2006,N_879,N_932);
or U2007 (N_2007,N_1043,N_1031);
nand U2008 (N_2008,N_1308,N_974);
nand U2009 (N_2009,N_895,N_1197);
nand U2010 (N_2010,N_1248,N_1035);
and U2011 (N_2011,N_1158,N_985);
or U2012 (N_2012,N_1107,N_904);
nand U2013 (N_2013,N_841,N_1492);
or U2014 (N_2014,N_1498,N_789);
and U2015 (N_2015,N_1383,N_800);
and U2016 (N_2016,N_847,N_1377);
nor U2017 (N_2017,N_839,N_1434);
nor U2018 (N_2018,N_829,N_1115);
or U2019 (N_2019,N_807,N_951);
nand U2020 (N_2020,N_1195,N_1087);
nor U2021 (N_2021,N_916,N_1109);
and U2022 (N_2022,N_816,N_1297);
and U2023 (N_2023,N_1439,N_1165);
or U2024 (N_2024,N_1408,N_982);
nand U2025 (N_2025,N_800,N_1413);
nand U2026 (N_2026,N_1011,N_986);
xnor U2027 (N_2027,N_857,N_1223);
or U2028 (N_2028,N_1343,N_1034);
nor U2029 (N_2029,N_999,N_1216);
or U2030 (N_2030,N_1384,N_1389);
and U2031 (N_2031,N_1309,N_771);
nor U2032 (N_2032,N_860,N_1389);
nand U2033 (N_2033,N_984,N_1263);
xnor U2034 (N_2034,N_1333,N_1058);
nand U2035 (N_2035,N_1427,N_1386);
or U2036 (N_2036,N_1055,N_1165);
nand U2037 (N_2037,N_1157,N_959);
and U2038 (N_2038,N_996,N_1124);
nand U2039 (N_2039,N_794,N_901);
xnor U2040 (N_2040,N_1261,N_841);
and U2041 (N_2041,N_1444,N_1306);
or U2042 (N_2042,N_1071,N_1460);
nand U2043 (N_2043,N_1198,N_1128);
nor U2044 (N_2044,N_1183,N_972);
nor U2045 (N_2045,N_1353,N_1082);
xor U2046 (N_2046,N_1360,N_988);
or U2047 (N_2047,N_863,N_1417);
xnor U2048 (N_2048,N_1341,N_1327);
nor U2049 (N_2049,N_1242,N_851);
xor U2050 (N_2050,N_1349,N_816);
nor U2051 (N_2051,N_1351,N_979);
nand U2052 (N_2052,N_971,N_765);
or U2053 (N_2053,N_996,N_1175);
nand U2054 (N_2054,N_882,N_1215);
nor U2055 (N_2055,N_848,N_805);
and U2056 (N_2056,N_1093,N_892);
and U2057 (N_2057,N_1272,N_841);
or U2058 (N_2058,N_1224,N_1289);
and U2059 (N_2059,N_1247,N_1257);
nor U2060 (N_2060,N_1039,N_864);
nand U2061 (N_2061,N_1326,N_942);
nor U2062 (N_2062,N_1282,N_863);
xor U2063 (N_2063,N_1002,N_1140);
or U2064 (N_2064,N_1383,N_777);
nand U2065 (N_2065,N_1419,N_899);
nand U2066 (N_2066,N_1393,N_1189);
nor U2067 (N_2067,N_1283,N_1046);
and U2068 (N_2068,N_1242,N_1174);
nor U2069 (N_2069,N_1203,N_772);
and U2070 (N_2070,N_1418,N_1002);
or U2071 (N_2071,N_1294,N_1237);
or U2072 (N_2072,N_860,N_1133);
or U2073 (N_2073,N_1120,N_791);
nor U2074 (N_2074,N_1104,N_1329);
nand U2075 (N_2075,N_1414,N_775);
nand U2076 (N_2076,N_1230,N_1478);
and U2077 (N_2077,N_1132,N_1226);
nand U2078 (N_2078,N_1264,N_1306);
or U2079 (N_2079,N_1415,N_1153);
and U2080 (N_2080,N_1487,N_1255);
nor U2081 (N_2081,N_1315,N_1488);
and U2082 (N_2082,N_1016,N_933);
or U2083 (N_2083,N_1333,N_1139);
and U2084 (N_2084,N_1378,N_1203);
xor U2085 (N_2085,N_983,N_1243);
or U2086 (N_2086,N_1285,N_1014);
nand U2087 (N_2087,N_1305,N_1344);
xor U2088 (N_2088,N_778,N_898);
nand U2089 (N_2089,N_1133,N_946);
nand U2090 (N_2090,N_1401,N_766);
xor U2091 (N_2091,N_1388,N_1276);
xnor U2092 (N_2092,N_989,N_1463);
nand U2093 (N_2093,N_869,N_1483);
nand U2094 (N_2094,N_906,N_1134);
and U2095 (N_2095,N_831,N_924);
or U2096 (N_2096,N_1152,N_965);
nor U2097 (N_2097,N_821,N_1032);
nor U2098 (N_2098,N_1217,N_889);
xnor U2099 (N_2099,N_1300,N_968);
nand U2100 (N_2100,N_978,N_1416);
nor U2101 (N_2101,N_954,N_854);
and U2102 (N_2102,N_1207,N_1386);
and U2103 (N_2103,N_1168,N_839);
or U2104 (N_2104,N_1154,N_1324);
xnor U2105 (N_2105,N_1198,N_1471);
and U2106 (N_2106,N_1063,N_1189);
or U2107 (N_2107,N_1311,N_1243);
and U2108 (N_2108,N_1109,N_864);
and U2109 (N_2109,N_928,N_794);
nor U2110 (N_2110,N_844,N_1089);
or U2111 (N_2111,N_934,N_1042);
nor U2112 (N_2112,N_1194,N_1101);
nand U2113 (N_2113,N_1485,N_986);
or U2114 (N_2114,N_1008,N_1387);
and U2115 (N_2115,N_977,N_1330);
and U2116 (N_2116,N_863,N_975);
or U2117 (N_2117,N_938,N_967);
nand U2118 (N_2118,N_1050,N_1284);
or U2119 (N_2119,N_1271,N_1446);
and U2120 (N_2120,N_1102,N_1447);
and U2121 (N_2121,N_884,N_960);
nand U2122 (N_2122,N_1339,N_1354);
xor U2123 (N_2123,N_1435,N_1362);
and U2124 (N_2124,N_904,N_1414);
nand U2125 (N_2125,N_1475,N_808);
nand U2126 (N_2126,N_1099,N_1285);
nor U2127 (N_2127,N_962,N_1179);
nand U2128 (N_2128,N_1069,N_1379);
nand U2129 (N_2129,N_1394,N_1265);
and U2130 (N_2130,N_983,N_1262);
or U2131 (N_2131,N_1367,N_1259);
xnor U2132 (N_2132,N_854,N_1083);
nand U2133 (N_2133,N_1485,N_1366);
or U2134 (N_2134,N_1132,N_768);
and U2135 (N_2135,N_829,N_1387);
and U2136 (N_2136,N_895,N_1321);
or U2137 (N_2137,N_1309,N_1446);
or U2138 (N_2138,N_1497,N_990);
and U2139 (N_2139,N_949,N_1207);
nand U2140 (N_2140,N_1113,N_1457);
nand U2141 (N_2141,N_1388,N_1476);
or U2142 (N_2142,N_1049,N_1218);
or U2143 (N_2143,N_934,N_796);
xor U2144 (N_2144,N_1099,N_1189);
nor U2145 (N_2145,N_985,N_849);
nor U2146 (N_2146,N_787,N_1074);
or U2147 (N_2147,N_1264,N_1316);
or U2148 (N_2148,N_1411,N_1080);
nand U2149 (N_2149,N_1118,N_962);
nand U2150 (N_2150,N_1439,N_1470);
nand U2151 (N_2151,N_954,N_883);
nor U2152 (N_2152,N_1111,N_1171);
and U2153 (N_2153,N_1383,N_1072);
or U2154 (N_2154,N_794,N_1041);
and U2155 (N_2155,N_841,N_1140);
or U2156 (N_2156,N_982,N_1462);
nand U2157 (N_2157,N_1455,N_1000);
nand U2158 (N_2158,N_917,N_1359);
or U2159 (N_2159,N_1247,N_1046);
and U2160 (N_2160,N_992,N_1425);
nor U2161 (N_2161,N_1354,N_1081);
xor U2162 (N_2162,N_833,N_1488);
nor U2163 (N_2163,N_1136,N_1120);
or U2164 (N_2164,N_924,N_1164);
nor U2165 (N_2165,N_1314,N_988);
and U2166 (N_2166,N_1355,N_1411);
and U2167 (N_2167,N_1083,N_1182);
nor U2168 (N_2168,N_976,N_1330);
and U2169 (N_2169,N_782,N_1178);
or U2170 (N_2170,N_1137,N_857);
and U2171 (N_2171,N_1496,N_1218);
and U2172 (N_2172,N_1362,N_1069);
nand U2173 (N_2173,N_1018,N_979);
and U2174 (N_2174,N_861,N_1441);
xnor U2175 (N_2175,N_989,N_771);
xnor U2176 (N_2176,N_1217,N_1349);
nand U2177 (N_2177,N_1116,N_874);
xnor U2178 (N_2178,N_1061,N_1432);
nor U2179 (N_2179,N_1046,N_1045);
xnor U2180 (N_2180,N_1171,N_891);
or U2181 (N_2181,N_1285,N_1323);
and U2182 (N_2182,N_1259,N_986);
and U2183 (N_2183,N_787,N_1254);
nor U2184 (N_2184,N_1379,N_1002);
nand U2185 (N_2185,N_1042,N_1306);
nor U2186 (N_2186,N_1023,N_1274);
and U2187 (N_2187,N_932,N_810);
or U2188 (N_2188,N_1020,N_1073);
nor U2189 (N_2189,N_1115,N_813);
nand U2190 (N_2190,N_1358,N_1254);
nand U2191 (N_2191,N_1097,N_879);
or U2192 (N_2192,N_1207,N_1076);
nand U2193 (N_2193,N_891,N_1472);
nor U2194 (N_2194,N_1048,N_910);
or U2195 (N_2195,N_1148,N_1173);
or U2196 (N_2196,N_1108,N_826);
nor U2197 (N_2197,N_1324,N_1066);
nand U2198 (N_2198,N_1330,N_1147);
and U2199 (N_2199,N_819,N_1454);
or U2200 (N_2200,N_1284,N_831);
and U2201 (N_2201,N_1163,N_815);
nor U2202 (N_2202,N_943,N_1344);
xor U2203 (N_2203,N_1324,N_880);
nor U2204 (N_2204,N_1488,N_792);
and U2205 (N_2205,N_1089,N_1308);
or U2206 (N_2206,N_898,N_888);
and U2207 (N_2207,N_1059,N_1472);
nand U2208 (N_2208,N_1164,N_960);
nor U2209 (N_2209,N_1256,N_952);
nor U2210 (N_2210,N_794,N_1150);
nor U2211 (N_2211,N_822,N_1088);
nand U2212 (N_2212,N_1222,N_1487);
and U2213 (N_2213,N_1320,N_1173);
or U2214 (N_2214,N_1367,N_1402);
and U2215 (N_2215,N_974,N_1121);
or U2216 (N_2216,N_849,N_831);
nor U2217 (N_2217,N_981,N_1038);
or U2218 (N_2218,N_1051,N_1095);
or U2219 (N_2219,N_902,N_1196);
nor U2220 (N_2220,N_1325,N_919);
and U2221 (N_2221,N_1397,N_1342);
xor U2222 (N_2222,N_1170,N_1411);
and U2223 (N_2223,N_1494,N_1366);
or U2224 (N_2224,N_1057,N_881);
xnor U2225 (N_2225,N_945,N_1328);
or U2226 (N_2226,N_893,N_1345);
nand U2227 (N_2227,N_1023,N_1394);
or U2228 (N_2228,N_1496,N_1090);
and U2229 (N_2229,N_1352,N_1334);
nor U2230 (N_2230,N_1123,N_925);
nor U2231 (N_2231,N_1100,N_1294);
or U2232 (N_2232,N_1128,N_1408);
and U2233 (N_2233,N_1234,N_1191);
nor U2234 (N_2234,N_1251,N_1381);
and U2235 (N_2235,N_1242,N_1070);
or U2236 (N_2236,N_762,N_983);
or U2237 (N_2237,N_1059,N_979);
nand U2238 (N_2238,N_1154,N_1230);
xor U2239 (N_2239,N_1012,N_1126);
or U2240 (N_2240,N_1359,N_1087);
or U2241 (N_2241,N_1270,N_862);
nand U2242 (N_2242,N_967,N_981);
and U2243 (N_2243,N_824,N_985);
nand U2244 (N_2244,N_1471,N_1084);
or U2245 (N_2245,N_757,N_1277);
and U2246 (N_2246,N_1192,N_996);
nand U2247 (N_2247,N_1251,N_832);
nor U2248 (N_2248,N_1371,N_977);
or U2249 (N_2249,N_1474,N_1353);
or U2250 (N_2250,N_2143,N_1627);
and U2251 (N_2251,N_1818,N_1588);
and U2252 (N_2252,N_1826,N_1608);
nor U2253 (N_2253,N_1925,N_1693);
or U2254 (N_2254,N_1986,N_1744);
nand U2255 (N_2255,N_1885,N_1918);
nor U2256 (N_2256,N_1539,N_1679);
or U2257 (N_2257,N_1635,N_1805);
nor U2258 (N_2258,N_1771,N_2171);
nand U2259 (N_2259,N_1565,N_1908);
nor U2260 (N_2260,N_1971,N_2185);
and U2261 (N_2261,N_2050,N_1589);
and U2262 (N_2262,N_1756,N_1522);
and U2263 (N_2263,N_1999,N_1894);
and U2264 (N_2264,N_1515,N_2152);
and U2265 (N_2265,N_2103,N_1776);
and U2266 (N_2266,N_1827,N_2058);
or U2267 (N_2267,N_2156,N_2230);
nor U2268 (N_2268,N_1692,N_1513);
nand U2269 (N_2269,N_1833,N_1912);
nand U2270 (N_2270,N_2003,N_2219);
xnor U2271 (N_2271,N_1860,N_1969);
nor U2272 (N_2272,N_1795,N_1648);
and U2273 (N_2273,N_1931,N_1753);
or U2274 (N_2274,N_2194,N_2061);
nand U2275 (N_2275,N_2119,N_1591);
nand U2276 (N_2276,N_1667,N_1766);
or U2277 (N_2277,N_2072,N_2024);
and U2278 (N_2278,N_1834,N_2111);
and U2279 (N_2279,N_2182,N_1717);
nand U2280 (N_2280,N_1720,N_1637);
nor U2281 (N_2281,N_1767,N_1956);
nand U2282 (N_2282,N_1857,N_1675);
nor U2283 (N_2283,N_1965,N_2064);
and U2284 (N_2284,N_1629,N_1760);
or U2285 (N_2285,N_1748,N_2159);
nor U2286 (N_2286,N_2225,N_1628);
xnor U2287 (N_2287,N_1829,N_2155);
and U2288 (N_2288,N_2224,N_1774);
nand U2289 (N_2289,N_2221,N_2222);
or U2290 (N_2290,N_2026,N_1689);
nand U2291 (N_2291,N_2184,N_2193);
nand U2292 (N_2292,N_1684,N_1509);
and U2293 (N_2293,N_1798,N_2117);
or U2294 (N_2294,N_1968,N_1558);
and U2295 (N_2295,N_1940,N_1561);
and U2296 (N_2296,N_1875,N_1524);
xnor U2297 (N_2297,N_1998,N_2084);
nand U2298 (N_2298,N_1987,N_1507);
and U2299 (N_2299,N_2128,N_1546);
or U2300 (N_2300,N_1709,N_1822);
or U2301 (N_2301,N_1523,N_2132);
and U2302 (N_2302,N_2076,N_2039);
xnor U2303 (N_2303,N_1884,N_2067);
or U2304 (N_2304,N_1859,N_1897);
nand U2305 (N_2305,N_1879,N_1994);
nand U2306 (N_2306,N_2075,N_2053);
and U2307 (N_2307,N_2055,N_1970);
nand U2308 (N_2308,N_2210,N_1701);
or U2309 (N_2309,N_1682,N_1806);
xnor U2310 (N_2310,N_2100,N_1581);
or U2311 (N_2311,N_1514,N_1520);
nand U2312 (N_2312,N_1848,N_1735);
nor U2313 (N_2313,N_1945,N_1721);
or U2314 (N_2314,N_1587,N_2052);
or U2315 (N_2315,N_2044,N_1584);
nor U2316 (N_2316,N_2195,N_2120);
and U2317 (N_2317,N_1896,N_1888);
nand U2318 (N_2318,N_1845,N_1775);
and U2319 (N_2319,N_2168,N_1611);
and U2320 (N_2320,N_1510,N_1892);
nand U2321 (N_2321,N_2147,N_1804);
nor U2322 (N_2322,N_1976,N_1758);
nand U2323 (N_2323,N_1670,N_1846);
and U2324 (N_2324,N_2022,N_2211);
or U2325 (N_2325,N_2089,N_1813);
nand U2326 (N_2326,N_2165,N_1501);
or U2327 (N_2327,N_2043,N_2137);
and U2328 (N_2328,N_2246,N_1828);
nor U2329 (N_2329,N_2006,N_1538);
or U2330 (N_2330,N_2231,N_1923);
or U2331 (N_2331,N_1697,N_2088);
xnor U2332 (N_2332,N_2037,N_2167);
and U2333 (N_2333,N_1723,N_1592);
and U2334 (N_2334,N_1855,N_1521);
and U2335 (N_2335,N_1935,N_1734);
xor U2336 (N_2336,N_1853,N_1733);
and U2337 (N_2337,N_1527,N_2032);
nor U2338 (N_2338,N_2106,N_2150);
and U2339 (N_2339,N_1893,N_1713);
or U2340 (N_2340,N_1762,N_2201);
nand U2341 (N_2341,N_2019,N_1719);
or U2342 (N_2342,N_1851,N_1618);
nand U2343 (N_2343,N_1516,N_1568);
nand U2344 (N_2344,N_1850,N_1506);
nand U2345 (N_2345,N_2093,N_2226);
and U2346 (N_2346,N_1549,N_1712);
nor U2347 (N_2347,N_1727,N_1955);
and U2348 (N_2348,N_1996,N_1557);
and U2349 (N_2349,N_2035,N_2070);
nand U2350 (N_2350,N_1903,N_2094);
and U2351 (N_2351,N_2216,N_1847);
and U2352 (N_2352,N_2213,N_1631);
or U2353 (N_2353,N_1708,N_2153);
xnor U2354 (N_2354,N_1570,N_1832);
and U2355 (N_2355,N_1674,N_1949);
nand U2356 (N_2356,N_1948,N_1728);
nor U2357 (N_2357,N_1671,N_1785);
nor U2358 (N_2358,N_1547,N_1541);
nor U2359 (N_2359,N_1505,N_1639);
xor U2360 (N_2360,N_1579,N_1919);
and U2361 (N_2361,N_1898,N_1901);
or U2362 (N_2362,N_1606,N_2099);
nand U2363 (N_2363,N_1946,N_2177);
or U2364 (N_2364,N_1612,N_1783);
xnor U2365 (N_2365,N_1761,N_1982);
nor U2366 (N_2366,N_2059,N_2115);
nand U2367 (N_2367,N_1820,N_1673);
nand U2368 (N_2368,N_1747,N_1602);
or U2369 (N_2369,N_1800,N_2158);
or U2370 (N_2370,N_2004,N_1525);
nand U2371 (N_2371,N_2057,N_1502);
nand U2372 (N_2372,N_1809,N_2002);
or U2373 (N_2373,N_1714,N_1984);
nand U2374 (N_2374,N_2172,N_2081);
xnor U2375 (N_2375,N_1656,N_1992);
nor U2376 (N_2376,N_1556,N_1622);
and U2377 (N_2377,N_1802,N_2001);
nor U2378 (N_2378,N_1858,N_1930);
or U2379 (N_2379,N_2060,N_1722);
and U2380 (N_2380,N_1595,N_1778);
nor U2381 (N_2381,N_2144,N_2233);
and U2382 (N_2382,N_2228,N_1927);
nand U2383 (N_2383,N_2105,N_1659);
or U2384 (N_2384,N_1967,N_2130);
nor U2385 (N_2385,N_1889,N_1989);
and U2386 (N_2386,N_1614,N_1812);
and U2387 (N_2387,N_1548,N_2097);
nand U2388 (N_2388,N_1545,N_2007);
xor U2389 (N_2389,N_1566,N_1890);
nand U2390 (N_2390,N_2197,N_2235);
xnor U2391 (N_2391,N_1921,N_1615);
and U2392 (N_2392,N_1696,N_1852);
and U2393 (N_2393,N_1621,N_1729);
nand U2394 (N_2394,N_2021,N_1958);
nor U2395 (N_2395,N_1594,N_1593);
nor U2396 (N_2396,N_1910,N_1691);
nand U2397 (N_2397,N_1640,N_1677);
or U2398 (N_2398,N_2175,N_2126);
nor U2399 (N_2399,N_2204,N_2247);
nor U2400 (N_2400,N_1687,N_1831);
nand U2401 (N_2401,N_1555,N_1873);
or U2402 (N_2402,N_1781,N_2123);
and U2403 (N_2403,N_1537,N_1928);
and U2404 (N_2404,N_2135,N_1601);
xor U2405 (N_2405,N_1862,N_2048);
and U2406 (N_2406,N_2096,N_2207);
or U2407 (N_2407,N_2218,N_2214);
and U2408 (N_2408,N_1634,N_2187);
xor U2409 (N_2409,N_1718,N_2133);
and U2410 (N_2410,N_1962,N_2078);
nand U2411 (N_2411,N_2149,N_1765);
xor U2412 (N_2412,N_1698,N_1799);
or U2413 (N_2413,N_2160,N_1796);
or U2414 (N_2414,N_1724,N_2178);
and U2415 (N_2415,N_2014,N_2095);
nor U2416 (N_2416,N_1768,N_2102);
nand U2417 (N_2417,N_1617,N_1934);
xor U2418 (N_2418,N_1926,N_1605);
or U2419 (N_2419,N_1500,N_2237);
or U2420 (N_2420,N_1743,N_1817);
nor U2421 (N_2421,N_2205,N_2011);
xnor U2422 (N_2422,N_1964,N_1835);
nor U2423 (N_2423,N_1902,N_2239);
xor U2424 (N_2424,N_1830,N_2206);
nand U2425 (N_2425,N_1844,N_1519);
and U2426 (N_2426,N_1562,N_1597);
or U2427 (N_2427,N_1534,N_2176);
and U2428 (N_2428,N_2173,N_1941);
nand U2429 (N_2429,N_1878,N_1609);
nand U2430 (N_2430,N_1808,N_2012);
or U2431 (N_2431,N_1825,N_1632);
nor U2432 (N_2432,N_1784,N_1993);
and U2433 (N_2433,N_1576,N_1567);
nand U2434 (N_2434,N_1624,N_2023);
nand U2435 (N_2435,N_1972,N_1690);
or U2436 (N_2436,N_2162,N_2065);
nor U2437 (N_2437,N_1867,N_1660);
or U2438 (N_2438,N_2101,N_1600);
nor U2439 (N_2439,N_2079,N_2045);
nor U2440 (N_2440,N_1819,N_1610);
and U2441 (N_2441,N_2074,N_1791);
and U2442 (N_2442,N_1988,N_1881);
nor U2443 (N_2443,N_1793,N_1957);
and U2444 (N_2444,N_1950,N_2116);
and U2445 (N_2445,N_1983,N_2217);
xor U2446 (N_2446,N_2046,N_1742);
xor U2447 (N_2447,N_1978,N_1598);
nand U2448 (N_2448,N_1954,N_1869);
and U2449 (N_2449,N_1536,N_1977);
xor U2450 (N_2450,N_2041,N_1990);
and U2451 (N_2451,N_1782,N_1552);
nand U2452 (N_2452,N_2009,N_1544);
nand U2453 (N_2453,N_1590,N_2245);
xor U2454 (N_2454,N_1870,N_1700);
nor U2455 (N_2455,N_1715,N_1877);
and U2456 (N_2456,N_2199,N_1961);
nor U2457 (N_2457,N_2179,N_2166);
nor U2458 (N_2458,N_1966,N_1563);
or U2459 (N_2459,N_2243,N_1653);
nor U2460 (N_2460,N_1790,N_2139);
or U2461 (N_2461,N_1650,N_2040);
xnor U2462 (N_2462,N_1779,N_2202);
or U2463 (N_2463,N_1574,N_1759);
nand U2464 (N_2464,N_1754,N_1705);
nand U2465 (N_2465,N_1803,N_1914);
or U2466 (N_2466,N_2203,N_1603);
nor U2467 (N_2467,N_1668,N_1749);
and U2468 (N_2468,N_1937,N_1751);
or U2469 (N_2469,N_1794,N_1939);
or U2470 (N_2470,N_1596,N_1572);
nor U2471 (N_2471,N_2073,N_2196);
and U2472 (N_2472,N_1543,N_1856);
nor U2473 (N_2473,N_2038,N_2118);
or U2474 (N_2474,N_1920,N_1681);
xor U2475 (N_2475,N_1787,N_2232);
or U2476 (N_2476,N_2062,N_2241);
or U2477 (N_2477,N_1985,N_1645);
nand U2478 (N_2478,N_1737,N_1676);
nor U2479 (N_2479,N_2170,N_1780);
nor U2480 (N_2480,N_2000,N_1854);
nor U2481 (N_2481,N_1849,N_1528);
nor U2482 (N_2482,N_1586,N_1625);
nor U2483 (N_2483,N_1883,N_1997);
nor U2484 (N_2484,N_2151,N_1953);
nor U2485 (N_2485,N_1732,N_1991);
nor U2486 (N_2486,N_1647,N_1944);
and U2487 (N_2487,N_2157,N_1731);
nand U2488 (N_2488,N_1633,N_2112);
nand U2489 (N_2489,N_1531,N_2161);
nand U2490 (N_2490,N_1569,N_1651);
or U2491 (N_2491,N_2140,N_2042);
nand U2492 (N_2492,N_1699,N_2181);
or U2493 (N_2493,N_1895,N_1932);
or U2494 (N_2494,N_2190,N_2107);
xor U2495 (N_2495,N_2015,N_1786);
nand U2496 (N_2496,N_1900,N_1707);
and U2497 (N_2497,N_1904,N_2227);
or U2498 (N_2498,N_1626,N_2141);
or U2499 (N_2499,N_1518,N_2028);
nand U2500 (N_2500,N_2234,N_1906);
xor U2501 (N_2501,N_2033,N_1642);
xor U2502 (N_2502,N_1613,N_2056);
nor U2503 (N_2503,N_2163,N_1535);
or U2504 (N_2504,N_1716,N_2136);
xor U2505 (N_2505,N_1909,N_1573);
and U2506 (N_2506,N_2122,N_1616);
nand U2507 (N_2507,N_2127,N_2129);
nand U2508 (N_2508,N_2198,N_1905);
and U2509 (N_2509,N_1980,N_1792);
or U2510 (N_2510,N_1788,N_2013);
and U2511 (N_2511,N_1951,N_1533);
nand U2512 (N_2512,N_2174,N_2082);
or U2513 (N_2513,N_2148,N_2240);
nor U2514 (N_2514,N_1503,N_2142);
nand U2515 (N_2515,N_1740,N_1532);
and U2516 (N_2516,N_2090,N_1745);
or U2517 (N_2517,N_1960,N_1599);
nand U2518 (N_2518,N_1880,N_1512);
nor U2519 (N_2519,N_1661,N_2191);
and U2520 (N_2520,N_2238,N_1652);
and U2521 (N_2521,N_1685,N_1553);
nor U2522 (N_2522,N_1876,N_2223);
nand U2523 (N_2523,N_1861,N_2029);
xnor U2524 (N_2524,N_2186,N_2063);
nor U2525 (N_2525,N_1739,N_1975);
nand U2526 (N_2526,N_1571,N_1665);
and U2527 (N_2527,N_1746,N_1511);
xnor U2528 (N_2528,N_1638,N_1672);
nor U2529 (N_2529,N_1836,N_1542);
nand U2530 (N_2530,N_2069,N_1736);
nand U2531 (N_2531,N_1959,N_1872);
nand U2532 (N_2532,N_1669,N_1702);
xor U2533 (N_2533,N_2083,N_1871);
and U2534 (N_2534,N_1947,N_1658);
or U2535 (N_2535,N_1620,N_2020);
or U2536 (N_2536,N_1868,N_2025);
nand U2537 (N_2537,N_1577,N_1560);
nor U2538 (N_2538,N_2010,N_2030);
xor U2539 (N_2539,N_1725,N_2027);
or U2540 (N_2540,N_1841,N_1824);
or U2541 (N_2541,N_1706,N_1839);
nor U2542 (N_2542,N_2086,N_1550);
nor U2543 (N_2543,N_1973,N_2180);
or U2544 (N_2544,N_2215,N_1936);
nand U2545 (N_2545,N_1630,N_1915);
or U2546 (N_2546,N_2209,N_1646);
or U2547 (N_2547,N_1559,N_1583);
and U2548 (N_2548,N_2054,N_1730);
and U2549 (N_2549,N_1695,N_2229);
nor U2550 (N_2550,N_2092,N_1666);
nor U2551 (N_2551,N_2110,N_1711);
nand U2552 (N_2552,N_1643,N_1763);
or U2553 (N_2553,N_2183,N_2047);
nand U2554 (N_2554,N_1604,N_1916);
and U2555 (N_2555,N_1526,N_1963);
or U2556 (N_2556,N_2036,N_2249);
nand U2557 (N_2557,N_1797,N_1755);
and U2558 (N_2558,N_1882,N_2248);
nor U2559 (N_2559,N_1694,N_1710);
nand U2560 (N_2560,N_2017,N_1952);
or U2561 (N_2561,N_1810,N_2236);
nor U2562 (N_2562,N_2145,N_1683);
xor U2563 (N_2563,N_1554,N_1911);
nand U2564 (N_2564,N_2049,N_1995);
xnor U2565 (N_2565,N_2124,N_2113);
and U2566 (N_2566,N_1821,N_1664);
or U2567 (N_2567,N_2031,N_1899);
and U2568 (N_2568,N_2131,N_2085);
or U2569 (N_2569,N_2091,N_1582);
nor U2570 (N_2570,N_1703,N_2071);
nand U2571 (N_2571,N_1770,N_1757);
or U2572 (N_2572,N_1704,N_1750);
nand U2573 (N_2573,N_1974,N_1738);
nand U2574 (N_2574,N_1789,N_1842);
or U2575 (N_2575,N_1654,N_1575);
nand U2576 (N_2576,N_1680,N_1843);
or U2577 (N_2577,N_1662,N_1607);
nand U2578 (N_2578,N_2220,N_1686);
nand U2579 (N_2579,N_1816,N_1741);
nand U2580 (N_2580,N_1891,N_2188);
nand U2581 (N_2581,N_1942,N_1864);
nor U2582 (N_2582,N_1663,N_1580);
nor U2583 (N_2583,N_2154,N_1641);
xnor U2584 (N_2584,N_2098,N_1807);
nand U2585 (N_2585,N_2244,N_2077);
and U2586 (N_2586,N_1508,N_1678);
or U2587 (N_2587,N_1837,N_1769);
nand U2588 (N_2588,N_1840,N_1649);
nor U2589 (N_2589,N_1726,N_1688);
nor U2590 (N_2590,N_2114,N_2034);
nor U2591 (N_2591,N_1657,N_2018);
nand U2592 (N_2592,N_2200,N_1772);
nand U2593 (N_2593,N_1517,N_2189);
and U2594 (N_2594,N_2164,N_2192);
nand U2595 (N_2595,N_2108,N_1764);
or U2596 (N_2596,N_1801,N_1924);
xor U2597 (N_2597,N_1933,N_2208);
and U2598 (N_2598,N_2008,N_2212);
or U2599 (N_2599,N_2109,N_1863);
nand U2600 (N_2600,N_1504,N_2087);
nor U2601 (N_2601,N_1917,N_1979);
or U2602 (N_2602,N_1773,N_2146);
nand U2603 (N_2603,N_1907,N_2242);
nand U2604 (N_2604,N_1529,N_2068);
and U2605 (N_2605,N_2125,N_1865);
or U2606 (N_2606,N_1886,N_1540);
xnor U2607 (N_2607,N_2134,N_1838);
nor U2608 (N_2608,N_1874,N_2016);
and U2609 (N_2609,N_1644,N_1887);
and U2610 (N_2610,N_2080,N_1623);
or U2611 (N_2611,N_1929,N_2121);
nand U2612 (N_2612,N_1655,N_1578);
nand U2613 (N_2613,N_1814,N_1913);
nand U2614 (N_2614,N_1943,N_1530);
nor U2615 (N_2615,N_1866,N_2138);
or U2616 (N_2616,N_1585,N_1981);
nor U2617 (N_2617,N_2104,N_2169);
nand U2618 (N_2618,N_1777,N_1752);
nand U2619 (N_2619,N_1636,N_2066);
xnor U2620 (N_2620,N_1564,N_1922);
and U2621 (N_2621,N_1811,N_1823);
or U2622 (N_2622,N_2005,N_1938);
xor U2623 (N_2623,N_1551,N_1619);
or U2624 (N_2624,N_1815,N_2051);
nor U2625 (N_2625,N_1821,N_1657);
nor U2626 (N_2626,N_1968,N_1634);
nor U2627 (N_2627,N_1890,N_1574);
nand U2628 (N_2628,N_2040,N_2116);
nor U2629 (N_2629,N_2142,N_2185);
nand U2630 (N_2630,N_2158,N_1579);
or U2631 (N_2631,N_2010,N_2181);
nand U2632 (N_2632,N_2093,N_1688);
or U2633 (N_2633,N_1597,N_1651);
nor U2634 (N_2634,N_1806,N_2246);
nand U2635 (N_2635,N_1640,N_1638);
nor U2636 (N_2636,N_2173,N_1744);
and U2637 (N_2637,N_1598,N_2200);
xor U2638 (N_2638,N_1879,N_1865);
nor U2639 (N_2639,N_2107,N_1683);
or U2640 (N_2640,N_1570,N_2074);
xnor U2641 (N_2641,N_1553,N_1835);
xor U2642 (N_2642,N_2230,N_2037);
nand U2643 (N_2643,N_1685,N_1981);
and U2644 (N_2644,N_1613,N_1556);
or U2645 (N_2645,N_1619,N_1911);
xor U2646 (N_2646,N_2077,N_1987);
nand U2647 (N_2647,N_1898,N_1845);
nand U2648 (N_2648,N_1650,N_1935);
nand U2649 (N_2649,N_2109,N_1546);
nand U2650 (N_2650,N_1993,N_1703);
nand U2651 (N_2651,N_1928,N_1503);
nor U2652 (N_2652,N_2075,N_2047);
and U2653 (N_2653,N_1654,N_1660);
nand U2654 (N_2654,N_1704,N_1638);
and U2655 (N_2655,N_1901,N_1836);
and U2656 (N_2656,N_2191,N_1533);
nand U2657 (N_2657,N_1547,N_1953);
and U2658 (N_2658,N_1850,N_1639);
or U2659 (N_2659,N_2000,N_2206);
nor U2660 (N_2660,N_1635,N_1878);
nand U2661 (N_2661,N_1972,N_1783);
and U2662 (N_2662,N_1828,N_1823);
or U2663 (N_2663,N_1604,N_2032);
and U2664 (N_2664,N_2222,N_1558);
nand U2665 (N_2665,N_2055,N_2200);
nand U2666 (N_2666,N_1570,N_2009);
and U2667 (N_2667,N_1952,N_1971);
nand U2668 (N_2668,N_2059,N_2203);
xor U2669 (N_2669,N_2141,N_1691);
or U2670 (N_2670,N_2030,N_2177);
or U2671 (N_2671,N_1935,N_1652);
nand U2672 (N_2672,N_1833,N_1612);
and U2673 (N_2673,N_1972,N_1502);
nor U2674 (N_2674,N_1510,N_1792);
or U2675 (N_2675,N_2132,N_1996);
nor U2676 (N_2676,N_1855,N_1534);
nor U2677 (N_2677,N_1612,N_2072);
nor U2678 (N_2678,N_1666,N_2111);
and U2679 (N_2679,N_1882,N_1636);
xnor U2680 (N_2680,N_2045,N_2229);
nand U2681 (N_2681,N_1565,N_1864);
nand U2682 (N_2682,N_1831,N_1859);
xnor U2683 (N_2683,N_1950,N_1693);
xor U2684 (N_2684,N_2218,N_1922);
or U2685 (N_2685,N_1729,N_2123);
nor U2686 (N_2686,N_1696,N_1509);
or U2687 (N_2687,N_2122,N_2012);
nand U2688 (N_2688,N_1561,N_2121);
nor U2689 (N_2689,N_1531,N_2232);
or U2690 (N_2690,N_2190,N_1606);
nor U2691 (N_2691,N_1640,N_1955);
or U2692 (N_2692,N_1873,N_1727);
and U2693 (N_2693,N_2120,N_1793);
nor U2694 (N_2694,N_2124,N_2236);
and U2695 (N_2695,N_1778,N_1776);
or U2696 (N_2696,N_1967,N_1937);
nand U2697 (N_2697,N_2222,N_1892);
nand U2698 (N_2698,N_1991,N_1731);
or U2699 (N_2699,N_1645,N_1637);
nand U2700 (N_2700,N_1619,N_1686);
nor U2701 (N_2701,N_2235,N_1872);
nand U2702 (N_2702,N_1866,N_2083);
nand U2703 (N_2703,N_2094,N_2226);
or U2704 (N_2704,N_1695,N_2217);
nor U2705 (N_2705,N_2248,N_1752);
or U2706 (N_2706,N_1616,N_2053);
or U2707 (N_2707,N_1781,N_1531);
or U2708 (N_2708,N_2060,N_1938);
and U2709 (N_2709,N_1548,N_2117);
nor U2710 (N_2710,N_2183,N_1619);
nand U2711 (N_2711,N_1598,N_2192);
nand U2712 (N_2712,N_2039,N_2227);
and U2713 (N_2713,N_1519,N_1687);
xnor U2714 (N_2714,N_2176,N_1789);
and U2715 (N_2715,N_1778,N_1915);
and U2716 (N_2716,N_2124,N_1994);
or U2717 (N_2717,N_1700,N_2020);
nand U2718 (N_2718,N_1510,N_2171);
or U2719 (N_2719,N_1846,N_2074);
or U2720 (N_2720,N_2071,N_1813);
and U2721 (N_2721,N_1557,N_1636);
and U2722 (N_2722,N_1613,N_2092);
and U2723 (N_2723,N_1703,N_1515);
nand U2724 (N_2724,N_1832,N_2047);
nor U2725 (N_2725,N_1519,N_1864);
and U2726 (N_2726,N_2205,N_1880);
xnor U2727 (N_2727,N_1543,N_1781);
nor U2728 (N_2728,N_1666,N_1534);
nand U2729 (N_2729,N_1642,N_1765);
nand U2730 (N_2730,N_1564,N_1605);
or U2731 (N_2731,N_1801,N_2111);
and U2732 (N_2732,N_1658,N_1918);
and U2733 (N_2733,N_1840,N_2076);
nand U2734 (N_2734,N_1751,N_1832);
nor U2735 (N_2735,N_2153,N_1772);
or U2736 (N_2736,N_2167,N_1721);
or U2737 (N_2737,N_1945,N_2088);
nor U2738 (N_2738,N_1712,N_1674);
and U2739 (N_2739,N_2030,N_1806);
xor U2740 (N_2740,N_1543,N_2178);
and U2741 (N_2741,N_1749,N_2008);
nor U2742 (N_2742,N_1969,N_2034);
xor U2743 (N_2743,N_1520,N_1989);
or U2744 (N_2744,N_2009,N_1529);
and U2745 (N_2745,N_2194,N_2156);
nor U2746 (N_2746,N_2095,N_1842);
nand U2747 (N_2747,N_1845,N_1938);
nand U2748 (N_2748,N_1950,N_1663);
and U2749 (N_2749,N_1592,N_1679);
or U2750 (N_2750,N_1774,N_1743);
and U2751 (N_2751,N_1901,N_1949);
and U2752 (N_2752,N_2120,N_1851);
and U2753 (N_2753,N_2215,N_1870);
and U2754 (N_2754,N_1526,N_2033);
and U2755 (N_2755,N_1763,N_2225);
nor U2756 (N_2756,N_2089,N_2127);
nor U2757 (N_2757,N_2144,N_1866);
nand U2758 (N_2758,N_1873,N_1560);
nor U2759 (N_2759,N_1648,N_1934);
nor U2760 (N_2760,N_1869,N_1905);
xnor U2761 (N_2761,N_1564,N_2052);
xnor U2762 (N_2762,N_1816,N_1940);
and U2763 (N_2763,N_1756,N_2044);
or U2764 (N_2764,N_2098,N_1820);
nor U2765 (N_2765,N_1928,N_1546);
nand U2766 (N_2766,N_1658,N_1700);
nor U2767 (N_2767,N_1878,N_1983);
or U2768 (N_2768,N_1992,N_1515);
nand U2769 (N_2769,N_2067,N_2096);
and U2770 (N_2770,N_2234,N_1594);
xor U2771 (N_2771,N_1574,N_2055);
and U2772 (N_2772,N_1563,N_2228);
or U2773 (N_2773,N_2044,N_1547);
xnor U2774 (N_2774,N_1602,N_1998);
nand U2775 (N_2775,N_1668,N_2124);
and U2776 (N_2776,N_1877,N_2091);
and U2777 (N_2777,N_1924,N_1665);
nand U2778 (N_2778,N_2129,N_2211);
or U2779 (N_2779,N_1511,N_1512);
nand U2780 (N_2780,N_1609,N_1662);
nor U2781 (N_2781,N_1523,N_1693);
or U2782 (N_2782,N_1520,N_1967);
or U2783 (N_2783,N_1947,N_2001);
nor U2784 (N_2784,N_2172,N_1737);
nand U2785 (N_2785,N_1740,N_1675);
or U2786 (N_2786,N_2070,N_2130);
nand U2787 (N_2787,N_1510,N_1551);
nand U2788 (N_2788,N_1868,N_1666);
and U2789 (N_2789,N_1528,N_1803);
nand U2790 (N_2790,N_1564,N_1578);
and U2791 (N_2791,N_2211,N_1651);
or U2792 (N_2792,N_1910,N_1570);
or U2793 (N_2793,N_2065,N_1974);
or U2794 (N_2794,N_1894,N_2102);
nor U2795 (N_2795,N_2201,N_1559);
or U2796 (N_2796,N_2138,N_1878);
or U2797 (N_2797,N_2021,N_1767);
or U2798 (N_2798,N_1583,N_1688);
nand U2799 (N_2799,N_1848,N_2113);
or U2800 (N_2800,N_2111,N_1563);
nor U2801 (N_2801,N_2012,N_2029);
nor U2802 (N_2802,N_1891,N_1815);
nand U2803 (N_2803,N_1961,N_2102);
nand U2804 (N_2804,N_2079,N_1506);
or U2805 (N_2805,N_1661,N_1985);
and U2806 (N_2806,N_1946,N_1767);
xnor U2807 (N_2807,N_1844,N_1630);
nand U2808 (N_2808,N_1654,N_1942);
or U2809 (N_2809,N_1706,N_1818);
nand U2810 (N_2810,N_1618,N_1765);
nand U2811 (N_2811,N_1538,N_2017);
or U2812 (N_2812,N_1690,N_1869);
and U2813 (N_2813,N_2179,N_1801);
nor U2814 (N_2814,N_1965,N_1505);
xor U2815 (N_2815,N_1957,N_1623);
and U2816 (N_2816,N_1673,N_2110);
nor U2817 (N_2817,N_1975,N_1790);
nor U2818 (N_2818,N_2103,N_1740);
and U2819 (N_2819,N_1632,N_1850);
nand U2820 (N_2820,N_1952,N_1976);
nand U2821 (N_2821,N_1719,N_1582);
or U2822 (N_2822,N_2056,N_1558);
nor U2823 (N_2823,N_1524,N_1645);
nor U2824 (N_2824,N_1703,N_2043);
nand U2825 (N_2825,N_1622,N_2122);
nor U2826 (N_2826,N_2206,N_2048);
nand U2827 (N_2827,N_1599,N_2214);
and U2828 (N_2828,N_2173,N_2196);
xor U2829 (N_2829,N_2160,N_2024);
and U2830 (N_2830,N_1912,N_1589);
nor U2831 (N_2831,N_2136,N_1725);
xor U2832 (N_2832,N_2103,N_1825);
nand U2833 (N_2833,N_2097,N_1896);
or U2834 (N_2834,N_2237,N_2037);
or U2835 (N_2835,N_2173,N_1886);
or U2836 (N_2836,N_2043,N_1882);
nand U2837 (N_2837,N_2040,N_1546);
or U2838 (N_2838,N_1590,N_2177);
or U2839 (N_2839,N_1605,N_1936);
or U2840 (N_2840,N_1847,N_1511);
and U2841 (N_2841,N_1684,N_1862);
nor U2842 (N_2842,N_2047,N_1513);
nand U2843 (N_2843,N_1515,N_1704);
nor U2844 (N_2844,N_1978,N_1842);
or U2845 (N_2845,N_2091,N_1936);
or U2846 (N_2846,N_2088,N_1507);
or U2847 (N_2847,N_1550,N_1906);
nand U2848 (N_2848,N_1533,N_1528);
or U2849 (N_2849,N_1872,N_1754);
xor U2850 (N_2850,N_2068,N_1676);
or U2851 (N_2851,N_1743,N_2072);
and U2852 (N_2852,N_1957,N_2218);
or U2853 (N_2853,N_1916,N_2028);
or U2854 (N_2854,N_2164,N_1734);
xnor U2855 (N_2855,N_1674,N_2178);
nor U2856 (N_2856,N_1713,N_1615);
and U2857 (N_2857,N_1900,N_1746);
or U2858 (N_2858,N_2124,N_1857);
nand U2859 (N_2859,N_1541,N_1511);
and U2860 (N_2860,N_2049,N_1700);
nand U2861 (N_2861,N_2061,N_1870);
and U2862 (N_2862,N_1843,N_1587);
nand U2863 (N_2863,N_1747,N_2153);
nor U2864 (N_2864,N_1776,N_2223);
nand U2865 (N_2865,N_1610,N_1827);
nor U2866 (N_2866,N_2174,N_1887);
nand U2867 (N_2867,N_2234,N_2037);
nand U2868 (N_2868,N_2145,N_2194);
nand U2869 (N_2869,N_1614,N_1634);
or U2870 (N_2870,N_2119,N_1920);
or U2871 (N_2871,N_1719,N_2223);
nand U2872 (N_2872,N_1893,N_1607);
nand U2873 (N_2873,N_2121,N_1831);
xnor U2874 (N_2874,N_1610,N_2228);
nand U2875 (N_2875,N_1617,N_2027);
or U2876 (N_2876,N_1575,N_2102);
xor U2877 (N_2877,N_1606,N_1834);
and U2878 (N_2878,N_1706,N_1705);
nand U2879 (N_2879,N_1614,N_1869);
or U2880 (N_2880,N_2222,N_1647);
or U2881 (N_2881,N_1893,N_1671);
and U2882 (N_2882,N_1708,N_1570);
xnor U2883 (N_2883,N_2053,N_2058);
nand U2884 (N_2884,N_1979,N_1906);
xor U2885 (N_2885,N_1574,N_1644);
xnor U2886 (N_2886,N_1950,N_1985);
or U2887 (N_2887,N_2181,N_2246);
and U2888 (N_2888,N_1724,N_2111);
or U2889 (N_2889,N_2002,N_1553);
nand U2890 (N_2890,N_1536,N_1647);
or U2891 (N_2891,N_1781,N_1587);
or U2892 (N_2892,N_1808,N_1618);
nor U2893 (N_2893,N_1756,N_1702);
and U2894 (N_2894,N_1782,N_1728);
nor U2895 (N_2895,N_2242,N_1738);
and U2896 (N_2896,N_1595,N_1726);
or U2897 (N_2897,N_1699,N_1574);
nor U2898 (N_2898,N_1914,N_2176);
nor U2899 (N_2899,N_1653,N_2118);
nor U2900 (N_2900,N_1951,N_1565);
nor U2901 (N_2901,N_2024,N_1889);
xor U2902 (N_2902,N_1936,N_1706);
nand U2903 (N_2903,N_1598,N_1980);
and U2904 (N_2904,N_1929,N_2171);
nor U2905 (N_2905,N_1762,N_2036);
nand U2906 (N_2906,N_2233,N_2245);
nand U2907 (N_2907,N_1850,N_2161);
nand U2908 (N_2908,N_1941,N_2210);
or U2909 (N_2909,N_1822,N_1500);
or U2910 (N_2910,N_1928,N_2033);
xnor U2911 (N_2911,N_1898,N_1843);
and U2912 (N_2912,N_2051,N_1701);
and U2913 (N_2913,N_2214,N_1698);
and U2914 (N_2914,N_1853,N_2194);
nor U2915 (N_2915,N_2064,N_1914);
nor U2916 (N_2916,N_1881,N_1509);
nand U2917 (N_2917,N_1502,N_1744);
nand U2918 (N_2918,N_1761,N_2062);
or U2919 (N_2919,N_1600,N_1915);
or U2920 (N_2920,N_1835,N_2068);
nand U2921 (N_2921,N_1534,N_1568);
or U2922 (N_2922,N_2152,N_1987);
nand U2923 (N_2923,N_1949,N_2093);
xnor U2924 (N_2924,N_2080,N_1785);
nor U2925 (N_2925,N_2029,N_2067);
and U2926 (N_2926,N_1881,N_2146);
and U2927 (N_2927,N_1927,N_1720);
or U2928 (N_2928,N_1539,N_1773);
nand U2929 (N_2929,N_1921,N_1599);
and U2930 (N_2930,N_2086,N_2004);
nor U2931 (N_2931,N_1949,N_1754);
or U2932 (N_2932,N_1834,N_1979);
and U2933 (N_2933,N_1967,N_1871);
nor U2934 (N_2934,N_1629,N_1877);
or U2935 (N_2935,N_1967,N_1847);
nor U2936 (N_2936,N_2009,N_1552);
and U2937 (N_2937,N_1809,N_1919);
and U2938 (N_2938,N_1970,N_1611);
nand U2939 (N_2939,N_1587,N_1599);
nor U2940 (N_2940,N_1770,N_1825);
nor U2941 (N_2941,N_1968,N_1714);
nor U2942 (N_2942,N_1933,N_2249);
nand U2943 (N_2943,N_1998,N_1562);
and U2944 (N_2944,N_2066,N_2015);
or U2945 (N_2945,N_1966,N_1926);
nor U2946 (N_2946,N_1862,N_1709);
and U2947 (N_2947,N_2016,N_2110);
nand U2948 (N_2948,N_2191,N_1888);
nor U2949 (N_2949,N_2078,N_1903);
and U2950 (N_2950,N_1540,N_2018);
nand U2951 (N_2951,N_1938,N_2202);
or U2952 (N_2952,N_2028,N_1770);
or U2953 (N_2953,N_1795,N_2229);
nand U2954 (N_2954,N_2072,N_1732);
and U2955 (N_2955,N_1998,N_1781);
nand U2956 (N_2956,N_1756,N_2216);
nor U2957 (N_2957,N_1857,N_1729);
and U2958 (N_2958,N_1946,N_1728);
nor U2959 (N_2959,N_2206,N_1776);
nand U2960 (N_2960,N_2192,N_1538);
and U2961 (N_2961,N_2241,N_1857);
or U2962 (N_2962,N_1978,N_1561);
nor U2963 (N_2963,N_1691,N_1920);
nand U2964 (N_2964,N_1677,N_2237);
nor U2965 (N_2965,N_1702,N_2173);
or U2966 (N_2966,N_2096,N_1923);
nor U2967 (N_2967,N_1808,N_2225);
and U2968 (N_2968,N_2035,N_1836);
nor U2969 (N_2969,N_1752,N_1524);
nand U2970 (N_2970,N_1539,N_1502);
nor U2971 (N_2971,N_2039,N_2157);
or U2972 (N_2972,N_1538,N_2019);
or U2973 (N_2973,N_2138,N_2119);
nor U2974 (N_2974,N_1859,N_1732);
nand U2975 (N_2975,N_1779,N_2132);
nor U2976 (N_2976,N_1640,N_2247);
nand U2977 (N_2977,N_1968,N_2205);
or U2978 (N_2978,N_2113,N_2123);
nand U2979 (N_2979,N_2103,N_2147);
nor U2980 (N_2980,N_1830,N_2207);
xor U2981 (N_2981,N_1814,N_2041);
nor U2982 (N_2982,N_2188,N_2175);
nor U2983 (N_2983,N_1709,N_2076);
and U2984 (N_2984,N_1707,N_1836);
and U2985 (N_2985,N_1584,N_1831);
nor U2986 (N_2986,N_1935,N_1799);
and U2987 (N_2987,N_1920,N_1559);
xor U2988 (N_2988,N_1802,N_2150);
or U2989 (N_2989,N_1607,N_1921);
and U2990 (N_2990,N_1575,N_2035);
nand U2991 (N_2991,N_1909,N_1934);
nand U2992 (N_2992,N_1960,N_2245);
nor U2993 (N_2993,N_2138,N_2156);
nor U2994 (N_2994,N_2006,N_2128);
or U2995 (N_2995,N_2181,N_1901);
nand U2996 (N_2996,N_2049,N_2219);
nand U2997 (N_2997,N_1880,N_1628);
and U2998 (N_2998,N_1532,N_1760);
nor U2999 (N_2999,N_1976,N_1765);
nor UO_0 (O_0,N_2403,N_2751);
nand UO_1 (O_1,N_2841,N_2357);
xor UO_2 (O_2,N_2254,N_2373);
nand UO_3 (O_3,N_2573,N_2265);
nor UO_4 (O_4,N_2398,N_2500);
and UO_5 (O_5,N_2526,N_2554);
nor UO_6 (O_6,N_2761,N_2396);
or UO_7 (O_7,N_2280,N_2728);
nand UO_8 (O_8,N_2452,N_2581);
or UO_9 (O_9,N_2287,N_2406);
nand UO_10 (O_10,N_2446,N_2772);
and UO_11 (O_11,N_2831,N_2474);
nand UO_12 (O_12,N_2683,N_2301);
nor UO_13 (O_13,N_2627,N_2976);
and UO_14 (O_14,N_2738,N_2495);
and UO_15 (O_15,N_2733,N_2777);
or UO_16 (O_16,N_2659,N_2596);
xnor UO_17 (O_17,N_2655,N_2444);
nand UO_18 (O_18,N_2578,N_2663);
nor UO_19 (O_19,N_2939,N_2887);
and UO_20 (O_20,N_2530,N_2984);
xor UO_21 (O_21,N_2970,N_2767);
nor UO_22 (O_22,N_2802,N_2670);
and UO_23 (O_23,N_2325,N_2516);
or UO_24 (O_24,N_2464,N_2525);
nor UO_25 (O_25,N_2730,N_2812);
or UO_26 (O_26,N_2508,N_2857);
xnor UO_27 (O_27,N_2645,N_2523);
nor UO_28 (O_28,N_2271,N_2756);
nor UO_29 (O_29,N_2296,N_2909);
nand UO_30 (O_30,N_2910,N_2443);
nand UO_31 (O_31,N_2992,N_2471);
xnor UO_32 (O_32,N_2690,N_2521);
or UO_33 (O_33,N_2954,N_2313);
or UO_34 (O_34,N_2441,N_2658);
nand UO_35 (O_35,N_2618,N_2652);
and UO_36 (O_36,N_2335,N_2413);
or UO_37 (O_37,N_2374,N_2358);
or UO_38 (O_38,N_2892,N_2987);
and UO_39 (O_39,N_2372,N_2983);
and UO_40 (O_40,N_2329,N_2380);
and UO_41 (O_41,N_2598,N_2896);
xnor UO_42 (O_42,N_2858,N_2447);
or UO_43 (O_43,N_2758,N_2964);
nand UO_44 (O_44,N_2996,N_2603);
xor UO_45 (O_45,N_2536,N_2883);
and UO_46 (O_46,N_2575,N_2846);
or UO_47 (O_47,N_2307,N_2929);
nor UO_48 (O_48,N_2469,N_2919);
or UO_49 (O_49,N_2366,N_2499);
and UO_50 (O_50,N_2449,N_2369);
nand UO_51 (O_51,N_2341,N_2590);
nor UO_52 (O_52,N_2453,N_2251);
and UO_53 (O_53,N_2537,N_2632);
nor UO_54 (O_54,N_2308,N_2486);
xnor UO_55 (O_55,N_2780,N_2750);
nand UO_56 (O_56,N_2926,N_2282);
nand UO_57 (O_57,N_2894,N_2807);
nand UO_58 (O_58,N_2975,N_2512);
nand UO_59 (O_59,N_2292,N_2545);
and UO_60 (O_60,N_2572,N_2799);
and UO_61 (O_61,N_2788,N_2724);
and UO_62 (O_62,N_2615,N_2813);
xnor UO_63 (O_63,N_2961,N_2672);
and UO_64 (O_64,N_2468,N_2888);
nor UO_65 (O_65,N_2700,N_2644);
nor UO_66 (O_66,N_2737,N_2640);
and UO_67 (O_67,N_2582,N_2747);
nor UO_68 (O_68,N_2462,N_2511);
nor UO_69 (O_69,N_2570,N_2790);
nor UO_70 (O_70,N_2560,N_2868);
nor UO_71 (O_71,N_2899,N_2819);
nand UO_72 (O_72,N_2520,N_2943);
nand UO_73 (O_73,N_2326,N_2533);
or UO_74 (O_74,N_2787,N_2876);
and UO_75 (O_75,N_2907,N_2740);
nand UO_76 (O_76,N_2707,N_2522);
or UO_77 (O_77,N_2956,N_2934);
and UO_78 (O_78,N_2829,N_2823);
and UO_79 (O_79,N_2753,N_2382);
nand UO_80 (O_80,N_2912,N_2998);
nor UO_81 (O_81,N_2255,N_2601);
nor UO_82 (O_82,N_2642,N_2354);
nand UO_83 (O_83,N_2990,N_2279);
nand UO_84 (O_84,N_2257,N_2597);
nand UO_85 (O_85,N_2490,N_2551);
nor UO_86 (O_86,N_2891,N_2338);
xnor UO_87 (O_87,N_2836,N_2681);
nand UO_88 (O_88,N_2631,N_2898);
xnor UO_89 (O_89,N_2874,N_2513);
or UO_90 (O_90,N_2386,N_2491);
and UO_91 (O_91,N_2774,N_2332);
nor UO_92 (O_92,N_2267,N_2978);
nor UO_93 (O_93,N_2701,N_2565);
and UO_94 (O_94,N_2922,N_2830);
nor UO_95 (O_95,N_2404,N_2930);
xor UO_96 (O_96,N_2626,N_2673);
xnor UO_97 (O_97,N_2370,N_2843);
and UO_98 (O_98,N_2960,N_2347);
nor UO_99 (O_99,N_2853,N_2743);
and UO_100 (O_100,N_2311,N_2872);
and UO_101 (O_101,N_2734,N_2465);
and UO_102 (O_102,N_2628,N_2320);
nand UO_103 (O_103,N_2412,N_2873);
and UO_104 (O_104,N_2262,N_2433);
nand UO_105 (O_105,N_2339,N_2826);
and UO_106 (O_106,N_2312,N_2540);
and UO_107 (O_107,N_2477,N_2387);
nand UO_108 (O_108,N_2483,N_2639);
xor UO_109 (O_109,N_2429,N_2726);
and UO_110 (O_110,N_2529,N_2967);
nand UO_111 (O_111,N_2869,N_2664);
and UO_112 (O_112,N_2427,N_2850);
or UO_113 (O_113,N_2507,N_2505);
nand UO_114 (O_114,N_2416,N_2949);
and UO_115 (O_115,N_2637,N_2344);
and UO_116 (O_116,N_2721,N_2771);
and UO_117 (O_117,N_2393,N_2454);
or UO_118 (O_118,N_2867,N_2902);
nor UO_119 (O_119,N_2293,N_2297);
nand UO_120 (O_120,N_2426,N_2343);
and UO_121 (O_121,N_2793,N_2256);
nand UO_122 (O_122,N_2784,N_2501);
and UO_123 (O_123,N_2608,N_2776);
and UO_124 (O_124,N_2671,N_2415);
nand UO_125 (O_125,N_2913,N_2834);
nand UO_126 (O_126,N_2363,N_2669);
and UO_127 (O_127,N_2379,N_2641);
and UO_128 (O_128,N_2622,N_2623);
and UO_129 (O_129,N_2588,N_2725);
or UO_130 (O_130,N_2971,N_2806);
or UO_131 (O_131,N_2745,N_2803);
nand UO_132 (O_132,N_2569,N_2835);
or UO_133 (O_133,N_2801,N_2440);
nor UO_134 (O_134,N_2274,N_2619);
nand UO_135 (O_135,N_2478,N_2268);
nor UO_136 (O_136,N_2804,N_2583);
nor UO_137 (O_137,N_2811,N_2317);
or UO_138 (O_138,N_2392,N_2364);
and UO_139 (O_139,N_2742,N_2283);
and UO_140 (O_140,N_2717,N_2821);
nand UO_141 (O_141,N_2861,N_2259);
or UO_142 (O_142,N_2918,N_2488);
nor UO_143 (O_143,N_2548,N_2924);
or UO_144 (O_144,N_2435,N_2845);
nor UO_145 (O_145,N_2617,N_2290);
or UO_146 (O_146,N_2880,N_2532);
nor UO_147 (O_147,N_2599,N_2385);
and UO_148 (O_148,N_2503,N_2824);
nand UO_149 (O_149,N_2306,N_2281);
and UO_150 (O_150,N_2436,N_2475);
nand UO_151 (O_151,N_2579,N_2557);
nor UO_152 (O_152,N_2410,N_2625);
xnor UO_153 (O_153,N_2263,N_2752);
or UO_154 (O_154,N_2527,N_2367);
nor UO_155 (O_155,N_2712,N_2482);
nand UO_156 (O_156,N_2968,N_2504);
and UO_157 (O_157,N_2542,N_2739);
nand UO_158 (O_158,N_2713,N_2849);
nor UO_159 (O_159,N_2871,N_2962);
and UO_160 (O_160,N_2350,N_2352);
and UO_161 (O_161,N_2999,N_2566);
and UO_162 (O_162,N_2825,N_2650);
and UO_163 (O_163,N_2820,N_2484);
nor UO_164 (O_164,N_2361,N_2269);
nand UO_165 (O_165,N_2792,N_2421);
nor UO_166 (O_166,N_2827,N_2252);
nand UO_167 (O_167,N_2714,N_2609);
and UO_168 (O_168,N_2679,N_2284);
xnor UO_169 (O_169,N_2286,N_2731);
xor UO_170 (O_170,N_2766,N_2794);
nand UO_171 (O_171,N_2559,N_2986);
nand UO_172 (O_172,N_2328,N_2316);
and UO_173 (O_173,N_2353,N_2305);
nor UO_174 (O_174,N_2715,N_2260);
or UO_175 (O_175,N_2321,N_2549);
nor UO_176 (O_176,N_2915,N_2895);
nand UO_177 (O_177,N_2727,N_2677);
or UO_178 (O_178,N_2764,N_2950);
and UO_179 (O_179,N_2675,N_2648);
nand UO_180 (O_180,N_2635,N_2381);
nand UO_181 (O_181,N_2594,N_2607);
xor UO_182 (O_182,N_2988,N_2921);
nand UO_183 (O_183,N_2535,N_2476);
and UO_184 (O_184,N_2275,N_2458);
and UO_185 (O_185,N_2318,N_2629);
nor UO_186 (O_186,N_2757,N_2732);
nand UO_187 (O_187,N_2839,N_2684);
nand UO_188 (O_188,N_2706,N_2917);
or UO_189 (O_189,N_2543,N_2748);
nand UO_190 (O_190,N_2779,N_2571);
and UO_191 (O_191,N_2408,N_2746);
or UO_192 (O_192,N_2345,N_2866);
and UO_193 (O_193,N_2833,N_2294);
nand UO_194 (O_194,N_2696,N_2704);
or UO_195 (O_195,N_2638,N_2711);
nand UO_196 (O_196,N_2762,N_2816);
nor UO_197 (O_197,N_2314,N_2291);
and UO_198 (O_198,N_2703,N_2550);
nor UO_199 (O_199,N_2562,N_2589);
or UO_200 (O_200,N_2304,N_2428);
or UO_201 (O_201,N_2616,N_2981);
and UO_202 (O_202,N_2266,N_2948);
and UO_203 (O_203,N_2765,N_2585);
and UO_204 (O_204,N_2665,N_2995);
nand UO_205 (O_205,N_2518,N_2974);
xnor UO_206 (O_206,N_2796,N_2510);
xnor UO_207 (O_207,N_2958,N_2502);
nor UO_208 (O_208,N_2591,N_2539);
and UO_209 (O_209,N_2994,N_2904);
xnor UO_210 (O_210,N_2815,N_2959);
or UO_211 (O_211,N_2937,N_2417);
nor UO_212 (O_212,N_2348,N_2362);
nor UO_213 (O_213,N_2310,N_2524);
and UO_214 (O_214,N_2678,N_2729);
nor UO_215 (O_215,N_2442,N_2997);
nand UO_216 (O_216,N_2933,N_2982);
nor UO_217 (O_217,N_2437,N_2276);
and UO_218 (O_218,N_2561,N_2553);
nor UO_219 (O_219,N_2384,N_2409);
xnor UO_220 (O_220,N_2870,N_2908);
and UO_221 (O_221,N_2558,N_2722);
or UO_222 (O_222,N_2351,N_2445);
or UO_223 (O_223,N_2587,N_2390);
nand UO_224 (O_224,N_2479,N_2461);
nand UO_225 (O_225,N_2250,N_2544);
and UO_226 (O_226,N_2837,N_2531);
or UO_227 (O_227,N_2697,N_2360);
xnor UO_228 (O_228,N_2319,N_2264);
and UO_229 (O_229,N_2528,N_2749);
nand UO_230 (O_230,N_2901,N_2346);
or UO_231 (O_231,N_2401,N_2755);
nor UO_232 (O_232,N_2480,N_2614);
nor UO_233 (O_233,N_2989,N_2333);
or UO_234 (O_234,N_2963,N_2840);
and UO_235 (O_235,N_2966,N_2782);
or UO_236 (O_236,N_2691,N_2969);
and UO_237 (O_237,N_2685,N_2977);
nand UO_238 (O_238,N_2315,N_2938);
nor UO_239 (O_239,N_2419,N_2927);
nand UO_240 (O_240,N_2633,N_2298);
nor UO_241 (O_241,N_2884,N_2580);
nand UO_242 (O_242,N_2710,N_2606);
and UO_243 (O_243,N_2568,N_2547);
nand UO_244 (O_244,N_2459,N_2340);
and UO_245 (O_245,N_2775,N_2705);
and UO_246 (O_246,N_2810,N_2770);
and UO_247 (O_247,N_2397,N_2916);
nand UO_248 (O_248,N_2947,N_2460);
nor UO_249 (O_249,N_2278,N_2388);
xor UO_250 (O_250,N_2688,N_2375);
nor UO_251 (O_251,N_2309,N_2498);
and UO_252 (O_252,N_2448,N_2514);
or UO_253 (O_253,N_2814,N_2719);
or UO_254 (O_254,N_2647,N_2768);
xor UO_255 (O_255,N_2695,N_2905);
nand UO_256 (O_256,N_2720,N_2928);
or UO_257 (O_257,N_2451,N_2931);
nand UO_258 (O_258,N_2646,N_2946);
or UO_259 (O_259,N_2923,N_2885);
and UO_260 (O_260,N_2337,N_2666);
nor UO_261 (O_261,N_2818,N_2649);
or UO_262 (O_262,N_2272,N_2359);
and UO_263 (O_263,N_2657,N_2651);
or UO_264 (O_264,N_2506,N_2661);
or UO_265 (O_265,N_2741,N_2791);
nor UO_266 (O_266,N_2330,N_2760);
and UO_267 (O_267,N_2759,N_2552);
or UO_268 (O_268,N_2630,N_2716);
nor UO_269 (O_269,N_2376,N_2723);
and UO_270 (O_270,N_2331,N_2420);
nand UO_271 (O_271,N_2405,N_2322);
nor UO_272 (O_272,N_2485,N_2694);
nand UO_273 (O_273,N_2430,N_2865);
nor UO_274 (O_274,N_2653,N_2920);
or UO_275 (O_275,N_2940,N_2854);
nor UO_276 (O_276,N_2334,N_2798);
or UO_277 (O_277,N_2680,N_2693);
and UO_278 (O_278,N_2431,N_2541);
and UO_279 (O_279,N_2261,N_2423);
and UO_280 (O_280,N_2686,N_2855);
or UO_281 (O_281,N_2487,N_2624);
and UO_282 (O_282,N_2538,N_2882);
nor UO_283 (O_283,N_2993,N_2941);
or UO_284 (O_284,N_2515,N_2481);
nand UO_285 (O_285,N_2809,N_2355);
nor UO_286 (O_286,N_2972,N_2991);
and UO_287 (O_287,N_2595,N_2844);
nor UO_288 (O_288,N_2832,N_2951);
nand UO_289 (O_289,N_2611,N_2494);
or UO_290 (O_290,N_2612,N_2473);
xnor UO_291 (O_291,N_2327,N_2273);
or UO_292 (O_292,N_2399,N_2593);
and UO_293 (O_293,N_2613,N_2323);
or UO_294 (O_294,N_2466,N_2875);
and UO_295 (O_295,N_2945,N_2600);
and UO_296 (O_296,N_2253,N_2258);
and UO_297 (O_297,N_2371,N_2735);
nor UO_298 (O_298,N_2556,N_2852);
or UO_299 (O_299,N_2708,N_2769);
nand UO_300 (O_300,N_2555,N_2288);
or UO_301 (O_301,N_2576,N_2592);
or UO_302 (O_302,N_2605,N_2878);
nor UO_303 (O_303,N_2795,N_2699);
and UO_304 (O_304,N_2944,N_2763);
nand UO_305 (O_305,N_2687,N_2942);
or UO_306 (O_306,N_2847,N_2604);
nor UO_307 (O_307,N_2324,N_2377);
or UO_308 (O_308,N_2395,N_2411);
xnor UO_309 (O_309,N_2965,N_2676);
and UO_310 (O_310,N_2574,N_2744);
or UO_311 (O_311,N_2973,N_2682);
or UO_312 (O_312,N_2509,N_2277);
or UO_313 (O_313,N_2467,N_2980);
and UO_314 (O_314,N_2620,N_2342);
or UO_315 (O_315,N_2879,N_2838);
or UO_316 (O_316,N_2952,N_2302);
and UO_317 (O_317,N_2698,N_2808);
nor UO_318 (O_318,N_2567,N_2425);
and UO_319 (O_319,N_2783,N_2654);
or UO_320 (O_320,N_2709,N_2881);
and UO_321 (O_321,N_2800,N_2295);
or UO_322 (O_322,N_2936,N_2414);
and UO_323 (O_323,N_2785,N_2389);
nor UO_324 (O_324,N_2434,N_2424);
nor UO_325 (O_325,N_2636,N_2356);
and UO_326 (O_326,N_2493,N_2667);
or UO_327 (O_327,N_2889,N_2817);
or UO_328 (O_328,N_2914,N_2497);
nor UO_329 (O_329,N_2336,N_2863);
nand UO_330 (O_330,N_2643,N_2668);
and UO_331 (O_331,N_2906,N_2584);
or UO_332 (O_332,N_2432,N_2903);
and UO_333 (O_333,N_2935,N_2455);
or UO_334 (O_334,N_2660,N_2985);
or UO_335 (O_335,N_2890,N_2692);
nor UO_336 (O_336,N_2900,N_2656);
or UO_337 (O_337,N_2450,N_2842);
nor UO_338 (O_338,N_2492,N_2862);
nand UO_339 (O_339,N_2407,N_2877);
and UO_340 (O_340,N_2289,N_2519);
nand UO_341 (O_341,N_2534,N_2270);
and UO_342 (O_342,N_2674,N_2953);
nor UO_343 (O_343,N_2299,N_2303);
or UO_344 (O_344,N_2564,N_2689);
nand UO_345 (O_345,N_2439,N_2402);
or UO_346 (O_346,N_2422,N_2463);
and UO_347 (O_347,N_2378,N_2859);
or UO_348 (O_348,N_2456,N_2472);
or UO_349 (O_349,N_2702,N_2955);
nor UO_350 (O_350,N_2349,N_2797);
or UO_351 (O_351,N_2860,N_2391);
or UO_352 (O_352,N_2781,N_2546);
xnor UO_353 (O_353,N_2864,N_2586);
or UO_354 (O_354,N_2621,N_2886);
nand UO_355 (O_355,N_2400,N_2932);
or UO_356 (O_356,N_2438,N_2470);
nor UO_357 (O_357,N_2718,N_2736);
nor UO_358 (O_358,N_2368,N_2418);
nor UO_359 (O_359,N_2489,N_2563);
and UO_360 (O_360,N_2925,N_2457);
or UO_361 (O_361,N_2848,N_2979);
or UO_362 (O_362,N_2365,N_2786);
nor UO_363 (O_363,N_2662,N_2394);
nand UO_364 (O_364,N_2828,N_2778);
nor UO_365 (O_365,N_2610,N_2517);
and UO_366 (O_366,N_2577,N_2856);
or UO_367 (O_367,N_2383,N_2634);
and UO_368 (O_368,N_2805,N_2822);
xor UO_369 (O_369,N_2893,N_2773);
or UO_370 (O_370,N_2602,N_2285);
and UO_371 (O_371,N_2851,N_2957);
nor UO_372 (O_372,N_2911,N_2754);
nor UO_373 (O_373,N_2897,N_2300);
and UO_374 (O_374,N_2789,N_2496);
or UO_375 (O_375,N_2463,N_2641);
nor UO_376 (O_376,N_2635,N_2719);
nand UO_377 (O_377,N_2941,N_2965);
or UO_378 (O_378,N_2676,N_2976);
nand UO_379 (O_379,N_2501,N_2804);
nand UO_380 (O_380,N_2725,N_2624);
nand UO_381 (O_381,N_2511,N_2756);
xor UO_382 (O_382,N_2696,N_2723);
nand UO_383 (O_383,N_2668,N_2943);
and UO_384 (O_384,N_2511,N_2339);
or UO_385 (O_385,N_2420,N_2510);
and UO_386 (O_386,N_2262,N_2735);
and UO_387 (O_387,N_2468,N_2687);
nor UO_388 (O_388,N_2814,N_2615);
xor UO_389 (O_389,N_2718,N_2396);
and UO_390 (O_390,N_2477,N_2687);
nor UO_391 (O_391,N_2488,N_2560);
or UO_392 (O_392,N_2438,N_2501);
and UO_393 (O_393,N_2397,N_2821);
nand UO_394 (O_394,N_2925,N_2330);
and UO_395 (O_395,N_2263,N_2253);
nand UO_396 (O_396,N_2995,N_2591);
and UO_397 (O_397,N_2743,N_2775);
and UO_398 (O_398,N_2750,N_2976);
nand UO_399 (O_399,N_2433,N_2392);
nand UO_400 (O_400,N_2777,N_2255);
and UO_401 (O_401,N_2385,N_2581);
xor UO_402 (O_402,N_2771,N_2353);
and UO_403 (O_403,N_2613,N_2917);
xor UO_404 (O_404,N_2717,N_2716);
nand UO_405 (O_405,N_2734,N_2975);
nand UO_406 (O_406,N_2741,N_2927);
and UO_407 (O_407,N_2462,N_2718);
nand UO_408 (O_408,N_2556,N_2883);
or UO_409 (O_409,N_2603,N_2264);
or UO_410 (O_410,N_2999,N_2401);
nor UO_411 (O_411,N_2529,N_2682);
nand UO_412 (O_412,N_2530,N_2794);
xor UO_413 (O_413,N_2712,N_2562);
nand UO_414 (O_414,N_2885,N_2449);
nand UO_415 (O_415,N_2676,N_2896);
nand UO_416 (O_416,N_2575,N_2746);
nor UO_417 (O_417,N_2854,N_2508);
nor UO_418 (O_418,N_2582,N_2489);
and UO_419 (O_419,N_2974,N_2816);
or UO_420 (O_420,N_2457,N_2478);
or UO_421 (O_421,N_2252,N_2880);
xor UO_422 (O_422,N_2308,N_2690);
nor UO_423 (O_423,N_2957,N_2788);
nor UO_424 (O_424,N_2623,N_2972);
xor UO_425 (O_425,N_2296,N_2623);
nor UO_426 (O_426,N_2327,N_2887);
nor UO_427 (O_427,N_2961,N_2543);
or UO_428 (O_428,N_2978,N_2662);
nand UO_429 (O_429,N_2735,N_2361);
nand UO_430 (O_430,N_2544,N_2480);
nor UO_431 (O_431,N_2761,N_2609);
nor UO_432 (O_432,N_2507,N_2394);
or UO_433 (O_433,N_2527,N_2955);
or UO_434 (O_434,N_2785,N_2426);
and UO_435 (O_435,N_2428,N_2958);
nor UO_436 (O_436,N_2835,N_2446);
xnor UO_437 (O_437,N_2845,N_2268);
and UO_438 (O_438,N_2673,N_2546);
or UO_439 (O_439,N_2524,N_2624);
xor UO_440 (O_440,N_2589,N_2899);
nor UO_441 (O_441,N_2883,N_2367);
xor UO_442 (O_442,N_2491,N_2273);
xor UO_443 (O_443,N_2519,N_2340);
nor UO_444 (O_444,N_2897,N_2821);
nand UO_445 (O_445,N_2380,N_2264);
or UO_446 (O_446,N_2290,N_2485);
nor UO_447 (O_447,N_2432,N_2626);
and UO_448 (O_448,N_2666,N_2653);
or UO_449 (O_449,N_2426,N_2916);
nor UO_450 (O_450,N_2367,N_2290);
nand UO_451 (O_451,N_2278,N_2384);
or UO_452 (O_452,N_2944,N_2777);
nand UO_453 (O_453,N_2787,N_2674);
nand UO_454 (O_454,N_2836,N_2570);
nor UO_455 (O_455,N_2449,N_2589);
xnor UO_456 (O_456,N_2847,N_2704);
and UO_457 (O_457,N_2383,N_2350);
and UO_458 (O_458,N_2793,N_2626);
and UO_459 (O_459,N_2729,N_2620);
or UO_460 (O_460,N_2304,N_2435);
nor UO_461 (O_461,N_2373,N_2401);
and UO_462 (O_462,N_2811,N_2399);
nand UO_463 (O_463,N_2887,N_2882);
and UO_464 (O_464,N_2760,N_2344);
nand UO_465 (O_465,N_2894,N_2293);
xor UO_466 (O_466,N_2655,N_2768);
and UO_467 (O_467,N_2955,N_2592);
nor UO_468 (O_468,N_2435,N_2460);
or UO_469 (O_469,N_2264,N_2574);
nand UO_470 (O_470,N_2668,N_2761);
nor UO_471 (O_471,N_2276,N_2715);
nor UO_472 (O_472,N_2262,N_2397);
nor UO_473 (O_473,N_2759,N_2549);
nand UO_474 (O_474,N_2337,N_2635);
nor UO_475 (O_475,N_2662,N_2268);
nor UO_476 (O_476,N_2652,N_2633);
nand UO_477 (O_477,N_2543,N_2261);
nand UO_478 (O_478,N_2636,N_2451);
nor UO_479 (O_479,N_2745,N_2912);
nand UO_480 (O_480,N_2952,N_2556);
and UO_481 (O_481,N_2966,N_2592);
or UO_482 (O_482,N_2604,N_2250);
nand UO_483 (O_483,N_2700,N_2763);
nor UO_484 (O_484,N_2862,N_2766);
nand UO_485 (O_485,N_2863,N_2561);
and UO_486 (O_486,N_2589,N_2996);
or UO_487 (O_487,N_2456,N_2698);
nand UO_488 (O_488,N_2804,N_2939);
or UO_489 (O_489,N_2262,N_2510);
xor UO_490 (O_490,N_2304,N_2701);
nor UO_491 (O_491,N_2873,N_2445);
xnor UO_492 (O_492,N_2554,N_2970);
or UO_493 (O_493,N_2298,N_2961);
nand UO_494 (O_494,N_2394,N_2719);
and UO_495 (O_495,N_2832,N_2742);
or UO_496 (O_496,N_2754,N_2919);
and UO_497 (O_497,N_2581,N_2954);
or UO_498 (O_498,N_2476,N_2953);
nor UO_499 (O_499,N_2863,N_2989);
endmodule