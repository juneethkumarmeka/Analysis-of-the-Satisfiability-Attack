module basic_750_5000_1000_2_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2510,N_2511,N_2512,N_2514,N_2516,N_2517,N_2518,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2537,N_2538,N_2539,N_2540,N_2541,N_2543,N_2544,N_2545,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2562,N_2564,N_2565,N_2567,N_2568,N_2569,N_2570,N_2571,N_2573,N_2574,N_2575,N_2576,N_2578,N_2579,N_2580,N_2581,N_2583,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2611,N_2612,N_2613,N_2615,N_2616,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2659,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2685,N_2686,N_2687,N_2688,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2738,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2757,N_2758,N_2760,N_2762,N_2763,N_2765,N_2766,N_2767,N_2768,N_2769,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2782,N_2784,N_2785,N_2787,N_2788,N_2790,N_2791,N_2792,N_2793,N_2795,N_2796,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2806,N_2807,N_2808,N_2809,N_2812,N_2813,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2832,N_2833,N_2834,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2855,N_2856,N_2857,N_2859,N_2860,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2911,N_2912,N_2913,N_2914,N_2916,N_2918,N_2920,N_2922,N_2923,N_2924,N_2925,N_2926,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2945,N_2946,N_2947,N_2950,N_2951,N_2952,N_2954,N_2955,N_2957,N_2958,N_2959,N_2961,N_2962,N_2963,N_2965,N_2966,N_2969,N_2970,N_2971,N_2972,N_2974,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2986,N_2988,N_2989,N_2990,N_2991,N_2992,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3013,N_3014,N_3015,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3033,N_3034,N_3035,N_3036,N_3037,N_3042,N_3043,N_3044,N_3045,N_3047,N_3048,N_3051,N_3052,N_3053,N_3055,N_3056,N_3057,N_3059,N_3061,N_3062,N_3063,N_3064,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3074,N_3077,N_3078,N_3079,N_3080,N_3081,N_3083,N_3084,N_3086,N_3087,N_3088,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3097,N_3098,N_3099,N_3100,N_3102,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3127,N_3129,N_3130,N_3131,N_3132,N_3134,N_3135,N_3136,N_3137,N_3138,N_3141,N_3142,N_3143,N_3144,N_3147,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3159,N_3160,N_3161,N_3162,N_3164,N_3165,N_3166,N_3167,N_3168,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3185,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3197,N_3199,N_3200,N_3201,N_3202,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3224,N_3225,N_3227,N_3228,N_3229,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3238,N_3239,N_3240,N_3241,N_3243,N_3246,N_3247,N_3248,N_3249,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3269,N_3270,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3282,N_3284,N_3285,N_3286,N_3287,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3302,N_3304,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3326,N_3327,N_3328,N_3329,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3342,N_3343,N_3345,N_3346,N_3347,N_3349,N_3350,N_3351,N_3352,N_3353,N_3355,N_3356,N_3357,N_3358,N_3359,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3378,N_3379,N_3380,N_3382,N_3383,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3394,N_3395,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3410,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3440,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3458,N_3459,N_3460,N_3462,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3471,N_3472,N_3473,N_3476,N_3478,N_3479,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3501,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3523,N_3524,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3535,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3545,N_3547,N_3548,N_3549,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3564,N_3565,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3583,N_3584,N_3585,N_3587,N_3589,N_3590,N_3591,N_3593,N_3594,N_3595,N_3597,N_3598,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3608,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3629,N_3630,N_3631,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3642,N_3644,N_3645,N_3646,N_3647,N_3648,N_3650,N_3651,N_3655,N_3656,N_3657,N_3658,N_3659,N_3661,N_3663,N_3664,N_3665,N_3666,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3680,N_3681,N_3682,N_3684,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3694,N_3695,N_3696,N_3698,N_3700,N_3701,N_3702,N_3703,N_3704,N_3706,N_3709,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3718,N_3719,N_3720,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3735,N_3737,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3747,N_3748,N_3749,N_3751,N_3752,N_3753,N_3754,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3767,N_3768,N_3769,N_3770,N_3772,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3782,N_3783,N_3784,N_3785,N_3786,N_3788,N_3789,N_3790,N_3791,N_3793,N_3797,N_3798,N_3799,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3814,N_3815,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3828,N_3829,N_3830,N_3832,N_3833,N_3834,N_3835,N_3837,N_3838,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3848,N_3849,N_3850,N_3851,N_3853,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3864,N_3865,N_3866,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3876,N_3877,N_3878,N_3880,N_3881,N_3882,N_3883,N_3886,N_3887,N_3889,N_3890,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3920,N_3921,N_3922,N_3923,N_3925,N_3928,N_3929,N_3930,N_3932,N_3933,N_3934,N_3935,N_3936,N_3939,N_3940,N_3941,N_3942,N_3944,N_3945,N_3946,N_3948,N_3949,N_3950,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3965,N_3966,N_3967,N_3972,N_3973,N_3974,N_3976,N_3977,N_3978,N_3980,N_3981,N_3982,N_3983,N_3984,N_3986,N_3987,N_3988,N_3989,N_3990,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4001,N_4002,N_4003,N_4004,N_4005,N_4007,N_4009,N_4010,N_4011,N_4012,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4039,N_4040,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4052,N_4053,N_4054,N_4055,N_4056,N_4059,N_4060,N_4063,N_4064,N_4067,N_4070,N_4072,N_4073,N_4074,N_4075,N_4076,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4111,N_4112,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4139,N_4140,N_4141,N_4143,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4153,N_4154,N_4155,N_4156,N_4158,N_4159,N_4160,N_4163,N_4164,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4177,N_4178,N_4179,N_4180,N_4181,N_4183,N_4184,N_4185,N_4186,N_4188,N_4189,N_4190,N_4191,N_4192,N_4194,N_4195,N_4196,N_4197,N_4200,N_4201,N_4202,N_4205,N_4206,N_4207,N_4209,N_4210,N_4211,N_4212,N_4213,N_4215,N_4217,N_4220,N_4221,N_4222,N_4223,N_4226,N_4227,N_4228,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4239,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4252,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4284,N_4285,N_4287,N_4290,N_4291,N_4293,N_4294,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4308,N_4310,N_4311,N_4312,N_4315,N_4316,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4345,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4354,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4366,N_4370,N_4371,N_4372,N_4373,N_4375,N_4376,N_4377,N_4379,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4393,N_4394,N_4395,N_4396,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4410,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4441,N_4443,N_4444,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4455,N_4456,N_4457,N_4460,N_4461,N_4462,N_4463,N_4465,N_4466,N_4469,N_4470,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4480,N_4481,N_4482,N_4484,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4495,N_4497,N_4499,N_4500,N_4501,N_4502,N_4504,N_4505,N_4506,N_4507,N_4510,N_4511,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4534,N_4535,N_4538,N_4539,N_4540,N_4541,N_4542,N_4544,N_4545,N_4546,N_4547,N_4549,N_4550,N_4551,N_4552,N_4554,N_4555,N_4557,N_4558,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4580,N_4581,N_4582,N_4584,N_4585,N_4586,N_4589,N_4591,N_4593,N_4594,N_4595,N_4598,N_4599,N_4601,N_4602,N_4603,N_4605,N_4607,N_4609,N_4612,N_4616,N_4617,N_4618,N_4619,N_4620,N_4622,N_4623,N_4624,N_4625,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4640,N_4641,N_4642,N_4643,N_4644,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4671,N_4672,N_4673,N_4674,N_4675,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4729,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4740,N_4741,N_4742,N_4744,N_4746,N_4747,N_4748,N_4750,N_4751,N_4752,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4764,N_4766,N_4767,N_4768,N_4770,N_4771,N_4773,N_4774,N_4777,N_4779,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4810,N_4812,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4844,N_4845,N_4847,N_4848,N_4849,N_4850,N_4852,N_4854,N_4855,N_4857,N_4858,N_4860,N_4861,N_4862,N_4864,N_4865,N_4867,N_4868,N_4870,N_4871,N_4872,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4881,N_4882,N_4883,N_4884,N_4886,N_4887,N_4890,N_4891,N_4892,N_4893,N_4895,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4925,N_4927,N_4928,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4953,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4963,N_4964,N_4965,N_4966,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4975,N_4978,N_4979,N_4980,N_4982,N_4983,N_4984,N_4985,N_4986,N_4989,N_4990,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_343,In_96);
nor U1 (N_1,In_390,In_404);
or U2 (N_2,In_560,In_428);
nand U3 (N_3,In_97,In_498);
nor U4 (N_4,In_522,In_639);
or U5 (N_5,In_393,In_319);
or U6 (N_6,In_504,In_570);
nor U7 (N_7,In_77,In_188);
xor U8 (N_8,In_241,In_174);
and U9 (N_9,In_274,In_526);
nand U10 (N_10,In_383,In_662);
and U11 (N_11,In_253,In_466);
xor U12 (N_12,In_328,In_746);
nand U13 (N_13,In_537,In_603);
nand U14 (N_14,In_739,In_42);
or U15 (N_15,In_376,In_239);
nor U16 (N_16,In_267,In_304);
xnor U17 (N_17,In_39,In_748);
nand U18 (N_18,In_702,In_622);
nor U19 (N_19,In_184,In_568);
or U20 (N_20,In_501,In_714);
nor U21 (N_21,In_62,In_250);
or U22 (N_22,In_75,In_679);
nand U23 (N_23,In_580,In_332);
or U24 (N_24,In_397,In_337);
xnor U25 (N_25,In_50,In_497);
nor U26 (N_26,In_191,In_690);
xnor U27 (N_27,In_730,In_102);
and U28 (N_28,In_146,In_584);
nand U29 (N_29,In_661,In_152);
xor U30 (N_30,In_516,In_417);
or U31 (N_31,In_104,In_732);
and U32 (N_32,In_557,In_442);
xor U33 (N_33,In_602,In_309);
nor U34 (N_34,In_133,In_43);
nor U35 (N_35,In_57,In_599);
nand U36 (N_36,In_230,In_348);
and U37 (N_37,In_190,In_644);
and U38 (N_38,In_206,In_481);
nor U39 (N_39,In_617,In_694);
nor U40 (N_40,In_699,In_243);
nand U41 (N_41,In_632,In_388);
or U42 (N_42,In_478,In_423);
or U43 (N_43,In_524,In_299);
nor U44 (N_44,In_384,In_727);
and U45 (N_45,In_216,In_704);
and U46 (N_46,In_643,In_60);
and U47 (N_47,In_252,In_31);
nand U48 (N_48,In_717,In_439);
nor U49 (N_49,In_2,In_186);
nor U50 (N_50,In_673,In_605);
xor U51 (N_51,In_531,In_13);
nor U52 (N_52,In_456,In_116);
nand U53 (N_53,In_449,In_483);
and U54 (N_54,In_78,In_346);
xor U55 (N_55,In_322,In_597);
nor U56 (N_56,In_462,In_223);
nor U57 (N_57,In_324,In_467);
xor U58 (N_58,In_113,In_548);
xnor U59 (N_59,In_621,In_36);
and U60 (N_60,In_373,In_619);
nor U61 (N_61,In_203,In_11);
and U62 (N_62,In_364,In_740);
nand U63 (N_63,In_187,In_499);
nand U64 (N_64,In_111,In_436);
or U65 (N_65,In_604,In_251);
nor U66 (N_66,In_294,In_68);
nand U67 (N_67,In_170,In_138);
or U68 (N_68,In_335,In_656);
and U69 (N_69,In_121,In_106);
xnor U70 (N_70,In_189,In_99);
nor U71 (N_71,In_379,In_698);
or U72 (N_72,In_520,In_496);
nor U73 (N_73,In_738,In_264);
or U74 (N_74,In_527,In_173);
xnor U75 (N_75,In_590,In_220);
or U76 (N_76,In_231,In_34);
and U77 (N_77,In_400,In_378);
or U78 (N_78,In_321,In_514);
nor U79 (N_79,In_687,In_678);
nor U80 (N_80,In_674,In_553);
or U81 (N_81,In_547,In_305);
and U82 (N_82,In_244,In_572);
or U83 (N_83,In_443,In_513);
or U84 (N_84,In_192,In_508);
nor U85 (N_85,In_525,In_28);
nor U86 (N_86,In_445,In_544);
xnor U87 (N_87,In_246,In_17);
nor U88 (N_88,In_66,In_433);
or U89 (N_89,In_82,In_281);
and U90 (N_90,In_79,In_144);
xor U91 (N_91,In_161,In_35);
nor U92 (N_92,In_720,In_367);
nand U93 (N_93,In_427,In_49);
or U94 (N_94,In_724,In_726);
nand U95 (N_95,In_598,In_234);
and U96 (N_96,In_616,In_100);
or U97 (N_97,In_405,In_53);
and U98 (N_98,In_519,In_196);
nand U99 (N_99,In_517,In_680);
and U100 (N_100,In_289,In_145);
nor U101 (N_101,In_124,In_539);
nor U102 (N_102,In_625,In_180);
nand U103 (N_103,In_648,In_708);
nand U104 (N_104,In_7,In_256);
or U105 (N_105,In_199,In_705);
nor U106 (N_106,In_471,In_167);
or U107 (N_107,In_683,In_147);
xor U108 (N_108,In_407,In_618);
and U109 (N_109,In_314,In_403);
and U110 (N_110,In_15,In_610);
xor U111 (N_111,In_94,In_394);
or U112 (N_112,In_172,In_26);
or U113 (N_113,In_612,In_658);
or U114 (N_114,In_691,In_503);
nand U115 (N_115,In_464,In_744);
nor U116 (N_116,In_58,In_292);
xor U117 (N_117,In_293,In_511);
nand U118 (N_118,In_391,In_709);
nand U119 (N_119,In_685,In_83);
nand U120 (N_120,In_606,In_255);
nand U121 (N_121,In_95,In_197);
nand U122 (N_122,In_715,In_600);
xor U123 (N_123,In_465,In_723);
nor U124 (N_124,In_472,In_358);
nor U125 (N_125,In_236,In_139);
nand U126 (N_126,In_89,In_453);
nand U127 (N_127,In_578,In_159);
xnor U128 (N_128,In_30,In_582);
xnor U129 (N_129,In_575,In_502);
or U130 (N_130,In_569,In_642);
nor U131 (N_131,In_14,In_81);
and U132 (N_132,In_657,In_178);
or U133 (N_133,In_733,In_312);
nor U134 (N_134,In_19,In_583);
xnor U135 (N_135,In_392,In_608);
xnor U136 (N_136,In_536,In_248);
and U137 (N_137,In_410,In_432);
nor U138 (N_138,In_684,In_668);
xor U139 (N_139,In_596,In_316);
xnor U140 (N_140,In_611,In_463);
or U141 (N_141,In_375,In_47);
or U142 (N_142,In_361,In_207);
nor U143 (N_143,In_490,In_577);
nor U144 (N_144,In_288,In_131);
nand U145 (N_145,In_129,In_412);
or U146 (N_146,In_218,In_22);
xor U147 (N_147,In_117,In_72);
nand U148 (N_148,In_444,In_574);
xnor U149 (N_149,In_438,In_645);
nor U150 (N_150,In_651,In_205);
or U151 (N_151,In_265,In_710);
nand U152 (N_152,In_480,In_385);
and U153 (N_153,In_647,In_226);
nand U154 (N_154,In_655,In_487);
nand U155 (N_155,In_562,In_166);
nor U156 (N_156,In_214,In_719);
xor U157 (N_157,In_512,In_308);
and U158 (N_158,In_576,In_209);
xor U159 (N_159,In_112,In_347);
nor U160 (N_160,In_352,In_46);
and U161 (N_161,In_165,In_283);
and U162 (N_162,In_118,In_493);
xor U163 (N_163,In_195,In_395);
or U164 (N_164,In_374,In_413);
and U165 (N_165,In_136,In_80);
xnor U166 (N_166,In_93,In_185);
xor U167 (N_167,In_132,In_747);
xnor U168 (N_168,In_329,In_105);
nor U169 (N_169,In_148,In_242);
and U170 (N_170,In_201,In_369);
nand U171 (N_171,In_401,In_507);
nor U172 (N_172,In_635,In_98);
xor U173 (N_173,In_317,In_240);
xnor U174 (N_174,In_85,In_424);
or U175 (N_175,In_10,In_182);
and U176 (N_176,In_591,In_276);
nor U177 (N_177,In_224,In_500);
and U178 (N_178,In_1,In_646);
xnor U179 (N_179,In_330,In_273);
or U180 (N_180,In_667,In_0);
nor U181 (N_181,In_71,In_446);
or U182 (N_182,In_441,In_233);
and U183 (N_183,In_725,In_183);
or U184 (N_184,In_212,In_65);
nor U185 (N_185,In_333,In_227);
or U186 (N_186,In_101,In_366);
nor U187 (N_187,In_134,In_495);
nor U188 (N_188,In_415,In_469);
nand U189 (N_189,In_27,In_734);
nand U190 (N_190,In_345,In_713);
nand U191 (N_191,In_677,In_505);
xnor U192 (N_192,In_33,In_566);
nand U193 (N_193,In_545,In_45);
nand U194 (N_194,In_556,In_682);
xor U195 (N_195,In_125,In_636);
nor U196 (N_196,In_592,In_641);
and U197 (N_197,In_671,In_549);
and U198 (N_198,In_198,In_247);
and U199 (N_199,In_235,In_538);
and U200 (N_200,In_84,In_67);
xor U201 (N_201,In_659,In_86);
or U202 (N_202,In_155,In_363);
xnor U203 (N_203,In_425,In_721);
nor U204 (N_204,In_286,In_302);
nor U205 (N_205,In_565,In_204);
xnor U206 (N_206,In_455,In_295);
nor U207 (N_207,In_735,In_8);
or U208 (N_208,In_638,In_257);
nor U209 (N_209,In_399,In_546);
or U210 (N_210,In_601,In_270);
or U211 (N_211,In_181,In_63);
and U212 (N_212,In_551,In_135);
and U213 (N_213,In_620,In_594);
nand U214 (N_214,In_342,In_211);
or U215 (N_215,In_74,In_217);
nand U216 (N_216,In_736,In_381);
xor U217 (N_217,In_411,In_664);
xnor U218 (N_218,In_114,In_126);
and U219 (N_219,In_225,In_540);
and U220 (N_220,In_277,In_108);
or U221 (N_221,In_711,In_589);
or U222 (N_222,In_272,In_269);
or U223 (N_223,In_485,In_238);
and U224 (N_224,In_663,In_567);
nor U225 (N_225,In_326,In_701);
nand U226 (N_226,In_419,In_303);
nor U227 (N_227,In_157,In_169);
xnor U228 (N_228,In_372,In_123);
and U229 (N_229,In_688,In_437);
xor U230 (N_230,In_543,In_630);
and U231 (N_231,In_149,In_676);
and U232 (N_232,In_473,In_115);
nand U233 (N_233,In_362,In_32);
nand U234 (N_234,In_73,In_703);
or U235 (N_235,In_509,In_237);
nor U236 (N_236,In_440,In_581);
and U237 (N_237,In_334,In_588);
nand U238 (N_238,In_731,In_722);
nand U239 (N_239,In_222,In_54);
xor U240 (N_240,In_406,In_450);
nor U241 (N_241,In_629,In_20);
nand U242 (N_242,In_408,In_354);
and U243 (N_243,In_482,In_380);
xnor U244 (N_244,In_491,In_258);
xnor U245 (N_245,In_488,In_128);
nor U246 (N_246,In_349,In_70);
xnor U247 (N_247,In_451,In_414);
nor U248 (N_248,In_282,In_672);
nor U249 (N_249,In_355,In_398);
nand U250 (N_250,In_529,In_494);
nor U251 (N_251,In_16,In_249);
or U252 (N_252,In_586,In_692);
or U253 (N_253,In_542,In_626);
nor U254 (N_254,In_533,In_460);
and U255 (N_255,In_245,In_457);
and U256 (N_256,In_44,In_340);
xor U257 (N_257,In_593,In_595);
xor U258 (N_258,In_142,In_154);
or U259 (N_259,In_541,In_300);
xnor U260 (N_260,In_3,In_229);
nor U261 (N_261,In_175,In_654);
nor U262 (N_262,In_176,In_12);
nor U263 (N_263,In_4,In_103);
xnor U264 (N_264,In_561,In_163);
or U265 (N_265,In_271,In_344);
or U266 (N_266,In_56,In_447);
xnor U267 (N_267,In_696,In_515);
nor U268 (N_268,In_420,In_200);
and U269 (N_269,In_479,In_558);
or U270 (N_270,In_331,In_21);
nand U271 (N_271,In_306,In_554);
nand U272 (N_272,In_634,In_351);
nor U273 (N_273,In_278,In_371);
xor U274 (N_274,In_266,In_37);
nand U275 (N_275,In_215,In_370);
nor U276 (N_276,In_631,In_219);
xor U277 (N_277,In_652,In_728);
nand U278 (N_278,In_448,In_127);
or U279 (N_279,In_458,In_279);
nor U280 (N_280,In_232,In_143);
nor U281 (N_281,In_23,In_649);
and U282 (N_282,In_459,In_61);
and U283 (N_283,In_742,In_164);
nor U284 (N_284,In_486,In_310);
or U285 (N_285,In_76,In_313);
nand U286 (N_286,In_280,In_5);
nor U287 (N_287,In_301,In_29);
nand U288 (N_288,In_359,In_743);
nand U289 (N_289,In_697,In_91);
nor U290 (N_290,In_418,In_559);
xor U291 (N_291,In_311,In_700);
xor U292 (N_292,In_627,In_290);
or U293 (N_293,In_477,In_637);
or U294 (N_294,In_377,In_396);
xnor U295 (N_295,In_429,In_119);
and U296 (N_296,In_51,In_552);
or U297 (N_297,In_357,In_263);
nor U298 (N_298,In_421,In_741);
and U299 (N_299,In_365,In_268);
xnor U300 (N_300,In_338,In_532);
nor U301 (N_301,In_208,In_693);
nor U302 (N_302,In_613,In_523);
or U303 (N_303,In_107,In_528);
or U304 (N_304,In_607,In_609);
or U305 (N_305,In_660,In_535);
nand U306 (N_306,In_402,In_137);
or U307 (N_307,In_262,In_474);
and U308 (N_308,In_284,In_573);
xor U309 (N_309,In_158,In_489);
xor U310 (N_310,In_506,In_275);
nand U311 (N_311,In_615,In_434);
or U312 (N_312,In_261,In_686);
nand U313 (N_313,In_555,In_476);
or U314 (N_314,In_382,In_670);
xor U315 (N_315,In_315,In_130);
and U316 (N_316,In_221,In_475);
or U317 (N_317,In_259,In_210);
and U318 (N_318,In_120,In_454);
xor U319 (N_319,In_325,In_571);
nor U320 (N_320,In_614,In_695);
nand U321 (N_321,In_563,In_153);
and U322 (N_322,In_254,In_534);
nor U323 (N_323,In_296,In_628);
and U324 (N_324,In_323,In_18);
nand U325 (N_325,In_160,In_9);
xnor U326 (N_326,In_387,In_6);
nand U327 (N_327,In_24,In_48);
and U328 (N_328,In_38,In_202);
nand U329 (N_329,In_64,In_162);
and U330 (N_330,In_90,In_177);
nand U331 (N_331,In_297,In_452);
xnor U332 (N_332,In_194,In_422);
or U333 (N_333,In_69,In_665);
nand U334 (N_334,In_287,In_88);
and U335 (N_335,In_470,In_431);
and U336 (N_336,In_52,In_707);
nor U337 (N_337,In_461,In_151);
or U338 (N_338,In_518,In_675);
or U339 (N_339,In_749,In_336);
nand U340 (N_340,In_587,In_681);
nand U341 (N_341,In_468,In_633);
or U342 (N_342,In_92,In_360);
xor U343 (N_343,In_339,In_171);
and U344 (N_344,In_213,In_318);
xnor U345 (N_345,In_298,In_666);
nor U346 (N_346,In_386,In_320);
nor U347 (N_347,In_59,In_55);
or U348 (N_348,In_260,In_745);
or U349 (N_349,In_141,In_737);
xnor U350 (N_350,In_150,In_228);
nor U351 (N_351,In_716,In_623);
xnor U352 (N_352,In_510,In_109);
or U353 (N_353,In_368,In_327);
nand U354 (N_354,In_140,In_356);
nor U355 (N_355,In_712,In_579);
nor U356 (N_356,In_40,In_25);
nor U357 (N_357,In_285,In_350);
nand U358 (N_358,In_291,In_484);
xnor U359 (N_359,In_585,In_168);
and U360 (N_360,In_409,In_307);
and U361 (N_361,In_435,In_156);
xnor U362 (N_362,In_426,In_341);
nor U363 (N_363,In_718,In_87);
or U364 (N_364,In_492,In_669);
or U365 (N_365,In_624,In_416);
and U366 (N_366,In_729,In_530);
nor U367 (N_367,In_193,In_689);
or U368 (N_368,In_389,In_550);
xnor U369 (N_369,In_179,In_706);
or U370 (N_370,In_353,In_640);
nor U371 (N_371,In_122,In_650);
nand U372 (N_372,In_430,In_564);
or U373 (N_373,In_110,In_41);
nor U374 (N_374,In_521,In_653);
and U375 (N_375,In_717,In_657);
and U376 (N_376,In_101,In_257);
nor U377 (N_377,In_95,In_81);
or U378 (N_378,In_20,In_355);
nor U379 (N_379,In_549,In_144);
nor U380 (N_380,In_699,In_587);
or U381 (N_381,In_445,In_80);
nor U382 (N_382,In_604,In_441);
nor U383 (N_383,In_66,In_674);
or U384 (N_384,In_14,In_582);
xnor U385 (N_385,In_219,In_270);
nand U386 (N_386,In_310,In_657);
or U387 (N_387,In_410,In_119);
nor U388 (N_388,In_408,In_208);
or U389 (N_389,In_254,In_440);
nand U390 (N_390,In_544,In_747);
or U391 (N_391,In_234,In_353);
and U392 (N_392,In_418,In_5);
or U393 (N_393,In_219,In_466);
and U394 (N_394,In_526,In_179);
nor U395 (N_395,In_359,In_515);
xnor U396 (N_396,In_203,In_448);
xnor U397 (N_397,In_159,In_633);
or U398 (N_398,In_264,In_182);
nand U399 (N_399,In_361,In_718);
nand U400 (N_400,In_266,In_404);
and U401 (N_401,In_229,In_331);
xnor U402 (N_402,In_263,In_680);
or U403 (N_403,In_227,In_327);
xor U404 (N_404,In_460,In_639);
nand U405 (N_405,In_176,In_590);
nand U406 (N_406,In_203,In_27);
xor U407 (N_407,In_210,In_107);
and U408 (N_408,In_187,In_389);
or U409 (N_409,In_237,In_724);
nor U410 (N_410,In_726,In_85);
nand U411 (N_411,In_0,In_691);
or U412 (N_412,In_109,In_328);
or U413 (N_413,In_725,In_311);
xor U414 (N_414,In_201,In_24);
or U415 (N_415,In_355,In_36);
nor U416 (N_416,In_574,In_118);
nor U417 (N_417,In_327,In_668);
and U418 (N_418,In_352,In_552);
nand U419 (N_419,In_622,In_444);
and U420 (N_420,In_626,In_474);
nor U421 (N_421,In_173,In_668);
nor U422 (N_422,In_660,In_35);
nand U423 (N_423,In_597,In_630);
nor U424 (N_424,In_338,In_55);
nor U425 (N_425,In_334,In_566);
nand U426 (N_426,In_636,In_1);
and U427 (N_427,In_262,In_4);
nor U428 (N_428,In_656,In_269);
xor U429 (N_429,In_691,In_360);
nor U430 (N_430,In_125,In_276);
or U431 (N_431,In_180,In_43);
and U432 (N_432,In_602,In_260);
xnor U433 (N_433,In_423,In_32);
xnor U434 (N_434,In_394,In_475);
nand U435 (N_435,In_58,In_236);
nand U436 (N_436,In_68,In_35);
or U437 (N_437,In_7,In_445);
xnor U438 (N_438,In_377,In_142);
or U439 (N_439,In_219,In_643);
and U440 (N_440,In_600,In_300);
xor U441 (N_441,In_543,In_296);
nand U442 (N_442,In_94,In_325);
nor U443 (N_443,In_529,In_311);
nor U444 (N_444,In_73,In_41);
nand U445 (N_445,In_558,In_601);
nor U446 (N_446,In_546,In_749);
or U447 (N_447,In_52,In_146);
nor U448 (N_448,In_222,In_173);
xnor U449 (N_449,In_224,In_569);
nor U450 (N_450,In_96,In_617);
nand U451 (N_451,In_173,In_555);
xor U452 (N_452,In_743,In_526);
nand U453 (N_453,In_15,In_269);
nor U454 (N_454,In_100,In_635);
and U455 (N_455,In_730,In_395);
and U456 (N_456,In_602,In_600);
nor U457 (N_457,In_567,In_89);
xnor U458 (N_458,In_19,In_45);
nor U459 (N_459,In_196,In_371);
xor U460 (N_460,In_155,In_458);
xor U461 (N_461,In_749,In_488);
xor U462 (N_462,In_440,In_549);
or U463 (N_463,In_76,In_139);
xor U464 (N_464,In_655,In_501);
and U465 (N_465,In_748,In_636);
and U466 (N_466,In_512,In_485);
nand U467 (N_467,In_512,In_168);
and U468 (N_468,In_530,In_264);
nand U469 (N_469,In_544,In_552);
nand U470 (N_470,In_490,In_470);
or U471 (N_471,In_127,In_672);
nand U472 (N_472,In_593,In_612);
nor U473 (N_473,In_141,In_644);
and U474 (N_474,In_444,In_338);
or U475 (N_475,In_51,In_607);
nor U476 (N_476,In_379,In_744);
nor U477 (N_477,In_732,In_182);
or U478 (N_478,In_662,In_326);
nor U479 (N_479,In_658,In_6);
nor U480 (N_480,In_302,In_475);
xnor U481 (N_481,In_487,In_153);
nand U482 (N_482,In_426,In_356);
and U483 (N_483,In_457,In_491);
nor U484 (N_484,In_356,In_52);
or U485 (N_485,In_388,In_405);
or U486 (N_486,In_537,In_136);
nor U487 (N_487,In_688,In_252);
and U488 (N_488,In_34,In_662);
nand U489 (N_489,In_269,In_727);
xnor U490 (N_490,In_578,In_36);
and U491 (N_491,In_283,In_94);
nand U492 (N_492,In_425,In_369);
nand U493 (N_493,In_44,In_14);
nor U494 (N_494,In_701,In_50);
nor U495 (N_495,In_602,In_556);
or U496 (N_496,In_580,In_629);
nand U497 (N_497,In_593,In_178);
xnor U498 (N_498,In_247,In_416);
nand U499 (N_499,In_295,In_410);
nand U500 (N_500,In_115,In_536);
and U501 (N_501,In_473,In_558);
nor U502 (N_502,In_63,In_118);
or U503 (N_503,In_402,In_117);
or U504 (N_504,In_645,In_361);
and U505 (N_505,In_461,In_255);
nand U506 (N_506,In_333,In_576);
and U507 (N_507,In_0,In_420);
nor U508 (N_508,In_574,In_249);
or U509 (N_509,In_38,In_553);
nor U510 (N_510,In_723,In_211);
nand U511 (N_511,In_590,In_336);
or U512 (N_512,In_702,In_377);
or U513 (N_513,In_210,In_483);
nand U514 (N_514,In_298,In_337);
xor U515 (N_515,In_605,In_100);
or U516 (N_516,In_302,In_735);
nand U517 (N_517,In_561,In_660);
nor U518 (N_518,In_407,In_78);
nand U519 (N_519,In_333,In_389);
nand U520 (N_520,In_738,In_490);
xnor U521 (N_521,In_138,In_483);
and U522 (N_522,In_733,In_217);
nor U523 (N_523,In_700,In_674);
nand U524 (N_524,In_631,In_220);
nand U525 (N_525,In_295,In_660);
xnor U526 (N_526,In_727,In_152);
or U527 (N_527,In_370,In_447);
xor U528 (N_528,In_19,In_74);
nor U529 (N_529,In_588,In_545);
or U530 (N_530,In_304,In_265);
and U531 (N_531,In_348,In_642);
xnor U532 (N_532,In_458,In_167);
nand U533 (N_533,In_200,In_359);
nand U534 (N_534,In_444,In_640);
and U535 (N_535,In_504,In_566);
nor U536 (N_536,In_161,In_103);
or U537 (N_537,In_334,In_378);
xnor U538 (N_538,In_415,In_70);
xnor U539 (N_539,In_532,In_495);
nor U540 (N_540,In_129,In_216);
xor U541 (N_541,In_602,In_525);
nor U542 (N_542,In_67,In_310);
or U543 (N_543,In_185,In_39);
nand U544 (N_544,In_464,In_163);
nand U545 (N_545,In_497,In_328);
xor U546 (N_546,In_47,In_377);
nand U547 (N_547,In_623,In_560);
or U548 (N_548,In_14,In_158);
or U549 (N_549,In_111,In_246);
or U550 (N_550,In_14,In_82);
xor U551 (N_551,In_599,In_165);
xor U552 (N_552,In_736,In_178);
or U553 (N_553,In_508,In_278);
nor U554 (N_554,In_564,In_100);
nand U555 (N_555,In_558,In_34);
and U556 (N_556,In_477,In_431);
nand U557 (N_557,In_690,In_543);
nor U558 (N_558,In_309,In_78);
nand U559 (N_559,In_351,In_663);
nor U560 (N_560,In_54,In_256);
xor U561 (N_561,In_663,In_648);
nand U562 (N_562,In_220,In_185);
nand U563 (N_563,In_405,In_571);
nor U564 (N_564,In_377,In_31);
nand U565 (N_565,In_94,In_484);
and U566 (N_566,In_280,In_46);
xnor U567 (N_567,In_106,In_123);
nand U568 (N_568,In_73,In_723);
or U569 (N_569,In_537,In_681);
xor U570 (N_570,In_443,In_99);
nor U571 (N_571,In_383,In_545);
xor U572 (N_572,In_629,In_554);
or U573 (N_573,In_482,In_472);
nor U574 (N_574,In_594,In_103);
xor U575 (N_575,In_490,In_70);
nand U576 (N_576,In_590,In_67);
nor U577 (N_577,In_47,In_686);
nor U578 (N_578,In_456,In_109);
nor U579 (N_579,In_448,In_61);
xnor U580 (N_580,In_676,In_215);
or U581 (N_581,In_7,In_328);
xor U582 (N_582,In_134,In_9);
or U583 (N_583,In_413,In_310);
nor U584 (N_584,In_444,In_14);
nand U585 (N_585,In_532,In_380);
nor U586 (N_586,In_126,In_41);
nand U587 (N_587,In_354,In_512);
nor U588 (N_588,In_99,In_631);
xnor U589 (N_589,In_634,In_256);
xor U590 (N_590,In_153,In_336);
nand U591 (N_591,In_304,In_742);
or U592 (N_592,In_254,In_297);
xor U593 (N_593,In_360,In_602);
nand U594 (N_594,In_144,In_11);
or U595 (N_595,In_170,In_137);
or U596 (N_596,In_74,In_469);
or U597 (N_597,In_687,In_742);
xor U598 (N_598,In_541,In_392);
xnor U599 (N_599,In_248,In_297);
or U600 (N_600,In_602,In_739);
or U601 (N_601,In_435,In_28);
xnor U602 (N_602,In_274,In_501);
or U603 (N_603,In_199,In_480);
and U604 (N_604,In_223,In_434);
nor U605 (N_605,In_407,In_336);
nand U606 (N_606,In_320,In_339);
nor U607 (N_607,In_358,In_443);
xor U608 (N_608,In_158,In_411);
xor U609 (N_609,In_358,In_274);
or U610 (N_610,In_348,In_503);
nand U611 (N_611,In_435,In_241);
nand U612 (N_612,In_729,In_1);
nand U613 (N_613,In_175,In_260);
nor U614 (N_614,In_219,In_111);
xnor U615 (N_615,In_283,In_563);
xor U616 (N_616,In_233,In_72);
nand U617 (N_617,In_722,In_420);
xnor U618 (N_618,In_138,In_726);
and U619 (N_619,In_731,In_698);
nand U620 (N_620,In_53,In_681);
nand U621 (N_621,In_537,In_253);
xnor U622 (N_622,In_696,In_471);
nor U623 (N_623,In_90,In_104);
nor U624 (N_624,In_50,In_77);
or U625 (N_625,In_34,In_284);
nor U626 (N_626,In_531,In_503);
or U627 (N_627,In_9,In_605);
xor U628 (N_628,In_227,In_185);
nor U629 (N_629,In_205,In_581);
and U630 (N_630,In_170,In_464);
xnor U631 (N_631,In_393,In_702);
nand U632 (N_632,In_524,In_610);
nor U633 (N_633,In_655,In_536);
nor U634 (N_634,In_638,In_410);
or U635 (N_635,In_269,In_567);
and U636 (N_636,In_656,In_423);
or U637 (N_637,In_169,In_343);
nand U638 (N_638,In_118,In_346);
or U639 (N_639,In_504,In_639);
nand U640 (N_640,In_356,In_473);
or U641 (N_641,In_339,In_661);
and U642 (N_642,In_301,In_485);
nand U643 (N_643,In_621,In_628);
nor U644 (N_644,In_672,In_101);
nand U645 (N_645,In_359,In_560);
and U646 (N_646,In_317,In_738);
and U647 (N_647,In_627,In_385);
nand U648 (N_648,In_385,In_474);
nand U649 (N_649,In_97,In_81);
xnor U650 (N_650,In_742,In_671);
or U651 (N_651,In_170,In_191);
nor U652 (N_652,In_749,In_413);
nand U653 (N_653,In_198,In_608);
or U654 (N_654,In_129,In_318);
or U655 (N_655,In_557,In_475);
nand U656 (N_656,In_394,In_648);
or U657 (N_657,In_422,In_524);
or U658 (N_658,In_86,In_198);
nor U659 (N_659,In_535,In_19);
nand U660 (N_660,In_374,In_682);
xnor U661 (N_661,In_432,In_592);
or U662 (N_662,In_171,In_518);
nor U663 (N_663,In_412,In_440);
or U664 (N_664,In_181,In_606);
nand U665 (N_665,In_673,In_621);
xnor U666 (N_666,In_173,In_127);
nor U667 (N_667,In_20,In_26);
or U668 (N_668,In_38,In_11);
xor U669 (N_669,In_467,In_209);
and U670 (N_670,In_613,In_410);
or U671 (N_671,In_748,In_541);
or U672 (N_672,In_399,In_15);
nor U673 (N_673,In_548,In_500);
nand U674 (N_674,In_646,In_492);
xnor U675 (N_675,In_131,In_597);
xnor U676 (N_676,In_232,In_1);
and U677 (N_677,In_429,In_668);
and U678 (N_678,In_475,In_241);
xnor U679 (N_679,In_254,In_413);
nor U680 (N_680,In_486,In_199);
nor U681 (N_681,In_67,In_391);
nor U682 (N_682,In_365,In_484);
or U683 (N_683,In_624,In_368);
and U684 (N_684,In_409,In_396);
nor U685 (N_685,In_490,In_308);
nor U686 (N_686,In_236,In_271);
xor U687 (N_687,In_494,In_89);
or U688 (N_688,In_747,In_323);
or U689 (N_689,In_82,In_59);
xor U690 (N_690,In_39,In_238);
nor U691 (N_691,In_648,In_93);
nor U692 (N_692,In_593,In_326);
or U693 (N_693,In_484,In_245);
nand U694 (N_694,In_356,In_674);
nor U695 (N_695,In_140,In_734);
and U696 (N_696,In_427,In_452);
nand U697 (N_697,In_684,In_61);
nand U698 (N_698,In_442,In_144);
nand U699 (N_699,In_20,In_229);
xnor U700 (N_700,In_527,In_295);
nor U701 (N_701,In_105,In_489);
or U702 (N_702,In_585,In_287);
or U703 (N_703,In_138,In_84);
or U704 (N_704,In_65,In_295);
nand U705 (N_705,In_185,In_374);
nand U706 (N_706,In_478,In_208);
xor U707 (N_707,In_649,In_53);
or U708 (N_708,In_23,In_131);
and U709 (N_709,In_132,In_429);
and U710 (N_710,In_432,In_94);
or U711 (N_711,In_568,In_315);
and U712 (N_712,In_661,In_507);
or U713 (N_713,In_700,In_218);
and U714 (N_714,In_649,In_232);
or U715 (N_715,In_728,In_120);
and U716 (N_716,In_105,In_464);
nor U717 (N_717,In_555,In_741);
or U718 (N_718,In_55,In_480);
nor U719 (N_719,In_708,In_733);
xnor U720 (N_720,In_704,In_85);
and U721 (N_721,In_398,In_625);
or U722 (N_722,In_648,In_641);
xnor U723 (N_723,In_545,In_198);
nor U724 (N_724,In_154,In_467);
and U725 (N_725,In_279,In_682);
and U726 (N_726,In_443,In_749);
nor U727 (N_727,In_346,In_742);
or U728 (N_728,In_414,In_661);
or U729 (N_729,In_114,In_600);
and U730 (N_730,In_164,In_466);
xnor U731 (N_731,In_62,In_151);
and U732 (N_732,In_559,In_676);
nor U733 (N_733,In_572,In_447);
nor U734 (N_734,In_47,In_715);
or U735 (N_735,In_310,In_375);
or U736 (N_736,In_335,In_639);
nor U737 (N_737,In_35,In_426);
nand U738 (N_738,In_24,In_714);
xnor U739 (N_739,In_155,In_397);
nand U740 (N_740,In_35,In_92);
nand U741 (N_741,In_458,In_699);
nor U742 (N_742,In_291,In_326);
and U743 (N_743,In_95,In_74);
xor U744 (N_744,In_88,In_274);
and U745 (N_745,In_742,In_275);
xor U746 (N_746,In_62,In_610);
nor U747 (N_747,In_47,In_183);
and U748 (N_748,In_731,In_170);
and U749 (N_749,In_272,In_282);
nor U750 (N_750,In_300,In_559);
or U751 (N_751,In_683,In_717);
nand U752 (N_752,In_99,In_321);
xnor U753 (N_753,In_266,In_488);
nor U754 (N_754,In_655,In_523);
and U755 (N_755,In_507,In_732);
nor U756 (N_756,In_349,In_249);
xnor U757 (N_757,In_338,In_272);
and U758 (N_758,In_562,In_1);
and U759 (N_759,In_321,In_580);
nand U760 (N_760,In_70,In_249);
nand U761 (N_761,In_604,In_576);
nand U762 (N_762,In_693,In_71);
or U763 (N_763,In_21,In_568);
nor U764 (N_764,In_495,In_534);
nand U765 (N_765,In_225,In_359);
xnor U766 (N_766,In_730,In_233);
or U767 (N_767,In_297,In_231);
and U768 (N_768,In_93,In_398);
xor U769 (N_769,In_44,In_525);
nand U770 (N_770,In_696,In_531);
xor U771 (N_771,In_65,In_465);
and U772 (N_772,In_13,In_273);
or U773 (N_773,In_81,In_435);
and U774 (N_774,In_447,In_468);
and U775 (N_775,In_54,In_153);
and U776 (N_776,In_170,In_355);
and U777 (N_777,In_125,In_12);
xnor U778 (N_778,In_88,In_272);
xor U779 (N_779,In_277,In_265);
xnor U780 (N_780,In_476,In_654);
or U781 (N_781,In_633,In_39);
nor U782 (N_782,In_521,In_629);
xnor U783 (N_783,In_272,In_596);
or U784 (N_784,In_569,In_125);
xor U785 (N_785,In_301,In_432);
xor U786 (N_786,In_57,In_0);
or U787 (N_787,In_12,In_73);
xor U788 (N_788,In_638,In_35);
nor U789 (N_789,In_476,In_661);
nand U790 (N_790,In_495,In_196);
nand U791 (N_791,In_412,In_395);
and U792 (N_792,In_31,In_700);
or U793 (N_793,In_551,In_68);
nand U794 (N_794,In_720,In_104);
and U795 (N_795,In_138,In_72);
nor U796 (N_796,In_425,In_661);
or U797 (N_797,In_369,In_450);
xnor U798 (N_798,In_588,In_678);
or U799 (N_799,In_157,In_35);
nor U800 (N_800,In_671,In_229);
xor U801 (N_801,In_467,In_736);
nand U802 (N_802,In_226,In_123);
or U803 (N_803,In_630,In_646);
xor U804 (N_804,In_201,In_50);
xnor U805 (N_805,In_158,In_42);
and U806 (N_806,In_201,In_550);
nand U807 (N_807,In_413,In_115);
nor U808 (N_808,In_462,In_219);
nand U809 (N_809,In_379,In_307);
nor U810 (N_810,In_376,In_563);
nand U811 (N_811,In_265,In_712);
and U812 (N_812,In_706,In_100);
or U813 (N_813,In_133,In_52);
xor U814 (N_814,In_528,In_638);
or U815 (N_815,In_604,In_166);
nor U816 (N_816,In_355,In_270);
and U817 (N_817,In_354,In_394);
xnor U818 (N_818,In_372,In_640);
xnor U819 (N_819,In_549,In_126);
nand U820 (N_820,In_460,In_56);
or U821 (N_821,In_80,In_696);
and U822 (N_822,In_464,In_346);
or U823 (N_823,In_38,In_113);
and U824 (N_824,In_704,In_472);
nand U825 (N_825,In_77,In_346);
nor U826 (N_826,In_285,In_665);
nor U827 (N_827,In_734,In_96);
and U828 (N_828,In_204,In_363);
xnor U829 (N_829,In_159,In_642);
or U830 (N_830,In_527,In_676);
nor U831 (N_831,In_555,In_729);
or U832 (N_832,In_425,In_376);
or U833 (N_833,In_257,In_118);
or U834 (N_834,In_169,In_495);
nand U835 (N_835,In_150,In_627);
or U836 (N_836,In_210,In_672);
or U837 (N_837,In_737,In_365);
or U838 (N_838,In_272,In_695);
or U839 (N_839,In_378,In_89);
or U840 (N_840,In_174,In_231);
nand U841 (N_841,In_144,In_233);
and U842 (N_842,In_745,In_741);
nand U843 (N_843,In_488,In_20);
xnor U844 (N_844,In_684,In_370);
or U845 (N_845,In_126,In_613);
nor U846 (N_846,In_2,In_448);
and U847 (N_847,In_349,In_705);
xor U848 (N_848,In_182,In_659);
nand U849 (N_849,In_52,In_412);
and U850 (N_850,In_500,In_282);
or U851 (N_851,In_258,In_456);
nand U852 (N_852,In_31,In_696);
nor U853 (N_853,In_662,In_371);
xnor U854 (N_854,In_580,In_540);
xor U855 (N_855,In_133,In_670);
or U856 (N_856,In_448,In_250);
nor U857 (N_857,In_355,In_196);
or U858 (N_858,In_418,In_417);
xnor U859 (N_859,In_265,In_223);
nand U860 (N_860,In_391,In_485);
nor U861 (N_861,In_484,In_722);
and U862 (N_862,In_509,In_652);
and U863 (N_863,In_396,In_30);
or U864 (N_864,In_3,In_62);
nand U865 (N_865,In_598,In_241);
nor U866 (N_866,In_473,In_620);
xnor U867 (N_867,In_467,In_268);
and U868 (N_868,In_404,In_183);
nand U869 (N_869,In_257,In_273);
and U870 (N_870,In_447,In_329);
xnor U871 (N_871,In_46,In_385);
xnor U872 (N_872,In_153,In_695);
nand U873 (N_873,In_439,In_104);
or U874 (N_874,In_718,In_120);
and U875 (N_875,In_677,In_666);
and U876 (N_876,In_454,In_679);
nand U877 (N_877,In_185,In_695);
xnor U878 (N_878,In_193,In_69);
and U879 (N_879,In_486,In_79);
and U880 (N_880,In_373,In_202);
or U881 (N_881,In_135,In_136);
nand U882 (N_882,In_202,In_174);
nand U883 (N_883,In_726,In_82);
nor U884 (N_884,In_83,In_143);
nand U885 (N_885,In_372,In_504);
and U886 (N_886,In_540,In_579);
nand U887 (N_887,In_556,In_246);
and U888 (N_888,In_652,In_266);
nand U889 (N_889,In_287,In_279);
or U890 (N_890,In_64,In_747);
nor U891 (N_891,In_729,In_251);
nor U892 (N_892,In_724,In_282);
nor U893 (N_893,In_669,In_144);
or U894 (N_894,In_364,In_725);
xnor U895 (N_895,In_162,In_417);
nor U896 (N_896,In_745,In_10);
xor U897 (N_897,In_424,In_453);
or U898 (N_898,In_113,In_573);
nor U899 (N_899,In_446,In_60);
nor U900 (N_900,In_9,In_348);
xnor U901 (N_901,In_739,In_329);
nor U902 (N_902,In_534,In_563);
and U903 (N_903,In_134,In_402);
or U904 (N_904,In_244,In_371);
xnor U905 (N_905,In_602,In_66);
and U906 (N_906,In_108,In_567);
nor U907 (N_907,In_671,In_731);
xor U908 (N_908,In_616,In_667);
nand U909 (N_909,In_354,In_683);
xor U910 (N_910,In_144,In_626);
nand U911 (N_911,In_174,In_157);
xnor U912 (N_912,In_487,In_72);
or U913 (N_913,In_461,In_580);
or U914 (N_914,In_287,In_465);
nor U915 (N_915,In_440,In_599);
and U916 (N_916,In_187,In_443);
nand U917 (N_917,In_48,In_75);
nor U918 (N_918,In_318,In_283);
or U919 (N_919,In_242,In_388);
or U920 (N_920,In_577,In_536);
or U921 (N_921,In_586,In_428);
nor U922 (N_922,In_622,In_690);
and U923 (N_923,In_246,In_168);
nand U924 (N_924,In_209,In_729);
xor U925 (N_925,In_67,In_527);
xnor U926 (N_926,In_319,In_571);
nor U927 (N_927,In_680,In_471);
nor U928 (N_928,In_70,In_381);
nand U929 (N_929,In_328,In_87);
and U930 (N_930,In_264,In_560);
or U931 (N_931,In_347,In_582);
or U932 (N_932,In_427,In_676);
or U933 (N_933,In_145,In_436);
xnor U934 (N_934,In_717,In_499);
xor U935 (N_935,In_368,In_280);
or U936 (N_936,In_690,In_617);
nand U937 (N_937,In_221,In_286);
and U938 (N_938,In_551,In_685);
nor U939 (N_939,In_480,In_417);
or U940 (N_940,In_384,In_339);
or U941 (N_941,In_453,In_700);
nand U942 (N_942,In_551,In_461);
xnor U943 (N_943,In_1,In_289);
and U944 (N_944,In_364,In_261);
or U945 (N_945,In_472,In_589);
xor U946 (N_946,In_277,In_40);
nand U947 (N_947,In_16,In_78);
nand U948 (N_948,In_235,In_126);
xor U949 (N_949,In_280,In_556);
nor U950 (N_950,In_622,In_434);
nor U951 (N_951,In_688,In_415);
or U952 (N_952,In_284,In_241);
or U953 (N_953,In_163,In_433);
xnor U954 (N_954,In_469,In_122);
and U955 (N_955,In_276,In_449);
nor U956 (N_956,In_694,In_22);
nor U957 (N_957,In_467,In_742);
xor U958 (N_958,In_508,In_276);
nor U959 (N_959,In_615,In_626);
or U960 (N_960,In_206,In_221);
nor U961 (N_961,In_599,In_622);
or U962 (N_962,In_715,In_61);
or U963 (N_963,In_628,In_216);
xnor U964 (N_964,In_225,In_249);
and U965 (N_965,In_524,In_246);
xor U966 (N_966,In_719,In_239);
and U967 (N_967,In_42,In_86);
or U968 (N_968,In_652,In_686);
nand U969 (N_969,In_669,In_653);
nor U970 (N_970,In_582,In_740);
nor U971 (N_971,In_14,In_731);
and U972 (N_972,In_348,In_625);
xnor U973 (N_973,In_70,In_247);
or U974 (N_974,In_286,In_159);
or U975 (N_975,In_457,In_181);
and U976 (N_976,In_50,In_197);
and U977 (N_977,In_350,In_507);
nor U978 (N_978,In_490,In_69);
or U979 (N_979,In_530,In_366);
nand U980 (N_980,In_546,In_612);
nor U981 (N_981,In_336,In_733);
nor U982 (N_982,In_12,In_119);
nand U983 (N_983,In_214,In_667);
nor U984 (N_984,In_22,In_0);
nand U985 (N_985,In_588,In_432);
nand U986 (N_986,In_403,In_509);
or U987 (N_987,In_226,In_132);
xnor U988 (N_988,In_325,In_697);
nor U989 (N_989,In_288,In_279);
nor U990 (N_990,In_685,In_352);
nand U991 (N_991,In_542,In_30);
or U992 (N_992,In_87,In_522);
nand U993 (N_993,In_335,In_432);
or U994 (N_994,In_77,In_236);
nand U995 (N_995,In_598,In_452);
and U996 (N_996,In_235,In_699);
nand U997 (N_997,In_484,In_306);
nor U998 (N_998,In_19,In_683);
nand U999 (N_999,In_286,In_483);
nor U1000 (N_1000,In_529,In_314);
and U1001 (N_1001,In_112,In_581);
nor U1002 (N_1002,In_291,In_366);
or U1003 (N_1003,In_361,In_52);
xor U1004 (N_1004,In_639,In_327);
xnor U1005 (N_1005,In_206,In_121);
nand U1006 (N_1006,In_184,In_587);
nor U1007 (N_1007,In_728,In_209);
nand U1008 (N_1008,In_265,In_733);
nand U1009 (N_1009,In_294,In_246);
and U1010 (N_1010,In_140,In_78);
xor U1011 (N_1011,In_652,In_376);
nand U1012 (N_1012,In_662,In_406);
nor U1013 (N_1013,In_179,In_392);
nand U1014 (N_1014,In_661,In_325);
nor U1015 (N_1015,In_224,In_13);
nor U1016 (N_1016,In_139,In_704);
xnor U1017 (N_1017,In_330,In_391);
xnor U1018 (N_1018,In_370,In_201);
or U1019 (N_1019,In_346,In_17);
and U1020 (N_1020,In_670,In_482);
xnor U1021 (N_1021,In_529,In_115);
or U1022 (N_1022,In_571,In_523);
xor U1023 (N_1023,In_206,In_225);
nor U1024 (N_1024,In_25,In_411);
nor U1025 (N_1025,In_657,In_55);
nand U1026 (N_1026,In_426,In_78);
and U1027 (N_1027,In_720,In_189);
xnor U1028 (N_1028,In_486,In_171);
and U1029 (N_1029,In_231,In_567);
nor U1030 (N_1030,In_448,In_351);
nand U1031 (N_1031,In_261,In_431);
and U1032 (N_1032,In_574,In_229);
nor U1033 (N_1033,In_687,In_178);
and U1034 (N_1034,In_517,In_327);
nand U1035 (N_1035,In_331,In_44);
or U1036 (N_1036,In_135,In_587);
or U1037 (N_1037,In_169,In_706);
nand U1038 (N_1038,In_501,In_725);
nor U1039 (N_1039,In_499,In_157);
nor U1040 (N_1040,In_460,In_406);
nand U1041 (N_1041,In_511,In_30);
nor U1042 (N_1042,In_725,In_43);
nand U1043 (N_1043,In_138,In_206);
xor U1044 (N_1044,In_255,In_714);
and U1045 (N_1045,In_273,In_200);
and U1046 (N_1046,In_299,In_177);
nand U1047 (N_1047,In_525,In_434);
and U1048 (N_1048,In_198,In_507);
nand U1049 (N_1049,In_385,In_47);
and U1050 (N_1050,In_486,In_513);
and U1051 (N_1051,In_615,In_127);
nor U1052 (N_1052,In_148,In_436);
nand U1053 (N_1053,In_121,In_445);
xnor U1054 (N_1054,In_463,In_609);
nor U1055 (N_1055,In_528,In_227);
xor U1056 (N_1056,In_555,In_376);
or U1057 (N_1057,In_427,In_503);
nor U1058 (N_1058,In_708,In_256);
nand U1059 (N_1059,In_477,In_436);
nor U1060 (N_1060,In_572,In_517);
or U1061 (N_1061,In_437,In_665);
xor U1062 (N_1062,In_129,In_639);
and U1063 (N_1063,In_627,In_544);
or U1064 (N_1064,In_353,In_319);
nand U1065 (N_1065,In_196,In_132);
nand U1066 (N_1066,In_324,In_116);
nor U1067 (N_1067,In_47,In_436);
and U1068 (N_1068,In_163,In_603);
xnor U1069 (N_1069,In_40,In_678);
nor U1070 (N_1070,In_102,In_260);
and U1071 (N_1071,In_635,In_217);
nand U1072 (N_1072,In_286,In_530);
or U1073 (N_1073,In_95,In_86);
and U1074 (N_1074,In_476,In_511);
xor U1075 (N_1075,In_579,In_206);
or U1076 (N_1076,In_136,In_236);
nand U1077 (N_1077,In_557,In_574);
and U1078 (N_1078,In_508,In_154);
nand U1079 (N_1079,In_693,In_702);
nor U1080 (N_1080,In_130,In_8);
nand U1081 (N_1081,In_65,In_619);
nor U1082 (N_1082,In_533,In_568);
nor U1083 (N_1083,In_66,In_103);
nand U1084 (N_1084,In_316,In_197);
nor U1085 (N_1085,In_19,In_194);
nand U1086 (N_1086,In_583,In_422);
or U1087 (N_1087,In_745,In_105);
xnor U1088 (N_1088,In_113,In_571);
and U1089 (N_1089,In_273,In_466);
xor U1090 (N_1090,In_56,In_164);
xnor U1091 (N_1091,In_404,In_405);
nor U1092 (N_1092,In_588,In_711);
and U1093 (N_1093,In_577,In_96);
and U1094 (N_1094,In_667,In_338);
and U1095 (N_1095,In_377,In_663);
or U1096 (N_1096,In_220,In_46);
xor U1097 (N_1097,In_733,In_690);
and U1098 (N_1098,In_487,In_351);
xor U1099 (N_1099,In_267,In_371);
xor U1100 (N_1100,In_470,In_17);
nand U1101 (N_1101,In_246,In_55);
xnor U1102 (N_1102,In_213,In_269);
nor U1103 (N_1103,In_31,In_408);
xnor U1104 (N_1104,In_445,In_428);
nand U1105 (N_1105,In_531,In_42);
nor U1106 (N_1106,In_103,In_584);
xor U1107 (N_1107,In_427,In_596);
nand U1108 (N_1108,In_13,In_716);
nor U1109 (N_1109,In_624,In_583);
xor U1110 (N_1110,In_384,In_263);
and U1111 (N_1111,In_443,In_58);
xor U1112 (N_1112,In_143,In_489);
or U1113 (N_1113,In_650,In_102);
xnor U1114 (N_1114,In_492,In_82);
nor U1115 (N_1115,In_86,In_269);
or U1116 (N_1116,In_415,In_276);
and U1117 (N_1117,In_201,In_191);
nand U1118 (N_1118,In_448,In_211);
nand U1119 (N_1119,In_213,In_742);
and U1120 (N_1120,In_419,In_215);
or U1121 (N_1121,In_179,In_91);
xor U1122 (N_1122,In_516,In_105);
nand U1123 (N_1123,In_85,In_357);
xnor U1124 (N_1124,In_207,In_153);
nor U1125 (N_1125,In_733,In_634);
or U1126 (N_1126,In_165,In_616);
and U1127 (N_1127,In_614,In_203);
xnor U1128 (N_1128,In_656,In_516);
xor U1129 (N_1129,In_24,In_545);
nand U1130 (N_1130,In_421,In_475);
nor U1131 (N_1131,In_62,In_7);
nand U1132 (N_1132,In_363,In_573);
nor U1133 (N_1133,In_105,In_692);
and U1134 (N_1134,In_160,In_432);
and U1135 (N_1135,In_682,In_175);
nand U1136 (N_1136,In_523,In_740);
nand U1137 (N_1137,In_576,In_664);
or U1138 (N_1138,In_439,In_76);
nor U1139 (N_1139,In_329,In_207);
xnor U1140 (N_1140,In_447,In_186);
xnor U1141 (N_1141,In_584,In_716);
or U1142 (N_1142,In_552,In_492);
and U1143 (N_1143,In_343,In_110);
or U1144 (N_1144,In_516,In_282);
or U1145 (N_1145,In_159,In_445);
and U1146 (N_1146,In_241,In_647);
or U1147 (N_1147,In_644,In_270);
and U1148 (N_1148,In_128,In_374);
nand U1149 (N_1149,In_485,In_118);
xnor U1150 (N_1150,In_574,In_119);
nand U1151 (N_1151,In_267,In_550);
and U1152 (N_1152,In_120,In_573);
nand U1153 (N_1153,In_310,In_255);
xor U1154 (N_1154,In_534,In_443);
nand U1155 (N_1155,In_298,In_321);
nand U1156 (N_1156,In_560,In_10);
nand U1157 (N_1157,In_458,In_160);
nand U1158 (N_1158,In_730,In_474);
or U1159 (N_1159,In_595,In_508);
or U1160 (N_1160,In_719,In_617);
nand U1161 (N_1161,In_514,In_546);
xnor U1162 (N_1162,In_493,In_655);
and U1163 (N_1163,In_521,In_528);
and U1164 (N_1164,In_469,In_221);
and U1165 (N_1165,In_731,In_342);
and U1166 (N_1166,In_649,In_30);
xnor U1167 (N_1167,In_749,In_423);
and U1168 (N_1168,In_741,In_346);
and U1169 (N_1169,In_67,In_272);
and U1170 (N_1170,In_498,In_473);
and U1171 (N_1171,In_603,In_635);
nor U1172 (N_1172,In_746,In_196);
nand U1173 (N_1173,In_255,In_272);
and U1174 (N_1174,In_79,In_440);
or U1175 (N_1175,In_139,In_285);
xnor U1176 (N_1176,In_40,In_721);
nor U1177 (N_1177,In_278,In_651);
nand U1178 (N_1178,In_18,In_452);
or U1179 (N_1179,In_453,In_440);
nor U1180 (N_1180,In_346,In_59);
xor U1181 (N_1181,In_604,In_519);
or U1182 (N_1182,In_501,In_645);
nand U1183 (N_1183,In_233,In_642);
nor U1184 (N_1184,In_17,In_51);
nor U1185 (N_1185,In_662,In_55);
xor U1186 (N_1186,In_381,In_40);
or U1187 (N_1187,In_543,In_3);
xnor U1188 (N_1188,In_645,In_406);
nor U1189 (N_1189,In_699,In_485);
nand U1190 (N_1190,In_393,In_245);
xor U1191 (N_1191,In_162,In_531);
nand U1192 (N_1192,In_352,In_140);
or U1193 (N_1193,In_222,In_336);
nor U1194 (N_1194,In_473,In_694);
nand U1195 (N_1195,In_299,In_477);
xnor U1196 (N_1196,In_362,In_158);
nand U1197 (N_1197,In_577,In_411);
xnor U1198 (N_1198,In_165,In_187);
or U1199 (N_1199,In_503,In_50);
or U1200 (N_1200,In_675,In_447);
nand U1201 (N_1201,In_119,In_582);
xnor U1202 (N_1202,In_188,In_692);
or U1203 (N_1203,In_216,In_656);
nor U1204 (N_1204,In_360,In_195);
xor U1205 (N_1205,In_303,In_610);
or U1206 (N_1206,In_657,In_659);
or U1207 (N_1207,In_272,In_687);
xnor U1208 (N_1208,In_579,In_24);
and U1209 (N_1209,In_673,In_512);
xnor U1210 (N_1210,In_96,In_73);
nand U1211 (N_1211,In_293,In_278);
nor U1212 (N_1212,In_67,In_732);
and U1213 (N_1213,In_545,In_527);
or U1214 (N_1214,In_252,In_410);
or U1215 (N_1215,In_535,In_733);
nand U1216 (N_1216,In_323,In_177);
nand U1217 (N_1217,In_321,In_693);
nor U1218 (N_1218,In_152,In_518);
or U1219 (N_1219,In_90,In_195);
or U1220 (N_1220,In_601,In_479);
or U1221 (N_1221,In_184,In_444);
xor U1222 (N_1222,In_82,In_571);
or U1223 (N_1223,In_563,In_282);
xor U1224 (N_1224,In_150,In_563);
or U1225 (N_1225,In_329,In_161);
and U1226 (N_1226,In_451,In_203);
nor U1227 (N_1227,In_696,In_170);
nand U1228 (N_1228,In_725,In_570);
and U1229 (N_1229,In_189,In_85);
or U1230 (N_1230,In_143,In_275);
and U1231 (N_1231,In_583,In_607);
or U1232 (N_1232,In_587,In_276);
or U1233 (N_1233,In_580,In_645);
and U1234 (N_1234,In_321,In_665);
or U1235 (N_1235,In_576,In_504);
or U1236 (N_1236,In_455,In_712);
and U1237 (N_1237,In_41,In_49);
or U1238 (N_1238,In_95,In_12);
or U1239 (N_1239,In_566,In_238);
nand U1240 (N_1240,In_371,In_139);
or U1241 (N_1241,In_486,In_108);
xor U1242 (N_1242,In_404,In_715);
nor U1243 (N_1243,In_326,In_605);
nand U1244 (N_1244,In_478,In_3);
or U1245 (N_1245,In_415,In_369);
and U1246 (N_1246,In_244,In_337);
nor U1247 (N_1247,In_232,In_577);
xor U1248 (N_1248,In_106,In_481);
nand U1249 (N_1249,In_280,In_113);
nand U1250 (N_1250,In_406,In_432);
or U1251 (N_1251,In_696,In_680);
xnor U1252 (N_1252,In_59,In_180);
and U1253 (N_1253,In_249,In_298);
or U1254 (N_1254,In_684,In_120);
and U1255 (N_1255,In_143,In_736);
or U1256 (N_1256,In_132,In_145);
or U1257 (N_1257,In_746,In_229);
or U1258 (N_1258,In_248,In_235);
or U1259 (N_1259,In_459,In_692);
nand U1260 (N_1260,In_355,In_675);
or U1261 (N_1261,In_310,In_615);
nor U1262 (N_1262,In_463,In_329);
xor U1263 (N_1263,In_659,In_602);
nor U1264 (N_1264,In_163,In_418);
and U1265 (N_1265,In_19,In_97);
xnor U1266 (N_1266,In_503,In_290);
and U1267 (N_1267,In_410,In_266);
nand U1268 (N_1268,In_683,In_595);
xnor U1269 (N_1269,In_34,In_494);
and U1270 (N_1270,In_123,In_197);
nand U1271 (N_1271,In_361,In_455);
nand U1272 (N_1272,In_305,In_340);
nand U1273 (N_1273,In_463,In_280);
nor U1274 (N_1274,In_436,In_549);
nand U1275 (N_1275,In_285,In_695);
or U1276 (N_1276,In_544,In_174);
xnor U1277 (N_1277,In_234,In_167);
nor U1278 (N_1278,In_729,In_166);
or U1279 (N_1279,In_178,In_56);
xnor U1280 (N_1280,In_311,In_211);
or U1281 (N_1281,In_343,In_591);
nor U1282 (N_1282,In_374,In_317);
and U1283 (N_1283,In_573,In_615);
or U1284 (N_1284,In_443,In_318);
nor U1285 (N_1285,In_249,In_67);
xor U1286 (N_1286,In_412,In_58);
nor U1287 (N_1287,In_436,In_459);
nor U1288 (N_1288,In_657,In_554);
nand U1289 (N_1289,In_277,In_239);
nand U1290 (N_1290,In_623,In_55);
or U1291 (N_1291,In_91,In_674);
or U1292 (N_1292,In_47,In_693);
nand U1293 (N_1293,In_375,In_323);
nor U1294 (N_1294,In_288,In_678);
xnor U1295 (N_1295,In_548,In_250);
or U1296 (N_1296,In_722,In_499);
nor U1297 (N_1297,In_744,In_4);
or U1298 (N_1298,In_733,In_311);
nand U1299 (N_1299,In_475,In_52);
xor U1300 (N_1300,In_218,In_482);
or U1301 (N_1301,In_229,In_139);
or U1302 (N_1302,In_266,In_51);
nor U1303 (N_1303,In_373,In_642);
xnor U1304 (N_1304,In_528,In_425);
and U1305 (N_1305,In_2,In_232);
or U1306 (N_1306,In_398,In_718);
or U1307 (N_1307,In_226,In_355);
nor U1308 (N_1308,In_633,In_95);
xor U1309 (N_1309,In_201,In_738);
or U1310 (N_1310,In_626,In_699);
nand U1311 (N_1311,In_394,In_290);
nand U1312 (N_1312,In_590,In_95);
and U1313 (N_1313,In_160,In_83);
and U1314 (N_1314,In_550,In_252);
or U1315 (N_1315,In_731,In_673);
xor U1316 (N_1316,In_185,In_497);
and U1317 (N_1317,In_447,In_217);
or U1318 (N_1318,In_137,In_246);
or U1319 (N_1319,In_27,In_635);
nor U1320 (N_1320,In_185,In_103);
nor U1321 (N_1321,In_352,In_171);
or U1322 (N_1322,In_348,In_727);
and U1323 (N_1323,In_343,In_75);
xnor U1324 (N_1324,In_451,In_723);
nor U1325 (N_1325,In_163,In_683);
xor U1326 (N_1326,In_648,In_554);
nand U1327 (N_1327,In_618,In_281);
nor U1328 (N_1328,In_301,In_398);
xor U1329 (N_1329,In_349,In_732);
nand U1330 (N_1330,In_383,In_666);
xnor U1331 (N_1331,In_378,In_377);
or U1332 (N_1332,In_330,In_590);
nand U1333 (N_1333,In_287,In_516);
nor U1334 (N_1334,In_452,In_614);
nor U1335 (N_1335,In_389,In_313);
xor U1336 (N_1336,In_381,In_601);
or U1337 (N_1337,In_365,In_445);
nand U1338 (N_1338,In_596,In_255);
nand U1339 (N_1339,In_618,In_426);
nand U1340 (N_1340,In_261,In_483);
nor U1341 (N_1341,In_425,In_717);
xnor U1342 (N_1342,In_404,In_378);
xnor U1343 (N_1343,In_631,In_693);
nand U1344 (N_1344,In_293,In_193);
or U1345 (N_1345,In_691,In_580);
nand U1346 (N_1346,In_234,In_349);
xor U1347 (N_1347,In_170,In_78);
nor U1348 (N_1348,In_694,In_403);
nand U1349 (N_1349,In_634,In_251);
or U1350 (N_1350,In_208,In_260);
or U1351 (N_1351,In_268,In_492);
nor U1352 (N_1352,In_610,In_311);
xor U1353 (N_1353,In_467,In_615);
nand U1354 (N_1354,In_638,In_405);
xnor U1355 (N_1355,In_182,In_231);
nand U1356 (N_1356,In_229,In_500);
nor U1357 (N_1357,In_544,In_545);
nand U1358 (N_1358,In_647,In_339);
xor U1359 (N_1359,In_330,In_287);
xnor U1360 (N_1360,In_194,In_22);
nor U1361 (N_1361,In_351,In_707);
nor U1362 (N_1362,In_739,In_735);
and U1363 (N_1363,In_208,In_467);
or U1364 (N_1364,In_60,In_163);
nand U1365 (N_1365,In_556,In_135);
xnor U1366 (N_1366,In_395,In_494);
nand U1367 (N_1367,In_87,In_461);
nand U1368 (N_1368,In_539,In_449);
or U1369 (N_1369,In_590,In_245);
nor U1370 (N_1370,In_612,In_731);
nand U1371 (N_1371,In_233,In_528);
and U1372 (N_1372,In_535,In_147);
xnor U1373 (N_1373,In_5,In_406);
and U1374 (N_1374,In_467,In_179);
xor U1375 (N_1375,In_238,In_516);
nor U1376 (N_1376,In_551,In_431);
or U1377 (N_1377,In_737,In_591);
xor U1378 (N_1378,In_557,In_317);
or U1379 (N_1379,In_448,In_143);
and U1380 (N_1380,In_137,In_292);
nand U1381 (N_1381,In_412,In_209);
nor U1382 (N_1382,In_612,In_332);
and U1383 (N_1383,In_245,In_9);
nand U1384 (N_1384,In_648,In_144);
nand U1385 (N_1385,In_594,In_494);
nand U1386 (N_1386,In_440,In_723);
nor U1387 (N_1387,In_88,In_524);
or U1388 (N_1388,In_233,In_383);
nand U1389 (N_1389,In_79,In_550);
and U1390 (N_1390,In_62,In_564);
nand U1391 (N_1391,In_374,In_625);
or U1392 (N_1392,In_738,In_609);
nand U1393 (N_1393,In_202,In_77);
and U1394 (N_1394,In_648,In_660);
xor U1395 (N_1395,In_632,In_494);
xnor U1396 (N_1396,In_683,In_104);
xnor U1397 (N_1397,In_632,In_558);
or U1398 (N_1398,In_608,In_220);
and U1399 (N_1399,In_468,In_749);
nand U1400 (N_1400,In_104,In_417);
and U1401 (N_1401,In_550,In_285);
nor U1402 (N_1402,In_66,In_280);
nor U1403 (N_1403,In_315,In_577);
and U1404 (N_1404,In_635,In_106);
or U1405 (N_1405,In_383,In_649);
xnor U1406 (N_1406,In_638,In_451);
or U1407 (N_1407,In_126,In_523);
nor U1408 (N_1408,In_191,In_413);
or U1409 (N_1409,In_357,In_411);
or U1410 (N_1410,In_598,In_632);
nor U1411 (N_1411,In_89,In_563);
xor U1412 (N_1412,In_655,In_733);
or U1413 (N_1413,In_496,In_431);
or U1414 (N_1414,In_692,In_425);
and U1415 (N_1415,In_104,In_412);
and U1416 (N_1416,In_46,In_66);
and U1417 (N_1417,In_636,In_489);
xor U1418 (N_1418,In_246,In_157);
and U1419 (N_1419,In_659,In_311);
nor U1420 (N_1420,In_365,In_615);
or U1421 (N_1421,In_735,In_139);
nand U1422 (N_1422,In_403,In_384);
xnor U1423 (N_1423,In_356,In_491);
and U1424 (N_1424,In_312,In_87);
xor U1425 (N_1425,In_33,In_340);
or U1426 (N_1426,In_466,In_63);
nand U1427 (N_1427,In_178,In_253);
nand U1428 (N_1428,In_400,In_710);
xor U1429 (N_1429,In_295,In_323);
and U1430 (N_1430,In_628,In_686);
and U1431 (N_1431,In_34,In_155);
nand U1432 (N_1432,In_595,In_583);
or U1433 (N_1433,In_95,In_717);
nand U1434 (N_1434,In_744,In_214);
and U1435 (N_1435,In_736,In_257);
nor U1436 (N_1436,In_355,In_14);
and U1437 (N_1437,In_325,In_411);
and U1438 (N_1438,In_455,In_414);
nand U1439 (N_1439,In_372,In_79);
xnor U1440 (N_1440,In_185,In_180);
nand U1441 (N_1441,In_459,In_428);
nand U1442 (N_1442,In_405,In_570);
xor U1443 (N_1443,In_118,In_739);
nor U1444 (N_1444,In_72,In_463);
xor U1445 (N_1445,In_353,In_193);
nand U1446 (N_1446,In_53,In_116);
xor U1447 (N_1447,In_539,In_509);
or U1448 (N_1448,In_614,In_94);
xnor U1449 (N_1449,In_288,In_295);
nor U1450 (N_1450,In_652,In_118);
or U1451 (N_1451,In_411,In_484);
and U1452 (N_1452,In_295,In_166);
nand U1453 (N_1453,In_156,In_63);
or U1454 (N_1454,In_594,In_334);
nor U1455 (N_1455,In_98,In_247);
xnor U1456 (N_1456,In_10,In_214);
and U1457 (N_1457,In_205,In_304);
xor U1458 (N_1458,In_578,In_344);
nor U1459 (N_1459,In_513,In_714);
nand U1460 (N_1460,In_117,In_480);
nor U1461 (N_1461,In_128,In_725);
xor U1462 (N_1462,In_632,In_523);
or U1463 (N_1463,In_604,In_210);
xor U1464 (N_1464,In_315,In_676);
xor U1465 (N_1465,In_349,In_402);
nor U1466 (N_1466,In_18,In_670);
or U1467 (N_1467,In_621,In_181);
and U1468 (N_1468,In_560,In_409);
xnor U1469 (N_1469,In_538,In_683);
xor U1470 (N_1470,In_335,In_600);
and U1471 (N_1471,In_25,In_621);
nand U1472 (N_1472,In_692,In_667);
nor U1473 (N_1473,In_236,In_408);
nand U1474 (N_1474,In_682,In_244);
or U1475 (N_1475,In_253,In_732);
nor U1476 (N_1476,In_511,In_557);
and U1477 (N_1477,In_80,In_78);
and U1478 (N_1478,In_357,In_313);
and U1479 (N_1479,In_25,In_261);
nor U1480 (N_1480,In_563,In_614);
nand U1481 (N_1481,In_442,In_741);
xor U1482 (N_1482,In_663,In_338);
xor U1483 (N_1483,In_296,In_548);
and U1484 (N_1484,In_188,In_276);
or U1485 (N_1485,In_547,In_206);
or U1486 (N_1486,In_345,In_440);
and U1487 (N_1487,In_385,In_405);
and U1488 (N_1488,In_454,In_18);
or U1489 (N_1489,In_410,In_471);
nor U1490 (N_1490,In_477,In_290);
or U1491 (N_1491,In_736,In_316);
and U1492 (N_1492,In_637,In_434);
or U1493 (N_1493,In_642,In_421);
or U1494 (N_1494,In_82,In_560);
nor U1495 (N_1495,In_500,In_92);
and U1496 (N_1496,In_465,In_319);
or U1497 (N_1497,In_585,In_173);
or U1498 (N_1498,In_29,In_197);
nor U1499 (N_1499,In_169,In_524);
or U1500 (N_1500,In_271,In_246);
nor U1501 (N_1501,In_683,In_314);
nand U1502 (N_1502,In_564,In_461);
and U1503 (N_1503,In_541,In_405);
and U1504 (N_1504,In_252,In_197);
or U1505 (N_1505,In_357,In_676);
and U1506 (N_1506,In_341,In_354);
xor U1507 (N_1507,In_480,In_251);
nand U1508 (N_1508,In_486,In_429);
nand U1509 (N_1509,In_81,In_190);
nor U1510 (N_1510,In_619,In_289);
nand U1511 (N_1511,In_238,In_732);
or U1512 (N_1512,In_473,In_385);
or U1513 (N_1513,In_517,In_693);
nand U1514 (N_1514,In_642,In_742);
xor U1515 (N_1515,In_689,In_17);
nand U1516 (N_1516,In_293,In_173);
xnor U1517 (N_1517,In_397,In_744);
xnor U1518 (N_1518,In_371,In_345);
nand U1519 (N_1519,In_733,In_615);
nor U1520 (N_1520,In_213,In_384);
or U1521 (N_1521,In_84,In_498);
nor U1522 (N_1522,In_308,In_160);
nor U1523 (N_1523,In_330,In_525);
xor U1524 (N_1524,In_335,In_518);
nor U1525 (N_1525,In_542,In_393);
or U1526 (N_1526,In_5,In_543);
xor U1527 (N_1527,In_470,In_262);
xor U1528 (N_1528,In_548,In_538);
nor U1529 (N_1529,In_517,In_527);
or U1530 (N_1530,In_558,In_648);
and U1531 (N_1531,In_200,In_324);
xnor U1532 (N_1532,In_183,In_384);
xor U1533 (N_1533,In_524,In_727);
or U1534 (N_1534,In_4,In_471);
nand U1535 (N_1535,In_376,In_100);
or U1536 (N_1536,In_715,In_717);
nor U1537 (N_1537,In_209,In_268);
nor U1538 (N_1538,In_522,In_389);
nand U1539 (N_1539,In_142,In_132);
and U1540 (N_1540,In_588,In_385);
and U1541 (N_1541,In_125,In_156);
or U1542 (N_1542,In_17,In_685);
xnor U1543 (N_1543,In_462,In_191);
or U1544 (N_1544,In_586,In_138);
and U1545 (N_1545,In_536,In_75);
nand U1546 (N_1546,In_295,In_281);
nor U1547 (N_1547,In_171,In_236);
nor U1548 (N_1548,In_396,In_37);
nor U1549 (N_1549,In_19,In_38);
and U1550 (N_1550,In_722,In_634);
xor U1551 (N_1551,In_400,In_419);
nor U1552 (N_1552,In_388,In_271);
xnor U1553 (N_1553,In_14,In_675);
or U1554 (N_1554,In_613,In_690);
and U1555 (N_1555,In_684,In_86);
or U1556 (N_1556,In_72,In_289);
and U1557 (N_1557,In_551,In_405);
nor U1558 (N_1558,In_625,In_605);
xor U1559 (N_1559,In_278,In_568);
xor U1560 (N_1560,In_372,In_665);
xor U1561 (N_1561,In_11,In_719);
and U1562 (N_1562,In_82,In_200);
xnor U1563 (N_1563,In_324,In_711);
nor U1564 (N_1564,In_181,In_450);
or U1565 (N_1565,In_604,In_195);
and U1566 (N_1566,In_713,In_85);
or U1567 (N_1567,In_636,In_697);
or U1568 (N_1568,In_340,In_106);
nand U1569 (N_1569,In_324,In_288);
xor U1570 (N_1570,In_127,In_208);
nor U1571 (N_1571,In_83,In_349);
and U1572 (N_1572,In_406,In_373);
xor U1573 (N_1573,In_437,In_606);
and U1574 (N_1574,In_519,In_726);
nand U1575 (N_1575,In_131,In_293);
or U1576 (N_1576,In_25,In_648);
xor U1577 (N_1577,In_115,In_434);
xor U1578 (N_1578,In_555,In_166);
and U1579 (N_1579,In_86,In_494);
or U1580 (N_1580,In_188,In_702);
or U1581 (N_1581,In_213,In_351);
nor U1582 (N_1582,In_730,In_654);
and U1583 (N_1583,In_107,In_382);
nand U1584 (N_1584,In_748,In_728);
or U1585 (N_1585,In_496,In_19);
xnor U1586 (N_1586,In_540,In_261);
nor U1587 (N_1587,In_290,In_517);
nor U1588 (N_1588,In_741,In_124);
xor U1589 (N_1589,In_185,In_237);
or U1590 (N_1590,In_220,In_432);
xor U1591 (N_1591,In_88,In_530);
or U1592 (N_1592,In_149,In_437);
and U1593 (N_1593,In_117,In_399);
nand U1594 (N_1594,In_274,In_451);
xnor U1595 (N_1595,In_8,In_261);
xor U1596 (N_1596,In_421,In_439);
nor U1597 (N_1597,In_441,In_227);
xor U1598 (N_1598,In_722,In_53);
xnor U1599 (N_1599,In_408,In_685);
and U1600 (N_1600,In_533,In_118);
nand U1601 (N_1601,In_576,In_676);
nand U1602 (N_1602,In_120,In_509);
or U1603 (N_1603,In_174,In_357);
xor U1604 (N_1604,In_727,In_580);
or U1605 (N_1605,In_514,In_224);
xor U1606 (N_1606,In_467,In_452);
and U1607 (N_1607,In_432,In_386);
or U1608 (N_1608,In_737,In_298);
nand U1609 (N_1609,In_207,In_282);
and U1610 (N_1610,In_178,In_61);
nand U1611 (N_1611,In_128,In_698);
nand U1612 (N_1612,In_458,In_156);
nor U1613 (N_1613,In_568,In_386);
and U1614 (N_1614,In_482,In_595);
or U1615 (N_1615,In_26,In_112);
xnor U1616 (N_1616,In_681,In_366);
or U1617 (N_1617,In_317,In_191);
nor U1618 (N_1618,In_472,In_136);
nor U1619 (N_1619,In_728,In_338);
or U1620 (N_1620,In_462,In_702);
and U1621 (N_1621,In_737,In_12);
xnor U1622 (N_1622,In_485,In_744);
or U1623 (N_1623,In_678,In_280);
and U1624 (N_1624,In_351,In_540);
or U1625 (N_1625,In_112,In_651);
xor U1626 (N_1626,In_294,In_463);
nand U1627 (N_1627,In_178,In_17);
xnor U1628 (N_1628,In_80,In_526);
and U1629 (N_1629,In_588,In_736);
or U1630 (N_1630,In_660,In_70);
nor U1631 (N_1631,In_444,In_591);
or U1632 (N_1632,In_251,In_625);
or U1633 (N_1633,In_533,In_347);
nor U1634 (N_1634,In_352,In_714);
xnor U1635 (N_1635,In_538,In_298);
or U1636 (N_1636,In_299,In_696);
and U1637 (N_1637,In_297,In_600);
or U1638 (N_1638,In_709,In_57);
and U1639 (N_1639,In_266,In_589);
nor U1640 (N_1640,In_232,In_215);
or U1641 (N_1641,In_683,In_224);
nand U1642 (N_1642,In_70,In_4);
nor U1643 (N_1643,In_177,In_375);
nand U1644 (N_1644,In_641,In_203);
xor U1645 (N_1645,In_431,In_394);
nor U1646 (N_1646,In_509,In_117);
and U1647 (N_1647,In_76,In_56);
nand U1648 (N_1648,In_565,In_148);
and U1649 (N_1649,In_328,In_563);
and U1650 (N_1650,In_45,In_435);
or U1651 (N_1651,In_493,In_351);
nor U1652 (N_1652,In_149,In_340);
nor U1653 (N_1653,In_557,In_509);
xnor U1654 (N_1654,In_262,In_93);
or U1655 (N_1655,In_147,In_375);
nor U1656 (N_1656,In_582,In_84);
or U1657 (N_1657,In_368,In_627);
xor U1658 (N_1658,In_670,In_535);
nand U1659 (N_1659,In_288,In_594);
nor U1660 (N_1660,In_365,In_360);
xor U1661 (N_1661,In_300,In_198);
or U1662 (N_1662,In_559,In_573);
and U1663 (N_1663,In_110,In_310);
xnor U1664 (N_1664,In_267,In_444);
nand U1665 (N_1665,In_234,In_480);
nor U1666 (N_1666,In_433,In_249);
and U1667 (N_1667,In_360,In_612);
nor U1668 (N_1668,In_286,In_346);
xnor U1669 (N_1669,In_172,In_676);
nor U1670 (N_1670,In_93,In_674);
nor U1671 (N_1671,In_123,In_36);
or U1672 (N_1672,In_54,In_676);
and U1673 (N_1673,In_222,In_43);
nor U1674 (N_1674,In_233,In_135);
nand U1675 (N_1675,In_748,In_248);
nand U1676 (N_1676,In_368,In_311);
nand U1677 (N_1677,In_315,In_208);
or U1678 (N_1678,In_244,In_32);
and U1679 (N_1679,In_15,In_600);
nor U1680 (N_1680,In_537,In_629);
nand U1681 (N_1681,In_88,In_496);
nor U1682 (N_1682,In_443,In_605);
nand U1683 (N_1683,In_304,In_521);
nor U1684 (N_1684,In_720,In_439);
nand U1685 (N_1685,In_46,In_253);
and U1686 (N_1686,In_496,In_393);
nor U1687 (N_1687,In_339,In_165);
and U1688 (N_1688,In_497,In_95);
xnor U1689 (N_1689,In_279,In_715);
nand U1690 (N_1690,In_463,In_606);
or U1691 (N_1691,In_424,In_492);
nand U1692 (N_1692,In_586,In_217);
xnor U1693 (N_1693,In_680,In_241);
nor U1694 (N_1694,In_425,In_34);
or U1695 (N_1695,In_110,In_293);
xnor U1696 (N_1696,In_225,In_535);
nand U1697 (N_1697,In_532,In_672);
or U1698 (N_1698,In_342,In_584);
or U1699 (N_1699,In_339,In_450);
nand U1700 (N_1700,In_124,In_305);
xor U1701 (N_1701,In_41,In_494);
nand U1702 (N_1702,In_686,In_271);
nor U1703 (N_1703,In_568,In_326);
xnor U1704 (N_1704,In_318,In_623);
or U1705 (N_1705,In_566,In_296);
xnor U1706 (N_1706,In_236,In_170);
xor U1707 (N_1707,In_110,In_474);
or U1708 (N_1708,In_151,In_320);
xor U1709 (N_1709,In_727,In_732);
xnor U1710 (N_1710,In_339,In_173);
or U1711 (N_1711,In_594,In_343);
xnor U1712 (N_1712,In_26,In_501);
or U1713 (N_1713,In_505,In_625);
and U1714 (N_1714,In_341,In_675);
or U1715 (N_1715,In_621,In_75);
nand U1716 (N_1716,In_24,In_481);
xnor U1717 (N_1717,In_593,In_78);
and U1718 (N_1718,In_88,In_609);
or U1719 (N_1719,In_708,In_583);
nand U1720 (N_1720,In_60,In_354);
xnor U1721 (N_1721,In_350,In_641);
or U1722 (N_1722,In_74,In_248);
and U1723 (N_1723,In_490,In_59);
nor U1724 (N_1724,In_529,In_239);
and U1725 (N_1725,In_106,In_356);
and U1726 (N_1726,In_551,In_558);
nor U1727 (N_1727,In_390,In_91);
nand U1728 (N_1728,In_478,In_26);
and U1729 (N_1729,In_718,In_216);
nand U1730 (N_1730,In_578,In_26);
xor U1731 (N_1731,In_25,In_680);
nor U1732 (N_1732,In_616,In_452);
xnor U1733 (N_1733,In_619,In_217);
and U1734 (N_1734,In_675,In_318);
nand U1735 (N_1735,In_460,In_126);
nand U1736 (N_1736,In_170,In_721);
nor U1737 (N_1737,In_46,In_204);
and U1738 (N_1738,In_238,In_272);
nand U1739 (N_1739,In_651,In_474);
nor U1740 (N_1740,In_2,In_738);
nor U1741 (N_1741,In_351,In_536);
nor U1742 (N_1742,In_737,In_557);
and U1743 (N_1743,In_533,In_514);
xor U1744 (N_1744,In_390,In_272);
nand U1745 (N_1745,In_634,In_264);
and U1746 (N_1746,In_630,In_101);
nand U1747 (N_1747,In_579,In_455);
nand U1748 (N_1748,In_661,In_20);
xor U1749 (N_1749,In_187,In_397);
nor U1750 (N_1750,In_278,In_619);
and U1751 (N_1751,In_419,In_404);
and U1752 (N_1752,In_327,In_36);
nor U1753 (N_1753,In_721,In_710);
xnor U1754 (N_1754,In_573,In_556);
and U1755 (N_1755,In_329,In_248);
or U1756 (N_1756,In_231,In_184);
or U1757 (N_1757,In_137,In_363);
nand U1758 (N_1758,In_19,In_292);
nor U1759 (N_1759,In_675,In_212);
nor U1760 (N_1760,In_486,In_667);
or U1761 (N_1761,In_111,In_527);
and U1762 (N_1762,In_421,In_249);
nand U1763 (N_1763,In_349,In_544);
nand U1764 (N_1764,In_107,In_301);
and U1765 (N_1765,In_211,In_232);
nor U1766 (N_1766,In_609,In_625);
nor U1767 (N_1767,In_149,In_721);
nor U1768 (N_1768,In_241,In_695);
nor U1769 (N_1769,In_296,In_687);
nand U1770 (N_1770,In_27,In_66);
or U1771 (N_1771,In_74,In_515);
nor U1772 (N_1772,In_440,In_268);
and U1773 (N_1773,In_64,In_487);
xnor U1774 (N_1774,In_562,In_701);
nand U1775 (N_1775,In_582,In_266);
nor U1776 (N_1776,In_592,In_454);
or U1777 (N_1777,In_743,In_97);
nand U1778 (N_1778,In_110,In_608);
and U1779 (N_1779,In_573,In_673);
nor U1780 (N_1780,In_56,In_513);
or U1781 (N_1781,In_335,In_659);
and U1782 (N_1782,In_376,In_317);
nand U1783 (N_1783,In_424,In_203);
and U1784 (N_1784,In_153,In_749);
xor U1785 (N_1785,In_273,In_724);
or U1786 (N_1786,In_335,In_296);
or U1787 (N_1787,In_147,In_662);
nand U1788 (N_1788,In_560,In_316);
or U1789 (N_1789,In_258,In_493);
or U1790 (N_1790,In_23,In_652);
xor U1791 (N_1791,In_523,In_134);
or U1792 (N_1792,In_662,In_434);
nor U1793 (N_1793,In_437,In_470);
and U1794 (N_1794,In_722,In_18);
nand U1795 (N_1795,In_278,In_33);
xnor U1796 (N_1796,In_0,In_45);
nand U1797 (N_1797,In_129,In_102);
nand U1798 (N_1798,In_99,In_505);
nor U1799 (N_1799,In_165,In_168);
xor U1800 (N_1800,In_658,In_667);
nand U1801 (N_1801,In_269,In_68);
nand U1802 (N_1802,In_690,In_237);
nand U1803 (N_1803,In_739,In_291);
or U1804 (N_1804,In_481,In_66);
or U1805 (N_1805,In_596,In_448);
or U1806 (N_1806,In_529,In_56);
or U1807 (N_1807,In_345,In_246);
nor U1808 (N_1808,In_593,In_546);
or U1809 (N_1809,In_476,In_615);
and U1810 (N_1810,In_390,In_745);
nand U1811 (N_1811,In_340,In_240);
and U1812 (N_1812,In_39,In_433);
nand U1813 (N_1813,In_317,In_399);
and U1814 (N_1814,In_360,In_343);
xnor U1815 (N_1815,In_159,In_246);
and U1816 (N_1816,In_615,In_184);
and U1817 (N_1817,In_573,In_337);
and U1818 (N_1818,In_564,In_379);
nor U1819 (N_1819,In_435,In_683);
and U1820 (N_1820,In_703,In_452);
nand U1821 (N_1821,In_494,In_271);
nor U1822 (N_1822,In_288,In_449);
nor U1823 (N_1823,In_743,In_63);
or U1824 (N_1824,In_338,In_207);
nand U1825 (N_1825,In_610,In_141);
and U1826 (N_1826,In_279,In_639);
or U1827 (N_1827,In_272,In_620);
nor U1828 (N_1828,In_692,In_703);
nand U1829 (N_1829,In_378,In_30);
or U1830 (N_1830,In_79,In_575);
nor U1831 (N_1831,In_304,In_226);
nand U1832 (N_1832,In_259,In_255);
xor U1833 (N_1833,In_701,In_485);
nand U1834 (N_1834,In_569,In_442);
xor U1835 (N_1835,In_268,In_703);
or U1836 (N_1836,In_289,In_641);
nor U1837 (N_1837,In_657,In_515);
and U1838 (N_1838,In_87,In_127);
or U1839 (N_1839,In_607,In_498);
or U1840 (N_1840,In_605,In_204);
and U1841 (N_1841,In_403,In_256);
and U1842 (N_1842,In_707,In_647);
or U1843 (N_1843,In_133,In_650);
nor U1844 (N_1844,In_668,In_721);
and U1845 (N_1845,In_416,In_125);
nand U1846 (N_1846,In_479,In_545);
xnor U1847 (N_1847,In_491,In_664);
nand U1848 (N_1848,In_501,In_608);
nor U1849 (N_1849,In_611,In_745);
nand U1850 (N_1850,In_11,In_153);
xnor U1851 (N_1851,In_347,In_459);
and U1852 (N_1852,In_288,In_334);
xor U1853 (N_1853,In_213,In_660);
or U1854 (N_1854,In_243,In_247);
nor U1855 (N_1855,In_281,In_142);
nor U1856 (N_1856,In_307,In_452);
and U1857 (N_1857,In_260,In_365);
xor U1858 (N_1858,In_604,In_704);
or U1859 (N_1859,In_510,In_747);
nor U1860 (N_1860,In_640,In_613);
nand U1861 (N_1861,In_587,In_477);
xnor U1862 (N_1862,In_691,In_439);
nand U1863 (N_1863,In_106,In_638);
nor U1864 (N_1864,In_603,In_621);
nand U1865 (N_1865,In_373,In_402);
xor U1866 (N_1866,In_25,In_476);
and U1867 (N_1867,In_393,In_251);
xnor U1868 (N_1868,In_510,In_451);
nand U1869 (N_1869,In_707,In_500);
or U1870 (N_1870,In_358,In_74);
nor U1871 (N_1871,In_515,In_181);
nand U1872 (N_1872,In_674,In_488);
nand U1873 (N_1873,In_360,In_392);
nand U1874 (N_1874,In_135,In_132);
or U1875 (N_1875,In_218,In_185);
nand U1876 (N_1876,In_57,In_663);
or U1877 (N_1877,In_78,In_721);
nand U1878 (N_1878,In_203,In_42);
or U1879 (N_1879,In_658,In_700);
xor U1880 (N_1880,In_89,In_223);
or U1881 (N_1881,In_481,In_503);
and U1882 (N_1882,In_647,In_499);
nor U1883 (N_1883,In_654,In_293);
nor U1884 (N_1884,In_55,In_242);
nand U1885 (N_1885,In_175,In_293);
and U1886 (N_1886,In_52,In_668);
xnor U1887 (N_1887,In_238,In_56);
and U1888 (N_1888,In_178,In_310);
nor U1889 (N_1889,In_580,In_305);
nand U1890 (N_1890,In_230,In_557);
or U1891 (N_1891,In_22,In_507);
or U1892 (N_1892,In_331,In_95);
nor U1893 (N_1893,In_554,In_327);
or U1894 (N_1894,In_676,In_33);
and U1895 (N_1895,In_303,In_437);
nand U1896 (N_1896,In_409,In_40);
nand U1897 (N_1897,In_674,In_515);
xnor U1898 (N_1898,In_82,In_603);
nand U1899 (N_1899,In_559,In_526);
and U1900 (N_1900,In_8,In_49);
xnor U1901 (N_1901,In_1,In_343);
or U1902 (N_1902,In_231,In_679);
nand U1903 (N_1903,In_522,In_679);
nand U1904 (N_1904,In_226,In_265);
xor U1905 (N_1905,In_60,In_383);
nor U1906 (N_1906,In_739,In_703);
xnor U1907 (N_1907,In_671,In_563);
and U1908 (N_1908,In_682,In_741);
nand U1909 (N_1909,In_447,In_630);
xor U1910 (N_1910,In_124,In_47);
nand U1911 (N_1911,In_463,In_559);
or U1912 (N_1912,In_182,In_551);
nor U1913 (N_1913,In_338,In_296);
and U1914 (N_1914,In_1,In_213);
nor U1915 (N_1915,In_394,In_638);
or U1916 (N_1916,In_511,In_748);
or U1917 (N_1917,In_696,In_135);
or U1918 (N_1918,In_203,In_545);
xnor U1919 (N_1919,In_392,In_331);
xnor U1920 (N_1920,In_178,In_391);
xnor U1921 (N_1921,In_464,In_256);
nor U1922 (N_1922,In_663,In_512);
xor U1923 (N_1923,In_577,In_597);
xor U1924 (N_1924,In_398,In_28);
nor U1925 (N_1925,In_265,In_63);
or U1926 (N_1926,In_66,In_245);
nor U1927 (N_1927,In_135,In_314);
and U1928 (N_1928,In_30,In_418);
xnor U1929 (N_1929,In_23,In_395);
nand U1930 (N_1930,In_593,In_447);
nor U1931 (N_1931,In_616,In_678);
nand U1932 (N_1932,In_32,In_41);
and U1933 (N_1933,In_516,In_627);
xnor U1934 (N_1934,In_58,In_652);
nand U1935 (N_1935,In_519,In_143);
and U1936 (N_1936,In_279,In_704);
nand U1937 (N_1937,In_747,In_321);
nor U1938 (N_1938,In_640,In_359);
xor U1939 (N_1939,In_746,In_111);
xnor U1940 (N_1940,In_705,In_516);
xor U1941 (N_1941,In_404,In_572);
and U1942 (N_1942,In_451,In_225);
nor U1943 (N_1943,In_202,In_396);
or U1944 (N_1944,In_307,In_345);
nand U1945 (N_1945,In_546,In_738);
nand U1946 (N_1946,In_53,In_68);
or U1947 (N_1947,In_468,In_609);
or U1948 (N_1948,In_503,In_255);
nand U1949 (N_1949,In_361,In_584);
nor U1950 (N_1950,In_158,In_248);
and U1951 (N_1951,In_540,In_714);
and U1952 (N_1952,In_610,In_253);
nand U1953 (N_1953,In_684,In_543);
nor U1954 (N_1954,In_266,In_630);
and U1955 (N_1955,In_47,In_32);
or U1956 (N_1956,In_607,In_726);
and U1957 (N_1957,In_363,In_311);
xor U1958 (N_1958,In_256,In_273);
xnor U1959 (N_1959,In_262,In_747);
nand U1960 (N_1960,In_37,In_146);
nor U1961 (N_1961,In_497,In_629);
or U1962 (N_1962,In_21,In_499);
nor U1963 (N_1963,In_189,In_580);
or U1964 (N_1964,In_183,In_171);
nor U1965 (N_1965,In_397,In_110);
nor U1966 (N_1966,In_320,In_596);
and U1967 (N_1967,In_588,In_206);
and U1968 (N_1968,In_22,In_83);
nand U1969 (N_1969,In_456,In_665);
nor U1970 (N_1970,In_375,In_319);
nor U1971 (N_1971,In_730,In_146);
nand U1972 (N_1972,In_152,In_270);
or U1973 (N_1973,In_104,In_502);
xor U1974 (N_1974,In_30,In_621);
nor U1975 (N_1975,In_539,In_377);
nor U1976 (N_1976,In_534,In_633);
xnor U1977 (N_1977,In_5,In_488);
and U1978 (N_1978,In_259,In_583);
and U1979 (N_1979,In_193,In_422);
nand U1980 (N_1980,In_125,In_470);
or U1981 (N_1981,In_482,In_549);
xnor U1982 (N_1982,In_318,In_701);
or U1983 (N_1983,In_239,In_200);
and U1984 (N_1984,In_306,In_75);
xor U1985 (N_1985,In_626,In_574);
or U1986 (N_1986,In_372,In_5);
nand U1987 (N_1987,In_621,In_217);
nand U1988 (N_1988,In_216,In_356);
xor U1989 (N_1989,In_429,In_24);
nand U1990 (N_1990,In_471,In_83);
xor U1991 (N_1991,In_465,In_356);
xnor U1992 (N_1992,In_459,In_575);
or U1993 (N_1993,In_71,In_264);
xor U1994 (N_1994,In_311,In_372);
xnor U1995 (N_1995,In_147,In_672);
nor U1996 (N_1996,In_396,In_55);
or U1997 (N_1997,In_453,In_354);
nor U1998 (N_1998,In_70,In_545);
or U1999 (N_1999,In_54,In_187);
nand U2000 (N_2000,In_505,In_259);
or U2001 (N_2001,In_216,In_468);
and U2002 (N_2002,In_354,In_242);
nand U2003 (N_2003,In_517,In_323);
nand U2004 (N_2004,In_295,In_92);
nor U2005 (N_2005,In_481,In_507);
nand U2006 (N_2006,In_213,In_738);
and U2007 (N_2007,In_39,In_440);
nand U2008 (N_2008,In_431,In_480);
or U2009 (N_2009,In_184,In_691);
and U2010 (N_2010,In_575,In_462);
nand U2011 (N_2011,In_636,In_439);
nand U2012 (N_2012,In_103,In_220);
nand U2013 (N_2013,In_723,In_627);
or U2014 (N_2014,In_332,In_472);
or U2015 (N_2015,In_83,In_462);
and U2016 (N_2016,In_495,In_715);
nor U2017 (N_2017,In_241,In_398);
nand U2018 (N_2018,In_630,In_565);
xor U2019 (N_2019,In_681,In_631);
nand U2020 (N_2020,In_208,In_476);
or U2021 (N_2021,In_545,In_264);
and U2022 (N_2022,In_256,In_235);
xnor U2023 (N_2023,In_64,In_734);
and U2024 (N_2024,In_450,In_26);
xnor U2025 (N_2025,In_42,In_398);
or U2026 (N_2026,In_504,In_520);
nand U2027 (N_2027,In_709,In_333);
nor U2028 (N_2028,In_724,In_61);
and U2029 (N_2029,In_379,In_15);
nand U2030 (N_2030,In_217,In_92);
and U2031 (N_2031,In_300,In_72);
nor U2032 (N_2032,In_586,In_400);
or U2033 (N_2033,In_736,In_136);
xor U2034 (N_2034,In_50,In_744);
xnor U2035 (N_2035,In_226,In_241);
nand U2036 (N_2036,In_61,In_62);
nand U2037 (N_2037,In_379,In_36);
nand U2038 (N_2038,In_559,In_69);
or U2039 (N_2039,In_463,In_651);
nor U2040 (N_2040,In_434,In_687);
nor U2041 (N_2041,In_8,In_535);
and U2042 (N_2042,In_393,In_33);
or U2043 (N_2043,In_504,In_358);
and U2044 (N_2044,In_619,In_132);
and U2045 (N_2045,In_593,In_70);
nand U2046 (N_2046,In_24,In_123);
nand U2047 (N_2047,In_118,In_475);
xnor U2048 (N_2048,In_492,In_731);
xor U2049 (N_2049,In_175,In_473);
or U2050 (N_2050,In_628,In_500);
xor U2051 (N_2051,In_246,In_674);
and U2052 (N_2052,In_288,In_75);
nor U2053 (N_2053,In_740,In_141);
nor U2054 (N_2054,In_129,In_500);
and U2055 (N_2055,In_203,In_485);
and U2056 (N_2056,In_390,In_239);
nand U2057 (N_2057,In_583,In_81);
nand U2058 (N_2058,In_171,In_153);
or U2059 (N_2059,In_612,In_664);
and U2060 (N_2060,In_294,In_521);
nor U2061 (N_2061,In_137,In_331);
nand U2062 (N_2062,In_622,In_588);
nor U2063 (N_2063,In_169,In_105);
nand U2064 (N_2064,In_186,In_415);
nor U2065 (N_2065,In_199,In_616);
nand U2066 (N_2066,In_422,In_398);
nand U2067 (N_2067,In_682,In_691);
or U2068 (N_2068,In_350,In_212);
nor U2069 (N_2069,In_672,In_400);
nand U2070 (N_2070,In_521,In_105);
or U2071 (N_2071,In_241,In_146);
or U2072 (N_2072,In_155,In_354);
or U2073 (N_2073,In_528,In_287);
and U2074 (N_2074,In_643,In_89);
nand U2075 (N_2075,In_697,In_499);
or U2076 (N_2076,In_479,In_554);
or U2077 (N_2077,In_428,In_34);
xnor U2078 (N_2078,In_372,In_580);
xor U2079 (N_2079,In_268,In_663);
or U2080 (N_2080,In_483,In_76);
nand U2081 (N_2081,In_605,In_476);
or U2082 (N_2082,In_423,In_610);
xnor U2083 (N_2083,In_584,In_87);
nor U2084 (N_2084,In_546,In_690);
and U2085 (N_2085,In_469,In_740);
nor U2086 (N_2086,In_83,In_660);
or U2087 (N_2087,In_99,In_50);
or U2088 (N_2088,In_691,In_400);
xnor U2089 (N_2089,In_277,In_552);
xnor U2090 (N_2090,In_674,In_468);
or U2091 (N_2091,In_102,In_669);
xnor U2092 (N_2092,In_136,In_432);
xnor U2093 (N_2093,In_324,In_96);
and U2094 (N_2094,In_173,In_502);
xnor U2095 (N_2095,In_501,In_153);
nor U2096 (N_2096,In_258,In_390);
or U2097 (N_2097,In_432,In_733);
or U2098 (N_2098,In_33,In_599);
or U2099 (N_2099,In_726,In_623);
and U2100 (N_2100,In_243,In_41);
or U2101 (N_2101,In_520,In_225);
and U2102 (N_2102,In_406,In_56);
nand U2103 (N_2103,In_604,In_646);
and U2104 (N_2104,In_35,In_28);
nor U2105 (N_2105,In_131,In_480);
or U2106 (N_2106,In_328,In_215);
or U2107 (N_2107,In_462,In_517);
and U2108 (N_2108,In_475,In_18);
or U2109 (N_2109,In_42,In_74);
xor U2110 (N_2110,In_668,In_431);
nor U2111 (N_2111,In_95,In_702);
nand U2112 (N_2112,In_53,In_189);
and U2113 (N_2113,In_707,In_6);
and U2114 (N_2114,In_479,In_208);
xnor U2115 (N_2115,In_555,In_334);
nor U2116 (N_2116,In_485,In_309);
and U2117 (N_2117,In_313,In_534);
nand U2118 (N_2118,In_372,In_381);
nor U2119 (N_2119,In_432,In_615);
or U2120 (N_2120,In_374,In_51);
or U2121 (N_2121,In_641,In_198);
xnor U2122 (N_2122,In_197,In_363);
xnor U2123 (N_2123,In_384,In_631);
nor U2124 (N_2124,In_167,In_734);
nor U2125 (N_2125,In_547,In_666);
and U2126 (N_2126,In_111,In_472);
nor U2127 (N_2127,In_59,In_22);
nand U2128 (N_2128,In_468,In_689);
and U2129 (N_2129,In_355,In_612);
nor U2130 (N_2130,In_678,In_670);
and U2131 (N_2131,In_8,In_47);
xnor U2132 (N_2132,In_283,In_204);
xnor U2133 (N_2133,In_745,In_594);
and U2134 (N_2134,In_376,In_511);
or U2135 (N_2135,In_149,In_616);
or U2136 (N_2136,In_698,In_592);
nand U2137 (N_2137,In_370,In_661);
or U2138 (N_2138,In_559,In_591);
nand U2139 (N_2139,In_311,In_726);
nand U2140 (N_2140,In_139,In_742);
nor U2141 (N_2141,In_342,In_608);
nand U2142 (N_2142,In_294,In_458);
or U2143 (N_2143,In_496,In_328);
and U2144 (N_2144,In_688,In_308);
nand U2145 (N_2145,In_635,In_578);
nor U2146 (N_2146,In_546,In_545);
or U2147 (N_2147,In_235,In_232);
nand U2148 (N_2148,In_293,In_412);
nand U2149 (N_2149,In_544,In_512);
or U2150 (N_2150,In_203,In_725);
nor U2151 (N_2151,In_574,In_129);
xor U2152 (N_2152,In_727,In_326);
nand U2153 (N_2153,In_454,In_76);
or U2154 (N_2154,In_201,In_425);
or U2155 (N_2155,In_748,In_684);
and U2156 (N_2156,In_414,In_360);
or U2157 (N_2157,In_184,In_287);
or U2158 (N_2158,In_742,In_694);
nand U2159 (N_2159,In_275,In_346);
and U2160 (N_2160,In_236,In_387);
xor U2161 (N_2161,In_383,In_464);
xor U2162 (N_2162,In_216,In_637);
nor U2163 (N_2163,In_343,In_658);
xnor U2164 (N_2164,In_152,In_618);
or U2165 (N_2165,In_494,In_627);
and U2166 (N_2166,In_665,In_562);
nor U2167 (N_2167,In_726,In_354);
nor U2168 (N_2168,In_518,In_195);
and U2169 (N_2169,In_702,In_433);
nor U2170 (N_2170,In_432,In_602);
nor U2171 (N_2171,In_684,In_624);
nor U2172 (N_2172,In_510,In_191);
or U2173 (N_2173,In_571,In_649);
xnor U2174 (N_2174,In_2,In_255);
nor U2175 (N_2175,In_47,In_539);
nor U2176 (N_2176,In_161,In_313);
or U2177 (N_2177,In_329,In_437);
xor U2178 (N_2178,In_381,In_503);
or U2179 (N_2179,In_43,In_68);
or U2180 (N_2180,In_150,In_114);
xor U2181 (N_2181,In_360,In_716);
nand U2182 (N_2182,In_446,In_671);
nand U2183 (N_2183,In_614,In_52);
or U2184 (N_2184,In_568,In_288);
nor U2185 (N_2185,In_478,In_555);
nand U2186 (N_2186,In_235,In_533);
nor U2187 (N_2187,In_425,In_217);
and U2188 (N_2188,In_395,In_743);
or U2189 (N_2189,In_262,In_670);
xor U2190 (N_2190,In_333,In_687);
nor U2191 (N_2191,In_192,In_412);
xor U2192 (N_2192,In_147,In_723);
xor U2193 (N_2193,In_384,In_734);
xor U2194 (N_2194,In_169,In_604);
or U2195 (N_2195,In_53,In_671);
or U2196 (N_2196,In_329,In_382);
nand U2197 (N_2197,In_57,In_735);
xnor U2198 (N_2198,In_550,In_109);
and U2199 (N_2199,In_112,In_453);
nor U2200 (N_2200,In_417,In_122);
and U2201 (N_2201,In_213,In_609);
nand U2202 (N_2202,In_714,In_444);
nor U2203 (N_2203,In_22,In_51);
nor U2204 (N_2204,In_683,In_573);
nand U2205 (N_2205,In_724,In_210);
xnor U2206 (N_2206,In_79,In_92);
xnor U2207 (N_2207,In_124,In_349);
or U2208 (N_2208,In_402,In_711);
nand U2209 (N_2209,In_710,In_90);
nand U2210 (N_2210,In_194,In_621);
nand U2211 (N_2211,In_563,In_412);
nor U2212 (N_2212,In_746,In_17);
or U2213 (N_2213,In_426,In_684);
and U2214 (N_2214,In_582,In_417);
nor U2215 (N_2215,In_592,In_325);
or U2216 (N_2216,In_22,In_139);
nand U2217 (N_2217,In_34,In_367);
xor U2218 (N_2218,In_287,In_390);
and U2219 (N_2219,In_641,In_638);
or U2220 (N_2220,In_367,In_78);
or U2221 (N_2221,In_722,In_575);
nand U2222 (N_2222,In_398,In_303);
and U2223 (N_2223,In_390,In_531);
or U2224 (N_2224,In_488,In_412);
xnor U2225 (N_2225,In_610,In_624);
xnor U2226 (N_2226,In_303,In_115);
nor U2227 (N_2227,In_715,In_143);
xor U2228 (N_2228,In_253,In_115);
and U2229 (N_2229,In_594,In_640);
or U2230 (N_2230,In_688,In_191);
xnor U2231 (N_2231,In_361,In_83);
and U2232 (N_2232,In_149,In_499);
or U2233 (N_2233,In_468,In_422);
or U2234 (N_2234,In_337,In_384);
and U2235 (N_2235,In_108,In_44);
xor U2236 (N_2236,In_494,In_258);
and U2237 (N_2237,In_0,In_150);
xnor U2238 (N_2238,In_255,In_398);
and U2239 (N_2239,In_304,In_144);
xnor U2240 (N_2240,In_540,In_9);
nand U2241 (N_2241,In_367,In_275);
nand U2242 (N_2242,In_726,In_609);
xnor U2243 (N_2243,In_286,In_84);
nand U2244 (N_2244,In_601,In_628);
nand U2245 (N_2245,In_550,In_399);
nor U2246 (N_2246,In_655,In_646);
or U2247 (N_2247,In_307,In_217);
nor U2248 (N_2248,In_553,In_542);
nand U2249 (N_2249,In_275,In_723);
and U2250 (N_2250,In_349,In_545);
nor U2251 (N_2251,In_26,In_326);
nand U2252 (N_2252,In_100,In_550);
nand U2253 (N_2253,In_66,In_464);
or U2254 (N_2254,In_512,In_344);
or U2255 (N_2255,In_656,In_221);
and U2256 (N_2256,In_499,In_32);
and U2257 (N_2257,In_258,In_255);
nand U2258 (N_2258,In_152,In_397);
and U2259 (N_2259,In_342,In_404);
nand U2260 (N_2260,In_713,In_521);
nand U2261 (N_2261,In_1,In_709);
or U2262 (N_2262,In_342,In_166);
and U2263 (N_2263,In_689,In_473);
or U2264 (N_2264,In_736,In_450);
xor U2265 (N_2265,In_597,In_143);
nor U2266 (N_2266,In_639,In_216);
nor U2267 (N_2267,In_584,In_37);
or U2268 (N_2268,In_360,In_73);
nor U2269 (N_2269,In_305,In_706);
or U2270 (N_2270,In_331,In_696);
nand U2271 (N_2271,In_260,In_107);
or U2272 (N_2272,In_170,In_657);
or U2273 (N_2273,In_68,In_567);
xnor U2274 (N_2274,In_645,In_694);
and U2275 (N_2275,In_655,In_632);
or U2276 (N_2276,In_153,In_249);
or U2277 (N_2277,In_667,In_404);
nor U2278 (N_2278,In_423,In_387);
nor U2279 (N_2279,In_544,In_432);
xnor U2280 (N_2280,In_523,In_291);
nand U2281 (N_2281,In_200,In_717);
nand U2282 (N_2282,In_746,In_735);
xnor U2283 (N_2283,In_266,In_290);
or U2284 (N_2284,In_451,In_543);
or U2285 (N_2285,In_686,In_274);
nand U2286 (N_2286,In_249,In_222);
and U2287 (N_2287,In_159,In_299);
or U2288 (N_2288,In_713,In_539);
xnor U2289 (N_2289,In_617,In_302);
nor U2290 (N_2290,In_19,In_395);
or U2291 (N_2291,In_56,In_224);
and U2292 (N_2292,In_53,In_377);
or U2293 (N_2293,In_408,In_740);
nor U2294 (N_2294,In_611,In_615);
or U2295 (N_2295,In_399,In_614);
nor U2296 (N_2296,In_463,In_396);
or U2297 (N_2297,In_67,In_63);
or U2298 (N_2298,In_330,In_2);
or U2299 (N_2299,In_461,In_497);
or U2300 (N_2300,In_555,In_38);
nor U2301 (N_2301,In_326,In_424);
and U2302 (N_2302,In_150,In_269);
xnor U2303 (N_2303,In_523,In_55);
nand U2304 (N_2304,In_47,In_614);
and U2305 (N_2305,In_280,In_487);
nor U2306 (N_2306,In_744,In_75);
nor U2307 (N_2307,In_311,In_305);
nand U2308 (N_2308,In_314,In_59);
nand U2309 (N_2309,In_255,In_207);
xnor U2310 (N_2310,In_347,In_636);
nand U2311 (N_2311,In_156,In_201);
and U2312 (N_2312,In_426,In_520);
or U2313 (N_2313,In_212,In_657);
nand U2314 (N_2314,In_123,In_597);
nand U2315 (N_2315,In_741,In_338);
nor U2316 (N_2316,In_212,In_554);
xor U2317 (N_2317,In_50,In_171);
and U2318 (N_2318,In_131,In_60);
or U2319 (N_2319,In_198,In_534);
and U2320 (N_2320,In_543,In_220);
and U2321 (N_2321,In_504,In_688);
xor U2322 (N_2322,In_676,In_737);
nand U2323 (N_2323,In_377,In_715);
nand U2324 (N_2324,In_677,In_44);
and U2325 (N_2325,In_210,In_163);
and U2326 (N_2326,In_166,In_584);
nand U2327 (N_2327,In_513,In_209);
or U2328 (N_2328,In_309,In_50);
and U2329 (N_2329,In_121,In_624);
or U2330 (N_2330,In_497,In_598);
xor U2331 (N_2331,In_93,In_445);
and U2332 (N_2332,In_14,In_602);
and U2333 (N_2333,In_532,In_464);
or U2334 (N_2334,In_22,In_274);
and U2335 (N_2335,In_488,In_470);
and U2336 (N_2336,In_742,In_324);
and U2337 (N_2337,In_586,In_168);
and U2338 (N_2338,In_376,In_412);
nand U2339 (N_2339,In_232,In_185);
and U2340 (N_2340,In_333,In_471);
xor U2341 (N_2341,In_742,In_415);
or U2342 (N_2342,In_258,In_744);
xnor U2343 (N_2343,In_626,In_33);
nand U2344 (N_2344,In_426,In_451);
and U2345 (N_2345,In_454,In_622);
xnor U2346 (N_2346,In_476,In_467);
nand U2347 (N_2347,In_437,In_169);
or U2348 (N_2348,In_209,In_152);
xnor U2349 (N_2349,In_75,In_381);
and U2350 (N_2350,In_710,In_160);
and U2351 (N_2351,In_201,In_581);
nor U2352 (N_2352,In_443,In_679);
xnor U2353 (N_2353,In_177,In_114);
nor U2354 (N_2354,In_379,In_274);
or U2355 (N_2355,In_84,In_187);
or U2356 (N_2356,In_585,In_618);
and U2357 (N_2357,In_264,In_691);
xnor U2358 (N_2358,In_452,In_651);
and U2359 (N_2359,In_120,In_611);
nand U2360 (N_2360,In_672,In_418);
xnor U2361 (N_2361,In_58,In_106);
nor U2362 (N_2362,In_76,In_214);
nand U2363 (N_2363,In_75,In_175);
and U2364 (N_2364,In_592,In_63);
and U2365 (N_2365,In_90,In_470);
and U2366 (N_2366,In_122,In_276);
and U2367 (N_2367,In_724,In_675);
or U2368 (N_2368,In_411,In_2);
and U2369 (N_2369,In_400,In_631);
or U2370 (N_2370,In_91,In_456);
nand U2371 (N_2371,In_696,In_197);
nand U2372 (N_2372,In_366,In_369);
nand U2373 (N_2373,In_631,In_302);
and U2374 (N_2374,In_733,In_157);
and U2375 (N_2375,In_543,In_329);
and U2376 (N_2376,In_720,In_403);
or U2377 (N_2377,In_239,In_393);
xor U2378 (N_2378,In_389,In_104);
nor U2379 (N_2379,In_14,In_222);
nor U2380 (N_2380,In_90,In_212);
nand U2381 (N_2381,In_684,In_281);
xnor U2382 (N_2382,In_664,In_214);
nor U2383 (N_2383,In_130,In_584);
xor U2384 (N_2384,In_164,In_451);
nor U2385 (N_2385,In_664,In_107);
xnor U2386 (N_2386,In_88,In_156);
xor U2387 (N_2387,In_336,In_564);
xnor U2388 (N_2388,In_400,In_274);
or U2389 (N_2389,In_639,In_222);
or U2390 (N_2390,In_150,In_617);
xnor U2391 (N_2391,In_470,In_94);
nor U2392 (N_2392,In_334,In_141);
nand U2393 (N_2393,In_749,In_290);
and U2394 (N_2394,In_365,In_33);
nand U2395 (N_2395,In_702,In_640);
or U2396 (N_2396,In_623,In_196);
xnor U2397 (N_2397,In_303,In_55);
nor U2398 (N_2398,In_581,In_578);
xor U2399 (N_2399,In_486,In_720);
or U2400 (N_2400,In_210,In_100);
nor U2401 (N_2401,In_47,In_477);
nand U2402 (N_2402,In_122,In_298);
and U2403 (N_2403,In_438,In_542);
xnor U2404 (N_2404,In_568,In_44);
or U2405 (N_2405,In_323,In_48);
nand U2406 (N_2406,In_585,In_157);
nand U2407 (N_2407,In_507,In_266);
and U2408 (N_2408,In_323,In_244);
or U2409 (N_2409,In_457,In_175);
nor U2410 (N_2410,In_729,In_489);
or U2411 (N_2411,In_141,In_584);
or U2412 (N_2412,In_651,In_236);
nor U2413 (N_2413,In_638,In_395);
nand U2414 (N_2414,In_678,In_644);
and U2415 (N_2415,In_394,In_480);
nor U2416 (N_2416,In_259,In_205);
xor U2417 (N_2417,In_33,In_155);
and U2418 (N_2418,In_625,In_158);
and U2419 (N_2419,In_529,In_42);
nor U2420 (N_2420,In_513,In_280);
nor U2421 (N_2421,In_128,In_394);
nand U2422 (N_2422,In_147,In_429);
xnor U2423 (N_2423,In_87,In_246);
xnor U2424 (N_2424,In_451,In_186);
nor U2425 (N_2425,In_570,In_548);
nand U2426 (N_2426,In_49,In_437);
nand U2427 (N_2427,In_674,In_13);
nor U2428 (N_2428,In_684,In_587);
and U2429 (N_2429,In_66,In_652);
xor U2430 (N_2430,In_145,In_137);
or U2431 (N_2431,In_86,In_711);
xnor U2432 (N_2432,In_700,In_323);
nor U2433 (N_2433,In_546,In_153);
nor U2434 (N_2434,In_401,In_407);
and U2435 (N_2435,In_397,In_615);
nand U2436 (N_2436,In_58,In_351);
or U2437 (N_2437,In_187,In_336);
and U2438 (N_2438,In_362,In_353);
nor U2439 (N_2439,In_658,In_719);
and U2440 (N_2440,In_714,In_391);
nor U2441 (N_2441,In_204,In_716);
xor U2442 (N_2442,In_597,In_526);
and U2443 (N_2443,In_725,In_555);
or U2444 (N_2444,In_400,In_180);
xnor U2445 (N_2445,In_645,In_507);
and U2446 (N_2446,In_673,In_480);
xnor U2447 (N_2447,In_554,In_428);
nand U2448 (N_2448,In_334,In_181);
xor U2449 (N_2449,In_298,In_597);
and U2450 (N_2450,In_645,In_513);
and U2451 (N_2451,In_338,In_221);
nand U2452 (N_2452,In_337,In_463);
or U2453 (N_2453,In_147,In_44);
or U2454 (N_2454,In_334,In_258);
and U2455 (N_2455,In_604,In_456);
and U2456 (N_2456,In_266,In_584);
nand U2457 (N_2457,In_304,In_1);
and U2458 (N_2458,In_536,In_741);
xnor U2459 (N_2459,In_413,In_711);
and U2460 (N_2460,In_667,In_142);
xnor U2461 (N_2461,In_452,In_260);
and U2462 (N_2462,In_49,In_674);
or U2463 (N_2463,In_176,In_309);
or U2464 (N_2464,In_587,In_13);
nand U2465 (N_2465,In_236,In_503);
xor U2466 (N_2466,In_212,In_119);
and U2467 (N_2467,In_661,In_722);
xnor U2468 (N_2468,In_465,In_427);
or U2469 (N_2469,In_85,In_552);
nor U2470 (N_2470,In_421,In_218);
nand U2471 (N_2471,In_381,In_137);
nor U2472 (N_2472,In_428,In_350);
nand U2473 (N_2473,In_270,In_446);
or U2474 (N_2474,In_525,In_459);
or U2475 (N_2475,In_253,In_214);
nand U2476 (N_2476,In_374,In_570);
xnor U2477 (N_2477,In_682,In_678);
xor U2478 (N_2478,In_653,In_403);
xnor U2479 (N_2479,In_313,In_662);
nor U2480 (N_2480,In_158,In_62);
nor U2481 (N_2481,In_207,In_604);
or U2482 (N_2482,In_619,In_182);
nor U2483 (N_2483,In_42,In_223);
nand U2484 (N_2484,In_596,In_744);
nand U2485 (N_2485,In_464,In_182);
nand U2486 (N_2486,In_78,In_456);
xnor U2487 (N_2487,In_553,In_608);
or U2488 (N_2488,In_718,In_387);
xnor U2489 (N_2489,In_124,In_432);
and U2490 (N_2490,In_102,In_470);
or U2491 (N_2491,In_726,In_596);
nand U2492 (N_2492,In_389,In_361);
nor U2493 (N_2493,In_680,In_469);
nand U2494 (N_2494,In_611,In_38);
xor U2495 (N_2495,In_208,In_571);
nor U2496 (N_2496,In_75,In_157);
and U2497 (N_2497,In_693,In_340);
or U2498 (N_2498,In_399,In_655);
and U2499 (N_2499,In_205,In_706);
or U2500 (N_2500,N_25,N_1012);
and U2501 (N_2501,N_531,N_198);
nand U2502 (N_2502,N_305,N_433);
xor U2503 (N_2503,N_1376,N_1570);
or U2504 (N_2504,N_455,N_345);
and U2505 (N_2505,N_553,N_529);
or U2506 (N_2506,N_2473,N_955);
nor U2507 (N_2507,N_845,N_1545);
or U2508 (N_2508,N_986,N_1756);
and U2509 (N_2509,N_1574,N_2358);
xor U2510 (N_2510,N_662,N_1506);
nand U2511 (N_2511,N_772,N_925);
and U2512 (N_2512,N_549,N_1922);
nor U2513 (N_2513,N_213,N_2097);
and U2514 (N_2514,N_1523,N_2045);
nor U2515 (N_2515,N_2411,N_1924);
or U2516 (N_2516,N_1009,N_1901);
and U2517 (N_2517,N_1881,N_231);
nor U2518 (N_2518,N_1710,N_1737);
xnor U2519 (N_2519,N_1507,N_1160);
or U2520 (N_2520,N_664,N_2039);
nor U2521 (N_2521,N_2116,N_1417);
xor U2522 (N_2522,N_1800,N_2338);
and U2523 (N_2523,N_534,N_1589);
nor U2524 (N_2524,N_494,N_1086);
or U2525 (N_2525,N_1220,N_1459);
nand U2526 (N_2526,N_655,N_851);
nor U2527 (N_2527,N_1436,N_1662);
nor U2528 (N_2528,N_295,N_255);
nand U2529 (N_2529,N_2173,N_735);
and U2530 (N_2530,N_1107,N_2110);
nand U2531 (N_2531,N_436,N_2264);
nor U2532 (N_2532,N_536,N_2459);
nor U2533 (N_2533,N_1972,N_2288);
nand U2534 (N_2534,N_942,N_2197);
and U2535 (N_2535,N_2008,N_149);
and U2536 (N_2536,N_896,N_475);
or U2537 (N_2537,N_604,N_2133);
or U2538 (N_2538,N_828,N_2200);
nor U2539 (N_2539,N_374,N_600);
nand U2540 (N_2540,N_2191,N_1460);
nand U2541 (N_2541,N_856,N_430);
or U2542 (N_2542,N_2034,N_2095);
nor U2543 (N_2543,N_1556,N_2463);
or U2544 (N_2544,N_163,N_1213);
xor U2545 (N_2545,N_912,N_882);
and U2546 (N_2546,N_1612,N_770);
xor U2547 (N_2547,N_2451,N_1394);
and U2548 (N_2548,N_339,N_2027);
nor U2549 (N_2549,N_1375,N_1030);
or U2550 (N_2550,N_510,N_593);
xor U2551 (N_2551,N_2483,N_139);
xor U2552 (N_2552,N_1920,N_2438);
nand U2553 (N_2553,N_425,N_680);
xnor U2554 (N_2554,N_607,N_519);
and U2555 (N_2555,N_1027,N_1419);
xnor U2556 (N_2556,N_91,N_1351);
or U2557 (N_2557,N_1004,N_825);
nor U2558 (N_2558,N_903,N_1156);
nor U2559 (N_2559,N_623,N_1127);
and U2560 (N_2560,N_109,N_785);
nand U2561 (N_2561,N_787,N_799);
nor U2562 (N_2562,N_818,N_2377);
xnor U2563 (N_2563,N_2328,N_2449);
or U2564 (N_2564,N_1807,N_1008);
or U2565 (N_2565,N_1536,N_2131);
or U2566 (N_2566,N_1289,N_2482);
or U2567 (N_2567,N_2370,N_1784);
nand U2568 (N_2568,N_489,N_611);
xor U2569 (N_2569,N_394,N_1532);
nor U2570 (N_2570,N_1644,N_621);
xnor U2571 (N_2571,N_186,N_2431);
and U2572 (N_2572,N_471,N_1108);
or U2573 (N_2573,N_2006,N_724);
and U2574 (N_2574,N_68,N_413);
xnor U2575 (N_2575,N_2219,N_1795);
nand U2576 (N_2576,N_2074,N_2147);
xor U2577 (N_2577,N_863,N_86);
or U2578 (N_2578,N_1251,N_316);
xor U2579 (N_2579,N_308,N_225);
xnor U2580 (N_2580,N_188,N_1699);
and U2581 (N_2581,N_2189,N_2426);
xor U2582 (N_2582,N_628,N_892);
xor U2583 (N_2583,N_1392,N_2235);
nor U2584 (N_2584,N_1828,N_1391);
nand U2585 (N_2585,N_382,N_364);
nor U2586 (N_2586,N_1063,N_1905);
or U2587 (N_2587,N_314,N_377);
and U2588 (N_2588,N_1346,N_826);
and U2589 (N_2589,N_1073,N_2321);
and U2590 (N_2590,N_2151,N_199);
nor U2591 (N_2591,N_775,N_1447);
xor U2592 (N_2592,N_741,N_2170);
or U2593 (N_2593,N_1007,N_2367);
and U2594 (N_2594,N_2193,N_997);
and U2595 (N_2595,N_954,N_2041);
xor U2596 (N_2596,N_1455,N_1087);
and U2597 (N_2597,N_792,N_2013);
nand U2598 (N_2598,N_1553,N_507);
or U2599 (N_2599,N_1898,N_1379);
or U2600 (N_2600,N_1718,N_1162);
and U2601 (N_2601,N_114,N_85);
nor U2602 (N_2602,N_2194,N_1918);
and U2603 (N_2603,N_2030,N_6);
and U2604 (N_2604,N_798,N_51);
or U2605 (N_2605,N_645,N_2399);
nand U2606 (N_2606,N_1785,N_411);
and U2607 (N_2607,N_281,N_5);
nand U2608 (N_2608,N_1735,N_597);
and U2609 (N_2609,N_2100,N_448);
nor U2610 (N_2610,N_594,N_1040);
and U2611 (N_2611,N_2232,N_635);
nand U2612 (N_2612,N_1979,N_28);
nand U2613 (N_2613,N_166,N_2401);
and U2614 (N_2614,N_216,N_1407);
and U2615 (N_2615,N_2249,N_1401);
nor U2616 (N_2616,N_690,N_2055);
xnor U2617 (N_2617,N_1762,N_2089);
nand U2618 (N_2618,N_1457,N_151);
nand U2619 (N_2619,N_1701,N_921);
and U2620 (N_2620,N_95,N_1902);
or U2621 (N_2621,N_1712,N_1695);
nor U2622 (N_2622,N_1148,N_627);
nand U2623 (N_2623,N_1554,N_379);
and U2624 (N_2624,N_524,N_910);
nand U2625 (N_2625,N_2282,N_1981);
and U2626 (N_2626,N_1907,N_323);
nor U2627 (N_2627,N_1431,N_2098);
xor U2628 (N_2628,N_2428,N_36);
nor U2629 (N_2629,N_1858,N_1912);
nor U2630 (N_2630,N_1282,N_2277);
nand U2631 (N_2631,N_218,N_839);
or U2632 (N_2632,N_1229,N_1094);
or U2633 (N_2633,N_2016,N_282);
nand U2634 (N_2634,N_602,N_69);
and U2635 (N_2635,N_1781,N_1477);
nand U2636 (N_2636,N_2169,N_2032);
nor U2637 (N_2637,N_234,N_505);
nor U2638 (N_2638,N_1999,N_2036);
xnor U2639 (N_2639,N_486,N_1950);
xnor U2640 (N_2640,N_205,N_22);
or U2641 (N_2641,N_306,N_1505);
nand U2642 (N_2642,N_965,N_1432);
nor U2643 (N_2643,N_1512,N_802);
xor U2644 (N_2644,N_1958,N_487);
and U2645 (N_2645,N_19,N_2260);
nor U2646 (N_2646,N_2261,N_2429);
and U2647 (N_2647,N_1497,N_1631);
nor U2648 (N_2648,N_1855,N_484);
or U2649 (N_2649,N_878,N_7);
and U2650 (N_2650,N_267,N_1703);
or U2651 (N_2651,N_1759,N_1362);
or U2652 (N_2652,N_778,N_195);
or U2653 (N_2653,N_117,N_1615);
nand U2654 (N_2654,N_2237,N_367);
xor U2655 (N_2655,N_1060,N_657);
nor U2656 (N_2656,N_477,N_1622);
nor U2657 (N_2657,N_2091,N_12);
and U2658 (N_2658,N_667,N_2295);
nand U2659 (N_2659,N_460,N_2205);
or U2660 (N_2660,N_1332,N_665);
xnor U2661 (N_2661,N_1441,N_1716);
nor U2662 (N_2662,N_1177,N_2405);
xor U2663 (N_2663,N_2172,N_1215);
and U2664 (N_2664,N_2332,N_516);
nand U2665 (N_2665,N_1890,N_937);
and U2666 (N_2666,N_2102,N_840);
and U2667 (N_2667,N_1371,N_2289);
nor U2668 (N_2668,N_1452,N_2479);
nand U2669 (N_2669,N_1204,N_1264);
nor U2670 (N_2670,N_1373,N_1608);
xor U2671 (N_2671,N_722,N_1696);
or U2672 (N_2672,N_1592,N_1549);
or U2673 (N_2673,N_294,N_1402);
nor U2674 (N_2674,N_1633,N_2047);
nand U2675 (N_2675,N_608,N_2268);
nor U2676 (N_2676,N_313,N_265);
xor U2677 (N_2677,N_2222,N_16);
xnor U2678 (N_2678,N_649,N_2085);
nand U2679 (N_2679,N_1011,N_1643);
xor U2680 (N_2680,N_2478,N_1363);
nor U2681 (N_2681,N_179,N_1867);
or U2682 (N_2682,N_1492,N_2413);
and U2683 (N_2683,N_1276,N_2033);
xor U2684 (N_2684,N_709,N_1036);
and U2685 (N_2685,N_836,N_1664);
nor U2686 (N_2686,N_351,N_1952);
and U2687 (N_2687,N_241,N_846);
or U2688 (N_2688,N_753,N_1397);
nand U2689 (N_2689,N_1680,N_1181);
and U2690 (N_2690,N_206,N_2273);
xor U2691 (N_2691,N_497,N_1797);
xor U2692 (N_2692,N_1439,N_1487);
nand U2693 (N_2693,N_2115,N_2175);
xor U2694 (N_2694,N_426,N_1021);
and U2695 (N_2695,N_287,N_2373);
or U2696 (N_2696,N_589,N_913);
or U2697 (N_2697,N_715,N_1640);
nor U2698 (N_2698,N_2466,N_1734);
nor U2699 (N_2699,N_780,N_1575);
nor U2700 (N_2700,N_122,N_1138);
nor U2701 (N_2701,N_482,N_1951);
nor U2702 (N_2702,N_699,N_2319);
nand U2703 (N_2703,N_318,N_196);
or U2704 (N_2704,N_1968,N_8);
nand U2705 (N_2705,N_418,N_1100);
nor U2706 (N_2706,N_634,N_742);
nor U2707 (N_2707,N_1947,N_2225);
xor U2708 (N_2708,N_1655,N_1225);
or U2709 (N_2709,N_644,N_1124);
xnor U2710 (N_2710,N_1051,N_2094);
nand U2711 (N_2711,N_1562,N_2035);
nand U2712 (N_2712,N_52,N_2375);
or U2713 (N_2713,N_528,N_733);
nor U2714 (N_2714,N_1179,N_570);
and U2715 (N_2715,N_1634,N_2212);
nor U2716 (N_2716,N_1121,N_2093);
and U2717 (N_2717,N_2203,N_1923);
nand U2718 (N_2718,N_328,N_1047);
nand U2719 (N_2719,N_976,N_424);
and U2720 (N_2720,N_1185,N_1805);
or U2721 (N_2721,N_1223,N_2347);
or U2722 (N_2722,N_848,N_551);
xor U2723 (N_2723,N_1061,N_1911);
nand U2724 (N_2724,N_1724,N_2427);
and U2725 (N_2725,N_564,N_2216);
nor U2726 (N_2726,N_1572,N_156);
xor U2727 (N_2727,N_469,N_310);
xnor U2728 (N_2728,N_1050,N_847);
and U2729 (N_2729,N_578,N_978);
or U2730 (N_2730,N_2121,N_273);
or U2731 (N_2731,N_427,N_599);
nor U2732 (N_2732,N_1930,N_1769);
xnor U2733 (N_2733,N_1058,N_1939);
nor U2734 (N_2734,N_1262,N_2185);
and U2735 (N_2735,N_50,N_2283);
nand U2736 (N_2736,N_508,N_76);
and U2737 (N_2737,N_2031,N_694);
and U2738 (N_2738,N_1269,N_1739);
nor U2739 (N_2739,N_2066,N_2470);
nand U2740 (N_2740,N_2207,N_734);
nand U2741 (N_2741,N_981,N_1421);
nor U2742 (N_2742,N_1675,N_669);
and U2743 (N_2743,N_492,N_1817);
and U2744 (N_2744,N_829,N_2388);
or U2745 (N_2745,N_1601,N_1428);
nand U2746 (N_2746,N_2424,N_1728);
xnor U2747 (N_2747,N_2383,N_745);
or U2748 (N_2748,N_1463,N_454);
nand U2749 (N_2749,N_746,N_1222);
and U2750 (N_2750,N_1365,N_217);
nor U2751 (N_2751,N_1842,N_1435);
nor U2752 (N_2752,N_1164,N_1015);
xor U2753 (N_2753,N_1228,N_2215);
and U2754 (N_2754,N_366,N_880);
nor U2755 (N_2755,N_133,N_1767);
and U2756 (N_2756,N_1184,N_2071);
and U2757 (N_2757,N_2099,N_1422);
xnor U2758 (N_2758,N_478,N_1141);
and U2759 (N_2759,N_521,N_2214);
and U2760 (N_2760,N_1883,N_811);
nor U2761 (N_2761,N_1456,N_105);
xnor U2762 (N_2762,N_1374,N_1515);
or U2763 (N_2763,N_340,N_691);
nor U2764 (N_2764,N_843,N_1420);
nand U2765 (N_2765,N_577,N_1687);
xor U2766 (N_2766,N_1773,N_901);
and U2767 (N_2767,N_2298,N_760);
and U2768 (N_2768,N_1216,N_1168);
nor U2769 (N_2769,N_399,N_1518);
xnor U2770 (N_2770,N_584,N_2234);
nor U2771 (N_2771,N_1861,N_1763);
and U2772 (N_2772,N_391,N_1731);
nand U2773 (N_2773,N_2391,N_1743);
and U2774 (N_2774,N_1409,N_2472);
or U2775 (N_2775,N_1064,N_203);
xnor U2776 (N_2776,N_1651,N_1281);
nand U2777 (N_2777,N_1565,N_1587);
nor U2778 (N_2778,N_1437,N_279);
xor U2779 (N_2779,N_782,N_1607);
or U2780 (N_2780,N_1450,N_1338);
and U2781 (N_2781,N_776,N_1768);
nand U2782 (N_2782,N_659,N_271);
and U2783 (N_2783,N_325,N_964);
xor U2784 (N_2784,N_974,N_159);
nand U2785 (N_2785,N_2302,N_495);
or U2786 (N_2786,N_1688,N_966);
or U2787 (N_2787,N_1559,N_739);
nand U2788 (N_2788,N_2192,N_2318);
nor U2789 (N_2789,N_1387,N_800);
nor U2790 (N_2790,N_1585,N_2226);
nor U2791 (N_2791,N_2351,N_1105);
nor U2792 (N_2792,N_1588,N_701);
nor U2793 (N_2793,N_1674,N_1927);
or U2794 (N_2794,N_242,N_1333);
and U2795 (N_2795,N_1789,N_1956);
or U2796 (N_2796,N_1042,N_1411);
xnor U2797 (N_2797,N_750,N_1353);
and U2798 (N_2798,N_237,N_2186);
xnor U2799 (N_2799,N_462,N_1090);
or U2800 (N_2800,N_1296,N_689);
xor U2801 (N_2801,N_2160,N_1823);
xnor U2802 (N_2802,N_2334,N_1410);
and U2803 (N_2803,N_1705,N_184);
or U2804 (N_2804,N_884,N_1329);
and U2805 (N_2805,N_1458,N_360);
nor U2806 (N_2806,N_1513,N_2010);
xor U2807 (N_2807,N_1535,N_2244);
nand U2808 (N_2808,N_985,N_372);
or U2809 (N_2809,N_2297,N_215);
nor U2810 (N_2810,N_1539,N_1840);
or U2811 (N_2811,N_889,N_1366);
xor U2812 (N_2812,N_1698,N_1316);
and U2813 (N_2813,N_1874,N_1961);
nor U2814 (N_2814,N_481,N_88);
and U2815 (N_2815,N_2112,N_353);
nand U2816 (N_2816,N_1793,N_1189);
nor U2817 (N_2817,N_2360,N_1445);
and U2818 (N_2818,N_1786,N_2162);
nor U2819 (N_2819,N_1197,N_990);
nor U2820 (N_2820,N_1826,N_2054);
and U2821 (N_2821,N_1234,N_1089);
xnor U2822 (N_2822,N_1537,N_1158);
or U2823 (N_2823,N_1226,N_784);
and U2824 (N_2824,N_1246,N_1654);
or U2825 (N_2825,N_2352,N_767);
and U2826 (N_2826,N_1285,N_66);
nand U2827 (N_2827,N_75,N_1736);
xor U2828 (N_2828,N_9,N_2171);
xnor U2829 (N_2829,N_2355,N_1151);
or U2830 (N_2830,N_407,N_1043);
nor U2831 (N_2831,N_1405,N_1624);
nand U2832 (N_2832,N_2143,N_697);
xor U2833 (N_2833,N_2471,N_130);
nor U2834 (N_2834,N_875,N_1238);
and U2835 (N_2835,N_290,N_1893);
nand U2836 (N_2836,N_1480,N_2402);
xor U2837 (N_2837,N_2307,N_2181);
and U2838 (N_2838,N_201,N_1097);
and U2839 (N_2839,N_613,N_1621);
xnor U2840 (N_2840,N_2259,N_855);
nand U2841 (N_2841,N_1746,N_758);
nor U2842 (N_2842,N_1929,N_1590);
nor U2843 (N_2843,N_1469,N_1006);
xor U2844 (N_2844,N_1290,N_1941);
and U2845 (N_2845,N_361,N_77);
or U2846 (N_2846,N_2275,N_2210);
nand U2847 (N_2847,N_1685,N_1741);
or U2848 (N_2848,N_2046,N_148);
and U2849 (N_2849,N_209,N_2231);
or U2850 (N_2850,N_1335,N_29);
xnor U2851 (N_2851,N_517,N_1261);
or U2852 (N_2852,N_124,N_1494);
or U2853 (N_2853,N_2294,N_270);
and U2854 (N_2854,N_1959,N_1862);
or U2855 (N_2855,N_939,N_1713);
and U2856 (N_2856,N_1209,N_2490);
nand U2857 (N_2857,N_1336,N_150);
nand U2858 (N_2858,N_685,N_342);
nor U2859 (N_2859,N_140,N_1501);
xnor U2860 (N_2860,N_1242,N_1853);
xnor U2861 (N_2861,N_2204,N_1758);
and U2862 (N_2862,N_632,N_1940);
or U2863 (N_2863,N_1331,N_2433);
nor U2864 (N_2864,N_2496,N_359);
or U2865 (N_2865,N_1122,N_1665);
xnor U2866 (N_2866,N_740,N_1103);
nand U2867 (N_2867,N_1399,N_1482);
and U2868 (N_2868,N_730,N_1174);
and U2869 (N_2869,N_1082,N_676);
nor U2870 (N_2870,N_1879,N_1875);
and U2871 (N_2871,N_1081,N_2380);
and U2872 (N_2872,N_708,N_500);
nor U2873 (N_2873,N_905,N_1292);
xor U2874 (N_2874,N_1418,N_2064);
xnor U2875 (N_2875,N_1300,N_931);
and U2876 (N_2876,N_1673,N_995);
and U2877 (N_2877,N_2484,N_769);
and U2878 (N_2878,N_1514,N_1057);
xnor U2879 (N_2879,N_2304,N_1991);
and U2880 (N_2880,N_2366,N_2323);
or U2881 (N_2881,N_2311,N_2293);
nand U2882 (N_2882,N_2245,N_2300);
and U2883 (N_2883,N_2368,N_941);
xor U2884 (N_2884,N_40,N_1339);
nor U2885 (N_2885,N_1866,N_2291);
or U2886 (N_2886,N_2043,N_1288);
or U2887 (N_2887,N_943,N_2442);
nand U2888 (N_2888,N_1322,N_539);
xnor U2889 (N_2889,N_2477,N_652);
or U2890 (N_2890,N_1311,N_1369);
or U2891 (N_2891,N_473,N_1344);
nor U2892 (N_2892,N_2003,N_1489);
nand U2893 (N_2893,N_1208,N_2336);
nor U2894 (N_2894,N_1367,N_1462);
nor U2895 (N_2895,N_1686,N_2096);
and U2896 (N_2896,N_2418,N_2004);
and U2897 (N_2897,N_1852,N_532);
nand U2898 (N_2898,N_1843,N_563);
and U2899 (N_2899,N_2270,N_142);
or U2900 (N_2900,N_842,N_2480);
or U2901 (N_2901,N_2209,N_2267);
or U2902 (N_2902,N_869,N_1304);
nor U2903 (N_2903,N_579,N_2410);
xnor U2904 (N_2904,N_2497,N_2365);
nor U2905 (N_2905,N_804,N_1798);
nor U2906 (N_2906,N_98,N_390);
nand U2907 (N_2907,N_2048,N_1041);
and U2908 (N_2908,N_2007,N_751);
and U2909 (N_2909,N_1440,N_1803);
or U2910 (N_2910,N_2213,N_874);
or U2911 (N_2911,N_356,N_1953);
and U2912 (N_2912,N_1844,N_89);
xnor U2913 (N_2913,N_1014,N_1312);
or U2914 (N_2914,N_1567,N_548);
or U2915 (N_2915,N_1119,N_11);
xnor U2916 (N_2916,N_2475,N_173);
xor U2917 (N_2917,N_587,N_283);
and U2918 (N_2918,N_1591,N_2345);
nand U2919 (N_2919,N_2243,N_642);
or U2920 (N_2920,N_550,N_830);
nand U2921 (N_2921,N_1217,N_2395);
nand U2922 (N_2922,N_1689,N_565);
or U2923 (N_2923,N_886,N_1577);
xnor U2924 (N_2924,N_2448,N_513);
xor U2925 (N_2925,N_1053,N_414);
or U2926 (N_2926,N_396,N_2078);
nor U2927 (N_2927,N_2156,N_115);
or U2928 (N_2928,N_392,N_284);
and U2929 (N_2929,N_2263,N_311);
nand U2930 (N_2930,N_864,N_397);
and U2931 (N_2931,N_1582,N_1906);
nor U2932 (N_2932,N_2038,N_1183);
or U2933 (N_2933,N_1069,N_1877);
or U2934 (N_2934,N_970,N_761);
and U2935 (N_2935,N_1002,N_181);
xnor U2936 (N_2936,N_585,N_2422);
and U2937 (N_2937,N_326,N_609);
nand U2938 (N_2938,N_716,N_1794);
xor U2939 (N_2939,N_289,N_2187);
and U2940 (N_2940,N_1982,N_1023);
nand U2941 (N_2941,N_193,N_916);
and U2942 (N_2942,N_2128,N_1812);
xnor U2943 (N_2943,N_1986,N_1239);
nor U2944 (N_2944,N_320,N_1093);
xnor U2945 (N_2945,N_1948,N_244);
nand U2946 (N_2946,N_726,N_395);
nor U2947 (N_2947,N_1860,N_1738);
nor U2948 (N_2948,N_1221,N_1670);
or U2949 (N_2949,N_1980,N_24);
or U2950 (N_2950,N_1308,N_169);
and U2951 (N_2951,N_2241,N_334);
and U2952 (N_2952,N_1919,N_459);
nand U2953 (N_2953,N_1835,N_269);
or U2954 (N_2954,N_768,N_1632);
nand U2955 (N_2955,N_1722,N_386);
nor U2956 (N_2956,N_540,N_174);
nand U2957 (N_2957,N_1995,N_1237);
or U2958 (N_2958,N_1140,N_1137);
xnor U2959 (N_2959,N_152,N_1382);
and U2960 (N_2960,N_2494,N_100);
nor U2961 (N_2961,N_123,N_1413);
or U2962 (N_2962,N_1871,N_881);
xnor U2963 (N_2963,N_719,N_247);
nand U2964 (N_2964,N_2385,N_2233);
and U2965 (N_2965,N_651,N_210);
and U2966 (N_2966,N_1484,N_1171);
and U2967 (N_2967,N_1530,N_2157);
nor U2968 (N_2968,N_327,N_654);
nor U2969 (N_2969,N_2015,N_2265);
or U2970 (N_2970,N_1707,N_835);
nand U2971 (N_2971,N_1580,N_1196);
xor U2972 (N_2972,N_1975,N_1055);
xnor U2973 (N_2973,N_791,N_718);
or U2974 (N_2974,N_1978,N_44);
and U2975 (N_2975,N_1493,N_1671);
xor U2976 (N_2976,N_387,N_819);
and U2977 (N_2977,N_204,N_647);
xor U2978 (N_2978,N_329,N_230);
nor U2979 (N_2979,N_1819,N_2272);
and U2980 (N_2980,N_1443,N_491);
and U2981 (N_2981,N_677,N_401);
xor U2982 (N_2982,N_951,N_1149);
nand U2983 (N_2983,N_1325,N_1679);
and U2984 (N_2984,N_422,N_2148);
nor U2985 (N_2985,N_1697,N_879);
and U2986 (N_2986,N_1870,N_922);
nand U2987 (N_2987,N_1780,N_432);
or U2988 (N_2988,N_1080,N_1849);
nor U2989 (N_2989,N_1555,N_1444);
nand U2990 (N_2990,N_960,N_969);
nor U2991 (N_2991,N_2404,N_1172);
or U2992 (N_2992,N_1123,N_810);
nor U2993 (N_2993,N_1065,N_2198);
nor U2994 (N_2994,N_132,N_598);
and U2995 (N_2995,N_2165,N_1816);
nand U2996 (N_2996,N_393,N_1730);
nor U2997 (N_2997,N_837,N_2119);
nand U2998 (N_2998,N_660,N_1314);
or U2999 (N_2999,N_975,N_99);
nand U3000 (N_3000,N_872,N_2026);
and U3001 (N_3001,N_1013,N_1997);
nor U3002 (N_3002,N_562,N_591);
and U3003 (N_3003,N_1748,N_1200);
and U3004 (N_3004,N_1566,N_42);
and U3005 (N_3005,N_1129,N_2489);
nor U3006 (N_3006,N_362,N_520);
nand U3007 (N_3007,N_404,N_1681);
xnor U3008 (N_3008,N_1846,N_658);
or U3009 (N_3009,N_1752,N_64);
nand U3010 (N_3010,N_1415,N_2236);
xnor U3011 (N_3011,N_2349,N_605);
nor U3012 (N_3012,N_618,N_1295);
and U3013 (N_3013,N_1193,N_1502);
nand U3014 (N_3014,N_348,N_766);
nand U3015 (N_3015,N_376,N_1019);
and U3016 (N_3016,N_1668,N_1438);
and U3017 (N_3017,N_2104,N_498);
nand U3018 (N_3018,N_347,N_2286);
xor U3019 (N_3019,N_1499,N_542);
or U3020 (N_3020,N_929,N_1751);
and U3021 (N_3021,N_1814,N_309);
nor U3022 (N_3022,N_212,N_949);
and U3023 (N_3023,N_1490,N_1667);
nor U3024 (N_3024,N_1528,N_67);
nor U3025 (N_3025,N_1791,N_299);
and U3026 (N_3026,N_1750,N_1259);
xor U3027 (N_3027,N_891,N_1965);
and U3028 (N_3028,N_857,N_474);
nand U3029 (N_3029,N_2423,N_1468);
nor U3030 (N_3030,N_850,N_412);
or U3031 (N_3031,N_2386,N_1663);
and U3032 (N_3032,N_1297,N_1777);
nand U3033 (N_3033,N_333,N_1962);
and U3034 (N_3034,N_1943,N_1386);
or U3035 (N_3035,N_1203,N_1301);
xor U3036 (N_3036,N_678,N_2042);
nor U3037 (N_3037,N_1232,N_1287);
or U3038 (N_3038,N_276,N_1776);
or U3039 (N_3039,N_1702,N_1859);
nand U3040 (N_3040,N_1099,N_2465);
nand U3041 (N_3041,N_1109,N_1888);
xnor U3042 (N_3042,N_671,N_1025);
nor U3043 (N_3043,N_1825,N_1909);
and U3044 (N_3044,N_762,N_702);
nor U3045 (N_3045,N_304,N_2229);
nor U3046 (N_3046,N_2142,N_1578);
xnor U3047 (N_3047,N_1133,N_932);
xor U3048 (N_3048,N_725,N_363);
nor U3049 (N_3049,N_2127,N_2384);
nand U3050 (N_3050,N_1257,N_547);
nand U3051 (N_3051,N_2,N_820);
nand U3052 (N_3052,N_2416,N_1725);
or U3053 (N_3053,N_1519,N_1054);
xnor U3054 (N_3054,N_266,N_1481);
or U3055 (N_3055,N_1267,N_1579);
and U3056 (N_3056,N_2444,N_1178);
nand U3057 (N_3057,N_2255,N_2230);
or U3058 (N_3058,N_197,N_2320);
xnor U3059 (N_3059,N_1101,N_814);
nor U3060 (N_3060,N_1552,N_1241);
nor U3061 (N_3061,N_71,N_232);
nor U3062 (N_3062,N_1960,N_447);
nand U3063 (N_3063,N_330,N_300);
nor U3064 (N_3064,N_2011,N_1284);
and U3065 (N_3065,N_182,N_859);
nor U3066 (N_3066,N_883,N_1256);
xor U3067 (N_3067,N_2341,N_79);
nand U3068 (N_3068,N_1700,N_0);
xnor U3069 (N_3069,N_2350,N_1810);
and U3070 (N_3070,N_1678,N_275);
nor U3071 (N_3071,N_1446,N_906);
nor U3072 (N_3072,N_1692,N_1569);
and U3073 (N_3073,N_1694,N_357);
nand U3074 (N_3074,N_2247,N_1603);
nand U3075 (N_3075,N_890,N_2113);
nor U3076 (N_3076,N_2056,N_1098);
or U3077 (N_3077,N_1534,N_1973);
and U3078 (N_3078,N_344,N_1361);
and U3079 (N_3079,N_33,N_832);
or U3080 (N_3080,N_240,N_1521);
and U3081 (N_3081,N_2257,N_470);
and U3082 (N_3082,N_2258,N_1182);
or U3083 (N_3083,N_1084,N_1563);
nor U3084 (N_3084,N_43,N_1598);
and U3085 (N_3085,N_1983,N_1620);
xnor U3086 (N_3086,N_1568,N_2062);
or U3087 (N_3087,N_1984,N_1328);
xnor U3088 (N_3088,N_2457,N_1236);
or U3089 (N_3089,N_118,N_2221);
xor U3090 (N_3090,N_146,N_2461);
nand U3091 (N_3091,N_1610,N_639);
and U3092 (N_3092,N_1190,N_2149);
nand U3093 (N_3093,N_2109,N_1733);
nand U3094 (N_3094,N_1254,N_2276);
xnor U3095 (N_3095,N_2279,N_793);
and U3096 (N_3096,N_321,N_2072);
and U3097 (N_3097,N_1334,N_1388);
xnor U3098 (N_3098,N_2114,N_261);
and U3099 (N_3099,N_2335,N_663);
or U3100 (N_3100,N_202,N_120);
nor U3101 (N_3101,N_1377,N_622);
xnor U3102 (N_3102,N_619,N_429);
and U3103 (N_3103,N_1273,N_1326);
or U3104 (N_3104,N_1719,N_53);
xnor U3105 (N_3105,N_1152,N_32);
or U3106 (N_3106,N_58,N_781);
nor U3107 (N_3107,N_1593,N_1205);
nor U3108 (N_3108,N_902,N_2409);
and U3109 (N_3109,N_557,N_1268);
and U3110 (N_3110,N_1202,N_461);
nor U3111 (N_3111,N_743,N_1661);
xor U3112 (N_3112,N_1474,N_1110);
nand U3113 (N_3113,N_1944,N_650);
or U3114 (N_3114,N_1896,N_2374);
nand U3115 (N_3115,N_1165,N_60);
nor U3116 (N_3116,N_160,N_194);
or U3117 (N_3117,N_278,N_220);
xnor U3118 (N_3118,N_1994,N_1766);
and U3119 (N_3119,N_1595,N_403);
xnor U3120 (N_3120,N_1250,N_472);
or U3121 (N_3121,N_838,N_235);
or U3122 (N_3122,N_1253,N_1934);
xnor U3123 (N_3123,N_560,N_157);
or U3124 (N_3124,N_1118,N_617);
xnor U3125 (N_3125,N_23,N_259);
nand U3126 (N_3126,N_796,N_381);
and U3127 (N_3127,N_439,N_2126);
and U3128 (N_3128,N_1914,N_10);
or U3129 (N_3129,N_2107,N_2464);
xnor U3130 (N_3130,N_1646,N_2329);
or U3131 (N_3131,N_21,N_1676);
nand U3132 (N_3132,N_675,N_992);
or U3133 (N_3133,N_335,N_1154);
and U3134 (N_3134,N_808,N_833);
nor U3135 (N_3135,N_1075,N_2390);
and U3136 (N_3136,N_92,N_2153);
xnor U3137 (N_3137,N_1597,N_2379);
xnor U3138 (N_3138,N_2387,N_503);
and U3139 (N_3139,N_756,N_280);
and U3140 (N_3140,N_1740,N_2087);
nand U3141 (N_3141,N_2452,N_94);
nor U3142 (N_3142,N_2453,N_338);
nand U3143 (N_3143,N_1157,N_341);
nor U3144 (N_3144,N_34,N_1029);
nor U3145 (N_3145,N_1128,N_2389);
or U3146 (N_3146,N_1318,N_2487);
or U3147 (N_3147,N_586,N_1755);
nand U3148 (N_3148,N_759,N_1693);
nand U3149 (N_3149,N_65,N_479);
nor U3150 (N_3150,N_1479,N_358);
and U3151 (N_3151,N_1244,N_1275);
nor U3152 (N_3152,N_523,N_2017);
and U3153 (N_3153,N_2086,N_2299);
or U3154 (N_3154,N_250,N_2174);
xor U3155 (N_3155,N_398,N_2146);
xnor U3156 (N_3156,N_2359,N_1599);
xnor U3157 (N_3157,N_2179,N_312);
or U3158 (N_3158,N_2009,N_1957);
xor U3159 (N_3159,N_423,N_688);
or U3160 (N_3160,N_2238,N_1645);
and U3161 (N_3161,N_2476,N_977);
xor U3162 (N_3162,N_2124,N_2362);
xor U3163 (N_3163,N_1303,N_421);
and U3164 (N_3164,N_1850,N_511);
nor U3165 (N_3165,N_991,N_980);
nor U3166 (N_3166,N_96,N_443);
nand U3167 (N_3167,N_15,N_2092);
nand U3168 (N_3168,N_1543,N_2493);
and U3169 (N_3169,N_684,N_1884);
and U3170 (N_3170,N_1142,N_572);
nor U3171 (N_3171,N_670,N_2180);
and U3172 (N_3172,N_668,N_1641);
nor U3173 (N_3173,N_2022,N_2018);
nor U3174 (N_3174,N_1464,N_1210);
or U3175 (N_3175,N_1765,N_2381);
and U3176 (N_3176,N_1271,N_2201);
xnor U3177 (N_3177,N_440,N_2266);
nor U3178 (N_3178,N_119,N_365);
nand U3179 (N_3179,N_1245,N_467);
or U3180 (N_3180,N_512,N_1771);
and U3181 (N_3181,N_2450,N_998);
or U3182 (N_3182,N_1485,N_493);
xor U3183 (N_3183,N_2284,N_80);
and U3184 (N_3184,N_1745,N_601);
nand U3185 (N_3185,N_2308,N_729);
xnor U3186 (N_3186,N_2005,N_813);
nand U3187 (N_3187,N_580,N_2129);
and U3188 (N_3188,N_1544,N_1887);
and U3189 (N_3189,N_509,N_853);
nor U3190 (N_3190,N_958,N_1188);
and U3191 (N_3191,N_526,N_1963);
nor U3192 (N_3192,N_1841,N_2152);
and U3193 (N_3193,N_1472,N_2285);
nor U3194 (N_3194,N_807,N_2061);
nand U3195 (N_3195,N_626,N_1600);
nand U3196 (N_3196,N_779,N_590);
or U3197 (N_3197,N_1876,N_2460);
or U3198 (N_3198,N_900,N_1619);
nor U3199 (N_3199,N_389,N_373);
xnor U3200 (N_3200,N_1854,N_999);
or U3201 (N_3201,N_102,N_674);
or U3202 (N_3202,N_303,N_238);
nand U3203 (N_3203,N_1163,N_541);
nand U3204 (N_3204,N_483,N_1211);
nand U3205 (N_3205,N_1195,N_87);
or U3206 (N_3206,N_2166,N_90);
nand U3207 (N_3207,N_1992,N_1509);
and U3208 (N_3208,N_243,N_2420);
nand U3209 (N_3209,N_1625,N_2040);
nor U3210 (N_3210,N_1754,N_435);
nor U3211 (N_3211,N_1977,N_1126);
xor U3212 (N_3212,N_2135,N_434);
nor U3213 (N_3213,N_865,N_2485);
or U3214 (N_3214,N_1258,N_1265);
nor U3215 (N_3215,N_933,N_78);
nor U3216 (N_3216,N_2070,N_1998);
nand U3217 (N_3217,N_1144,N_1690);
or U3218 (N_3218,N_1199,N_1380);
nor U3219 (N_3219,N_615,N_683);
xnor U3220 (N_3220,N_686,N_1932);
or U3221 (N_3221,N_1845,N_172);
xnor U3222 (N_3222,N_908,N_1478);
and U3223 (N_3223,N_774,N_2068);
nor U3224 (N_3224,N_2292,N_1942);
xnor U3225 (N_3225,N_2118,N_867);
nand U3226 (N_3226,N_264,N_2144);
and U3227 (N_3227,N_70,N_82);
xor U3228 (N_3228,N_973,N_714);
or U3229 (N_3229,N_164,N_127);
and U3230 (N_3230,N_248,N_1503);
nor U3231 (N_3231,N_1851,N_502);
or U3232 (N_3232,N_831,N_2253);
xnor U3233 (N_3233,N_1092,N_2076);
and U3234 (N_3234,N_322,N_57);
or U3235 (N_3235,N_614,N_1760);
nor U3236 (N_3236,N_2106,N_168);
xor U3237 (N_3237,N_298,N_31);
xnor U3238 (N_3238,N_1400,N_2330);
nor U3239 (N_3239,N_1001,N_866);
nor U3240 (N_3240,N_2440,N_2051);
xnor U3241 (N_3241,N_1433,N_907);
or U3242 (N_3242,N_816,N_1916);
and U3243 (N_3243,N_1219,N_1938);
nor U3244 (N_3244,N_982,N_2246);
or U3245 (N_3245,N_1475,N_47);
or U3246 (N_3246,N_794,N_2361);
nor U3247 (N_3247,N_245,N_1669);
and U3248 (N_3248,N_1802,N_887);
or U3249 (N_3249,N_161,N_1954);
or U3250 (N_3250,N_111,N_595);
nand U3251 (N_3251,N_496,N_221);
and U3252 (N_3252,N_2155,N_2090);
or U3253 (N_3253,N_1891,N_2305);
and U3254 (N_3254,N_1470,N_2371);
nand U3255 (N_3255,N_55,N_773);
nand U3256 (N_3256,N_844,N_465);
nand U3257 (N_3257,N_1937,N_1788);
nor U3258 (N_3258,N_1483,N_2498);
nand U3259 (N_3259,N_2343,N_870);
nor U3260 (N_3260,N_384,N_2393);
or U3261 (N_3261,N_1639,N_545);
nand U3262 (N_3262,N_286,N_1811);
and U3263 (N_3263,N_1018,N_2177);
xnor U3264 (N_3264,N_789,N_1024);
nor U3265 (N_3265,N_2250,N_1207);
or U3266 (N_3266,N_2325,N_409);
xnor U3267 (N_3267,N_445,N_629);
and U3268 (N_3268,N_1606,N_928);
nor U3269 (N_3269,N_501,N_612);
nor U3270 (N_3270,N_1547,N_821);
xor U3271 (N_3271,N_1143,N_1635);
or U3272 (N_3272,N_1538,N_45);
xnor U3273 (N_3273,N_1175,N_1037);
nand U3274 (N_3274,N_2053,N_1471);
nand U3275 (N_3275,N_2372,N_1594);
nand U3276 (N_3276,N_1372,N_569);
nor U3277 (N_3277,N_1278,N_2354);
xnor U3278 (N_3278,N_153,N_2199);
and U3279 (N_3279,N_1302,N_1167);
nand U3280 (N_3280,N_1653,N_812);
nor U3281 (N_3281,N_2023,N_1837);
xor U3282 (N_3282,N_227,N_1111);
nor U3283 (N_3283,N_698,N_588);
or U3284 (N_3284,N_1224,N_817);
and U3285 (N_3285,N_1442,N_187);
xnor U3286 (N_3286,N_2178,N_868);
and U3287 (N_3287,N_2363,N_1120);
nor U3288 (N_3288,N_1404,N_2301);
and U3289 (N_3289,N_2316,N_638);
xnor U3290 (N_3290,N_1790,N_1323);
xnor U3291 (N_3291,N_1116,N_1039);
nor U3292 (N_3292,N_1517,N_480);
or U3293 (N_3293,N_419,N_26);
or U3294 (N_3294,N_1032,N_1076);
xnor U3295 (N_3295,N_1864,N_4);
xor U3296 (N_3296,N_2474,N_988);
xor U3297 (N_3297,N_713,N_1616);
and U3298 (N_3298,N_2002,N_251);
nand U3299 (N_3299,N_144,N_2348);
and U3300 (N_3300,N_192,N_566);
or U3301 (N_3301,N_1546,N_554);
xnor U3302 (N_3302,N_450,N_324);
xor U3303 (N_3303,N_1623,N_1406);
xor U3304 (N_3304,N_1026,N_518);
nor U3305 (N_3305,N_1135,N_911);
nand U3306 (N_3306,N_1666,N_2020);
nor U3307 (N_3307,N_226,N_1827);
and U3308 (N_3308,N_464,N_573);
nor U3309 (N_3309,N_1747,N_2059);
xnor U3310 (N_3310,N_301,N_2028);
nand U3311 (N_3311,N_81,N_1017);
nand U3312 (N_3312,N_2312,N_1390);
nand U3313 (N_3313,N_1430,N_349);
nor U3314 (N_3314,N_383,N_555);
and U3315 (N_3315,N_1586,N_1749);
xor U3316 (N_3316,N_1247,N_46);
nand U3317 (N_3317,N_1764,N_1408);
nand U3318 (N_3318,N_2050,N_506);
and U3319 (N_3319,N_1112,N_74);
or U3320 (N_3320,N_352,N_945);
nor U3321 (N_3321,N_963,N_1341);
and U3322 (N_3322,N_236,N_1976);
and U3323 (N_3323,N_62,N_1252);
xor U3324 (N_3324,N_1581,N_1520);
and U3325 (N_3325,N_63,N_490);
or U3326 (N_3326,N_1330,N_695);
xnor U3327 (N_3327,N_596,N_2081);
nand U3328 (N_3328,N_2310,N_2037);
or U3329 (N_3329,N_2168,N_1872);
or U3330 (N_3330,N_1838,N_1542);
nor U3331 (N_3331,N_1783,N_1714);
nand U3332 (N_3332,N_871,N_452);
nor U3333 (N_3333,N_1020,N_993);
nand U3334 (N_3334,N_1044,N_211);
xnor U3335 (N_3335,N_1005,N_1270);
and U3336 (N_3336,N_1279,N_457);
nand U3337 (N_3337,N_1974,N_207);
xor U3338 (N_3338,N_2000,N_961);
nor U3339 (N_3339,N_1310,N_1272);
nand U3340 (N_3340,N_1618,N_1550);
and U3341 (N_3341,N_291,N_2134);
and U3342 (N_3342,N_1658,N_2077);
or U3343 (N_3343,N_1145,N_446);
xor U3344 (N_3344,N_1465,N_1571);
and U3345 (N_3345,N_823,N_2407);
and U3346 (N_3346,N_897,N_1873);
xor U3347 (N_3347,N_530,N_971);
nor U3348 (N_3348,N_2188,N_661);
and U3349 (N_3349,N_1056,N_1704);
xnor U3350 (N_3350,N_1091,N_346);
nor U3351 (N_3351,N_354,N_2306);
nand U3352 (N_3352,N_1880,N_1067);
nor U3353 (N_3353,N_575,N_1723);
nor U3354 (N_3354,N_1508,N_1820);
or U3355 (N_3355,N_1354,N_2164);
xnor U3356 (N_3356,N_2049,N_809);
nand U3357 (N_3357,N_1573,N_1946);
nor U3358 (N_3358,N_1772,N_2356);
xor U3359 (N_3359,N_125,N_1192);
nor U3360 (N_3360,N_2447,N_223);
nor U3361 (N_3361,N_1709,N_178);
and U3362 (N_3362,N_2239,N_1636);
or U3363 (N_3363,N_2499,N_2103);
nand U3364 (N_3364,N_1046,N_292);
and U3365 (N_3365,N_948,N_1921);
or U3366 (N_3366,N_777,N_388);
and U3367 (N_3367,N_2251,N_1677);
xnor U3368 (N_3368,N_2315,N_1863);
nor U3369 (N_3369,N_1286,N_2111);
or U3370 (N_3370,N_728,N_525);
or U3371 (N_3371,N_260,N_2406);
or U3372 (N_3372,N_1897,N_860);
nor U3373 (N_3373,N_537,N_2083);
nand U3374 (N_3374,N_2314,N_1000);
xor U3375 (N_3375,N_2396,N_1359);
nand U3376 (N_3376,N_790,N_1804);
nor U3377 (N_3377,N_987,N_246);
nor U3378 (N_3378,N_514,N_214);
xor U3379 (N_3379,N_2084,N_1650);
and U3380 (N_3380,N_1949,N_801);
or U3381 (N_3381,N_640,N_1931);
nor U3382 (N_3382,N_2105,N_27);
or U3383 (N_3383,N_1155,N_1062);
nand U3384 (N_3384,N_155,N_656);
nand U3385 (N_3385,N_369,N_2120);
and U3386 (N_3386,N_1393,N_2412);
nor U3387 (N_3387,N_2382,N_672);
or U3388 (N_3388,N_355,N_1899);
nor U3389 (N_3389,N_927,N_876);
nand U3390 (N_3390,N_1987,N_979);
and U3391 (N_3391,N_1832,N_1925);
nand U3392 (N_3392,N_1052,N_2252);
and U3393 (N_3393,N_1691,N_1357);
xnor U3394 (N_3394,N_1637,N_1180);
and U3395 (N_3395,N_1806,N_1904);
or U3396 (N_3396,N_918,N_755);
and U3397 (N_3397,N_1235,N_1260);
and U3398 (N_3398,N_926,N_1642);
nand U3399 (N_3399,N_2456,N_1830);
nor U3400 (N_3400,N_1233,N_1900);
nor U3401 (N_3401,N_1449,N_984);
and U3402 (N_3402,N_1970,N_1034);
nand U3403 (N_3403,N_108,N_1720);
xor U3404 (N_3404,N_2138,N_1801);
xor U3405 (N_3405,N_1596,N_175);
and U3406 (N_3406,N_2176,N_1829);
xor U3407 (N_3407,N_1306,N_1398);
nor U3408 (N_3408,N_666,N_1218);
xor U3409 (N_3409,N_2132,N_1077);
xnor U3410 (N_3410,N_1147,N_1648);
nor U3411 (N_3411,N_485,N_2437);
nand U3412 (N_3412,N_131,N_2357);
nand U3413 (N_3413,N_935,N_2167);
and U3414 (N_3414,N_1136,N_1385);
and U3415 (N_3415,N_1451,N_442);
or U3416 (N_3416,N_167,N_1266);
xnor U3417 (N_3417,N_2159,N_2455);
or U3418 (N_3418,N_1280,N_1857);
or U3419 (N_3419,N_1059,N_1917);
and U3420 (N_3420,N_1074,N_1248);
nor U3421 (N_3421,N_1774,N_748);
nand U3422 (N_3422,N_370,N_946);
nor U3423 (N_3423,N_1910,N_93);
nand U3424 (N_3424,N_315,N_1307);
nand U3425 (N_3425,N_1313,N_1352);
nand U3426 (N_3426,N_2309,N_1529);
nand U3427 (N_3427,N_1647,N_180);
and U3428 (N_3428,N_2400,N_1971);
and U3429 (N_3429,N_2227,N_2122);
nor U3430 (N_3430,N_648,N_2271);
nor U3431 (N_3431,N_625,N_416);
or U3432 (N_3432,N_1757,N_1198);
nor U3433 (N_3433,N_1969,N_1630);
xnor U3434 (N_3434,N_2065,N_2495);
or U3435 (N_3435,N_256,N_1293);
xor U3436 (N_3436,N_2435,N_1083);
xor U3437 (N_3437,N_431,N_2224);
nand U3438 (N_3438,N_1496,N_533);
nand U3439 (N_3439,N_2462,N_1159);
xor U3440 (N_3440,N_707,N_1309);
and U3441 (N_3441,N_2344,N_2069);
xnor U3442 (N_3442,N_1176,N_13);
nor U3443 (N_3443,N_145,N_696);
or U3444 (N_3444,N_3,N_110);
nor U3445 (N_3445,N_682,N_930);
nor U3446 (N_3446,N_463,N_1263);
and U3447 (N_3447,N_1527,N_862);
xor U3448 (N_3448,N_141,N_834);
nor U3449 (N_3449,N_915,N_1584);
nand U3450 (N_3450,N_1045,N_371);
xnor U3451 (N_3451,N_1936,N_113);
and U3452 (N_3452,N_1033,N_2353);
nand U3453 (N_3453,N_1990,N_1070);
or U3454 (N_3454,N_1822,N_1340);
and U3455 (N_3455,N_936,N_2063);
or U3456 (N_3456,N_1885,N_1461);
xor U3457 (N_3457,N_1511,N_2052);
and U3458 (N_3458,N_1277,N_2468);
nor U3459 (N_3459,N_2469,N_827);
xnor U3460 (N_3460,N_950,N_1319);
or U3461 (N_3461,N_2082,N_1403);
nor U3462 (N_3462,N_1495,N_272);
nor U3463 (N_3463,N_1602,N_449);
xnor U3464 (N_3464,N_1933,N_1146);
nor U3465 (N_3465,N_736,N_2408);
xnor U3466 (N_3466,N_1255,N_1291);
and U3467 (N_3467,N_765,N_302);
nand U3468 (N_3468,N_1815,N_1869);
xnor U3469 (N_3469,N_2421,N_307);
nand U3470 (N_3470,N_996,N_2057);
or U3471 (N_3471,N_408,N_1524);
nor U3472 (N_3472,N_1113,N_2342);
and U3473 (N_3473,N_582,N_968);
xor U3474 (N_3474,N_1583,N_983);
nand U3475 (N_3475,N_2080,N_643);
nor U3476 (N_3476,N_1732,N_126);
nand U3477 (N_3477,N_288,N_1358);
xor U3478 (N_3478,N_692,N_2458);
or U3479 (N_3479,N_888,N_2441);
nor U3480 (N_3480,N_1321,N_673);
nand U3481 (N_3481,N_1711,N_2163);
nand U3482 (N_3482,N_2217,N_263);
nand U3483 (N_3483,N_343,N_1169);
xor U3484 (N_3484,N_106,N_1383);
and U3485 (N_3485,N_285,N_1865);
nor U3486 (N_3486,N_2141,N_1926);
and U3487 (N_3487,N_1775,N_957);
and U3488 (N_3488,N_1049,N_2262);
or U3489 (N_3489,N_1609,N_1068);
or U3490 (N_3490,N_576,N_2430);
nor U3491 (N_3491,N_185,N_54);
nand U3492 (N_3492,N_1096,N_2024);
or U3493 (N_3493,N_2206,N_350);
and U3494 (N_3494,N_2088,N_704);
nor U3495 (N_3495,N_2269,N_2281);
or U3496 (N_3496,N_2333,N_2101);
nand U3497 (N_3497,N_538,N_1230);
or U3498 (N_3498,N_1453,N_1130);
xnor U3499 (N_3499,N_535,N_603);
and U3500 (N_3500,N_727,N_104);
or U3501 (N_3501,N_189,N_2079);
nor U3502 (N_3502,N_2376,N_653);
and U3503 (N_3503,N_417,N_400);
and U3504 (N_3504,N_747,N_1454);
or U3505 (N_3505,N_710,N_556);
xor U3506 (N_3506,N_2190,N_1491);
nor U3507 (N_3507,N_854,N_723);
and U3508 (N_3508,N_592,N_466);
and U3509 (N_3509,N_1095,N_2280);
or U3510 (N_3510,N_752,N_1355);
nor U3511 (N_3511,N_1378,N_1659);
nor U3512 (N_3512,N_877,N_121);
xnor U3513 (N_3513,N_1201,N_1315);
nor U3514 (N_3514,N_1726,N_1395);
and U3515 (N_3515,N_1560,N_2154);
or U3516 (N_3516,N_2058,N_806);
nand U3517 (N_3517,N_402,N_1558);
nor U3518 (N_3518,N_858,N_641);
and U3519 (N_3519,N_41,N_458);
or U3520 (N_3520,N_630,N_1214);
xor U3521 (N_3521,N_451,N_861);
xor U3522 (N_3522,N_1721,N_1324);
nor U3523 (N_3523,N_940,N_39);
and U3524 (N_3524,N_1102,N_38);
nor U3525 (N_3525,N_899,N_456);
or U3526 (N_3526,N_2364,N_720);
nand U3527 (N_3527,N_1384,N_1903);
nor U3528 (N_3528,N_128,N_1787);
xor U3529 (N_3529,N_561,N_2019);
or U3530 (N_3530,N_191,N_952);
nor U3531 (N_3531,N_165,N_252);
or U3532 (N_3532,N_1038,N_2195);
nor U3533 (N_3533,N_1770,N_1424);
xor U3534 (N_3534,N_1429,N_646);
and U3535 (N_3535,N_1500,N_2290);
nand U3536 (N_3536,N_1227,N_2130);
xor U3537 (N_3537,N_420,N_239);
nor U3538 (N_3538,N_637,N_546);
and U3539 (N_3539,N_208,N_258);
nand U3540 (N_3540,N_1186,N_1848);
nand U3541 (N_3541,N_1889,N_1072);
and U3542 (N_3542,N_1360,N_177);
nor U3543 (N_3543,N_1320,N_2491);
or U3544 (N_3544,N_296,N_2123);
nand U3545 (N_3545,N_2012,N_1913);
xnor U3546 (N_3546,N_17,N_2436);
and U3547 (N_3547,N_56,N_895);
xor U3548 (N_3548,N_1249,N_297);
nand U3549 (N_3549,N_2278,N_1821);
nand U3550 (N_3550,N_129,N_1066);
or U3551 (N_3551,N_1967,N_137);
nand U3552 (N_3552,N_441,N_705);
nor U3553 (N_3553,N_2145,N_1989);
xor U3554 (N_3554,N_1966,N_2196);
or U3555 (N_3555,N_1088,N_721);
nor U3556 (N_3556,N_1153,N_2202);
xor U3557 (N_3557,N_1985,N_1048);
or U3558 (N_3558,N_610,N_1);
xnor U3559 (N_3559,N_1139,N_1488);
and U3560 (N_3560,N_1104,N_706);
xnor U3561 (N_3561,N_14,N_254);
nor U3562 (N_3562,N_1892,N_972);
nor U3563 (N_3563,N_944,N_1427);
or U3564 (N_3564,N_331,N_1298);
nand U3565 (N_3565,N_73,N_1847);
nand U3566 (N_3566,N_1106,N_1031);
nor U3567 (N_3567,N_1856,N_2117);
and U3568 (N_3568,N_97,N_1945);
xnor U3569 (N_3569,N_1656,N_1657);
nor U3570 (N_3570,N_994,N_1988);
and U3571 (N_3571,N_2182,N_1617);
or U3572 (N_3572,N_162,N_59);
and U3573 (N_3573,N_1796,N_2161);
xnor U3574 (N_3574,N_1416,N_293);
and U3575 (N_3575,N_1626,N_1370);
and U3576 (N_3576,N_1525,N_35);
or U3577 (N_3577,N_18,N_815);
and U3578 (N_3578,N_1299,N_2228);
or U3579 (N_3579,N_107,N_893);
and U3580 (N_3580,N_1706,N_2158);
and U3581 (N_3581,N_2136,N_1744);
and U3582 (N_3582,N_2322,N_1212);
nand U3583 (N_3583,N_2211,N_2317);
nand U3584 (N_3584,N_2331,N_437);
or U3585 (N_3585,N_1548,N_1425);
nand U3586 (N_3586,N_158,N_154);
nor U3587 (N_3587,N_1389,N_543);
xor U3588 (N_3588,N_1327,N_2067);
or U3589 (N_3589,N_1541,N_1708);
xnor U3590 (N_3590,N_1396,N_2303);
xor U3591 (N_3591,N_1868,N_428);
xnor U3592 (N_3592,N_1839,N_1078);
nand U3593 (N_3593,N_919,N_317);
and U3594 (N_3594,N_606,N_2029);
nor U3595 (N_3595,N_967,N_1510);
and U3596 (N_3596,N_2296,N_200);
and U3597 (N_3597,N_904,N_2208);
nand U3598 (N_3598,N_631,N_2415);
nor U3599 (N_3599,N_1649,N_171);
xor U3600 (N_3600,N_1522,N_1561);
or U3601 (N_3601,N_1349,N_1628);
nor U3602 (N_3602,N_406,N_2274);
or U3603 (N_3603,N_917,N_83);
nand U3604 (N_3604,N_1187,N_1368);
nor U3605 (N_3605,N_1834,N_1727);
xor U3606 (N_3606,N_914,N_1466);
nand U3607 (N_3607,N_711,N_1964);
and U3608 (N_3608,N_249,N_544);
xnor U3609 (N_3609,N_2432,N_1652);
nor U3610 (N_3610,N_873,N_1614);
or U3611 (N_3611,N_453,N_228);
xor U3612 (N_3612,N_2425,N_2481);
xor U3613 (N_3613,N_1028,N_378);
xor U3614 (N_3614,N_1125,N_1779);
nand U3615 (N_3615,N_1170,N_1955);
nor U3616 (N_3616,N_522,N_336);
nand U3617 (N_3617,N_147,N_1627);
nand U3618 (N_3618,N_1531,N_37);
or U3619 (N_3619,N_732,N_1016);
nand U3620 (N_3620,N_1381,N_170);
and U3621 (N_3621,N_2240,N_852);
xnor U3622 (N_3622,N_61,N_679);
or U3623 (N_3623,N_176,N_135);
xor U3624 (N_3624,N_2184,N_2439);
or U3625 (N_3625,N_253,N_319);
nor U3626 (N_3626,N_1114,N_1206);
nand U3627 (N_3627,N_1717,N_574);
or U3628 (N_3628,N_797,N_552);
nand U3629 (N_3629,N_1605,N_2467);
and U3630 (N_3630,N_138,N_712);
and U3631 (N_3631,N_1150,N_1753);
nand U3632 (N_3632,N_1426,N_84);
xnor U3633 (N_3633,N_788,N_731);
and U3634 (N_3634,N_1423,N_183);
nand U3635 (N_3635,N_1824,N_527);
nand U3636 (N_3636,N_1194,N_616);
xnor U3637 (N_3637,N_885,N_1498);
nand U3638 (N_3638,N_620,N_700);
nand U3639 (N_3639,N_229,N_738);
nor U3640 (N_3640,N_1894,N_1345);
xnor U3641 (N_3641,N_2417,N_1231);
nand U3642 (N_3642,N_2445,N_49);
nor U3643 (N_3643,N_1448,N_636);
and U3644 (N_3644,N_2287,N_959);
nor U3645 (N_3645,N_962,N_2254);
xnor U3646 (N_3646,N_1808,N_1161);
nor U3647 (N_3647,N_257,N_1557);
xnor U3648 (N_3648,N_783,N_2001);
xnor U3649 (N_3649,N_2446,N_1882);
and U3650 (N_3650,N_633,N_805);
or U3651 (N_3651,N_136,N_771);
xor U3652 (N_3652,N_1684,N_1240);
nor U3653 (N_3653,N_1660,N_1831);
and U3654 (N_3654,N_101,N_488);
or U3655 (N_3655,N_841,N_558);
nor U3656 (N_3656,N_624,N_757);
and U3657 (N_3657,N_1347,N_2139);
or U3658 (N_3658,N_2337,N_2486);
or U3659 (N_3659,N_380,N_1836);
and U3660 (N_3660,N_504,N_568);
or U3661 (N_3661,N_1915,N_1540);
xnor U3662 (N_3662,N_1792,N_749);
xor U3663 (N_3663,N_274,N_1928);
xnor U3664 (N_3664,N_571,N_1294);
or U3665 (N_3665,N_1878,N_222);
nor U3666 (N_3666,N_415,N_1526);
nor U3667 (N_3667,N_1364,N_803);
nor U3668 (N_3668,N_1348,N_2454);
and U3669 (N_3669,N_2183,N_1611);
or U3670 (N_3670,N_567,N_1473);
nand U3671 (N_3671,N_1022,N_224);
nand U3672 (N_3672,N_410,N_1761);
or U3673 (N_3673,N_1564,N_1895);
nand U3674 (N_3674,N_262,N_190);
nor U3675 (N_3675,N_1010,N_2025);
nand U3676 (N_3676,N_717,N_468);
nor U3677 (N_3677,N_1516,N_1134);
nand U3678 (N_3678,N_2242,N_2137);
and U3679 (N_3679,N_989,N_1317);
and U3680 (N_3680,N_375,N_681);
nor U3681 (N_3681,N_2073,N_693);
or U3682 (N_3682,N_2014,N_2324);
nand U3683 (N_3683,N_2414,N_2313);
nor U3684 (N_3684,N_1132,N_2394);
nor U3685 (N_3685,N_1533,N_103);
or U3686 (N_3686,N_924,N_1085);
xor U3687 (N_3687,N_2218,N_1131);
and U3688 (N_3688,N_476,N_934);
or U3689 (N_3689,N_764,N_438);
or U3690 (N_3690,N_332,N_1356);
or U3691 (N_3691,N_2346,N_30);
and U3692 (N_3692,N_1191,N_1173);
nor U3693 (N_3693,N_1035,N_2075);
nor U3694 (N_3694,N_1799,N_795);
nor U3695 (N_3695,N_1504,N_956);
and U3696 (N_3696,N_1551,N_909);
xnor U3697 (N_3697,N_337,N_786);
or U3698 (N_3698,N_1935,N_233);
xnor U3699 (N_3699,N_1342,N_219);
nor U3700 (N_3700,N_1809,N_1629);
nor U3701 (N_3701,N_2021,N_1343);
nor U3702 (N_3702,N_824,N_953);
or U3703 (N_3703,N_2369,N_277);
and U3704 (N_3704,N_1729,N_559);
or U3705 (N_3705,N_1467,N_1115);
nor U3706 (N_3706,N_1079,N_1715);
nand U3707 (N_3707,N_2223,N_1166);
xnor U3708 (N_3708,N_1117,N_2398);
nand U3709 (N_3709,N_20,N_1993);
nor U3710 (N_3710,N_1283,N_1003);
nand U3711 (N_3711,N_444,N_2125);
nand U3712 (N_3712,N_1833,N_822);
or U3713 (N_3713,N_2403,N_2340);
nand U3714 (N_3714,N_143,N_744);
xor U3715 (N_3715,N_1672,N_1576);
nor U3716 (N_3716,N_1274,N_687);
nand U3717 (N_3717,N_368,N_515);
and U3718 (N_3718,N_1742,N_1412);
nor U3719 (N_3719,N_1996,N_1350);
or U3720 (N_3720,N_1071,N_48);
xor U3721 (N_3721,N_2044,N_920);
and U3722 (N_3722,N_1434,N_2434);
or U3723 (N_3723,N_1337,N_894);
nand U3724 (N_3724,N_2492,N_754);
xor U3725 (N_3725,N_1486,N_1908);
nand U3726 (N_3726,N_2327,N_1604);
nand U3727 (N_3727,N_405,N_1476);
nand U3728 (N_3728,N_2339,N_1683);
nand U3729 (N_3729,N_2248,N_1682);
nand U3730 (N_3730,N_112,N_938);
nor U3731 (N_3731,N_1813,N_947);
xnor U3732 (N_3732,N_581,N_1778);
xor U3733 (N_3733,N_2443,N_1305);
xnor U3734 (N_3734,N_1414,N_134);
or U3735 (N_3735,N_737,N_1243);
and U3736 (N_3736,N_2150,N_116);
nor U3737 (N_3737,N_1886,N_849);
or U3738 (N_3738,N_72,N_2392);
xnor U3739 (N_3739,N_268,N_2326);
xor U3740 (N_3740,N_2140,N_2108);
xor U3741 (N_3741,N_2397,N_898);
nand U3742 (N_3742,N_2256,N_2378);
xnor U3743 (N_3743,N_1818,N_499);
and U3744 (N_3744,N_923,N_2488);
nor U3745 (N_3745,N_1782,N_583);
nand U3746 (N_3746,N_763,N_2419);
nand U3747 (N_3747,N_1613,N_2220);
xnor U3748 (N_3748,N_703,N_2060);
and U3749 (N_3749,N_385,N_1638);
nand U3750 (N_3750,N_570,N_1704);
xnor U3751 (N_3751,N_15,N_572);
nand U3752 (N_3752,N_462,N_1487);
nand U3753 (N_3753,N_1362,N_63);
nor U3754 (N_3754,N_196,N_2304);
xnor U3755 (N_3755,N_1533,N_192);
nand U3756 (N_3756,N_1018,N_866);
or U3757 (N_3757,N_1701,N_2303);
xnor U3758 (N_3758,N_2298,N_491);
xnor U3759 (N_3759,N_2441,N_1514);
nand U3760 (N_3760,N_2408,N_1865);
xor U3761 (N_3761,N_1205,N_468);
or U3762 (N_3762,N_1942,N_1113);
xor U3763 (N_3763,N_50,N_2165);
xnor U3764 (N_3764,N_1459,N_2054);
or U3765 (N_3765,N_1035,N_2387);
or U3766 (N_3766,N_1722,N_2269);
nor U3767 (N_3767,N_118,N_976);
or U3768 (N_3768,N_216,N_305);
nor U3769 (N_3769,N_886,N_2210);
and U3770 (N_3770,N_1678,N_1652);
and U3771 (N_3771,N_1176,N_1841);
nor U3772 (N_3772,N_2204,N_706);
or U3773 (N_3773,N_379,N_111);
and U3774 (N_3774,N_1270,N_1248);
or U3775 (N_3775,N_400,N_697);
or U3776 (N_3776,N_1814,N_1221);
nand U3777 (N_3777,N_1957,N_2042);
and U3778 (N_3778,N_1144,N_1511);
nand U3779 (N_3779,N_1771,N_1431);
nand U3780 (N_3780,N_280,N_538);
or U3781 (N_3781,N_1766,N_1666);
xnor U3782 (N_3782,N_843,N_2136);
nand U3783 (N_3783,N_2134,N_1030);
nand U3784 (N_3784,N_423,N_39);
or U3785 (N_3785,N_1531,N_277);
nor U3786 (N_3786,N_2147,N_1973);
xor U3787 (N_3787,N_916,N_1175);
nand U3788 (N_3788,N_826,N_750);
nor U3789 (N_3789,N_643,N_98);
nor U3790 (N_3790,N_352,N_125);
nand U3791 (N_3791,N_1740,N_1252);
nor U3792 (N_3792,N_1570,N_790);
xor U3793 (N_3793,N_2319,N_820);
and U3794 (N_3794,N_801,N_2499);
and U3795 (N_3795,N_2186,N_2472);
xor U3796 (N_3796,N_1739,N_493);
xnor U3797 (N_3797,N_880,N_1018);
nand U3798 (N_3798,N_1556,N_1501);
and U3799 (N_3799,N_1283,N_321);
nand U3800 (N_3800,N_1564,N_688);
nand U3801 (N_3801,N_2149,N_128);
or U3802 (N_3802,N_167,N_2365);
nor U3803 (N_3803,N_419,N_1635);
nor U3804 (N_3804,N_130,N_801);
and U3805 (N_3805,N_164,N_559);
xnor U3806 (N_3806,N_1780,N_623);
xnor U3807 (N_3807,N_1071,N_1955);
xnor U3808 (N_3808,N_1554,N_1911);
nand U3809 (N_3809,N_638,N_769);
and U3810 (N_3810,N_1563,N_1971);
nand U3811 (N_3811,N_42,N_1155);
xor U3812 (N_3812,N_1971,N_900);
or U3813 (N_3813,N_2087,N_172);
and U3814 (N_3814,N_945,N_576);
nand U3815 (N_3815,N_1611,N_2073);
nand U3816 (N_3816,N_2229,N_2354);
or U3817 (N_3817,N_1265,N_1366);
or U3818 (N_3818,N_37,N_23);
or U3819 (N_3819,N_2498,N_132);
or U3820 (N_3820,N_1969,N_1766);
nand U3821 (N_3821,N_1339,N_655);
xor U3822 (N_3822,N_2270,N_1594);
nand U3823 (N_3823,N_2240,N_1960);
nand U3824 (N_3824,N_212,N_1091);
or U3825 (N_3825,N_1364,N_810);
or U3826 (N_3826,N_2057,N_2157);
or U3827 (N_3827,N_1064,N_1445);
or U3828 (N_3828,N_38,N_1805);
and U3829 (N_3829,N_2481,N_508);
and U3830 (N_3830,N_1535,N_465);
and U3831 (N_3831,N_1400,N_1324);
xnor U3832 (N_3832,N_1463,N_2331);
or U3833 (N_3833,N_224,N_254);
nand U3834 (N_3834,N_1667,N_1419);
or U3835 (N_3835,N_59,N_1031);
or U3836 (N_3836,N_1309,N_1086);
xnor U3837 (N_3837,N_976,N_880);
nand U3838 (N_3838,N_853,N_1830);
xnor U3839 (N_3839,N_208,N_2144);
nor U3840 (N_3840,N_1527,N_203);
or U3841 (N_3841,N_1237,N_1784);
nand U3842 (N_3842,N_2458,N_1621);
or U3843 (N_3843,N_1435,N_2491);
and U3844 (N_3844,N_1130,N_1519);
xor U3845 (N_3845,N_245,N_1336);
or U3846 (N_3846,N_2437,N_522);
nand U3847 (N_3847,N_1409,N_695);
nand U3848 (N_3848,N_581,N_1930);
xor U3849 (N_3849,N_1110,N_890);
and U3850 (N_3850,N_977,N_1877);
nand U3851 (N_3851,N_1222,N_133);
nand U3852 (N_3852,N_1144,N_1940);
xnor U3853 (N_3853,N_1407,N_485);
xnor U3854 (N_3854,N_2492,N_1680);
nand U3855 (N_3855,N_1905,N_1831);
nand U3856 (N_3856,N_1868,N_1454);
or U3857 (N_3857,N_2313,N_1836);
or U3858 (N_3858,N_1146,N_1936);
nor U3859 (N_3859,N_898,N_175);
nor U3860 (N_3860,N_1758,N_731);
nor U3861 (N_3861,N_1095,N_823);
nand U3862 (N_3862,N_1866,N_685);
and U3863 (N_3863,N_2094,N_673);
xor U3864 (N_3864,N_1898,N_485);
xor U3865 (N_3865,N_747,N_2345);
nand U3866 (N_3866,N_1164,N_159);
xnor U3867 (N_3867,N_619,N_1716);
or U3868 (N_3868,N_319,N_2417);
or U3869 (N_3869,N_1657,N_669);
nor U3870 (N_3870,N_145,N_2024);
nand U3871 (N_3871,N_1294,N_453);
xor U3872 (N_3872,N_1359,N_480);
and U3873 (N_3873,N_617,N_2138);
and U3874 (N_3874,N_394,N_1834);
nand U3875 (N_3875,N_206,N_1001);
and U3876 (N_3876,N_753,N_901);
and U3877 (N_3877,N_90,N_1505);
nor U3878 (N_3878,N_2433,N_528);
nor U3879 (N_3879,N_627,N_1614);
and U3880 (N_3880,N_1048,N_126);
or U3881 (N_3881,N_1337,N_1688);
and U3882 (N_3882,N_2170,N_1828);
nor U3883 (N_3883,N_786,N_1242);
nand U3884 (N_3884,N_510,N_1649);
nor U3885 (N_3885,N_1550,N_2202);
nor U3886 (N_3886,N_771,N_1959);
and U3887 (N_3887,N_377,N_375);
nor U3888 (N_3888,N_305,N_2266);
nand U3889 (N_3889,N_600,N_78);
xor U3890 (N_3890,N_2362,N_1762);
nand U3891 (N_3891,N_2217,N_1254);
and U3892 (N_3892,N_1779,N_2029);
xor U3893 (N_3893,N_1126,N_2247);
and U3894 (N_3894,N_1271,N_1430);
and U3895 (N_3895,N_1934,N_906);
and U3896 (N_3896,N_2266,N_1160);
nand U3897 (N_3897,N_1518,N_1808);
nand U3898 (N_3898,N_2401,N_1311);
or U3899 (N_3899,N_1001,N_2380);
or U3900 (N_3900,N_1855,N_223);
nor U3901 (N_3901,N_1350,N_2177);
and U3902 (N_3902,N_846,N_2155);
and U3903 (N_3903,N_548,N_1655);
nor U3904 (N_3904,N_2455,N_1699);
nand U3905 (N_3905,N_1476,N_1174);
and U3906 (N_3906,N_2104,N_410);
nor U3907 (N_3907,N_1754,N_335);
or U3908 (N_3908,N_1776,N_12);
and U3909 (N_3909,N_1270,N_1521);
or U3910 (N_3910,N_1495,N_2470);
and U3911 (N_3911,N_1002,N_494);
nor U3912 (N_3912,N_1367,N_333);
xnor U3913 (N_3913,N_2158,N_1443);
and U3914 (N_3914,N_1166,N_2363);
nor U3915 (N_3915,N_734,N_1852);
xnor U3916 (N_3916,N_2048,N_1836);
nand U3917 (N_3917,N_1151,N_2346);
nor U3918 (N_3918,N_1889,N_1137);
nor U3919 (N_3919,N_2418,N_174);
xnor U3920 (N_3920,N_198,N_2014);
nand U3921 (N_3921,N_1323,N_678);
nand U3922 (N_3922,N_2173,N_1414);
and U3923 (N_3923,N_784,N_209);
and U3924 (N_3924,N_2,N_682);
or U3925 (N_3925,N_379,N_389);
nor U3926 (N_3926,N_1124,N_1819);
nor U3927 (N_3927,N_1007,N_1820);
nor U3928 (N_3928,N_2023,N_1732);
nand U3929 (N_3929,N_1031,N_1317);
nor U3930 (N_3930,N_937,N_2300);
nand U3931 (N_3931,N_775,N_2391);
nand U3932 (N_3932,N_345,N_193);
nor U3933 (N_3933,N_152,N_1366);
or U3934 (N_3934,N_2093,N_1697);
nor U3935 (N_3935,N_2081,N_594);
and U3936 (N_3936,N_1151,N_141);
or U3937 (N_3937,N_1775,N_104);
nor U3938 (N_3938,N_1814,N_1859);
or U3939 (N_3939,N_103,N_1909);
nand U3940 (N_3940,N_1264,N_107);
xor U3941 (N_3941,N_1070,N_268);
xnor U3942 (N_3942,N_338,N_1278);
and U3943 (N_3943,N_1580,N_2154);
and U3944 (N_3944,N_2439,N_1651);
and U3945 (N_3945,N_920,N_2360);
xnor U3946 (N_3946,N_2300,N_2094);
and U3947 (N_3947,N_1599,N_1073);
or U3948 (N_3948,N_383,N_1500);
nor U3949 (N_3949,N_146,N_1365);
and U3950 (N_3950,N_1406,N_298);
xnor U3951 (N_3951,N_1955,N_1387);
nor U3952 (N_3952,N_1578,N_1659);
and U3953 (N_3953,N_1200,N_1835);
nor U3954 (N_3954,N_1704,N_181);
or U3955 (N_3955,N_371,N_2245);
and U3956 (N_3956,N_2393,N_1761);
or U3957 (N_3957,N_2322,N_704);
nor U3958 (N_3958,N_2011,N_906);
xnor U3959 (N_3959,N_987,N_1807);
nand U3960 (N_3960,N_726,N_357);
nand U3961 (N_3961,N_2380,N_915);
nor U3962 (N_3962,N_1342,N_802);
nor U3963 (N_3963,N_2156,N_682);
nor U3964 (N_3964,N_2074,N_1209);
nand U3965 (N_3965,N_971,N_1805);
nand U3966 (N_3966,N_1577,N_488);
or U3967 (N_3967,N_933,N_1656);
or U3968 (N_3968,N_209,N_51);
nor U3969 (N_3969,N_1983,N_216);
nand U3970 (N_3970,N_476,N_1597);
nand U3971 (N_3971,N_71,N_1023);
nand U3972 (N_3972,N_2110,N_327);
nor U3973 (N_3973,N_34,N_955);
or U3974 (N_3974,N_2061,N_1155);
nor U3975 (N_3975,N_142,N_560);
and U3976 (N_3976,N_1227,N_1330);
xor U3977 (N_3977,N_2308,N_1324);
nor U3978 (N_3978,N_867,N_2134);
and U3979 (N_3979,N_920,N_244);
and U3980 (N_3980,N_982,N_1671);
nand U3981 (N_3981,N_1745,N_845);
nand U3982 (N_3982,N_1934,N_2329);
xnor U3983 (N_3983,N_1886,N_1989);
or U3984 (N_3984,N_916,N_1022);
or U3985 (N_3985,N_657,N_675);
xor U3986 (N_3986,N_9,N_1579);
xor U3987 (N_3987,N_285,N_1436);
xor U3988 (N_3988,N_353,N_314);
xor U3989 (N_3989,N_1426,N_3);
nor U3990 (N_3990,N_1182,N_2017);
or U3991 (N_3991,N_932,N_1503);
nor U3992 (N_3992,N_905,N_1908);
and U3993 (N_3993,N_113,N_1183);
or U3994 (N_3994,N_1205,N_1937);
xnor U3995 (N_3995,N_34,N_2355);
nand U3996 (N_3996,N_1366,N_2075);
or U3997 (N_3997,N_480,N_2310);
or U3998 (N_3998,N_1059,N_30);
nand U3999 (N_3999,N_113,N_1489);
and U4000 (N_4000,N_1951,N_180);
or U4001 (N_4001,N_2208,N_2495);
or U4002 (N_4002,N_859,N_1976);
nor U4003 (N_4003,N_2119,N_39);
nor U4004 (N_4004,N_266,N_1412);
nor U4005 (N_4005,N_1949,N_1303);
or U4006 (N_4006,N_1490,N_1177);
or U4007 (N_4007,N_454,N_767);
or U4008 (N_4008,N_1136,N_820);
xor U4009 (N_4009,N_2147,N_1716);
or U4010 (N_4010,N_1854,N_487);
and U4011 (N_4011,N_2447,N_2062);
and U4012 (N_4012,N_2199,N_342);
nand U4013 (N_4013,N_1126,N_214);
or U4014 (N_4014,N_1994,N_176);
nand U4015 (N_4015,N_943,N_1981);
nand U4016 (N_4016,N_375,N_2172);
nor U4017 (N_4017,N_717,N_1569);
nor U4018 (N_4018,N_2283,N_389);
nor U4019 (N_4019,N_2159,N_618);
or U4020 (N_4020,N_2170,N_2091);
or U4021 (N_4021,N_1765,N_991);
nand U4022 (N_4022,N_24,N_1551);
nor U4023 (N_4023,N_1425,N_1442);
or U4024 (N_4024,N_658,N_925);
or U4025 (N_4025,N_64,N_81);
and U4026 (N_4026,N_635,N_1352);
xor U4027 (N_4027,N_890,N_2265);
nand U4028 (N_4028,N_1320,N_1182);
nand U4029 (N_4029,N_2293,N_1202);
or U4030 (N_4030,N_1300,N_2392);
or U4031 (N_4031,N_2303,N_1760);
or U4032 (N_4032,N_1746,N_112);
xnor U4033 (N_4033,N_1868,N_1161);
nor U4034 (N_4034,N_163,N_391);
and U4035 (N_4035,N_1631,N_1820);
xor U4036 (N_4036,N_290,N_1372);
or U4037 (N_4037,N_2453,N_1798);
nand U4038 (N_4038,N_1022,N_1609);
xor U4039 (N_4039,N_2075,N_1414);
nand U4040 (N_4040,N_1260,N_2258);
nor U4041 (N_4041,N_2211,N_1070);
or U4042 (N_4042,N_1907,N_1263);
or U4043 (N_4043,N_1054,N_161);
and U4044 (N_4044,N_1520,N_836);
nor U4045 (N_4045,N_1060,N_132);
and U4046 (N_4046,N_160,N_1594);
and U4047 (N_4047,N_349,N_2216);
xnor U4048 (N_4048,N_595,N_97);
xor U4049 (N_4049,N_1232,N_1600);
nor U4050 (N_4050,N_1841,N_197);
nand U4051 (N_4051,N_19,N_2029);
nor U4052 (N_4052,N_475,N_2169);
xnor U4053 (N_4053,N_1667,N_822);
nand U4054 (N_4054,N_1286,N_413);
xnor U4055 (N_4055,N_135,N_920);
nand U4056 (N_4056,N_1241,N_1571);
nand U4057 (N_4057,N_617,N_2064);
nor U4058 (N_4058,N_1608,N_880);
xnor U4059 (N_4059,N_531,N_698);
or U4060 (N_4060,N_731,N_1335);
nand U4061 (N_4061,N_738,N_548);
xnor U4062 (N_4062,N_1080,N_2350);
or U4063 (N_4063,N_1713,N_1945);
xnor U4064 (N_4064,N_1553,N_1754);
nand U4065 (N_4065,N_1015,N_2243);
or U4066 (N_4066,N_649,N_891);
or U4067 (N_4067,N_200,N_1163);
and U4068 (N_4068,N_907,N_1871);
nand U4069 (N_4069,N_1265,N_2122);
xnor U4070 (N_4070,N_1565,N_1108);
or U4071 (N_4071,N_1111,N_125);
nor U4072 (N_4072,N_2304,N_600);
nand U4073 (N_4073,N_1565,N_1159);
and U4074 (N_4074,N_1242,N_1977);
or U4075 (N_4075,N_687,N_1764);
xnor U4076 (N_4076,N_839,N_2391);
and U4077 (N_4077,N_1830,N_1813);
xor U4078 (N_4078,N_1044,N_2318);
nor U4079 (N_4079,N_951,N_633);
nor U4080 (N_4080,N_1778,N_1730);
or U4081 (N_4081,N_814,N_1267);
nand U4082 (N_4082,N_1543,N_285);
xor U4083 (N_4083,N_1376,N_1065);
or U4084 (N_4084,N_753,N_711);
nand U4085 (N_4085,N_1782,N_2451);
xnor U4086 (N_4086,N_244,N_2038);
nor U4087 (N_4087,N_1982,N_2121);
or U4088 (N_4088,N_2233,N_941);
nand U4089 (N_4089,N_387,N_696);
and U4090 (N_4090,N_250,N_679);
nor U4091 (N_4091,N_764,N_2310);
nand U4092 (N_4092,N_1432,N_896);
and U4093 (N_4093,N_2051,N_87);
nor U4094 (N_4094,N_2175,N_1508);
or U4095 (N_4095,N_1999,N_2179);
or U4096 (N_4096,N_2214,N_472);
and U4097 (N_4097,N_2147,N_2137);
xor U4098 (N_4098,N_1187,N_380);
nand U4099 (N_4099,N_1591,N_1613);
nand U4100 (N_4100,N_2412,N_2243);
or U4101 (N_4101,N_878,N_564);
xor U4102 (N_4102,N_1411,N_76);
xnor U4103 (N_4103,N_1433,N_704);
nor U4104 (N_4104,N_1221,N_1157);
xor U4105 (N_4105,N_346,N_601);
or U4106 (N_4106,N_291,N_2194);
xor U4107 (N_4107,N_878,N_327);
and U4108 (N_4108,N_1960,N_2087);
and U4109 (N_4109,N_122,N_1995);
xor U4110 (N_4110,N_2134,N_571);
nor U4111 (N_4111,N_2222,N_1786);
xnor U4112 (N_4112,N_2059,N_352);
nor U4113 (N_4113,N_706,N_2256);
nand U4114 (N_4114,N_146,N_1098);
xnor U4115 (N_4115,N_1765,N_354);
and U4116 (N_4116,N_1239,N_1493);
or U4117 (N_4117,N_113,N_715);
nand U4118 (N_4118,N_465,N_38);
nand U4119 (N_4119,N_1811,N_2365);
xor U4120 (N_4120,N_964,N_71);
and U4121 (N_4121,N_2299,N_2140);
or U4122 (N_4122,N_669,N_504);
nor U4123 (N_4123,N_1804,N_967);
nor U4124 (N_4124,N_1059,N_692);
or U4125 (N_4125,N_42,N_2075);
nor U4126 (N_4126,N_285,N_2277);
or U4127 (N_4127,N_2306,N_1369);
nand U4128 (N_4128,N_291,N_2269);
nor U4129 (N_4129,N_1342,N_2384);
or U4130 (N_4130,N_2462,N_2219);
nor U4131 (N_4131,N_636,N_1580);
xnor U4132 (N_4132,N_796,N_1591);
nor U4133 (N_4133,N_434,N_1255);
or U4134 (N_4134,N_1490,N_38);
and U4135 (N_4135,N_629,N_2132);
and U4136 (N_4136,N_1673,N_1880);
and U4137 (N_4137,N_2228,N_82);
nor U4138 (N_4138,N_2282,N_2154);
xor U4139 (N_4139,N_1086,N_2135);
nor U4140 (N_4140,N_299,N_1784);
or U4141 (N_4141,N_105,N_2468);
nor U4142 (N_4142,N_1414,N_1690);
nor U4143 (N_4143,N_1644,N_2335);
nor U4144 (N_4144,N_1659,N_479);
nor U4145 (N_4145,N_867,N_695);
and U4146 (N_4146,N_370,N_1976);
xnor U4147 (N_4147,N_1601,N_1337);
xor U4148 (N_4148,N_1035,N_1290);
nand U4149 (N_4149,N_2394,N_2082);
xnor U4150 (N_4150,N_1567,N_1452);
and U4151 (N_4151,N_1215,N_2079);
xnor U4152 (N_4152,N_1557,N_1224);
nand U4153 (N_4153,N_2005,N_1374);
xor U4154 (N_4154,N_2468,N_990);
xor U4155 (N_4155,N_533,N_1451);
nand U4156 (N_4156,N_2099,N_1262);
nor U4157 (N_4157,N_912,N_340);
xnor U4158 (N_4158,N_752,N_1);
nor U4159 (N_4159,N_1263,N_572);
nand U4160 (N_4160,N_2295,N_2349);
nor U4161 (N_4161,N_1170,N_464);
nor U4162 (N_4162,N_253,N_2049);
nor U4163 (N_4163,N_927,N_1967);
or U4164 (N_4164,N_472,N_117);
xnor U4165 (N_4165,N_1231,N_245);
nor U4166 (N_4166,N_1964,N_199);
nand U4167 (N_4167,N_2472,N_49);
xnor U4168 (N_4168,N_482,N_1055);
and U4169 (N_4169,N_1249,N_2135);
nand U4170 (N_4170,N_796,N_1545);
nor U4171 (N_4171,N_1287,N_271);
and U4172 (N_4172,N_2434,N_1969);
xor U4173 (N_4173,N_182,N_241);
nand U4174 (N_4174,N_1851,N_1435);
and U4175 (N_4175,N_1384,N_1712);
xor U4176 (N_4176,N_1066,N_206);
and U4177 (N_4177,N_1649,N_2442);
or U4178 (N_4178,N_1035,N_2220);
nor U4179 (N_4179,N_1445,N_2148);
or U4180 (N_4180,N_2426,N_669);
nor U4181 (N_4181,N_571,N_338);
xnor U4182 (N_4182,N_985,N_2055);
and U4183 (N_4183,N_1358,N_343);
or U4184 (N_4184,N_1159,N_353);
nor U4185 (N_4185,N_1790,N_2435);
nand U4186 (N_4186,N_853,N_2401);
and U4187 (N_4187,N_1698,N_1838);
xor U4188 (N_4188,N_2474,N_1907);
or U4189 (N_4189,N_1593,N_1964);
or U4190 (N_4190,N_935,N_127);
nand U4191 (N_4191,N_2100,N_1203);
xnor U4192 (N_4192,N_240,N_1100);
nand U4193 (N_4193,N_1574,N_635);
nand U4194 (N_4194,N_2183,N_1990);
nor U4195 (N_4195,N_2476,N_273);
xor U4196 (N_4196,N_598,N_2476);
and U4197 (N_4197,N_2422,N_2095);
nand U4198 (N_4198,N_418,N_111);
xnor U4199 (N_4199,N_84,N_595);
nand U4200 (N_4200,N_2392,N_1689);
nor U4201 (N_4201,N_1266,N_767);
nor U4202 (N_4202,N_2336,N_1608);
nor U4203 (N_4203,N_1802,N_999);
xnor U4204 (N_4204,N_177,N_418);
and U4205 (N_4205,N_100,N_1166);
nand U4206 (N_4206,N_1770,N_1372);
and U4207 (N_4207,N_656,N_1002);
xnor U4208 (N_4208,N_2062,N_397);
xor U4209 (N_4209,N_1152,N_849);
and U4210 (N_4210,N_505,N_939);
xnor U4211 (N_4211,N_427,N_934);
nor U4212 (N_4212,N_2467,N_1813);
nor U4213 (N_4213,N_1313,N_1641);
xor U4214 (N_4214,N_2454,N_1748);
nand U4215 (N_4215,N_1849,N_2306);
nor U4216 (N_4216,N_1864,N_1030);
and U4217 (N_4217,N_387,N_919);
and U4218 (N_4218,N_16,N_2263);
nor U4219 (N_4219,N_1582,N_1503);
nand U4220 (N_4220,N_1364,N_2289);
nand U4221 (N_4221,N_70,N_1292);
and U4222 (N_4222,N_1168,N_691);
nand U4223 (N_4223,N_1965,N_1903);
nand U4224 (N_4224,N_934,N_1165);
and U4225 (N_4225,N_2164,N_985);
xnor U4226 (N_4226,N_308,N_1435);
nor U4227 (N_4227,N_1793,N_1017);
and U4228 (N_4228,N_1903,N_947);
nand U4229 (N_4229,N_1902,N_1732);
nor U4230 (N_4230,N_564,N_2425);
and U4231 (N_4231,N_2153,N_696);
and U4232 (N_4232,N_442,N_2033);
nor U4233 (N_4233,N_1139,N_2487);
and U4234 (N_4234,N_264,N_167);
or U4235 (N_4235,N_1512,N_217);
xnor U4236 (N_4236,N_660,N_995);
xnor U4237 (N_4237,N_2494,N_1349);
nand U4238 (N_4238,N_1962,N_538);
nor U4239 (N_4239,N_1696,N_568);
nand U4240 (N_4240,N_1988,N_1942);
and U4241 (N_4241,N_184,N_285);
nand U4242 (N_4242,N_1303,N_436);
xor U4243 (N_4243,N_989,N_404);
nor U4244 (N_4244,N_2041,N_286);
or U4245 (N_4245,N_2091,N_1075);
and U4246 (N_4246,N_2392,N_2368);
nand U4247 (N_4247,N_773,N_1928);
xor U4248 (N_4248,N_1107,N_1720);
nor U4249 (N_4249,N_2074,N_178);
and U4250 (N_4250,N_1711,N_2008);
and U4251 (N_4251,N_2168,N_297);
nand U4252 (N_4252,N_782,N_1606);
or U4253 (N_4253,N_527,N_2429);
nand U4254 (N_4254,N_1806,N_1558);
or U4255 (N_4255,N_2237,N_575);
and U4256 (N_4256,N_878,N_940);
or U4257 (N_4257,N_63,N_919);
nand U4258 (N_4258,N_2154,N_378);
or U4259 (N_4259,N_2179,N_2081);
nor U4260 (N_4260,N_972,N_484);
nor U4261 (N_4261,N_833,N_1940);
nor U4262 (N_4262,N_214,N_198);
nand U4263 (N_4263,N_1825,N_2329);
nor U4264 (N_4264,N_690,N_1535);
nand U4265 (N_4265,N_1573,N_1840);
xor U4266 (N_4266,N_2340,N_2346);
nor U4267 (N_4267,N_1051,N_1485);
nor U4268 (N_4268,N_1900,N_331);
nor U4269 (N_4269,N_1211,N_1715);
and U4270 (N_4270,N_1458,N_1942);
and U4271 (N_4271,N_1016,N_2362);
nor U4272 (N_4272,N_1809,N_1663);
xnor U4273 (N_4273,N_1472,N_2359);
nand U4274 (N_4274,N_944,N_249);
nand U4275 (N_4275,N_998,N_1002);
nand U4276 (N_4276,N_2106,N_556);
or U4277 (N_4277,N_2113,N_237);
nor U4278 (N_4278,N_383,N_105);
and U4279 (N_4279,N_2217,N_2440);
nor U4280 (N_4280,N_1076,N_923);
nand U4281 (N_4281,N_2143,N_1967);
or U4282 (N_4282,N_165,N_2297);
and U4283 (N_4283,N_730,N_726);
and U4284 (N_4284,N_1193,N_66);
or U4285 (N_4285,N_604,N_2039);
nand U4286 (N_4286,N_2298,N_335);
nand U4287 (N_4287,N_677,N_676);
or U4288 (N_4288,N_2273,N_1836);
nor U4289 (N_4289,N_875,N_1932);
or U4290 (N_4290,N_2154,N_111);
and U4291 (N_4291,N_419,N_69);
xnor U4292 (N_4292,N_1073,N_667);
nor U4293 (N_4293,N_1679,N_2298);
nor U4294 (N_4294,N_2029,N_805);
or U4295 (N_4295,N_2137,N_500);
nand U4296 (N_4296,N_2268,N_1247);
xnor U4297 (N_4297,N_829,N_1938);
nor U4298 (N_4298,N_37,N_501);
and U4299 (N_4299,N_45,N_1704);
xor U4300 (N_4300,N_328,N_1237);
xnor U4301 (N_4301,N_490,N_1739);
and U4302 (N_4302,N_839,N_608);
or U4303 (N_4303,N_558,N_1341);
or U4304 (N_4304,N_705,N_903);
xor U4305 (N_4305,N_1013,N_1770);
nor U4306 (N_4306,N_809,N_2263);
xnor U4307 (N_4307,N_1956,N_1024);
nor U4308 (N_4308,N_1316,N_1201);
xor U4309 (N_4309,N_2040,N_1623);
and U4310 (N_4310,N_1457,N_568);
nor U4311 (N_4311,N_2297,N_27);
and U4312 (N_4312,N_2159,N_62);
nor U4313 (N_4313,N_1886,N_60);
or U4314 (N_4314,N_2031,N_240);
nor U4315 (N_4315,N_225,N_882);
and U4316 (N_4316,N_2029,N_410);
nand U4317 (N_4317,N_2044,N_1916);
or U4318 (N_4318,N_1532,N_1623);
nand U4319 (N_4319,N_173,N_122);
nor U4320 (N_4320,N_1842,N_839);
and U4321 (N_4321,N_723,N_364);
nand U4322 (N_4322,N_264,N_358);
nor U4323 (N_4323,N_2344,N_1094);
nand U4324 (N_4324,N_2050,N_956);
nand U4325 (N_4325,N_2499,N_2132);
nor U4326 (N_4326,N_96,N_1463);
nand U4327 (N_4327,N_432,N_1211);
or U4328 (N_4328,N_716,N_149);
nor U4329 (N_4329,N_117,N_1805);
nand U4330 (N_4330,N_574,N_1383);
and U4331 (N_4331,N_241,N_248);
or U4332 (N_4332,N_2371,N_993);
and U4333 (N_4333,N_945,N_122);
xnor U4334 (N_4334,N_2477,N_1039);
nor U4335 (N_4335,N_2463,N_1408);
and U4336 (N_4336,N_2222,N_136);
nand U4337 (N_4337,N_624,N_1332);
xnor U4338 (N_4338,N_2455,N_2238);
nor U4339 (N_4339,N_564,N_80);
or U4340 (N_4340,N_765,N_1493);
nor U4341 (N_4341,N_73,N_2035);
nor U4342 (N_4342,N_313,N_785);
and U4343 (N_4343,N_1384,N_1414);
xor U4344 (N_4344,N_516,N_1540);
nand U4345 (N_4345,N_1311,N_1647);
and U4346 (N_4346,N_79,N_2142);
nand U4347 (N_4347,N_62,N_1072);
xnor U4348 (N_4348,N_698,N_1968);
or U4349 (N_4349,N_516,N_2336);
and U4350 (N_4350,N_1016,N_744);
xnor U4351 (N_4351,N_976,N_956);
xor U4352 (N_4352,N_285,N_1014);
and U4353 (N_4353,N_890,N_1401);
xor U4354 (N_4354,N_1041,N_1445);
and U4355 (N_4355,N_1931,N_823);
nand U4356 (N_4356,N_1724,N_1455);
nand U4357 (N_4357,N_586,N_516);
and U4358 (N_4358,N_2407,N_1836);
and U4359 (N_4359,N_1933,N_346);
and U4360 (N_4360,N_1718,N_734);
or U4361 (N_4361,N_764,N_144);
or U4362 (N_4362,N_814,N_1694);
nor U4363 (N_4363,N_1564,N_1288);
nand U4364 (N_4364,N_1812,N_2380);
or U4365 (N_4365,N_119,N_693);
and U4366 (N_4366,N_2133,N_2178);
or U4367 (N_4367,N_758,N_2267);
xor U4368 (N_4368,N_274,N_1402);
or U4369 (N_4369,N_1972,N_238);
or U4370 (N_4370,N_1168,N_357);
xor U4371 (N_4371,N_1716,N_1561);
nand U4372 (N_4372,N_1262,N_1081);
nor U4373 (N_4373,N_691,N_80);
or U4374 (N_4374,N_2219,N_595);
nand U4375 (N_4375,N_259,N_2078);
or U4376 (N_4376,N_893,N_2023);
nor U4377 (N_4377,N_1162,N_2435);
xor U4378 (N_4378,N_1850,N_987);
nor U4379 (N_4379,N_1909,N_1955);
nor U4380 (N_4380,N_1109,N_1848);
and U4381 (N_4381,N_2325,N_2324);
and U4382 (N_4382,N_858,N_1503);
or U4383 (N_4383,N_2194,N_2341);
or U4384 (N_4384,N_2003,N_27);
and U4385 (N_4385,N_1461,N_1859);
nor U4386 (N_4386,N_88,N_1408);
nand U4387 (N_4387,N_1547,N_511);
or U4388 (N_4388,N_1970,N_1907);
nor U4389 (N_4389,N_1155,N_1203);
nor U4390 (N_4390,N_1712,N_1416);
or U4391 (N_4391,N_765,N_2083);
nand U4392 (N_4392,N_865,N_236);
or U4393 (N_4393,N_2286,N_2431);
xor U4394 (N_4394,N_463,N_2347);
or U4395 (N_4395,N_1206,N_489);
and U4396 (N_4396,N_1113,N_853);
or U4397 (N_4397,N_2162,N_1317);
and U4398 (N_4398,N_777,N_939);
nor U4399 (N_4399,N_2405,N_1426);
xor U4400 (N_4400,N_1797,N_1471);
or U4401 (N_4401,N_898,N_514);
and U4402 (N_4402,N_971,N_279);
or U4403 (N_4403,N_916,N_1300);
nor U4404 (N_4404,N_1796,N_1933);
or U4405 (N_4405,N_55,N_65);
or U4406 (N_4406,N_337,N_1349);
nor U4407 (N_4407,N_1304,N_1711);
or U4408 (N_4408,N_2345,N_887);
xnor U4409 (N_4409,N_477,N_2176);
xnor U4410 (N_4410,N_2089,N_1715);
xnor U4411 (N_4411,N_2231,N_2449);
and U4412 (N_4412,N_402,N_134);
nand U4413 (N_4413,N_1540,N_2491);
and U4414 (N_4414,N_131,N_140);
or U4415 (N_4415,N_2115,N_2233);
nand U4416 (N_4416,N_234,N_1021);
xor U4417 (N_4417,N_1177,N_30);
and U4418 (N_4418,N_2177,N_1671);
nor U4419 (N_4419,N_1025,N_1121);
nand U4420 (N_4420,N_1892,N_1475);
and U4421 (N_4421,N_160,N_120);
xnor U4422 (N_4422,N_1854,N_1189);
nand U4423 (N_4423,N_2388,N_2472);
and U4424 (N_4424,N_1480,N_1442);
nand U4425 (N_4425,N_824,N_1847);
nor U4426 (N_4426,N_1015,N_1171);
nand U4427 (N_4427,N_562,N_359);
nor U4428 (N_4428,N_2248,N_1072);
nand U4429 (N_4429,N_1075,N_448);
or U4430 (N_4430,N_266,N_1662);
and U4431 (N_4431,N_1026,N_266);
xor U4432 (N_4432,N_147,N_57);
nor U4433 (N_4433,N_2404,N_1023);
nand U4434 (N_4434,N_332,N_60);
nor U4435 (N_4435,N_859,N_2131);
or U4436 (N_4436,N_1374,N_2119);
or U4437 (N_4437,N_4,N_486);
nor U4438 (N_4438,N_2034,N_1810);
xnor U4439 (N_4439,N_122,N_56);
xor U4440 (N_4440,N_1922,N_357);
and U4441 (N_4441,N_806,N_198);
nand U4442 (N_4442,N_2041,N_718);
nand U4443 (N_4443,N_1673,N_1805);
nand U4444 (N_4444,N_884,N_1945);
xor U4445 (N_4445,N_1621,N_1417);
nand U4446 (N_4446,N_220,N_1827);
or U4447 (N_4447,N_818,N_1790);
nor U4448 (N_4448,N_2117,N_2131);
or U4449 (N_4449,N_2148,N_1580);
nor U4450 (N_4450,N_2405,N_773);
nor U4451 (N_4451,N_637,N_1382);
and U4452 (N_4452,N_2361,N_1413);
nand U4453 (N_4453,N_1839,N_1588);
nor U4454 (N_4454,N_2443,N_2325);
nand U4455 (N_4455,N_1206,N_745);
and U4456 (N_4456,N_1951,N_1250);
xnor U4457 (N_4457,N_244,N_761);
or U4458 (N_4458,N_1342,N_1388);
and U4459 (N_4459,N_2424,N_2058);
nor U4460 (N_4460,N_588,N_1045);
nand U4461 (N_4461,N_1712,N_966);
or U4462 (N_4462,N_2264,N_655);
nor U4463 (N_4463,N_1367,N_269);
nor U4464 (N_4464,N_2366,N_685);
nand U4465 (N_4465,N_160,N_623);
xnor U4466 (N_4466,N_1114,N_1652);
and U4467 (N_4467,N_1486,N_1167);
and U4468 (N_4468,N_1049,N_887);
nor U4469 (N_4469,N_41,N_877);
and U4470 (N_4470,N_350,N_2221);
nor U4471 (N_4471,N_697,N_287);
nor U4472 (N_4472,N_874,N_1907);
and U4473 (N_4473,N_2464,N_280);
xnor U4474 (N_4474,N_387,N_160);
xor U4475 (N_4475,N_1898,N_1963);
and U4476 (N_4476,N_612,N_1352);
nand U4477 (N_4477,N_150,N_1783);
nand U4478 (N_4478,N_1688,N_2201);
xnor U4479 (N_4479,N_192,N_135);
nor U4480 (N_4480,N_418,N_811);
or U4481 (N_4481,N_99,N_833);
and U4482 (N_4482,N_1958,N_2199);
nor U4483 (N_4483,N_2315,N_935);
or U4484 (N_4484,N_1756,N_746);
xor U4485 (N_4485,N_2146,N_1862);
nand U4486 (N_4486,N_2218,N_2443);
and U4487 (N_4487,N_2172,N_2499);
xor U4488 (N_4488,N_1334,N_28);
xor U4489 (N_4489,N_1652,N_2140);
nor U4490 (N_4490,N_2486,N_449);
nand U4491 (N_4491,N_2260,N_572);
nor U4492 (N_4492,N_97,N_732);
or U4493 (N_4493,N_1139,N_1727);
xnor U4494 (N_4494,N_1234,N_2004);
and U4495 (N_4495,N_1038,N_40);
nand U4496 (N_4496,N_975,N_700);
and U4497 (N_4497,N_972,N_39);
xnor U4498 (N_4498,N_1233,N_1644);
xnor U4499 (N_4499,N_2136,N_1529);
nor U4500 (N_4500,N_272,N_30);
nand U4501 (N_4501,N_617,N_2488);
xnor U4502 (N_4502,N_465,N_2044);
xor U4503 (N_4503,N_2483,N_485);
or U4504 (N_4504,N_295,N_1500);
or U4505 (N_4505,N_510,N_166);
nand U4506 (N_4506,N_215,N_736);
nor U4507 (N_4507,N_1273,N_432);
and U4508 (N_4508,N_51,N_67);
nand U4509 (N_4509,N_2278,N_98);
or U4510 (N_4510,N_1134,N_1294);
nand U4511 (N_4511,N_930,N_474);
nand U4512 (N_4512,N_1780,N_175);
nand U4513 (N_4513,N_487,N_1945);
nor U4514 (N_4514,N_886,N_876);
and U4515 (N_4515,N_2111,N_1586);
xor U4516 (N_4516,N_871,N_2140);
and U4517 (N_4517,N_806,N_1496);
or U4518 (N_4518,N_1656,N_2029);
xor U4519 (N_4519,N_2282,N_2066);
nand U4520 (N_4520,N_129,N_1156);
xor U4521 (N_4521,N_1534,N_2387);
xnor U4522 (N_4522,N_2071,N_2349);
nand U4523 (N_4523,N_2293,N_294);
nand U4524 (N_4524,N_2425,N_2185);
nor U4525 (N_4525,N_85,N_1993);
nor U4526 (N_4526,N_1124,N_461);
nand U4527 (N_4527,N_2333,N_2317);
or U4528 (N_4528,N_2480,N_960);
and U4529 (N_4529,N_1389,N_1289);
xor U4530 (N_4530,N_633,N_467);
nor U4531 (N_4531,N_592,N_2090);
nand U4532 (N_4532,N_1868,N_2367);
nand U4533 (N_4533,N_1282,N_2304);
nand U4534 (N_4534,N_1467,N_728);
and U4535 (N_4535,N_24,N_2408);
nand U4536 (N_4536,N_1224,N_783);
xor U4537 (N_4537,N_2016,N_389);
xnor U4538 (N_4538,N_82,N_1107);
or U4539 (N_4539,N_242,N_2298);
nor U4540 (N_4540,N_2318,N_1364);
or U4541 (N_4541,N_1793,N_1270);
or U4542 (N_4542,N_1756,N_1133);
nand U4543 (N_4543,N_119,N_1135);
xnor U4544 (N_4544,N_2298,N_2006);
nor U4545 (N_4545,N_1311,N_2439);
xnor U4546 (N_4546,N_315,N_156);
nand U4547 (N_4547,N_1131,N_461);
and U4548 (N_4548,N_741,N_47);
nor U4549 (N_4549,N_491,N_2464);
nand U4550 (N_4550,N_2081,N_1153);
nand U4551 (N_4551,N_689,N_260);
xnor U4552 (N_4552,N_2111,N_2413);
and U4553 (N_4553,N_2097,N_2396);
and U4554 (N_4554,N_1526,N_2000);
xor U4555 (N_4555,N_1985,N_1376);
or U4556 (N_4556,N_119,N_115);
and U4557 (N_4557,N_1006,N_2002);
xor U4558 (N_4558,N_1420,N_1477);
nor U4559 (N_4559,N_1051,N_630);
and U4560 (N_4560,N_1628,N_463);
nand U4561 (N_4561,N_734,N_575);
and U4562 (N_4562,N_287,N_1620);
and U4563 (N_4563,N_1601,N_1974);
or U4564 (N_4564,N_1238,N_1682);
and U4565 (N_4565,N_733,N_35);
and U4566 (N_4566,N_588,N_2029);
and U4567 (N_4567,N_543,N_696);
xor U4568 (N_4568,N_692,N_12);
xnor U4569 (N_4569,N_490,N_2203);
nor U4570 (N_4570,N_747,N_1815);
nor U4571 (N_4571,N_1954,N_2450);
or U4572 (N_4572,N_2157,N_2417);
nand U4573 (N_4573,N_1397,N_167);
nand U4574 (N_4574,N_2104,N_1743);
xnor U4575 (N_4575,N_1775,N_1857);
or U4576 (N_4576,N_1349,N_2225);
xnor U4577 (N_4577,N_2387,N_1734);
xor U4578 (N_4578,N_59,N_522);
or U4579 (N_4579,N_2252,N_989);
or U4580 (N_4580,N_2170,N_2445);
nand U4581 (N_4581,N_18,N_1896);
or U4582 (N_4582,N_1614,N_14);
nor U4583 (N_4583,N_1697,N_1263);
nor U4584 (N_4584,N_2028,N_543);
or U4585 (N_4585,N_0,N_644);
or U4586 (N_4586,N_2484,N_2455);
or U4587 (N_4587,N_874,N_972);
nand U4588 (N_4588,N_1812,N_2269);
nor U4589 (N_4589,N_1737,N_607);
nor U4590 (N_4590,N_2216,N_28);
nor U4591 (N_4591,N_1963,N_762);
xor U4592 (N_4592,N_2306,N_711);
or U4593 (N_4593,N_463,N_1600);
and U4594 (N_4594,N_1875,N_1814);
nand U4595 (N_4595,N_2009,N_1848);
nand U4596 (N_4596,N_2267,N_881);
xnor U4597 (N_4597,N_847,N_1974);
and U4598 (N_4598,N_389,N_224);
nand U4599 (N_4599,N_2105,N_1025);
and U4600 (N_4600,N_183,N_1588);
or U4601 (N_4601,N_1690,N_2171);
or U4602 (N_4602,N_1667,N_1270);
nor U4603 (N_4603,N_1881,N_1263);
xor U4604 (N_4604,N_851,N_1952);
and U4605 (N_4605,N_2426,N_994);
and U4606 (N_4606,N_1556,N_1366);
or U4607 (N_4607,N_88,N_1168);
xnor U4608 (N_4608,N_2309,N_1148);
or U4609 (N_4609,N_306,N_1738);
or U4610 (N_4610,N_859,N_217);
or U4611 (N_4611,N_617,N_70);
xor U4612 (N_4612,N_718,N_157);
nor U4613 (N_4613,N_1392,N_759);
nand U4614 (N_4614,N_1264,N_1818);
nor U4615 (N_4615,N_475,N_2114);
xnor U4616 (N_4616,N_1701,N_1679);
xnor U4617 (N_4617,N_1480,N_2032);
and U4618 (N_4618,N_790,N_1108);
or U4619 (N_4619,N_2497,N_1287);
or U4620 (N_4620,N_1510,N_1155);
and U4621 (N_4621,N_2449,N_1654);
xnor U4622 (N_4622,N_1734,N_250);
nand U4623 (N_4623,N_1788,N_521);
and U4624 (N_4624,N_531,N_1809);
nand U4625 (N_4625,N_1491,N_1567);
xnor U4626 (N_4626,N_832,N_657);
or U4627 (N_4627,N_1000,N_1688);
xnor U4628 (N_4628,N_701,N_2401);
xnor U4629 (N_4629,N_66,N_2453);
xnor U4630 (N_4630,N_1554,N_1872);
xnor U4631 (N_4631,N_37,N_2029);
xnor U4632 (N_4632,N_674,N_789);
and U4633 (N_4633,N_2317,N_897);
nand U4634 (N_4634,N_2404,N_1789);
xnor U4635 (N_4635,N_1162,N_1279);
nor U4636 (N_4636,N_1389,N_1036);
xor U4637 (N_4637,N_1671,N_1892);
or U4638 (N_4638,N_383,N_519);
nor U4639 (N_4639,N_469,N_804);
or U4640 (N_4640,N_1560,N_669);
nor U4641 (N_4641,N_588,N_1297);
nor U4642 (N_4642,N_1034,N_2300);
or U4643 (N_4643,N_2056,N_2346);
and U4644 (N_4644,N_50,N_858);
or U4645 (N_4645,N_12,N_1062);
nor U4646 (N_4646,N_885,N_671);
or U4647 (N_4647,N_2437,N_2447);
nand U4648 (N_4648,N_42,N_1177);
nand U4649 (N_4649,N_2014,N_1192);
nor U4650 (N_4650,N_1803,N_778);
nand U4651 (N_4651,N_1063,N_1515);
nor U4652 (N_4652,N_2103,N_606);
nor U4653 (N_4653,N_143,N_1239);
xnor U4654 (N_4654,N_242,N_344);
or U4655 (N_4655,N_1361,N_1202);
and U4656 (N_4656,N_2332,N_314);
or U4657 (N_4657,N_1450,N_603);
nand U4658 (N_4658,N_2050,N_882);
or U4659 (N_4659,N_660,N_933);
nand U4660 (N_4660,N_548,N_1047);
nand U4661 (N_4661,N_366,N_632);
xor U4662 (N_4662,N_2221,N_1218);
xor U4663 (N_4663,N_330,N_1363);
and U4664 (N_4664,N_1825,N_1465);
nor U4665 (N_4665,N_506,N_201);
and U4666 (N_4666,N_1005,N_8);
and U4667 (N_4667,N_2248,N_1800);
or U4668 (N_4668,N_581,N_941);
nand U4669 (N_4669,N_1161,N_924);
xor U4670 (N_4670,N_1192,N_2093);
or U4671 (N_4671,N_1900,N_1248);
nand U4672 (N_4672,N_488,N_2100);
or U4673 (N_4673,N_1620,N_1377);
and U4674 (N_4674,N_1164,N_541);
or U4675 (N_4675,N_2474,N_2089);
nand U4676 (N_4676,N_1638,N_1410);
nor U4677 (N_4677,N_639,N_1394);
nand U4678 (N_4678,N_62,N_2134);
or U4679 (N_4679,N_1951,N_800);
xor U4680 (N_4680,N_1626,N_2480);
xor U4681 (N_4681,N_1664,N_1912);
or U4682 (N_4682,N_2471,N_463);
or U4683 (N_4683,N_2469,N_1321);
or U4684 (N_4684,N_605,N_2376);
and U4685 (N_4685,N_1019,N_1895);
and U4686 (N_4686,N_2260,N_1990);
or U4687 (N_4687,N_2225,N_2264);
nand U4688 (N_4688,N_185,N_256);
nand U4689 (N_4689,N_1185,N_369);
nand U4690 (N_4690,N_2465,N_801);
xnor U4691 (N_4691,N_2010,N_161);
or U4692 (N_4692,N_161,N_2194);
xnor U4693 (N_4693,N_2270,N_2192);
and U4694 (N_4694,N_543,N_622);
and U4695 (N_4695,N_567,N_1490);
xnor U4696 (N_4696,N_890,N_1805);
or U4697 (N_4697,N_937,N_82);
nor U4698 (N_4698,N_234,N_675);
or U4699 (N_4699,N_658,N_1708);
xnor U4700 (N_4700,N_1724,N_1980);
and U4701 (N_4701,N_603,N_943);
nand U4702 (N_4702,N_225,N_100);
nor U4703 (N_4703,N_2355,N_1788);
and U4704 (N_4704,N_323,N_2447);
or U4705 (N_4705,N_2417,N_2115);
and U4706 (N_4706,N_343,N_164);
nand U4707 (N_4707,N_1675,N_803);
nand U4708 (N_4708,N_1337,N_316);
nand U4709 (N_4709,N_1303,N_178);
nand U4710 (N_4710,N_1804,N_2040);
xnor U4711 (N_4711,N_2392,N_839);
nand U4712 (N_4712,N_827,N_477);
and U4713 (N_4713,N_1347,N_1935);
nand U4714 (N_4714,N_1700,N_305);
nand U4715 (N_4715,N_602,N_1629);
or U4716 (N_4716,N_2323,N_1254);
or U4717 (N_4717,N_1058,N_507);
and U4718 (N_4718,N_2196,N_31);
or U4719 (N_4719,N_2096,N_1208);
or U4720 (N_4720,N_301,N_394);
nand U4721 (N_4721,N_1967,N_832);
xor U4722 (N_4722,N_1410,N_1122);
xnor U4723 (N_4723,N_1502,N_1942);
or U4724 (N_4724,N_529,N_319);
nor U4725 (N_4725,N_1708,N_430);
and U4726 (N_4726,N_1769,N_676);
nor U4727 (N_4727,N_2256,N_833);
nand U4728 (N_4728,N_1802,N_106);
and U4729 (N_4729,N_460,N_1539);
or U4730 (N_4730,N_1747,N_315);
or U4731 (N_4731,N_754,N_1201);
xor U4732 (N_4732,N_1625,N_193);
xnor U4733 (N_4733,N_375,N_1961);
or U4734 (N_4734,N_1758,N_139);
xor U4735 (N_4735,N_1830,N_2003);
or U4736 (N_4736,N_567,N_395);
and U4737 (N_4737,N_107,N_65);
nand U4738 (N_4738,N_32,N_1741);
nand U4739 (N_4739,N_234,N_1478);
and U4740 (N_4740,N_506,N_1680);
nor U4741 (N_4741,N_1857,N_1048);
xnor U4742 (N_4742,N_2208,N_2079);
nor U4743 (N_4743,N_1851,N_2024);
or U4744 (N_4744,N_2170,N_1836);
and U4745 (N_4745,N_153,N_1469);
nor U4746 (N_4746,N_1835,N_44);
nand U4747 (N_4747,N_1179,N_422);
nor U4748 (N_4748,N_898,N_1364);
nor U4749 (N_4749,N_2291,N_73);
or U4750 (N_4750,N_545,N_1697);
xnor U4751 (N_4751,N_605,N_945);
xnor U4752 (N_4752,N_1572,N_479);
nand U4753 (N_4753,N_1035,N_2071);
or U4754 (N_4754,N_879,N_2163);
xnor U4755 (N_4755,N_2221,N_2417);
nand U4756 (N_4756,N_1722,N_48);
nor U4757 (N_4757,N_1016,N_1995);
nand U4758 (N_4758,N_2404,N_2230);
xnor U4759 (N_4759,N_2313,N_661);
nand U4760 (N_4760,N_1022,N_1925);
or U4761 (N_4761,N_1376,N_1522);
and U4762 (N_4762,N_2033,N_790);
xor U4763 (N_4763,N_1723,N_2413);
and U4764 (N_4764,N_2278,N_1194);
xor U4765 (N_4765,N_1192,N_2007);
or U4766 (N_4766,N_1599,N_2491);
and U4767 (N_4767,N_637,N_1626);
nand U4768 (N_4768,N_2087,N_283);
xnor U4769 (N_4769,N_165,N_1341);
nand U4770 (N_4770,N_2041,N_2427);
nor U4771 (N_4771,N_105,N_320);
nand U4772 (N_4772,N_1579,N_902);
and U4773 (N_4773,N_1701,N_1849);
or U4774 (N_4774,N_1613,N_2147);
and U4775 (N_4775,N_842,N_1080);
xnor U4776 (N_4776,N_960,N_1674);
and U4777 (N_4777,N_2216,N_1529);
and U4778 (N_4778,N_1059,N_1593);
or U4779 (N_4779,N_1469,N_1480);
nor U4780 (N_4780,N_869,N_2021);
and U4781 (N_4781,N_1793,N_394);
xnor U4782 (N_4782,N_368,N_2266);
or U4783 (N_4783,N_953,N_2439);
or U4784 (N_4784,N_536,N_1018);
or U4785 (N_4785,N_469,N_67);
nand U4786 (N_4786,N_2127,N_1862);
and U4787 (N_4787,N_23,N_2471);
nand U4788 (N_4788,N_2332,N_663);
and U4789 (N_4789,N_1403,N_2117);
and U4790 (N_4790,N_729,N_2361);
and U4791 (N_4791,N_2187,N_2381);
nand U4792 (N_4792,N_2060,N_1934);
xor U4793 (N_4793,N_2182,N_799);
xnor U4794 (N_4794,N_105,N_2115);
and U4795 (N_4795,N_1924,N_1810);
and U4796 (N_4796,N_1446,N_1475);
xor U4797 (N_4797,N_1507,N_35);
and U4798 (N_4798,N_509,N_1617);
xnor U4799 (N_4799,N_1104,N_1179);
nand U4800 (N_4800,N_2455,N_1723);
xnor U4801 (N_4801,N_726,N_1660);
xor U4802 (N_4802,N_2280,N_1836);
nand U4803 (N_4803,N_341,N_2323);
or U4804 (N_4804,N_1218,N_216);
nand U4805 (N_4805,N_865,N_2098);
xnor U4806 (N_4806,N_2320,N_1419);
or U4807 (N_4807,N_2139,N_1805);
nand U4808 (N_4808,N_386,N_592);
or U4809 (N_4809,N_2360,N_2363);
or U4810 (N_4810,N_116,N_2220);
or U4811 (N_4811,N_602,N_1636);
xnor U4812 (N_4812,N_41,N_472);
nor U4813 (N_4813,N_882,N_2349);
nor U4814 (N_4814,N_1277,N_1991);
nor U4815 (N_4815,N_2238,N_2185);
xor U4816 (N_4816,N_1230,N_1436);
and U4817 (N_4817,N_1874,N_677);
and U4818 (N_4818,N_1722,N_832);
nor U4819 (N_4819,N_643,N_2115);
xor U4820 (N_4820,N_1567,N_1402);
and U4821 (N_4821,N_37,N_1614);
nor U4822 (N_4822,N_1381,N_1415);
xnor U4823 (N_4823,N_222,N_1566);
nor U4824 (N_4824,N_29,N_1395);
and U4825 (N_4825,N_570,N_1446);
xor U4826 (N_4826,N_2487,N_2308);
nand U4827 (N_4827,N_953,N_1723);
or U4828 (N_4828,N_1720,N_2182);
or U4829 (N_4829,N_413,N_1627);
and U4830 (N_4830,N_1024,N_1623);
xnor U4831 (N_4831,N_1480,N_2047);
xnor U4832 (N_4832,N_1716,N_998);
or U4833 (N_4833,N_2042,N_522);
nor U4834 (N_4834,N_1676,N_844);
nor U4835 (N_4835,N_480,N_2207);
xor U4836 (N_4836,N_1521,N_790);
nor U4837 (N_4837,N_926,N_2081);
nand U4838 (N_4838,N_512,N_1341);
nor U4839 (N_4839,N_2403,N_2218);
and U4840 (N_4840,N_2282,N_1924);
nand U4841 (N_4841,N_1995,N_1209);
or U4842 (N_4842,N_1157,N_1237);
or U4843 (N_4843,N_1379,N_1853);
xor U4844 (N_4844,N_1119,N_348);
and U4845 (N_4845,N_429,N_1824);
nor U4846 (N_4846,N_506,N_2182);
and U4847 (N_4847,N_842,N_417);
and U4848 (N_4848,N_372,N_385);
nand U4849 (N_4849,N_1070,N_165);
xnor U4850 (N_4850,N_504,N_849);
and U4851 (N_4851,N_2160,N_280);
or U4852 (N_4852,N_1877,N_1657);
xor U4853 (N_4853,N_1094,N_2279);
nand U4854 (N_4854,N_903,N_948);
and U4855 (N_4855,N_1921,N_2374);
or U4856 (N_4856,N_2353,N_635);
and U4857 (N_4857,N_1170,N_2436);
or U4858 (N_4858,N_800,N_1999);
xor U4859 (N_4859,N_240,N_658);
nor U4860 (N_4860,N_369,N_1824);
or U4861 (N_4861,N_2235,N_1802);
nand U4862 (N_4862,N_1148,N_1439);
and U4863 (N_4863,N_431,N_1331);
xor U4864 (N_4864,N_730,N_1888);
nor U4865 (N_4865,N_906,N_2294);
and U4866 (N_4866,N_2165,N_1233);
and U4867 (N_4867,N_1166,N_2023);
nor U4868 (N_4868,N_274,N_1701);
and U4869 (N_4869,N_659,N_1470);
nand U4870 (N_4870,N_1707,N_443);
nand U4871 (N_4871,N_733,N_195);
nor U4872 (N_4872,N_665,N_1593);
nor U4873 (N_4873,N_370,N_781);
nand U4874 (N_4874,N_646,N_1623);
or U4875 (N_4875,N_2416,N_2048);
and U4876 (N_4876,N_1372,N_1910);
and U4877 (N_4877,N_1113,N_674);
or U4878 (N_4878,N_435,N_880);
and U4879 (N_4879,N_1906,N_2341);
or U4880 (N_4880,N_915,N_352);
nand U4881 (N_4881,N_2155,N_516);
and U4882 (N_4882,N_429,N_2157);
nor U4883 (N_4883,N_257,N_553);
and U4884 (N_4884,N_533,N_1591);
nor U4885 (N_4885,N_91,N_678);
and U4886 (N_4886,N_2369,N_2154);
nor U4887 (N_4887,N_2078,N_2410);
nor U4888 (N_4888,N_2302,N_1986);
nand U4889 (N_4889,N_1938,N_941);
or U4890 (N_4890,N_590,N_1623);
xnor U4891 (N_4891,N_1496,N_1704);
xor U4892 (N_4892,N_703,N_1119);
nand U4893 (N_4893,N_2031,N_1180);
or U4894 (N_4894,N_2200,N_2083);
xnor U4895 (N_4895,N_1193,N_2014);
nand U4896 (N_4896,N_16,N_2030);
nor U4897 (N_4897,N_2160,N_387);
xnor U4898 (N_4898,N_1110,N_891);
or U4899 (N_4899,N_2094,N_1916);
or U4900 (N_4900,N_1641,N_427);
nor U4901 (N_4901,N_2455,N_2423);
nor U4902 (N_4902,N_2425,N_1660);
and U4903 (N_4903,N_1035,N_2133);
nor U4904 (N_4904,N_829,N_1516);
nor U4905 (N_4905,N_906,N_2322);
nand U4906 (N_4906,N_157,N_1260);
or U4907 (N_4907,N_59,N_1145);
and U4908 (N_4908,N_2288,N_1484);
xnor U4909 (N_4909,N_47,N_2003);
xor U4910 (N_4910,N_1288,N_1380);
and U4911 (N_4911,N_287,N_171);
nor U4912 (N_4912,N_337,N_451);
nand U4913 (N_4913,N_1709,N_362);
or U4914 (N_4914,N_1510,N_2148);
nand U4915 (N_4915,N_1770,N_1854);
and U4916 (N_4916,N_2442,N_2116);
nand U4917 (N_4917,N_1304,N_1203);
and U4918 (N_4918,N_2163,N_1154);
nand U4919 (N_4919,N_929,N_1444);
xnor U4920 (N_4920,N_987,N_1444);
and U4921 (N_4921,N_1852,N_1061);
or U4922 (N_4922,N_2039,N_1711);
and U4923 (N_4923,N_1611,N_1);
or U4924 (N_4924,N_507,N_469);
and U4925 (N_4925,N_841,N_575);
nand U4926 (N_4926,N_994,N_922);
nand U4927 (N_4927,N_2197,N_903);
or U4928 (N_4928,N_414,N_2015);
and U4929 (N_4929,N_783,N_2452);
xnor U4930 (N_4930,N_282,N_2138);
xnor U4931 (N_4931,N_1770,N_1986);
and U4932 (N_4932,N_1034,N_913);
xor U4933 (N_4933,N_94,N_1782);
and U4934 (N_4934,N_2108,N_1623);
nor U4935 (N_4935,N_2381,N_2000);
or U4936 (N_4936,N_1613,N_2159);
or U4937 (N_4937,N_559,N_2362);
nand U4938 (N_4938,N_1593,N_1748);
xnor U4939 (N_4939,N_2436,N_2155);
xnor U4940 (N_4940,N_1422,N_2491);
or U4941 (N_4941,N_2460,N_357);
and U4942 (N_4942,N_1437,N_629);
and U4943 (N_4943,N_562,N_267);
and U4944 (N_4944,N_1614,N_2427);
nand U4945 (N_4945,N_2089,N_947);
and U4946 (N_4946,N_1232,N_1340);
xor U4947 (N_4947,N_1184,N_2194);
xor U4948 (N_4948,N_2074,N_1002);
and U4949 (N_4949,N_561,N_2364);
xnor U4950 (N_4950,N_1975,N_1247);
nor U4951 (N_4951,N_2201,N_1694);
nand U4952 (N_4952,N_293,N_424);
nand U4953 (N_4953,N_2023,N_2265);
and U4954 (N_4954,N_929,N_110);
nand U4955 (N_4955,N_1249,N_1021);
xor U4956 (N_4956,N_1315,N_380);
or U4957 (N_4957,N_1154,N_2238);
xnor U4958 (N_4958,N_248,N_1672);
nand U4959 (N_4959,N_231,N_498);
or U4960 (N_4960,N_1294,N_2434);
nor U4961 (N_4961,N_905,N_146);
or U4962 (N_4962,N_2299,N_1172);
nand U4963 (N_4963,N_1990,N_2293);
nor U4964 (N_4964,N_287,N_2288);
nor U4965 (N_4965,N_1909,N_1675);
nor U4966 (N_4966,N_1513,N_731);
nor U4967 (N_4967,N_633,N_338);
and U4968 (N_4968,N_1359,N_436);
or U4969 (N_4969,N_479,N_1411);
or U4970 (N_4970,N_638,N_1109);
xnor U4971 (N_4971,N_456,N_753);
nor U4972 (N_4972,N_1063,N_1510);
and U4973 (N_4973,N_421,N_2115);
nand U4974 (N_4974,N_2320,N_1370);
or U4975 (N_4975,N_388,N_1188);
and U4976 (N_4976,N_625,N_770);
xnor U4977 (N_4977,N_270,N_584);
nor U4978 (N_4978,N_1054,N_1651);
nand U4979 (N_4979,N_714,N_155);
and U4980 (N_4980,N_1334,N_271);
nand U4981 (N_4981,N_1654,N_2353);
xnor U4982 (N_4982,N_1089,N_1766);
or U4983 (N_4983,N_1531,N_394);
nand U4984 (N_4984,N_2429,N_1814);
and U4985 (N_4985,N_441,N_1635);
and U4986 (N_4986,N_2475,N_1282);
and U4987 (N_4987,N_1744,N_424);
and U4988 (N_4988,N_219,N_1191);
nor U4989 (N_4989,N_714,N_1134);
nor U4990 (N_4990,N_2496,N_850);
or U4991 (N_4991,N_501,N_1396);
xnor U4992 (N_4992,N_1697,N_878);
or U4993 (N_4993,N_558,N_1668);
nor U4994 (N_4994,N_1140,N_1466);
or U4995 (N_4995,N_969,N_1163);
xor U4996 (N_4996,N_982,N_2458);
nor U4997 (N_4997,N_2082,N_2179);
xnor U4998 (N_4998,N_1943,N_832);
nor U4999 (N_4999,N_1525,N_404);
and UO_0 (O_0,N_4734,N_4419);
nand UO_1 (O_1,N_3729,N_3832);
nor UO_2 (O_2,N_3253,N_3170);
nor UO_3 (O_3,N_4870,N_3895);
nand UO_4 (O_4,N_3865,N_4434);
xnor UO_5 (O_5,N_2834,N_3877);
nand UO_6 (O_6,N_3672,N_2892);
nand UO_7 (O_7,N_3748,N_4441);
or UO_8 (O_8,N_4582,N_2923);
and UO_9 (O_9,N_3187,N_2952);
nand UO_10 (O_10,N_3903,N_4209);
xor UO_11 (O_11,N_3595,N_4546);
or UO_12 (O_12,N_2701,N_3193);
or UO_13 (O_13,N_2725,N_3511);
nand UO_14 (O_14,N_3791,N_3608);
or UO_15 (O_15,N_4391,N_2802);
or UO_16 (O_16,N_4423,N_3210);
nor UO_17 (O_17,N_2819,N_4886);
or UO_18 (O_18,N_2635,N_2875);
nor UO_19 (O_19,N_3718,N_4207);
nor UO_20 (O_20,N_4347,N_3922);
xor UO_21 (O_21,N_2512,N_2651);
and UO_22 (O_22,N_2742,N_3157);
xor UO_23 (O_23,N_3821,N_4666);
xor UO_24 (O_24,N_3633,N_3703);
xnor UO_25 (O_25,N_2578,N_4430);
nor UO_26 (O_26,N_4770,N_3772);
nor UO_27 (O_27,N_4644,N_4744);
and UO_28 (O_28,N_3280,N_3572);
nand UO_29 (O_29,N_4618,N_3848);
nor UO_30 (O_30,N_4173,N_3130);
xnor UO_31 (O_31,N_3334,N_3232);
xor UO_32 (O_32,N_3753,N_3912);
or UO_33 (O_33,N_4460,N_3684);
or UO_34 (O_34,N_3487,N_4336);
nor UO_35 (O_35,N_4872,N_2607);
xnor UO_36 (O_36,N_4569,N_4010);
xnor UO_37 (O_37,N_3820,N_3491);
and UO_38 (O_38,N_4842,N_3757);
or UO_39 (O_39,N_3709,N_3008);
or UO_40 (O_40,N_3798,N_4449);
xor UO_41 (O_41,N_2762,N_4116);
or UO_42 (O_42,N_3651,N_4308);
nor UO_43 (O_43,N_2568,N_3518);
or UO_44 (O_44,N_4890,N_4617);
or UO_45 (O_45,N_3257,N_2690);
or UO_46 (O_46,N_2533,N_4697);
nand UO_47 (O_47,N_3067,N_3982);
and UO_48 (O_48,N_4303,N_3902);
nand UO_49 (O_49,N_4146,N_2669);
nand UO_50 (O_50,N_3647,N_4100);
nor UO_51 (O_51,N_3219,N_2768);
xor UO_52 (O_52,N_4966,N_4312);
nor UO_53 (O_53,N_2521,N_3297);
xor UO_54 (O_54,N_2901,N_4281);
and UO_55 (O_55,N_3137,N_4534);
nand UO_56 (O_56,N_4447,N_2924);
nor UO_57 (O_57,N_2816,N_4320);
and UO_58 (O_58,N_4335,N_3337);
nand UO_59 (O_59,N_2895,N_2981);
or UO_60 (O_60,N_2755,N_4541);
nand UO_61 (O_61,N_3368,N_4837);
nand UO_62 (O_62,N_4761,N_3455);
nand UO_63 (O_63,N_3197,N_4833);
and UO_64 (O_64,N_4622,N_3627);
and UO_65 (O_65,N_3581,N_2569);
and UO_66 (O_66,N_3842,N_2851);
nor UO_67 (O_67,N_4425,N_2947);
xnor UO_68 (O_68,N_3068,N_4528);
or UO_69 (O_69,N_3775,N_3100);
xor UO_70 (O_70,N_2809,N_4825);
nand UO_71 (O_71,N_4884,N_3055);
or UO_72 (O_72,N_2988,N_4034);
or UO_73 (O_73,N_3620,N_3571);
and UO_74 (O_74,N_4422,N_4530);
or UO_75 (O_75,N_4767,N_2586);
xnor UO_76 (O_76,N_3819,N_4262);
and UO_77 (O_77,N_3425,N_4020);
nor UO_78 (O_78,N_3663,N_4341);
xor UO_79 (O_79,N_3314,N_3510);
nor UO_80 (O_80,N_4278,N_4701);
nand UO_81 (O_81,N_2776,N_3695);
or UO_82 (O_82,N_4003,N_2696);
and UO_83 (O_83,N_3084,N_2567);
nor UO_84 (O_84,N_4994,N_4111);
nand UO_85 (O_85,N_2792,N_3835);
xor UO_86 (O_86,N_4861,N_3866);
nand UO_87 (O_87,N_3611,N_2717);
and UO_88 (O_88,N_2591,N_4630);
xnor UO_89 (O_89,N_4197,N_3097);
or UO_90 (O_90,N_2587,N_4659);
or UO_91 (O_91,N_4046,N_4643);
xnor UO_92 (O_92,N_3287,N_4118);
or UO_93 (O_93,N_2632,N_4348);
and UO_94 (O_94,N_4291,N_3352);
nor UO_95 (O_95,N_3272,N_2619);
xnor UO_96 (O_96,N_4603,N_2500);
nor UO_97 (O_97,N_3029,N_4654);
nor UO_98 (O_98,N_3509,N_2551);
xnor UO_99 (O_99,N_3427,N_4032);
nand UO_100 (O_100,N_4797,N_4554);
or UO_101 (O_101,N_3747,N_2857);
nor UO_102 (O_102,N_3388,N_4527);
or UO_103 (O_103,N_3657,N_3715);
xnor UO_104 (O_104,N_4511,N_4651);
nor UO_105 (O_105,N_3053,N_4267);
nand UO_106 (O_106,N_2878,N_4089);
nand UO_107 (O_107,N_3883,N_4306);
or UO_108 (O_108,N_2608,N_4403);
xor UO_109 (O_109,N_3767,N_4390);
nor UO_110 (O_110,N_4881,N_3876);
and UO_111 (O_111,N_4404,N_4752);
xnor UO_112 (O_112,N_3929,N_3355);
xor UO_113 (O_113,N_4545,N_2940);
and UO_114 (O_114,N_4220,N_4660);
and UO_115 (O_115,N_3700,N_4708);
or UO_116 (O_116,N_4180,N_4192);
nor UO_117 (O_117,N_3448,N_4480);
xnor UO_118 (O_118,N_4414,N_3451);
nand UO_119 (O_119,N_2868,N_3003);
and UO_120 (O_120,N_3814,N_3241);
nand UO_121 (O_121,N_3999,N_3589);
xnor UO_122 (O_122,N_3765,N_3122);
and UO_123 (O_123,N_4393,N_4631);
xnor UO_124 (O_124,N_3552,N_3892);
xor UO_125 (O_125,N_3687,N_3415);
or UO_126 (O_126,N_3006,N_4993);
nand UO_127 (O_127,N_3732,N_3310);
xnor UO_128 (O_128,N_3701,N_4812);
or UO_129 (O_129,N_4371,N_4167);
nand UO_130 (O_130,N_3059,N_3333);
xor UO_131 (O_131,N_4864,N_4462);
or UO_132 (O_132,N_2604,N_3070);
and UO_133 (O_133,N_3735,N_3972);
and UO_134 (O_134,N_3890,N_4027);
and UO_135 (O_135,N_2990,N_4495);
nand UO_136 (O_136,N_4083,N_3307);
nand UO_137 (O_137,N_2715,N_2803);
and UO_138 (O_138,N_3335,N_2800);
nand UO_139 (O_139,N_4457,N_4932);
or UO_140 (O_140,N_2833,N_3258);
and UO_141 (O_141,N_3472,N_3167);
and UO_142 (O_142,N_3490,N_2896);
nor UO_143 (O_143,N_2541,N_3164);
xor UO_144 (O_144,N_3298,N_4839);
and UO_145 (O_145,N_3156,N_4437);
xor UO_146 (O_146,N_3071,N_3279);
xnor UO_147 (O_147,N_3806,N_3222);
nor UO_148 (O_148,N_2508,N_4080);
nand UO_149 (O_149,N_3665,N_3976);
nand UO_150 (O_150,N_4995,N_3664);
nand UO_151 (O_151,N_3135,N_2822);
nor UO_152 (O_152,N_3569,N_4756);
and UO_153 (O_153,N_3824,N_3512);
or UO_154 (O_154,N_4426,N_3142);
nand UO_155 (O_155,N_2745,N_3669);
and UO_156 (O_156,N_3209,N_4633);
xor UO_157 (O_157,N_4268,N_3119);
or UO_158 (O_158,N_2929,N_4448);
xor UO_159 (O_159,N_3990,N_3332);
or UO_160 (O_160,N_4092,N_3066);
xor UO_161 (O_161,N_2864,N_2907);
and UO_162 (O_162,N_2823,N_2594);
nand UO_163 (O_163,N_3690,N_3247);
and UO_164 (O_164,N_2662,N_4366);
and UO_165 (O_165,N_2879,N_2850);
xnor UO_166 (O_166,N_4677,N_2708);
or UO_167 (O_167,N_3399,N_3688);
or UO_168 (O_168,N_3961,N_3954);
xor UO_169 (O_169,N_3243,N_3580);
nor UO_170 (O_170,N_2722,N_4081);
nand UO_171 (O_171,N_3051,N_4407);
and UO_172 (O_172,N_3471,N_3661);
nand UO_173 (O_173,N_3486,N_2785);
nor UO_174 (O_174,N_4624,N_4538);
xor UO_175 (O_175,N_2784,N_3273);
or UO_176 (O_176,N_2853,N_4274);
or UO_177 (O_177,N_4215,N_3719);
nor UO_178 (O_178,N_3005,N_2698);
and UO_179 (O_179,N_4120,N_3398);
nand UO_180 (O_180,N_3967,N_4710);
nand UO_181 (O_181,N_2711,N_3030);
nor UO_182 (O_182,N_3104,N_3846);
xnor UO_183 (O_183,N_4175,N_4595);
nor UO_184 (O_184,N_3072,N_3111);
nand UO_185 (O_185,N_4245,N_3950);
xor UO_186 (O_186,N_4505,N_3549);
or UO_187 (O_187,N_4913,N_2687);
or UO_188 (O_188,N_4087,N_4101);
or UO_189 (O_189,N_4713,N_3930);
nand UO_190 (O_190,N_2659,N_3642);
or UO_191 (O_191,N_4189,N_4299);
nand UO_192 (O_192,N_3565,N_3900);
or UO_193 (O_193,N_4915,N_3422);
nor UO_194 (O_194,N_2621,N_4005);
and UO_195 (O_195,N_3321,N_3240);
and UO_196 (O_196,N_2626,N_2980);
nand UO_197 (O_197,N_2695,N_4035);
nor UO_198 (O_198,N_2517,N_4918);
and UO_199 (O_199,N_4850,N_4158);
and UO_200 (O_200,N_4104,N_4017);
xor UO_201 (O_201,N_4927,N_4056);
nor UO_202 (O_202,N_3102,N_3992);
nor UO_203 (O_203,N_3177,N_4009);
nor UO_204 (O_204,N_4916,N_3027);
nor UO_205 (O_205,N_4269,N_3044);
or UO_206 (O_206,N_4359,N_2970);
and UO_207 (O_207,N_3594,N_4712);
xor UO_208 (O_208,N_4515,N_4834);
and UO_209 (O_209,N_4979,N_3916);
and UO_210 (O_210,N_2771,N_2763);
or UO_211 (O_211,N_3452,N_3389);
and UO_212 (O_212,N_4097,N_3624);
and UO_213 (O_213,N_3026,N_4661);
and UO_214 (O_214,N_3365,N_2653);
nor UO_215 (O_215,N_3980,N_2746);
or UO_216 (O_216,N_2535,N_2652);
xor UO_217 (O_217,N_4729,N_3276);
and UO_218 (O_218,N_2939,N_3837);
and UO_219 (O_219,N_4518,N_2713);
xor UO_220 (O_220,N_3300,N_4902);
and UO_221 (O_221,N_4827,N_3372);
nor UO_222 (O_222,N_4424,N_3376);
and UO_223 (O_223,N_2562,N_3113);
or UO_224 (O_224,N_4085,N_4031);
nand UO_225 (O_225,N_4573,N_4784);
nand UO_226 (O_226,N_2958,N_3911);
nand UO_227 (O_227,N_2821,N_3727);
xnor UO_228 (O_228,N_3694,N_2998);
xor UO_229 (O_229,N_2681,N_3007);
nand UO_230 (O_230,N_3034,N_4679);
and UO_231 (O_231,N_3617,N_4326);
nand UO_232 (O_232,N_3405,N_3459);
nand UO_233 (O_233,N_4304,N_2824);
nor UO_234 (O_234,N_4547,N_4736);
xor UO_235 (O_235,N_3249,N_3416);
or UO_236 (O_236,N_4698,N_4510);
nand UO_237 (O_237,N_4748,N_3898);
xor UO_238 (O_238,N_2691,N_4264);
and UO_239 (O_239,N_4724,N_4657);
and UO_240 (O_240,N_2796,N_2959);
nor UO_241 (O_241,N_2693,N_2994);
nand UO_242 (O_242,N_3004,N_3134);
nor UO_243 (O_243,N_3311,N_4986);
xor UO_244 (O_244,N_3412,N_4914);
nor UO_245 (O_245,N_2510,N_2815);
nor UO_246 (O_246,N_4576,N_2706);
nand UO_247 (O_247,N_4364,N_2571);
or UO_248 (O_248,N_4802,N_4271);
nand UO_249 (O_249,N_2596,N_4164);
and UO_250 (O_250,N_3269,N_4322);
xor UO_251 (O_251,N_2986,N_3373);
nor UO_252 (O_252,N_2775,N_3932);
xnor UO_253 (O_253,N_4760,N_4357);
or UO_254 (O_254,N_3286,N_3751);
or UO_255 (O_255,N_2634,N_4658);
nand UO_256 (O_256,N_3532,N_4774);
and UO_257 (O_257,N_4696,N_4210);
nor UO_258 (O_258,N_2898,N_3691);
xnor UO_259 (O_259,N_4726,N_4506);
nor UO_260 (O_260,N_4128,N_3634);
nor UO_261 (O_261,N_2925,N_2527);
nand UO_262 (O_262,N_2734,N_3385);
xnor UO_263 (O_263,N_3442,N_4593);
nor UO_264 (O_264,N_3575,N_4689);
nand UO_265 (O_265,N_4064,N_4841);
nand UO_266 (O_266,N_3294,N_2649);
xor UO_267 (O_267,N_2881,N_4112);
or UO_268 (O_268,N_3987,N_4805);
or UO_269 (O_269,N_4951,N_3000);
and UO_270 (O_270,N_4566,N_4102);
xnor UO_271 (O_271,N_3506,N_4477);
or UO_272 (O_272,N_2657,N_3585);
nor UO_273 (O_273,N_3720,N_3754);
nor UO_274 (O_274,N_2997,N_3656);
or UO_275 (O_275,N_3414,N_2740);
nor UO_276 (O_276,N_2860,N_4568);
or UO_277 (O_277,N_4857,N_3897);
nor UO_278 (O_278,N_3213,N_4149);
or UO_279 (O_279,N_2518,N_3495);
xnor UO_280 (O_280,N_4715,N_3523);
xnor UO_281 (O_281,N_4800,N_4302);
or UO_282 (O_282,N_3935,N_2766);
nor UO_283 (O_283,N_3221,N_4398);
and UO_284 (O_284,N_3869,N_3022);
and UO_285 (O_285,N_4594,N_4628);
or UO_286 (O_286,N_4882,N_4682);
and UO_287 (O_287,N_4849,N_2609);
or UO_288 (O_288,N_3317,N_2570);
xor UO_289 (O_289,N_2544,N_2631);
nand UO_290 (O_290,N_3304,N_3419);
or UO_291 (O_291,N_3677,N_3176);
or UO_292 (O_292,N_3559,N_4574);
nor UO_293 (O_293,N_3347,N_2991);
or UO_294 (O_294,N_4244,N_4318);
or UO_295 (O_295,N_3864,N_2530);
nand UO_296 (O_296,N_3218,N_3844);
nand UO_297 (O_297,N_4463,N_3136);
and UO_298 (O_298,N_3692,N_2644);
nand UO_299 (O_299,N_3778,N_3957);
xnor UO_300 (O_300,N_4860,N_3162);
or UO_301 (O_301,N_3645,N_3395);
xor UO_302 (O_302,N_3154,N_4996);
nor UO_303 (O_303,N_4261,N_2579);
xor UO_304 (O_304,N_3155,N_4147);
nand UO_305 (O_305,N_4095,N_4362);
xor UO_306 (O_306,N_3390,N_4648);
or UO_307 (O_307,N_3469,N_3584);
nand UO_308 (O_308,N_4421,N_4970);
nor UO_309 (O_309,N_3783,N_3849);
and UO_310 (O_310,N_4777,N_4808);
or UO_311 (O_311,N_4755,N_4943);
or UO_312 (O_312,N_4602,N_3622);
and UO_313 (O_313,N_4279,N_3578);
nand UO_314 (O_314,N_3371,N_4939);
xnor UO_315 (O_315,N_4170,N_2655);
nand UO_316 (O_316,N_4334,N_3944);
or UO_317 (O_317,N_4612,N_2843);
or UO_318 (O_318,N_3785,N_3637);
nor UO_319 (O_319,N_2716,N_3850);
xnor UO_320 (O_320,N_2951,N_4280);
and UO_321 (O_321,N_3949,N_2772);
nor UO_322 (O_322,N_3263,N_4206);
nand UO_323 (O_323,N_3855,N_4925);
or UO_324 (O_324,N_2979,N_3295);
nor UO_325 (O_325,N_2641,N_2782);
nor UO_326 (O_326,N_2559,N_4664);
and UO_327 (O_327,N_4563,N_3567);
nand UO_328 (O_328,N_3141,N_2799);
nand UO_329 (O_329,N_3542,N_2849);
and UO_330 (O_330,N_3843,N_3092);
nand UO_331 (O_331,N_3181,N_2955);
nor UO_332 (O_332,N_3973,N_3322);
and UO_333 (O_333,N_3638,N_3099);
xnor UO_334 (O_334,N_3098,N_2909);
or UO_335 (O_335,N_4840,N_2842);
nand UO_336 (O_336,N_4443,N_3318);
nor UO_337 (O_337,N_2962,N_3417);
xnor UO_338 (O_338,N_4782,N_4687);
or UO_339 (O_339,N_2912,N_3217);
nand UO_340 (O_340,N_3291,N_2507);
and UO_341 (O_341,N_4039,N_4384);
xnor UO_342 (O_342,N_4921,N_3988);
and UO_343 (O_343,N_3953,N_4804);
xnor UO_344 (O_344,N_4181,N_4329);
nand UO_345 (O_345,N_3933,N_2751);
nor UO_346 (O_346,N_4798,N_4903);
xnor UO_347 (O_347,N_4938,N_2777);
xor UO_348 (O_348,N_3986,N_4023);
and UO_349 (O_349,N_4950,N_3153);
nand UO_350 (O_350,N_4340,N_2904);
nor UO_351 (O_351,N_4990,N_3826);
xor UO_352 (O_352,N_4387,N_3201);
nand UO_353 (O_353,N_4917,N_4072);
nand UO_354 (O_354,N_4999,N_3668);
nand UO_355 (O_355,N_4188,N_3117);
xor UO_356 (O_356,N_3501,N_4738);
nor UO_357 (O_357,N_2585,N_3605);
nand UO_358 (O_358,N_4502,N_4956);
nand UO_359 (O_359,N_2774,N_3604);
nand UO_360 (O_360,N_2887,N_4436);
xnor UO_361 (O_361,N_4036,N_2931);
nand UO_362 (O_362,N_4119,N_4106);
xor UO_363 (O_363,N_4022,N_4001);
nand UO_364 (O_364,N_3945,N_3613);
nand UO_365 (O_365,N_3960,N_4942);
nand UO_366 (O_366,N_3182,N_3028);
nor UO_367 (O_367,N_4681,N_2911);
or UO_368 (O_368,N_2589,N_2963);
and UO_369 (O_369,N_4212,N_4786);
or UO_370 (O_370,N_4721,N_3234);
nor UO_371 (O_371,N_3799,N_3714);
and UO_372 (O_372,N_4227,N_3447);
or UO_373 (O_373,N_4004,N_4815);
nand UO_374 (O_374,N_3650,N_4131);
xnor UO_375 (O_375,N_4845,N_4810);
or UO_376 (O_376,N_2950,N_3015);
nand UO_377 (O_377,N_4349,N_4803);
nand UO_378 (O_378,N_3106,N_3252);
xor UO_379 (O_379,N_2856,N_4823);
xor UO_380 (O_380,N_2540,N_3675);
or UO_381 (O_381,N_3020,N_2611);
and UO_382 (O_382,N_2900,N_4632);
or UO_383 (O_383,N_2618,N_3043);
or UO_384 (O_384,N_3872,N_4552);
and UO_385 (O_385,N_4200,N_4099);
and UO_386 (O_386,N_4237,N_4042);
nor UO_387 (O_387,N_2920,N_4202);
xnor UO_388 (O_388,N_2954,N_4732);
and UO_389 (O_389,N_4693,N_4324);
or UO_390 (O_390,N_4746,N_3517);
and UO_391 (O_391,N_2869,N_2828);
or UO_392 (O_392,N_3282,N_2932);
xor UO_393 (O_393,N_4048,N_4452);
or UO_394 (O_394,N_4195,N_2847);
and UO_395 (O_395,N_3941,N_4817);
xnor UO_396 (O_396,N_3636,N_2966);
or UO_397 (O_397,N_3878,N_4580);
nand UO_398 (O_398,N_4363,N_3936);
xor UO_399 (O_399,N_4232,N_2730);
nor UO_400 (O_400,N_2654,N_2913);
and UO_401 (O_401,N_3993,N_2752);
xnor UO_402 (O_402,N_4490,N_4300);
or UO_403 (O_403,N_2889,N_4294);
nor UO_404 (O_404,N_3631,N_3220);
and UO_405 (O_405,N_4720,N_4155);
xor UO_406 (O_406,N_4801,N_3306);
or UO_407 (O_407,N_3265,N_3593);
and UO_408 (O_408,N_4172,N_4584);
xor UO_409 (O_409,N_3095,N_3758);
or UO_410 (O_410,N_4968,N_3516);
xnor UO_411 (O_411,N_3648,N_4372);
and UO_412 (O_412,N_2807,N_3454);
xnor UO_413 (O_413,N_3410,N_4961);
xnor UO_414 (O_414,N_3383,N_3423);
nor UO_415 (O_415,N_4213,N_4507);
nor UO_416 (O_416,N_2989,N_4727);
or UO_417 (O_417,N_3387,N_3401);
xnor UO_418 (O_418,N_4539,N_3770);
or UO_419 (O_419,N_4828,N_2664);
and UO_420 (O_420,N_4821,N_3845);
nor UO_421 (O_421,N_4143,N_3984);
nor UO_422 (O_422,N_4751,N_3671);
nor UO_423 (O_423,N_4735,N_3553);
xnor UO_424 (O_424,N_3983,N_2671);
nand UO_425 (O_425,N_4328,N_4169);
and UO_426 (O_426,N_2741,N_4785);
xor UO_427 (O_427,N_3434,N_4382);
or UO_428 (O_428,N_4521,N_3144);
xor UO_429 (O_429,N_2902,N_2801);
nor UO_430 (O_430,N_4868,N_4855);
and UO_431 (O_431,N_2829,N_4358);
nor UO_432 (O_432,N_3438,N_3568);
xnor UO_433 (O_433,N_4417,N_3315);
or UO_434 (O_434,N_3179,N_4562);
or UO_435 (O_435,N_3851,N_4026);
nand UO_436 (O_436,N_3918,N_4234);
or UO_437 (O_437,N_4565,N_2806);
xor UO_438 (O_438,N_2930,N_4653);
nor UO_439 (O_439,N_4297,N_4768);
or UO_440 (O_440,N_2665,N_4375);
or UO_441 (O_441,N_4470,N_4500);
nand UO_442 (O_442,N_2976,N_3404);
nand UO_443 (O_443,N_3336,N_3363);
nor UO_444 (O_444,N_4647,N_2538);
nor UO_445 (O_445,N_3204,N_3997);
and UO_446 (O_446,N_4386,N_4270);
or UO_447 (O_447,N_3435,N_4413);
xor UO_448 (O_448,N_4105,N_3640);
or UO_449 (O_449,N_2862,N_3309);
xor UO_450 (O_450,N_3323,N_3893);
xor UO_451 (O_451,N_4469,N_3786);
and UO_452 (O_452,N_3236,N_2686);
xnor UO_453 (O_453,N_4290,N_3610);
nor UO_454 (O_454,N_4783,N_4088);
or UO_455 (O_455,N_3917,N_4723);
or UO_456 (O_456,N_4050,N_4028);
xor UO_457 (O_457,N_4492,N_3833);
xnor UO_458 (O_458,N_3150,N_3426);
or UO_459 (O_459,N_3551,N_4114);
nand UO_460 (O_460,N_4959,N_3696);
and UO_461 (O_461,N_3989,N_4965);
nor UO_462 (O_462,N_3382,N_3524);
nand UO_463 (O_463,N_4650,N_4456);
and UO_464 (O_464,N_4263,N_4799);
nand UO_465 (O_465,N_3428,N_2922);
nor UO_466 (O_466,N_4620,N_2590);
nand UO_467 (O_467,N_4862,N_3299);
nand UO_468 (O_468,N_4455,N_3958);
or UO_469 (O_469,N_4905,N_3208);
nor UO_470 (O_470,N_3206,N_4920);
or UO_471 (O_471,N_4499,N_4781);
xnor UO_472 (O_472,N_4501,N_3035);
nand UO_473 (O_473,N_2514,N_3995);
xnor UO_474 (O_474,N_4867,N_4895);
nor UO_475 (O_475,N_2606,N_3598);
xor UO_476 (O_476,N_2599,N_4084);
nor UO_477 (O_477,N_3562,N_4504);
or UO_478 (O_478,N_4123,N_4242);
or UO_479 (O_479,N_3172,N_3822);
xor UO_480 (O_480,N_4476,N_3124);
xnor UO_481 (O_481,N_3074,N_3573);
xnor UO_482 (O_482,N_3614,N_4226);
nor UO_483 (O_483,N_4497,N_4816);
nand UO_484 (O_484,N_3112,N_4338);
nand UO_485 (O_485,N_4758,N_3231);
xor UO_486 (O_486,N_3238,N_3939);
nor UO_487 (O_487,N_4305,N_2612);
and UO_488 (O_488,N_3259,N_4636);
nand UO_489 (O_489,N_4018,N_2511);
xnor UO_490 (O_490,N_3357,N_3492);
and UO_491 (O_491,N_4233,N_4402);
nor UO_492 (O_492,N_4982,N_4055);
or UO_493 (O_493,N_3227,N_4874);
xor UO_494 (O_494,N_3762,N_3977);
nor UO_495 (O_495,N_4060,N_3202);
nor UO_496 (O_496,N_4955,N_4174);
xnor UO_497 (O_497,N_4514,N_2812);
and UO_498 (O_498,N_3752,N_3557);
and UO_499 (O_499,N_4540,N_2867);
xnor UO_500 (O_500,N_4021,N_4139);
nor UO_501 (O_501,N_4984,N_4875);
nand UO_502 (O_502,N_3270,N_4716);
nand UO_503 (O_503,N_3519,N_4794);
nand UO_504 (O_504,N_2526,N_3036);
and UO_505 (O_505,N_3621,N_3597);
and UO_506 (O_506,N_2855,N_2735);
nand UO_507 (O_507,N_3782,N_4714);
or UO_508 (O_508,N_3031,N_4711);
nand UO_509 (O_509,N_3174,N_3560);
nor UO_510 (O_510,N_2760,N_2539);
nand UO_511 (O_511,N_2971,N_2863);
xnor UO_512 (O_512,N_4091,N_2531);
xnor UO_513 (O_513,N_3358,N_4985);
xor UO_514 (O_514,N_4236,N_2817);
nand UO_515 (O_515,N_3545,N_3793);
xor UO_516 (O_516,N_3616,N_3513);
xnor UO_517 (O_517,N_3339,N_4796);
and UO_518 (O_518,N_3840,N_3639);
nand UO_519 (O_519,N_4079,N_4395);
nor UO_520 (O_520,N_4829,N_4779);
and UO_521 (O_521,N_3655,N_3533);
and UO_522 (O_522,N_3125,N_3625);
nor UO_523 (O_523,N_2961,N_2905);
or UO_524 (O_524,N_3952,N_4581);
nor UO_525 (O_525,N_3630,N_3108);
nor UO_526 (O_526,N_3725,N_4700);
nand UO_527 (O_527,N_3940,N_3577);
xnor UO_528 (O_528,N_4063,N_4121);
nand UO_529 (O_529,N_3094,N_4561);
and UO_530 (O_530,N_4016,N_3615);
or UO_531 (O_531,N_4906,N_4228);
xor UO_532 (O_532,N_3996,N_3407);
xor UO_533 (O_533,N_3229,N_2573);
and UO_534 (O_534,N_3576,N_4989);
xor UO_535 (O_535,N_4641,N_4656);
and UO_536 (O_536,N_3366,N_2682);
xnor UO_537 (O_537,N_3450,N_2504);
or UO_538 (O_538,N_3090,N_3255);
nand UO_539 (O_539,N_4879,N_4978);
and UO_540 (O_540,N_2791,N_2874);
or UO_541 (O_541,N_3374,N_4394);
xor UO_542 (O_542,N_4339,N_4704);
nor UO_543 (O_543,N_2648,N_2859);
nand UO_544 (O_544,N_4190,N_3324);
xnor UO_545 (O_545,N_3400,N_3504);
and UO_546 (O_546,N_3583,N_3200);
nand UO_547 (O_547,N_4473,N_3686);
or UO_548 (O_548,N_4688,N_2719);
xor UO_549 (O_549,N_4446,N_3760);
nand UO_550 (O_550,N_2852,N_4012);
nor UO_551 (O_551,N_3659,N_4272);
or UO_552 (O_552,N_4258,N_4680);
xor UO_553 (O_553,N_3178,N_3737);
xnor UO_554 (O_554,N_3731,N_4482);
nor UO_555 (O_555,N_2575,N_4675);
or UO_556 (O_556,N_2576,N_4273);
or UO_557 (O_557,N_3346,N_4002);
nand UO_558 (O_558,N_3923,N_2557);
nor UO_559 (O_559,N_3284,N_4707);
nand UO_560 (O_560,N_4019,N_4221);
and UO_561 (O_561,N_3681,N_4287);
or UO_562 (O_562,N_4807,N_4887);
or UO_563 (O_563,N_4075,N_3702);
or UO_564 (O_564,N_4564,N_4053);
and UO_565 (O_565,N_4379,N_2773);
nand UO_566 (O_566,N_3955,N_2999);
and UO_567 (O_567,N_2670,N_2965);
nand UO_568 (O_568,N_3350,N_3394);
xor UO_569 (O_569,N_4361,N_3380);
or UO_570 (O_570,N_4625,N_4793);
and UO_571 (O_571,N_4438,N_3853);
nand UO_572 (O_572,N_3143,N_3804);
or UO_573 (O_573,N_4040,N_4558);
xnor UO_574 (O_574,N_2616,N_2598);
xor UO_575 (O_575,N_3756,N_3277);
or UO_576 (O_576,N_3803,N_2754);
nand UO_577 (O_577,N_4525,N_3828);
nor UO_578 (O_578,N_3777,N_4876);
and UO_579 (O_579,N_4773,N_2685);
nor UO_580 (O_580,N_3402,N_3788);
or UO_581 (O_581,N_4185,N_3761);
nor UO_582 (O_582,N_3345,N_2882);
and UO_583 (O_583,N_4360,N_4891);
or UO_584 (O_584,N_3467,N_3823);
nand UO_585 (O_585,N_4259,N_2880);
nor UO_586 (O_586,N_2790,N_4526);
nand UO_587 (O_587,N_4549,N_3809);
nor UO_588 (O_588,N_3429,N_4356);
xnor UO_589 (O_589,N_4858,N_2702);
nand UO_590 (O_590,N_3019,N_3290);
and UO_591 (O_591,N_2636,N_3706);
or UO_592 (O_592,N_4140,N_2942);
xnor UO_593 (O_593,N_3319,N_2873);
or UO_594 (O_594,N_3496,N_2767);
or UO_595 (O_595,N_2605,N_2732);
nand UO_596 (O_596,N_2972,N_3460);
and UO_597 (O_597,N_4316,N_4239);
nor UO_598 (O_598,N_2624,N_3152);
or UO_599 (O_599,N_3882,N_3121);
xnor UO_600 (O_600,N_3726,N_2622);
nand UO_601 (O_601,N_3424,N_3602);
and UO_602 (O_602,N_3716,N_4788);
nand UO_603 (O_603,N_2543,N_2558);
xor UO_604 (O_604,N_4865,N_2872);
and UO_605 (O_605,N_2704,N_4179);
or UO_606 (O_606,N_3887,N_4255);
xnor UO_607 (O_607,N_3086,N_2703);
or UO_608 (O_608,N_3861,N_3449);
xnor UO_609 (O_609,N_3445,N_4029);
or UO_610 (O_610,N_2628,N_3539);
xor UO_611 (O_611,N_3579,N_4388);
nand UO_612 (O_612,N_3025,N_3769);
xnor UO_613 (O_613,N_4912,N_2712);
nand UO_614 (O_614,N_4493,N_4922);
nor UO_615 (O_615,N_4045,N_4519);
and UO_616 (O_616,N_4427,N_3351);
xor UO_617 (O_617,N_4136,N_4132);
and UO_618 (O_618,N_4591,N_4054);
and UO_619 (O_619,N_2888,N_2841);
xor UO_620 (O_620,N_4694,N_4963);
xnor UO_621 (O_621,N_3779,N_4750);
and UO_622 (O_622,N_4487,N_4043);
nor UO_623 (O_623,N_2556,N_4718);
xnor UO_624 (O_624,N_2903,N_4333);
or UO_625 (O_625,N_4376,N_2656);
nand UO_626 (O_626,N_4908,N_3342);
xor UO_627 (O_627,N_4898,N_3488);
nor UO_628 (O_628,N_3856,N_4293);
nand UO_629 (O_629,N_4323,N_3254);
nor UO_630 (O_630,N_4678,N_4652);
and UO_631 (O_631,N_3313,N_3673);
nor UO_632 (O_632,N_3275,N_4820);
nor UO_633 (O_633,N_2593,N_4577);
nor UO_634 (O_634,N_2705,N_4669);
xnor UO_635 (O_635,N_3749,N_3062);
and UO_636 (O_636,N_4640,N_4649);
or UO_637 (O_637,N_3948,N_4465);
or UO_638 (O_638,N_2721,N_2506);
or UO_639 (O_639,N_4844,N_3834);
nand UO_640 (O_640,N_2977,N_2753);
and UO_641 (O_641,N_3626,N_2505);
nor UO_642 (O_642,N_4766,N_3159);
nand UO_643 (O_643,N_4094,N_3138);
xor UO_644 (O_644,N_3807,N_4466);
nor UO_645 (O_645,N_3894,N_4877);
nand UO_646 (O_646,N_4742,N_4159);
and UO_647 (O_647,N_4517,N_4408);
or UO_648 (O_648,N_3080,N_3635);
nor UO_649 (O_649,N_3666,N_3338);
nor UO_650 (O_650,N_3722,N_3479);
nand UO_651 (O_651,N_3129,N_4150);
xor UO_652 (O_652,N_4429,N_4184);
nand UO_653 (O_653,N_4975,N_2758);
nor UO_654 (O_654,N_3261,N_2750);
nand UO_655 (O_655,N_4265,N_4243);
nor UO_656 (O_656,N_3235,N_4997);
and UO_657 (O_657,N_3498,N_4960);
xnor UO_658 (O_658,N_3391,N_3789);
or UO_659 (O_659,N_4141,N_4683);
and UO_660 (O_660,N_2661,N_4325);
nor UO_661 (O_661,N_4899,N_3013);
or UO_662 (O_662,N_3002,N_3045);
nand UO_663 (O_663,N_3123,N_3436);
or UO_664 (O_664,N_3056,N_2765);
or UO_665 (O_665,N_2525,N_4531);
nor UO_666 (O_666,N_4148,N_3962);
nor UO_667 (O_667,N_4301,N_3768);
nand UO_668 (O_668,N_4352,N_4972);
nand UO_669 (O_669,N_4211,N_3784);
or UO_670 (O_670,N_2623,N_4074);
nor UO_671 (O_671,N_3001,N_3406);
and UO_672 (O_672,N_4156,N_4607);
xor UO_673 (O_673,N_4909,N_2726);
and UO_674 (O_674,N_4733,N_3507);
or UO_675 (O_675,N_3528,N_4699);
or UO_676 (O_676,N_3505,N_3830);
nand UO_677 (O_677,N_4067,N_2937);
nand UO_678 (O_678,N_3362,N_4848);
nand UO_679 (O_679,N_3260,N_4623);
and UO_680 (O_680,N_4771,N_3131);
or UO_681 (O_681,N_2643,N_2733);
or UO_682 (O_682,N_4415,N_2503);
nor UO_683 (O_683,N_2630,N_2629);
or UO_684 (O_684,N_2697,N_4252);
or UO_685 (O_685,N_3285,N_3343);
or UO_686 (O_686,N_4103,N_4832);
and UO_687 (O_687,N_3473,N_4217);
nor UO_688 (O_688,N_3361,N_4586);
and UO_689 (O_689,N_3904,N_4248);
or UO_690 (O_690,N_3871,N_4575);
nand UO_691 (O_691,N_4605,N_3289);
nor UO_692 (O_692,N_3205,N_2637);
nand UO_693 (O_693,N_3493,N_3485);
and UO_694 (O_694,N_4667,N_4177);
nand UO_695 (O_695,N_4722,N_2996);
nor UO_696 (O_696,N_4754,N_3320);
xnor UO_697 (O_697,N_3790,N_3858);
or UO_698 (O_698,N_3239,N_4059);
nand UO_699 (O_699,N_3811,N_2844);
nor UO_700 (O_700,N_4741,N_4481);
nand UO_701 (O_701,N_3711,N_2866);
xnor UO_702 (O_702,N_3704,N_3744);
nand UO_703 (O_703,N_3375,N_3712);
or UO_704 (O_704,N_4183,N_3120);
nor UO_705 (O_705,N_2769,N_4524);
or UO_706 (O_706,N_3359,N_4824);
nand UO_707 (O_707,N_4560,N_3541);
xor UO_708 (O_708,N_4383,N_2808);
or UO_709 (O_709,N_3548,N_3966);
nand UO_710 (O_710,N_4310,N_4052);
nand UO_711 (O_711,N_3190,N_4163);
and UO_712 (O_712,N_2891,N_2846);
xor UO_713 (O_713,N_2679,N_4818);
or UO_714 (O_714,N_4491,N_3743);
nand UO_715 (O_715,N_2674,N_4635);
nand UO_716 (O_716,N_2710,N_2883);
xnor UO_717 (O_717,N_4201,N_2633);
nand UO_718 (O_718,N_4516,N_3194);
or UO_719 (O_719,N_4168,N_4907);
or UO_720 (O_720,N_2943,N_3601);
or UO_721 (O_721,N_4078,N_2827);
and UO_722 (O_722,N_2995,N_2876);
and UO_723 (O_723,N_4789,N_4690);
nand UO_724 (O_724,N_2700,N_4936);
xnor UO_725 (O_725,N_3740,N_3212);
nand UO_726 (O_726,N_4637,N_3191);
nand UO_727 (O_727,N_3327,N_2545);
or UO_728 (O_728,N_4957,N_3908);
nor UO_729 (O_729,N_3674,N_3476);
and UO_730 (O_730,N_4854,N_2688);
or UO_731 (O_731,N_3161,N_3118);
nand UO_732 (O_732,N_3910,N_3433);
or UO_733 (O_733,N_2663,N_3808);
xnor UO_734 (O_734,N_2871,N_3812);
nor UO_735 (O_735,N_3114,N_3033);
or UO_736 (O_736,N_3482,N_3603);
or UO_737 (O_737,N_4125,N_3017);
xnor UO_738 (O_738,N_4737,N_2678);
and UO_739 (O_739,N_3981,N_4472);
xnor UO_740 (O_740,N_2982,N_3195);
and UO_741 (O_741,N_3256,N_3998);
or UO_742 (O_742,N_3538,N_3021);
and UO_743 (O_743,N_4673,N_4747);
or UO_744 (O_744,N_4847,N_3207);
or UO_745 (O_745,N_4420,N_2778);
nor UO_746 (O_746,N_3956,N_3520);
or UO_747 (O_747,N_2793,N_4076);
xnor UO_748 (O_748,N_2779,N_3014);
nand UO_749 (O_749,N_3188,N_3558);
nor UO_750 (O_750,N_3899,N_2906);
nand UO_751 (O_751,N_3047,N_4901);
nor UO_752 (O_752,N_3081,N_3959);
or UO_753 (O_753,N_3057,N_2673);
and UO_754 (O_754,N_2941,N_2804);
xor UO_755 (O_755,N_4134,N_4033);
nand UO_756 (O_756,N_2554,N_3540);
and UO_757 (O_757,N_3180,N_4171);
nor UO_758 (O_758,N_2588,N_3228);
nand UO_759 (O_759,N_4911,N_3886);
xor UO_760 (O_760,N_3379,N_2707);
and UO_761 (O_761,N_3088,N_3091);
xnor UO_762 (O_762,N_4015,N_4377);
xnor UO_763 (O_763,N_4399,N_4488);
and UO_764 (O_764,N_3742,N_3211);
xnor UO_765 (O_765,N_4706,N_4285);
and UO_766 (O_766,N_4601,N_4826);
xnor UO_767 (O_767,N_4090,N_3464);
nor UO_768 (O_768,N_3151,N_3420);
and UO_769 (O_769,N_3042,N_4634);
nand UO_770 (O_770,N_2625,N_3224);
or UO_771 (O_771,N_3083,N_3946);
and UO_772 (O_772,N_2914,N_3233);
nor UO_773 (O_773,N_4740,N_2523);
xor UO_774 (O_774,N_3292,N_2672);
or UO_775 (O_775,N_4277,N_3745);
nor UO_776 (O_776,N_2692,N_2757);
xnor UO_777 (O_777,N_4971,N_4513);
and UO_778 (O_778,N_4642,N_4806);
nor UO_779 (O_779,N_3296,N_4373);
or UO_780 (O_780,N_3913,N_3024);
or UO_781 (O_781,N_4717,N_4629);
and UO_782 (O_782,N_4250,N_3730);
and UO_783 (O_783,N_4014,N_3763);
and UO_784 (O_784,N_4934,N_4572);
nand UO_785 (O_785,N_3199,N_4949);
nor UO_786 (O_786,N_4599,N_4638);
or UO_787 (O_787,N_3531,N_3048);
xnor UO_788 (O_788,N_4830,N_4822);
nor UO_789 (O_789,N_3349,N_4431);
or UO_790 (O_790,N_4223,N_3353);
nor UO_791 (O_791,N_3543,N_2749);
xor UO_792 (O_792,N_2583,N_4194);
xnor UO_793 (O_793,N_4070,N_4433);
or UO_794 (O_794,N_2780,N_4196);
or UO_795 (O_795,N_2666,N_3369);
nand UO_796 (O_796,N_4671,N_3440);
xor UO_797 (O_797,N_3116,N_2938);
and UO_798 (O_798,N_3774,N_2848);
nand UO_799 (O_799,N_4665,N_3340);
xnor UO_800 (O_800,N_3994,N_4257);
and UO_801 (O_801,N_3109,N_2918);
xnor UO_802 (O_802,N_4401,N_4249);
and UO_803 (O_803,N_3698,N_4992);
nand UO_804 (O_804,N_3776,N_3942);
nor UO_805 (O_805,N_3444,N_3367);
or UO_806 (O_806,N_3646,N_4444);
nor UO_807 (O_807,N_3418,N_4082);
xnor UO_808 (O_808,N_3189,N_2908);
nand UO_809 (O_809,N_3266,N_3386);
and UO_810 (O_810,N_4222,N_4948);
nor UO_811 (O_811,N_4919,N_4145);
or UO_812 (O_812,N_2595,N_3978);
nand UO_813 (O_813,N_2714,N_4073);
nor UO_814 (O_814,N_4567,N_2933);
or UO_815 (O_815,N_2946,N_4684);
nor UO_816 (O_816,N_3801,N_4535);
nor UO_817 (O_817,N_3925,N_3965);
and UO_818 (O_818,N_4247,N_2709);
nor UO_819 (O_819,N_4973,N_2818);
xnor UO_820 (O_820,N_4354,N_4451);
and UO_821 (O_821,N_2581,N_3530);
nor UO_822 (O_822,N_3590,N_3262);
and UO_823 (O_823,N_4315,N_3489);
xnor UO_824 (O_824,N_2813,N_3529);
or UO_825 (O_825,N_4570,N_2537);
nand UO_826 (O_826,N_4589,N_3521);
or UO_827 (O_827,N_2890,N_4935);
or UO_828 (O_828,N_3308,N_3914);
or UO_829 (O_829,N_3246,N_2957);
and UO_830 (O_830,N_4662,N_2826);
xnor UO_831 (O_831,N_4235,N_3078);
nand UO_832 (O_832,N_2720,N_4663);
nor UO_833 (O_833,N_4191,N_4672);
and UO_834 (O_834,N_2646,N_2845);
xnor UO_835 (O_835,N_3554,N_4160);
nor UO_836 (O_836,N_2795,N_4246);
xor UO_837 (O_837,N_3484,N_4115);
nor UO_838 (O_838,N_2884,N_3468);
or UO_839 (O_839,N_2743,N_3921);
nor UO_840 (O_840,N_3149,N_3168);
nand UO_841 (O_841,N_3293,N_4619);
or UO_842 (O_842,N_2620,N_3570);
nor UO_843 (O_843,N_3274,N_4616);
nand UO_844 (O_844,N_2820,N_3873);
or UO_845 (O_845,N_3430,N_4343);
nand UO_846 (O_846,N_3166,N_2524);
or UO_847 (O_847,N_3739,N_2677);
or UO_848 (O_848,N_3556,N_3587);
xor UO_849 (O_849,N_3069,N_3115);
nand UO_850 (O_850,N_3802,N_2877);
nand UO_851 (O_851,N_3723,N_3160);
nand UO_852 (O_852,N_4703,N_3815);
nand UO_853 (O_853,N_4321,N_3248);
nand UO_854 (O_854,N_4953,N_3920);
and UO_855 (O_855,N_4969,N_4557);
or UO_856 (O_856,N_4178,N_2580);
nor UO_857 (O_857,N_4686,N_3764);
xnor UO_858 (O_858,N_3413,N_2926);
nand UO_859 (O_859,N_3874,N_2603);
xor UO_860 (O_860,N_4551,N_3644);
nand UO_861 (O_861,N_2738,N_4937);
or UO_862 (O_862,N_4892,N_4439);
and UO_863 (O_863,N_4400,N_3527);
and UO_864 (O_864,N_2564,N_4410);
or UO_865 (O_865,N_3600,N_4154);
xor UO_866 (O_866,N_4049,N_3907);
nor UO_867 (O_867,N_4489,N_2520);
and UO_868 (O_868,N_4674,N_3264);
nand UO_869 (O_869,N_2574,N_3443);
xnor UO_870 (O_870,N_2694,N_2787);
and UO_871 (O_871,N_4725,N_3810);
or UO_872 (O_872,N_2885,N_4428);
and UO_873 (O_873,N_3728,N_4520);
and UO_874 (O_874,N_3192,N_4298);
nand UO_875 (O_875,N_4475,N_3857);
nor UO_876 (O_876,N_4980,N_4093);
nand UO_877 (O_877,N_3105,N_3535);
xor UO_878 (O_878,N_4900,N_3670);
and UO_879 (O_879,N_4947,N_2718);
and UO_880 (O_880,N_4691,N_3458);
xor UO_881 (O_881,N_3018,N_3432);
or UO_882 (O_882,N_2832,N_3713);
xor UO_883 (O_883,N_2916,N_3370);
nand UO_884 (O_884,N_3915,N_4276);
or UO_885 (O_885,N_3127,N_2825);
and UO_886 (O_886,N_4107,N_3063);
xnor UO_887 (O_887,N_2728,N_3508);
nand UO_888 (O_888,N_3147,N_3838);
or UO_889 (O_889,N_3077,N_4759);
nand UO_890 (O_890,N_4370,N_3278);
nor UO_891 (O_891,N_4941,N_4332);
and UO_892 (O_892,N_2969,N_4350);
nor UO_893 (O_893,N_3171,N_4836);
or UO_894 (O_894,N_2747,N_2893);
nor UO_895 (O_895,N_3547,N_3676);
and UO_896 (O_896,N_2865,N_4838);
nand UO_897 (O_897,N_4450,N_3478);
and UO_898 (O_898,N_4124,N_3421);
and UO_899 (O_899,N_3733,N_4416);
and UO_900 (O_900,N_2945,N_4044);
or UO_901 (O_901,N_4435,N_4787);
and UO_902 (O_902,N_3185,N_4047);
or UO_903 (O_903,N_4958,N_4266);
nor UO_904 (O_904,N_3555,N_2934);
nand UO_905 (O_905,N_3741,N_3483);
or UO_906 (O_906,N_4923,N_4351);
and UO_907 (O_907,N_3499,N_3564);
nand UO_908 (O_908,N_4461,N_3859);
nand UO_909 (O_909,N_4135,N_2724);
nor UO_910 (O_910,N_3403,N_2731);
xor UO_911 (O_911,N_4030,N_3868);
nand UO_912 (O_912,N_3328,N_4127);
or UO_913 (O_913,N_3909,N_3326);
xnor UO_914 (O_914,N_2748,N_2565);
nor UO_915 (O_915,N_4484,N_4284);
xor UO_916 (O_916,N_2788,N_3841);
and UO_917 (O_917,N_4331,N_3682);
nor UO_918 (O_918,N_3165,N_4928);
nor UO_919 (O_919,N_3724,N_3173);
and UO_920 (O_920,N_2532,N_4319);
and UO_921 (O_921,N_4878,N_3107);
xnor UO_922 (O_922,N_2553,N_4709);
and UO_923 (O_923,N_4011,N_3132);
and UO_924 (O_924,N_4790,N_2516);
nand UO_925 (O_925,N_3689,N_3302);
xor UO_926 (O_926,N_4256,N_3896);
and UO_927 (O_927,N_3446,N_4086);
and UO_928 (O_928,N_3494,N_4186);
and UO_929 (O_929,N_4153,N_4883);
xnor UO_930 (O_930,N_2522,N_2983);
nand UO_931 (O_931,N_2899,N_4555);
nand UO_932 (O_932,N_3064,N_3526);
nand UO_933 (O_933,N_2935,N_4389);
and UO_934 (O_934,N_4007,N_4705);
or UO_935 (O_935,N_4983,N_4254);
nand UO_936 (O_936,N_3087,N_2647);
and UO_937 (O_937,N_4345,N_3680);
xor UO_938 (O_938,N_2613,N_2615);
nor UO_939 (O_939,N_3974,N_4609);
or UO_940 (O_940,N_2676,N_2645);
nor UO_941 (O_941,N_4122,N_3175);
or UO_942 (O_942,N_4685,N_4342);
nor UO_943 (O_943,N_3356,N_3829);
or UO_944 (O_944,N_4964,N_2550);
nand UO_945 (O_945,N_4814,N_3619);
and UO_946 (O_946,N_4792,N_3037);
and UO_947 (O_947,N_4542,N_4406);
or UO_948 (O_948,N_3503,N_3881);
and UO_949 (O_949,N_4757,N_4550);
nor UO_950 (O_950,N_3023,N_3825);
nor UO_951 (O_951,N_3797,N_2744);
or UO_952 (O_952,N_3329,N_4109);
or UO_953 (O_953,N_3591,N_4852);
nor UO_954 (O_954,N_3183,N_3678);
and UO_955 (O_955,N_3606,N_2978);
or UO_956 (O_956,N_3093,N_4598);
xnor UO_957 (O_957,N_4695,N_4098);
nand UO_958 (O_958,N_4819,N_4998);
and UO_959 (O_959,N_4275,N_2642);
nand UO_960 (O_960,N_4791,N_4311);
nor UO_961 (O_961,N_4897,N_4544);
xor UO_962 (O_962,N_4946,N_2974);
or UO_963 (O_963,N_3061,N_4933);
and UO_964 (O_964,N_2992,N_3928);
nor UO_965 (O_965,N_4904,N_4412);
nor UO_966 (O_966,N_3870,N_3934);
or UO_967 (O_967,N_3623,N_2597);
or UO_968 (O_968,N_4762,N_3889);
xor UO_969 (O_969,N_2897,N_4893);
and UO_970 (O_970,N_4385,N_2683);
and UO_971 (O_971,N_2501,N_4646);
nand UO_972 (O_972,N_2534,N_3612);
nor UO_973 (O_973,N_2555,N_2723);
and UO_974 (O_974,N_4231,N_3392);
or UO_975 (O_975,N_3658,N_3312);
nand UO_976 (O_976,N_4405,N_4330);
nand UO_977 (O_977,N_3225,N_4396);
xnor UO_978 (O_978,N_2680,N_4944);
xor UO_979 (O_979,N_4529,N_3079);
or UO_980 (O_980,N_4108,N_3880);
xnor UO_981 (O_981,N_2886,N_4474);
nand UO_982 (O_982,N_3364,N_3561);
xnor UO_983 (O_983,N_4381,N_3214);
nand UO_984 (O_984,N_4831,N_4133);
xnor UO_985 (O_985,N_4945,N_4835);
nor UO_986 (O_986,N_3905,N_3378);
xnor UO_987 (O_987,N_2936,N_2552);
xnor UO_988 (O_988,N_4702,N_3629);
xnor UO_989 (O_989,N_2549,N_4260);
or UO_990 (O_990,N_4126,N_3431);
and UO_991 (O_991,N_4585,N_4764);
nand UO_992 (O_992,N_3052,N_4668);
and UO_993 (O_993,N_3466,N_4871);
and UO_994 (O_994,N_2727,N_3906);
nand UO_995 (O_995,N_3462,N_3805);
xor UO_996 (O_996,N_3497,N_3453);
nand UO_997 (O_997,N_3901,N_4117);
nor UO_998 (O_998,N_3759,N_4296);
xor UO_999 (O_999,N_3465,N_4205);
endmodule