module basic_500_3000_500_15_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_85,In_495);
and U1 (N_1,In_421,In_325);
and U2 (N_2,In_418,In_396);
and U3 (N_3,In_1,In_38);
nor U4 (N_4,In_130,In_7);
xor U5 (N_5,In_8,In_267);
nor U6 (N_6,In_382,In_19);
or U7 (N_7,In_84,In_18);
nand U8 (N_8,In_333,In_24);
xnor U9 (N_9,In_434,In_385);
and U10 (N_10,In_33,In_304);
or U11 (N_11,In_457,In_11);
nand U12 (N_12,In_363,In_209);
or U13 (N_13,In_136,In_307);
or U14 (N_14,In_192,In_237);
nor U15 (N_15,In_365,In_378);
and U16 (N_16,In_171,In_452);
or U17 (N_17,In_331,In_224);
and U18 (N_18,In_187,In_42);
and U19 (N_19,In_47,In_108);
nor U20 (N_20,In_334,In_362);
and U21 (N_21,In_262,In_266);
or U22 (N_22,In_99,In_290);
nand U23 (N_23,In_299,In_355);
or U24 (N_24,In_463,In_249);
xor U25 (N_25,In_359,In_183);
or U26 (N_26,In_121,In_79);
nor U27 (N_27,In_52,In_459);
nor U28 (N_28,In_427,In_32);
or U29 (N_29,In_155,In_438);
and U30 (N_30,In_408,In_360);
and U31 (N_31,In_301,In_88);
and U32 (N_32,In_94,In_356);
nor U33 (N_33,In_309,In_219);
nand U34 (N_34,In_461,In_257);
and U35 (N_35,In_291,In_156);
nor U36 (N_36,In_428,In_244);
or U37 (N_37,In_71,In_12);
nor U38 (N_38,In_345,In_271);
or U39 (N_39,In_195,In_473);
nand U40 (N_40,In_37,In_150);
or U41 (N_41,In_90,In_14);
or U42 (N_42,In_404,In_200);
nand U43 (N_43,In_313,In_422);
nor U44 (N_44,In_339,In_120);
and U45 (N_45,In_62,In_319);
or U46 (N_46,In_321,In_269);
and U47 (N_47,In_26,In_369);
nor U48 (N_48,In_83,In_31);
nand U49 (N_49,In_186,In_435);
and U50 (N_50,In_391,In_45);
and U51 (N_51,In_161,In_188);
and U52 (N_52,In_53,In_380);
nor U53 (N_53,In_185,In_194);
and U54 (N_54,In_276,In_476);
and U55 (N_55,In_167,In_118);
nand U56 (N_56,In_207,In_253);
and U57 (N_57,In_481,In_450);
nand U58 (N_58,In_328,In_420);
nor U59 (N_59,In_112,In_160);
nand U60 (N_60,In_223,In_446);
and U61 (N_61,In_462,In_116);
or U62 (N_62,In_451,In_371);
nand U63 (N_63,In_117,In_104);
nor U64 (N_64,In_379,In_179);
and U65 (N_65,In_381,In_20);
nand U66 (N_66,In_89,In_289);
nand U67 (N_67,In_281,In_165);
and U68 (N_68,In_341,In_443);
nand U69 (N_69,In_139,In_402);
or U70 (N_70,In_412,In_211);
and U71 (N_71,In_105,In_425);
nor U72 (N_72,In_305,In_140);
nor U73 (N_73,In_372,In_449);
and U74 (N_74,In_335,In_256);
nor U75 (N_75,In_115,In_270);
or U76 (N_76,In_190,In_230);
nor U77 (N_77,In_357,In_338);
nand U78 (N_78,In_125,In_35);
or U79 (N_79,In_22,In_431);
or U80 (N_80,In_184,In_212);
nor U81 (N_81,In_3,In_407);
nor U82 (N_82,In_275,In_478);
nor U83 (N_83,In_36,In_370);
and U84 (N_84,In_133,In_92);
nand U85 (N_85,In_13,In_264);
nor U86 (N_86,In_352,In_86);
nor U87 (N_87,In_292,In_484);
nand U88 (N_88,In_245,In_152);
and U89 (N_89,In_166,In_241);
or U90 (N_90,In_469,In_197);
or U91 (N_91,In_260,In_274);
and U92 (N_92,In_442,In_231);
and U93 (N_93,In_43,In_168);
or U94 (N_94,In_318,In_100);
and U95 (N_95,In_220,In_398);
or U96 (N_96,In_440,In_426);
and U97 (N_97,In_263,In_388);
nand U98 (N_98,In_377,In_173);
xnor U99 (N_99,In_413,In_448);
and U100 (N_100,In_98,In_323);
nor U101 (N_101,In_49,In_272);
or U102 (N_102,In_122,In_393);
and U103 (N_103,In_399,In_466);
and U104 (N_104,In_21,In_460);
nand U105 (N_105,In_491,In_222);
or U106 (N_106,In_114,In_154);
nand U107 (N_107,In_251,In_170);
nor U108 (N_108,In_87,In_454);
or U109 (N_109,In_475,In_479);
or U110 (N_110,In_445,In_236);
and U111 (N_111,In_178,In_169);
nand U112 (N_112,In_401,In_347);
nand U113 (N_113,In_293,In_193);
nor U114 (N_114,In_483,In_308);
nand U115 (N_115,In_181,In_414);
nand U116 (N_116,In_282,In_390);
nand U117 (N_117,In_409,In_10);
and U118 (N_118,In_471,In_158);
and U119 (N_119,In_430,In_239);
nand U120 (N_120,In_59,In_214);
and U121 (N_121,In_280,In_141);
nand U122 (N_122,In_488,In_238);
nor U123 (N_123,In_261,In_278);
nand U124 (N_124,In_374,In_157);
or U125 (N_125,In_68,In_288);
nand U126 (N_126,In_327,In_135);
and U127 (N_127,In_227,In_392);
and U128 (N_128,In_375,In_74);
or U129 (N_129,In_101,In_72);
or U130 (N_130,In_66,In_23);
or U131 (N_131,In_265,In_436);
nand U132 (N_132,In_480,In_386);
nor U133 (N_133,In_298,In_148);
nor U134 (N_134,In_73,In_444);
or U135 (N_135,In_247,In_39);
and U136 (N_136,In_410,In_204);
nand U137 (N_137,In_138,In_0);
and U138 (N_138,In_326,In_492);
nand U139 (N_139,In_416,In_180);
or U140 (N_140,In_348,In_102);
nor U141 (N_141,In_40,In_486);
nand U142 (N_142,In_317,In_162);
nor U143 (N_143,In_343,In_128);
or U144 (N_144,In_234,In_346);
nor U145 (N_145,In_489,In_127);
and U146 (N_146,In_332,In_342);
and U147 (N_147,In_60,In_6);
nand U148 (N_148,In_9,In_417);
nor U149 (N_149,In_2,In_191);
or U150 (N_150,In_55,In_294);
nand U151 (N_151,In_78,In_351);
and U152 (N_152,In_210,In_350);
nor U153 (N_153,In_225,In_70);
or U154 (N_154,In_499,In_497);
nor U155 (N_155,In_424,In_322);
nor U156 (N_156,In_103,In_297);
and U157 (N_157,In_163,In_217);
and U158 (N_158,In_69,In_295);
nor U159 (N_159,In_64,In_429);
or U160 (N_160,In_50,In_406);
nor U161 (N_161,In_306,In_67);
or U162 (N_162,In_354,In_56);
or U163 (N_163,In_373,In_151);
or U164 (N_164,In_51,In_34);
nor U165 (N_165,In_496,In_455);
or U166 (N_166,In_252,In_330);
nor U167 (N_167,In_432,In_441);
nand U168 (N_168,In_411,In_196);
and U169 (N_169,In_199,In_397);
nand U170 (N_170,In_93,In_44);
or U171 (N_171,In_254,In_361);
nor U172 (N_172,In_405,In_389);
nor U173 (N_173,In_240,In_81);
and U174 (N_174,In_123,In_95);
or U175 (N_175,In_329,In_477);
and U176 (N_176,In_176,In_437);
and U177 (N_177,In_364,In_233);
nand U178 (N_178,In_498,In_229);
and U179 (N_179,In_485,In_259);
nor U180 (N_180,In_46,In_54);
or U181 (N_181,In_4,In_284);
nor U182 (N_182,In_113,In_320);
nor U183 (N_183,In_96,In_464);
nor U184 (N_184,In_232,In_358);
or U185 (N_185,In_16,In_387);
nand U186 (N_186,In_403,In_311);
and U187 (N_187,In_91,In_41);
nor U188 (N_188,In_340,In_344);
and U189 (N_189,In_48,In_134);
nand U190 (N_190,In_28,In_336);
nand U191 (N_191,In_246,In_303);
or U192 (N_192,In_147,In_146);
nand U193 (N_193,In_243,In_137);
nand U194 (N_194,In_142,In_76);
nor U195 (N_195,In_235,In_205);
nand U196 (N_196,In_175,In_143);
and U197 (N_197,In_415,In_129);
nand U198 (N_198,In_474,In_17);
and U199 (N_199,In_494,In_61);
and U200 (N_200,In_250,N_14);
nand U201 (N_201,N_46,N_143);
and U202 (N_202,N_84,In_164);
nor U203 (N_203,N_101,In_242);
nor U204 (N_204,In_106,N_115);
nand U205 (N_205,In_107,N_30);
nand U206 (N_206,In_423,N_156);
and U207 (N_207,N_178,In_458);
nor U208 (N_208,N_90,In_433);
nor U209 (N_209,In_110,N_78);
nor U210 (N_210,In_201,In_149);
or U211 (N_211,N_99,N_50);
nand U212 (N_212,In_248,In_490);
xor U213 (N_213,N_92,In_258);
and U214 (N_214,In_285,N_62);
nor U215 (N_215,N_174,In_111);
or U216 (N_216,In_215,N_11);
or U217 (N_217,In_487,N_120);
and U218 (N_218,N_98,In_226);
nor U219 (N_219,N_144,In_63);
nor U220 (N_220,In_315,N_100);
nor U221 (N_221,N_102,N_121);
nor U222 (N_222,N_44,In_172);
and U223 (N_223,In_376,N_187);
nand U224 (N_224,N_198,N_83);
nor U225 (N_225,N_20,In_57);
and U226 (N_226,In_216,N_199);
and U227 (N_227,N_190,N_97);
and U228 (N_228,In_5,In_97);
or U229 (N_229,N_41,N_103);
and U230 (N_230,N_33,In_177);
or U231 (N_231,In_153,N_189);
or U232 (N_232,In_447,In_174);
nand U233 (N_233,N_35,N_76);
or U234 (N_234,N_162,N_150);
xor U235 (N_235,In_126,N_123);
nand U236 (N_236,In_75,N_81);
nand U237 (N_237,N_141,In_132);
or U238 (N_238,N_166,In_316);
or U239 (N_239,In_65,In_419);
nor U240 (N_240,N_63,N_0);
nor U241 (N_241,N_65,N_155);
nand U242 (N_242,N_9,N_180);
nand U243 (N_243,N_96,N_154);
nand U244 (N_244,In_302,N_127);
nand U245 (N_245,N_8,In_384);
nand U246 (N_246,N_85,N_148);
nor U247 (N_247,N_147,N_136);
or U248 (N_248,N_184,N_59);
or U249 (N_249,N_181,N_47);
or U250 (N_250,In_456,In_394);
or U251 (N_251,N_23,In_29);
or U252 (N_252,N_122,N_4);
and U253 (N_253,N_108,In_273);
and U254 (N_254,N_38,N_93);
and U255 (N_255,N_107,N_43);
and U256 (N_256,In_310,In_296);
nor U257 (N_257,N_48,N_87);
and U258 (N_258,N_188,N_12);
or U259 (N_259,N_28,In_213);
or U260 (N_260,N_6,In_368);
or U261 (N_261,In_189,In_27);
and U262 (N_262,N_70,In_25);
and U263 (N_263,In_383,In_124);
and U264 (N_264,In_202,In_277);
or U265 (N_265,N_168,N_138);
nand U266 (N_266,N_131,N_149);
nand U267 (N_267,In_286,N_146);
nor U268 (N_268,N_36,N_183);
and U269 (N_269,N_128,N_119);
nand U270 (N_270,In_82,N_52);
nor U271 (N_271,N_179,In_198);
nand U272 (N_272,N_194,N_137);
nand U273 (N_273,In_353,N_22);
or U274 (N_274,N_110,In_395);
nor U275 (N_275,In_255,N_130);
and U276 (N_276,N_1,N_32);
and U277 (N_277,N_77,N_54);
nand U278 (N_278,N_134,N_24);
or U279 (N_279,N_151,N_56);
or U280 (N_280,N_18,N_112);
nand U281 (N_281,N_167,N_177);
nand U282 (N_282,N_89,N_152);
nor U283 (N_283,N_49,N_163);
and U284 (N_284,N_71,N_19);
or U285 (N_285,In_349,In_470);
nor U286 (N_286,N_126,N_133);
and U287 (N_287,N_53,In_400);
or U288 (N_288,N_79,N_16);
nand U289 (N_289,In_287,N_27);
nor U290 (N_290,N_2,N_191);
or U291 (N_291,N_171,N_67);
and U292 (N_292,N_64,In_159);
or U293 (N_293,N_34,In_366);
nand U294 (N_294,N_195,In_80);
or U295 (N_295,In_482,In_218);
nand U296 (N_296,N_170,N_109);
nand U297 (N_297,In_467,N_186);
nor U298 (N_298,N_10,N_91);
or U299 (N_299,N_15,N_135);
nor U300 (N_300,N_196,N_55);
nand U301 (N_301,N_192,N_95);
and U302 (N_302,N_42,In_119);
or U303 (N_303,N_153,In_468);
nor U304 (N_304,N_25,N_82);
nand U305 (N_305,N_37,In_283);
nand U306 (N_306,N_69,N_5);
nor U307 (N_307,In_472,N_193);
or U308 (N_308,N_31,N_51);
nand U309 (N_309,N_139,In_145);
or U310 (N_310,In_439,N_173);
and U311 (N_311,In_324,N_172);
nor U312 (N_312,In_367,In_221);
and U313 (N_313,In_465,N_80);
nor U314 (N_314,In_109,N_169);
or U315 (N_315,N_68,In_206);
and U316 (N_316,In_77,In_58);
nand U317 (N_317,N_26,N_113);
nor U318 (N_318,N_13,In_15);
and U319 (N_319,N_165,In_314);
or U320 (N_320,N_39,In_144);
nand U321 (N_321,In_203,N_105);
and U322 (N_322,In_131,N_114);
and U323 (N_323,N_111,N_94);
and U324 (N_324,N_116,N_182);
or U325 (N_325,N_3,N_175);
and U326 (N_326,N_72,N_106);
nor U327 (N_327,N_7,N_88);
or U328 (N_328,N_58,N_21);
or U329 (N_329,N_75,N_158);
or U330 (N_330,N_124,In_228);
and U331 (N_331,N_117,N_86);
nand U332 (N_332,N_60,N_73);
nand U333 (N_333,N_57,N_29);
nand U334 (N_334,N_132,N_197);
and U335 (N_335,N_125,N_185);
nor U336 (N_336,N_159,N_142);
and U337 (N_337,N_45,N_17);
nor U338 (N_338,In_493,N_145);
nor U339 (N_339,N_118,In_182);
nand U340 (N_340,N_160,In_208);
nor U341 (N_341,N_164,N_74);
and U342 (N_342,In_30,N_161);
and U343 (N_343,In_453,N_66);
nand U344 (N_344,N_104,N_140);
nor U345 (N_345,N_157,In_337);
or U346 (N_346,In_312,In_300);
nor U347 (N_347,N_40,N_61);
and U348 (N_348,In_268,In_279);
nand U349 (N_349,N_176,N_129);
nand U350 (N_350,In_250,In_149);
or U351 (N_351,N_85,N_189);
nand U352 (N_352,N_65,In_215);
nor U353 (N_353,N_93,N_128);
and U354 (N_354,N_67,N_83);
and U355 (N_355,N_61,N_2);
and U356 (N_356,N_107,N_72);
or U357 (N_357,N_118,N_14);
and U358 (N_358,N_184,N_45);
nor U359 (N_359,N_82,N_196);
and U360 (N_360,N_62,N_69);
or U361 (N_361,N_2,In_97);
nand U362 (N_362,In_470,N_42);
nor U363 (N_363,N_161,N_182);
or U364 (N_364,N_147,N_6);
or U365 (N_365,N_55,In_216);
nand U366 (N_366,In_172,N_140);
and U367 (N_367,N_197,In_423);
and U368 (N_368,N_79,N_28);
and U369 (N_369,N_76,N_176);
or U370 (N_370,In_65,In_493);
and U371 (N_371,N_160,In_472);
nand U372 (N_372,In_255,N_198);
nand U373 (N_373,N_49,In_80);
nor U374 (N_374,In_470,N_180);
or U375 (N_375,N_63,N_110);
nand U376 (N_376,In_433,N_105);
nand U377 (N_377,N_58,N_91);
nand U378 (N_378,N_150,N_106);
nor U379 (N_379,N_169,In_153);
or U380 (N_380,N_176,In_353);
or U381 (N_381,N_93,In_400);
or U382 (N_382,N_32,In_177);
or U383 (N_383,N_186,N_199);
nand U384 (N_384,In_453,In_470);
and U385 (N_385,N_97,In_124);
nand U386 (N_386,In_423,N_88);
nand U387 (N_387,In_302,In_472);
nand U388 (N_388,N_120,N_133);
and U389 (N_389,N_75,N_128);
nand U390 (N_390,In_456,In_131);
nand U391 (N_391,In_285,N_50);
nand U392 (N_392,N_52,In_218);
nand U393 (N_393,N_45,N_23);
nand U394 (N_394,N_129,N_184);
nor U395 (N_395,In_349,N_176);
nand U396 (N_396,N_59,N_75);
and U397 (N_397,N_108,In_286);
nand U398 (N_398,N_17,N_197);
nand U399 (N_399,N_131,N_12);
and U400 (N_400,N_340,N_284);
nor U401 (N_401,N_258,N_399);
nand U402 (N_402,N_275,N_252);
and U403 (N_403,N_280,N_323);
and U404 (N_404,N_299,N_298);
and U405 (N_405,N_362,N_350);
nor U406 (N_406,N_364,N_259);
nand U407 (N_407,N_303,N_244);
nor U408 (N_408,N_234,N_334);
or U409 (N_409,N_328,N_349);
nor U410 (N_410,N_333,N_365);
nor U411 (N_411,N_326,N_344);
and U412 (N_412,N_287,N_216);
or U413 (N_413,N_207,N_373);
nor U414 (N_414,N_354,N_255);
or U415 (N_415,N_290,N_223);
nor U416 (N_416,N_208,N_210);
or U417 (N_417,N_225,N_227);
nor U418 (N_418,N_308,N_200);
nor U419 (N_419,N_337,N_268);
nand U420 (N_420,N_397,N_236);
nor U421 (N_421,N_237,N_246);
nand U422 (N_422,N_204,N_209);
and U423 (N_423,N_243,N_359);
nor U424 (N_424,N_331,N_267);
or U425 (N_425,N_294,N_296);
nand U426 (N_426,N_222,N_379);
or U427 (N_427,N_261,N_235);
nor U428 (N_428,N_322,N_324);
and U429 (N_429,N_387,N_274);
or U430 (N_430,N_249,N_277);
nor U431 (N_431,N_272,N_218);
and U432 (N_432,N_355,N_247);
nor U433 (N_433,N_229,N_394);
and U434 (N_434,N_219,N_366);
nor U435 (N_435,N_297,N_378);
or U436 (N_436,N_314,N_313);
nand U437 (N_437,N_319,N_385);
or U438 (N_438,N_302,N_241);
or U439 (N_439,N_266,N_220);
or U440 (N_440,N_346,N_339);
nor U441 (N_441,N_372,N_206);
or U442 (N_442,N_292,N_276);
or U443 (N_443,N_291,N_264);
and U444 (N_444,N_392,N_332);
nor U445 (N_445,N_257,N_383);
or U446 (N_446,N_305,N_317);
and U447 (N_447,N_212,N_369);
nor U448 (N_448,N_254,N_321);
and U449 (N_449,N_232,N_384);
nor U450 (N_450,N_293,N_233);
nand U451 (N_451,N_318,N_370);
and U452 (N_452,N_380,N_320);
nor U453 (N_453,N_300,N_398);
or U454 (N_454,N_338,N_221);
or U455 (N_455,N_203,N_368);
or U456 (N_456,N_304,N_310);
and U457 (N_457,N_329,N_393);
nand U458 (N_458,N_390,N_341);
or U459 (N_459,N_361,N_285);
and U460 (N_460,N_226,N_357);
or U461 (N_461,N_214,N_283);
and U462 (N_462,N_377,N_396);
nand U463 (N_463,N_381,N_217);
nand U464 (N_464,N_262,N_248);
nor U465 (N_465,N_391,N_279);
or U466 (N_466,N_386,N_289);
or U467 (N_467,N_260,N_351);
and U468 (N_468,N_240,N_309);
or U469 (N_469,N_376,N_315);
and U470 (N_470,N_202,N_327);
nand U471 (N_471,N_271,N_231);
and U472 (N_472,N_213,N_374);
or U473 (N_473,N_363,N_281);
nand U474 (N_474,N_356,N_360);
and U475 (N_475,N_306,N_224);
nor U476 (N_476,N_345,N_336);
nor U477 (N_477,N_253,N_311);
nand U478 (N_478,N_270,N_388);
and U479 (N_479,N_316,N_286);
and U480 (N_480,N_251,N_278);
and U481 (N_481,N_295,N_375);
nor U482 (N_482,N_211,N_307);
nor U483 (N_483,N_215,N_312);
nand U484 (N_484,N_205,N_238);
nor U485 (N_485,N_325,N_371);
nand U486 (N_486,N_395,N_353);
or U487 (N_487,N_352,N_342);
xnor U488 (N_488,N_358,N_343);
or U489 (N_489,N_273,N_242);
and U490 (N_490,N_288,N_201);
nand U491 (N_491,N_263,N_256);
or U492 (N_492,N_282,N_269);
or U493 (N_493,N_230,N_301);
or U494 (N_494,N_330,N_335);
nor U495 (N_495,N_389,N_239);
nor U496 (N_496,N_382,N_245);
nor U497 (N_497,N_367,N_228);
and U498 (N_498,N_347,N_265);
nand U499 (N_499,N_250,N_348);
nor U500 (N_500,N_302,N_265);
nor U501 (N_501,N_245,N_385);
or U502 (N_502,N_202,N_342);
and U503 (N_503,N_295,N_258);
and U504 (N_504,N_268,N_211);
nand U505 (N_505,N_357,N_333);
or U506 (N_506,N_377,N_307);
nand U507 (N_507,N_268,N_295);
or U508 (N_508,N_377,N_261);
xor U509 (N_509,N_209,N_276);
nand U510 (N_510,N_393,N_388);
nand U511 (N_511,N_377,N_244);
nand U512 (N_512,N_262,N_272);
and U513 (N_513,N_329,N_300);
nand U514 (N_514,N_374,N_365);
and U515 (N_515,N_293,N_230);
nand U516 (N_516,N_247,N_368);
xor U517 (N_517,N_258,N_382);
and U518 (N_518,N_263,N_364);
or U519 (N_519,N_201,N_298);
or U520 (N_520,N_317,N_296);
or U521 (N_521,N_349,N_297);
xnor U522 (N_522,N_208,N_268);
nor U523 (N_523,N_229,N_338);
and U524 (N_524,N_262,N_252);
or U525 (N_525,N_378,N_392);
nand U526 (N_526,N_237,N_290);
or U527 (N_527,N_294,N_320);
and U528 (N_528,N_214,N_398);
or U529 (N_529,N_348,N_279);
or U530 (N_530,N_203,N_235);
nand U531 (N_531,N_240,N_363);
nor U532 (N_532,N_283,N_355);
nor U533 (N_533,N_329,N_232);
and U534 (N_534,N_310,N_356);
and U535 (N_535,N_233,N_229);
and U536 (N_536,N_376,N_359);
nor U537 (N_537,N_270,N_273);
nor U538 (N_538,N_348,N_258);
and U539 (N_539,N_382,N_276);
nand U540 (N_540,N_219,N_265);
nand U541 (N_541,N_347,N_388);
nor U542 (N_542,N_266,N_268);
nand U543 (N_543,N_279,N_323);
and U544 (N_544,N_281,N_301);
nand U545 (N_545,N_288,N_381);
nand U546 (N_546,N_241,N_380);
and U547 (N_547,N_304,N_293);
and U548 (N_548,N_264,N_259);
nor U549 (N_549,N_267,N_207);
and U550 (N_550,N_372,N_290);
or U551 (N_551,N_245,N_327);
or U552 (N_552,N_372,N_213);
nand U553 (N_553,N_313,N_232);
nor U554 (N_554,N_338,N_396);
nand U555 (N_555,N_265,N_226);
and U556 (N_556,N_317,N_287);
nor U557 (N_557,N_398,N_289);
or U558 (N_558,N_309,N_229);
and U559 (N_559,N_341,N_392);
nor U560 (N_560,N_207,N_332);
and U561 (N_561,N_348,N_204);
nand U562 (N_562,N_344,N_318);
or U563 (N_563,N_372,N_356);
nor U564 (N_564,N_322,N_213);
or U565 (N_565,N_251,N_271);
or U566 (N_566,N_260,N_281);
and U567 (N_567,N_307,N_339);
nor U568 (N_568,N_389,N_205);
and U569 (N_569,N_380,N_222);
nand U570 (N_570,N_246,N_228);
or U571 (N_571,N_384,N_250);
nor U572 (N_572,N_280,N_306);
nand U573 (N_573,N_240,N_368);
nand U574 (N_574,N_244,N_299);
or U575 (N_575,N_381,N_388);
nor U576 (N_576,N_258,N_224);
nand U577 (N_577,N_314,N_381);
nand U578 (N_578,N_333,N_262);
nand U579 (N_579,N_293,N_312);
or U580 (N_580,N_247,N_397);
or U581 (N_581,N_371,N_329);
nor U582 (N_582,N_306,N_391);
nor U583 (N_583,N_314,N_351);
nand U584 (N_584,N_246,N_342);
and U585 (N_585,N_212,N_398);
nor U586 (N_586,N_279,N_398);
nand U587 (N_587,N_237,N_242);
nor U588 (N_588,N_333,N_256);
nand U589 (N_589,N_207,N_396);
and U590 (N_590,N_261,N_325);
or U591 (N_591,N_251,N_252);
nor U592 (N_592,N_362,N_351);
and U593 (N_593,N_301,N_237);
xor U594 (N_594,N_357,N_243);
or U595 (N_595,N_287,N_347);
or U596 (N_596,N_260,N_314);
nor U597 (N_597,N_317,N_208);
or U598 (N_598,N_334,N_216);
nand U599 (N_599,N_293,N_366);
nor U600 (N_600,N_437,N_451);
and U601 (N_601,N_421,N_588);
nand U602 (N_602,N_449,N_491);
and U603 (N_603,N_501,N_484);
nor U604 (N_604,N_567,N_568);
and U605 (N_605,N_429,N_573);
and U606 (N_606,N_518,N_438);
and U607 (N_607,N_494,N_507);
nor U608 (N_608,N_516,N_550);
nor U609 (N_609,N_462,N_452);
and U610 (N_610,N_548,N_478);
or U611 (N_611,N_475,N_461);
and U612 (N_612,N_570,N_579);
and U613 (N_613,N_436,N_569);
and U614 (N_614,N_416,N_598);
xor U615 (N_615,N_497,N_464);
nor U616 (N_616,N_595,N_422);
or U617 (N_617,N_407,N_537);
and U618 (N_618,N_492,N_534);
and U619 (N_619,N_456,N_420);
nand U620 (N_620,N_417,N_405);
nand U621 (N_621,N_559,N_561);
and U622 (N_622,N_474,N_447);
and U623 (N_623,N_535,N_586);
nor U624 (N_624,N_508,N_528);
nor U625 (N_625,N_571,N_448);
or U626 (N_626,N_521,N_582);
nand U627 (N_627,N_546,N_425);
or U628 (N_628,N_587,N_412);
nand U629 (N_629,N_583,N_434);
or U630 (N_630,N_402,N_409);
nor U631 (N_631,N_498,N_514);
or U632 (N_632,N_444,N_431);
or U633 (N_633,N_538,N_556);
and U634 (N_634,N_496,N_504);
or U635 (N_635,N_511,N_515);
and U636 (N_636,N_530,N_581);
or U637 (N_637,N_499,N_467);
or U638 (N_638,N_460,N_472);
nand U639 (N_639,N_566,N_589);
and U640 (N_640,N_541,N_562);
or U641 (N_641,N_505,N_560);
or U642 (N_642,N_572,N_458);
nand U643 (N_643,N_533,N_432);
nand U644 (N_644,N_457,N_552);
or U645 (N_645,N_590,N_476);
nor U646 (N_646,N_591,N_424);
or U647 (N_647,N_563,N_413);
and U648 (N_648,N_418,N_427);
and U649 (N_649,N_465,N_482);
or U650 (N_650,N_426,N_488);
nand U651 (N_651,N_578,N_489);
and U652 (N_652,N_529,N_593);
or U653 (N_653,N_439,N_525);
and U654 (N_654,N_400,N_596);
or U655 (N_655,N_404,N_487);
and U656 (N_656,N_410,N_543);
and U657 (N_657,N_473,N_428);
nor U658 (N_658,N_446,N_554);
or U659 (N_659,N_527,N_577);
nand U660 (N_660,N_553,N_479);
nand U661 (N_661,N_502,N_544);
or U662 (N_662,N_558,N_463);
and U663 (N_663,N_403,N_443);
nand U664 (N_664,N_584,N_406);
or U665 (N_665,N_539,N_423);
nor U666 (N_666,N_470,N_574);
and U667 (N_667,N_549,N_592);
nor U668 (N_668,N_408,N_455);
or U669 (N_669,N_526,N_555);
and U670 (N_670,N_414,N_551);
or U671 (N_671,N_520,N_468);
and U672 (N_672,N_480,N_440);
nor U673 (N_673,N_450,N_401);
nand U674 (N_674,N_540,N_441);
nor U675 (N_675,N_599,N_481);
or U676 (N_676,N_575,N_459);
and U677 (N_677,N_486,N_564);
nand U678 (N_678,N_415,N_454);
or U679 (N_679,N_597,N_509);
and U680 (N_680,N_411,N_419);
nand U681 (N_681,N_477,N_585);
nor U682 (N_682,N_485,N_576);
or U683 (N_683,N_469,N_517);
xor U684 (N_684,N_506,N_500);
and U685 (N_685,N_557,N_493);
nand U686 (N_686,N_495,N_580);
and U687 (N_687,N_519,N_453);
or U688 (N_688,N_433,N_483);
and U689 (N_689,N_442,N_532);
and U690 (N_690,N_490,N_545);
and U691 (N_691,N_524,N_565);
nor U692 (N_692,N_542,N_522);
nor U693 (N_693,N_510,N_503);
or U694 (N_694,N_512,N_594);
or U695 (N_695,N_531,N_547);
and U696 (N_696,N_523,N_430);
and U697 (N_697,N_513,N_466);
nor U698 (N_698,N_445,N_536);
nor U699 (N_699,N_435,N_471);
and U700 (N_700,N_444,N_568);
or U701 (N_701,N_410,N_508);
and U702 (N_702,N_467,N_460);
and U703 (N_703,N_412,N_568);
or U704 (N_704,N_485,N_509);
or U705 (N_705,N_491,N_584);
and U706 (N_706,N_430,N_589);
and U707 (N_707,N_557,N_433);
nor U708 (N_708,N_452,N_514);
nand U709 (N_709,N_535,N_510);
nor U710 (N_710,N_471,N_400);
nor U711 (N_711,N_500,N_561);
nor U712 (N_712,N_449,N_585);
and U713 (N_713,N_446,N_512);
or U714 (N_714,N_565,N_555);
nand U715 (N_715,N_592,N_505);
nor U716 (N_716,N_436,N_529);
nand U717 (N_717,N_574,N_543);
xnor U718 (N_718,N_592,N_485);
and U719 (N_719,N_549,N_562);
nor U720 (N_720,N_510,N_579);
nand U721 (N_721,N_406,N_417);
nand U722 (N_722,N_457,N_487);
xor U723 (N_723,N_496,N_511);
and U724 (N_724,N_580,N_589);
or U725 (N_725,N_429,N_436);
nor U726 (N_726,N_462,N_523);
nand U727 (N_727,N_426,N_588);
xor U728 (N_728,N_521,N_549);
nand U729 (N_729,N_472,N_594);
or U730 (N_730,N_525,N_543);
nor U731 (N_731,N_550,N_498);
nor U732 (N_732,N_471,N_437);
nand U733 (N_733,N_539,N_430);
or U734 (N_734,N_514,N_524);
and U735 (N_735,N_427,N_471);
nand U736 (N_736,N_482,N_467);
and U737 (N_737,N_516,N_499);
or U738 (N_738,N_423,N_491);
and U739 (N_739,N_569,N_595);
or U740 (N_740,N_561,N_405);
and U741 (N_741,N_531,N_508);
and U742 (N_742,N_555,N_434);
nand U743 (N_743,N_581,N_520);
or U744 (N_744,N_587,N_509);
nand U745 (N_745,N_468,N_548);
nand U746 (N_746,N_474,N_599);
and U747 (N_747,N_475,N_480);
and U748 (N_748,N_568,N_507);
xnor U749 (N_749,N_451,N_536);
nor U750 (N_750,N_479,N_556);
and U751 (N_751,N_559,N_469);
nand U752 (N_752,N_466,N_441);
and U753 (N_753,N_424,N_471);
nor U754 (N_754,N_514,N_446);
nor U755 (N_755,N_444,N_450);
and U756 (N_756,N_582,N_528);
xnor U757 (N_757,N_563,N_568);
or U758 (N_758,N_562,N_479);
and U759 (N_759,N_491,N_526);
nand U760 (N_760,N_489,N_440);
and U761 (N_761,N_400,N_572);
nand U762 (N_762,N_573,N_474);
nor U763 (N_763,N_421,N_519);
nor U764 (N_764,N_521,N_496);
and U765 (N_765,N_488,N_482);
nor U766 (N_766,N_528,N_570);
and U767 (N_767,N_402,N_561);
or U768 (N_768,N_456,N_540);
or U769 (N_769,N_561,N_550);
nand U770 (N_770,N_458,N_585);
nor U771 (N_771,N_533,N_486);
or U772 (N_772,N_485,N_409);
or U773 (N_773,N_443,N_576);
or U774 (N_774,N_493,N_495);
nand U775 (N_775,N_400,N_436);
and U776 (N_776,N_531,N_589);
and U777 (N_777,N_437,N_492);
nor U778 (N_778,N_444,N_449);
xnor U779 (N_779,N_526,N_505);
nand U780 (N_780,N_515,N_596);
nand U781 (N_781,N_468,N_446);
nand U782 (N_782,N_438,N_464);
nor U783 (N_783,N_532,N_538);
and U784 (N_784,N_477,N_485);
or U785 (N_785,N_522,N_475);
nor U786 (N_786,N_506,N_534);
or U787 (N_787,N_533,N_574);
and U788 (N_788,N_541,N_599);
or U789 (N_789,N_473,N_515);
or U790 (N_790,N_563,N_507);
nand U791 (N_791,N_548,N_444);
nor U792 (N_792,N_578,N_576);
and U793 (N_793,N_573,N_581);
or U794 (N_794,N_509,N_503);
nand U795 (N_795,N_495,N_497);
xor U796 (N_796,N_586,N_461);
nand U797 (N_797,N_422,N_597);
nor U798 (N_798,N_466,N_475);
or U799 (N_799,N_457,N_522);
nand U800 (N_800,N_668,N_641);
or U801 (N_801,N_644,N_712);
nor U802 (N_802,N_687,N_773);
and U803 (N_803,N_669,N_629);
nand U804 (N_804,N_661,N_701);
and U805 (N_805,N_610,N_720);
and U806 (N_806,N_672,N_797);
nor U807 (N_807,N_649,N_748);
nor U808 (N_808,N_702,N_774);
and U809 (N_809,N_777,N_628);
nor U810 (N_810,N_783,N_731);
nand U811 (N_811,N_686,N_634);
nor U812 (N_812,N_654,N_733);
and U813 (N_813,N_689,N_758);
nor U814 (N_814,N_751,N_630);
and U815 (N_815,N_770,N_618);
nand U816 (N_816,N_767,N_694);
nor U817 (N_817,N_740,N_625);
and U818 (N_818,N_724,N_747);
nor U819 (N_819,N_743,N_650);
nand U820 (N_820,N_648,N_678);
nor U821 (N_821,N_787,N_732);
nand U822 (N_822,N_713,N_780);
nand U823 (N_823,N_744,N_667);
nand U824 (N_824,N_789,N_734);
or U825 (N_825,N_652,N_794);
nand U826 (N_826,N_616,N_710);
and U827 (N_827,N_736,N_635);
nand U828 (N_828,N_714,N_742);
nor U829 (N_829,N_674,N_764);
nand U830 (N_830,N_754,N_623);
and U831 (N_831,N_706,N_603);
nand U832 (N_832,N_752,N_760);
and U833 (N_833,N_798,N_725);
and U834 (N_834,N_624,N_782);
and U835 (N_835,N_658,N_703);
nor U836 (N_836,N_788,N_757);
nor U837 (N_837,N_643,N_699);
or U838 (N_838,N_612,N_671);
or U839 (N_839,N_682,N_716);
or U840 (N_840,N_642,N_781);
or U841 (N_841,N_670,N_615);
and U842 (N_842,N_721,N_684);
nand U843 (N_843,N_775,N_795);
and U844 (N_844,N_659,N_605);
and U845 (N_845,N_756,N_651);
and U846 (N_846,N_768,N_704);
nand U847 (N_847,N_680,N_692);
or U848 (N_848,N_719,N_750);
nand U849 (N_849,N_664,N_614);
nor U850 (N_850,N_785,N_679);
nand U851 (N_851,N_685,N_639);
and U852 (N_852,N_791,N_741);
nand U853 (N_853,N_620,N_691);
and U854 (N_854,N_695,N_793);
and U855 (N_855,N_772,N_613);
nor U856 (N_856,N_753,N_778);
and U857 (N_857,N_640,N_681);
and U858 (N_858,N_796,N_727);
and U859 (N_859,N_677,N_786);
or U860 (N_860,N_601,N_609);
and U861 (N_861,N_604,N_662);
nor U862 (N_862,N_700,N_745);
nand U863 (N_863,N_632,N_715);
nor U864 (N_864,N_693,N_707);
and U865 (N_865,N_600,N_645);
or U866 (N_866,N_763,N_607);
or U867 (N_867,N_738,N_647);
nor U868 (N_868,N_749,N_737);
nand U869 (N_869,N_755,N_606);
nor U870 (N_870,N_759,N_735);
and U871 (N_871,N_697,N_790);
and U872 (N_872,N_711,N_638);
nor U873 (N_873,N_784,N_688);
and U874 (N_874,N_769,N_728);
and U875 (N_875,N_602,N_766);
or U876 (N_876,N_799,N_726);
nand U877 (N_877,N_617,N_666);
or U878 (N_878,N_771,N_653);
nor U879 (N_879,N_730,N_637);
or U880 (N_880,N_646,N_673);
nand U881 (N_881,N_729,N_657);
nand U882 (N_882,N_675,N_631);
nor U883 (N_883,N_705,N_636);
nand U884 (N_884,N_792,N_676);
xnor U885 (N_885,N_665,N_739);
or U886 (N_886,N_746,N_708);
nand U887 (N_887,N_762,N_655);
or U888 (N_888,N_656,N_765);
nand U889 (N_889,N_621,N_690);
nor U890 (N_890,N_608,N_718);
and U891 (N_891,N_663,N_619);
and U892 (N_892,N_698,N_696);
nor U893 (N_893,N_723,N_779);
nand U894 (N_894,N_709,N_611);
and U895 (N_895,N_683,N_622);
or U896 (N_896,N_627,N_722);
or U897 (N_897,N_660,N_717);
or U898 (N_898,N_776,N_761);
nand U899 (N_899,N_633,N_626);
or U900 (N_900,N_684,N_640);
nand U901 (N_901,N_774,N_620);
or U902 (N_902,N_754,N_784);
nor U903 (N_903,N_640,N_611);
nand U904 (N_904,N_675,N_719);
nand U905 (N_905,N_666,N_628);
and U906 (N_906,N_768,N_754);
and U907 (N_907,N_726,N_791);
nor U908 (N_908,N_693,N_630);
and U909 (N_909,N_632,N_762);
or U910 (N_910,N_722,N_686);
nor U911 (N_911,N_711,N_712);
nor U912 (N_912,N_622,N_650);
nand U913 (N_913,N_622,N_728);
nand U914 (N_914,N_638,N_745);
nand U915 (N_915,N_625,N_687);
nand U916 (N_916,N_727,N_695);
or U917 (N_917,N_759,N_610);
and U918 (N_918,N_736,N_653);
nor U919 (N_919,N_707,N_673);
nand U920 (N_920,N_604,N_602);
nor U921 (N_921,N_738,N_645);
nor U922 (N_922,N_687,N_782);
or U923 (N_923,N_607,N_693);
and U924 (N_924,N_720,N_679);
nand U925 (N_925,N_666,N_694);
nand U926 (N_926,N_744,N_722);
nand U927 (N_927,N_629,N_700);
nand U928 (N_928,N_621,N_671);
nor U929 (N_929,N_671,N_625);
or U930 (N_930,N_778,N_662);
and U931 (N_931,N_659,N_761);
nand U932 (N_932,N_746,N_713);
or U933 (N_933,N_773,N_749);
or U934 (N_934,N_621,N_606);
or U935 (N_935,N_626,N_661);
and U936 (N_936,N_754,N_781);
and U937 (N_937,N_781,N_728);
nand U938 (N_938,N_709,N_635);
nor U939 (N_939,N_650,N_684);
or U940 (N_940,N_740,N_762);
nand U941 (N_941,N_620,N_697);
nand U942 (N_942,N_635,N_795);
nor U943 (N_943,N_658,N_632);
nor U944 (N_944,N_653,N_764);
nand U945 (N_945,N_619,N_609);
or U946 (N_946,N_701,N_664);
or U947 (N_947,N_615,N_684);
and U948 (N_948,N_769,N_714);
nor U949 (N_949,N_773,N_748);
or U950 (N_950,N_744,N_605);
and U951 (N_951,N_684,N_636);
and U952 (N_952,N_659,N_635);
and U953 (N_953,N_758,N_631);
xor U954 (N_954,N_771,N_742);
or U955 (N_955,N_704,N_710);
nand U956 (N_956,N_787,N_600);
and U957 (N_957,N_601,N_781);
nand U958 (N_958,N_702,N_626);
nand U959 (N_959,N_724,N_602);
or U960 (N_960,N_711,N_786);
nor U961 (N_961,N_743,N_645);
nand U962 (N_962,N_660,N_621);
and U963 (N_963,N_734,N_674);
nand U964 (N_964,N_693,N_675);
nor U965 (N_965,N_729,N_772);
nand U966 (N_966,N_715,N_699);
or U967 (N_967,N_781,N_623);
nor U968 (N_968,N_799,N_703);
nor U969 (N_969,N_753,N_726);
nand U970 (N_970,N_799,N_621);
nand U971 (N_971,N_672,N_703);
and U972 (N_972,N_602,N_705);
and U973 (N_973,N_794,N_691);
or U974 (N_974,N_650,N_635);
or U975 (N_975,N_678,N_726);
and U976 (N_976,N_725,N_686);
and U977 (N_977,N_616,N_670);
or U978 (N_978,N_746,N_611);
and U979 (N_979,N_757,N_659);
and U980 (N_980,N_749,N_668);
or U981 (N_981,N_689,N_682);
nor U982 (N_982,N_644,N_785);
xor U983 (N_983,N_639,N_740);
and U984 (N_984,N_718,N_696);
nand U985 (N_985,N_751,N_794);
nor U986 (N_986,N_777,N_629);
nor U987 (N_987,N_643,N_600);
or U988 (N_988,N_703,N_685);
or U989 (N_989,N_626,N_674);
nand U990 (N_990,N_615,N_673);
and U991 (N_991,N_693,N_618);
nand U992 (N_992,N_648,N_685);
or U993 (N_993,N_630,N_632);
and U994 (N_994,N_744,N_779);
and U995 (N_995,N_756,N_797);
or U996 (N_996,N_659,N_636);
and U997 (N_997,N_621,N_744);
and U998 (N_998,N_714,N_627);
and U999 (N_999,N_702,N_728);
and U1000 (N_1000,N_958,N_802);
and U1001 (N_1001,N_920,N_936);
nor U1002 (N_1002,N_971,N_948);
nand U1003 (N_1003,N_821,N_883);
or U1004 (N_1004,N_912,N_914);
nand U1005 (N_1005,N_988,N_878);
and U1006 (N_1006,N_855,N_831);
nand U1007 (N_1007,N_982,N_856);
xnor U1008 (N_1008,N_853,N_818);
nor U1009 (N_1009,N_946,N_979);
or U1010 (N_1010,N_808,N_842);
nand U1011 (N_1011,N_800,N_973);
nor U1012 (N_1012,N_823,N_944);
and U1013 (N_1013,N_943,N_811);
xor U1014 (N_1014,N_891,N_886);
nand U1015 (N_1015,N_838,N_935);
nand U1016 (N_1016,N_919,N_922);
and U1017 (N_1017,N_933,N_969);
nor U1018 (N_1018,N_926,N_862);
or U1019 (N_1019,N_816,N_807);
nor U1020 (N_1020,N_999,N_998);
or U1021 (N_1021,N_848,N_830);
nand U1022 (N_1022,N_810,N_822);
and U1023 (N_1023,N_897,N_834);
nor U1024 (N_1024,N_918,N_825);
nand U1025 (N_1025,N_903,N_869);
nor U1026 (N_1026,N_877,N_980);
nor U1027 (N_1027,N_925,N_941);
and U1028 (N_1028,N_904,N_937);
nand U1029 (N_1029,N_962,N_801);
nor U1030 (N_1030,N_993,N_892);
and U1031 (N_1031,N_870,N_956);
nand U1032 (N_1032,N_910,N_985);
nor U1033 (N_1033,N_876,N_945);
nor U1034 (N_1034,N_879,N_929);
and U1035 (N_1035,N_888,N_916);
and U1036 (N_1036,N_970,N_826);
nand U1037 (N_1037,N_898,N_986);
nand U1038 (N_1038,N_871,N_815);
or U1039 (N_1039,N_865,N_857);
or U1040 (N_1040,N_867,N_809);
or U1041 (N_1041,N_952,N_851);
and U1042 (N_1042,N_872,N_806);
nand U1043 (N_1043,N_875,N_906);
nor U1044 (N_1044,N_968,N_913);
and U1045 (N_1045,N_817,N_899);
or U1046 (N_1046,N_804,N_894);
and U1047 (N_1047,N_832,N_928);
or U1048 (N_1048,N_896,N_957);
nand U1049 (N_1049,N_964,N_864);
nor U1050 (N_1050,N_835,N_847);
or U1051 (N_1051,N_953,N_880);
nor U1052 (N_1052,N_874,N_967);
and U1053 (N_1053,N_893,N_976);
nand U1054 (N_1054,N_991,N_997);
and U1055 (N_1055,N_887,N_917);
or U1056 (N_1056,N_931,N_949);
nor U1057 (N_1057,N_930,N_989);
and U1058 (N_1058,N_939,N_965);
and U1059 (N_1059,N_955,N_824);
nand U1060 (N_1060,N_996,N_981);
nor U1061 (N_1061,N_895,N_961);
nor U1062 (N_1062,N_960,N_995);
or U1063 (N_1063,N_947,N_905);
nor U1064 (N_1064,N_923,N_849);
nand U1065 (N_1065,N_889,N_940);
nor U1066 (N_1066,N_908,N_977);
and U1067 (N_1067,N_854,N_846);
or U1068 (N_1068,N_805,N_843);
nand U1069 (N_1069,N_839,N_963);
nand U1070 (N_1070,N_978,N_959);
and U1071 (N_1071,N_833,N_924);
or U1072 (N_1072,N_966,N_882);
or U1073 (N_1073,N_860,N_840);
and U1074 (N_1074,N_927,N_829);
and U1075 (N_1075,N_820,N_902);
or U1076 (N_1076,N_915,N_828);
or U1077 (N_1077,N_950,N_858);
or U1078 (N_1078,N_866,N_992);
nor U1079 (N_1079,N_827,N_881);
nor U1080 (N_1080,N_994,N_850);
or U1081 (N_1081,N_974,N_934);
nor U1082 (N_1082,N_907,N_911);
nor U1083 (N_1083,N_814,N_885);
nand U1084 (N_1084,N_863,N_884);
nand U1085 (N_1085,N_972,N_812);
or U1086 (N_1086,N_951,N_819);
nand U1087 (N_1087,N_890,N_901);
and U1088 (N_1088,N_844,N_987);
and U1089 (N_1089,N_942,N_861);
and U1090 (N_1090,N_984,N_900);
nor U1091 (N_1091,N_852,N_836);
or U1092 (N_1092,N_845,N_837);
nor U1093 (N_1093,N_859,N_975);
and U1094 (N_1094,N_868,N_932);
and U1095 (N_1095,N_873,N_841);
nand U1096 (N_1096,N_909,N_803);
and U1097 (N_1097,N_983,N_921);
or U1098 (N_1098,N_813,N_954);
and U1099 (N_1099,N_990,N_938);
and U1100 (N_1100,N_822,N_828);
nor U1101 (N_1101,N_806,N_971);
nor U1102 (N_1102,N_804,N_837);
and U1103 (N_1103,N_987,N_877);
and U1104 (N_1104,N_846,N_880);
or U1105 (N_1105,N_811,N_853);
nor U1106 (N_1106,N_934,N_918);
nand U1107 (N_1107,N_937,N_947);
and U1108 (N_1108,N_904,N_836);
nand U1109 (N_1109,N_940,N_941);
and U1110 (N_1110,N_867,N_983);
or U1111 (N_1111,N_981,N_924);
nor U1112 (N_1112,N_851,N_905);
nor U1113 (N_1113,N_910,N_918);
and U1114 (N_1114,N_826,N_886);
nor U1115 (N_1115,N_983,N_952);
or U1116 (N_1116,N_923,N_865);
nand U1117 (N_1117,N_905,N_840);
nor U1118 (N_1118,N_977,N_925);
nand U1119 (N_1119,N_998,N_806);
nand U1120 (N_1120,N_910,N_877);
xnor U1121 (N_1121,N_890,N_871);
nand U1122 (N_1122,N_818,N_878);
and U1123 (N_1123,N_896,N_982);
xnor U1124 (N_1124,N_913,N_818);
nand U1125 (N_1125,N_889,N_865);
or U1126 (N_1126,N_910,N_814);
and U1127 (N_1127,N_952,N_999);
nor U1128 (N_1128,N_905,N_854);
and U1129 (N_1129,N_896,N_824);
and U1130 (N_1130,N_810,N_981);
or U1131 (N_1131,N_859,N_800);
nand U1132 (N_1132,N_851,N_808);
and U1133 (N_1133,N_949,N_942);
nand U1134 (N_1134,N_867,N_918);
nor U1135 (N_1135,N_935,N_842);
xor U1136 (N_1136,N_991,N_934);
or U1137 (N_1137,N_946,N_885);
nor U1138 (N_1138,N_999,N_927);
and U1139 (N_1139,N_959,N_997);
and U1140 (N_1140,N_969,N_900);
nand U1141 (N_1141,N_916,N_838);
or U1142 (N_1142,N_905,N_843);
and U1143 (N_1143,N_953,N_936);
or U1144 (N_1144,N_868,N_873);
nand U1145 (N_1145,N_848,N_996);
and U1146 (N_1146,N_866,N_831);
or U1147 (N_1147,N_948,N_918);
nand U1148 (N_1148,N_831,N_847);
and U1149 (N_1149,N_830,N_865);
or U1150 (N_1150,N_982,N_909);
or U1151 (N_1151,N_963,N_934);
nand U1152 (N_1152,N_927,N_897);
or U1153 (N_1153,N_961,N_834);
nand U1154 (N_1154,N_956,N_998);
nand U1155 (N_1155,N_940,N_964);
or U1156 (N_1156,N_873,N_837);
or U1157 (N_1157,N_878,N_846);
or U1158 (N_1158,N_831,N_807);
or U1159 (N_1159,N_985,N_849);
nand U1160 (N_1160,N_847,N_925);
or U1161 (N_1161,N_936,N_855);
and U1162 (N_1162,N_925,N_860);
and U1163 (N_1163,N_908,N_924);
nor U1164 (N_1164,N_977,N_916);
and U1165 (N_1165,N_837,N_974);
nand U1166 (N_1166,N_939,N_823);
nand U1167 (N_1167,N_947,N_810);
and U1168 (N_1168,N_899,N_978);
nor U1169 (N_1169,N_919,N_913);
or U1170 (N_1170,N_811,N_904);
nand U1171 (N_1171,N_997,N_972);
or U1172 (N_1172,N_837,N_863);
nand U1173 (N_1173,N_965,N_820);
xor U1174 (N_1174,N_969,N_982);
nor U1175 (N_1175,N_929,N_928);
or U1176 (N_1176,N_851,N_842);
or U1177 (N_1177,N_940,N_902);
or U1178 (N_1178,N_911,N_935);
or U1179 (N_1179,N_898,N_885);
nor U1180 (N_1180,N_809,N_881);
or U1181 (N_1181,N_819,N_864);
and U1182 (N_1182,N_991,N_819);
and U1183 (N_1183,N_877,N_816);
and U1184 (N_1184,N_839,N_989);
and U1185 (N_1185,N_858,N_800);
and U1186 (N_1186,N_912,N_873);
or U1187 (N_1187,N_819,N_925);
and U1188 (N_1188,N_943,N_978);
nand U1189 (N_1189,N_982,N_853);
and U1190 (N_1190,N_851,N_805);
and U1191 (N_1191,N_812,N_807);
or U1192 (N_1192,N_945,N_937);
or U1193 (N_1193,N_938,N_855);
and U1194 (N_1194,N_975,N_902);
or U1195 (N_1195,N_840,N_977);
or U1196 (N_1196,N_917,N_962);
and U1197 (N_1197,N_839,N_834);
and U1198 (N_1198,N_955,N_828);
or U1199 (N_1199,N_958,N_909);
nand U1200 (N_1200,N_1152,N_1192);
or U1201 (N_1201,N_1144,N_1157);
or U1202 (N_1202,N_1129,N_1100);
nor U1203 (N_1203,N_1003,N_1089);
nand U1204 (N_1204,N_1166,N_1037);
nand U1205 (N_1205,N_1140,N_1088);
nand U1206 (N_1206,N_1029,N_1188);
and U1207 (N_1207,N_1022,N_1102);
or U1208 (N_1208,N_1014,N_1048);
nor U1209 (N_1209,N_1001,N_1197);
and U1210 (N_1210,N_1039,N_1020);
and U1211 (N_1211,N_1198,N_1094);
nand U1212 (N_1212,N_1175,N_1090);
nor U1213 (N_1213,N_1004,N_1118);
nor U1214 (N_1214,N_1196,N_1116);
and U1215 (N_1215,N_1171,N_1121);
nor U1216 (N_1216,N_1151,N_1050);
or U1217 (N_1217,N_1106,N_1011);
or U1218 (N_1218,N_1136,N_1124);
or U1219 (N_1219,N_1123,N_1109);
nor U1220 (N_1220,N_1169,N_1059);
nand U1221 (N_1221,N_1016,N_1135);
nand U1222 (N_1222,N_1078,N_1111);
or U1223 (N_1223,N_1097,N_1165);
and U1224 (N_1224,N_1126,N_1062);
nand U1225 (N_1225,N_1036,N_1132);
and U1226 (N_1226,N_1045,N_1052);
and U1227 (N_1227,N_1079,N_1194);
or U1228 (N_1228,N_1110,N_1173);
and U1229 (N_1229,N_1178,N_1019);
nor U1230 (N_1230,N_1139,N_1038);
nand U1231 (N_1231,N_1033,N_1160);
nor U1232 (N_1232,N_1164,N_1064);
nand U1233 (N_1233,N_1007,N_1098);
nor U1234 (N_1234,N_1080,N_1112);
nand U1235 (N_1235,N_1172,N_1096);
nor U1236 (N_1236,N_1095,N_1163);
and U1237 (N_1237,N_1083,N_1081);
nand U1238 (N_1238,N_1181,N_1108);
nor U1239 (N_1239,N_1026,N_1184);
nand U1240 (N_1240,N_1074,N_1115);
or U1241 (N_1241,N_1133,N_1055);
nand U1242 (N_1242,N_1187,N_1141);
nor U1243 (N_1243,N_1008,N_1161);
and U1244 (N_1244,N_1068,N_1190);
or U1245 (N_1245,N_1195,N_1137);
nor U1246 (N_1246,N_1066,N_1076);
and U1247 (N_1247,N_1051,N_1149);
nor U1248 (N_1248,N_1056,N_1035);
nor U1249 (N_1249,N_1049,N_1041);
or U1250 (N_1250,N_1138,N_1134);
nand U1251 (N_1251,N_1009,N_1180);
and U1252 (N_1252,N_1176,N_1170);
or U1253 (N_1253,N_1005,N_1073);
nor U1254 (N_1254,N_1077,N_1099);
nor U1255 (N_1255,N_1156,N_1069);
and U1256 (N_1256,N_1189,N_1027);
nor U1257 (N_1257,N_1183,N_1044);
and U1258 (N_1258,N_1128,N_1082);
nand U1259 (N_1259,N_1006,N_1017);
or U1260 (N_1260,N_1046,N_1150);
or U1261 (N_1261,N_1075,N_1168);
nand U1262 (N_1262,N_1167,N_1158);
nand U1263 (N_1263,N_1155,N_1065);
nand U1264 (N_1264,N_1182,N_1114);
or U1265 (N_1265,N_1072,N_1087);
or U1266 (N_1266,N_1030,N_1130);
or U1267 (N_1267,N_1058,N_1021);
nor U1268 (N_1268,N_1120,N_1040);
nor U1269 (N_1269,N_1053,N_1104);
nor U1270 (N_1270,N_1032,N_1148);
or U1271 (N_1271,N_1147,N_1012);
nor U1272 (N_1272,N_1131,N_1119);
nand U1273 (N_1273,N_1093,N_1057);
or U1274 (N_1274,N_1103,N_1146);
nor U1275 (N_1275,N_1043,N_1107);
nand U1276 (N_1276,N_1042,N_1070);
nor U1277 (N_1277,N_1177,N_1063);
or U1278 (N_1278,N_1060,N_1000);
xor U1279 (N_1279,N_1143,N_1142);
nand U1280 (N_1280,N_1199,N_1125);
and U1281 (N_1281,N_1092,N_1159);
or U1282 (N_1282,N_1031,N_1024);
nor U1283 (N_1283,N_1018,N_1015);
nor U1284 (N_1284,N_1154,N_1162);
nor U1285 (N_1285,N_1193,N_1145);
or U1286 (N_1286,N_1086,N_1153);
nor U1287 (N_1287,N_1101,N_1113);
nand U1288 (N_1288,N_1185,N_1084);
and U1289 (N_1289,N_1122,N_1023);
nand U1290 (N_1290,N_1071,N_1067);
or U1291 (N_1291,N_1127,N_1028);
nand U1292 (N_1292,N_1091,N_1085);
and U1293 (N_1293,N_1117,N_1013);
and U1294 (N_1294,N_1186,N_1179);
nand U1295 (N_1295,N_1061,N_1054);
nand U1296 (N_1296,N_1002,N_1010);
and U1297 (N_1297,N_1025,N_1191);
nor U1298 (N_1298,N_1047,N_1105);
or U1299 (N_1299,N_1034,N_1174);
nand U1300 (N_1300,N_1098,N_1091);
and U1301 (N_1301,N_1166,N_1196);
nor U1302 (N_1302,N_1093,N_1038);
and U1303 (N_1303,N_1115,N_1199);
and U1304 (N_1304,N_1163,N_1047);
nand U1305 (N_1305,N_1127,N_1154);
nor U1306 (N_1306,N_1037,N_1109);
and U1307 (N_1307,N_1094,N_1197);
nor U1308 (N_1308,N_1058,N_1124);
nor U1309 (N_1309,N_1186,N_1134);
or U1310 (N_1310,N_1061,N_1148);
and U1311 (N_1311,N_1163,N_1032);
xor U1312 (N_1312,N_1073,N_1039);
or U1313 (N_1313,N_1152,N_1198);
and U1314 (N_1314,N_1107,N_1123);
nor U1315 (N_1315,N_1101,N_1008);
nand U1316 (N_1316,N_1112,N_1021);
and U1317 (N_1317,N_1126,N_1176);
nand U1318 (N_1318,N_1128,N_1070);
nor U1319 (N_1319,N_1174,N_1021);
or U1320 (N_1320,N_1188,N_1089);
and U1321 (N_1321,N_1103,N_1125);
or U1322 (N_1322,N_1127,N_1022);
nand U1323 (N_1323,N_1050,N_1041);
or U1324 (N_1324,N_1173,N_1114);
and U1325 (N_1325,N_1169,N_1174);
and U1326 (N_1326,N_1039,N_1127);
nor U1327 (N_1327,N_1148,N_1001);
nor U1328 (N_1328,N_1132,N_1042);
nand U1329 (N_1329,N_1113,N_1073);
or U1330 (N_1330,N_1032,N_1075);
nor U1331 (N_1331,N_1060,N_1108);
and U1332 (N_1332,N_1127,N_1010);
or U1333 (N_1333,N_1058,N_1139);
and U1334 (N_1334,N_1131,N_1182);
and U1335 (N_1335,N_1091,N_1160);
nand U1336 (N_1336,N_1107,N_1165);
and U1337 (N_1337,N_1042,N_1143);
nand U1338 (N_1338,N_1131,N_1080);
or U1339 (N_1339,N_1189,N_1033);
nand U1340 (N_1340,N_1155,N_1073);
nor U1341 (N_1341,N_1108,N_1151);
nor U1342 (N_1342,N_1174,N_1047);
and U1343 (N_1343,N_1198,N_1113);
nor U1344 (N_1344,N_1109,N_1113);
nor U1345 (N_1345,N_1019,N_1063);
or U1346 (N_1346,N_1197,N_1185);
nand U1347 (N_1347,N_1046,N_1031);
or U1348 (N_1348,N_1044,N_1068);
nor U1349 (N_1349,N_1151,N_1060);
or U1350 (N_1350,N_1052,N_1029);
or U1351 (N_1351,N_1127,N_1125);
nor U1352 (N_1352,N_1190,N_1188);
nand U1353 (N_1353,N_1172,N_1140);
nand U1354 (N_1354,N_1060,N_1090);
nor U1355 (N_1355,N_1121,N_1029);
or U1356 (N_1356,N_1125,N_1063);
and U1357 (N_1357,N_1068,N_1148);
nor U1358 (N_1358,N_1036,N_1160);
or U1359 (N_1359,N_1171,N_1118);
or U1360 (N_1360,N_1064,N_1113);
or U1361 (N_1361,N_1025,N_1178);
or U1362 (N_1362,N_1066,N_1181);
xor U1363 (N_1363,N_1066,N_1118);
nor U1364 (N_1364,N_1087,N_1019);
nor U1365 (N_1365,N_1060,N_1109);
nand U1366 (N_1366,N_1077,N_1183);
or U1367 (N_1367,N_1199,N_1181);
and U1368 (N_1368,N_1097,N_1128);
and U1369 (N_1369,N_1112,N_1152);
and U1370 (N_1370,N_1025,N_1066);
nand U1371 (N_1371,N_1021,N_1090);
nand U1372 (N_1372,N_1012,N_1022);
nor U1373 (N_1373,N_1174,N_1178);
and U1374 (N_1374,N_1183,N_1137);
nor U1375 (N_1375,N_1160,N_1090);
nor U1376 (N_1376,N_1123,N_1144);
and U1377 (N_1377,N_1057,N_1062);
and U1378 (N_1378,N_1097,N_1197);
or U1379 (N_1379,N_1157,N_1085);
or U1380 (N_1380,N_1012,N_1132);
or U1381 (N_1381,N_1102,N_1160);
nand U1382 (N_1382,N_1084,N_1127);
nor U1383 (N_1383,N_1133,N_1147);
or U1384 (N_1384,N_1078,N_1116);
or U1385 (N_1385,N_1130,N_1196);
or U1386 (N_1386,N_1070,N_1149);
or U1387 (N_1387,N_1179,N_1086);
nor U1388 (N_1388,N_1159,N_1143);
and U1389 (N_1389,N_1094,N_1178);
and U1390 (N_1390,N_1004,N_1103);
nand U1391 (N_1391,N_1047,N_1008);
nand U1392 (N_1392,N_1047,N_1082);
or U1393 (N_1393,N_1034,N_1127);
and U1394 (N_1394,N_1056,N_1097);
and U1395 (N_1395,N_1019,N_1112);
nand U1396 (N_1396,N_1090,N_1195);
nand U1397 (N_1397,N_1065,N_1054);
and U1398 (N_1398,N_1146,N_1067);
nand U1399 (N_1399,N_1011,N_1020);
and U1400 (N_1400,N_1290,N_1241);
nor U1401 (N_1401,N_1206,N_1232);
and U1402 (N_1402,N_1243,N_1384);
and U1403 (N_1403,N_1276,N_1287);
or U1404 (N_1404,N_1246,N_1391);
nor U1405 (N_1405,N_1274,N_1208);
or U1406 (N_1406,N_1305,N_1271);
nand U1407 (N_1407,N_1318,N_1263);
and U1408 (N_1408,N_1307,N_1297);
nor U1409 (N_1409,N_1380,N_1265);
nor U1410 (N_1410,N_1349,N_1352);
or U1411 (N_1411,N_1226,N_1239);
nand U1412 (N_1412,N_1293,N_1337);
and U1413 (N_1413,N_1238,N_1209);
or U1414 (N_1414,N_1205,N_1254);
or U1415 (N_1415,N_1366,N_1341);
and U1416 (N_1416,N_1291,N_1317);
nand U1417 (N_1417,N_1396,N_1388);
nor U1418 (N_1418,N_1220,N_1332);
and U1419 (N_1419,N_1218,N_1365);
nand U1420 (N_1420,N_1370,N_1210);
nand U1421 (N_1421,N_1255,N_1236);
or U1422 (N_1422,N_1338,N_1336);
nor U1423 (N_1423,N_1237,N_1377);
or U1424 (N_1424,N_1357,N_1354);
nor U1425 (N_1425,N_1294,N_1267);
or U1426 (N_1426,N_1269,N_1387);
or U1427 (N_1427,N_1345,N_1356);
and U1428 (N_1428,N_1323,N_1343);
nor U1429 (N_1429,N_1266,N_1249);
or U1430 (N_1430,N_1368,N_1311);
nor U1431 (N_1431,N_1224,N_1322);
nor U1432 (N_1432,N_1277,N_1214);
nor U1433 (N_1433,N_1228,N_1285);
nand U1434 (N_1434,N_1248,N_1328);
nor U1435 (N_1435,N_1222,N_1325);
nor U1436 (N_1436,N_1344,N_1273);
nor U1437 (N_1437,N_1286,N_1299);
or U1438 (N_1438,N_1367,N_1264);
or U1439 (N_1439,N_1284,N_1397);
or U1440 (N_1440,N_1288,N_1330);
or U1441 (N_1441,N_1221,N_1378);
and U1442 (N_1442,N_1262,N_1207);
nand U1443 (N_1443,N_1353,N_1240);
nand U1444 (N_1444,N_1363,N_1303);
or U1445 (N_1445,N_1358,N_1348);
and U1446 (N_1446,N_1326,N_1355);
nand U1447 (N_1447,N_1316,N_1217);
and U1448 (N_1448,N_1320,N_1389);
and U1449 (N_1449,N_1329,N_1270);
and U1450 (N_1450,N_1394,N_1379);
nand U1451 (N_1451,N_1324,N_1201);
or U1452 (N_1452,N_1295,N_1260);
or U1453 (N_1453,N_1257,N_1300);
nand U1454 (N_1454,N_1234,N_1242);
nor U1455 (N_1455,N_1256,N_1351);
and U1456 (N_1456,N_1250,N_1200);
nor U1457 (N_1457,N_1335,N_1296);
and U1458 (N_1458,N_1219,N_1229);
or U1459 (N_1459,N_1261,N_1314);
nand U1460 (N_1460,N_1360,N_1334);
or U1461 (N_1461,N_1292,N_1342);
or U1462 (N_1462,N_1302,N_1306);
nor U1463 (N_1463,N_1372,N_1251);
nand U1464 (N_1464,N_1398,N_1227);
nor U1465 (N_1465,N_1359,N_1385);
or U1466 (N_1466,N_1369,N_1321);
and U1467 (N_1467,N_1399,N_1279);
nand U1468 (N_1468,N_1319,N_1392);
or U1469 (N_1469,N_1364,N_1247);
xor U1470 (N_1470,N_1390,N_1204);
or U1471 (N_1471,N_1202,N_1282);
or U1472 (N_1472,N_1346,N_1230);
nand U1473 (N_1473,N_1382,N_1374);
or U1474 (N_1474,N_1381,N_1339);
or U1475 (N_1475,N_1215,N_1289);
and U1476 (N_1476,N_1272,N_1386);
and U1477 (N_1477,N_1312,N_1281);
or U1478 (N_1478,N_1340,N_1233);
nor U1479 (N_1479,N_1373,N_1253);
and U1480 (N_1480,N_1245,N_1347);
and U1481 (N_1481,N_1225,N_1252);
and U1482 (N_1482,N_1231,N_1309);
and U1483 (N_1483,N_1350,N_1283);
nor U1484 (N_1484,N_1223,N_1216);
or U1485 (N_1485,N_1308,N_1268);
nor U1486 (N_1486,N_1393,N_1371);
nand U1487 (N_1487,N_1301,N_1304);
and U1488 (N_1488,N_1376,N_1313);
or U1489 (N_1489,N_1362,N_1235);
nor U1490 (N_1490,N_1331,N_1327);
or U1491 (N_1491,N_1203,N_1212);
or U1492 (N_1492,N_1259,N_1275);
nor U1493 (N_1493,N_1375,N_1244);
nor U1494 (N_1494,N_1278,N_1315);
nand U1495 (N_1495,N_1280,N_1333);
nand U1496 (N_1496,N_1298,N_1310);
or U1497 (N_1497,N_1211,N_1258);
nand U1498 (N_1498,N_1361,N_1383);
and U1499 (N_1499,N_1395,N_1213);
nand U1500 (N_1500,N_1345,N_1260);
nand U1501 (N_1501,N_1293,N_1355);
and U1502 (N_1502,N_1205,N_1387);
nor U1503 (N_1503,N_1226,N_1203);
nand U1504 (N_1504,N_1390,N_1359);
and U1505 (N_1505,N_1345,N_1275);
nand U1506 (N_1506,N_1201,N_1275);
nor U1507 (N_1507,N_1204,N_1355);
nand U1508 (N_1508,N_1219,N_1396);
nand U1509 (N_1509,N_1373,N_1222);
nor U1510 (N_1510,N_1393,N_1337);
or U1511 (N_1511,N_1382,N_1222);
or U1512 (N_1512,N_1349,N_1301);
or U1513 (N_1513,N_1238,N_1302);
or U1514 (N_1514,N_1374,N_1394);
nand U1515 (N_1515,N_1252,N_1313);
nor U1516 (N_1516,N_1222,N_1337);
or U1517 (N_1517,N_1334,N_1244);
nor U1518 (N_1518,N_1298,N_1293);
and U1519 (N_1519,N_1348,N_1293);
nor U1520 (N_1520,N_1295,N_1378);
nand U1521 (N_1521,N_1230,N_1365);
nand U1522 (N_1522,N_1244,N_1327);
or U1523 (N_1523,N_1333,N_1300);
nor U1524 (N_1524,N_1385,N_1260);
or U1525 (N_1525,N_1206,N_1377);
nand U1526 (N_1526,N_1332,N_1222);
and U1527 (N_1527,N_1207,N_1366);
or U1528 (N_1528,N_1331,N_1253);
nand U1529 (N_1529,N_1276,N_1356);
or U1530 (N_1530,N_1255,N_1296);
nand U1531 (N_1531,N_1210,N_1247);
nor U1532 (N_1532,N_1226,N_1323);
and U1533 (N_1533,N_1374,N_1222);
nor U1534 (N_1534,N_1225,N_1306);
and U1535 (N_1535,N_1332,N_1382);
nand U1536 (N_1536,N_1388,N_1258);
nand U1537 (N_1537,N_1349,N_1271);
nand U1538 (N_1538,N_1213,N_1231);
nand U1539 (N_1539,N_1354,N_1256);
nor U1540 (N_1540,N_1291,N_1331);
nor U1541 (N_1541,N_1398,N_1387);
or U1542 (N_1542,N_1378,N_1212);
and U1543 (N_1543,N_1241,N_1316);
or U1544 (N_1544,N_1236,N_1226);
or U1545 (N_1545,N_1297,N_1340);
nand U1546 (N_1546,N_1215,N_1279);
or U1547 (N_1547,N_1353,N_1304);
nor U1548 (N_1548,N_1358,N_1207);
and U1549 (N_1549,N_1301,N_1230);
nand U1550 (N_1550,N_1218,N_1351);
nand U1551 (N_1551,N_1348,N_1386);
nor U1552 (N_1552,N_1335,N_1323);
nor U1553 (N_1553,N_1365,N_1248);
and U1554 (N_1554,N_1330,N_1382);
nor U1555 (N_1555,N_1233,N_1309);
and U1556 (N_1556,N_1385,N_1292);
nand U1557 (N_1557,N_1245,N_1372);
nand U1558 (N_1558,N_1257,N_1301);
nand U1559 (N_1559,N_1241,N_1332);
and U1560 (N_1560,N_1230,N_1322);
nor U1561 (N_1561,N_1250,N_1321);
and U1562 (N_1562,N_1297,N_1377);
xor U1563 (N_1563,N_1225,N_1386);
and U1564 (N_1564,N_1381,N_1342);
nand U1565 (N_1565,N_1386,N_1338);
or U1566 (N_1566,N_1223,N_1312);
nor U1567 (N_1567,N_1354,N_1258);
or U1568 (N_1568,N_1268,N_1381);
nand U1569 (N_1569,N_1292,N_1361);
or U1570 (N_1570,N_1248,N_1312);
or U1571 (N_1571,N_1371,N_1239);
and U1572 (N_1572,N_1200,N_1340);
nor U1573 (N_1573,N_1320,N_1258);
nor U1574 (N_1574,N_1291,N_1332);
nor U1575 (N_1575,N_1275,N_1278);
and U1576 (N_1576,N_1323,N_1307);
nand U1577 (N_1577,N_1347,N_1337);
nand U1578 (N_1578,N_1201,N_1257);
nand U1579 (N_1579,N_1302,N_1284);
nor U1580 (N_1580,N_1288,N_1263);
nand U1581 (N_1581,N_1247,N_1386);
or U1582 (N_1582,N_1384,N_1270);
nand U1583 (N_1583,N_1351,N_1386);
or U1584 (N_1584,N_1298,N_1395);
nand U1585 (N_1585,N_1365,N_1380);
or U1586 (N_1586,N_1393,N_1382);
and U1587 (N_1587,N_1334,N_1268);
nor U1588 (N_1588,N_1331,N_1344);
and U1589 (N_1589,N_1254,N_1371);
nor U1590 (N_1590,N_1256,N_1225);
and U1591 (N_1591,N_1320,N_1294);
and U1592 (N_1592,N_1261,N_1382);
or U1593 (N_1593,N_1250,N_1368);
and U1594 (N_1594,N_1392,N_1323);
nand U1595 (N_1595,N_1225,N_1270);
and U1596 (N_1596,N_1229,N_1221);
and U1597 (N_1597,N_1387,N_1376);
nand U1598 (N_1598,N_1281,N_1396);
and U1599 (N_1599,N_1379,N_1376);
nand U1600 (N_1600,N_1480,N_1589);
nor U1601 (N_1601,N_1556,N_1577);
and U1602 (N_1602,N_1426,N_1494);
or U1603 (N_1603,N_1486,N_1575);
and U1604 (N_1604,N_1415,N_1544);
or U1605 (N_1605,N_1401,N_1460);
and U1606 (N_1606,N_1402,N_1412);
nor U1607 (N_1607,N_1411,N_1591);
and U1608 (N_1608,N_1525,N_1418);
or U1609 (N_1609,N_1536,N_1454);
nor U1610 (N_1610,N_1573,N_1441);
nand U1611 (N_1611,N_1523,N_1554);
nor U1612 (N_1612,N_1457,N_1564);
or U1613 (N_1613,N_1429,N_1500);
and U1614 (N_1614,N_1546,N_1482);
and U1615 (N_1615,N_1407,N_1528);
and U1616 (N_1616,N_1541,N_1485);
or U1617 (N_1617,N_1459,N_1537);
and U1618 (N_1618,N_1474,N_1484);
nand U1619 (N_1619,N_1581,N_1592);
nor U1620 (N_1620,N_1462,N_1543);
or U1621 (N_1621,N_1493,N_1571);
and U1622 (N_1622,N_1532,N_1508);
and U1623 (N_1623,N_1425,N_1538);
nor U1624 (N_1624,N_1467,N_1568);
or U1625 (N_1625,N_1522,N_1550);
nand U1626 (N_1626,N_1535,N_1434);
nor U1627 (N_1627,N_1489,N_1451);
or U1628 (N_1628,N_1582,N_1405);
nand U1629 (N_1629,N_1507,N_1468);
nor U1630 (N_1630,N_1501,N_1566);
nor U1631 (N_1631,N_1512,N_1587);
nand U1632 (N_1632,N_1513,N_1437);
and U1633 (N_1633,N_1560,N_1553);
and U1634 (N_1634,N_1479,N_1403);
and U1635 (N_1635,N_1400,N_1455);
nor U1636 (N_1636,N_1511,N_1406);
nor U1637 (N_1637,N_1574,N_1533);
nor U1638 (N_1638,N_1481,N_1471);
nor U1639 (N_1639,N_1516,N_1586);
nand U1640 (N_1640,N_1469,N_1510);
and U1641 (N_1641,N_1408,N_1440);
and U1642 (N_1642,N_1521,N_1472);
nor U1643 (N_1643,N_1476,N_1514);
xnor U1644 (N_1644,N_1596,N_1428);
nor U1645 (N_1645,N_1475,N_1583);
nand U1646 (N_1646,N_1595,N_1593);
nor U1647 (N_1647,N_1404,N_1545);
and U1648 (N_1648,N_1442,N_1561);
nand U1649 (N_1649,N_1549,N_1584);
nand U1650 (N_1650,N_1558,N_1435);
nor U1651 (N_1651,N_1436,N_1423);
nor U1652 (N_1652,N_1557,N_1519);
and U1653 (N_1653,N_1420,N_1509);
and U1654 (N_1654,N_1430,N_1416);
and U1655 (N_1655,N_1433,N_1456);
nand U1656 (N_1656,N_1579,N_1413);
and U1657 (N_1657,N_1539,N_1518);
and U1658 (N_1658,N_1470,N_1599);
nor U1659 (N_1659,N_1542,N_1450);
nand U1660 (N_1660,N_1520,N_1515);
or U1661 (N_1661,N_1424,N_1438);
nand U1662 (N_1662,N_1414,N_1491);
and U1663 (N_1663,N_1547,N_1463);
nor U1664 (N_1664,N_1567,N_1458);
and U1665 (N_1665,N_1597,N_1580);
nor U1666 (N_1666,N_1529,N_1540);
nor U1667 (N_1667,N_1443,N_1452);
nor U1668 (N_1668,N_1551,N_1530);
nor U1669 (N_1669,N_1502,N_1505);
and U1670 (N_1670,N_1496,N_1478);
nand U1671 (N_1671,N_1570,N_1444);
nand U1672 (N_1672,N_1439,N_1598);
and U1673 (N_1673,N_1431,N_1449);
nor U1674 (N_1674,N_1562,N_1465);
and U1675 (N_1675,N_1422,N_1563);
and U1676 (N_1676,N_1531,N_1448);
and U1677 (N_1677,N_1588,N_1477);
xor U1678 (N_1678,N_1572,N_1504);
or U1679 (N_1679,N_1578,N_1499);
and U1680 (N_1680,N_1534,N_1461);
and U1681 (N_1681,N_1552,N_1421);
nand U1682 (N_1682,N_1569,N_1576);
nor U1683 (N_1683,N_1585,N_1432);
nor U1684 (N_1684,N_1410,N_1487);
nand U1685 (N_1685,N_1492,N_1506);
or U1686 (N_1686,N_1464,N_1526);
nor U1687 (N_1687,N_1548,N_1565);
nand U1688 (N_1688,N_1594,N_1503);
and U1689 (N_1689,N_1498,N_1473);
nor U1690 (N_1690,N_1417,N_1427);
and U1691 (N_1691,N_1447,N_1490);
and U1692 (N_1692,N_1517,N_1497);
and U1693 (N_1693,N_1559,N_1555);
and U1694 (N_1694,N_1527,N_1488);
or U1695 (N_1695,N_1446,N_1453);
and U1696 (N_1696,N_1590,N_1419);
and U1697 (N_1697,N_1445,N_1409);
or U1698 (N_1698,N_1524,N_1483);
nor U1699 (N_1699,N_1466,N_1495);
and U1700 (N_1700,N_1495,N_1462);
nor U1701 (N_1701,N_1508,N_1510);
nand U1702 (N_1702,N_1546,N_1439);
nand U1703 (N_1703,N_1465,N_1555);
nand U1704 (N_1704,N_1431,N_1577);
nor U1705 (N_1705,N_1552,N_1488);
and U1706 (N_1706,N_1574,N_1592);
and U1707 (N_1707,N_1499,N_1563);
and U1708 (N_1708,N_1450,N_1575);
nand U1709 (N_1709,N_1580,N_1450);
or U1710 (N_1710,N_1503,N_1455);
or U1711 (N_1711,N_1459,N_1596);
or U1712 (N_1712,N_1576,N_1467);
and U1713 (N_1713,N_1559,N_1502);
or U1714 (N_1714,N_1521,N_1450);
nand U1715 (N_1715,N_1568,N_1448);
nor U1716 (N_1716,N_1503,N_1541);
or U1717 (N_1717,N_1595,N_1579);
and U1718 (N_1718,N_1509,N_1480);
nand U1719 (N_1719,N_1544,N_1455);
nor U1720 (N_1720,N_1583,N_1507);
nand U1721 (N_1721,N_1419,N_1463);
nand U1722 (N_1722,N_1506,N_1416);
and U1723 (N_1723,N_1582,N_1542);
nor U1724 (N_1724,N_1496,N_1406);
or U1725 (N_1725,N_1481,N_1540);
and U1726 (N_1726,N_1558,N_1481);
or U1727 (N_1727,N_1539,N_1479);
nor U1728 (N_1728,N_1420,N_1438);
and U1729 (N_1729,N_1423,N_1460);
and U1730 (N_1730,N_1579,N_1424);
or U1731 (N_1731,N_1426,N_1428);
and U1732 (N_1732,N_1463,N_1505);
nand U1733 (N_1733,N_1557,N_1570);
and U1734 (N_1734,N_1443,N_1434);
nor U1735 (N_1735,N_1410,N_1400);
and U1736 (N_1736,N_1516,N_1423);
nand U1737 (N_1737,N_1555,N_1497);
or U1738 (N_1738,N_1553,N_1430);
nor U1739 (N_1739,N_1493,N_1543);
nor U1740 (N_1740,N_1564,N_1430);
nor U1741 (N_1741,N_1463,N_1531);
nand U1742 (N_1742,N_1548,N_1457);
nor U1743 (N_1743,N_1434,N_1530);
and U1744 (N_1744,N_1526,N_1572);
or U1745 (N_1745,N_1587,N_1563);
and U1746 (N_1746,N_1532,N_1418);
or U1747 (N_1747,N_1459,N_1534);
xor U1748 (N_1748,N_1556,N_1562);
nor U1749 (N_1749,N_1545,N_1501);
nor U1750 (N_1750,N_1526,N_1556);
nand U1751 (N_1751,N_1471,N_1442);
and U1752 (N_1752,N_1455,N_1541);
and U1753 (N_1753,N_1490,N_1555);
nand U1754 (N_1754,N_1595,N_1493);
and U1755 (N_1755,N_1542,N_1428);
and U1756 (N_1756,N_1520,N_1565);
nand U1757 (N_1757,N_1444,N_1587);
nor U1758 (N_1758,N_1415,N_1455);
nor U1759 (N_1759,N_1456,N_1551);
and U1760 (N_1760,N_1468,N_1461);
nand U1761 (N_1761,N_1413,N_1553);
nor U1762 (N_1762,N_1477,N_1573);
and U1763 (N_1763,N_1525,N_1453);
and U1764 (N_1764,N_1500,N_1592);
nand U1765 (N_1765,N_1402,N_1468);
nand U1766 (N_1766,N_1476,N_1426);
xnor U1767 (N_1767,N_1534,N_1570);
and U1768 (N_1768,N_1570,N_1490);
and U1769 (N_1769,N_1447,N_1577);
nor U1770 (N_1770,N_1443,N_1571);
and U1771 (N_1771,N_1476,N_1418);
nor U1772 (N_1772,N_1562,N_1498);
or U1773 (N_1773,N_1459,N_1597);
nor U1774 (N_1774,N_1539,N_1492);
nand U1775 (N_1775,N_1459,N_1575);
and U1776 (N_1776,N_1458,N_1459);
nor U1777 (N_1777,N_1407,N_1595);
nor U1778 (N_1778,N_1594,N_1489);
or U1779 (N_1779,N_1464,N_1555);
and U1780 (N_1780,N_1587,N_1562);
nor U1781 (N_1781,N_1411,N_1422);
and U1782 (N_1782,N_1513,N_1507);
nor U1783 (N_1783,N_1541,N_1578);
nor U1784 (N_1784,N_1480,N_1547);
nor U1785 (N_1785,N_1455,N_1569);
xor U1786 (N_1786,N_1586,N_1485);
nor U1787 (N_1787,N_1511,N_1585);
and U1788 (N_1788,N_1437,N_1583);
nor U1789 (N_1789,N_1505,N_1418);
or U1790 (N_1790,N_1426,N_1438);
or U1791 (N_1791,N_1425,N_1470);
nand U1792 (N_1792,N_1409,N_1427);
nor U1793 (N_1793,N_1584,N_1489);
nand U1794 (N_1794,N_1421,N_1409);
nor U1795 (N_1795,N_1540,N_1578);
nor U1796 (N_1796,N_1496,N_1429);
and U1797 (N_1797,N_1543,N_1498);
xor U1798 (N_1798,N_1411,N_1534);
or U1799 (N_1799,N_1431,N_1521);
and U1800 (N_1800,N_1757,N_1665);
and U1801 (N_1801,N_1775,N_1784);
and U1802 (N_1802,N_1673,N_1790);
nand U1803 (N_1803,N_1752,N_1716);
nand U1804 (N_1804,N_1638,N_1772);
and U1805 (N_1805,N_1660,N_1612);
nand U1806 (N_1806,N_1602,N_1605);
or U1807 (N_1807,N_1780,N_1652);
nor U1808 (N_1808,N_1656,N_1798);
nor U1809 (N_1809,N_1649,N_1789);
and U1810 (N_1810,N_1704,N_1733);
or U1811 (N_1811,N_1648,N_1601);
nand U1812 (N_1812,N_1619,N_1632);
nand U1813 (N_1813,N_1712,N_1725);
nor U1814 (N_1814,N_1754,N_1771);
and U1815 (N_1815,N_1669,N_1753);
and U1816 (N_1816,N_1685,N_1688);
nor U1817 (N_1817,N_1709,N_1626);
nor U1818 (N_1818,N_1639,N_1615);
nor U1819 (N_1819,N_1779,N_1692);
or U1820 (N_1820,N_1710,N_1631);
nand U1821 (N_1821,N_1668,N_1676);
nand U1822 (N_1822,N_1751,N_1647);
or U1823 (N_1823,N_1707,N_1706);
or U1824 (N_1824,N_1726,N_1698);
nor U1825 (N_1825,N_1607,N_1654);
or U1826 (N_1826,N_1799,N_1682);
or U1827 (N_1827,N_1610,N_1611);
and U1828 (N_1828,N_1658,N_1614);
or U1829 (N_1829,N_1756,N_1613);
or U1830 (N_1830,N_1791,N_1641);
nor U1831 (N_1831,N_1618,N_1686);
and U1832 (N_1832,N_1655,N_1730);
nor U1833 (N_1833,N_1623,N_1739);
or U1834 (N_1834,N_1770,N_1731);
nand U1835 (N_1835,N_1696,N_1732);
or U1836 (N_1836,N_1759,N_1636);
nor U1837 (N_1837,N_1720,N_1643);
nor U1838 (N_1838,N_1690,N_1748);
or U1839 (N_1839,N_1785,N_1721);
or U1840 (N_1840,N_1747,N_1620);
nand U1841 (N_1841,N_1627,N_1633);
or U1842 (N_1842,N_1600,N_1761);
nand U1843 (N_1843,N_1793,N_1760);
nor U1844 (N_1844,N_1650,N_1765);
and U1845 (N_1845,N_1794,N_1738);
nand U1846 (N_1846,N_1746,N_1603);
nor U1847 (N_1847,N_1745,N_1637);
and U1848 (N_1848,N_1608,N_1702);
and U1849 (N_1849,N_1727,N_1781);
nand U1850 (N_1850,N_1767,N_1737);
nand U1851 (N_1851,N_1679,N_1674);
nand U1852 (N_1852,N_1606,N_1773);
nor U1853 (N_1853,N_1792,N_1677);
or U1854 (N_1854,N_1689,N_1640);
and U1855 (N_1855,N_1635,N_1742);
and U1856 (N_1856,N_1699,N_1651);
nor U1857 (N_1857,N_1796,N_1675);
nor U1858 (N_1858,N_1769,N_1678);
nor U1859 (N_1859,N_1680,N_1728);
nor U1860 (N_1860,N_1684,N_1788);
and U1861 (N_1861,N_1735,N_1630);
and U1862 (N_1862,N_1695,N_1642);
nor U1863 (N_1863,N_1703,N_1740);
and U1864 (N_1864,N_1729,N_1661);
or U1865 (N_1865,N_1717,N_1722);
nand U1866 (N_1866,N_1755,N_1750);
nor U1867 (N_1867,N_1604,N_1663);
and U1868 (N_1868,N_1758,N_1718);
and U1869 (N_1869,N_1624,N_1719);
nor U1870 (N_1870,N_1736,N_1659);
and U1871 (N_1871,N_1700,N_1713);
nand U1872 (N_1872,N_1671,N_1694);
and U1873 (N_1873,N_1776,N_1708);
nor U1874 (N_1874,N_1646,N_1657);
nand U1875 (N_1875,N_1634,N_1778);
or U1876 (N_1876,N_1666,N_1697);
nor U1877 (N_1877,N_1711,N_1714);
and U1878 (N_1878,N_1724,N_1687);
and U1879 (N_1879,N_1629,N_1644);
nand U1880 (N_1880,N_1616,N_1681);
and U1881 (N_1881,N_1723,N_1701);
or U1882 (N_1882,N_1783,N_1777);
nand U1883 (N_1883,N_1628,N_1795);
and U1884 (N_1884,N_1672,N_1762);
or U1885 (N_1885,N_1609,N_1797);
and U1886 (N_1886,N_1774,N_1763);
nor U1887 (N_1887,N_1766,N_1653);
and U1888 (N_1888,N_1741,N_1625);
or U1889 (N_1889,N_1787,N_1670);
and U1890 (N_1890,N_1645,N_1743);
nand U1891 (N_1891,N_1621,N_1683);
and U1892 (N_1892,N_1617,N_1764);
nor U1893 (N_1893,N_1786,N_1667);
and U1894 (N_1894,N_1768,N_1662);
nor U1895 (N_1895,N_1664,N_1749);
or U1896 (N_1896,N_1734,N_1693);
xor U1897 (N_1897,N_1782,N_1691);
and U1898 (N_1898,N_1705,N_1744);
nand U1899 (N_1899,N_1622,N_1715);
nor U1900 (N_1900,N_1650,N_1715);
nor U1901 (N_1901,N_1612,N_1649);
or U1902 (N_1902,N_1654,N_1717);
nand U1903 (N_1903,N_1797,N_1674);
nor U1904 (N_1904,N_1674,N_1716);
nand U1905 (N_1905,N_1603,N_1659);
nor U1906 (N_1906,N_1786,N_1603);
nor U1907 (N_1907,N_1718,N_1705);
xor U1908 (N_1908,N_1636,N_1766);
nor U1909 (N_1909,N_1763,N_1726);
or U1910 (N_1910,N_1625,N_1646);
or U1911 (N_1911,N_1716,N_1604);
or U1912 (N_1912,N_1780,N_1624);
or U1913 (N_1913,N_1638,N_1699);
and U1914 (N_1914,N_1770,N_1695);
or U1915 (N_1915,N_1622,N_1781);
nor U1916 (N_1916,N_1709,N_1747);
nor U1917 (N_1917,N_1610,N_1649);
and U1918 (N_1918,N_1625,N_1616);
nor U1919 (N_1919,N_1626,N_1686);
and U1920 (N_1920,N_1605,N_1747);
and U1921 (N_1921,N_1711,N_1689);
and U1922 (N_1922,N_1672,N_1724);
nor U1923 (N_1923,N_1654,N_1621);
nand U1924 (N_1924,N_1713,N_1621);
and U1925 (N_1925,N_1701,N_1691);
xnor U1926 (N_1926,N_1619,N_1729);
or U1927 (N_1927,N_1701,N_1625);
and U1928 (N_1928,N_1618,N_1615);
nor U1929 (N_1929,N_1619,N_1695);
nor U1930 (N_1930,N_1617,N_1719);
nand U1931 (N_1931,N_1792,N_1682);
or U1932 (N_1932,N_1621,N_1712);
and U1933 (N_1933,N_1763,N_1718);
or U1934 (N_1934,N_1621,N_1701);
and U1935 (N_1935,N_1616,N_1632);
or U1936 (N_1936,N_1674,N_1607);
and U1937 (N_1937,N_1753,N_1799);
nor U1938 (N_1938,N_1662,N_1777);
and U1939 (N_1939,N_1616,N_1786);
nor U1940 (N_1940,N_1769,N_1786);
and U1941 (N_1941,N_1677,N_1745);
and U1942 (N_1942,N_1720,N_1653);
nor U1943 (N_1943,N_1600,N_1699);
nor U1944 (N_1944,N_1755,N_1741);
and U1945 (N_1945,N_1776,N_1756);
or U1946 (N_1946,N_1606,N_1623);
nand U1947 (N_1947,N_1744,N_1624);
and U1948 (N_1948,N_1643,N_1740);
nor U1949 (N_1949,N_1692,N_1634);
or U1950 (N_1950,N_1762,N_1669);
nor U1951 (N_1951,N_1670,N_1663);
and U1952 (N_1952,N_1786,N_1687);
or U1953 (N_1953,N_1749,N_1759);
or U1954 (N_1954,N_1727,N_1675);
nand U1955 (N_1955,N_1796,N_1700);
nand U1956 (N_1956,N_1673,N_1683);
nand U1957 (N_1957,N_1749,N_1642);
and U1958 (N_1958,N_1697,N_1664);
nand U1959 (N_1959,N_1611,N_1765);
nor U1960 (N_1960,N_1785,N_1745);
or U1961 (N_1961,N_1648,N_1702);
nand U1962 (N_1962,N_1739,N_1652);
or U1963 (N_1963,N_1672,N_1630);
and U1964 (N_1964,N_1781,N_1616);
nand U1965 (N_1965,N_1688,N_1756);
or U1966 (N_1966,N_1622,N_1796);
nand U1967 (N_1967,N_1783,N_1782);
nand U1968 (N_1968,N_1745,N_1797);
nor U1969 (N_1969,N_1657,N_1659);
nor U1970 (N_1970,N_1741,N_1731);
nor U1971 (N_1971,N_1768,N_1757);
nor U1972 (N_1972,N_1762,N_1784);
nor U1973 (N_1973,N_1614,N_1666);
or U1974 (N_1974,N_1774,N_1666);
or U1975 (N_1975,N_1785,N_1759);
or U1976 (N_1976,N_1669,N_1731);
nor U1977 (N_1977,N_1738,N_1752);
nand U1978 (N_1978,N_1739,N_1752);
nor U1979 (N_1979,N_1650,N_1772);
and U1980 (N_1980,N_1615,N_1672);
or U1981 (N_1981,N_1637,N_1771);
and U1982 (N_1982,N_1785,N_1647);
nand U1983 (N_1983,N_1619,N_1629);
or U1984 (N_1984,N_1672,N_1613);
nand U1985 (N_1985,N_1753,N_1762);
and U1986 (N_1986,N_1724,N_1773);
or U1987 (N_1987,N_1681,N_1691);
or U1988 (N_1988,N_1662,N_1602);
or U1989 (N_1989,N_1750,N_1679);
nand U1990 (N_1990,N_1644,N_1657);
nor U1991 (N_1991,N_1776,N_1686);
or U1992 (N_1992,N_1701,N_1764);
and U1993 (N_1993,N_1694,N_1685);
or U1994 (N_1994,N_1693,N_1714);
nand U1995 (N_1995,N_1760,N_1676);
or U1996 (N_1996,N_1785,N_1662);
and U1997 (N_1997,N_1725,N_1668);
and U1998 (N_1998,N_1674,N_1733);
nor U1999 (N_1999,N_1716,N_1782);
nand U2000 (N_2000,N_1965,N_1980);
and U2001 (N_2001,N_1967,N_1916);
nand U2002 (N_2002,N_1816,N_1819);
nor U2003 (N_2003,N_1820,N_1925);
nor U2004 (N_2004,N_1898,N_1912);
nand U2005 (N_2005,N_1988,N_1983);
nor U2006 (N_2006,N_1871,N_1861);
nand U2007 (N_2007,N_1917,N_1963);
nand U2008 (N_2008,N_1902,N_1866);
and U2009 (N_2009,N_1811,N_1937);
nand U2010 (N_2010,N_1973,N_1952);
nand U2011 (N_2011,N_1878,N_1998);
and U2012 (N_2012,N_1985,N_1882);
and U2013 (N_2013,N_1885,N_1807);
nor U2014 (N_2014,N_1859,N_1897);
nand U2015 (N_2015,N_1913,N_1884);
and U2016 (N_2016,N_1954,N_1883);
nand U2017 (N_2017,N_1945,N_1947);
and U2018 (N_2018,N_1975,N_1972);
or U2019 (N_2019,N_1818,N_1924);
and U2020 (N_2020,N_1932,N_1931);
nand U2021 (N_2021,N_1854,N_1817);
or U2022 (N_2022,N_1872,N_1837);
nor U2023 (N_2023,N_1930,N_1961);
nand U2024 (N_2024,N_1939,N_1891);
or U2025 (N_2025,N_1844,N_1944);
nor U2026 (N_2026,N_1896,N_1946);
nor U2027 (N_2027,N_1823,N_1888);
nor U2028 (N_2028,N_1969,N_1836);
nand U2029 (N_2029,N_1886,N_1832);
or U2030 (N_2030,N_1941,N_1949);
or U2031 (N_2031,N_1846,N_1852);
and U2032 (N_2032,N_1953,N_1959);
nand U2033 (N_2033,N_1922,N_1848);
nand U2034 (N_2034,N_1986,N_1976);
nor U2035 (N_2035,N_1813,N_1831);
nand U2036 (N_2036,N_1920,N_1803);
nand U2037 (N_2037,N_1869,N_1905);
nand U2038 (N_2038,N_1996,N_1857);
and U2039 (N_2039,N_1995,N_1870);
nor U2040 (N_2040,N_1858,N_1970);
or U2041 (N_2041,N_1933,N_1966);
or U2042 (N_2042,N_1929,N_1971);
nand U2043 (N_2043,N_1950,N_1877);
nor U2044 (N_2044,N_1994,N_1951);
nor U2045 (N_2045,N_1802,N_1801);
nand U2046 (N_2046,N_1907,N_1982);
and U2047 (N_2047,N_1825,N_1847);
and U2048 (N_2048,N_1915,N_1958);
and U2049 (N_2049,N_1838,N_1806);
or U2050 (N_2050,N_1923,N_1873);
and U2051 (N_2051,N_1899,N_1892);
nor U2052 (N_2052,N_1979,N_1853);
or U2053 (N_2053,N_1865,N_1812);
and U2054 (N_2054,N_1955,N_1850);
nand U2055 (N_2055,N_1936,N_1978);
nand U2056 (N_2056,N_1908,N_1867);
and U2057 (N_2057,N_1889,N_1822);
nand U2058 (N_2058,N_1828,N_1809);
and U2059 (N_2059,N_1943,N_1834);
and U2060 (N_2060,N_1993,N_1842);
nor U2061 (N_2061,N_1957,N_1999);
nor U2062 (N_2062,N_1938,N_1981);
and U2063 (N_2063,N_1826,N_1879);
or U2064 (N_2064,N_1868,N_1926);
nand U2065 (N_2065,N_1841,N_1855);
xor U2066 (N_2066,N_1962,N_1845);
or U2067 (N_2067,N_1942,N_1821);
nand U2068 (N_2068,N_1840,N_1856);
nand U2069 (N_2069,N_1843,N_1895);
and U2070 (N_2070,N_1989,N_1928);
nor U2071 (N_2071,N_1991,N_1824);
and U2072 (N_2072,N_1997,N_1956);
and U2073 (N_2073,N_1919,N_1910);
nand U2074 (N_2074,N_1880,N_1992);
nand U2075 (N_2075,N_1934,N_1906);
nand U2076 (N_2076,N_1827,N_1968);
or U2077 (N_2077,N_1881,N_1876);
and U2078 (N_2078,N_1875,N_1890);
nand U2079 (N_2079,N_1833,N_1990);
and U2080 (N_2080,N_1808,N_1805);
or U2081 (N_2081,N_1804,N_1810);
nor U2082 (N_2082,N_1911,N_1901);
nand U2083 (N_2083,N_1940,N_1948);
or U2084 (N_2084,N_1849,N_1830);
nor U2085 (N_2085,N_1887,N_1862);
or U2086 (N_2086,N_1863,N_1800);
nor U2087 (N_2087,N_1894,N_1977);
nor U2088 (N_2088,N_1914,N_1904);
and U2089 (N_2089,N_1984,N_1974);
nand U2090 (N_2090,N_1851,N_1829);
nand U2091 (N_2091,N_1903,N_1874);
or U2092 (N_2092,N_1860,N_1839);
and U2093 (N_2093,N_1814,N_1835);
and U2094 (N_2094,N_1918,N_1893);
and U2095 (N_2095,N_1900,N_1987);
or U2096 (N_2096,N_1921,N_1960);
nand U2097 (N_2097,N_1909,N_1815);
or U2098 (N_2098,N_1964,N_1935);
and U2099 (N_2099,N_1927,N_1864);
nor U2100 (N_2100,N_1969,N_1944);
or U2101 (N_2101,N_1989,N_1923);
or U2102 (N_2102,N_1986,N_1876);
or U2103 (N_2103,N_1970,N_1867);
nand U2104 (N_2104,N_1956,N_1938);
xor U2105 (N_2105,N_1991,N_1915);
and U2106 (N_2106,N_1954,N_1921);
nand U2107 (N_2107,N_1946,N_1892);
nand U2108 (N_2108,N_1824,N_1930);
or U2109 (N_2109,N_1913,N_1911);
nor U2110 (N_2110,N_1961,N_1871);
nor U2111 (N_2111,N_1993,N_1869);
nand U2112 (N_2112,N_1924,N_1896);
xor U2113 (N_2113,N_1862,N_1872);
or U2114 (N_2114,N_1988,N_1986);
nor U2115 (N_2115,N_1860,N_1906);
or U2116 (N_2116,N_1902,N_1940);
or U2117 (N_2117,N_1920,N_1979);
nand U2118 (N_2118,N_1884,N_1994);
or U2119 (N_2119,N_1957,N_1844);
or U2120 (N_2120,N_1878,N_1814);
or U2121 (N_2121,N_1856,N_1926);
and U2122 (N_2122,N_1913,N_1854);
nand U2123 (N_2123,N_1931,N_1907);
nor U2124 (N_2124,N_1959,N_1873);
nor U2125 (N_2125,N_1885,N_1827);
nor U2126 (N_2126,N_1962,N_1924);
and U2127 (N_2127,N_1965,N_1882);
and U2128 (N_2128,N_1861,N_1998);
or U2129 (N_2129,N_1897,N_1930);
nor U2130 (N_2130,N_1931,N_1910);
or U2131 (N_2131,N_1810,N_1935);
or U2132 (N_2132,N_1859,N_1962);
and U2133 (N_2133,N_1818,N_1816);
or U2134 (N_2134,N_1977,N_1852);
or U2135 (N_2135,N_1825,N_1990);
or U2136 (N_2136,N_1816,N_1886);
and U2137 (N_2137,N_1835,N_1930);
nand U2138 (N_2138,N_1851,N_1803);
and U2139 (N_2139,N_1969,N_1921);
nand U2140 (N_2140,N_1818,N_1960);
nand U2141 (N_2141,N_1992,N_1998);
nand U2142 (N_2142,N_1862,N_1987);
and U2143 (N_2143,N_1830,N_1913);
and U2144 (N_2144,N_1928,N_1941);
nand U2145 (N_2145,N_1855,N_1833);
and U2146 (N_2146,N_1930,N_1872);
or U2147 (N_2147,N_1998,N_1909);
nand U2148 (N_2148,N_1852,N_1955);
or U2149 (N_2149,N_1841,N_1922);
and U2150 (N_2150,N_1921,N_1823);
nand U2151 (N_2151,N_1867,N_1844);
nor U2152 (N_2152,N_1922,N_1995);
or U2153 (N_2153,N_1810,N_1862);
nor U2154 (N_2154,N_1948,N_1931);
or U2155 (N_2155,N_1974,N_1811);
and U2156 (N_2156,N_1964,N_1986);
or U2157 (N_2157,N_1903,N_1918);
nand U2158 (N_2158,N_1955,N_1976);
nor U2159 (N_2159,N_1942,N_1977);
nor U2160 (N_2160,N_1965,N_1899);
nor U2161 (N_2161,N_1839,N_1928);
xnor U2162 (N_2162,N_1835,N_1947);
and U2163 (N_2163,N_1873,N_1861);
nor U2164 (N_2164,N_1830,N_1867);
nor U2165 (N_2165,N_1966,N_1928);
nand U2166 (N_2166,N_1862,N_1823);
and U2167 (N_2167,N_1971,N_1993);
or U2168 (N_2168,N_1972,N_1875);
or U2169 (N_2169,N_1833,N_1808);
or U2170 (N_2170,N_1821,N_1841);
nor U2171 (N_2171,N_1821,N_1950);
and U2172 (N_2172,N_1956,N_1817);
or U2173 (N_2173,N_1909,N_1910);
nor U2174 (N_2174,N_1958,N_1840);
and U2175 (N_2175,N_1942,N_1816);
or U2176 (N_2176,N_1997,N_1904);
xor U2177 (N_2177,N_1950,N_1905);
nand U2178 (N_2178,N_1890,N_1828);
or U2179 (N_2179,N_1933,N_1890);
nor U2180 (N_2180,N_1964,N_1924);
or U2181 (N_2181,N_1858,N_1881);
or U2182 (N_2182,N_1984,N_1824);
nor U2183 (N_2183,N_1932,N_1933);
and U2184 (N_2184,N_1874,N_1844);
nand U2185 (N_2185,N_1996,N_1914);
and U2186 (N_2186,N_1824,N_1968);
or U2187 (N_2187,N_1920,N_1928);
xnor U2188 (N_2188,N_1849,N_1862);
nand U2189 (N_2189,N_1892,N_1873);
or U2190 (N_2190,N_1984,N_1808);
or U2191 (N_2191,N_1974,N_1897);
nand U2192 (N_2192,N_1986,N_1925);
nand U2193 (N_2193,N_1894,N_1984);
nor U2194 (N_2194,N_1848,N_1963);
and U2195 (N_2195,N_1987,N_1997);
and U2196 (N_2196,N_1900,N_1891);
and U2197 (N_2197,N_1962,N_1919);
or U2198 (N_2198,N_1948,N_1880);
or U2199 (N_2199,N_1808,N_1968);
nor U2200 (N_2200,N_2011,N_2002);
nor U2201 (N_2201,N_2054,N_2154);
nor U2202 (N_2202,N_2185,N_2194);
or U2203 (N_2203,N_2089,N_2127);
and U2204 (N_2204,N_2019,N_2048);
and U2205 (N_2205,N_2016,N_2168);
and U2206 (N_2206,N_2085,N_2138);
nand U2207 (N_2207,N_2001,N_2075);
or U2208 (N_2208,N_2195,N_2040);
nor U2209 (N_2209,N_2162,N_2056);
nor U2210 (N_2210,N_2028,N_2047);
or U2211 (N_2211,N_2009,N_2081);
nand U2212 (N_2212,N_2037,N_2105);
or U2213 (N_2213,N_2083,N_2036);
xnor U2214 (N_2214,N_2023,N_2114);
xor U2215 (N_2215,N_2174,N_2058);
nand U2216 (N_2216,N_2147,N_2141);
nand U2217 (N_2217,N_2169,N_2070);
or U2218 (N_2218,N_2167,N_2156);
nand U2219 (N_2219,N_2178,N_2007);
or U2220 (N_2220,N_2066,N_2181);
and U2221 (N_2221,N_2175,N_2038);
nor U2222 (N_2222,N_2145,N_2057);
nor U2223 (N_2223,N_2015,N_2000);
and U2224 (N_2224,N_2088,N_2098);
nand U2225 (N_2225,N_2163,N_2152);
and U2226 (N_2226,N_2123,N_2031);
nor U2227 (N_2227,N_2153,N_2193);
nand U2228 (N_2228,N_2026,N_2133);
and U2229 (N_2229,N_2039,N_2188);
and U2230 (N_2230,N_2155,N_2130);
nand U2231 (N_2231,N_2131,N_2069);
or U2232 (N_2232,N_2139,N_2021);
nand U2233 (N_2233,N_2120,N_2003);
and U2234 (N_2234,N_2022,N_2191);
nand U2235 (N_2235,N_2074,N_2182);
or U2236 (N_2236,N_2080,N_2055);
or U2237 (N_2237,N_2136,N_2128);
nor U2238 (N_2238,N_2198,N_2045);
or U2239 (N_2239,N_2052,N_2084);
or U2240 (N_2240,N_2125,N_2094);
or U2241 (N_2241,N_2116,N_2041);
and U2242 (N_2242,N_2097,N_2192);
nor U2243 (N_2243,N_2106,N_2095);
nor U2244 (N_2244,N_2183,N_2100);
nor U2245 (N_2245,N_2060,N_2117);
and U2246 (N_2246,N_2137,N_2112);
or U2247 (N_2247,N_2024,N_2101);
and U2248 (N_2248,N_2046,N_2176);
or U2249 (N_2249,N_2018,N_2146);
nor U2250 (N_2250,N_2108,N_2087);
and U2251 (N_2251,N_2160,N_2115);
nand U2252 (N_2252,N_2171,N_2149);
and U2253 (N_2253,N_2032,N_2025);
nor U2254 (N_2254,N_2014,N_2006);
or U2255 (N_2255,N_2049,N_2170);
and U2256 (N_2256,N_2102,N_2068);
or U2257 (N_2257,N_2118,N_2093);
or U2258 (N_2258,N_2079,N_2113);
nor U2259 (N_2259,N_2065,N_2062);
nor U2260 (N_2260,N_2142,N_2059);
and U2261 (N_2261,N_2042,N_2148);
or U2262 (N_2262,N_2135,N_2179);
and U2263 (N_2263,N_2186,N_2050);
nand U2264 (N_2264,N_2110,N_2073);
nand U2265 (N_2265,N_2035,N_2122);
nand U2266 (N_2266,N_2027,N_2103);
and U2267 (N_2267,N_2033,N_2099);
nor U2268 (N_2268,N_2067,N_2180);
or U2269 (N_2269,N_2187,N_2020);
and U2270 (N_2270,N_2177,N_2132);
nand U2271 (N_2271,N_2034,N_2017);
and U2272 (N_2272,N_2077,N_2082);
nand U2273 (N_2273,N_2064,N_2159);
nand U2274 (N_2274,N_2008,N_2165);
and U2275 (N_2275,N_2109,N_2030);
and U2276 (N_2276,N_2119,N_2121);
and U2277 (N_2277,N_2190,N_2053);
nand U2278 (N_2278,N_2004,N_2072);
nand U2279 (N_2279,N_2129,N_2158);
nand U2280 (N_2280,N_2164,N_2071);
and U2281 (N_2281,N_2090,N_2029);
or U2282 (N_2282,N_2124,N_2086);
nor U2283 (N_2283,N_2173,N_2076);
nand U2284 (N_2284,N_2012,N_2140);
nand U2285 (N_2285,N_2189,N_2107);
nand U2286 (N_2286,N_2134,N_2144);
nor U2287 (N_2287,N_2197,N_2091);
and U2288 (N_2288,N_2013,N_2161);
or U2289 (N_2289,N_2051,N_2092);
nor U2290 (N_2290,N_2126,N_2044);
or U2291 (N_2291,N_2111,N_2096);
nor U2292 (N_2292,N_2043,N_2184);
nor U2293 (N_2293,N_2150,N_2199);
or U2294 (N_2294,N_2104,N_2005);
and U2295 (N_2295,N_2143,N_2157);
or U2296 (N_2296,N_2010,N_2151);
nand U2297 (N_2297,N_2196,N_2166);
nand U2298 (N_2298,N_2061,N_2078);
or U2299 (N_2299,N_2063,N_2172);
nor U2300 (N_2300,N_2011,N_2187);
nor U2301 (N_2301,N_2112,N_2085);
nor U2302 (N_2302,N_2127,N_2054);
or U2303 (N_2303,N_2088,N_2172);
nand U2304 (N_2304,N_2189,N_2055);
nand U2305 (N_2305,N_2188,N_2098);
and U2306 (N_2306,N_2003,N_2143);
and U2307 (N_2307,N_2181,N_2140);
nand U2308 (N_2308,N_2006,N_2147);
and U2309 (N_2309,N_2122,N_2121);
nand U2310 (N_2310,N_2140,N_2032);
nand U2311 (N_2311,N_2130,N_2089);
nor U2312 (N_2312,N_2115,N_2067);
and U2313 (N_2313,N_2056,N_2075);
and U2314 (N_2314,N_2035,N_2169);
and U2315 (N_2315,N_2179,N_2043);
or U2316 (N_2316,N_2086,N_2166);
nand U2317 (N_2317,N_2001,N_2033);
nand U2318 (N_2318,N_2062,N_2140);
and U2319 (N_2319,N_2158,N_2124);
or U2320 (N_2320,N_2122,N_2147);
and U2321 (N_2321,N_2163,N_2167);
nand U2322 (N_2322,N_2048,N_2191);
nand U2323 (N_2323,N_2056,N_2199);
and U2324 (N_2324,N_2192,N_2160);
nand U2325 (N_2325,N_2068,N_2143);
nor U2326 (N_2326,N_2033,N_2164);
nor U2327 (N_2327,N_2159,N_2004);
or U2328 (N_2328,N_2069,N_2024);
nand U2329 (N_2329,N_2073,N_2037);
and U2330 (N_2330,N_2164,N_2119);
and U2331 (N_2331,N_2178,N_2063);
and U2332 (N_2332,N_2061,N_2051);
or U2333 (N_2333,N_2035,N_2148);
and U2334 (N_2334,N_2088,N_2045);
or U2335 (N_2335,N_2060,N_2183);
or U2336 (N_2336,N_2046,N_2061);
nand U2337 (N_2337,N_2131,N_2138);
nor U2338 (N_2338,N_2130,N_2073);
nor U2339 (N_2339,N_2173,N_2019);
nor U2340 (N_2340,N_2077,N_2075);
nand U2341 (N_2341,N_2068,N_2161);
or U2342 (N_2342,N_2199,N_2109);
or U2343 (N_2343,N_2151,N_2183);
nor U2344 (N_2344,N_2017,N_2058);
nor U2345 (N_2345,N_2043,N_2004);
nor U2346 (N_2346,N_2024,N_2034);
nand U2347 (N_2347,N_2132,N_2191);
nand U2348 (N_2348,N_2165,N_2036);
and U2349 (N_2349,N_2194,N_2125);
nor U2350 (N_2350,N_2026,N_2040);
nor U2351 (N_2351,N_2141,N_2144);
nor U2352 (N_2352,N_2085,N_2081);
and U2353 (N_2353,N_2107,N_2020);
nand U2354 (N_2354,N_2086,N_2125);
and U2355 (N_2355,N_2152,N_2105);
and U2356 (N_2356,N_2162,N_2186);
or U2357 (N_2357,N_2103,N_2149);
or U2358 (N_2358,N_2015,N_2063);
or U2359 (N_2359,N_2073,N_2135);
nand U2360 (N_2360,N_2019,N_2172);
and U2361 (N_2361,N_2086,N_2049);
nand U2362 (N_2362,N_2041,N_2039);
nand U2363 (N_2363,N_2091,N_2171);
nor U2364 (N_2364,N_2143,N_2066);
and U2365 (N_2365,N_2118,N_2199);
or U2366 (N_2366,N_2181,N_2012);
nor U2367 (N_2367,N_2062,N_2072);
and U2368 (N_2368,N_2089,N_2195);
or U2369 (N_2369,N_2049,N_2051);
nor U2370 (N_2370,N_2176,N_2173);
or U2371 (N_2371,N_2064,N_2168);
and U2372 (N_2372,N_2175,N_2132);
nand U2373 (N_2373,N_2129,N_2197);
and U2374 (N_2374,N_2030,N_2128);
nor U2375 (N_2375,N_2006,N_2049);
and U2376 (N_2376,N_2096,N_2131);
nand U2377 (N_2377,N_2100,N_2133);
nor U2378 (N_2378,N_2038,N_2018);
nand U2379 (N_2379,N_2063,N_2113);
nand U2380 (N_2380,N_2137,N_2010);
or U2381 (N_2381,N_2192,N_2181);
or U2382 (N_2382,N_2013,N_2086);
nand U2383 (N_2383,N_2072,N_2006);
nor U2384 (N_2384,N_2112,N_2076);
and U2385 (N_2385,N_2127,N_2148);
or U2386 (N_2386,N_2180,N_2086);
nor U2387 (N_2387,N_2196,N_2107);
nor U2388 (N_2388,N_2061,N_2055);
xnor U2389 (N_2389,N_2101,N_2157);
and U2390 (N_2390,N_2152,N_2145);
nor U2391 (N_2391,N_2039,N_2077);
nor U2392 (N_2392,N_2002,N_2178);
nand U2393 (N_2393,N_2046,N_2002);
xor U2394 (N_2394,N_2118,N_2097);
or U2395 (N_2395,N_2164,N_2123);
nand U2396 (N_2396,N_2071,N_2041);
or U2397 (N_2397,N_2009,N_2149);
nor U2398 (N_2398,N_2055,N_2171);
nand U2399 (N_2399,N_2107,N_2054);
xnor U2400 (N_2400,N_2391,N_2383);
and U2401 (N_2401,N_2251,N_2362);
nor U2402 (N_2402,N_2379,N_2228);
nand U2403 (N_2403,N_2217,N_2336);
nor U2404 (N_2404,N_2222,N_2308);
nor U2405 (N_2405,N_2244,N_2320);
and U2406 (N_2406,N_2325,N_2381);
nand U2407 (N_2407,N_2343,N_2385);
nor U2408 (N_2408,N_2395,N_2327);
or U2409 (N_2409,N_2278,N_2234);
or U2410 (N_2410,N_2282,N_2322);
nand U2411 (N_2411,N_2269,N_2202);
or U2412 (N_2412,N_2214,N_2271);
nand U2413 (N_2413,N_2352,N_2287);
or U2414 (N_2414,N_2306,N_2293);
or U2415 (N_2415,N_2297,N_2284);
or U2416 (N_2416,N_2241,N_2212);
or U2417 (N_2417,N_2236,N_2230);
nand U2418 (N_2418,N_2210,N_2305);
nor U2419 (N_2419,N_2372,N_2351);
and U2420 (N_2420,N_2288,N_2220);
or U2421 (N_2421,N_2283,N_2247);
and U2422 (N_2422,N_2216,N_2356);
nand U2423 (N_2423,N_2359,N_2295);
and U2424 (N_2424,N_2317,N_2258);
or U2425 (N_2425,N_2279,N_2393);
or U2426 (N_2426,N_2355,N_2272);
and U2427 (N_2427,N_2350,N_2312);
nand U2428 (N_2428,N_2201,N_2398);
and U2429 (N_2429,N_2315,N_2219);
nand U2430 (N_2430,N_2218,N_2328);
and U2431 (N_2431,N_2208,N_2231);
nor U2432 (N_2432,N_2307,N_2341);
nand U2433 (N_2433,N_2246,N_2365);
and U2434 (N_2434,N_2361,N_2239);
or U2435 (N_2435,N_2399,N_2298);
or U2436 (N_2436,N_2267,N_2285);
nand U2437 (N_2437,N_2302,N_2321);
nor U2438 (N_2438,N_2318,N_2299);
nor U2439 (N_2439,N_2252,N_2311);
and U2440 (N_2440,N_2370,N_2266);
nand U2441 (N_2441,N_2237,N_2382);
nor U2442 (N_2442,N_2274,N_2229);
nor U2443 (N_2443,N_2227,N_2215);
or U2444 (N_2444,N_2335,N_2257);
or U2445 (N_2445,N_2323,N_2289);
nand U2446 (N_2446,N_2324,N_2358);
or U2447 (N_2447,N_2316,N_2376);
nand U2448 (N_2448,N_2276,N_2373);
nand U2449 (N_2449,N_2260,N_2225);
nand U2450 (N_2450,N_2205,N_2255);
and U2451 (N_2451,N_2268,N_2243);
nor U2452 (N_2452,N_2290,N_2349);
nand U2453 (N_2453,N_2374,N_2378);
or U2454 (N_2454,N_2242,N_2347);
or U2455 (N_2455,N_2390,N_2329);
or U2456 (N_2456,N_2249,N_2334);
nor U2457 (N_2457,N_2265,N_2256);
or U2458 (N_2458,N_2338,N_2232);
nor U2459 (N_2459,N_2238,N_2348);
nor U2460 (N_2460,N_2339,N_2377);
and U2461 (N_2461,N_2332,N_2333);
nor U2462 (N_2462,N_2368,N_2363);
or U2463 (N_2463,N_2270,N_2226);
nor U2464 (N_2464,N_2342,N_2206);
nor U2465 (N_2465,N_2262,N_2345);
nor U2466 (N_2466,N_2275,N_2364);
nor U2467 (N_2467,N_2366,N_2280);
or U2468 (N_2468,N_2375,N_2207);
or U2469 (N_2469,N_2300,N_2309);
or U2470 (N_2470,N_2277,N_2397);
and U2471 (N_2471,N_2326,N_2340);
and U2472 (N_2472,N_2292,N_2254);
nand U2473 (N_2473,N_2245,N_2389);
nor U2474 (N_2474,N_2301,N_2346);
nor U2475 (N_2475,N_2394,N_2224);
nand U2476 (N_2476,N_2240,N_2367);
nand U2477 (N_2477,N_2330,N_2392);
nor U2478 (N_2478,N_2263,N_2235);
nor U2479 (N_2479,N_2369,N_2371);
or U2480 (N_2480,N_2233,N_2213);
nand U2481 (N_2481,N_2354,N_2331);
nor U2482 (N_2482,N_2380,N_2221);
and U2483 (N_2483,N_2387,N_2303);
and U2484 (N_2484,N_2259,N_2314);
nand U2485 (N_2485,N_2253,N_2360);
xnor U2486 (N_2486,N_2204,N_2223);
and U2487 (N_2487,N_2310,N_2353);
nand U2488 (N_2488,N_2203,N_2281);
xor U2489 (N_2489,N_2337,N_2209);
and U2490 (N_2490,N_2273,N_2319);
nand U2491 (N_2491,N_2304,N_2286);
or U2492 (N_2492,N_2261,N_2264);
nand U2493 (N_2493,N_2248,N_2384);
nor U2494 (N_2494,N_2313,N_2396);
nand U2495 (N_2495,N_2344,N_2357);
and U2496 (N_2496,N_2200,N_2211);
nand U2497 (N_2497,N_2388,N_2250);
nand U2498 (N_2498,N_2296,N_2291);
nor U2499 (N_2499,N_2294,N_2386);
nor U2500 (N_2500,N_2227,N_2259);
nand U2501 (N_2501,N_2308,N_2340);
or U2502 (N_2502,N_2360,N_2222);
or U2503 (N_2503,N_2320,N_2212);
nor U2504 (N_2504,N_2317,N_2356);
nor U2505 (N_2505,N_2323,N_2205);
xor U2506 (N_2506,N_2257,N_2380);
or U2507 (N_2507,N_2216,N_2394);
nand U2508 (N_2508,N_2296,N_2263);
and U2509 (N_2509,N_2349,N_2315);
nor U2510 (N_2510,N_2267,N_2302);
and U2511 (N_2511,N_2255,N_2387);
and U2512 (N_2512,N_2274,N_2307);
nor U2513 (N_2513,N_2246,N_2275);
xnor U2514 (N_2514,N_2247,N_2373);
nand U2515 (N_2515,N_2335,N_2399);
and U2516 (N_2516,N_2249,N_2387);
xnor U2517 (N_2517,N_2369,N_2342);
and U2518 (N_2518,N_2340,N_2367);
and U2519 (N_2519,N_2248,N_2243);
nand U2520 (N_2520,N_2330,N_2216);
and U2521 (N_2521,N_2297,N_2280);
nor U2522 (N_2522,N_2246,N_2349);
xor U2523 (N_2523,N_2387,N_2250);
nor U2524 (N_2524,N_2382,N_2294);
or U2525 (N_2525,N_2390,N_2357);
and U2526 (N_2526,N_2330,N_2249);
nand U2527 (N_2527,N_2231,N_2247);
nand U2528 (N_2528,N_2391,N_2212);
and U2529 (N_2529,N_2364,N_2210);
nand U2530 (N_2530,N_2230,N_2360);
or U2531 (N_2531,N_2233,N_2250);
nand U2532 (N_2532,N_2283,N_2330);
nor U2533 (N_2533,N_2279,N_2378);
nor U2534 (N_2534,N_2287,N_2311);
and U2535 (N_2535,N_2346,N_2245);
and U2536 (N_2536,N_2335,N_2269);
nand U2537 (N_2537,N_2301,N_2295);
nor U2538 (N_2538,N_2231,N_2337);
nand U2539 (N_2539,N_2231,N_2278);
nand U2540 (N_2540,N_2260,N_2277);
nand U2541 (N_2541,N_2261,N_2347);
nand U2542 (N_2542,N_2246,N_2297);
nor U2543 (N_2543,N_2368,N_2357);
nand U2544 (N_2544,N_2237,N_2376);
nand U2545 (N_2545,N_2282,N_2346);
nor U2546 (N_2546,N_2261,N_2236);
nor U2547 (N_2547,N_2359,N_2331);
nor U2548 (N_2548,N_2370,N_2200);
nand U2549 (N_2549,N_2328,N_2268);
nor U2550 (N_2550,N_2395,N_2200);
and U2551 (N_2551,N_2207,N_2237);
or U2552 (N_2552,N_2363,N_2340);
nor U2553 (N_2553,N_2257,N_2363);
and U2554 (N_2554,N_2251,N_2386);
nor U2555 (N_2555,N_2233,N_2248);
or U2556 (N_2556,N_2233,N_2288);
nor U2557 (N_2557,N_2348,N_2388);
or U2558 (N_2558,N_2273,N_2363);
nor U2559 (N_2559,N_2232,N_2373);
or U2560 (N_2560,N_2249,N_2388);
nand U2561 (N_2561,N_2338,N_2243);
or U2562 (N_2562,N_2302,N_2345);
and U2563 (N_2563,N_2325,N_2292);
or U2564 (N_2564,N_2303,N_2250);
and U2565 (N_2565,N_2285,N_2355);
nand U2566 (N_2566,N_2276,N_2305);
or U2567 (N_2567,N_2337,N_2225);
nand U2568 (N_2568,N_2263,N_2342);
nand U2569 (N_2569,N_2329,N_2228);
or U2570 (N_2570,N_2285,N_2254);
or U2571 (N_2571,N_2325,N_2315);
nor U2572 (N_2572,N_2234,N_2211);
nor U2573 (N_2573,N_2370,N_2337);
nand U2574 (N_2574,N_2292,N_2243);
nand U2575 (N_2575,N_2390,N_2395);
nor U2576 (N_2576,N_2347,N_2325);
or U2577 (N_2577,N_2237,N_2203);
or U2578 (N_2578,N_2299,N_2397);
and U2579 (N_2579,N_2334,N_2346);
nand U2580 (N_2580,N_2313,N_2200);
nor U2581 (N_2581,N_2205,N_2272);
nor U2582 (N_2582,N_2248,N_2271);
or U2583 (N_2583,N_2371,N_2213);
nand U2584 (N_2584,N_2276,N_2335);
and U2585 (N_2585,N_2287,N_2260);
nor U2586 (N_2586,N_2263,N_2369);
or U2587 (N_2587,N_2276,N_2384);
and U2588 (N_2588,N_2221,N_2230);
nor U2589 (N_2589,N_2329,N_2356);
nor U2590 (N_2590,N_2398,N_2373);
and U2591 (N_2591,N_2396,N_2384);
or U2592 (N_2592,N_2338,N_2278);
and U2593 (N_2593,N_2366,N_2393);
nor U2594 (N_2594,N_2223,N_2210);
or U2595 (N_2595,N_2388,N_2299);
and U2596 (N_2596,N_2394,N_2240);
and U2597 (N_2597,N_2399,N_2349);
and U2598 (N_2598,N_2331,N_2270);
nand U2599 (N_2599,N_2234,N_2363);
nand U2600 (N_2600,N_2556,N_2532);
or U2601 (N_2601,N_2402,N_2422);
and U2602 (N_2602,N_2419,N_2409);
nand U2603 (N_2603,N_2491,N_2400);
or U2604 (N_2604,N_2524,N_2516);
nand U2605 (N_2605,N_2464,N_2465);
nand U2606 (N_2606,N_2561,N_2545);
nor U2607 (N_2607,N_2435,N_2505);
and U2608 (N_2608,N_2534,N_2401);
or U2609 (N_2609,N_2565,N_2560);
or U2610 (N_2610,N_2518,N_2550);
nor U2611 (N_2611,N_2544,N_2459);
or U2612 (N_2612,N_2451,N_2488);
and U2613 (N_2613,N_2474,N_2551);
or U2614 (N_2614,N_2442,N_2448);
nand U2615 (N_2615,N_2579,N_2526);
and U2616 (N_2616,N_2415,N_2509);
and U2617 (N_2617,N_2423,N_2414);
nand U2618 (N_2618,N_2520,N_2522);
nand U2619 (N_2619,N_2478,N_2500);
nand U2620 (N_2620,N_2501,N_2519);
nand U2621 (N_2621,N_2508,N_2456);
and U2622 (N_2622,N_2525,N_2429);
nand U2623 (N_2623,N_2591,N_2590);
nand U2624 (N_2624,N_2460,N_2553);
nand U2625 (N_2625,N_2572,N_2530);
or U2626 (N_2626,N_2506,N_2587);
or U2627 (N_2627,N_2425,N_2597);
or U2628 (N_2628,N_2595,N_2430);
nand U2629 (N_2629,N_2443,N_2510);
and U2630 (N_2630,N_2540,N_2535);
nand U2631 (N_2631,N_2542,N_2581);
nand U2632 (N_2632,N_2447,N_2469);
and U2633 (N_2633,N_2417,N_2571);
nand U2634 (N_2634,N_2489,N_2404);
nor U2635 (N_2635,N_2547,N_2497);
nand U2636 (N_2636,N_2521,N_2476);
nand U2637 (N_2637,N_2596,N_2405);
nand U2638 (N_2638,N_2554,N_2475);
and U2639 (N_2639,N_2586,N_2408);
and U2640 (N_2640,N_2481,N_2480);
or U2641 (N_2641,N_2453,N_2483);
or U2642 (N_2642,N_2562,N_2439);
nor U2643 (N_2643,N_2598,N_2416);
or U2644 (N_2644,N_2575,N_2445);
nor U2645 (N_2645,N_2484,N_2427);
or U2646 (N_2646,N_2428,N_2461);
or U2647 (N_2647,N_2494,N_2558);
and U2648 (N_2648,N_2503,N_2441);
and U2649 (N_2649,N_2432,N_2454);
nor U2650 (N_2650,N_2450,N_2537);
and U2651 (N_2651,N_2436,N_2589);
nor U2652 (N_2652,N_2493,N_2463);
nor U2653 (N_2653,N_2564,N_2552);
nand U2654 (N_2654,N_2411,N_2559);
nand U2655 (N_2655,N_2594,N_2468);
nand U2656 (N_2656,N_2569,N_2502);
or U2657 (N_2657,N_2437,N_2573);
and U2658 (N_2658,N_2473,N_2549);
nand U2659 (N_2659,N_2444,N_2574);
or U2660 (N_2660,N_2511,N_2563);
or U2661 (N_2661,N_2539,N_2536);
nand U2662 (N_2662,N_2514,N_2543);
nor U2663 (N_2663,N_2566,N_2455);
or U2664 (N_2664,N_2548,N_2583);
and U2665 (N_2665,N_2407,N_2434);
or U2666 (N_2666,N_2541,N_2496);
nor U2667 (N_2667,N_2527,N_2438);
and U2668 (N_2668,N_2412,N_2466);
or U2669 (N_2669,N_2578,N_2467);
and U2670 (N_2670,N_2470,N_2458);
nor U2671 (N_2671,N_2504,N_2570);
and U2672 (N_2672,N_2406,N_2431);
or U2673 (N_2673,N_2515,N_2592);
nor U2674 (N_2674,N_2528,N_2420);
or U2675 (N_2675,N_2477,N_2580);
xnor U2676 (N_2676,N_2585,N_2426);
nor U2677 (N_2677,N_2499,N_2584);
nand U2678 (N_2678,N_2449,N_2588);
and U2679 (N_2679,N_2421,N_2567);
or U2680 (N_2680,N_2568,N_2582);
nor U2681 (N_2681,N_2403,N_2512);
nand U2682 (N_2682,N_2495,N_2531);
nor U2683 (N_2683,N_2471,N_2446);
or U2684 (N_2684,N_2546,N_2538);
nor U2685 (N_2685,N_2599,N_2533);
or U2686 (N_2686,N_2413,N_2517);
and U2687 (N_2687,N_2485,N_2486);
and U2688 (N_2688,N_2418,N_2523);
and U2689 (N_2689,N_2490,N_2452);
nor U2690 (N_2690,N_2507,N_2440);
and U2691 (N_2691,N_2410,N_2555);
and U2692 (N_2692,N_2482,N_2577);
nand U2693 (N_2693,N_2557,N_2492);
and U2694 (N_2694,N_2462,N_2513);
nand U2695 (N_2695,N_2529,N_2457);
or U2696 (N_2696,N_2498,N_2433);
nor U2697 (N_2697,N_2593,N_2472);
or U2698 (N_2698,N_2576,N_2424);
nand U2699 (N_2699,N_2479,N_2487);
and U2700 (N_2700,N_2559,N_2509);
or U2701 (N_2701,N_2558,N_2480);
nand U2702 (N_2702,N_2484,N_2524);
nand U2703 (N_2703,N_2514,N_2515);
nor U2704 (N_2704,N_2469,N_2598);
and U2705 (N_2705,N_2421,N_2470);
nor U2706 (N_2706,N_2563,N_2554);
or U2707 (N_2707,N_2565,N_2427);
nor U2708 (N_2708,N_2446,N_2448);
nor U2709 (N_2709,N_2472,N_2534);
nor U2710 (N_2710,N_2588,N_2597);
and U2711 (N_2711,N_2401,N_2540);
nand U2712 (N_2712,N_2517,N_2558);
nor U2713 (N_2713,N_2476,N_2487);
nor U2714 (N_2714,N_2553,N_2515);
nor U2715 (N_2715,N_2426,N_2579);
nand U2716 (N_2716,N_2457,N_2563);
nand U2717 (N_2717,N_2476,N_2413);
nand U2718 (N_2718,N_2530,N_2450);
and U2719 (N_2719,N_2518,N_2427);
or U2720 (N_2720,N_2413,N_2586);
nand U2721 (N_2721,N_2527,N_2593);
nand U2722 (N_2722,N_2519,N_2509);
and U2723 (N_2723,N_2488,N_2523);
and U2724 (N_2724,N_2504,N_2520);
nand U2725 (N_2725,N_2550,N_2507);
nand U2726 (N_2726,N_2519,N_2414);
nor U2727 (N_2727,N_2543,N_2564);
and U2728 (N_2728,N_2482,N_2506);
nor U2729 (N_2729,N_2494,N_2567);
nand U2730 (N_2730,N_2422,N_2461);
nor U2731 (N_2731,N_2504,N_2445);
or U2732 (N_2732,N_2582,N_2563);
or U2733 (N_2733,N_2488,N_2496);
and U2734 (N_2734,N_2599,N_2473);
nor U2735 (N_2735,N_2428,N_2564);
and U2736 (N_2736,N_2561,N_2472);
nor U2737 (N_2737,N_2417,N_2453);
or U2738 (N_2738,N_2545,N_2572);
or U2739 (N_2739,N_2518,N_2591);
nand U2740 (N_2740,N_2575,N_2570);
and U2741 (N_2741,N_2512,N_2439);
nor U2742 (N_2742,N_2517,N_2545);
nand U2743 (N_2743,N_2549,N_2564);
and U2744 (N_2744,N_2470,N_2560);
nor U2745 (N_2745,N_2501,N_2593);
nand U2746 (N_2746,N_2473,N_2516);
nand U2747 (N_2747,N_2597,N_2439);
nor U2748 (N_2748,N_2418,N_2531);
or U2749 (N_2749,N_2454,N_2474);
nor U2750 (N_2750,N_2418,N_2498);
or U2751 (N_2751,N_2426,N_2465);
nand U2752 (N_2752,N_2504,N_2590);
or U2753 (N_2753,N_2530,N_2477);
nor U2754 (N_2754,N_2553,N_2487);
nor U2755 (N_2755,N_2528,N_2478);
nand U2756 (N_2756,N_2565,N_2529);
nor U2757 (N_2757,N_2456,N_2594);
nand U2758 (N_2758,N_2536,N_2505);
nor U2759 (N_2759,N_2528,N_2487);
nor U2760 (N_2760,N_2522,N_2504);
nand U2761 (N_2761,N_2421,N_2496);
nor U2762 (N_2762,N_2462,N_2405);
nor U2763 (N_2763,N_2474,N_2570);
xnor U2764 (N_2764,N_2563,N_2477);
and U2765 (N_2765,N_2479,N_2417);
xnor U2766 (N_2766,N_2507,N_2545);
and U2767 (N_2767,N_2548,N_2469);
and U2768 (N_2768,N_2413,N_2498);
nor U2769 (N_2769,N_2563,N_2555);
nand U2770 (N_2770,N_2468,N_2501);
xnor U2771 (N_2771,N_2413,N_2524);
nand U2772 (N_2772,N_2572,N_2463);
and U2773 (N_2773,N_2524,N_2447);
nor U2774 (N_2774,N_2423,N_2549);
nand U2775 (N_2775,N_2405,N_2493);
nand U2776 (N_2776,N_2591,N_2494);
or U2777 (N_2777,N_2414,N_2478);
nor U2778 (N_2778,N_2493,N_2550);
nand U2779 (N_2779,N_2490,N_2598);
or U2780 (N_2780,N_2461,N_2413);
nand U2781 (N_2781,N_2585,N_2420);
nand U2782 (N_2782,N_2523,N_2407);
or U2783 (N_2783,N_2519,N_2430);
nand U2784 (N_2784,N_2496,N_2497);
or U2785 (N_2785,N_2466,N_2555);
or U2786 (N_2786,N_2415,N_2404);
or U2787 (N_2787,N_2420,N_2480);
and U2788 (N_2788,N_2521,N_2414);
and U2789 (N_2789,N_2567,N_2471);
nand U2790 (N_2790,N_2550,N_2490);
or U2791 (N_2791,N_2596,N_2418);
nor U2792 (N_2792,N_2586,N_2439);
nand U2793 (N_2793,N_2536,N_2583);
nand U2794 (N_2794,N_2470,N_2556);
nor U2795 (N_2795,N_2530,N_2447);
nor U2796 (N_2796,N_2467,N_2518);
nor U2797 (N_2797,N_2555,N_2585);
nor U2798 (N_2798,N_2494,N_2451);
xnor U2799 (N_2799,N_2555,N_2436);
or U2800 (N_2800,N_2761,N_2724);
and U2801 (N_2801,N_2737,N_2627);
and U2802 (N_2802,N_2640,N_2729);
nand U2803 (N_2803,N_2781,N_2604);
nand U2804 (N_2804,N_2658,N_2689);
nand U2805 (N_2805,N_2635,N_2657);
or U2806 (N_2806,N_2608,N_2600);
or U2807 (N_2807,N_2722,N_2676);
nand U2808 (N_2808,N_2690,N_2698);
nor U2809 (N_2809,N_2631,N_2768);
or U2810 (N_2810,N_2636,N_2672);
and U2811 (N_2811,N_2610,N_2663);
or U2812 (N_2812,N_2673,N_2692);
or U2813 (N_2813,N_2686,N_2682);
and U2814 (N_2814,N_2766,N_2638);
and U2815 (N_2815,N_2799,N_2725);
nor U2816 (N_2816,N_2785,N_2797);
and U2817 (N_2817,N_2671,N_2626);
and U2818 (N_2818,N_2650,N_2739);
or U2819 (N_2819,N_2751,N_2699);
or U2820 (N_2820,N_2648,N_2745);
and U2821 (N_2821,N_2755,N_2633);
or U2822 (N_2822,N_2717,N_2760);
or U2823 (N_2823,N_2656,N_2701);
and U2824 (N_2824,N_2696,N_2661);
or U2825 (N_2825,N_2670,N_2607);
nand U2826 (N_2826,N_2778,N_2651);
nand U2827 (N_2827,N_2779,N_2660);
nand U2828 (N_2828,N_2791,N_2728);
nand U2829 (N_2829,N_2691,N_2623);
or U2830 (N_2830,N_2617,N_2616);
nor U2831 (N_2831,N_2789,N_2795);
or U2832 (N_2832,N_2709,N_2712);
or U2833 (N_2833,N_2619,N_2652);
and U2834 (N_2834,N_2685,N_2615);
nand U2835 (N_2835,N_2622,N_2681);
and U2836 (N_2836,N_2603,N_2639);
or U2837 (N_2837,N_2787,N_2625);
nor U2838 (N_2838,N_2675,N_2783);
nand U2839 (N_2839,N_2613,N_2769);
nor U2840 (N_2840,N_2637,N_2702);
nand U2841 (N_2841,N_2777,N_2782);
nor U2842 (N_2842,N_2644,N_2684);
nand U2843 (N_2843,N_2736,N_2649);
nor U2844 (N_2844,N_2704,N_2602);
nand U2845 (N_2845,N_2764,N_2731);
and U2846 (N_2846,N_2752,N_2700);
or U2847 (N_2847,N_2723,N_2662);
and U2848 (N_2848,N_2727,N_2741);
or U2849 (N_2849,N_2746,N_2618);
or U2850 (N_2850,N_2601,N_2767);
and U2851 (N_2851,N_2611,N_2770);
and U2852 (N_2852,N_2740,N_2679);
nor U2853 (N_2853,N_2747,N_2634);
nand U2854 (N_2854,N_2655,N_2706);
and U2855 (N_2855,N_2659,N_2645);
or U2856 (N_2856,N_2757,N_2732);
or U2857 (N_2857,N_2756,N_2620);
and U2858 (N_2858,N_2776,N_2688);
and U2859 (N_2859,N_2788,N_2612);
nand U2860 (N_2860,N_2667,N_2753);
or U2861 (N_2861,N_2703,N_2668);
or U2862 (N_2862,N_2628,N_2605);
and U2863 (N_2863,N_2707,N_2718);
or U2864 (N_2864,N_2643,N_2687);
nor U2865 (N_2865,N_2646,N_2624);
or U2866 (N_2866,N_2711,N_2754);
nand U2867 (N_2867,N_2710,N_2694);
or U2868 (N_2868,N_2733,N_2748);
or U2869 (N_2869,N_2677,N_2730);
nor U2870 (N_2870,N_2715,N_2647);
and U2871 (N_2871,N_2792,N_2720);
and U2872 (N_2872,N_2784,N_2609);
nor U2873 (N_2873,N_2697,N_2775);
nor U2874 (N_2874,N_2796,N_2641);
nand U2875 (N_2875,N_2716,N_2743);
or U2876 (N_2876,N_2693,N_2678);
nor U2877 (N_2877,N_2780,N_2749);
nand U2878 (N_2878,N_2735,N_2630);
and U2879 (N_2879,N_2705,N_2744);
nand U2880 (N_2880,N_2759,N_2664);
and U2881 (N_2881,N_2653,N_2629);
and U2882 (N_2882,N_2798,N_2680);
nor U2883 (N_2883,N_2758,N_2793);
and U2884 (N_2884,N_2683,N_2674);
and U2885 (N_2885,N_2614,N_2774);
and U2886 (N_2886,N_2669,N_2742);
or U2887 (N_2887,N_2786,N_2750);
nand U2888 (N_2888,N_2714,N_2734);
or U2889 (N_2889,N_2765,N_2719);
and U2890 (N_2890,N_2666,N_2762);
nand U2891 (N_2891,N_2606,N_2713);
or U2892 (N_2892,N_2665,N_2642);
nand U2893 (N_2893,N_2794,N_2738);
nand U2894 (N_2894,N_2632,N_2790);
nor U2895 (N_2895,N_2763,N_2654);
nand U2896 (N_2896,N_2726,N_2772);
nand U2897 (N_2897,N_2773,N_2771);
nor U2898 (N_2898,N_2695,N_2721);
or U2899 (N_2899,N_2708,N_2621);
nor U2900 (N_2900,N_2774,N_2718);
or U2901 (N_2901,N_2667,N_2671);
nor U2902 (N_2902,N_2742,N_2640);
nand U2903 (N_2903,N_2743,N_2795);
or U2904 (N_2904,N_2694,N_2689);
nand U2905 (N_2905,N_2711,N_2666);
nand U2906 (N_2906,N_2602,N_2667);
and U2907 (N_2907,N_2603,N_2740);
and U2908 (N_2908,N_2768,N_2626);
and U2909 (N_2909,N_2797,N_2625);
or U2910 (N_2910,N_2651,N_2693);
and U2911 (N_2911,N_2690,N_2624);
xor U2912 (N_2912,N_2732,N_2780);
and U2913 (N_2913,N_2725,N_2750);
and U2914 (N_2914,N_2701,N_2720);
and U2915 (N_2915,N_2743,N_2722);
or U2916 (N_2916,N_2671,N_2654);
nand U2917 (N_2917,N_2655,N_2639);
nand U2918 (N_2918,N_2702,N_2771);
nor U2919 (N_2919,N_2734,N_2689);
nand U2920 (N_2920,N_2799,N_2732);
or U2921 (N_2921,N_2721,N_2718);
nor U2922 (N_2922,N_2782,N_2750);
nand U2923 (N_2923,N_2687,N_2745);
nand U2924 (N_2924,N_2607,N_2669);
nand U2925 (N_2925,N_2666,N_2631);
or U2926 (N_2926,N_2682,N_2697);
nor U2927 (N_2927,N_2641,N_2762);
or U2928 (N_2928,N_2643,N_2799);
nand U2929 (N_2929,N_2795,N_2625);
and U2930 (N_2930,N_2720,N_2762);
nor U2931 (N_2931,N_2667,N_2771);
or U2932 (N_2932,N_2796,N_2624);
nand U2933 (N_2933,N_2775,N_2638);
nand U2934 (N_2934,N_2752,N_2751);
and U2935 (N_2935,N_2743,N_2721);
nand U2936 (N_2936,N_2721,N_2770);
or U2937 (N_2937,N_2776,N_2791);
and U2938 (N_2938,N_2695,N_2629);
and U2939 (N_2939,N_2745,N_2715);
nand U2940 (N_2940,N_2636,N_2778);
nor U2941 (N_2941,N_2640,N_2607);
nor U2942 (N_2942,N_2622,N_2780);
nand U2943 (N_2943,N_2661,N_2681);
and U2944 (N_2944,N_2664,N_2617);
or U2945 (N_2945,N_2774,N_2712);
nand U2946 (N_2946,N_2730,N_2799);
or U2947 (N_2947,N_2673,N_2660);
nor U2948 (N_2948,N_2754,N_2628);
or U2949 (N_2949,N_2634,N_2715);
or U2950 (N_2950,N_2712,N_2777);
nor U2951 (N_2951,N_2612,N_2602);
nand U2952 (N_2952,N_2650,N_2610);
nor U2953 (N_2953,N_2748,N_2774);
and U2954 (N_2954,N_2635,N_2627);
and U2955 (N_2955,N_2648,N_2658);
or U2956 (N_2956,N_2729,N_2735);
nand U2957 (N_2957,N_2677,N_2634);
and U2958 (N_2958,N_2679,N_2782);
and U2959 (N_2959,N_2729,N_2717);
or U2960 (N_2960,N_2790,N_2785);
nor U2961 (N_2961,N_2767,N_2652);
nand U2962 (N_2962,N_2614,N_2613);
and U2963 (N_2963,N_2678,N_2618);
or U2964 (N_2964,N_2734,N_2765);
xnor U2965 (N_2965,N_2759,N_2661);
nand U2966 (N_2966,N_2654,N_2647);
and U2967 (N_2967,N_2656,N_2684);
or U2968 (N_2968,N_2755,N_2646);
and U2969 (N_2969,N_2729,N_2688);
or U2970 (N_2970,N_2753,N_2675);
and U2971 (N_2971,N_2756,N_2681);
or U2972 (N_2972,N_2750,N_2766);
and U2973 (N_2973,N_2708,N_2692);
or U2974 (N_2974,N_2678,N_2798);
nor U2975 (N_2975,N_2663,N_2799);
or U2976 (N_2976,N_2606,N_2766);
nand U2977 (N_2977,N_2765,N_2608);
nand U2978 (N_2978,N_2782,N_2793);
or U2979 (N_2979,N_2785,N_2740);
or U2980 (N_2980,N_2688,N_2702);
nand U2981 (N_2981,N_2654,N_2747);
nor U2982 (N_2982,N_2667,N_2608);
or U2983 (N_2983,N_2699,N_2797);
nor U2984 (N_2984,N_2747,N_2764);
nor U2985 (N_2985,N_2705,N_2686);
and U2986 (N_2986,N_2661,N_2658);
nand U2987 (N_2987,N_2673,N_2759);
nor U2988 (N_2988,N_2607,N_2697);
and U2989 (N_2989,N_2753,N_2608);
or U2990 (N_2990,N_2656,N_2779);
or U2991 (N_2991,N_2609,N_2698);
nor U2992 (N_2992,N_2708,N_2779);
nand U2993 (N_2993,N_2682,N_2707);
nand U2994 (N_2994,N_2676,N_2741);
or U2995 (N_2995,N_2786,N_2617);
nand U2996 (N_2996,N_2608,N_2716);
or U2997 (N_2997,N_2761,N_2706);
nand U2998 (N_2998,N_2678,N_2630);
nand U2999 (N_2999,N_2710,N_2631);
and UO_0 (O_0,N_2988,N_2997);
nor UO_1 (O_1,N_2951,N_2991);
xnor UO_2 (O_2,N_2969,N_2865);
nor UO_3 (O_3,N_2854,N_2968);
or UO_4 (O_4,N_2814,N_2842);
and UO_5 (O_5,N_2879,N_2850);
nor UO_6 (O_6,N_2931,N_2994);
nand UO_7 (O_7,N_2928,N_2880);
nor UO_8 (O_8,N_2885,N_2985);
nor UO_9 (O_9,N_2826,N_2904);
nand UO_10 (O_10,N_2962,N_2851);
and UO_11 (O_11,N_2906,N_2803);
nor UO_12 (O_12,N_2903,N_2907);
nor UO_13 (O_13,N_2864,N_2832);
nor UO_14 (O_14,N_2897,N_2943);
or UO_15 (O_15,N_2805,N_2810);
nor UO_16 (O_16,N_2986,N_2960);
and UO_17 (O_17,N_2957,N_2873);
nor UO_18 (O_18,N_2866,N_2937);
or UO_19 (O_19,N_2976,N_2820);
or UO_20 (O_20,N_2990,N_2902);
nand UO_21 (O_21,N_2899,N_2895);
and UO_22 (O_22,N_2843,N_2953);
and UO_23 (O_23,N_2952,N_2927);
or UO_24 (O_24,N_2966,N_2970);
nor UO_25 (O_25,N_2901,N_2972);
nand UO_26 (O_26,N_2930,N_2841);
nor UO_27 (O_27,N_2961,N_2973);
nor UO_28 (O_28,N_2905,N_2827);
nor UO_29 (O_29,N_2975,N_2844);
nand UO_30 (O_30,N_2861,N_2913);
xnor UO_31 (O_31,N_2878,N_2802);
nor UO_32 (O_32,N_2889,N_2932);
and UO_33 (O_33,N_2979,N_2918);
nor UO_34 (O_34,N_2910,N_2884);
or UO_35 (O_35,N_2870,N_2967);
or UO_36 (O_36,N_2817,N_2806);
or UO_37 (O_37,N_2888,N_2944);
nand UO_38 (O_38,N_2893,N_2881);
or UO_39 (O_39,N_2971,N_2845);
nand UO_40 (O_40,N_2922,N_2894);
nor UO_41 (O_41,N_2896,N_2846);
and UO_42 (O_42,N_2950,N_2874);
nor UO_43 (O_43,N_2812,N_2933);
nand UO_44 (O_44,N_2839,N_2956);
or UO_45 (O_45,N_2987,N_2958);
and UO_46 (O_46,N_2929,N_2942);
nand UO_47 (O_47,N_2816,N_2995);
and UO_48 (O_48,N_2886,N_2916);
xnor UO_49 (O_49,N_2871,N_2811);
and UO_50 (O_50,N_2852,N_2813);
nand UO_51 (O_51,N_2829,N_2882);
or UO_52 (O_52,N_2868,N_2984);
nor UO_53 (O_53,N_2980,N_2921);
nand UO_54 (O_54,N_2911,N_2831);
nor UO_55 (O_55,N_2949,N_2848);
and UO_56 (O_56,N_2822,N_2989);
nand UO_57 (O_57,N_2982,N_2856);
and UO_58 (O_58,N_2858,N_2996);
and UO_59 (O_59,N_2946,N_2919);
or UO_60 (O_60,N_2925,N_2892);
or UO_61 (O_61,N_2837,N_2804);
and UO_62 (O_62,N_2974,N_2876);
nor UO_63 (O_63,N_2912,N_2983);
nor UO_64 (O_64,N_2828,N_2891);
or UO_65 (O_65,N_2830,N_2887);
nor UO_66 (O_66,N_2877,N_2862);
nor UO_67 (O_67,N_2954,N_2923);
nand UO_68 (O_68,N_2908,N_2917);
nand UO_69 (O_69,N_2940,N_2964);
nor UO_70 (O_70,N_2825,N_2935);
or UO_71 (O_71,N_2898,N_2945);
nand UO_72 (O_72,N_2847,N_2875);
nand UO_73 (O_73,N_2924,N_2938);
nor UO_74 (O_74,N_2836,N_2872);
nand UO_75 (O_75,N_2939,N_2978);
nor UO_76 (O_76,N_2883,N_2840);
and UO_77 (O_77,N_2992,N_2819);
nor UO_78 (O_78,N_2909,N_2948);
or UO_79 (O_79,N_2818,N_2853);
and UO_80 (O_80,N_2807,N_2947);
or UO_81 (O_81,N_2900,N_2833);
or UO_82 (O_82,N_2955,N_2926);
and UO_83 (O_83,N_2965,N_2824);
nand UO_84 (O_84,N_2869,N_2863);
or UO_85 (O_85,N_2801,N_2860);
nand UO_86 (O_86,N_2981,N_2809);
nand UO_87 (O_87,N_2859,N_2936);
or UO_88 (O_88,N_2849,N_2959);
and UO_89 (O_89,N_2838,N_2815);
or UO_90 (O_90,N_2941,N_2808);
and UO_91 (O_91,N_2977,N_2999);
or UO_92 (O_92,N_2867,N_2834);
and UO_93 (O_93,N_2821,N_2915);
or UO_94 (O_94,N_2857,N_2914);
or UO_95 (O_95,N_2963,N_2998);
or UO_96 (O_96,N_2835,N_2890);
nor UO_97 (O_97,N_2920,N_2800);
nor UO_98 (O_98,N_2934,N_2993);
nor UO_99 (O_99,N_2855,N_2823);
nand UO_100 (O_100,N_2831,N_2899);
nand UO_101 (O_101,N_2883,N_2805);
and UO_102 (O_102,N_2859,N_2963);
nand UO_103 (O_103,N_2820,N_2993);
or UO_104 (O_104,N_2911,N_2857);
nand UO_105 (O_105,N_2865,N_2963);
or UO_106 (O_106,N_2872,N_2990);
and UO_107 (O_107,N_2945,N_2981);
nand UO_108 (O_108,N_2885,N_2852);
and UO_109 (O_109,N_2968,N_2964);
nor UO_110 (O_110,N_2896,N_2927);
nor UO_111 (O_111,N_2903,N_2983);
and UO_112 (O_112,N_2953,N_2812);
nand UO_113 (O_113,N_2838,N_2893);
xor UO_114 (O_114,N_2914,N_2818);
and UO_115 (O_115,N_2835,N_2830);
nand UO_116 (O_116,N_2845,N_2909);
nand UO_117 (O_117,N_2904,N_2885);
nor UO_118 (O_118,N_2915,N_2914);
and UO_119 (O_119,N_2845,N_2981);
and UO_120 (O_120,N_2818,N_2820);
or UO_121 (O_121,N_2837,N_2927);
nand UO_122 (O_122,N_2886,N_2852);
or UO_123 (O_123,N_2967,N_2975);
or UO_124 (O_124,N_2848,N_2999);
and UO_125 (O_125,N_2968,N_2922);
nand UO_126 (O_126,N_2942,N_2919);
nand UO_127 (O_127,N_2997,N_2803);
or UO_128 (O_128,N_2868,N_2806);
nor UO_129 (O_129,N_2869,N_2819);
or UO_130 (O_130,N_2998,N_2833);
nor UO_131 (O_131,N_2971,N_2854);
nand UO_132 (O_132,N_2853,N_2858);
or UO_133 (O_133,N_2897,N_2908);
and UO_134 (O_134,N_2974,N_2918);
and UO_135 (O_135,N_2857,N_2848);
nor UO_136 (O_136,N_2918,N_2881);
nand UO_137 (O_137,N_2965,N_2967);
or UO_138 (O_138,N_2898,N_2821);
nor UO_139 (O_139,N_2944,N_2829);
nand UO_140 (O_140,N_2884,N_2923);
nor UO_141 (O_141,N_2911,N_2890);
nor UO_142 (O_142,N_2830,N_2882);
or UO_143 (O_143,N_2986,N_2825);
xnor UO_144 (O_144,N_2973,N_2970);
nor UO_145 (O_145,N_2894,N_2888);
nand UO_146 (O_146,N_2807,N_2905);
or UO_147 (O_147,N_2952,N_2877);
nor UO_148 (O_148,N_2926,N_2961);
or UO_149 (O_149,N_2845,N_2924);
and UO_150 (O_150,N_2921,N_2835);
and UO_151 (O_151,N_2894,N_2910);
nand UO_152 (O_152,N_2916,N_2908);
nor UO_153 (O_153,N_2962,N_2877);
nand UO_154 (O_154,N_2944,N_2988);
nor UO_155 (O_155,N_2928,N_2819);
nor UO_156 (O_156,N_2874,N_2945);
nand UO_157 (O_157,N_2962,N_2871);
and UO_158 (O_158,N_2836,N_2952);
nand UO_159 (O_159,N_2851,N_2854);
nor UO_160 (O_160,N_2981,N_2953);
nand UO_161 (O_161,N_2807,N_2857);
or UO_162 (O_162,N_2899,N_2911);
nor UO_163 (O_163,N_2945,N_2802);
nand UO_164 (O_164,N_2865,N_2835);
nand UO_165 (O_165,N_2881,N_2941);
nor UO_166 (O_166,N_2922,N_2931);
nor UO_167 (O_167,N_2929,N_2814);
nand UO_168 (O_168,N_2911,N_2933);
and UO_169 (O_169,N_2885,N_2838);
or UO_170 (O_170,N_2891,N_2898);
and UO_171 (O_171,N_2845,N_2926);
nand UO_172 (O_172,N_2865,N_2930);
and UO_173 (O_173,N_2878,N_2910);
nor UO_174 (O_174,N_2854,N_2802);
nor UO_175 (O_175,N_2961,N_2841);
or UO_176 (O_176,N_2965,N_2895);
nor UO_177 (O_177,N_2894,N_2861);
and UO_178 (O_178,N_2970,N_2944);
or UO_179 (O_179,N_2840,N_2901);
nand UO_180 (O_180,N_2918,N_2831);
nand UO_181 (O_181,N_2816,N_2862);
and UO_182 (O_182,N_2865,N_2809);
and UO_183 (O_183,N_2956,N_2814);
nor UO_184 (O_184,N_2822,N_2987);
and UO_185 (O_185,N_2851,N_2874);
or UO_186 (O_186,N_2843,N_2814);
nand UO_187 (O_187,N_2910,N_2843);
or UO_188 (O_188,N_2840,N_2972);
and UO_189 (O_189,N_2832,N_2952);
nand UO_190 (O_190,N_2815,N_2875);
or UO_191 (O_191,N_2988,N_2855);
nor UO_192 (O_192,N_2865,N_2881);
or UO_193 (O_193,N_2986,N_2812);
and UO_194 (O_194,N_2946,N_2986);
or UO_195 (O_195,N_2912,N_2964);
nand UO_196 (O_196,N_2847,N_2942);
nor UO_197 (O_197,N_2826,N_2919);
and UO_198 (O_198,N_2860,N_2880);
nor UO_199 (O_199,N_2865,N_2806);
and UO_200 (O_200,N_2900,N_2987);
nand UO_201 (O_201,N_2914,N_2918);
or UO_202 (O_202,N_2966,N_2876);
nand UO_203 (O_203,N_2922,N_2856);
or UO_204 (O_204,N_2898,N_2878);
or UO_205 (O_205,N_2909,N_2994);
and UO_206 (O_206,N_2830,N_2875);
or UO_207 (O_207,N_2957,N_2959);
nand UO_208 (O_208,N_2899,N_2964);
or UO_209 (O_209,N_2971,N_2949);
or UO_210 (O_210,N_2971,N_2955);
nor UO_211 (O_211,N_2808,N_2860);
or UO_212 (O_212,N_2896,N_2842);
nand UO_213 (O_213,N_2876,N_2843);
nor UO_214 (O_214,N_2881,N_2946);
and UO_215 (O_215,N_2858,N_2965);
nand UO_216 (O_216,N_2831,N_2959);
nor UO_217 (O_217,N_2883,N_2952);
nand UO_218 (O_218,N_2851,N_2967);
nand UO_219 (O_219,N_2963,N_2921);
nor UO_220 (O_220,N_2911,N_2905);
or UO_221 (O_221,N_2957,N_2818);
and UO_222 (O_222,N_2845,N_2910);
and UO_223 (O_223,N_2891,N_2847);
or UO_224 (O_224,N_2864,N_2964);
nand UO_225 (O_225,N_2833,N_2884);
or UO_226 (O_226,N_2916,N_2813);
or UO_227 (O_227,N_2976,N_2828);
and UO_228 (O_228,N_2942,N_2908);
nor UO_229 (O_229,N_2908,N_2890);
nor UO_230 (O_230,N_2802,N_2899);
and UO_231 (O_231,N_2956,N_2812);
nand UO_232 (O_232,N_2938,N_2962);
and UO_233 (O_233,N_2999,N_2891);
nand UO_234 (O_234,N_2863,N_2844);
nor UO_235 (O_235,N_2959,N_2834);
nor UO_236 (O_236,N_2862,N_2859);
and UO_237 (O_237,N_2834,N_2902);
and UO_238 (O_238,N_2801,N_2933);
nor UO_239 (O_239,N_2893,N_2803);
nand UO_240 (O_240,N_2869,N_2943);
and UO_241 (O_241,N_2853,N_2932);
nor UO_242 (O_242,N_2949,N_2840);
nand UO_243 (O_243,N_2815,N_2918);
xnor UO_244 (O_244,N_2828,N_2865);
nor UO_245 (O_245,N_2979,N_2961);
nand UO_246 (O_246,N_2886,N_2806);
nor UO_247 (O_247,N_2900,N_2890);
nor UO_248 (O_248,N_2974,N_2839);
nor UO_249 (O_249,N_2976,N_2939);
or UO_250 (O_250,N_2925,N_2936);
and UO_251 (O_251,N_2927,N_2871);
nand UO_252 (O_252,N_2912,N_2940);
or UO_253 (O_253,N_2862,N_2939);
and UO_254 (O_254,N_2999,N_2960);
nor UO_255 (O_255,N_2927,N_2973);
or UO_256 (O_256,N_2960,N_2969);
or UO_257 (O_257,N_2834,N_2842);
or UO_258 (O_258,N_2859,N_2839);
or UO_259 (O_259,N_2975,N_2987);
nor UO_260 (O_260,N_2823,N_2994);
or UO_261 (O_261,N_2852,N_2831);
nand UO_262 (O_262,N_2877,N_2979);
or UO_263 (O_263,N_2854,N_2976);
nor UO_264 (O_264,N_2996,N_2922);
and UO_265 (O_265,N_2902,N_2800);
or UO_266 (O_266,N_2972,N_2811);
nand UO_267 (O_267,N_2806,N_2846);
or UO_268 (O_268,N_2891,N_2805);
nor UO_269 (O_269,N_2881,N_2820);
nor UO_270 (O_270,N_2857,N_2829);
or UO_271 (O_271,N_2943,N_2904);
nor UO_272 (O_272,N_2993,N_2940);
and UO_273 (O_273,N_2985,N_2816);
nor UO_274 (O_274,N_2902,N_2980);
and UO_275 (O_275,N_2921,N_2912);
nor UO_276 (O_276,N_2875,N_2945);
and UO_277 (O_277,N_2815,N_2901);
or UO_278 (O_278,N_2856,N_2965);
nand UO_279 (O_279,N_2950,N_2980);
nor UO_280 (O_280,N_2951,N_2937);
nand UO_281 (O_281,N_2865,N_2841);
and UO_282 (O_282,N_2970,N_2943);
or UO_283 (O_283,N_2915,N_2814);
and UO_284 (O_284,N_2998,N_2811);
and UO_285 (O_285,N_2898,N_2877);
and UO_286 (O_286,N_2830,N_2968);
or UO_287 (O_287,N_2828,N_2859);
and UO_288 (O_288,N_2826,N_2819);
nor UO_289 (O_289,N_2918,N_2933);
nor UO_290 (O_290,N_2970,N_2984);
nand UO_291 (O_291,N_2911,N_2825);
or UO_292 (O_292,N_2887,N_2960);
nand UO_293 (O_293,N_2962,N_2933);
nand UO_294 (O_294,N_2981,N_2880);
and UO_295 (O_295,N_2955,N_2813);
nor UO_296 (O_296,N_2936,N_2991);
nor UO_297 (O_297,N_2906,N_2830);
nand UO_298 (O_298,N_2926,N_2848);
or UO_299 (O_299,N_2933,N_2803);
and UO_300 (O_300,N_2851,N_2943);
and UO_301 (O_301,N_2900,N_2845);
nor UO_302 (O_302,N_2856,N_2906);
xnor UO_303 (O_303,N_2821,N_2822);
and UO_304 (O_304,N_2814,N_2901);
or UO_305 (O_305,N_2905,N_2971);
and UO_306 (O_306,N_2811,N_2989);
nand UO_307 (O_307,N_2831,N_2815);
or UO_308 (O_308,N_2853,N_2828);
or UO_309 (O_309,N_2926,N_2806);
nor UO_310 (O_310,N_2951,N_2810);
nand UO_311 (O_311,N_2999,N_2988);
or UO_312 (O_312,N_2841,N_2830);
or UO_313 (O_313,N_2958,N_2959);
and UO_314 (O_314,N_2966,N_2988);
nand UO_315 (O_315,N_2815,N_2949);
or UO_316 (O_316,N_2858,N_2910);
and UO_317 (O_317,N_2903,N_2979);
or UO_318 (O_318,N_2823,N_2971);
and UO_319 (O_319,N_2903,N_2841);
and UO_320 (O_320,N_2832,N_2820);
nand UO_321 (O_321,N_2959,N_2942);
or UO_322 (O_322,N_2829,N_2878);
nor UO_323 (O_323,N_2892,N_2949);
nor UO_324 (O_324,N_2914,N_2920);
or UO_325 (O_325,N_2853,N_2869);
nor UO_326 (O_326,N_2921,N_2988);
and UO_327 (O_327,N_2815,N_2857);
nor UO_328 (O_328,N_2838,N_2821);
nor UO_329 (O_329,N_2876,N_2855);
and UO_330 (O_330,N_2946,N_2970);
nand UO_331 (O_331,N_2968,N_2872);
nor UO_332 (O_332,N_2908,N_2906);
or UO_333 (O_333,N_2978,N_2832);
nor UO_334 (O_334,N_2980,N_2919);
nor UO_335 (O_335,N_2923,N_2966);
or UO_336 (O_336,N_2975,N_2828);
nand UO_337 (O_337,N_2895,N_2956);
nor UO_338 (O_338,N_2850,N_2843);
and UO_339 (O_339,N_2971,N_2919);
nor UO_340 (O_340,N_2951,N_2840);
nor UO_341 (O_341,N_2884,N_2969);
nor UO_342 (O_342,N_2832,N_2835);
nand UO_343 (O_343,N_2888,N_2964);
nand UO_344 (O_344,N_2988,N_2907);
and UO_345 (O_345,N_2908,N_2861);
and UO_346 (O_346,N_2831,N_2817);
nand UO_347 (O_347,N_2955,N_2867);
and UO_348 (O_348,N_2879,N_2875);
or UO_349 (O_349,N_2812,N_2985);
and UO_350 (O_350,N_2896,N_2833);
and UO_351 (O_351,N_2862,N_2995);
and UO_352 (O_352,N_2804,N_2925);
nand UO_353 (O_353,N_2998,N_2926);
nand UO_354 (O_354,N_2960,N_2930);
and UO_355 (O_355,N_2850,N_2816);
nor UO_356 (O_356,N_2867,N_2877);
nand UO_357 (O_357,N_2835,N_2855);
nor UO_358 (O_358,N_2977,N_2857);
and UO_359 (O_359,N_2876,N_2834);
nor UO_360 (O_360,N_2827,N_2815);
nand UO_361 (O_361,N_2991,N_2814);
and UO_362 (O_362,N_2891,N_2856);
or UO_363 (O_363,N_2844,N_2906);
nand UO_364 (O_364,N_2943,N_2821);
nand UO_365 (O_365,N_2988,N_2987);
or UO_366 (O_366,N_2835,N_2996);
or UO_367 (O_367,N_2991,N_2877);
nor UO_368 (O_368,N_2924,N_2892);
nor UO_369 (O_369,N_2912,N_2939);
nand UO_370 (O_370,N_2811,N_2851);
nand UO_371 (O_371,N_2992,N_2988);
and UO_372 (O_372,N_2948,N_2897);
nand UO_373 (O_373,N_2920,N_2872);
and UO_374 (O_374,N_2979,N_2999);
and UO_375 (O_375,N_2930,N_2955);
nor UO_376 (O_376,N_2831,N_2969);
or UO_377 (O_377,N_2813,N_2856);
nor UO_378 (O_378,N_2954,N_2914);
nor UO_379 (O_379,N_2812,N_2949);
or UO_380 (O_380,N_2813,N_2800);
nand UO_381 (O_381,N_2831,N_2822);
or UO_382 (O_382,N_2899,N_2901);
and UO_383 (O_383,N_2850,N_2906);
nor UO_384 (O_384,N_2889,N_2918);
and UO_385 (O_385,N_2878,N_2897);
nand UO_386 (O_386,N_2965,N_2904);
nand UO_387 (O_387,N_2946,N_2909);
nand UO_388 (O_388,N_2980,N_2816);
nor UO_389 (O_389,N_2859,N_2892);
or UO_390 (O_390,N_2896,N_2892);
and UO_391 (O_391,N_2867,N_2809);
and UO_392 (O_392,N_2984,N_2866);
nand UO_393 (O_393,N_2925,N_2825);
or UO_394 (O_394,N_2933,N_2848);
and UO_395 (O_395,N_2924,N_2985);
nor UO_396 (O_396,N_2946,N_2913);
and UO_397 (O_397,N_2879,N_2865);
or UO_398 (O_398,N_2960,N_2828);
nor UO_399 (O_399,N_2836,N_2968);
or UO_400 (O_400,N_2889,N_2849);
and UO_401 (O_401,N_2923,N_2922);
nor UO_402 (O_402,N_2998,N_2819);
nand UO_403 (O_403,N_2852,N_2983);
nand UO_404 (O_404,N_2932,N_2921);
nor UO_405 (O_405,N_2999,N_2967);
and UO_406 (O_406,N_2975,N_2896);
or UO_407 (O_407,N_2940,N_2983);
and UO_408 (O_408,N_2958,N_2907);
nor UO_409 (O_409,N_2830,N_2986);
and UO_410 (O_410,N_2805,N_2836);
nor UO_411 (O_411,N_2821,N_2928);
nand UO_412 (O_412,N_2899,N_2992);
nor UO_413 (O_413,N_2822,N_2859);
or UO_414 (O_414,N_2915,N_2895);
or UO_415 (O_415,N_2976,N_2885);
nor UO_416 (O_416,N_2862,N_2812);
or UO_417 (O_417,N_2980,N_2874);
or UO_418 (O_418,N_2945,N_2941);
or UO_419 (O_419,N_2991,N_2824);
nor UO_420 (O_420,N_2892,N_2818);
and UO_421 (O_421,N_2824,N_2979);
and UO_422 (O_422,N_2963,N_2900);
nand UO_423 (O_423,N_2898,N_2991);
or UO_424 (O_424,N_2919,N_2809);
or UO_425 (O_425,N_2997,N_2986);
or UO_426 (O_426,N_2907,N_2924);
nand UO_427 (O_427,N_2874,N_2863);
nor UO_428 (O_428,N_2959,N_2863);
nor UO_429 (O_429,N_2947,N_2892);
nor UO_430 (O_430,N_2933,N_2872);
or UO_431 (O_431,N_2965,N_2948);
nand UO_432 (O_432,N_2818,N_2810);
nand UO_433 (O_433,N_2990,N_2888);
nand UO_434 (O_434,N_2853,N_2877);
or UO_435 (O_435,N_2909,N_2938);
nor UO_436 (O_436,N_2999,N_2837);
and UO_437 (O_437,N_2870,N_2846);
or UO_438 (O_438,N_2918,N_2978);
nor UO_439 (O_439,N_2951,N_2930);
nand UO_440 (O_440,N_2846,N_2912);
nor UO_441 (O_441,N_2868,N_2962);
nor UO_442 (O_442,N_2967,N_2957);
nor UO_443 (O_443,N_2805,N_2914);
nor UO_444 (O_444,N_2906,N_2864);
nand UO_445 (O_445,N_2910,N_2861);
nand UO_446 (O_446,N_2807,N_2941);
and UO_447 (O_447,N_2860,N_2970);
nor UO_448 (O_448,N_2891,N_2832);
nand UO_449 (O_449,N_2983,N_2812);
nor UO_450 (O_450,N_2924,N_2959);
nand UO_451 (O_451,N_2969,N_2978);
or UO_452 (O_452,N_2921,N_2926);
or UO_453 (O_453,N_2852,N_2989);
nand UO_454 (O_454,N_2942,N_2968);
or UO_455 (O_455,N_2935,N_2849);
or UO_456 (O_456,N_2928,N_2905);
nand UO_457 (O_457,N_2972,N_2834);
or UO_458 (O_458,N_2828,N_2904);
nand UO_459 (O_459,N_2903,N_2847);
or UO_460 (O_460,N_2874,N_2852);
nand UO_461 (O_461,N_2909,N_2933);
nand UO_462 (O_462,N_2834,N_2810);
nor UO_463 (O_463,N_2913,N_2959);
nor UO_464 (O_464,N_2925,N_2897);
nand UO_465 (O_465,N_2920,N_2885);
nor UO_466 (O_466,N_2806,N_2922);
or UO_467 (O_467,N_2821,N_2815);
nand UO_468 (O_468,N_2979,N_2884);
or UO_469 (O_469,N_2913,N_2836);
and UO_470 (O_470,N_2852,N_2901);
and UO_471 (O_471,N_2963,N_2880);
or UO_472 (O_472,N_2966,N_2817);
and UO_473 (O_473,N_2968,N_2871);
nor UO_474 (O_474,N_2968,N_2932);
and UO_475 (O_475,N_2928,N_2993);
and UO_476 (O_476,N_2926,N_2929);
and UO_477 (O_477,N_2922,N_2902);
and UO_478 (O_478,N_2886,N_2835);
or UO_479 (O_479,N_2962,N_2926);
nand UO_480 (O_480,N_2825,N_2930);
nand UO_481 (O_481,N_2910,N_2814);
or UO_482 (O_482,N_2837,N_2864);
or UO_483 (O_483,N_2887,N_2878);
or UO_484 (O_484,N_2924,N_2817);
and UO_485 (O_485,N_2980,N_2952);
and UO_486 (O_486,N_2924,N_2956);
or UO_487 (O_487,N_2965,N_2836);
nand UO_488 (O_488,N_2968,N_2930);
nor UO_489 (O_489,N_2900,N_2824);
and UO_490 (O_490,N_2867,N_2946);
or UO_491 (O_491,N_2992,N_2853);
nor UO_492 (O_492,N_2819,N_2923);
nor UO_493 (O_493,N_2985,N_2839);
or UO_494 (O_494,N_2835,N_2937);
and UO_495 (O_495,N_2871,N_2878);
nand UO_496 (O_496,N_2850,N_2878);
or UO_497 (O_497,N_2974,N_2938);
or UO_498 (O_498,N_2959,N_2995);
xor UO_499 (O_499,N_2924,N_2827);
endmodule