module basic_500_3000_500_50_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_32,In_13);
nand U1 (N_1,In_313,In_252);
xnor U2 (N_2,In_426,In_2);
and U3 (N_3,In_101,In_428);
and U4 (N_4,In_231,In_230);
and U5 (N_5,In_169,In_491);
nor U6 (N_6,In_0,In_353);
nor U7 (N_7,In_373,In_406);
or U8 (N_8,In_47,In_415);
nor U9 (N_9,In_223,In_298);
nand U10 (N_10,In_89,In_235);
xor U11 (N_11,In_454,In_289);
xor U12 (N_12,In_55,In_418);
nor U13 (N_13,In_149,In_268);
nand U14 (N_14,In_63,In_411);
and U15 (N_15,In_151,In_237);
and U16 (N_16,In_293,In_239);
and U17 (N_17,In_109,In_332);
nor U18 (N_18,In_20,In_163);
nor U19 (N_19,In_74,In_115);
nor U20 (N_20,In_470,In_215);
nor U21 (N_21,In_106,In_233);
and U22 (N_22,In_127,In_202);
nand U23 (N_23,In_383,In_460);
or U24 (N_24,In_262,In_108);
and U25 (N_25,In_245,In_376);
and U26 (N_26,In_93,In_322);
or U27 (N_27,In_105,In_483);
nand U28 (N_28,In_170,In_422);
xnor U29 (N_29,In_375,In_261);
or U30 (N_30,In_441,In_389);
and U31 (N_31,In_140,In_193);
or U32 (N_32,In_302,In_278);
nand U33 (N_33,In_180,In_340);
or U34 (N_34,In_338,In_33);
nand U35 (N_35,In_161,In_145);
or U36 (N_36,In_366,In_431);
and U37 (N_37,In_394,In_306);
nor U38 (N_38,In_59,In_378);
or U39 (N_39,In_22,In_143);
and U40 (N_40,In_80,In_166);
nor U41 (N_41,In_5,In_144);
nand U42 (N_42,In_232,In_294);
nor U43 (N_43,In_167,In_334);
and U44 (N_44,In_153,In_485);
nor U45 (N_45,In_317,In_410);
nand U46 (N_46,In_67,In_210);
nor U47 (N_47,In_205,In_16);
or U48 (N_48,In_444,In_323);
nand U49 (N_49,In_346,In_284);
and U50 (N_50,In_92,In_416);
or U51 (N_51,In_464,In_374);
nand U52 (N_52,In_31,In_466);
and U53 (N_53,In_94,In_489);
nor U54 (N_54,In_365,In_190);
and U55 (N_55,In_225,In_188);
and U56 (N_56,In_421,In_453);
or U57 (N_57,In_295,In_157);
nand U58 (N_58,In_120,In_456);
or U59 (N_59,In_69,In_312);
nand U60 (N_60,In_357,In_8);
or U61 (N_61,N_29,In_176);
nand U62 (N_62,In_240,In_221);
nor U63 (N_63,N_34,In_321);
nor U64 (N_64,In_222,In_164);
or U65 (N_65,In_459,In_212);
nor U66 (N_66,In_326,In_452);
nand U67 (N_67,In_427,In_354);
nor U68 (N_68,In_402,In_17);
nand U69 (N_69,In_97,In_303);
and U70 (N_70,In_76,In_341);
or U71 (N_71,In_95,In_479);
nor U72 (N_72,In_248,In_238);
nor U73 (N_73,In_247,N_46);
nand U74 (N_74,N_13,In_260);
nor U75 (N_75,In_25,In_177);
or U76 (N_76,N_43,In_49);
nor U77 (N_77,In_436,In_121);
and U78 (N_78,In_39,In_116);
or U79 (N_79,In_150,In_325);
and U80 (N_80,In_372,In_156);
xnor U81 (N_81,In_280,N_49);
nor U82 (N_82,In_276,In_184);
and U83 (N_83,In_10,In_440);
or U84 (N_84,In_496,In_327);
and U85 (N_85,In_198,In_102);
nor U86 (N_86,In_86,In_371);
or U87 (N_87,In_467,In_175);
nor U88 (N_88,In_490,In_336);
or U89 (N_89,In_12,In_152);
nand U90 (N_90,In_296,N_52);
nor U91 (N_91,In_70,In_314);
or U92 (N_92,In_301,In_348);
nor U93 (N_93,In_85,In_124);
and U94 (N_94,In_228,In_64);
nor U95 (N_95,In_409,In_253);
nor U96 (N_96,In_213,In_342);
and U97 (N_97,In_259,In_192);
nor U98 (N_98,In_83,In_291);
or U99 (N_99,In_356,In_172);
nor U100 (N_100,In_54,In_494);
nand U101 (N_101,In_424,N_15);
or U102 (N_102,In_419,In_51);
nand U103 (N_103,In_335,N_14);
or U104 (N_104,In_407,In_380);
and U105 (N_105,N_12,N_57);
nand U106 (N_106,In_495,In_52);
nand U107 (N_107,In_183,In_226);
nor U108 (N_108,In_497,In_35);
or U109 (N_109,In_279,In_448);
nand U110 (N_110,In_160,In_285);
nand U111 (N_111,In_24,In_206);
nor U112 (N_112,In_111,N_5);
or U113 (N_113,In_417,In_382);
and U114 (N_114,In_300,In_320);
nor U115 (N_115,In_36,In_242);
nor U116 (N_116,In_201,N_38);
and U117 (N_117,In_481,In_488);
or U118 (N_118,In_395,In_107);
nor U119 (N_119,In_256,In_200);
nor U120 (N_120,In_267,In_385);
nand U121 (N_121,In_360,N_85);
nor U122 (N_122,N_96,In_251);
and U123 (N_123,In_139,In_480);
nand U124 (N_124,N_4,In_412);
nand U125 (N_125,N_94,N_97);
and U126 (N_126,In_171,N_51);
or U127 (N_127,N_11,N_3);
nand U128 (N_128,N_65,In_399);
nor U129 (N_129,In_135,In_339);
nor U130 (N_130,In_71,In_297);
nand U131 (N_131,N_101,N_111);
nor U132 (N_132,N_31,In_492);
and U133 (N_133,N_114,N_79);
nand U134 (N_134,N_27,In_405);
or U135 (N_135,In_393,In_78);
xor U136 (N_136,N_19,In_103);
nor U137 (N_137,In_305,In_203);
and U138 (N_138,N_110,In_288);
or U139 (N_139,In_81,In_246);
or U140 (N_140,In_28,N_105);
or U141 (N_141,In_46,In_119);
or U142 (N_142,N_77,N_60);
nand U143 (N_143,N_68,In_182);
nand U144 (N_144,In_272,In_439);
nor U145 (N_145,N_35,N_99);
nand U146 (N_146,In_61,In_333);
or U147 (N_147,In_62,In_56);
nand U148 (N_148,In_19,In_65);
nor U149 (N_149,In_58,In_82);
nor U150 (N_150,In_110,In_162);
nor U151 (N_151,In_337,In_482);
nor U152 (N_152,In_45,In_128);
or U153 (N_153,In_462,In_7);
or U154 (N_154,In_315,In_403);
nor U155 (N_155,In_73,In_447);
and U156 (N_156,In_18,In_329);
nor U157 (N_157,In_282,N_100);
nand U158 (N_158,N_115,In_208);
or U159 (N_159,In_75,N_40);
nand U160 (N_160,In_219,In_141);
or U161 (N_161,In_361,In_344);
and U162 (N_162,In_234,In_457);
or U163 (N_163,In_487,N_21);
or U164 (N_164,In_478,N_54);
nand U165 (N_165,N_69,In_474);
or U166 (N_166,In_352,N_17);
nand U167 (N_167,In_48,In_271);
nor U168 (N_168,In_132,In_430);
nand U169 (N_169,In_189,In_493);
nor U170 (N_170,In_472,In_217);
nand U171 (N_171,In_138,In_181);
and U172 (N_172,In_324,N_88);
or U173 (N_173,In_350,N_44);
nand U174 (N_174,N_112,In_21);
nor U175 (N_175,N_22,In_290);
or U176 (N_176,N_25,N_24);
and U177 (N_177,In_429,N_10);
nor U178 (N_178,N_50,In_244);
and U179 (N_179,In_186,In_174);
nor U180 (N_180,N_59,In_434);
nor U181 (N_181,In_122,N_1);
and U182 (N_182,In_41,In_147);
and U183 (N_183,In_68,In_270);
or U184 (N_184,In_178,In_34);
and U185 (N_185,N_159,N_158);
and U186 (N_186,In_29,N_61);
and U187 (N_187,N_86,N_48);
and U188 (N_188,In_4,In_43);
and U189 (N_189,N_16,In_209);
nand U190 (N_190,N_42,N_95);
or U191 (N_191,N_125,In_194);
or U192 (N_192,In_216,In_437);
and U193 (N_193,N_179,In_1);
nand U194 (N_194,N_122,In_40);
or U195 (N_195,In_400,In_100);
and U196 (N_196,In_264,In_377);
nor U197 (N_197,N_103,N_132);
nor U198 (N_198,In_257,In_438);
or U199 (N_199,N_161,In_220);
nor U200 (N_200,N_176,N_104);
or U201 (N_201,In_158,In_218);
nor U202 (N_202,In_443,In_369);
or U203 (N_203,N_142,N_164);
nor U204 (N_204,In_465,In_258);
nand U205 (N_205,In_44,In_392);
nand U206 (N_206,N_55,N_87);
or U207 (N_207,In_53,N_137);
nand U208 (N_208,In_386,In_196);
and U209 (N_209,In_98,In_458);
or U210 (N_210,N_63,In_319);
or U211 (N_211,In_423,In_126);
and U212 (N_212,N_106,In_250);
nor U213 (N_213,N_143,In_273);
nor U214 (N_214,N_134,N_148);
and U215 (N_215,In_397,N_74);
xor U216 (N_216,In_286,In_330);
and U217 (N_217,In_299,In_207);
nor U218 (N_218,In_292,N_136);
nand U219 (N_219,In_475,In_463);
and U220 (N_220,In_137,In_351);
nor U221 (N_221,In_404,N_83);
nand U222 (N_222,N_127,N_173);
nand U223 (N_223,In_125,N_149);
or U224 (N_224,In_118,N_153);
or U225 (N_225,In_26,N_167);
nand U226 (N_226,N_108,N_157);
or U227 (N_227,N_30,N_75);
and U228 (N_228,In_249,N_6);
nand U229 (N_229,N_71,In_455);
nor U230 (N_230,N_102,In_471);
nand U231 (N_231,N_154,N_72);
nand U232 (N_232,In_287,N_168);
and U233 (N_233,N_147,N_20);
nor U234 (N_234,In_461,N_109);
or U235 (N_235,In_499,In_425);
nand U236 (N_236,In_384,N_113);
nor U237 (N_237,N_169,In_433);
nand U238 (N_238,N_172,N_36);
nor U239 (N_239,In_281,N_7);
and U240 (N_240,N_67,In_155);
xor U241 (N_241,N_209,In_476);
nor U242 (N_242,In_311,N_138);
nand U243 (N_243,In_187,N_203);
nor U244 (N_244,In_328,N_47);
or U245 (N_245,In_173,In_224);
or U246 (N_246,In_136,N_129);
and U247 (N_247,N_165,N_217);
nor U248 (N_248,N_231,N_80);
and U249 (N_249,N_175,In_129);
xnor U250 (N_250,In_42,N_214);
xor U251 (N_251,N_152,In_304);
or U252 (N_252,In_266,N_76);
or U253 (N_253,N_236,In_331);
nand U254 (N_254,In_390,In_214);
and U255 (N_255,N_118,N_205);
and U256 (N_256,In_391,In_368);
or U257 (N_257,In_381,In_30);
nand U258 (N_258,N_58,N_128);
and U259 (N_259,N_123,In_367);
and U260 (N_260,N_234,N_39);
nand U261 (N_261,In_473,N_171);
nand U262 (N_262,In_130,N_201);
and U263 (N_263,In_117,N_198);
or U264 (N_264,In_435,In_274);
nand U265 (N_265,In_195,N_41);
or U266 (N_266,N_91,N_62);
nor U267 (N_267,In_442,In_359);
and U268 (N_268,N_199,N_124);
nand U269 (N_269,In_269,N_121);
nand U270 (N_270,In_142,N_183);
and U271 (N_271,In_414,In_309);
or U272 (N_272,In_477,In_358);
or U273 (N_273,N_187,In_316);
nand U274 (N_274,In_37,N_56);
nand U275 (N_275,N_200,N_166);
and U276 (N_276,In_379,N_223);
nand U277 (N_277,In_449,In_227);
xor U278 (N_278,In_432,In_146);
nor U279 (N_279,N_117,N_120);
nand U280 (N_280,In_11,In_84);
or U281 (N_281,In_349,N_215);
or U282 (N_282,In_91,In_446);
and U283 (N_283,N_193,N_163);
nor U284 (N_284,In_451,In_486);
nand U285 (N_285,N_230,In_277);
nor U286 (N_286,In_179,N_186);
and U287 (N_287,N_84,N_98);
nand U288 (N_288,N_93,In_199);
or U289 (N_289,In_14,In_104);
nand U290 (N_290,N_227,N_216);
nand U291 (N_291,N_229,N_145);
nor U292 (N_292,N_82,N_197);
or U293 (N_293,In_362,N_177);
xnor U294 (N_294,N_81,N_218);
nor U295 (N_295,N_23,N_211);
xnor U296 (N_296,N_228,N_238);
or U297 (N_297,In_388,In_112);
nor U298 (N_298,In_72,In_204);
nand U299 (N_299,N_146,N_196);
nor U300 (N_300,In_263,N_210);
nor U301 (N_301,In_283,N_45);
nor U302 (N_302,N_206,In_343);
xnor U303 (N_303,N_73,N_254);
and U304 (N_304,N_284,In_87);
and U305 (N_305,N_8,N_194);
nand U306 (N_306,N_89,N_248);
nor U307 (N_307,N_251,N_271);
nor U308 (N_308,N_178,N_283);
nor U309 (N_309,N_277,N_92);
and U310 (N_310,N_33,In_347);
nor U311 (N_311,N_219,N_66);
and U312 (N_312,In_310,In_229);
nor U313 (N_313,N_297,In_408);
nand U314 (N_314,In_307,N_207);
or U315 (N_315,In_114,N_288);
or U316 (N_316,In_401,N_139);
nand U317 (N_317,N_2,In_96);
nand U318 (N_318,N_170,N_239);
or U319 (N_319,N_64,N_151);
nand U320 (N_320,N_220,N_293);
and U321 (N_321,In_79,N_225);
and U322 (N_322,In_318,In_148);
nand U323 (N_323,N_290,N_150);
or U324 (N_324,In_241,N_282);
and U325 (N_325,In_113,In_60);
or U326 (N_326,In_243,N_162);
nor U327 (N_327,N_237,N_272);
nor U328 (N_328,N_245,N_299);
nand U329 (N_329,N_241,N_262);
nor U330 (N_330,N_202,N_292);
xor U331 (N_331,N_26,In_197);
nor U332 (N_332,N_295,N_28);
and U333 (N_333,In_168,In_345);
nor U334 (N_334,N_235,N_213);
nor U335 (N_335,N_182,N_222);
or U336 (N_336,N_192,N_208);
nand U337 (N_337,N_133,N_298);
nor U338 (N_338,N_252,N_180);
nand U339 (N_339,N_258,In_88);
nand U340 (N_340,In_398,N_280);
and U341 (N_341,In_159,N_185);
nor U342 (N_342,N_285,In_50);
or U343 (N_343,N_131,N_244);
nand U344 (N_344,In_27,In_185);
xnor U345 (N_345,N_250,N_221);
nor U346 (N_346,N_32,N_226);
and U347 (N_347,In_191,N_184);
and U348 (N_348,N_135,In_413);
and U349 (N_349,In_364,N_281);
nand U350 (N_350,N_273,In_123);
or U351 (N_351,N_256,N_261);
or U352 (N_352,N_119,In_396);
nor U353 (N_353,N_266,In_9);
nand U354 (N_354,In_255,N_276);
or U355 (N_355,N_275,N_9);
nor U356 (N_356,N_18,In_498);
and U357 (N_357,N_191,N_286);
or U358 (N_358,N_90,N_296);
nor U359 (N_359,In_134,In_99);
and U360 (N_360,N_257,N_212);
or U361 (N_361,N_318,In_57);
nor U362 (N_362,In_468,In_90);
nor U363 (N_363,N_310,In_308);
and U364 (N_364,N_311,N_332);
nor U365 (N_365,N_309,N_204);
or U366 (N_366,N_346,N_326);
or U367 (N_367,N_263,N_337);
xor U368 (N_368,In_154,N_352);
nand U369 (N_369,N_358,N_289);
nor U370 (N_370,N_313,N_350);
nand U371 (N_371,N_316,N_156);
and U372 (N_372,N_287,N_340);
nor U373 (N_373,N_37,N_344);
nor U374 (N_374,N_307,N_351);
and U375 (N_375,In_420,N_247);
and U376 (N_376,In_265,N_356);
and U377 (N_377,N_224,In_133);
nand U378 (N_378,N_334,In_77);
nor U379 (N_379,In_254,In_15);
nand U380 (N_380,N_126,N_0);
and U381 (N_381,N_242,In_66);
and U382 (N_382,N_232,N_140);
nand U383 (N_383,N_144,N_312);
nor U384 (N_384,In_38,N_70);
nand U385 (N_385,N_347,N_53);
xor U386 (N_386,N_322,N_141);
or U387 (N_387,In_131,In_3);
and U388 (N_388,N_321,N_107);
nand U389 (N_389,N_315,N_243);
nand U390 (N_390,In_275,N_355);
nor U391 (N_391,N_188,N_274);
nor U392 (N_392,N_333,N_317);
nor U393 (N_393,N_301,N_116);
nor U394 (N_394,N_246,N_174);
nor U395 (N_395,N_328,N_339);
nand U396 (N_396,N_279,N_335);
nand U397 (N_397,N_314,N_324);
nor U398 (N_398,N_260,N_354);
and U399 (N_399,N_291,N_323);
or U400 (N_400,N_160,In_484);
nor U401 (N_401,In_450,In_211);
and U402 (N_402,N_306,N_195);
or U403 (N_403,N_181,N_327);
and U404 (N_404,N_343,N_357);
and U405 (N_405,N_342,N_345);
nor U406 (N_406,N_331,N_349);
nand U407 (N_407,N_330,N_305);
and U408 (N_408,N_338,N_264);
or U409 (N_409,N_78,In_165);
nand U410 (N_410,N_240,N_189);
and U411 (N_411,In_6,In_363);
and U412 (N_412,In_370,N_308);
and U413 (N_413,In_387,N_302);
or U414 (N_414,In_23,N_304);
and U415 (N_415,N_259,N_265);
or U416 (N_416,N_233,N_270);
nor U417 (N_417,N_359,In_445);
or U418 (N_418,N_353,N_300);
and U419 (N_419,N_341,N_336);
nor U420 (N_420,N_386,N_419);
xnor U421 (N_421,N_390,N_374);
and U422 (N_422,N_398,N_409);
nor U423 (N_423,N_408,N_377);
and U424 (N_424,N_404,N_394);
nand U425 (N_425,N_348,In_355);
or U426 (N_426,N_373,N_269);
nand U427 (N_427,N_405,N_414);
and U428 (N_428,N_411,N_389);
or U429 (N_429,N_367,N_400);
nor U430 (N_430,In_236,N_395);
nand U431 (N_431,N_416,N_294);
or U432 (N_432,N_376,N_368);
nor U433 (N_433,N_410,N_402);
or U434 (N_434,N_378,N_360);
and U435 (N_435,N_190,N_303);
and U436 (N_436,N_329,N_320);
and U437 (N_437,N_370,N_319);
xnor U438 (N_438,N_417,N_401);
nand U439 (N_439,N_325,N_249);
nor U440 (N_440,N_268,N_393);
nor U441 (N_441,N_418,N_399);
and U442 (N_442,N_364,N_371);
nor U443 (N_443,N_366,N_130);
or U444 (N_444,N_387,N_361);
or U445 (N_445,N_381,N_362);
or U446 (N_446,N_365,N_391);
nand U447 (N_447,N_406,N_375);
and U448 (N_448,N_372,N_407);
or U449 (N_449,N_155,N_385);
nor U450 (N_450,N_383,N_392);
or U451 (N_451,N_267,N_384);
and U452 (N_452,N_363,N_380);
and U453 (N_453,N_255,N_379);
or U454 (N_454,N_382,N_388);
and U455 (N_455,N_369,In_469);
and U456 (N_456,N_413,N_412);
nand U457 (N_457,N_278,N_403);
and U458 (N_458,N_253,N_415);
nand U459 (N_459,N_397,N_396);
and U460 (N_460,N_386,N_402);
and U461 (N_461,N_419,N_402);
and U462 (N_462,N_398,N_268);
nor U463 (N_463,N_408,N_392);
nand U464 (N_464,N_369,N_362);
nand U465 (N_465,N_411,N_378);
nand U466 (N_466,N_403,N_419);
xor U467 (N_467,N_399,N_249);
nor U468 (N_468,N_386,N_414);
nor U469 (N_469,N_303,N_372);
nand U470 (N_470,N_375,N_155);
and U471 (N_471,N_378,N_402);
or U472 (N_472,N_395,N_278);
and U473 (N_473,N_372,N_400);
and U474 (N_474,N_130,N_371);
or U475 (N_475,N_377,N_325);
nor U476 (N_476,N_382,N_255);
and U477 (N_477,N_390,In_355);
nor U478 (N_478,In_236,N_385);
nand U479 (N_479,N_369,N_348);
nand U480 (N_480,N_436,N_422);
or U481 (N_481,N_462,N_460);
nor U482 (N_482,N_435,N_457);
and U483 (N_483,N_431,N_439);
xnor U484 (N_484,N_474,N_456);
and U485 (N_485,N_468,N_466);
nor U486 (N_486,N_442,N_453);
nand U487 (N_487,N_424,N_441);
nand U488 (N_488,N_426,N_464);
or U489 (N_489,N_445,N_423);
or U490 (N_490,N_461,N_470);
and U491 (N_491,N_459,N_463);
and U492 (N_492,N_452,N_427);
xor U493 (N_493,N_476,N_432);
nand U494 (N_494,N_479,N_451);
or U495 (N_495,N_420,N_421);
or U496 (N_496,N_450,N_429);
nand U497 (N_497,N_446,N_472);
nor U498 (N_498,N_473,N_428);
nor U499 (N_499,N_469,N_467);
or U500 (N_500,N_425,N_438);
nor U501 (N_501,N_447,N_444);
nand U502 (N_502,N_454,N_443);
nor U503 (N_503,N_449,N_430);
nand U504 (N_504,N_478,N_433);
and U505 (N_505,N_477,N_434);
or U506 (N_506,N_458,N_437);
xor U507 (N_507,N_440,N_475);
or U508 (N_508,N_471,N_455);
xnor U509 (N_509,N_448,N_465);
xor U510 (N_510,N_465,N_429);
nor U511 (N_511,N_455,N_460);
and U512 (N_512,N_429,N_423);
nand U513 (N_513,N_462,N_429);
or U514 (N_514,N_478,N_420);
nor U515 (N_515,N_473,N_423);
or U516 (N_516,N_431,N_434);
or U517 (N_517,N_477,N_438);
nand U518 (N_518,N_438,N_474);
or U519 (N_519,N_432,N_447);
nand U520 (N_520,N_420,N_452);
or U521 (N_521,N_456,N_420);
nor U522 (N_522,N_479,N_454);
xor U523 (N_523,N_431,N_428);
or U524 (N_524,N_455,N_435);
nor U525 (N_525,N_465,N_430);
or U526 (N_526,N_423,N_420);
and U527 (N_527,N_447,N_429);
nand U528 (N_528,N_454,N_432);
nor U529 (N_529,N_439,N_473);
nand U530 (N_530,N_445,N_455);
nand U531 (N_531,N_428,N_433);
nor U532 (N_532,N_458,N_422);
xnor U533 (N_533,N_436,N_459);
and U534 (N_534,N_469,N_472);
nor U535 (N_535,N_427,N_473);
or U536 (N_536,N_469,N_434);
and U537 (N_537,N_467,N_439);
nor U538 (N_538,N_438,N_433);
and U539 (N_539,N_458,N_438);
nor U540 (N_540,N_512,N_520);
nand U541 (N_541,N_498,N_536);
nand U542 (N_542,N_504,N_484);
or U543 (N_543,N_493,N_495);
nand U544 (N_544,N_534,N_516);
and U545 (N_545,N_481,N_480);
nand U546 (N_546,N_527,N_509);
and U547 (N_547,N_526,N_502);
nand U548 (N_548,N_496,N_517);
nand U549 (N_549,N_490,N_497);
and U550 (N_550,N_486,N_488);
and U551 (N_551,N_503,N_494);
or U552 (N_552,N_500,N_514);
and U553 (N_553,N_524,N_532);
nor U554 (N_554,N_507,N_506);
nand U555 (N_555,N_528,N_533);
or U556 (N_556,N_499,N_539);
or U557 (N_557,N_522,N_531);
or U558 (N_558,N_492,N_483);
and U559 (N_559,N_511,N_538);
xor U560 (N_560,N_487,N_535);
or U561 (N_561,N_525,N_501);
nor U562 (N_562,N_523,N_489);
or U563 (N_563,N_529,N_530);
nand U564 (N_564,N_510,N_491);
and U565 (N_565,N_537,N_521);
or U566 (N_566,N_518,N_508);
and U567 (N_567,N_505,N_519);
or U568 (N_568,N_482,N_513);
xor U569 (N_569,N_485,N_515);
nand U570 (N_570,N_521,N_512);
and U571 (N_571,N_531,N_486);
and U572 (N_572,N_533,N_523);
or U573 (N_573,N_492,N_518);
xor U574 (N_574,N_511,N_527);
or U575 (N_575,N_539,N_497);
nand U576 (N_576,N_480,N_504);
nor U577 (N_577,N_500,N_496);
nand U578 (N_578,N_493,N_491);
and U579 (N_579,N_492,N_533);
nor U580 (N_580,N_539,N_520);
nor U581 (N_581,N_534,N_493);
nor U582 (N_582,N_522,N_528);
and U583 (N_583,N_502,N_497);
or U584 (N_584,N_508,N_516);
and U585 (N_585,N_524,N_526);
nor U586 (N_586,N_529,N_485);
nand U587 (N_587,N_528,N_507);
or U588 (N_588,N_529,N_514);
or U589 (N_589,N_494,N_524);
xnor U590 (N_590,N_501,N_538);
nor U591 (N_591,N_521,N_513);
nand U592 (N_592,N_504,N_510);
and U593 (N_593,N_522,N_484);
nor U594 (N_594,N_525,N_480);
nand U595 (N_595,N_498,N_502);
or U596 (N_596,N_535,N_515);
and U597 (N_597,N_510,N_536);
or U598 (N_598,N_516,N_522);
nand U599 (N_599,N_485,N_510);
and U600 (N_600,N_540,N_548);
and U601 (N_601,N_580,N_570);
and U602 (N_602,N_573,N_556);
nand U603 (N_603,N_561,N_587);
and U604 (N_604,N_560,N_575);
nor U605 (N_605,N_545,N_583);
and U606 (N_606,N_567,N_554);
nand U607 (N_607,N_557,N_581);
nand U608 (N_608,N_562,N_579);
and U609 (N_609,N_565,N_541);
nand U610 (N_610,N_596,N_571);
nor U611 (N_611,N_547,N_543);
and U612 (N_612,N_552,N_544);
nor U613 (N_613,N_551,N_564);
nor U614 (N_614,N_578,N_574);
or U615 (N_615,N_594,N_550);
nand U616 (N_616,N_586,N_566);
nor U617 (N_617,N_576,N_582);
or U618 (N_618,N_563,N_572);
and U619 (N_619,N_589,N_585);
nand U620 (N_620,N_588,N_553);
and U621 (N_621,N_568,N_590);
nor U622 (N_622,N_584,N_599);
and U623 (N_623,N_591,N_546);
nor U624 (N_624,N_597,N_558);
and U625 (N_625,N_595,N_549);
nand U626 (N_626,N_555,N_542);
nor U627 (N_627,N_577,N_598);
nand U628 (N_628,N_592,N_593);
and U629 (N_629,N_569,N_559);
nor U630 (N_630,N_564,N_558);
nand U631 (N_631,N_581,N_584);
or U632 (N_632,N_547,N_555);
and U633 (N_633,N_582,N_597);
and U634 (N_634,N_549,N_573);
nor U635 (N_635,N_558,N_590);
nand U636 (N_636,N_564,N_569);
or U637 (N_637,N_577,N_587);
and U638 (N_638,N_567,N_568);
and U639 (N_639,N_553,N_590);
and U640 (N_640,N_555,N_551);
or U641 (N_641,N_560,N_558);
or U642 (N_642,N_570,N_583);
nor U643 (N_643,N_595,N_585);
nor U644 (N_644,N_576,N_547);
nor U645 (N_645,N_572,N_574);
xor U646 (N_646,N_588,N_584);
nor U647 (N_647,N_562,N_594);
nand U648 (N_648,N_563,N_580);
nor U649 (N_649,N_551,N_544);
nor U650 (N_650,N_559,N_547);
nor U651 (N_651,N_587,N_596);
nor U652 (N_652,N_547,N_578);
or U653 (N_653,N_586,N_559);
nor U654 (N_654,N_541,N_594);
or U655 (N_655,N_560,N_562);
nand U656 (N_656,N_566,N_588);
nand U657 (N_657,N_545,N_548);
and U658 (N_658,N_593,N_575);
nand U659 (N_659,N_593,N_574);
and U660 (N_660,N_619,N_649);
nand U661 (N_661,N_655,N_650);
or U662 (N_662,N_625,N_634);
xor U663 (N_663,N_640,N_617);
or U664 (N_664,N_658,N_605);
or U665 (N_665,N_656,N_626);
nand U666 (N_666,N_633,N_635);
nand U667 (N_667,N_609,N_638);
or U668 (N_668,N_653,N_642);
nand U669 (N_669,N_603,N_639);
or U670 (N_670,N_630,N_641);
and U671 (N_671,N_621,N_607);
and U672 (N_672,N_602,N_613);
and U673 (N_673,N_636,N_632);
or U674 (N_674,N_646,N_651);
nand U675 (N_675,N_612,N_611);
and U676 (N_676,N_616,N_627);
or U677 (N_677,N_652,N_610);
and U678 (N_678,N_657,N_644);
nor U679 (N_679,N_623,N_618);
and U680 (N_680,N_622,N_637);
nand U681 (N_681,N_648,N_643);
or U682 (N_682,N_614,N_628);
or U683 (N_683,N_654,N_647);
nor U684 (N_684,N_624,N_608);
or U685 (N_685,N_659,N_629);
or U686 (N_686,N_606,N_600);
nor U687 (N_687,N_645,N_601);
or U688 (N_688,N_631,N_615);
or U689 (N_689,N_620,N_604);
nand U690 (N_690,N_610,N_602);
nor U691 (N_691,N_610,N_648);
and U692 (N_692,N_638,N_608);
nand U693 (N_693,N_631,N_642);
nor U694 (N_694,N_626,N_627);
nor U695 (N_695,N_617,N_603);
or U696 (N_696,N_632,N_618);
nor U697 (N_697,N_632,N_643);
nand U698 (N_698,N_659,N_643);
nand U699 (N_699,N_647,N_658);
or U700 (N_700,N_603,N_629);
nand U701 (N_701,N_631,N_613);
and U702 (N_702,N_607,N_645);
and U703 (N_703,N_644,N_618);
nand U704 (N_704,N_656,N_657);
and U705 (N_705,N_655,N_647);
and U706 (N_706,N_632,N_635);
or U707 (N_707,N_602,N_607);
nand U708 (N_708,N_655,N_636);
nand U709 (N_709,N_653,N_628);
and U710 (N_710,N_645,N_630);
nor U711 (N_711,N_617,N_638);
and U712 (N_712,N_636,N_601);
and U713 (N_713,N_600,N_638);
xor U714 (N_714,N_619,N_615);
nor U715 (N_715,N_648,N_608);
or U716 (N_716,N_646,N_637);
and U717 (N_717,N_619,N_650);
and U718 (N_718,N_644,N_645);
nand U719 (N_719,N_642,N_649);
or U720 (N_720,N_690,N_695);
nand U721 (N_721,N_696,N_706);
or U722 (N_722,N_673,N_663);
nand U723 (N_723,N_700,N_699);
or U724 (N_724,N_693,N_709);
nand U725 (N_725,N_698,N_717);
nand U726 (N_726,N_697,N_661);
nand U727 (N_727,N_713,N_716);
or U728 (N_728,N_715,N_684);
nor U729 (N_729,N_666,N_712);
or U730 (N_730,N_679,N_701);
nand U731 (N_731,N_670,N_674);
nand U732 (N_732,N_669,N_678);
or U733 (N_733,N_711,N_664);
nand U734 (N_734,N_708,N_704);
nor U735 (N_735,N_710,N_677);
nand U736 (N_736,N_687,N_692);
nor U737 (N_737,N_707,N_718);
nand U738 (N_738,N_703,N_672);
nand U739 (N_739,N_702,N_686);
and U740 (N_740,N_675,N_671);
nand U741 (N_741,N_719,N_665);
or U742 (N_742,N_660,N_681);
and U743 (N_743,N_705,N_668);
or U744 (N_744,N_662,N_694);
or U745 (N_745,N_683,N_714);
or U746 (N_746,N_667,N_680);
or U747 (N_747,N_689,N_688);
or U748 (N_748,N_682,N_685);
and U749 (N_749,N_691,N_676);
nor U750 (N_750,N_707,N_693);
and U751 (N_751,N_710,N_680);
nor U752 (N_752,N_688,N_663);
nand U753 (N_753,N_696,N_668);
nor U754 (N_754,N_677,N_679);
or U755 (N_755,N_676,N_684);
nand U756 (N_756,N_696,N_675);
and U757 (N_757,N_706,N_674);
or U758 (N_758,N_708,N_669);
and U759 (N_759,N_714,N_665);
and U760 (N_760,N_718,N_708);
and U761 (N_761,N_717,N_689);
nor U762 (N_762,N_699,N_706);
nand U763 (N_763,N_710,N_717);
nor U764 (N_764,N_698,N_688);
xor U765 (N_765,N_670,N_717);
nor U766 (N_766,N_708,N_661);
and U767 (N_767,N_717,N_707);
nand U768 (N_768,N_690,N_718);
nor U769 (N_769,N_694,N_664);
or U770 (N_770,N_685,N_675);
and U771 (N_771,N_682,N_694);
nor U772 (N_772,N_700,N_678);
or U773 (N_773,N_692,N_712);
nor U774 (N_774,N_673,N_670);
nand U775 (N_775,N_667,N_703);
or U776 (N_776,N_672,N_716);
and U777 (N_777,N_666,N_663);
and U778 (N_778,N_689,N_706);
and U779 (N_779,N_662,N_709);
and U780 (N_780,N_751,N_778);
xnor U781 (N_781,N_721,N_761);
or U782 (N_782,N_739,N_735);
nor U783 (N_783,N_757,N_747);
nor U784 (N_784,N_736,N_720);
nor U785 (N_785,N_776,N_762);
or U786 (N_786,N_766,N_734);
nand U787 (N_787,N_738,N_777);
nand U788 (N_788,N_726,N_752);
or U789 (N_789,N_754,N_774);
nor U790 (N_790,N_768,N_758);
nor U791 (N_791,N_750,N_760);
nor U792 (N_792,N_745,N_742);
nor U793 (N_793,N_779,N_755);
nor U794 (N_794,N_733,N_731);
and U795 (N_795,N_764,N_723);
nand U796 (N_796,N_753,N_737);
nor U797 (N_797,N_743,N_770);
and U798 (N_798,N_740,N_746);
or U799 (N_799,N_765,N_759);
nor U800 (N_800,N_725,N_748);
nor U801 (N_801,N_730,N_724);
and U802 (N_802,N_763,N_749);
and U803 (N_803,N_729,N_773);
or U804 (N_804,N_771,N_767);
xor U805 (N_805,N_775,N_756);
or U806 (N_806,N_744,N_769);
nand U807 (N_807,N_732,N_741);
nor U808 (N_808,N_728,N_772);
nand U809 (N_809,N_722,N_727);
or U810 (N_810,N_754,N_741);
nand U811 (N_811,N_730,N_740);
or U812 (N_812,N_732,N_759);
nor U813 (N_813,N_730,N_774);
nor U814 (N_814,N_778,N_741);
nand U815 (N_815,N_765,N_758);
nand U816 (N_816,N_775,N_746);
nor U817 (N_817,N_765,N_757);
nor U818 (N_818,N_737,N_773);
nand U819 (N_819,N_723,N_758);
nor U820 (N_820,N_721,N_770);
nand U821 (N_821,N_748,N_732);
nand U822 (N_822,N_773,N_735);
nor U823 (N_823,N_741,N_763);
nand U824 (N_824,N_767,N_752);
nand U825 (N_825,N_756,N_730);
nand U826 (N_826,N_749,N_753);
nor U827 (N_827,N_725,N_760);
nand U828 (N_828,N_730,N_771);
nor U829 (N_829,N_760,N_766);
or U830 (N_830,N_758,N_727);
nand U831 (N_831,N_748,N_775);
and U832 (N_832,N_731,N_754);
or U833 (N_833,N_735,N_731);
nand U834 (N_834,N_770,N_740);
nand U835 (N_835,N_742,N_759);
or U836 (N_836,N_774,N_732);
nor U837 (N_837,N_740,N_760);
nor U838 (N_838,N_728,N_742);
nor U839 (N_839,N_726,N_723);
nand U840 (N_840,N_835,N_836);
nor U841 (N_841,N_798,N_813);
and U842 (N_842,N_832,N_839);
or U843 (N_843,N_824,N_802);
nand U844 (N_844,N_796,N_793);
and U845 (N_845,N_826,N_794);
nor U846 (N_846,N_809,N_786);
or U847 (N_847,N_792,N_788);
nor U848 (N_848,N_816,N_817);
and U849 (N_849,N_827,N_781);
nor U850 (N_850,N_815,N_818);
or U851 (N_851,N_833,N_780);
or U852 (N_852,N_823,N_834);
nand U853 (N_853,N_821,N_811);
nor U854 (N_854,N_805,N_782);
or U855 (N_855,N_803,N_806);
or U856 (N_856,N_804,N_790);
or U857 (N_857,N_787,N_819);
and U858 (N_858,N_820,N_822);
and U859 (N_859,N_801,N_825);
nor U860 (N_860,N_785,N_791);
or U861 (N_861,N_810,N_812);
xor U862 (N_862,N_807,N_838);
or U863 (N_863,N_814,N_784);
or U864 (N_864,N_783,N_831);
and U865 (N_865,N_800,N_795);
or U866 (N_866,N_837,N_799);
nand U867 (N_867,N_828,N_808);
or U868 (N_868,N_797,N_789);
and U869 (N_869,N_829,N_830);
nor U870 (N_870,N_831,N_800);
or U871 (N_871,N_813,N_815);
nand U872 (N_872,N_803,N_801);
or U873 (N_873,N_831,N_808);
and U874 (N_874,N_812,N_816);
nor U875 (N_875,N_838,N_815);
or U876 (N_876,N_792,N_791);
nand U877 (N_877,N_804,N_795);
and U878 (N_878,N_828,N_826);
and U879 (N_879,N_821,N_805);
or U880 (N_880,N_822,N_792);
nor U881 (N_881,N_786,N_835);
nand U882 (N_882,N_800,N_811);
and U883 (N_883,N_807,N_827);
nor U884 (N_884,N_798,N_804);
nor U885 (N_885,N_811,N_803);
nor U886 (N_886,N_800,N_819);
or U887 (N_887,N_790,N_811);
nor U888 (N_888,N_838,N_793);
and U889 (N_889,N_806,N_789);
nand U890 (N_890,N_806,N_814);
nor U891 (N_891,N_780,N_827);
and U892 (N_892,N_825,N_824);
nor U893 (N_893,N_788,N_786);
and U894 (N_894,N_820,N_795);
or U895 (N_895,N_829,N_832);
nand U896 (N_896,N_801,N_822);
nor U897 (N_897,N_793,N_799);
nor U898 (N_898,N_801,N_815);
nor U899 (N_899,N_792,N_831);
nand U900 (N_900,N_891,N_850);
and U901 (N_901,N_862,N_884);
and U902 (N_902,N_883,N_849);
or U903 (N_903,N_897,N_865);
and U904 (N_904,N_845,N_878);
xor U905 (N_905,N_870,N_843);
and U906 (N_906,N_874,N_889);
or U907 (N_907,N_875,N_885);
nor U908 (N_908,N_877,N_867);
and U909 (N_909,N_859,N_840);
or U910 (N_910,N_860,N_855);
nand U911 (N_911,N_847,N_871);
nor U912 (N_912,N_842,N_882);
nor U913 (N_913,N_853,N_863);
nor U914 (N_914,N_846,N_899);
or U915 (N_915,N_866,N_881);
nor U916 (N_916,N_898,N_876);
or U917 (N_917,N_887,N_856);
nor U918 (N_918,N_880,N_852);
and U919 (N_919,N_864,N_857);
nor U920 (N_920,N_869,N_896);
and U921 (N_921,N_888,N_854);
nand U922 (N_922,N_844,N_848);
nor U923 (N_923,N_868,N_894);
nor U924 (N_924,N_895,N_890);
nor U925 (N_925,N_851,N_879);
nor U926 (N_926,N_886,N_892);
nand U927 (N_927,N_858,N_872);
or U928 (N_928,N_873,N_861);
nor U929 (N_929,N_893,N_841);
and U930 (N_930,N_844,N_860);
nor U931 (N_931,N_894,N_871);
nand U932 (N_932,N_848,N_894);
nand U933 (N_933,N_882,N_861);
and U934 (N_934,N_846,N_879);
and U935 (N_935,N_865,N_873);
nand U936 (N_936,N_886,N_848);
and U937 (N_937,N_855,N_866);
or U938 (N_938,N_879,N_862);
nor U939 (N_939,N_884,N_866);
nor U940 (N_940,N_899,N_863);
or U941 (N_941,N_852,N_872);
nor U942 (N_942,N_877,N_891);
nand U943 (N_943,N_894,N_880);
nand U944 (N_944,N_895,N_869);
or U945 (N_945,N_854,N_840);
or U946 (N_946,N_895,N_857);
nor U947 (N_947,N_845,N_877);
nor U948 (N_948,N_868,N_892);
and U949 (N_949,N_864,N_845);
and U950 (N_950,N_854,N_866);
nand U951 (N_951,N_840,N_846);
and U952 (N_952,N_878,N_884);
nand U953 (N_953,N_898,N_866);
nor U954 (N_954,N_850,N_896);
or U955 (N_955,N_878,N_859);
and U956 (N_956,N_890,N_882);
and U957 (N_957,N_881,N_899);
nand U958 (N_958,N_863,N_873);
and U959 (N_959,N_876,N_854);
nor U960 (N_960,N_925,N_919);
nand U961 (N_961,N_920,N_903);
or U962 (N_962,N_900,N_946);
nand U963 (N_963,N_958,N_908);
nor U964 (N_964,N_955,N_940);
nand U965 (N_965,N_951,N_915);
nand U966 (N_966,N_934,N_916);
nand U967 (N_967,N_912,N_932);
nor U968 (N_968,N_924,N_913);
nor U969 (N_969,N_957,N_905);
and U970 (N_970,N_933,N_927);
nand U971 (N_971,N_937,N_926);
or U972 (N_972,N_910,N_909);
or U973 (N_973,N_935,N_947);
nand U974 (N_974,N_930,N_952);
or U975 (N_975,N_901,N_917);
or U976 (N_976,N_954,N_942);
nor U977 (N_977,N_911,N_953);
nand U978 (N_978,N_928,N_922);
and U979 (N_979,N_943,N_938);
nand U980 (N_980,N_904,N_941);
nor U981 (N_981,N_918,N_929);
nor U982 (N_982,N_948,N_923);
xnor U983 (N_983,N_959,N_944);
nor U984 (N_984,N_949,N_906);
and U985 (N_985,N_956,N_902);
nand U986 (N_986,N_945,N_936);
or U987 (N_987,N_939,N_907);
or U988 (N_988,N_921,N_931);
nor U989 (N_989,N_950,N_914);
nand U990 (N_990,N_937,N_955);
or U991 (N_991,N_907,N_936);
nor U992 (N_992,N_954,N_957);
nand U993 (N_993,N_909,N_916);
or U994 (N_994,N_946,N_937);
nand U995 (N_995,N_913,N_901);
or U996 (N_996,N_930,N_916);
nand U997 (N_997,N_959,N_933);
and U998 (N_998,N_914,N_939);
nand U999 (N_999,N_951,N_938);
nand U1000 (N_1000,N_937,N_952);
or U1001 (N_1001,N_941,N_935);
nand U1002 (N_1002,N_953,N_937);
nand U1003 (N_1003,N_900,N_914);
nor U1004 (N_1004,N_924,N_904);
nand U1005 (N_1005,N_920,N_934);
nand U1006 (N_1006,N_946,N_902);
and U1007 (N_1007,N_923,N_927);
and U1008 (N_1008,N_953,N_957);
and U1009 (N_1009,N_946,N_915);
nor U1010 (N_1010,N_941,N_947);
nor U1011 (N_1011,N_904,N_923);
and U1012 (N_1012,N_922,N_930);
nor U1013 (N_1013,N_929,N_944);
or U1014 (N_1014,N_914,N_924);
or U1015 (N_1015,N_953,N_924);
nor U1016 (N_1016,N_945,N_907);
nor U1017 (N_1017,N_936,N_951);
nor U1018 (N_1018,N_929,N_921);
and U1019 (N_1019,N_939,N_944);
nand U1020 (N_1020,N_1001,N_1010);
or U1021 (N_1021,N_963,N_970);
and U1022 (N_1022,N_984,N_1003);
and U1023 (N_1023,N_973,N_1013);
nor U1024 (N_1024,N_1002,N_980);
or U1025 (N_1025,N_977,N_1011);
and U1026 (N_1026,N_962,N_992);
nand U1027 (N_1027,N_1000,N_1017);
or U1028 (N_1028,N_1005,N_987);
nand U1029 (N_1029,N_985,N_979);
nand U1030 (N_1030,N_1006,N_967);
or U1031 (N_1031,N_960,N_981);
nand U1032 (N_1032,N_1008,N_976);
nand U1033 (N_1033,N_975,N_988);
nor U1034 (N_1034,N_966,N_1016);
and U1035 (N_1035,N_961,N_999);
xnor U1036 (N_1036,N_971,N_997);
nand U1037 (N_1037,N_1009,N_986);
nor U1038 (N_1038,N_1014,N_978);
and U1039 (N_1039,N_1018,N_1012);
and U1040 (N_1040,N_993,N_995);
and U1041 (N_1041,N_1015,N_964);
and U1042 (N_1042,N_989,N_1019);
and U1043 (N_1043,N_991,N_1007);
nand U1044 (N_1044,N_972,N_974);
or U1045 (N_1045,N_998,N_990);
or U1046 (N_1046,N_983,N_965);
nor U1047 (N_1047,N_969,N_968);
nor U1048 (N_1048,N_994,N_1004);
and U1049 (N_1049,N_996,N_982);
nor U1050 (N_1050,N_960,N_1011);
and U1051 (N_1051,N_965,N_997);
or U1052 (N_1052,N_986,N_967);
nor U1053 (N_1053,N_975,N_1000);
or U1054 (N_1054,N_982,N_975);
nand U1055 (N_1055,N_1005,N_998);
and U1056 (N_1056,N_996,N_963);
nor U1057 (N_1057,N_973,N_1009);
nand U1058 (N_1058,N_991,N_993);
and U1059 (N_1059,N_1000,N_967);
and U1060 (N_1060,N_1016,N_967);
or U1061 (N_1061,N_1018,N_981);
nand U1062 (N_1062,N_965,N_976);
and U1063 (N_1063,N_971,N_1002);
xnor U1064 (N_1064,N_981,N_1011);
nor U1065 (N_1065,N_990,N_997);
nand U1066 (N_1066,N_981,N_988);
and U1067 (N_1067,N_967,N_990);
nand U1068 (N_1068,N_1017,N_993);
or U1069 (N_1069,N_1002,N_976);
nand U1070 (N_1070,N_964,N_1009);
nand U1071 (N_1071,N_987,N_1014);
xnor U1072 (N_1072,N_1004,N_969);
and U1073 (N_1073,N_974,N_997);
or U1074 (N_1074,N_985,N_989);
and U1075 (N_1075,N_967,N_996);
or U1076 (N_1076,N_1018,N_1019);
nor U1077 (N_1077,N_985,N_982);
and U1078 (N_1078,N_967,N_964);
or U1079 (N_1079,N_981,N_974);
and U1080 (N_1080,N_1023,N_1071);
and U1081 (N_1081,N_1050,N_1020);
nand U1082 (N_1082,N_1032,N_1022);
nor U1083 (N_1083,N_1024,N_1078);
and U1084 (N_1084,N_1030,N_1051);
or U1085 (N_1085,N_1044,N_1073);
and U1086 (N_1086,N_1068,N_1043);
nor U1087 (N_1087,N_1042,N_1027);
nor U1088 (N_1088,N_1045,N_1054);
or U1089 (N_1089,N_1061,N_1036);
or U1090 (N_1090,N_1029,N_1075);
and U1091 (N_1091,N_1065,N_1026);
or U1092 (N_1092,N_1074,N_1066);
nand U1093 (N_1093,N_1072,N_1039);
or U1094 (N_1094,N_1064,N_1057);
and U1095 (N_1095,N_1079,N_1041);
or U1096 (N_1096,N_1060,N_1031);
nand U1097 (N_1097,N_1025,N_1058);
nor U1098 (N_1098,N_1070,N_1034);
or U1099 (N_1099,N_1067,N_1076);
nor U1100 (N_1100,N_1077,N_1021);
and U1101 (N_1101,N_1048,N_1035);
nor U1102 (N_1102,N_1033,N_1028);
nor U1103 (N_1103,N_1037,N_1053);
or U1104 (N_1104,N_1055,N_1038);
or U1105 (N_1105,N_1047,N_1046);
xnor U1106 (N_1106,N_1069,N_1040);
or U1107 (N_1107,N_1062,N_1052);
or U1108 (N_1108,N_1059,N_1049);
and U1109 (N_1109,N_1063,N_1056);
nand U1110 (N_1110,N_1029,N_1058);
nand U1111 (N_1111,N_1074,N_1069);
nor U1112 (N_1112,N_1020,N_1069);
and U1113 (N_1113,N_1067,N_1069);
nor U1114 (N_1114,N_1068,N_1064);
nor U1115 (N_1115,N_1066,N_1043);
nand U1116 (N_1116,N_1025,N_1046);
and U1117 (N_1117,N_1043,N_1038);
and U1118 (N_1118,N_1057,N_1067);
and U1119 (N_1119,N_1069,N_1055);
or U1120 (N_1120,N_1046,N_1027);
nand U1121 (N_1121,N_1058,N_1067);
and U1122 (N_1122,N_1048,N_1076);
nor U1123 (N_1123,N_1078,N_1055);
xnor U1124 (N_1124,N_1057,N_1029);
nand U1125 (N_1125,N_1049,N_1048);
nor U1126 (N_1126,N_1070,N_1078);
or U1127 (N_1127,N_1033,N_1041);
nor U1128 (N_1128,N_1056,N_1067);
or U1129 (N_1129,N_1048,N_1039);
or U1130 (N_1130,N_1041,N_1023);
nor U1131 (N_1131,N_1041,N_1076);
or U1132 (N_1132,N_1077,N_1069);
or U1133 (N_1133,N_1066,N_1031);
and U1134 (N_1134,N_1029,N_1068);
nand U1135 (N_1135,N_1045,N_1068);
nand U1136 (N_1136,N_1044,N_1046);
nand U1137 (N_1137,N_1046,N_1036);
or U1138 (N_1138,N_1053,N_1041);
nand U1139 (N_1139,N_1068,N_1032);
or U1140 (N_1140,N_1108,N_1139);
and U1141 (N_1141,N_1124,N_1092);
and U1142 (N_1142,N_1112,N_1086);
xnor U1143 (N_1143,N_1091,N_1099);
nand U1144 (N_1144,N_1134,N_1085);
nor U1145 (N_1145,N_1120,N_1130);
nand U1146 (N_1146,N_1105,N_1117);
or U1147 (N_1147,N_1090,N_1089);
and U1148 (N_1148,N_1137,N_1135);
nand U1149 (N_1149,N_1100,N_1128);
and U1150 (N_1150,N_1122,N_1136);
or U1151 (N_1151,N_1132,N_1102);
and U1152 (N_1152,N_1129,N_1126);
and U1153 (N_1153,N_1084,N_1088);
or U1154 (N_1154,N_1107,N_1081);
nor U1155 (N_1155,N_1098,N_1138);
and U1156 (N_1156,N_1111,N_1121);
nand U1157 (N_1157,N_1116,N_1097);
or U1158 (N_1158,N_1104,N_1123);
and U1159 (N_1159,N_1106,N_1113);
and U1160 (N_1160,N_1118,N_1095);
nor U1161 (N_1161,N_1103,N_1127);
or U1162 (N_1162,N_1119,N_1094);
or U1163 (N_1163,N_1083,N_1080);
nand U1164 (N_1164,N_1115,N_1125);
nor U1165 (N_1165,N_1082,N_1114);
nand U1166 (N_1166,N_1096,N_1133);
nor U1167 (N_1167,N_1131,N_1093);
or U1168 (N_1168,N_1087,N_1110);
nand U1169 (N_1169,N_1109,N_1101);
and U1170 (N_1170,N_1090,N_1118);
and U1171 (N_1171,N_1080,N_1124);
and U1172 (N_1172,N_1128,N_1105);
and U1173 (N_1173,N_1124,N_1089);
or U1174 (N_1174,N_1134,N_1092);
and U1175 (N_1175,N_1080,N_1103);
nor U1176 (N_1176,N_1129,N_1084);
nor U1177 (N_1177,N_1103,N_1119);
nor U1178 (N_1178,N_1108,N_1125);
and U1179 (N_1179,N_1135,N_1127);
nand U1180 (N_1180,N_1131,N_1089);
nand U1181 (N_1181,N_1113,N_1132);
xor U1182 (N_1182,N_1091,N_1105);
or U1183 (N_1183,N_1123,N_1101);
nor U1184 (N_1184,N_1081,N_1116);
and U1185 (N_1185,N_1132,N_1105);
or U1186 (N_1186,N_1099,N_1097);
nor U1187 (N_1187,N_1082,N_1104);
nand U1188 (N_1188,N_1134,N_1086);
or U1189 (N_1189,N_1098,N_1127);
or U1190 (N_1190,N_1126,N_1095);
and U1191 (N_1191,N_1104,N_1099);
nor U1192 (N_1192,N_1094,N_1116);
or U1193 (N_1193,N_1086,N_1128);
nor U1194 (N_1194,N_1136,N_1135);
or U1195 (N_1195,N_1116,N_1096);
nor U1196 (N_1196,N_1099,N_1100);
and U1197 (N_1197,N_1083,N_1094);
or U1198 (N_1198,N_1104,N_1095);
or U1199 (N_1199,N_1125,N_1084);
xor U1200 (N_1200,N_1191,N_1167);
and U1201 (N_1201,N_1199,N_1169);
and U1202 (N_1202,N_1163,N_1171);
xnor U1203 (N_1203,N_1154,N_1175);
nand U1204 (N_1204,N_1141,N_1162);
nor U1205 (N_1205,N_1156,N_1165);
nor U1206 (N_1206,N_1146,N_1160);
and U1207 (N_1207,N_1153,N_1144);
and U1208 (N_1208,N_1149,N_1173);
and U1209 (N_1209,N_1177,N_1189);
or U1210 (N_1210,N_1186,N_1196);
nand U1211 (N_1211,N_1181,N_1185);
and U1212 (N_1212,N_1178,N_1182);
nand U1213 (N_1213,N_1170,N_1187);
and U1214 (N_1214,N_1183,N_1193);
nand U1215 (N_1215,N_1176,N_1155);
and U1216 (N_1216,N_1143,N_1180);
and U1217 (N_1217,N_1179,N_1190);
or U1218 (N_1218,N_1174,N_1140);
and U1219 (N_1219,N_1157,N_1150);
and U1220 (N_1220,N_1172,N_1198);
or U1221 (N_1221,N_1166,N_1195);
xnor U1222 (N_1222,N_1168,N_1192);
or U1223 (N_1223,N_1151,N_1159);
or U1224 (N_1224,N_1164,N_1197);
nand U1225 (N_1225,N_1158,N_1142);
and U1226 (N_1226,N_1188,N_1145);
or U1227 (N_1227,N_1161,N_1148);
and U1228 (N_1228,N_1147,N_1152);
and U1229 (N_1229,N_1184,N_1194);
and U1230 (N_1230,N_1143,N_1146);
nor U1231 (N_1231,N_1187,N_1148);
or U1232 (N_1232,N_1179,N_1191);
nand U1233 (N_1233,N_1140,N_1160);
nand U1234 (N_1234,N_1145,N_1153);
and U1235 (N_1235,N_1192,N_1180);
and U1236 (N_1236,N_1150,N_1191);
and U1237 (N_1237,N_1175,N_1165);
and U1238 (N_1238,N_1188,N_1180);
or U1239 (N_1239,N_1188,N_1146);
or U1240 (N_1240,N_1174,N_1187);
nor U1241 (N_1241,N_1163,N_1164);
nor U1242 (N_1242,N_1141,N_1164);
or U1243 (N_1243,N_1196,N_1162);
nor U1244 (N_1244,N_1195,N_1141);
xnor U1245 (N_1245,N_1144,N_1146);
or U1246 (N_1246,N_1153,N_1150);
nor U1247 (N_1247,N_1149,N_1153);
xor U1248 (N_1248,N_1154,N_1169);
nor U1249 (N_1249,N_1182,N_1156);
nor U1250 (N_1250,N_1173,N_1197);
xor U1251 (N_1251,N_1142,N_1174);
xnor U1252 (N_1252,N_1178,N_1142);
and U1253 (N_1253,N_1193,N_1195);
or U1254 (N_1254,N_1144,N_1196);
nand U1255 (N_1255,N_1183,N_1151);
or U1256 (N_1256,N_1166,N_1161);
or U1257 (N_1257,N_1189,N_1192);
nand U1258 (N_1258,N_1181,N_1194);
or U1259 (N_1259,N_1144,N_1186);
or U1260 (N_1260,N_1222,N_1258);
nand U1261 (N_1261,N_1218,N_1248);
nor U1262 (N_1262,N_1223,N_1209);
or U1263 (N_1263,N_1244,N_1259);
nand U1264 (N_1264,N_1247,N_1217);
or U1265 (N_1265,N_1215,N_1254);
nor U1266 (N_1266,N_1208,N_1242);
or U1267 (N_1267,N_1225,N_1255);
nor U1268 (N_1268,N_1220,N_1251);
nor U1269 (N_1269,N_1237,N_1224);
and U1270 (N_1270,N_1214,N_1232);
or U1271 (N_1271,N_1245,N_1204);
nand U1272 (N_1272,N_1202,N_1210);
nand U1273 (N_1273,N_1200,N_1229);
or U1274 (N_1274,N_1216,N_1256);
nand U1275 (N_1275,N_1253,N_1213);
nand U1276 (N_1276,N_1240,N_1234);
and U1277 (N_1277,N_1230,N_1231);
nor U1278 (N_1278,N_1241,N_1207);
nand U1279 (N_1279,N_1205,N_1250);
or U1280 (N_1280,N_1221,N_1239);
or U1281 (N_1281,N_1206,N_1252);
nor U1282 (N_1282,N_1235,N_1236);
and U1283 (N_1283,N_1226,N_1243);
nand U1284 (N_1284,N_1212,N_1227);
or U1285 (N_1285,N_1219,N_1246);
nand U1286 (N_1286,N_1257,N_1211);
nand U1287 (N_1287,N_1201,N_1249);
nor U1288 (N_1288,N_1233,N_1238);
or U1289 (N_1289,N_1203,N_1228);
and U1290 (N_1290,N_1259,N_1240);
nor U1291 (N_1291,N_1250,N_1244);
nor U1292 (N_1292,N_1259,N_1241);
nand U1293 (N_1293,N_1209,N_1217);
nor U1294 (N_1294,N_1204,N_1247);
or U1295 (N_1295,N_1231,N_1212);
and U1296 (N_1296,N_1255,N_1251);
nand U1297 (N_1297,N_1215,N_1216);
nand U1298 (N_1298,N_1245,N_1256);
nand U1299 (N_1299,N_1220,N_1216);
and U1300 (N_1300,N_1219,N_1200);
nor U1301 (N_1301,N_1241,N_1201);
nor U1302 (N_1302,N_1250,N_1237);
or U1303 (N_1303,N_1211,N_1205);
and U1304 (N_1304,N_1237,N_1218);
or U1305 (N_1305,N_1231,N_1233);
or U1306 (N_1306,N_1243,N_1249);
and U1307 (N_1307,N_1251,N_1206);
xor U1308 (N_1308,N_1249,N_1200);
or U1309 (N_1309,N_1243,N_1245);
nand U1310 (N_1310,N_1235,N_1217);
nand U1311 (N_1311,N_1231,N_1244);
and U1312 (N_1312,N_1204,N_1217);
or U1313 (N_1313,N_1246,N_1250);
and U1314 (N_1314,N_1201,N_1226);
nor U1315 (N_1315,N_1254,N_1226);
nor U1316 (N_1316,N_1242,N_1223);
and U1317 (N_1317,N_1209,N_1215);
and U1318 (N_1318,N_1258,N_1208);
nor U1319 (N_1319,N_1256,N_1249);
nor U1320 (N_1320,N_1266,N_1260);
and U1321 (N_1321,N_1289,N_1284);
nor U1322 (N_1322,N_1279,N_1280);
xor U1323 (N_1323,N_1261,N_1299);
or U1324 (N_1324,N_1296,N_1297);
nor U1325 (N_1325,N_1292,N_1298);
nand U1326 (N_1326,N_1272,N_1311);
xnor U1327 (N_1327,N_1306,N_1294);
or U1328 (N_1328,N_1293,N_1317);
and U1329 (N_1329,N_1278,N_1291);
nand U1330 (N_1330,N_1263,N_1267);
or U1331 (N_1331,N_1281,N_1307);
and U1332 (N_1332,N_1304,N_1276);
nand U1333 (N_1333,N_1312,N_1277);
nand U1334 (N_1334,N_1287,N_1316);
and U1335 (N_1335,N_1295,N_1271);
nand U1336 (N_1336,N_1282,N_1303);
nand U1337 (N_1337,N_1310,N_1269);
nor U1338 (N_1338,N_1308,N_1274);
nand U1339 (N_1339,N_1268,N_1285);
nand U1340 (N_1340,N_1302,N_1319);
nor U1341 (N_1341,N_1286,N_1315);
or U1342 (N_1342,N_1288,N_1262);
nand U1343 (N_1343,N_1264,N_1300);
and U1344 (N_1344,N_1273,N_1301);
nor U1345 (N_1345,N_1270,N_1290);
or U1346 (N_1346,N_1265,N_1305);
or U1347 (N_1347,N_1314,N_1318);
nor U1348 (N_1348,N_1309,N_1275);
and U1349 (N_1349,N_1313,N_1283);
nor U1350 (N_1350,N_1306,N_1309);
nand U1351 (N_1351,N_1261,N_1306);
nor U1352 (N_1352,N_1260,N_1261);
nor U1353 (N_1353,N_1305,N_1287);
and U1354 (N_1354,N_1315,N_1272);
or U1355 (N_1355,N_1316,N_1279);
and U1356 (N_1356,N_1288,N_1287);
xnor U1357 (N_1357,N_1277,N_1304);
or U1358 (N_1358,N_1294,N_1304);
and U1359 (N_1359,N_1270,N_1271);
nor U1360 (N_1360,N_1316,N_1305);
or U1361 (N_1361,N_1272,N_1268);
or U1362 (N_1362,N_1314,N_1303);
or U1363 (N_1363,N_1282,N_1300);
nand U1364 (N_1364,N_1289,N_1309);
and U1365 (N_1365,N_1314,N_1308);
and U1366 (N_1366,N_1286,N_1260);
nor U1367 (N_1367,N_1305,N_1269);
nand U1368 (N_1368,N_1301,N_1270);
nor U1369 (N_1369,N_1310,N_1295);
nor U1370 (N_1370,N_1282,N_1268);
and U1371 (N_1371,N_1307,N_1293);
nand U1372 (N_1372,N_1301,N_1282);
nand U1373 (N_1373,N_1282,N_1313);
nand U1374 (N_1374,N_1285,N_1317);
xor U1375 (N_1375,N_1290,N_1309);
or U1376 (N_1376,N_1283,N_1285);
nand U1377 (N_1377,N_1288,N_1302);
xnor U1378 (N_1378,N_1276,N_1293);
nand U1379 (N_1379,N_1288,N_1274);
and U1380 (N_1380,N_1352,N_1331);
nor U1381 (N_1381,N_1371,N_1351);
nand U1382 (N_1382,N_1346,N_1327);
nor U1383 (N_1383,N_1338,N_1337);
nand U1384 (N_1384,N_1377,N_1378);
nor U1385 (N_1385,N_1366,N_1335);
and U1386 (N_1386,N_1348,N_1355);
nor U1387 (N_1387,N_1336,N_1340);
nor U1388 (N_1388,N_1347,N_1325);
nor U1389 (N_1389,N_1342,N_1367);
nand U1390 (N_1390,N_1375,N_1344);
or U1391 (N_1391,N_1343,N_1334);
and U1392 (N_1392,N_1373,N_1322);
nor U1393 (N_1393,N_1324,N_1360);
nand U1394 (N_1394,N_1321,N_1323);
and U1395 (N_1395,N_1341,N_1333);
or U1396 (N_1396,N_1339,N_1329);
or U1397 (N_1397,N_1354,N_1363);
and U1398 (N_1398,N_1357,N_1356);
nor U1399 (N_1399,N_1372,N_1350);
xor U1400 (N_1400,N_1349,N_1368);
nor U1401 (N_1401,N_1376,N_1320);
or U1402 (N_1402,N_1345,N_1332);
or U1403 (N_1403,N_1364,N_1330);
nor U1404 (N_1404,N_1379,N_1361);
nand U1405 (N_1405,N_1369,N_1353);
or U1406 (N_1406,N_1358,N_1365);
or U1407 (N_1407,N_1362,N_1328);
nor U1408 (N_1408,N_1374,N_1359);
xnor U1409 (N_1409,N_1370,N_1326);
and U1410 (N_1410,N_1342,N_1371);
nand U1411 (N_1411,N_1332,N_1336);
and U1412 (N_1412,N_1364,N_1350);
nand U1413 (N_1413,N_1376,N_1352);
nor U1414 (N_1414,N_1366,N_1352);
or U1415 (N_1415,N_1340,N_1372);
nor U1416 (N_1416,N_1356,N_1328);
or U1417 (N_1417,N_1350,N_1353);
nand U1418 (N_1418,N_1373,N_1349);
nand U1419 (N_1419,N_1338,N_1340);
nor U1420 (N_1420,N_1351,N_1345);
and U1421 (N_1421,N_1369,N_1350);
or U1422 (N_1422,N_1365,N_1334);
nor U1423 (N_1423,N_1327,N_1355);
and U1424 (N_1424,N_1343,N_1371);
or U1425 (N_1425,N_1372,N_1325);
nand U1426 (N_1426,N_1343,N_1364);
or U1427 (N_1427,N_1363,N_1379);
or U1428 (N_1428,N_1344,N_1327);
or U1429 (N_1429,N_1372,N_1366);
and U1430 (N_1430,N_1335,N_1345);
xnor U1431 (N_1431,N_1329,N_1361);
nand U1432 (N_1432,N_1368,N_1379);
nand U1433 (N_1433,N_1373,N_1333);
or U1434 (N_1434,N_1350,N_1379);
nand U1435 (N_1435,N_1344,N_1361);
and U1436 (N_1436,N_1321,N_1322);
and U1437 (N_1437,N_1378,N_1329);
nor U1438 (N_1438,N_1359,N_1323);
and U1439 (N_1439,N_1378,N_1356);
nand U1440 (N_1440,N_1406,N_1387);
and U1441 (N_1441,N_1422,N_1380);
or U1442 (N_1442,N_1382,N_1411);
or U1443 (N_1443,N_1419,N_1416);
nand U1444 (N_1444,N_1393,N_1395);
or U1445 (N_1445,N_1381,N_1405);
nor U1446 (N_1446,N_1421,N_1385);
nand U1447 (N_1447,N_1407,N_1410);
nand U1448 (N_1448,N_1383,N_1397);
nand U1449 (N_1449,N_1435,N_1430);
or U1450 (N_1450,N_1408,N_1390);
and U1451 (N_1451,N_1386,N_1420);
nor U1452 (N_1452,N_1432,N_1412);
or U1453 (N_1453,N_1402,N_1431);
nor U1454 (N_1454,N_1404,N_1436);
nor U1455 (N_1455,N_1423,N_1414);
and U1456 (N_1456,N_1391,N_1427);
or U1457 (N_1457,N_1396,N_1400);
or U1458 (N_1458,N_1415,N_1398);
nand U1459 (N_1459,N_1438,N_1417);
nor U1460 (N_1460,N_1434,N_1439);
and U1461 (N_1461,N_1418,N_1413);
or U1462 (N_1462,N_1429,N_1409);
or U1463 (N_1463,N_1401,N_1392);
nor U1464 (N_1464,N_1424,N_1403);
or U1465 (N_1465,N_1426,N_1437);
or U1466 (N_1466,N_1399,N_1388);
or U1467 (N_1467,N_1433,N_1389);
or U1468 (N_1468,N_1384,N_1425);
or U1469 (N_1469,N_1428,N_1394);
nor U1470 (N_1470,N_1435,N_1393);
nand U1471 (N_1471,N_1383,N_1384);
and U1472 (N_1472,N_1396,N_1411);
and U1473 (N_1473,N_1410,N_1429);
and U1474 (N_1474,N_1381,N_1433);
and U1475 (N_1475,N_1406,N_1411);
nand U1476 (N_1476,N_1418,N_1384);
or U1477 (N_1477,N_1415,N_1430);
nor U1478 (N_1478,N_1394,N_1422);
nor U1479 (N_1479,N_1416,N_1402);
nand U1480 (N_1480,N_1394,N_1411);
and U1481 (N_1481,N_1437,N_1388);
nand U1482 (N_1482,N_1438,N_1432);
nand U1483 (N_1483,N_1420,N_1439);
nor U1484 (N_1484,N_1431,N_1436);
or U1485 (N_1485,N_1416,N_1386);
nor U1486 (N_1486,N_1386,N_1408);
nand U1487 (N_1487,N_1429,N_1414);
or U1488 (N_1488,N_1428,N_1423);
nand U1489 (N_1489,N_1399,N_1417);
nand U1490 (N_1490,N_1397,N_1402);
and U1491 (N_1491,N_1388,N_1426);
nand U1492 (N_1492,N_1433,N_1409);
nor U1493 (N_1493,N_1425,N_1421);
and U1494 (N_1494,N_1392,N_1398);
or U1495 (N_1495,N_1418,N_1382);
or U1496 (N_1496,N_1393,N_1418);
and U1497 (N_1497,N_1393,N_1394);
or U1498 (N_1498,N_1397,N_1400);
nand U1499 (N_1499,N_1433,N_1404);
nor U1500 (N_1500,N_1499,N_1474);
or U1501 (N_1501,N_1455,N_1480);
and U1502 (N_1502,N_1440,N_1475);
or U1503 (N_1503,N_1488,N_1461);
and U1504 (N_1504,N_1454,N_1494);
and U1505 (N_1505,N_1466,N_1449);
and U1506 (N_1506,N_1497,N_1492);
nand U1507 (N_1507,N_1446,N_1498);
and U1508 (N_1508,N_1441,N_1448);
or U1509 (N_1509,N_1486,N_1496);
nand U1510 (N_1510,N_1490,N_1487);
and U1511 (N_1511,N_1462,N_1442);
or U1512 (N_1512,N_1468,N_1495);
nor U1513 (N_1513,N_1452,N_1473);
xnor U1514 (N_1514,N_1464,N_1471);
or U1515 (N_1515,N_1493,N_1453);
nor U1516 (N_1516,N_1485,N_1476);
nor U1517 (N_1517,N_1459,N_1483);
nand U1518 (N_1518,N_1465,N_1484);
nor U1519 (N_1519,N_1467,N_1489);
and U1520 (N_1520,N_1478,N_1479);
or U1521 (N_1521,N_1477,N_1451);
or U1522 (N_1522,N_1445,N_1458);
nor U1523 (N_1523,N_1481,N_1447);
and U1524 (N_1524,N_1457,N_1460);
nand U1525 (N_1525,N_1463,N_1443);
and U1526 (N_1526,N_1491,N_1482);
or U1527 (N_1527,N_1469,N_1444);
or U1528 (N_1528,N_1470,N_1450);
nor U1529 (N_1529,N_1456,N_1472);
and U1530 (N_1530,N_1450,N_1494);
xnor U1531 (N_1531,N_1468,N_1466);
or U1532 (N_1532,N_1489,N_1460);
nor U1533 (N_1533,N_1488,N_1446);
or U1534 (N_1534,N_1443,N_1492);
nor U1535 (N_1535,N_1440,N_1484);
and U1536 (N_1536,N_1467,N_1476);
nand U1537 (N_1537,N_1461,N_1491);
or U1538 (N_1538,N_1484,N_1455);
nor U1539 (N_1539,N_1495,N_1451);
or U1540 (N_1540,N_1484,N_1481);
nand U1541 (N_1541,N_1441,N_1460);
and U1542 (N_1542,N_1471,N_1450);
nand U1543 (N_1543,N_1476,N_1480);
and U1544 (N_1544,N_1470,N_1472);
and U1545 (N_1545,N_1442,N_1486);
or U1546 (N_1546,N_1455,N_1446);
and U1547 (N_1547,N_1452,N_1498);
or U1548 (N_1548,N_1445,N_1467);
nor U1549 (N_1549,N_1481,N_1462);
nand U1550 (N_1550,N_1497,N_1454);
nor U1551 (N_1551,N_1464,N_1478);
nand U1552 (N_1552,N_1478,N_1488);
nand U1553 (N_1553,N_1498,N_1477);
or U1554 (N_1554,N_1477,N_1454);
nand U1555 (N_1555,N_1444,N_1453);
nand U1556 (N_1556,N_1465,N_1453);
or U1557 (N_1557,N_1461,N_1448);
and U1558 (N_1558,N_1481,N_1464);
or U1559 (N_1559,N_1465,N_1454);
nor U1560 (N_1560,N_1510,N_1532);
nand U1561 (N_1561,N_1556,N_1508);
nor U1562 (N_1562,N_1559,N_1551);
nor U1563 (N_1563,N_1517,N_1547);
or U1564 (N_1564,N_1537,N_1506);
or U1565 (N_1565,N_1522,N_1534);
and U1566 (N_1566,N_1545,N_1539);
and U1567 (N_1567,N_1535,N_1519);
and U1568 (N_1568,N_1505,N_1554);
nand U1569 (N_1569,N_1531,N_1538);
and U1570 (N_1570,N_1503,N_1530);
nand U1571 (N_1571,N_1536,N_1558);
nand U1572 (N_1572,N_1507,N_1548);
nor U1573 (N_1573,N_1512,N_1516);
nand U1574 (N_1574,N_1550,N_1518);
nor U1575 (N_1575,N_1526,N_1514);
or U1576 (N_1576,N_1524,N_1500);
or U1577 (N_1577,N_1542,N_1557);
nand U1578 (N_1578,N_1523,N_1504);
nor U1579 (N_1579,N_1515,N_1527);
nand U1580 (N_1580,N_1529,N_1502);
nand U1581 (N_1581,N_1544,N_1509);
nor U1582 (N_1582,N_1549,N_1553);
nor U1583 (N_1583,N_1543,N_1552);
nor U1584 (N_1584,N_1555,N_1546);
nor U1585 (N_1585,N_1541,N_1511);
nor U1586 (N_1586,N_1533,N_1540);
or U1587 (N_1587,N_1528,N_1520);
nor U1588 (N_1588,N_1513,N_1521);
or U1589 (N_1589,N_1501,N_1525);
or U1590 (N_1590,N_1510,N_1509);
nor U1591 (N_1591,N_1552,N_1544);
and U1592 (N_1592,N_1508,N_1505);
and U1593 (N_1593,N_1534,N_1530);
nand U1594 (N_1594,N_1530,N_1523);
nand U1595 (N_1595,N_1522,N_1507);
nand U1596 (N_1596,N_1504,N_1500);
or U1597 (N_1597,N_1533,N_1543);
nor U1598 (N_1598,N_1555,N_1543);
nand U1599 (N_1599,N_1533,N_1538);
and U1600 (N_1600,N_1510,N_1528);
and U1601 (N_1601,N_1519,N_1528);
and U1602 (N_1602,N_1530,N_1541);
and U1603 (N_1603,N_1557,N_1553);
and U1604 (N_1604,N_1507,N_1542);
nand U1605 (N_1605,N_1531,N_1529);
and U1606 (N_1606,N_1501,N_1532);
and U1607 (N_1607,N_1545,N_1503);
xnor U1608 (N_1608,N_1525,N_1515);
or U1609 (N_1609,N_1500,N_1518);
or U1610 (N_1610,N_1530,N_1516);
nor U1611 (N_1611,N_1525,N_1557);
nand U1612 (N_1612,N_1547,N_1511);
and U1613 (N_1613,N_1532,N_1500);
and U1614 (N_1614,N_1503,N_1556);
or U1615 (N_1615,N_1510,N_1501);
and U1616 (N_1616,N_1530,N_1510);
or U1617 (N_1617,N_1557,N_1534);
and U1618 (N_1618,N_1518,N_1503);
nor U1619 (N_1619,N_1527,N_1531);
or U1620 (N_1620,N_1601,N_1578);
nor U1621 (N_1621,N_1562,N_1571);
and U1622 (N_1622,N_1617,N_1586);
and U1623 (N_1623,N_1580,N_1611);
and U1624 (N_1624,N_1561,N_1568);
and U1625 (N_1625,N_1598,N_1604);
nor U1626 (N_1626,N_1572,N_1575);
nand U1627 (N_1627,N_1603,N_1590);
and U1628 (N_1628,N_1608,N_1565);
or U1629 (N_1629,N_1612,N_1560);
or U1630 (N_1630,N_1570,N_1574);
xnor U1631 (N_1631,N_1613,N_1589);
xnor U1632 (N_1632,N_1585,N_1600);
nand U1633 (N_1633,N_1576,N_1584);
or U1634 (N_1634,N_1591,N_1619);
or U1635 (N_1635,N_1587,N_1606);
and U1636 (N_1636,N_1599,N_1610);
or U1637 (N_1637,N_1616,N_1569);
nor U1638 (N_1638,N_1583,N_1577);
and U1639 (N_1639,N_1579,N_1607);
or U1640 (N_1640,N_1593,N_1567);
nor U1641 (N_1641,N_1605,N_1615);
and U1642 (N_1642,N_1596,N_1592);
nor U1643 (N_1643,N_1581,N_1602);
or U1644 (N_1644,N_1594,N_1595);
and U1645 (N_1645,N_1566,N_1609);
and U1646 (N_1646,N_1582,N_1597);
xor U1647 (N_1647,N_1618,N_1588);
or U1648 (N_1648,N_1573,N_1563);
nor U1649 (N_1649,N_1614,N_1564);
and U1650 (N_1650,N_1607,N_1572);
and U1651 (N_1651,N_1597,N_1585);
and U1652 (N_1652,N_1571,N_1575);
and U1653 (N_1653,N_1609,N_1565);
or U1654 (N_1654,N_1596,N_1605);
nor U1655 (N_1655,N_1602,N_1572);
or U1656 (N_1656,N_1603,N_1577);
or U1657 (N_1657,N_1615,N_1560);
or U1658 (N_1658,N_1579,N_1562);
nand U1659 (N_1659,N_1581,N_1578);
nor U1660 (N_1660,N_1596,N_1604);
nand U1661 (N_1661,N_1562,N_1606);
nand U1662 (N_1662,N_1589,N_1612);
or U1663 (N_1663,N_1612,N_1582);
and U1664 (N_1664,N_1608,N_1571);
nand U1665 (N_1665,N_1618,N_1575);
and U1666 (N_1666,N_1570,N_1588);
and U1667 (N_1667,N_1569,N_1586);
or U1668 (N_1668,N_1619,N_1570);
nor U1669 (N_1669,N_1604,N_1586);
or U1670 (N_1670,N_1605,N_1587);
nand U1671 (N_1671,N_1572,N_1600);
nand U1672 (N_1672,N_1569,N_1590);
and U1673 (N_1673,N_1585,N_1568);
nor U1674 (N_1674,N_1603,N_1586);
or U1675 (N_1675,N_1573,N_1579);
and U1676 (N_1676,N_1614,N_1571);
and U1677 (N_1677,N_1572,N_1619);
and U1678 (N_1678,N_1577,N_1565);
nand U1679 (N_1679,N_1609,N_1589);
or U1680 (N_1680,N_1645,N_1642);
nand U1681 (N_1681,N_1639,N_1623);
or U1682 (N_1682,N_1630,N_1675);
and U1683 (N_1683,N_1648,N_1668);
nand U1684 (N_1684,N_1672,N_1664);
and U1685 (N_1685,N_1634,N_1671);
or U1686 (N_1686,N_1627,N_1643);
and U1687 (N_1687,N_1673,N_1679);
or U1688 (N_1688,N_1652,N_1655);
nand U1689 (N_1689,N_1621,N_1658);
and U1690 (N_1690,N_1670,N_1676);
or U1691 (N_1691,N_1649,N_1651);
and U1692 (N_1692,N_1662,N_1632);
nor U1693 (N_1693,N_1625,N_1669);
or U1694 (N_1694,N_1644,N_1624);
nor U1695 (N_1695,N_1633,N_1663);
or U1696 (N_1696,N_1657,N_1665);
and U1697 (N_1697,N_1620,N_1637);
and U1698 (N_1698,N_1622,N_1678);
nand U1699 (N_1699,N_1667,N_1629);
or U1700 (N_1700,N_1674,N_1666);
nor U1701 (N_1701,N_1650,N_1659);
nand U1702 (N_1702,N_1640,N_1660);
nand U1703 (N_1703,N_1677,N_1626);
and U1704 (N_1704,N_1641,N_1636);
nand U1705 (N_1705,N_1656,N_1661);
nor U1706 (N_1706,N_1628,N_1635);
nor U1707 (N_1707,N_1638,N_1646);
and U1708 (N_1708,N_1647,N_1631);
nor U1709 (N_1709,N_1654,N_1653);
or U1710 (N_1710,N_1650,N_1663);
or U1711 (N_1711,N_1636,N_1626);
and U1712 (N_1712,N_1661,N_1657);
and U1713 (N_1713,N_1646,N_1664);
or U1714 (N_1714,N_1633,N_1628);
and U1715 (N_1715,N_1667,N_1635);
and U1716 (N_1716,N_1636,N_1668);
and U1717 (N_1717,N_1665,N_1642);
nor U1718 (N_1718,N_1657,N_1635);
nor U1719 (N_1719,N_1669,N_1646);
nor U1720 (N_1720,N_1631,N_1622);
or U1721 (N_1721,N_1636,N_1651);
nand U1722 (N_1722,N_1625,N_1650);
and U1723 (N_1723,N_1629,N_1675);
nor U1724 (N_1724,N_1676,N_1638);
or U1725 (N_1725,N_1670,N_1677);
xnor U1726 (N_1726,N_1647,N_1621);
nand U1727 (N_1727,N_1642,N_1660);
and U1728 (N_1728,N_1646,N_1662);
nor U1729 (N_1729,N_1664,N_1678);
nand U1730 (N_1730,N_1670,N_1644);
or U1731 (N_1731,N_1622,N_1667);
nand U1732 (N_1732,N_1642,N_1650);
nor U1733 (N_1733,N_1679,N_1672);
nand U1734 (N_1734,N_1627,N_1651);
or U1735 (N_1735,N_1636,N_1645);
nand U1736 (N_1736,N_1633,N_1662);
nand U1737 (N_1737,N_1669,N_1668);
or U1738 (N_1738,N_1632,N_1630);
and U1739 (N_1739,N_1642,N_1676);
and U1740 (N_1740,N_1709,N_1713);
and U1741 (N_1741,N_1723,N_1717);
or U1742 (N_1742,N_1694,N_1738);
and U1743 (N_1743,N_1684,N_1707);
or U1744 (N_1744,N_1729,N_1706);
or U1745 (N_1745,N_1682,N_1728);
or U1746 (N_1746,N_1692,N_1698);
nor U1747 (N_1747,N_1724,N_1720);
xor U1748 (N_1748,N_1686,N_1710);
or U1749 (N_1749,N_1730,N_1739);
or U1750 (N_1750,N_1704,N_1726);
nand U1751 (N_1751,N_1732,N_1727);
or U1752 (N_1752,N_1701,N_1685);
nand U1753 (N_1753,N_1696,N_1695);
and U1754 (N_1754,N_1689,N_1683);
nor U1755 (N_1755,N_1736,N_1725);
nor U1756 (N_1756,N_1722,N_1734);
or U1757 (N_1757,N_1737,N_1700);
nor U1758 (N_1758,N_1721,N_1731);
or U1759 (N_1759,N_1714,N_1687);
nand U1760 (N_1760,N_1688,N_1680);
or U1761 (N_1761,N_1697,N_1703);
nand U1762 (N_1762,N_1708,N_1699);
and U1763 (N_1763,N_1719,N_1702);
and U1764 (N_1764,N_1711,N_1690);
and U1765 (N_1765,N_1716,N_1712);
and U1766 (N_1766,N_1693,N_1715);
nor U1767 (N_1767,N_1681,N_1705);
nor U1768 (N_1768,N_1733,N_1718);
and U1769 (N_1769,N_1691,N_1735);
nor U1770 (N_1770,N_1707,N_1724);
nor U1771 (N_1771,N_1736,N_1712);
and U1772 (N_1772,N_1692,N_1730);
nand U1773 (N_1773,N_1736,N_1730);
or U1774 (N_1774,N_1696,N_1706);
nor U1775 (N_1775,N_1692,N_1739);
nor U1776 (N_1776,N_1719,N_1711);
nor U1777 (N_1777,N_1737,N_1682);
and U1778 (N_1778,N_1689,N_1711);
nand U1779 (N_1779,N_1694,N_1692);
and U1780 (N_1780,N_1696,N_1715);
and U1781 (N_1781,N_1733,N_1680);
nor U1782 (N_1782,N_1701,N_1715);
xor U1783 (N_1783,N_1712,N_1725);
or U1784 (N_1784,N_1719,N_1681);
nand U1785 (N_1785,N_1715,N_1713);
or U1786 (N_1786,N_1690,N_1700);
and U1787 (N_1787,N_1709,N_1723);
nor U1788 (N_1788,N_1711,N_1706);
or U1789 (N_1789,N_1691,N_1736);
and U1790 (N_1790,N_1708,N_1709);
or U1791 (N_1791,N_1703,N_1684);
nand U1792 (N_1792,N_1712,N_1738);
nand U1793 (N_1793,N_1694,N_1700);
nand U1794 (N_1794,N_1727,N_1684);
or U1795 (N_1795,N_1699,N_1736);
nand U1796 (N_1796,N_1728,N_1689);
xor U1797 (N_1797,N_1691,N_1695);
and U1798 (N_1798,N_1724,N_1710);
nand U1799 (N_1799,N_1709,N_1680);
and U1800 (N_1800,N_1796,N_1740);
nand U1801 (N_1801,N_1794,N_1757);
and U1802 (N_1802,N_1780,N_1787);
and U1803 (N_1803,N_1789,N_1758);
and U1804 (N_1804,N_1752,N_1768);
nor U1805 (N_1805,N_1763,N_1778);
nor U1806 (N_1806,N_1785,N_1793);
nor U1807 (N_1807,N_1765,N_1741);
nand U1808 (N_1808,N_1779,N_1770);
and U1809 (N_1809,N_1745,N_1754);
and U1810 (N_1810,N_1773,N_1759);
nor U1811 (N_1811,N_1767,N_1764);
nand U1812 (N_1812,N_1775,N_1755);
or U1813 (N_1813,N_1749,N_1795);
nand U1814 (N_1814,N_1751,N_1756);
and U1815 (N_1815,N_1784,N_1762);
and U1816 (N_1816,N_1799,N_1772);
or U1817 (N_1817,N_1774,N_1782);
or U1818 (N_1818,N_1791,N_1777);
nand U1819 (N_1819,N_1769,N_1742);
or U1820 (N_1820,N_1798,N_1776);
or U1821 (N_1821,N_1792,N_1797);
or U1822 (N_1822,N_1766,N_1747);
or U1823 (N_1823,N_1746,N_1786);
nor U1824 (N_1824,N_1788,N_1761);
or U1825 (N_1825,N_1743,N_1753);
nand U1826 (N_1826,N_1748,N_1744);
nand U1827 (N_1827,N_1781,N_1790);
nand U1828 (N_1828,N_1783,N_1760);
and U1829 (N_1829,N_1771,N_1750);
or U1830 (N_1830,N_1795,N_1747);
and U1831 (N_1831,N_1765,N_1761);
and U1832 (N_1832,N_1785,N_1753);
nor U1833 (N_1833,N_1786,N_1772);
and U1834 (N_1834,N_1747,N_1790);
or U1835 (N_1835,N_1740,N_1769);
or U1836 (N_1836,N_1780,N_1792);
and U1837 (N_1837,N_1788,N_1751);
nor U1838 (N_1838,N_1766,N_1762);
and U1839 (N_1839,N_1743,N_1758);
nand U1840 (N_1840,N_1753,N_1764);
nand U1841 (N_1841,N_1778,N_1773);
or U1842 (N_1842,N_1756,N_1777);
nor U1843 (N_1843,N_1750,N_1741);
nor U1844 (N_1844,N_1753,N_1797);
nor U1845 (N_1845,N_1743,N_1761);
nor U1846 (N_1846,N_1762,N_1796);
or U1847 (N_1847,N_1759,N_1741);
nor U1848 (N_1848,N_1753,N_1769);
or U1849 (N_1849,N_1741,N_1760);
and U1850 (N_1850,N_1775,N_1747);
nand U1851 (N_1851,N_1785,N_1741);
nand U1852 (N_1852,N_1743,N_1764);
and U1853 (N_1853,N_1796,N_1753);
nand U1854 (N_1854,N_1755,N_1758);
nor U1855 (N_1855,N_1798,N_1750);
or U1856 (N_1856,N_1766,N_1763);
or U1857 (N_1857,N_1763,N_1740);
nand U1858 (N_1858,N_1752,N_1775);
or U1859 (N_1859,N_1752,N_1784);
nand U1860 (N_1860,N_1834,N_1817);
and U1861 (N_1861,N_1850,N_1818);
nand U1862 (N_1862,N_1821,N_1838);
nand U1863 (N_1863,N_1815,N_1853);
or U1864 (N_1864,N_1810,N_1830);
or U1865 (N_1865,N_1811,N_1849);
nor U1866 (N_1866,N_1801,N_1828);
nor U1867 (N_1867,N_1808,N_1807);
nor U1868 (N_1868,N_1809,N_1842);
and U1869 (N_1869,N_1813,N_1824);
nor U1870 (N_1870,N_1841,N_1802);
nand U1871 (N_1871,N_1825,N_1833);
or U1872 (N_1872,N_1805,N_1827);
and U1873 (N_1873,N_1820,N_1839);
nand U1874 (N_1874,N_1823,N_1837);
and U1875 (N_1875,N_1800,N_1856);
and U1876 (N_1876,N_1832,N_1843);
nor U1877 (N_1877,N_1844,N_1806);
nand U1878 (N_1878,N_1835,N_1819);
nand U1879 (N_1879,N_1826,N_1816);
or U1880 (N_1880,N_1836,N_1851);
or U1881 (N_1881,N_1822,N_1857);
and U1882 (N_1882,N_1829,N_1831);
and U1883 (N_1883,N_1846,N_1859);
nor U1884 (N_1884,N_1852,N_1840);
xnor U1885 (N_1885,N_1848,N_1803);
and U1886 (N_1886,N_1855,N_1845);
nor U1887 (N_1887,N_1847,N_1814);
or U1888 (N_1888,N_1854,N_1858);
and U1889 (N_1889,N_1804,N_1812);
and U1890 (N_1890,N_1805,N_1850);
or U1891 (N_1891,N_1837,N_1849);
nand U1892 (N_1892,N_1831,N_1834);
nand U1893 (N_1893,N_1808,N_1809);
or U1894 (N_1894,N_1854,N_1838);
and U1895 (N_1895,N_1818,N_1801);
nand U1896 (N_1896,N_1840,N_1845);
nand U1897 (N_1897,N_1808,N_1830);
nor U1898 (N_1898,N_1816,N_1830);
nor U1899 (N_1899,N_1851,N_1833);
nor U1900 (N_1900,N_1804,N_1850);
and U1901 (N_1901,N_1850,N_1857);
or U1902 (N_1902,N_1854,N_1804);
nand U1903 (N_1903,N_1849,N_1821);
and U1904 (N_1904,N_1847,N_1806);
nor U1905 (N_1905,N_1825,N_1806);
nand U1906 (N_1906,N_1808,N_1845);
and U1907 (N_1907,N_1812,N_1856);
nand U1908 (N_1908,N_1850,N_1827);
nand U1909 (N_1909,N_1802,N_1822);
nand U1910 (N_1910,N_1859,N_1830);
and U1911 (N_1911,N_1828,N_1855);
nor U1912 (N_1912,N_1833,N_1830);
nor U1913 (N_1913,N_1801,N_1811);
nor U1914 (N_1914,N_1853,N_1829);
nand U1915 (N_1915,N_1846,N_1849);
and U1916 (N_1916,N_1807,N_1832);
nand U1917 (N_1917,N_1856,N_1823);
nor U1918 (N_1918,N_1845,N_1807);
nand U1919 (N_1919,N_1844,N_1810);
nor U1920 (N_1920,N_1878,N_1887);
nor U1921 (N_1921,N_1865,N_1883);
nor U1922 (N_1922,N_1909,N_1912);
xnor U1923 (N_1923,N_1884,N_1860);
and U1924 (N_1924,N_1863,N_1908);
and U1925 (N_1925,N_1874,N_1868);
nor U1926 (N_1926,N_1904,N_1873);
and U1927 (N_1927,N_1881,N_1876);
nor U1928 (N_1928,N_1886,N_1903);
nor U1929 (N_1929,N_1872,N_1880);
nand U1930 (N_1930,N_1861,N_1906);
nor U1931 (N_1931,N_1894,N_1899);
nor U1932 (N_1932,N_1867,N_1911);
or U1933 (N_1933,N_1882,N_1888);
or U1934 (N_1934,N_1896,N_1897);
nand U1935 (N_1935,N_1862,N_1877);
nand U1936 (N_1936,N_1915,N_1879);
nor U1937 (N_1937,N_1918,N_1898);
nand U1938 (N_1938,N_1891,N_1919);
and U1939 (N_1939,N_1885,N_1870);
and U1940 (N_1940,N_1917,N_1864);
nand U1941 (N_1941,N_1905,N_1889);
nand U1942 (N_1942,N_1902,N_1900);
or U1943 (N_1943,N_1916,N_1866);
or U1944 (N_1944,N_1914,N_1910);
or U1945 (N_1945,N_1871,N_1875);
and U1946 (N_1946,N_1895,N_1913);
nor U1947 (N_1947,N_1893,N_1892);
and U1948 (N_1948,N_1907,N_1890);
nand U1949 (N_1949,N_1901,N_1869);
nand U1950 (N_1950,N_1877,N_1885);
or U1951 (N_1951,N_1897,N_1877);
nand U1952 (N_1952,N_1872,N_1877);
or U1953 (N_1953,N_1901,N_1872);
or U1954 (N_1954,N_1879,N_1910);
and U1955 (N_1955,N_1917,N_1872);
and U1956 (N_1956,N_1866,N_1903);
nor U1957 (N_1957,N_1914,N_1867);
and U1958 (N_1958,N_1873,N_1905);
nor U1959 (N_1959,N_1898,N_1873);
or U1960 (N_1960,N_1866,N_1870);
nor U1961 (N_1961,N_1869,N_1861);
nor U1962 (N_1962,N_1864,N_1887);
nor U1963 (N_1963,N_1913,N_1874);
nand U1964 (N_1964,N_1869,N_1866);
nor U1965 (N_1965,N_1875,N_1908);
nand U1966 (N_1966,N_1912,N_1910);
or U1967 (N_1967,N_1909,N_1875);
nand U1968 (N_1968,N_1877,N_1914);
or U1969 (N_1969,N_1910,N_1894);
nand U1970 (N_1970,N_1901,N_1918);
and U1971 (N_1971,N_1894,N_1903);
and U1972 (N_1972,N_1903,N_1877);
and U1973 (N_1973,N_1882,N_1883);
and U1974 (N_1974,N_1865,N_1871);
nand U1975 (N_1975,N_1876,N_1860);
or U1976 (N_1976,N_1884,N_1909);
or U1977 (N_1977,N_1863,N_1916);
nand U1978 (N_1978,N_1905,N_1892);
and U1979 (N_1979,N_1871,N_1903);
nor U1980 (N_1980,N_1975,N_1959);
nor U1981 (N_1981,N_1955,N_1963);
nand U1982 (N_1982,N_1956,N_1969);
xor U1983 (N_1983,N_1951,N_1948);
and U1984 (N_1984,N_1946,N_1923);
and U1985 (N_1985,N_1925,N_1929);
nand U1986 (N_1986,N_1965,N_1924);
or U1987 (N_1987,N_1926,N_1932);
or U1988 (N_1988,N_1978,N_1979);
and U1989 (N_1989,N_1940,N_1939);
nor U1990 (N_1990,N_1957,N_1960);
nand U1991 (N_1991,N_1937,N_1936);
xor U1992 (N_1992,N_1943,N_1968);
nor U1993 (N_1993,N_1921,N_1972);
nand U1994 (N_1994,N_1961,N_1949);
and U1995 (N_1995,N_1933,N_1942);
or U1996 (N_1996,N_1920,N_1930);
or U1997 (N_1997,N_1964,N_1922);
or U1998 (N_1998,N_1944,N_1970);
nor U1999 (N_1999,N_1928,N_1941);
and U2000 (N_2000,N_1931,N_1974);
and U2001 (N_2001,N_1952,N_1958);
and U2002 (N_2002,N_1967,N_1977);
or U2003 (N_2003,N_1966,N_1938);
and U2004 (N_2004,N_1953,N_1934);
nand U2005 (N_2005,N_1976,N_1971);
and U2006 (N_2006,N_1962,N_1935);
and U2007 (N_2007,N_1954,N_1947);
and U2008 (N_2008,N_1945,N_1973);
nor U2009 (N_2009,N_1927,N_1950);
nand U2010 (N_2010,N_1956,N_1966);
nor U2011 (N_2011,N_1970,N_1927);
and U2012 (N_2012,N_1928,N_1939);
or U2013 (N_2013,N_1964,N_1940);
nor U2014 (N_2014,N_1928,N_1949);
nor U2015 (N_2015,N_1932,N_1950);
or U2016 (N_2016,N_1965,N_1949);
or U2017 (N_2017,N_1968,N_1959);
and U2018 (N_2018,N_1921,N_1946);
and U2019 (N_2019,N_1953,N_1945);
nand U2020 (N_2020,N_1978,N_1972);
or U2021 (N_2021,N_1955,N_1941);
or U2022 (N_2022,N_1948,N_1950);
nand U2023 (N_2023,N_1932,N_1925);
or U2024 (N_2024,N_1959,N_1925);
and U2025 (N_2025,N_1959,N_1972);
or U2026 (N_2026,N_1971,N_1937);
nor U2027 (N_2027,N_1957,N_1936);
nor U2028 (N_2028,N_1977,N_1969);
or U2029 (N_2029,N_1971,N_1978);
nand U2030 (N_2030,N_1921,N_1959);
or U2031 (N_2031,N_1935,N_1963);
nand U2032 (N_2032,N_1952,N_1964);
and U2033 (N_2033,N_1933,N_1938);
nor U2034 (N_2034,N_1973,N_1964);
or U2035 (N_2035,N_1964,N_1961);
nor U2036 (N_2036,N_1927,N_1965);
or U2037 (N_2037,N_1925,N_1946);
nor U2038 (N_2038,N_1945,N_1972);
and U2039 (N_2039,N_1930,N_1960);
or U2040 (N_2040,N_2017,N_1986);
and U2041 (N_2041,N_1980,N_1998);
nand U2042 (N_2042,N_2031,N_2007);
or U2043 (N_2043,N_2005,N_1996);
nor U2044 (N_2044,N_2015,N_1995);
nand U2045 (N_2045,N_1992,N_1990);
nor U2046 (N_2046,N_2025,N_2023);
and U2047 (N_2047,N_2001,N_2011);
nand U2048 (N_2048,N_1985,N_2033);
nand U2049 (N_2049,N_2032,N_2012);
nor U2050 (N_2050,N_2038,N_1994);
nand U2051 (N_2051,N_2026,N_2004);
nand U2052 (N_2052,N_1988,N_2021);
and U2053 (N_2053,N_2009,N_2013);
nor U2054 (N_2054,N_2030,N_2020);
nand U2055 (N_2055,N_1997,N_1999);
or U2056 (N_2056,N_1983,N_2037);
nor U2057 (N_2057,N_2034,N_2029);
nand U2058 (N_2058,N_2016,N_1993);
and U2059 (N_2059,N_2028,N_1982);
and U2060 (N_2060,N_2027,N_1991);
or U2061 (N_2061,N_2010,N_2018);
and U2062 (N_2062,N_2000,N_2003);
xor U2063 (N_2063,N_2002,N_2022);
nor U2064 (N_2064,N_2039,N_2024);
or U2065 (N_2065,N_2035,N_1981);
or U2066 (N_2066,N_1989,N_1984);
nand U2067 (N_2067,N_2006,N_2008);
nor U2068 (N_2068,N_2036,N_1987);
nor U2069 (N_2069,N_2014,N_2019);
or U2070 (N_2070,N_2006,N_1999);
nor U2071 (N_2071,N_2031,N_2039);
nor U2072 (N_2072,N_1983,N_2038);
nand U2073 (N_2073,N_1988,N_1995);
or U2074 (N_2074,N_2030,N_1980);
or U2075 (N_2075,N_2025,N_1986);
nor U2076 (N_2076,N_2006,N_2002);
nand U2077 (N_2077,N_2021,N_2005);
and U2078 (N_2078,N_1995,N_1982);
or U2079 (N_2079,N_2000,N_2007);
or U2080 (N_2080,N_1988,N_2029);
nand U2081 (N_2081,N_2008,N_1983);
and U2082 (N_2082,N_1994,N_2039);
xor U2083 (N_2083,N_2031,N_2028);
and U2084 (N_2084,N_2035,N_2002);
or U2085 (N_2085,N_2034,N_2020);
nor U2086 (N_2086,N_1998,N_1986);
nor U2087 (N_2087,N_2008,N_1987);
and U2088 (N_2088,N_2005,N_1985);
xnor U2089 (N_2089,N_1982,N_1980);
xor U2090 (N_2090,N_1998,N_2004);
nor U2091 (N_2091,N_2023,N_1989);
nor U2092 (N_2092,N_1996,N_2031);
nor U2093 (N_2093,N_2009,N_2020);
nor U2094 (N_2094,N_1985,N_2032);
and U2095 (N_2095,N_1983,N_2022);
nand U2096 (N_2096,N_1981,N_2014);
nor U2097 (N_2097,N_1987,N_2025);
nor U2098 (N_2098,N_2035,N_2000);
nor U2099 (N_2099,N_2006,N_1998);
nand U2100 (N_2100,N_2057,N_2063);
nand U2101 (N_2101,N_2084,N_2062);
xor U2102 (N_2102,N_2099,N_2066);
nand U2103 (N_2103,N_2070,N_2047);
nor U2104 (N_2104,N_2044,N_2040);
and U2105 (N_2105,N_2059,N_2043);
or U2106 (N_2106,N_2051,N_2042);
nor U2107 (N_2107,N_2098,N_2058);
or U2108 (N_2108,N_2046,N_2056);
or U2109 (N_2109,N_2086,N_2077);
or U2110 (N_2110,N_2045,N_2061);
nand U2111 (N_2111,N_2075,N_2073);
or U2112 (N_2112,N_2097,N_2053);
xnor U2113 (N_2113,N_2082,N_2094);
nor U2114 (N_2114,N_2049,N_2074);
nor U2115 (N_2115,N_2079,N_2080);
or U2116 (N_2116,N_2068,N_2050);
and U2117 (N_2117,N_2065,N_2087);
nand U2118 (N_2118,N_2067,N_2090);
nand U2119 (N_2119,N_2071,N_2089);
nor U2120 (N_2120,N_2078,N_2096);
or U2121 (N_2121,N_2052,N_2085);
nand U2122 (N_2122,N_2041,N_2069);
xor U2123 (N_2123,N_2088,N_2093);
or U2124 (N_2124,N_2054,N_2060);
or U2125 (N_2125,N_2095,N_2092);
or U2126 (N_2126,N_2083,N_2055);
nor U2127 (N_2127,N_2048,N_2072);
and U2128 (N_2128,N_2076,N_2091);
nand U2129 (N_2129,N_2081,N_2064);
nor U2130 (N_2130,N_2097,N_2065);
or U2131 (N_2131,N_2081,N_2087);
nand U2132 (N_2132,N_2079,N_2085);
and U2133 (N_2133,N_2098,N_2048);
or U2134 (N_2134,N_2054,N_2051);
or U2135 (N_2135,N_2055,N_2060);
and U2136 (N_2136,N_2041,N_2086);
nor U2137 (N_2137,N_2087,N_2060);
nor U2138 (N_2138,N_2072,N_2061);
and U2139 (N_2139,N_2067,N_2095);
nand U2140 (N_2140,N_2072,N_2096);
nand U2141 (N_2141,N_2063,N_2099);
and U2142 (N_2142,N_2096,N_2069);
xnor U2143 (N_2143,N_2055,N_2067);
nand U2144 (N_2144,N_2082,N_2065);
and U2145 (N_2145,N_2041,N_2065);
nor U2146 (N_2146,N_2052,N_2048);
nor U2147 (N_2147,N_2071,N_2040);
and U2148 (N_2148,N_2098,N_2085);
nor U2149 (N_2149,N_2046,N_2093);
or U2150 (N_2150,N_2050,N_2061);
nor U2151 (N_2151,N_2064,N_2043);
nor U2152 (N_2152,N_2047,N_2090);
or U2153 (N_2153,N_2083,N_2044);
nand U2154 (N_2154,N_2098,N_2041);
nand U2155 (N_2155,N_2070,N_2073);
nand U2156 (N_2156,N_2049,N_2063);
nor U2157 (N_2157,N_2072,N_2043);
nor U2158 (N_2158,N_2084,N_2090);
or U2159 (N_2159,N_2075,N_2061);
nor U2160 (N_2160,N_2113,N_2119);
and U2161 (N_2161,N_2157,N_2138);
nor U2162 (N_2162,N_2135,N_2133);
and U2163 (N_2163,N_2154,N_2137);
and U2164 (N_2164,N_2151,N_2112);
and U2165 (N_2165,N_2131,N_2115);
or U2166 (N_2166,N_2139,N_2126);
or U2167 (N_2167,N_2124,N_2148);
nor U2168 (N_2168,N_2144,N_2125);
nand U2169 (N_2169,N_2107,N_2105);
and U2170 (N_2170,N_2129,N_2101);
nand U2171 (N_2171,N_2142,N_2109);
nor U2172 (N_2172,N_2110,N_2152);
or U2173 (N_2173,N_2116,N_2103);
nor U2174 (N_2174,N_2136,N_2153);
and U2175 (N_2175,N_2128,N_2117);
or U2176 (N_2176,N_2102,N_2106);
or U2177 (N_2177,N_2140,N_2149);
and U2178 (N_2178,N_2118,N_2132);
and U2179 (N_2179,N_2122,N_2146);
nor U2180 (N_2180,N_2159,N_2147);
or U2181 (N_2181,N_2156,N_2111);
and U2182 (N_2182,N_2130,N_2150);
nor U2183 (N_2183,N_2141,N_2120);
nor U2184 (N_2184,N_2127,N_2123);
or U2185 (N_2185,N_2143,N_2114);
nor U2186 (N_2186,N_2155,N_2108);
nor U2187 (N_2187,N_2100,N_2145);
and U2188 (N_2188,N_2134,N_2121);
and U2189 (N_2189,N_2104,N_2158);
nor U2190 (N_2190,N_2114,N_2152);
nand U2191 (N_2191,N_2109,N_2156);
nand U2192 (N_2192,N_2108,N_2146);
nor U2193 (N_2193,N_2150,N_2154);
nor U2194 (N_2194,N_2106,N_2127);
nor U2195 (N_2195,N_2139,N_2123);
or U2196 (N_2196,N_2148,N_2137);
nand U2197 (N_2197,N_2151,N_2113);
nor U2198 (N_2198,N_2117,N_2109);
or U2199 (N_2199,N_2102,N_2156);
and U2200 (N_2200,N_2153,N_2101);
nor U2201 (N_2201,N_2152,N_2107);
nand U2202 (N_2202,N_2147,N_2151);
and U2203 (N_2203,N_2118,N_2108);
nor U2204 (N_2204,N_2118,N_2110);
nand U2205 (N_2205,N_2112,N_2123);
or U2206 (N_2206,N_2104,N_2147);
nor U2207 (N_2207,N_2152,N_2108);
nor U2208 (N_2208,N_2101,N_2128);
or U2209 (N_2209,N_2146,N_2138);
and U2210 (N_2210,N_2155,N_2135);
nor U2211 (N_2211,N_2150,N_2139);
nor U2212 (N_2212,N_2150,N_2120);
nor U2213 (N_2213,N_2140,N_2132);
and U2214 (N_2214,N_2119,N_2141);
nor U2215 (N_2215,N_2101,N_2126);
or U2216 (N_2216,N_2146,N_2107);
or U2217 (N_2217,N_2152,N_2140);
and U2218 (N_2218,N_2133,N_2155);
nor U2219 (N_2219,N_2106,N_2150);
and U2220 (N_2220,N_2183,N_2219);
nor U2221 (N_2221,N_2190,N_2189);
nor U2222 (N_2222,N_2160,N_2216);
nor U2223 (N_2223,N_2200,N_2162);
or U2224 (N_2224,N_2205,N_2185);
or U2225 (N_2225,N_2209,N_2186);
or U2226 (N_2226,N_2187,N_2207);
and U2227 (N_2227,N_2170,N_2181);
and U2228 (N_2228,N_2168,N_2188);
nor U2229 (N_2229,N_2179,N_2196);
or U2230 (N_2230,N_2210,N_2174);
or U2231 (N_2231,N_2178,N_2184);
or U2232 (N_2232,N_2167,N_2215);
nand U2233 (N_2233,N_2212,N_2182);
nor U2234 (N_2234,N_2169,N_2161);
or U2235 (N_2235,N_2176,N_2165);
or U2236 (N_2236,N_2194,N_2193);
nand U2237 (N_2237,N_2177,N_2204);
or U2238 (N_2238,N_2173,N_2203);
and U2239 (N_2239,N_2201,N_2172);
nand U2240 (N_2240,N_2164,N_2175);
nand U2241 (N_2241,N_2213,N_2191);
nor U2242 (N_2242,N_2171,N_2218);
and U2243 (N_2243,N_2199,N_2180);
and U2244 (N_2244,N_2198,N_2195);
nor U2245 (N_2245,N_2202,N_2217);
nor U2246 (N_2246,N_2166,N_2211);
or U2247 (N_2247,N_2206,N_2163);
nor U2248 (N_2248,N_2214,N_2197);
nor U2249 (N_2249,N_2192,N_2208);
and U2250 (N_2250,N_2197,N_2179);
nor U2251 (N_2251,N_2176,N_2162);
nand U2252 (N_2252,N_2178,N_2217);
or U2253 (N_2253,N_2178,N_2188);
and U2254 (N_2254,N_2194,N_2167);
nand U2255 (N_2255,N_2184,N_2180);
or U2256 (N_2256,N_2178,N_2219);
and U2257 (N_2257,N_2177,N_2219);
xnor U2258 (N_2258,N_2196,N_2184);
or U2259 (N_2259,N_2160,N_2208);
or U2260 (N_2260,N_2202,N_2172);
and U2261 (N_2261,N_2167,N_2160);
or U2262 (N_2262,N_2177,N_2191);
nand U2263 (N_2263,N_2210,N_2182);
or U2264 (N_2264,N_2190,N_2197);
and U2265 (N_2265,N_2173,N_2199);
nand U2266 (N_2266,N_2188,N_2200);
nand U2267 (N_2267,N_2168,N_2175);
and U2268 (N_2268,N_2194,N_2199);
or U2269 (N_2269,N_2183,N_2165);
nand U2270 (N_2270,N_2219,N_2215);
and U2271 (N_2271,N_2219,N_2194);
or U2272 (N_2272,N_2215,N_2201);
nor U2273 (N_2273,N_2166,N_2217);
and U2274 (N_2274,N_2183,N_2205);
nand U2275 (N_2275,N_2164,N_2210);
nor U2276 (N_2276,N_2204,N_2168);
or U2277 (N_2277,N_2173,N_2197);
nor U2278 (N_2278,N_2204,N_2189);
or U2279 (N_2279,N_2192,N_2198);
nor U2280 (N_2280,N_2268,N_2236);
nand U2281 (N_2281,N_2241,N_2264);
nor U2282 (N_2282,N_2262,N_2228);
and U2283 (N_2283,N_2237,N_2256);
nand U2284 (N_2284,N_2240,N_2257);
nor U2285 (N_2285,N_2259,N_2271);
or U2286 (N_2286,N_2276,N_2250);
or U2287 (N_2287,N_2242,N_2252);
xor U2288 (N_2288,N_2253,N_2266);
nor U2289 (N_2289,N_2225,N_2226);
xnor U2290 (N_2290,N_2230,N_2221);
and U2291 (N_2291,N_2247,N_2244);
nand U2292 (N_2292,N_2272,N_2270);
nand U2293 (N_2293,N_2254,N_2231);
or U2294 (N_2294,N_2234,N_2261);
nand U2295 (N_2295,N_2251,N_2279);
nand U2296 (N_2296,N_2220,N_2233);
nand U2297 (N_2297,N_2235,N_2245);
nand U2298 (N_2298,N_2260,N_2277);
nand U2299 (N_2299,N_2227,N_2232);
nor U2300 (N_2300,N_2224,N_2278);
nand U2301 (N_2301,N_2249,N_2243);
nand U2302 (N_2302,N_2267,N_2238);
nor U2303 (N_2303,N_2265,N_2274);
nand U2304 (N_2304,N_2263,N_2223);
or U2305 (N_2305,N_2246,N_2258);
and U2306 (N_2306,N_2239,N_2273);
and U2307 (N_2307,N_2229,N_2275);
and U2308 (N_2308,N_2248,N_2222);
nor U2309 (N_2309,N_2255,N_2269);
and U2310 (N_2310,N_2264,N_2250);
and U2311 (N_2311,N_2235,N_2222);
nand U2312 (N_2312,N_2260,N_2273);
nand U2313 (N_2313,N_2257,N_2241);
and U2314 (N_2314,N_2239,N_2241);
nor U2315 (N_2315,N_2245,N_2253);
and U2316 (N_2316,N_2266,N_2240);
and U2317 (N_2317,N_2242,N_2278);
nand U2318 (N_2318,N_2273,N_2267);
nor U2319 (N_2319,N_2277,N_2225);
or U2320 (N_2320,N_2256,N_2261);
and U2321 (N_2321,N_2247,N_2258);
xor U2322 (N_2322,N_2246,N_2229);
and U2323 (N_2323,N_2275,N_2241);
nand U2324 (N_2324,N_2246,N_2228);
or U2325 (N_2325,N_2232,N_2221);
and U2326 (N_2326,N_2231,N_2239);
or U2327 (N_2327,N_2242,N_2255);
or U2328 (N_2328,N_2261,N_2221);
nor U2329 (N_2329,N_2242,N_2234);
nand U2330 (N_2330,N_2241,N_2245);
or U2331 (N_2331,N_2268,N_2253);
or U2332 (N_2332,N_2273,N_2243);
and U2333 (N_2333,N_2233,N_2249);
nand U2334 (N_2334,N_2270,N_2228);
and U2335 (N_2335,N_2234,N_2249);
and U2336 (N_2336,N_2259,N_2236);
and U2337 (N_2337,N_2268,N_2242);
or U2338 (N_2338,N_2237,N_2230);
or U2339 (N_2339,N_2221,N_2273);
and U2340 (N_2340,N_2323,N_2332);
or U2341 (N_2341,N_2291,N_2327);
and U2342 (N_2342,N_2325,N_2285);
nand U2343 (N_2343,N_2338,N_2289);
xor U2344 (N_2344,N_2306,N_2281);
and U2345 (N_2345,N_2337,N_2298);
nor U2346 (N_2346,N_2334,N_2286);
nor U2347 (N_2347,N_2280,N_2317);
xnor U2348 (N_2348,N_2292,N_2318);
nand U2349 (N_2349,N_2296,N_2321);
or U2350 (N_2350,N_2283,N_2336);
nand U2351 (N_2351,N_2300,N_2313);
nor U2352 (N_2352,N_2299,N_2324);
nand U2353 (N_2353,N_2331,N_2303);
nor U2354 (N_2354,N_2311,N_2316);
nand U2355 (N_2355,N_2295,N_2293);
and U2356 (N_2356,N_2335,N_2309);
nand U2357 (N_2357,N_2302,N_2282);
or U2358 (N_2358,N_2326,N_2315);
nor U2359 (N_2359,N_2307,N_2314);
nand U2360 (N_2360,N_2339,N_2294);
nor U2361 (N_2361,N_2288,N_2322);
nand U2362 (N_2362,N_2301,N_2312);
and U2363 (N_2363,N_2319,N_2305);
nor U2364 (N_2364,N_2329,N_2328);
nor U2365 (N_2365,N_2287,N_2320);
or U2366 (N_2366,N_2290,N_2330);
or U2367 (N_2367,N_2310,N_2297);
nand U2368 (N_2368,N_2333,N_2308);
nand U2369 (N_2369,N_2284,N_2304);
or U2370 (N_2370,N_2286,N_2325);
and U2371 (N_2371,N_2318,N_2285);
and U2372 (N_2372,N_2288,N_2326);
nor U2373 (N_2373,N_2310,N_2315);
nand U2374 (N_2374,N_2285,N_2299);
nand U2375 (N_2375,N_2313,N_2296);
nor U2376 (N_2376,N_2318,N_2325);
nor U2377 (N_2377,N_2323,N_2312);
nor U2378 (N_2378,N_2326,N_2318);
or U2379 (N_2379,N_2333,N_2289);
and U2380 (N_2380,N_2303,N_2308);
or U2381 (N_2381,N_2300,N_2303);
nor U2382 (N_2382,N_2314,N_2293);
and U2383 (N_2383,N_2305,N_2337);
nor U2384 (N_2384,N_2331,N_2287);
or U2385 (N_2385,N_2317,N_2316);
and U2386 (N_2386,N_2333,N_2299);
and U2387 (N_2387,N_2294,N_2292);
and U2388 (N_2388,N_2317,N_2292);
nor U2389 (N_2389,N_2324,N_2331);
nand U2390 (N_2390,N_2326,N_2319);
nor U2391 (N_2391,N_2327,N_2326);
nor U2392 (N_2392,N_2298,N_2308);
nand U2393 (N_2393,N_2333,N_2284);
and U2394 (N_2394,N_2311,N_2339);
or U2395 (N_2395,N_2337,N_2335);
or U2396 (N_2396,N_2338,N_2336);
xnor U2397 (N_2397,N_2296,N_2310);
nor U2398 (N_2398,N_2299,N_2306);
nor U2399 (N_2399,N_2336,N_2312);
nor U2400 (N_2400,N_2346,N_2344);
or U2401 (N_2401,N_2348,N_2395);
and U2402 (N_2402,N_2398,N_2388);
or U2403 (N_2403,N_2381,N_2359);
nor U2404 (N_2404,N_2391,N_2396);
or U2405 (N_2405,N_2357,N_2340);
and U2406 (N_2406,N_2387,N_2377);
nand U2407 (N_2407,N_2342,N_2373);
nor U2408 (N_2408,N_2386,N_2361);
and U2409 (N_2409,N_2366,N_2369);
or U2410 (N_2410,N_2371,N_2341);
nand U2411 (N_2411,N_2363,N_2380);
and U2412 (N_2412,N_2358,N_2354);
nor U2413 (N_2413,N_2374,N_2360);
nor U2414 (N_2414,N_2350,N_2384);
nand U2415 (N_2415,N_2389,N_2343);
nand U2416 (N_2416,N_2368,N_2347);
and U2417 (N_2417,N_2397,N_2370);
and U2418 (N_2418,N_2392,N_2382);
or U2419 (N_2419,N_2349,N_2378);
nand U2420 (N_2420,N_2376,N_2393);
nand U2421 (N_2421,N_2367,N_2364);
nand U2422 (N_2422,N_2351,N_2390);
nor U2423 (N_2423,N_2362,N_2372);
and U2424 (N_2424,N_2356,N_2365);
and U2425 (N_2425,N_2399,N_2383);
or U2426 (N_2426,N_2394,N_2352);
nor U2427 (N_2427,N_2375,N_2355);
or U2428 (N_2428,N_2345,N_2353);
or U2429 (N_2429,N_2385,N_2379);
and U2430 (N_2430,N_2346,N_2384);
and U2431 (N_2431,N_2367,N_2383);
or U2432 (N_2432,N_2367,N_2388);
and U2433 (N_2433,N_2383,N_2359);
or U2434 (N_2434,N_2398,N_2361);
nand U2435 (N_2435,N_2368,N_2344);
nand U2436 (N_2436,N_2363,N_2345);
nor U2437 (N_2437,N_2342,N_2367);
and U2438 (N_2438,N_2374,N_2353);
and U2439 (N_2439,N_2350,N_2344);
nor U2440 (N_2440,N_2379,N_2386);
nand U2441 (N_2441,N_2391,N_2386);
and U2442 (N_2442,N_2340,N_2375);
and U2443 (N_2443,N_2368,N_2394);
or U2444 (N_2444,N_2383,N_2342);
nand U2445 (N_2445,N_2373,N_2369);
nand U2446 (N_2446,N_2368,N_2377);
nand U2447 (N_2447,N_2388,N_2399);
and U2448 (N_2448,N_2386,N_2369);
nand U2449 (N_2449,N_2379,N_2384);
and U2450 (N_2450,N_2393,N_2383);
nand U2451 (N_2451,N_2348,N_2341);
nand U2452 (N_2452,N_2377,N_2372);
or U2453 (N_2453,N_2368,N_2382);
nor U2454 (N_2454,N_2353,N_2363);
nand U2455 (N_2455,N_2387,N_2365);
or U2456 (N_2456,N_2343,N_2356);
and U2457 (N_2457,N_2399,N_2386);
nand U2458 (N_2458,N_2392,N_2388);
nor U2459 (N_2459,N_2371,N_2390);
or U2460 (N_2460,N_2452,N_2421);
xnor U2461 (N_2461,N_2424,N_2416);
nand U2462 (N_2462,N_2455,N_2439);
nand U2463 (N_2463,N_2426,N_2407);
nor U2464 (N_2464,N_2411,N_2403);
or U2465 (N_2465,N_2406,N_2429);
and U2466 (N_2466,N_2427,N_2431);
nand U2467 (N_2467,N_2402,N_2413);
and U2468 (N_2468,N_2459,N_2437);
xnor U2469 (N_2469,N_2438,N_2445);
nand U2470 (N_2470,N_2400,N_2441);
nor U2471 (N_2471,N_2454,N_2430);
nand U2472 (N_2472,N_2401,N_2446);
nand U2473 (N_2473,N_2448,N_2419);
nor U2474 (N_2474,N_2434,N_2435);
and U2475 (N_2475,N_2423,N_2422);
nor U2476 (N_2476,N_2451,N_2425);
nand U2477 (N_2477,N_2453,N_2440);
or U2478 (N_2478,N_2456,N_2405);
nor U2479 (N_2479,N_2457,N_2458);
nor U2480 (N_2480,N_2433,N_2444);
and U2481 (N_2481,N_2408,N_2449);
or U2482 (N_2482,N_2417,N_2404);
nand U2483 (N_2483,N_2450,N_2414);
nand U2484 (N_2484,N_2443,N_2436);
and U2485 (N_2485,N_2412,N_2432);
and U2486 (N_2486,N_2410,N_2409);
nor U2487 (N_2487,N_2418,N_2447);
or U2488 (N_2488,N_2420,N_2428);
nand U2489 (N_2489,N_2442,N_2415);
nor U2490 (N_2490,N_2455,N_2432);
nand U2491 (N_2491,N_2443,N_2446);
and U2492 (N_2492,N_2455,N_2458);
nand U2493 (N_2493,N_2448,N_2429);
and U2494 (N_2494,N_2421,N_2440);
nor U2495 (N_2495,N_2437,N_2450);
nor U2496 (N_2496,N_2402,N_2443);
nor U2497 (N_2497,N_2435,N_2451);
nor U2498 (N_2498,N_2444,N_2402);
xor U2499 (N_2499,N_2426,N_2412);
nand U2500 (N_2500,N_2401,N_2442);
nor U2501 (N_2501,N_2456,N_2438);
nor U2502 (N_2502,N_2423,N_2427);
nor U2503 (N_2503,N_2427,N_2426);
nor U2504 (N_2504,N_2450,N_2429);
or U2505 (N_2505,N_2443,N_2412);
or U2506 (N_2506,N_2446,N_2429);
nor U2507 (N_2507,N_2429,N_2428);
or U2508 (N_2508,N_2440,N_2409);
or U2509 (N_2509,N_2452,N_2420);
and U2510 (N_2510,N_2416,N_2412);
or U2511 (N_2511,N_2408,N_2454);
nor U2512 (N_2512,N_2448,N_2447);
and U2513 (N_2513,N_2451,N_2449);
and U2514 (N_2514,N_2434,N_2438);
or U2515 (N_2515,N_2401,N_2439);
and U2516 (N_2516,N_2427,N_2456);
or U2517 (N_2517,N_2430,N_2407);
and U2518 (N_2518,N_2434,N_2457);
nor U2519 (N_2519,N_2437,N_2444);
and U2520 (N_2520,N_2484,N_2462);
nand U2521 (N_2521,N_2469,N_2481);
or U2522 (N_2522,N_2468,N_2519);
or U2523 (N_2523,N_2512,N_2460);
and U2524 (N_2524,N_2471,N_2477);
nand U2525 (N_2525,N_2473,N_2514);
nand U2526 (N_2526,N_2500,N_2506);
or U2527 (N_2527,N_2502,N_2504);
nor U2528 (N_2528,N_2518,N_2501);
nand U2529 (N_2529,N_2507,N_2494);
nand U2530 (N_2530,N_2496,N_2510);
and U2531 (N_2531,N_2492,N_2516);
nand U2532 (N_2532,N_2491,N_2478);
and U2533 (N_2533,N_2511,N_2508);
and U2534 (N_2534,N_2517,N_2474);
and U2535 (N_2535,N_2515,N_2472);
and U2536 (N_2536,N_2488,N_2467);
and U2537 (N_2537,N_2498,N_2490);
nand U2538 (N_2538,N_2493,N_2485);
nand U2539 (N_2539,N_2483,N_2509);
nor U2540 (N_2540,N_2497,N_2480);
nor U2541 (N_2541,N_2487,N_2513);
nand U2542 (N_2542,N_2479,N_2476);
xor U2543 (N_2543,N_2475,N_2466);
or U2544 (N_2544,N_2495,N_2489);
nand U2545 (N_2545,N_2470,N_2486);
or U2546 (N_2546,N_2464,N_2503);
nand U2547 (N_2547,N_2499,N_2465);
xnor U2548 (N_2548,N_2482,N_2463);
and U2549 (N_2549,N_2505,N_2461);
nor U2550 (N_2550,N_2473,N_2516);
and U2551 (N_2551,N_2508,N_2474);
and U2552 (N_2552,N_2465,N_2462);
or U2553 (N_2553,N_2487,N_2466);
nand U2554 (N_2554,N_2467,N_2463);
nand U2555 (N_2555,N_2513,N_2510);
or U2556 (N_2556,N_2476,N_2512);
and U2557 (N_2557,N_2486,N_2467);
nor U2558 (N_2558,N_2506,N_2475);
and U2559 (N_2559,N_2508,N_2482);
nand U2560 (N_2560,N_2481,N_2468);
nor U2561 (N_2561,N_2489,N_2502);
nor U2562 (N_2562,N_2513,N_2486);
nand U2563 (N_2563,N_2513,N_2473);
and U2564 (N_2564,N_2477,N_2466);
nor U2565 (N_2565,N_2463,N_2507);
nand U2566 (N_2566,N_2498,N_2494);
and U2567 (N_2567,N_2499,N_2469);
nand U2568 (N_2568,N_2470,N_2504);
nand U2569 (N_2569,N_2466,N_2470);
nor U2570 (N_2570,N_2487,N_2503);
nor U2571 (N_2571,N_2471,N_2478);
or U2572 (N_2572,N_2515,N_2519);
or U2573 (N_2573,N_2471,N_2495);
and U2574 (N_2574,N_2481,N_2489);
xor U2575 (N_2575,N_2476,N_2472);
or U2576 (N_2576,N_2504,N_2469);
or U2577 (N_2577,N_2474,N_2514);
nor U2578 (N_2578,N_2480,N_2462);
and U2579 (N_2579,N_2467,N_2479);
nand U2580 (N_2580,N_2579,N_2544);
nor U2581 (N_2581,N_2530,N_2545);
or U2582 (N_2582,N_2537,N_2572);
nor U2583 (N_2583,N_2557,N_2566);
or U2584 (N_2584,N_2525,N_2555);
nor U2585 (N_2585,N_2553,N_2539);
nand U2586 (N_2586,N_2568,N_2560);
nor U2587 (N_2587,N_2559,N_2527);
and U2588 (N_2588,N_2577,N_2538);
nor U2589 (N_2589,N_2548,N_2542);
nand U2590 (N_2590,N_2526,N_2534);
nand U2591 (N_2591,N_2521,N_2573);
nand U2592 (N_2592,N_2524,N_2520);
and U2593 (N_2593,N_2565,N_2532);
nand U2594 (N_2594,N_2575,N_2533);
or U2595 (N_2595,N_2550,N_2523);
xor U2596 (N_2596,N_2569,N_2541);
nor U2597 (N_2597,N_2543,N_2536);
nand U2598 (N_2598,N_2546,N_2540);
nand U2599 (N_2599,N_2567,N_2578);
nor U2600 (N_2600,N_2571,N_2535);
or U2601 (N_2601,N_2522,N_2570);
nor U2602 (N_2602,N_2558,N_2551);
and U2603 (N_2603,N_2561,N_2564);
or U2604 (N_2604,N_2563,N_2574);
nor U2605 (N_2605,N_2556,N_2531);
nand U2606 (N_2606,N_2552,N_2549);
nor U2607 (N_2607,N_2547,N_2528);
nor U2608 (N_2608,N_2529,N_2562);
and U2609 (N_2609,N_2554,N_2576);
or U2610 (N_2610,N_2520,N_2570);
nand U2611 (N_2611,N_2557,N_2530);
or U2612 (N_2612,N_2570,N_2568);
nor U2613 (N_2613,N_2568,N_2546);
nor U2614 (N_2614,N_2534,N_2562);
and U2615 (N_2615,N_2526,N_2536);
nor U2616 (N_2616,N_2543,N_2528);
nor U2617 (N_2617,N_2555,N_2541);
nand U2618 (N_2618,N_2543,N_2575);
nand U2619 (N_2619,N_2533,N_2539);
nor U2620 (N_2620,N_2576,N_2549);
nor U2621 (N_2621,N_2521,N_2579);
xor U2622 (N_2622,N_2532,N_2539);
nor U2623 (N_2623,N_2526,N_2542);
nor U2624 (N_2624,N_2528,N_2576);
or U2625 (N_2625,N_2520,N_2548);
nand U2626 (N_2626,N_2554,N_2525);
and U2627 (N_2627,N_2532,N_2522);
or U2628 (N_2628,N_2578,N_2545);
nand U2629 (N_2629,N_2541,N_2525);
nand U2630 (N_2630,N_2576,N_2534);
nand U2631 (N_2631,N_2525,N_2567);
and U2632 (N_2632,N_2560,N_2522);
and U2633 (N_2633,N_2521,N_2562);
nand U2634 (N_2634,N_2525,N_2549);
or U2635 (N_2635,N_2545,N_2571);
and U2636 (N_2636,N_2544,N_2557);
or U2637 (N_2637,N_2576,N_2556);
nand U2638 (N_2638,N_2566,N_2576);
nor U2639 (N_2639,N_2564,N_2522);
or U2640 (N_2640,N_2601,N_2591);
and U2641 (N_2641,N_2611,N_2585);
and U2642 (N_2642,N_2632,N_2590);
and U2643 (N_2643,N_2604,N_2597);
nand U2644 (N_2644,N_2635,N_2603);
or U2645 (N_2645,N_2636,N_2615);
and U2646 (N_2646,N_2620,N_2633);
or U2647 (N_2647,N_2593,N_2582);
nand U2648 (N_2648,N_2602,N_2617);
or U2649 (N_2649,N_2592,N_2630);
or U2650 (N_2650,N_2619,N_2618);
and U2651 (N_2651,N_2606,N_2613);
and U2652 (N_2652,N_2587,N_2584);
xnor U2653 (N_2653,N_2638,N_2588);
and U2654 (N_2654,N_2628,N_2596);
nand U2655 (N_2655,N_2627,N_2634);
or U2656 (N_2656,N_2589,N_2605);
xnor U2657 (N_2657,N_2624,N_2622);
nor U2658 (N_2658,N_2608,N_2616);
nand U2659 (N_2659,N_2598,N_2583);
or U2660 (N_2660,N_2581,N_2612);
nor U2661 (N_2661,N_2631,N_2600);
and U2662 (N_2662,N_2607,N_2594);
xnor U2663 (N_2663,N_2637,N_2639);
and U2664 (N_2664,N_2580,N_2621);
nor U2665 (N_2665,N_2626,N_2614);
and U2666 (N_2666,N_2629,N_2595);
and U2667 (N_2667,N_2625,N_2586);
nand U2668 (N_2668,N_2610,N_2623);
and U2669 (N_2669,N_2609,N_2599);
xnor U2670 (N_2670,N_2633,N_2616);
nor U2671 (N_2671,N_2619,N_2603);
nand U2672 (N_2672,N_2604,N_2581);
or U2673 (N_2673,N_2616,N_2624);
nor U2674 (N_2674,N_2623,N_2637);
nor U2675 (N_2675,N_2613,N_2600);
nand U2676 (N_2676,N_2622,N_2607);
and U2677 (N_2677,N_2594,N_2627);
nor U2678 (N_2678,N_2618,N_2625);
and U2679 (N_2679,N_2608,N_2603);
xor U2680 (N_2680,N_2605,N_2625);
nor U2681 (N_2681,N_2582,N_2628);
and U2682 (N_2682,N_2596,N_2625);
nand U2683 (N_2683,N_2621,N_2613);
nand U2684 (N_2684,N_2587,N_2624);
nand U2685 (N_2685,N_2618,N_2610);
nor U2686 (N_2686,N_2597,N_2621);
or U2687 (N_2687,N_2613,N_2622);
nor U2688 (N_2688,N_2616,N_2591);
nand U2689 (N_2689,N_2631,N_2619);
nand U2690 (N_2690,N_2602,N_2631);
or U2691 (N_2691,N_2584,N_2595);
nand U2692 (N_2692,N_2637,N_2636);
nand U2693 (N_2693,N_2603,N_2606);
and U2694 (N_2694,N_2607,N_2616);
or U2695 (N_2695,N_2598,N_2591);
nand U2696 (N_2696,N_2593,N_2626);
xnor U2697 (N_2697,N_2620,N_2590);
nand U2698 (N_2698,N_2594,N_2635);
nand U2699 (N_2699,N_2623,N_2594);
and U2700 (N_2700,N_2677,N_2699);
and U2701 (N_2701,N_2660,N_2641);
and U2702 (N_2702,N_2643,N_2661);
and U2703 (N_2703,N_2696,N_2653);
and U2704 (N_2704,N_2646,N_2666);
nor U2705 (N_2705,N_2680,N_2648);
and U2706 (N_2706,N_2670,N_2668);
nand U2707 (N_2707,N_2692,N_2684);
or U2708 (N_2708,N_2694,N_2688);
nand U2709 (N_2709,N_2659,N_2664);
nor U2710 (N_2710,N_2691,N_2651);
and U2711 (N_2711,N_2678,N_2689);
or U2712 (N_2712,N_2652,N_2656);
and U2713 (N_2713,N_2673,N_2655);
nor U2714 (N_2714,N_2690,N_2650);
nand U2715 (N_2715,N_2686,N_2654);
or U2716 (N_2716,N_2682,N_2685);
xor U2717 (N_2717,N_2647,N_2662);
nand U2718 (N_2718,N_2681,N_2671);
nor U2719 (N_2719,N_2669,N_2645);
nand U2720 (N_2720,N_2644,N_2640);
or U2721 (N_2721,N_2658,N_2675);
or U2722 (N_2722,N_2698,N_2695);
nand U2723 (N_2723,N_2649,N_2674);
or U2724 (N_2724,N_2679,N_2683);
and U2725 (N_2725,N_2657,N_2665);
or U2726 (N_2726,N_2642,N_2687);
nand U2727 (N_2727,N_2663,N_2667);
nor U2728 (N_2728,N_2693,N_2697);
nor U2729 (N_2729,N_2672,N_2676);
or U2730 (N_2730,N_2695,N_2656);
nand U2731 (N_2731,N_2669,N_2675);
nor U2732 (N_2732,N_2661,N_2649);
and U2733 (N_2733,N_2687,N_2643);
nand U2734 (N_2734,N_2650,N_2666);
and U2735 (N_2735,N_2660,N_2689);
nand U2736 (N_2736,N_2643,N_2654);
nand U2737 (N_2737,N_2663,N_2691);
nand U2738 (N_2738,N_2694,N_2689);
or U2739 (N_2739,N_2644,N_2687);
nand U2740 (N_2740,N_2687,N_2650);
nor U2741 (N_2741,N_2646,N_2669);
or U2742 (N_2742,N_2677,N_2658);
or U2743 (N_2743,N_2654,N_2693);
nor U2744 (N_2744,N_2667,N_2652);
nor U2745 (N_2745,N_2679,N_2655);
nor U2746 (N_2746,N_2643,N_2670);
nand U2747 (N_2747,N_2669,N_2692);
nor U2748 (N_2748,N_2678,N_2674);
nor U2749 (N_2749,N_2670,N_2684);
and U2750 (N_2750,N_2642,N_2664);
and U2751 (N_2751,N_2650,N_2645);
nor U2752 (N_2752,N_2696,N_2649);
or U2753 (N_2753,N_2676,N_2687);
or U2754 (N_2754,N_2648,N_2663);
or U2755 (N_2755,N_2685,N_2660);
or U2756 (N_2756,N_2692,N_2679);
and U2757 (N_2757,N_2664,N_2645);
nor U2758 (N_2758,N_2671,N_2675);
and U2759 (N_2759,N_2641,N_2666);
and U2760 (N_2760,N_2737,N_2724);
or U2761 (N_2761,N_2706,N_2753);
nor U2762 (N_2762,N_2714,N_2748);
nor U2763 (N_2763,N_2715,N_2702);
xnor U2764 (N_2764,N_2739,N_2759);
nand U2765 (N_2765,N_2704,N_2722);
or U2766 (N_2766,N_2708,N_2743);
and U2767 (N_2767,N_2745,N_2735);
xor U2768 (N_2768,N_2710,N_2711);
or U2769 (N_2769,N_2754,N_2729);
and U2770 (N_2770,N_2725,N_2756);
or U2771 (N_2771,N_2738,N_2751);
nor U2772 (N_2772,N_2726,N_2744);
and U2773 (N_2773,N_2713,N_2727);
or U2774 (N_2774,N_2707,N_2705);
nand U2775 (N_2775,N_2747,N_2717);
nand U2776 (N_2776,N_2701,N_2740);
nand U2777 (N_2777,N_2741,N_2700);
nand U2778 (N_2778,N_2721,N_2733);
nand U2779 (N_2779,N_2746,N_2716);
or U2780 (N_2780,N_2718,N_2742);
or U2781 (N_2781,N_2728,N_2723);
nand U2782 (N_2782,N_2750,N_2731);
nor U2783 (N_2783,N_2732,N_2749);
or U2784 (N_2784,N_2734,N_2703);
nor U2785 (N_2785,N_2755,N_2719);
and U2786 (N_2786,N_2752,N_2709);
nor U2787 (N_2787,N_2730,N_2758);
or U2788 (N_2788,N_2712,N_2736);
nor U2789 (N_2789,N_2720,N_2757);
nand U2790 (N_2790,N_2745,N_2711);
xnor U2791 (N_2791,N_2743,N_2745);
nand U2792 (N_2792,N_2714,N_2738);
nor U2793 (N_2793,N_2754,N_2720);
nor U2794 (N_2794,N_2734,N_2733);
nor U2795 (N_2795,N_2707,N_2712);
and U2796 (N_2796,N_2707,N_2746);
nor U2797 (N_2797,N_2733,N_2740);
nand U2798 (N_2798,N_2741,N_2753);
nand U2799 (N_2799,N_2741,N_2723);
or U2800 (N_2800,N_2704,N_2752);
and U2801 (N_2801,N_2739,N_2711);
nand U2802 (N_2802,N_2722,N_2751);
and U2803 (N_2803,N_2726,N_2708);
and U2804 (N_2804,N_2707,N_2722);
nor U2805 (N_2805,N_2720,N_2733);
or U2806 (N_2806,N_2754,N_2716);
nor U2807 (N_2807,N_2728,N_2759);
and U2808 (N_2808,N_2735,N_2715);
nor U2809 (N_2809,N_2700,N_2759);
or U2810 (N_2810,N_2712,N_2721);
and U2811 (N_2811,N_2745,N_2719);
or U2812 (N_2812,N_2744,N_2755);
nand U2813 (N_2813,N_2738,N_2726);
or U2814 (N_2814,N_2701,N_2754);
nand U2815 (N_2815,N_2744,N_2743);
and U2816 (N_2816,N_2735,N_2738);
and U2817 (N_2817,N_2705,N_2728);
nor U2818 (N_2818,N_2709,N_2754);
nor U2819 (N_2819,N_2737,N_2709);
and U2820 (N_2820,N_2764,N_2791);
nor U2821 (N_2821,N_2801,N_2803);
and U2822 (N_2822,N_2799,N_2795);
or U2823 (N_2823,N_2774,N_2798);
nand U2824 (N_2824,N_2771,N_2778);
or U2825 (N_2825,N_2814,N_2782);
or U2826 (N_2826,N_2760,N_2805);
or U2827 (N_2827,N_2768,N_2813);
and U2828 (N_2828,N_2786,N_2815);
and U2829 (N_2829,N_2781,N_2806);
nor U2830 (N_2830,N_2796,N_2785);
and U2831 (N_2831,N_2800,N_2765);
nor U2832 (N_2832,N_2788,N_2787);
or U2833 (N_2833,N_2810,N_2770);
nand U2834 (N_2834,N_2776,N_2780);
nor U2835 (N_2835,N_2817,N_2793);
and U2836 (N_2836,N_2769,N_2804);
nand U2837 (N_2837,N_2816,N_2767);
and U2838 (N_2838,N_2783,N_2811);
and U2839 (N_2839,N_2789,N_2807);
and U2840 (N_2840,N_2773,N_2808);
nor U2841 (N_2841,N_2763,N_2818);
nand U2842 (N_2842,N_2819,N_2777);
and U2843 (N_2843,N_2772,N_2762);
nor U2844 (N_2844,N_2792,N_2766);
nand U2845 (N_2845,N_2784,N_2794);
and U2846 (N_2846,N_2779,N_2809);
nand U2847 (N_2847,N_2790,N_2812);
xnor U2848 (N_2848,N_2802,N_2775);
nand U2849 (N_2849,N_2761,N_2797);
nor U2850 (N_2850,N_2807,N_2797);
or U2851 (N_2851,N_2779,N_2818);
nand U2852 (N_2852,N_2788,N_2808);
and U2853 (N_2853,N_2760,N_2806);
or U2854 (N_2854,N_2783,N_2784);
nor U2855 (N_2855,N_2817,N_2770);
nor U2856 (N_2856,N_2805,N_2792);
nand U2857 (N_2857,N_2816,N_2776);
and U2858 (N_2858,N_2806,N_2779);
nand U2859 (N_2859,N_2777,N_2816);
and U2860 (N_2860,N_2781,N_2777);
and U2861 (N_2861,N_2812,N_2779);
or U2862 (N_2862,N_2764,N_2771);
xor U2863 (N_2863,N_2787,N_2791);
or U2864 (N_2864,N_2807,N_2795);
and U2865 (N_2865,N_2800,N_2811);
nand U2866 (N_2866,N_2803,N_2819);
and U2867 (N_2867,N_2781,N_2765);
and U2868 (N_2868,N_2807,N_2775);
and U2869 (N_2869,N_2808,N_2819);
nor U2870 (N_2870,N_2805,N_2788);
and U2871 (N_2871,N_2818,N_2765);
or U2872 (N_2872,N_2788,N_2762);
nand U2873 (N_2873,N_2802,N_2772);
nor U2874 (N_2874,N_2800,N_2817);
nor U2875 (N_2875,N_2783,N_2786);
xnor U2876 (N_2876,N_2807,N_2812);
xnor U2877 (N_2877,N_2795,N_2777);
nand U2878 (N_2878,N_2808,N_2799);
nand U2879 (N_2879,N_2814,N_2793);
nand U2880 (N_2880,N_2876,N_2860);
nor U2881 (N_2881,N_2854,N_2863);
nand U2882 (N_2882,N_2828,N_2832);
nand U2883 (N_2883,N_2871,N_2870);
or U2884 (N_2884,N_2850,N_2874);
nand U2885 (N_2885,N_2858,N_2820);
nor U2886 (N_2886,N_2864,N_2865);
and U2887 (N_2887,N_2878,N_2829);
and U2888 (N_2888,N_2867,N_2831);
and U2889 (N_2889,N_2847,N_2843);
or U2890 (N_2890,N_2835,N_2851);
nand U2891 (N_2891,N_2868,N_2857);
or U2892 (N_2892,N_2862,N_2872);
nand U2893 (N_2893,N_2845,N_2840);
and U2894 (N_2894,N_2856,N_2846);
nor U2895 (N_2895,N_2877,N_2837);
and U2896 (N_2896,N_2834,N_2824);
nand U2897 (N_2897,N_2833,N_2839);
or U2898 (N_2898,N_2852,N_2866);
or U2899 (N_2899,N_2848,N_2836);
nand U2900 (N_2900,N_2838,N_2849);
and U2901 (N_2901,N_2826,N_2875);
and U2902 (N_2902,N_2873,N_2821);
and U2903 (N_2903,N_2853,N_2830);
and U2904 (N_2904,N_2842,N_2869);
nor U2905 (N_2905,N_2827,N_2859);
nor U2906 (N_2906,N_2822,N_2823);
nor U2907 (N_2907,N_2879,N_2855);
and U2908 (N_2908,N_2825,N_2861);
nor U2909 (N_2909,N_2844,N_2841);
or U2910 (N_2910,N_2848,N_2872);
or U2911 (N_2911,N_2825,N_2866);
and U2912 (N_2912,N_2833,N_2878);
and U2913 (N_2913,N_2866,N_2828);
nand U2914 (N_2914,N_2831,N_2825);
or U2915 (N_2915,N_2870,N_2827);
and U2916 (N_2916,N_2847,N_2878);
xor U2917 (N_2917,N_2876,N_2872);
nand U2918 (N_2918,N_2876,N_2828);
nand U2919 (N_2919,N_2856,N_2840);
or U2920 (N_2920,N_2830,N_2858);
nand U2921 (N_2921,N_2864,N_2875);
nor U2922 (N_2922,N_2829,N_2867);
nand U2923 (N_2923,N_2851,N_2823);
and U2924 (N_2924,N_2843,N_2825);
and U2925 (N_2925,N_2848,N_2838);
nor U2926 (N_2926,N_2876,N_2877);
and U2927 (N_2927,N_2854,N_2875);
or U2928 (N_2928,N_2856,N_2828);
and U2929 (N_2929,N_2843,N_2855);
nand U2930 (N_2930,N_2829,N_2866);
nor U2931 (N_2931,N_2827,N_2846);
nor U2932 (N_2932,N_2836,N_2863);
nor U2933 (N_2933,N_2823,N_2853);
or U2934 (N_2934,N_2866,N_2876);
nor U2935 (N_2935,N_2852,N_2837);
and U2936 (N_2936,N_2857,N_2878);
nand U2937 (N_2937,N_2831,N_2824);
nor U2938 (N_2938,N_2864,N_2868);
and U2939 (N_2939,N_2824,N_2820);
xnor U2940 (N_2940,N_2909,N_2923);
nand U2941 (N_2941,N_2891,N_2926);
nand U2942 (N_2942,N_2934,N_2890);
nor U2943 (N_2943,N_2930,N_2902);
nand U2944 (N_2944,N_2903,N_2887);
nand U2945 (N_2945,N_2896,N_2911);
nor U2946 (N_2946,N_2888,N_2931);
nor U2947 (N_2947,N_2904,N_2915);
nand U2948 (N_2948,N_2917,N_2919);
and U2949 (N_2949,N_2937,N_2898);
or U2950 (N_2950,N_2921,N_2881);
or U2951 (N_2951,N_2916,N_2910);
or U2952 (N_2952,N_2907,N_2893);
nand U2953 (N_2953,N_2924,N_2929);
nand U2954 (N_2954,N_2883,N_2882);
nor U2955 (N_2955,N_2912,N_2894);
nand U2956 (N_2956,N_2938,N_2897);
or U2957 (N_2957,N_2928,N_2914);
or U2958 (N_2958,N_2901,N_2913);
nor U2959 (N_2959,N_2886,N_2922);
nor U2960 (N_2960,N_2889,N_2936);
and U2961 (N_2961,N_2892,N_2895);
nor U2962 (N_2962,N_2933,N_2918);
nor U2963 (N_2963,N_2906,N_2885);
nor U2964 (N_2964,N_2908,N_2900);
or U2965 (N_2965,N_2939,N_2899);
or U2966 (N_2966,N_2935,N_2920);
and U2967 (N_2967,N_2884,N_2925);
nand U2968 (N_2968,N_2932,N_2880);
nand U2969 (N_2969,N_2905,N_2927);
and U2970 (N_2970,N_2925,N_2906);
nand U2971 (N_2971,N_2909,N_2901);
or U2972 (N_2972,N_2907,N_2884);
nand U2973 (N_2973,N_2893,N_2932);
nand U2974 (N_2974,N_2907,N_2882);
and U2975 (N_2975,N_2902,N_2912);
nor U2976 (N_2976,N_2923,N_2935);
nor U2977 (N_2977,N_2912,N_2882);
and U2978 (N_2978,N_2921,N_2908);
and U2979 (N_2979,N_2911,N_2925);
nor U2980 (N_2980,N_2898,N_2897);
nand U2981 (N_2981,N_2926,N_2938);
nand U2982 (N_2982,N_2924,N_2902);
or U2983 (N_2983,N_2895,N_2921);
nand U2984 (N_2984,N_2901,N_2921);
nand U2985 (N_2985,N_2913,N_2914);
nor U2986 (N_2986,N_2935,N_2936);
nand U2987 (N_2987,N_2921,N_2927);
nand U2988 (N_2988,N_2895,N_2934);
and U2989 (N_2989,N_2903,N_2936);
nor U2990 (N_2990,N_2904,N_2884);
or U2991 (N_2991,N_2928,N_2921);
nand U2992 (N_2992,N_2909,N_2880);
nand U2993 (N_2993,N_2887,N_2905);
nor U2994 (N_2994,N_2923,N_2930);
nor U2995 (N_2995,N_2922,N_2929);
nand U2996 (N_2996,N_2929,N_2935);
nor U2997 (N_2997,N_2925,N_2890);
nor U2998 (N_2998,N_2920,N_2932);
nand U2999 (N_2999,N_2937,N_2933);
nand UO_0 (O_0,N_2997,N_2994);
nand UO_1 (O_1,N_2990,N_2993);
or UO_2 (O_2,N_2998,N_2961);
nor UO_3 (O_3,N_2952,N_2948);
nor UO_4 (O_4,N_2958,N_2955);
nand UO_5 (O_5,N_2968,N_2969);
nor UO_6 (O_6,N_2962,N_2959);
nand UO_7 (O_7,N_2940,N_2944);
and UO_8 (O_8,N_2995,N_2967);
xnor UO_9 (O_9,N_2970,N_2957);
or UO_10 (O_10,N_2991,N_2947);
and UO_11 (O_11,N_2981,N_2984);
or UO_12 (O_12,N_2996,N_2988);
nor UO_13 (O_13,N_2999,N_2943);
and UO_14 (O_14,N_2986,N_2964);
nand UO_15 (O_15,N_2976,N_2974);
or UO_16 (O_16,N_2945,N_2963);
nor UO_17 (O_17,N_2979,N_2949);
and UO_18 (O_18,N_2950,N_2978);
and UO_19 (O_19,N_2975,N_2953);
or UO_20 (O_20,N_2980,N_2965);
and UO_21 (O_21,N_2941,N_2942);
nor UO_22 (O_22,N_2956,N_2972);
or UO_23 (O_23,N_2982,N_2946);
nand UO_24 (O_24,N_2966,N_2960);
nand UO_25 (O_25,N_2983,N_2989);
or UO_26 (O_26,N_2985,N_2954);
nor UO_27 (O_27,N_2951,N_2977);
nor UO_28 (O_28,N_2992,N_2973);
nand UO_29 (O_29,N_2987,N_2971);
nand UO_30 (O_30,N_2997,N_2986);
or UO_31 (O_31,N_2957,N_2961);
or UO_32 (O_32,N_2940,N_2994);
and UO_33 (O_33,N_2961,N_2986);
and UO_34 (O_34,N_2979,N_2983);
or UO_35 (O_35,N_2988,N_2994);
xnor UO_36 (O_36,N_2988,N_2970);
or UO_37 (O_37,N_2968,N_2956);
or UO_38 (O_38,N_2982,N_2956);
xor UO_39 (O_39,N_2995,N_2952);
nor UO_40 (O_40,N_2973,N_2976);
nand UO_41 (O_41,N_2993,N_2967);
and UO_42 (O_42,N_2966,N_2962);
nor UO_43 (O_43,N_2972,N_2988);
nor UO_44 (O_44,N_2961,N_2943);
and UO_45 (O_45,N_2958,N_2961);
and UO_46 (O_46,N_2956,N_2940);
nor UO_47 (O_47,N_2985,N_2942);
nand UO_48 (O_48,N_2941,N_2983);
nor UO_49 (O_49,N_2944,N_2978);
nand UO_50 (O_50,N_2974,N_2943);
nand UO_51 (O_51,N_2958,N_2960);
or UO_52 (O_52,N_2955,N_2991);
nor UO_53 (O_53,N_2994,N_2973);
and UO_54 (O_54,N_2981,N_2966);
nor UO_55 (O_55,N_2943,N_2966);
nor UO_56 (O_56,N_2984,N_2977);
nor UO_57 (O_57,N_2971,N_2995);
or UO_58 (O_58,N_2998,N_2978);
nand UO_59 (O_59,N_2947,N_2965);
and UO_60 (O_60,N_2986,N_2984);
nand UO_61 (O_61,N_2956,N_2955);
or UO_62 (O_62,N_2955,N_2988);
or UO_63 (O_63,N_2975,N_2972);
nand UO_64 (O_64,N_2997,N_2984);
nand UO_65 (O_65,N_2969,N_2996);
nor UO_66 (O_66,N_2991,N_2961);
nand UO_67 (O_67,N_2945,N_2995);
nand UO_68 (O_68,N_2981,N_2940);
or UO_69 (O_69,N_2984,N_2985);
nand UO_70 (O_70,N_2969,N_2987);
or UO_71 (O_71,N_2986,N_2958);
and UO_72 (O_72,N_2941,N_2980);
and UO_73 (O_73,N_2940,N_2992);
or UO_74 (O_74,N_2964,N_2954);
nand UO_75 (O_75,N_2972,N_2989);
nand UO_76 (O_76,N_2995,N_2946);
or UO_77 (O_77,N_2972,N_2979);
and UO_78 (O_78,N_2988,N_2982);
and UO_79 (O_79,N_2993,N_2966);
or UO_80 (O_80,N_2948,N_2954);
or UO_81 (O_81,N_2985,N_2948);
nand UO_82 (O_82,N_2952,N_2940);
nand UO_83 (O_83,N_2992,N_2964);
nor UO_84 (O_84,N_2954,N_2988);
nand UO_85 (O_85,N_2955,N_2999);
nand UO_86 (O_86,N_2950,N_2976);
nand UO_87 (O_87,N_2962,N_2968);
nand UO_88 (O_88,N_2964,N_2969);
or UO_89 (O_89,N_2964,N_2950);
and UO_90 (O_90,N_2987,N_2996);
nand UO_91 (O_91,N_2999,N_2963);
or UO_92 (O_92,N_2960,N_2967);
or UO_93 (O_93,N_2971,N_2955);
or UO_94 (O_94,N_2967,N_2987);
nor UO_95 (O_95,N_2962,N_2960);
nor UO_96 (O_96,N_2946,N_2955);
and UO_97 (O_97,N_2961,N_2966);
or UO_98 (O_98,N_2943,N_2957);
or UO_99 (O_99,N_2956,N_2957);
and UO_100 (O_100,N_2948,N_2947);
or UO_101 (O_101,N_2958,N_2988);
nand UO_102 (O_102,N_2942,N_2965);
nor UO_103 (O_103,N_2975,N_2970);
or UO_104 (O_104,N_2966,N_2985);
or UO_105 (O_105,N_2985,N_2949);
and UO_106 (O_106,N_2943,N_2963);
or UO_107 (O_107,N_2954,N_2970);
and UO_108 (O_108,N_2970,N_2956);
and UO_109 (O_109,N_2972,N_2941);
or UO_110 (O_110,N_2982,N_2967);
or UO_111 (O_111,N_2953,N_2985);
nor UO_112 (O_112,N_2955,N_2940);
and UO_113 (O_113,N_2985,N_2995);
nor UO_114 (O_114,N_2996,N_2989);
nand UO_115 (O_115,N_2988,N_2997);
nor UO_116 (O_116,N_2955,N_2966);
and UO_117 (O_117,N_2990,N_2948);
nand UO_118 (O_118,N_2954,N_2978);
nand UO_119 (O_119,N_2952,N_2977);
nor UO_120 (O_120,N_2992,N_2999);
and UO_121 (O_121,N_2983,N_2975);
nand UO_122 (O_122,N_2984,N_2988);
or UO_123 (O_123,N_2979,N_2946);
and UO_124 (O_124,N_2960,N_2995);
nand UO_125 (O_125,N_2982,N_2995);
nor UO_126 (O_126,N_2943,N_2988);
and UO_127 (O_127,N_2944,N_2989);
or UO_128 (O_128,N_2978,N_2953);
and UO_129 (O_129,N_2952,N_2945);
nand UO_130 (O_130,N_2958,N_2959);
and UO_131 (O_131,N_2941,N_2951);
nor UO_132 (O_132,N_2940,N_2947);
and UO_133 (O_133,N_2942,N_2982);
and UO_134 (O_134,N_2982,N_2992);
and UO_135 (O_135,N_2956,N_2976);
and UO_136 (O_136,N_2955,N_2984);
nand UO_137 (O_137,N_2988,N_2978);
or UO_138 (O_138,N_2970,N_2966);
nor UO_139 (O_139,N_2963,N_2991);
nand UO_140 (O_140,N_2991,N_2957);
nand UO_141 (O_141,N_2986,N_2973);
and UO_142 (O_142,N_2949,N_2982);
xnor UO_143 (O_143,N_2964,N_2957);
nand UO_144 (O_144,N_2982,N_2962);
or UO_145 (O_145,N_2972,N_2997);
nor UO_146 (O_146,N_2974,N_2966);
or UO_147 (O_147,N_2991,N_2960);
nand UO_148 (O_148,N_2957,N_2966);
or UO_149 (O_149,N_2964,N_2978);
and UO_150 (O_150,N_2995,N_2943);
or UO_151 (O_151,N_2989,N_2975);
or UO_152 (O_152,N_2953,N_2967);
or UO_153 (O_153,N_2946,N_2947);
nand UO_154 (O_154,N_2961,N_2963);
and UO_155 (O_155,N_2964,N_2985);
nor UO_156 (O_156,N_2982,N_2943);
and UO_157 (O_157,N_2962,N_2994);
and UO_158 (O_158,N_2949,N_2948);
or UO_159 (O_159,N_2943,N_2959);
nand UO_160 (O_160,N_2967,N_2988);
nor UO_161 (O_161,N_2982,N_2994);
or UO_162 (O_162,N_2999,N_2962);
and UO_163 (O_163,N_2971,N_2986);
nand UO_164 (O_164,N_2941,N_2974);
xor UO_165 (O_165,N_2966,N_2988);
or UO_166 (O_166,N_2964,N_2962);
nand UO_167 (O_167,N_2987,N_2963);
or UO_168 (O_168,N_2940,N_2998);
and UO_169 (O_169,N_2959,N_2997);
or UO_170 (O_170,N_2956,N_2963);
and UO_171 (O_171,N_2947,N_2984);
and UO_172 (O_172,N_2952,N_2976);
nand UO_173 (O_173,N_2980,N_2956);
nor UO_174 (O_174,N_2981,N_2990);
nand UO_175 (O_175,N_2980,N_2988);
nor UO_176 (O_176,N_2987,N_2981);
nand UO_177 (O_177,N_2946,N_2957);
nor UO_178 (O_178,N_2940,N_2982);
nor UO_179 (O_179,N_2982,N_2959);
nand UO_180 (O_180,N_2985,N_2944);
nor UO_181 (O_181,N_2982,N_2961);
and UO_182 (O_182,N_2997,N_2975);
nand UO_183 (O_183,N_2991,N_2995);
nand UO_184 (O_184,N_2996,N_2941);
and UO_185 (O_185,N_2968,N_2974);
nand UO_186 (O_186,N_2963,N_2946);
or UO_187 (O_187,N_2976,N_2951);
nand UO_188 (O_188,N_2984,N_2975);
nor UO_189 (O_189,N_2942,N_2963);
and UO_190 (O_190,N_2984,N_2967);
nor UO_191 (O_191,N_2950,N_2971);
and UO_192 (O_192,N_2959,N_2999);
nor UO_193 (O_193,N_2978,N_2942);
nor UO_194 (O_194,N_2995,N_2956);
xnor UO_195 (O_195,N_2966,N_2956);
and UO_196 (O_196,N_2982,N_2998);
nand UO_197 (O_197,N_2969,N_2966);
and UO_198 (O_198,N_2942,N_2976);
and UO_199 (O_199,N_2944,N_2964);
xnor UO_200 (O_200,N_2997,N_2977);
nor UO_201 (O_201,N_2940,N_2991);
or UO_202 (O_202,N_2990,N_2949);
nor UO_203 (O_203,N_2947,N_2944);
and UO_204 (O_204,N_2975,N_2947);
or UO_205 (O_205,N_2987,N_2946);
nor UO_206 (O_206,N_2980,N_2940);
and UO_207 (O_207,N_2943,N_2990);
nand UO_208 (O_208,N_2975,N_2955);
xnor UO_209 (O_209,N_2972,N_2963);
nor UO_210 (O_210,N_2997,N_2998);
and UO_211 (O_211,N_2983,N_2971);
nor UO_212 (O_212,N_2986,N_2996);
and UO_213 (O_213,N_2986,N_2987);
nand UO_214 (O_214,N_2965,N_2946);
and UO_215 (O_215,N_2984,N_2972);
xor UO_216 (O_216,N_2991,N_2979);
and UO_217 (O_217,N_2986,N_2977);
nor UO_218 (O_218,N_2994,N_2958);
nand UO_219 (O_219,N_2957,N_2972);
nand UO_220 (O_220,N_2986,N_2981);
and UO_221 (O_221,N_2988,N_2961);
nand UO_222 (O_222,N_2996,N_2959);
and UO_223 (O_223,N_2966,N_2991);
or UO_224 (O_224,N_2984,N_2978);
or UO_225 (O_225,N_2972,N_2967);
and UO_226 (O_226,N_2951,N_2944);
nand UO_227 (O_227,N_2991,N_2973);
nor UO_228 (O_228,N_2942,N_2995);
nor UO_229 (O_229,N_2948,N_2991);
xor UO_230 (O_230,N_2980,N_2975);
nor UO_231 (O_231,N_2944,N_2946);
or UO_232 (O_232,N_2953,N_2949);
and UO_233 (O_233,N_2966,N_2975);
or UO_234 (O_234,N_2999,N_2970);
or UO_235 (O_235,N_2952,N_2971);
or UO_236 (O_236,N_2973,N_2980);
nor UO_237 (O_237,N_2965,N_2949);
or UO_238 (O_238,N_2983,N_2990);
nand UO_239 (O_239,N_2952,N_2998);
or UO_240 (O_240,N_2984,N_2970);
and UO_241 (O_241,N_2944,N_2974);
nor UO_242 (O_242,N_2967,N_2942);
nand UO_243 (O_243,N_2978,N_2992);
nand UO_244 (O_244,N_2979,N_2964);
and UO_245 (O_245,N_2971,N_2976);
or UO_246 (O_246,N_2946,N_2951);
or UO_247 (O_247,N_2977,N_2946);
nor UO_248 (O_248,N_2985,N_2992);
nor UO_249 (O_249,N_2978,N_2973);
nand UO_250 (O_250,N_2950,N_2940);
nor UO_251 (O_251,N_2949,N_2941);
nand UO_252 (O_252,N_2992,N_2991);
nand UO_253 (O_253,N_2956,N_2973);
nor UO_254 (O_254,N_2955,N_2980);
nand UO_255 (O_255,N_2941,N_2990);
or UO_256 (O_256,N_2978,N_2977);
or UO_257 (O_257,N_2991,N_2975);
or UO_258 (O_258,N_2972,N_2992);
nand UO_259 (O_259,N_2954,N_2955);
and UO_260 (O_260,N_2998,N_2994);
or UO_261 (O_261,N_2947,N_2969);
or UO_262 (O_262,N_2947,N_2968);
nor UO_263 (O_263,N_2994,N_2947);
and UO_264 (O_264,N_2999,N_2995);
nand UO_265 (O_265,N_2945,N_2979);
and UO_266 (O_266,N_2945,N_2973);
nor UO_267 (O_267,N_2975,N_2996);
nor UO_268 (O_268,N_2960,N_2953);
and UO_269 (O_269,N_2967,N_2986);
nor UO_270 (O_270,N_2974,N_2973);
nor UO_271 (O_271,N_2989,N_2965);
nor UO_272 (O_272,N_2942,N_2947);
nor UO_273 (O_273,N_2953,N_2951);
nand UO_274 (O_274,N_2992,N_2970);
nor UO_275 (O_275,N_2944,N_2996);
nand UO_276 (O_276,N_2956,N_2943);
nand UO_277 (O_277,N_2943,N_2950);
and UO_278 (O_278,N_2972,N_2947);
and UO_279 (O_279,N_2997,N_2949);
nor UO_280 (O_280,N_2995,N_2996);
nor UO_281 (O_281,N_2990,N_2989);
nand UO_282 (O_282,N_2982,N_2986);
nor UO_283 (O_283,N_2959,N_2961);
nor UO_284 (O_284,N_2940,N_2954);
or UO_285 (O_285,N_2955,N_2982);
nor UO_286 (O_286,N_2950,N_2981);
nand UO_287 (O_287,N_2986,N_2969);
xor UO_288 (O_288,N_2998,N_2957);
nor UO_289 (O_289,N_2998,N_2996);
and UO_290 (O_290,N_2994,N_2963);
nand UO_291 (O_291,N_2979,N_2989);
nor UO_292 (O_292,N_2983,N_2961);
and UO_293 (O_293,N_2964,N_2996);
nand UO_294 (O_294,N_2965,N_2969);
nor UO_295 (O_295,N_2967,N_2981);
nor UO_296 (O_296,N_2978,N_2971);
and UO_297 (O_297,N_2981,N_2999);
nand UO_298 (O_298,N_2972,N_2976);
and UO_299 (O_299,N_2968,N_2992);
and UO_300 (O_300,N_2977,N_2994);
and UO_301 (O_301,N_2987,N_2978);
or UO_302 (O_302,N_2980,N_2964);
nor UO_303 (O_303,N_2962,N_2958);
nor UO_304 (O_304,N_2950,N_2989);
nor UO_305 (O_305,N_2942,N_2960);
and UO_306 (O_306,N_2992,N_2971);
xor UO_307 (O_307,N_2950,N_2942);
nor UO_308 (O_308,N_2961,N_2978);
nand UO_309 (O_309,N_2966,N_2997);
and UO_310 (O_310,N_2997,N_2982);
and UO_311 (O_311,N_2968,N_2945);
and UO_312 (O_312,N_2995,N_2948);
and UO_313 (O_313,N_2943,N_2971);
nand UO_314 (O_314,N_2949,N_2976);
and UO_315 (O_315,N_2973,N_2998);
nor UO_316 (O_316,N_2986,N_2999);
and UO_317 (O_317,N_2959,N_2955);
and UO_318 (O_318,N_2958,N_2949);
xnor UO_319 (O_319,N_2973,N_2946);
nand UO_320 (O_320,N_2980,N_2958);
or UO_321 (O_321,N_2984,N_2954);
nor UO_322 (O_322,N_2953,N_2994);
nor UO_323 (O_323,N_2965,N_2966);
or UO_324 (O_324,N_2993,N_2998);
nand UO_325 (O_325,N_2973,N_2959);
or UO_326 (O_326,N_2951,N_2956);
and UO_327 (O_327,N_2963,N_2981);
nor UO_328 (O_328,N_2975,N_2961);
nand UO_329 (O_329,N_2993,N_2995);
nor UO_330 (O_330,N_2979,N_2981);
nor UO_331 (O_331,N_2954,N_2949);
nand UO_332 (O_332,N_2975,N_2998);
nor UO_333 (O_333,N_2955,N_2995);
nor UO_334 (O_334,N_2992,N_2996);
nand UO_335 (O_335,N_2982,N_2983);
nand UO_336 (O_336,N_2950,N_2969);
or UO_337 (O_337,N_2990,N_2966);
and UO_338 (O_338,N_2994,N_2941);
or UO_339 (O_339,N_2954,N_2974);
nand UO_340 (O_340,N_2996,N_2958);
or UO_341 (O_341,N_2957,N_2963);
or UO_342 (O_342,N_2965,N_2971);
nor UO_343 (O_343,N_2944,N_2980);
nand UO_344 (O_344,N_2988,N_2999);
nand UO_345 (O_345,N_2956,N_2986);
and UO_346 (O_346,N_2952,N_2982);
and UO_347 (O_347,N_2964,N_2970);
and UO_348 (O_348,N_2985,N_2962);
or UO_349 (O_349,N_2980,N_2995);
or UO_350 (O_350,N_2973,N_2951);
or UO_351 (O_351,N_2947,N_2949);
or UO_352 (O_352,N_2978,N_2983);
or UO_353 (O_353,N_2944,N_2977);
or UO_354 (O_354,N_2943,N_2949);
nand UO_355 (O_355,N_2950,N_2956);
nor UO_356 (O_356,N_2954,N_2993);
or UO_357 (O_357,N_2985,N_2987);
nand UO_358 (O_358,N_2940,N_2963);
or UO_359 (O_359,N_2949,N_2942);
or UO_360 (O_360,N_2972,N_2973);
nand UO_361 (O_361,N_2963,N_2952);
and UO_362 (O_362,N_2956,N_2948);
xor UO_363 (O_363,N_2978,N_2968);
or UO_364 (O_364,N_2946,N_2943);
nand UO_365 (O_365,N_2966,N_2948);
nor UO_366 (O_366,N_2985,N_2941);
nand UO_367 (O_367,N_2955,N_2951);
and UO_368 (O_368,N_2940,N_2942);
nor UO_369 (O_369,N_2968,N_2982);
or UO_370 (O_370,N_2940,N_2989);
nor UO_371 (O_371,N_2978,N_2963);
nand UO_372 (O_372,N_2979,N_2940);
nor UO_373 (O_373,N_2949,N_2992);
or UO_374 (O_374,N_2983,N_2997);
nand UO_375 (O_375,N_2976,N_2947);
nor UO_376 (O_376,N_2946,N_2942);
or UO_377 (O_377,N_2980,N_2949);
nand UO_378 (O_378,N_2973,N_2993);
and UO_379 (O_379,N_2980,N_2942);
and UO_380 (O_380,N_2994,N_2955);
nand UO_381 (O_381,N_2949,N_2951);
nand UO_382 (O_382,N_2959,N_2991);
nor UO_383 (O_383,N_2960,N_2978);
nor UO_384 (O_384,N_2993,N_2969);
or UO_385 (O_385,N_2948,N_2953);
nor UO_386 (O_386,N_2991,N_2983);
nor UO_387 (O_387,N_2975,N_2964);
and UO_388 (O_388,N_2945,N_2953);
or UO_389 (O_389,N_2968,N_2961);
and UO_390 (O_390,N_2949,N_2995);
nand UO_391 (O_391,N_2947,N_2958);
or UO_392 (O_392,N_2994,N_2961);
or UO_393 (O_393,N_2940,N_2988);
nor UO_394 (O_394,N_2999,N_2954);
or UO_395 (O_395,N_2989,N_2968);
nand UO_396 (O_396,N_2979,N_2999);
nor UO_397 (O_397,N_2951,N_2943);
or UO_398 (O_398,N_2976,N_2987);
nor UO_399 (O_399,N_2981,N_2989);
or UO_400 (O_400,N_2994,N_2966);
nor UO_401 (O_401,N_2963,N_2984);
and UO_402 (O_402,N_2974,N_2995);
or UO_403 (O_403,N_2947,N_2980);
nor UO_404 (O_404,N_2986,N_2952);
and UO_405 (O_405,N_2979,N_2990);
and UO_406 (O_406,N_2959,N_2945);
nor UO_407 (O_407,N_2940,N_2949);
and UO_408 (O_408,N_2966,N_2992);
or UO_409 (O_409,N_2997,N_2978);
nand UO_410 (O_410,N_2969,N_2943);
nand UO_411 (O_411,N_2945,N_2982);
nand UO_412 (O_412,N_2990,N_2942);
or UO_413 (O_413,N_2948,N_2958);
nor UO_414 (O_414,N_2951,N_2967);
or UO_415 (O_415,N_2952,N_2961);
or UO_416 (O_416,N_2953,N_2974);
nor UO_417 (O_417,N_2941,N_2944);
nand UO_418 (O_418,N_2961,N_2967);
nand UO_419 (O_419,N_2964,N_2948);
or UO_420 (O_420,N_2997,N_2976);
or UO_421 (O_421,N_2979,N_2954);
nand UO_422 (O_422,N_2941,N_2959);
nor UO_423 (O_423,N_2980,N_2972);
nand UO_424 (O_424,N_2978,N_2952);
nand UO_425 (O_425,N_2980,N_2998);
or UO_426 (O_426,N_2982,N_2964);
or UO_427 (O_427,N_2949,N_2960);
nor UO_428 (O_428,N_2953,N_2940);
or UO_429 (O_429,N_2996,N_2962);
and UO_430 (O_430,N_2954,N_2971);
or UO_431 (O_431,N_2993,N_2970);
nand UO_432 (O_432,N_2959,N_2946);
nand UO_433 (O_433,N_2974,N_2989);
and UO_434 (O_434,N_2962,N_2948);
or UO_435 (O_435,N_2954,N_2981);
or UO_436 (O_436,N_2989,N_2977);
nand UO_437 (O_437,N_2967,N_2971);
nand UO_438 (O_438,N_2993,N_2962);
nand UO_439 (O_439,N_2979,N_2978);
nand UO_440 (O_440,N_2967,N_2943);
and UO_441 (O_441,N_2944,N_2953);
xor UO_442 (O_442,N_2980,N_2981);
nor UO_443 (O_443,N_2967,N_2979);
nand UO_444 (O_444,N_2969,N_2984);
nand UO_445 (O_445,N_2944,N_2995);
nand UO_446 (O_446,N_2988,N_2944);
nand UO_447 (O_447,N_2952,N_2947);
nor UO_448 (O_448,N_2990,N_2963);
and UO_449 (O_449,N_2948,N_2989);
nand UO_450 (O_450,N_2980,N_2976);
nand UO_451 (O_451,N_2960,N_2992);
nand UO_452 (O_452,N_2964,N_2940);
nor UO_453 (O_453,N_2988,N_2950);
and UO_454 (O_454,N_2983,N_2994);
nand UO_455 (O_455,N_2944,N_2954);
nand UO_456 (O_456,N_2974,N_2946);
nor UO_457 (O_457,N_2965,N_2959);
or UO_458 (O_458,N_2971,N_2941);
or UO_459 (O_459,N_2981,N_2955);
or UO_460 (O_460,N_2948,N_2982);
and UO_461 (O_461,N_2955,N_2965);
and UO_462 (O_462,N_2999,N_2967);
nor UO_463 (O_463,N_2974,N_2988);
and UO_464 (O_464,N_2971,N_2979);
and UO_465 (O_465,N_2943,N_2989);
nor UO_466 (O_466,N_2958,N_2963);
and UO_467 (O_467,N_2955,N_2972);
nand UO_468 (O_468,N_2973,N_2967);
nand UO_469 (O_469,N_2964,N_2946);
and UO_470 (O_470,N_2945,N_2984);
nand UO_471 (O_471,N_2967,N_2975);
nor UO_472 (O_472,N_2988,N_2947);
nor UO_473 (O_473,N_2970,N_2944);
or UO_474 (O_474,N_2976,N_2977);
or UO_475 (O_475,N_2980,N_2957);
nand UO_476 (O_476,N_2956,N_2978);
and UO_477 (O_477,N_2965,N_2957);
or UO_478 (O_478,N_2967,N_2958);
nor UO_479 (O_479,N_2941,N_2952);
nor UO_480 (O_480,N_2961,N_2955);
and UO_481 (O_481,N_2985,N_2967);
or UO_482 (O_482,N_2965,N_2940);
nand UO_483 (O_483,N_2983,N_2955);
nor UO_484 (O_484,N_2998,N_2944);
xnor UO_485 (O_485,N_2971,N_2951);
nor UO_486 (O_486,N_2975,N_2963);
and UO_487 (O_487,N_2982,N_2984);
xnor UO_488 (O_488,N_2994,N_2954);
and UO_489 (O_489,N_2964,N_2942);
nand UO_490 (O_490,N_2983,N_2980);
nor UO_491 (O_491,N_2973,N_2958);
nor UO_492 (O_492,N_2940,N_2995);
nand UO_493 (O_493,N_2999,N_2997);
nor UO_494 (O_494,N_2940,N_2967);
nor UO_495 (O_495,N_2957,N_2985);
or UO_496 (O_496,N_2955,N_2996);
or UO_497 (O_497,N_2978,N_2972);
or UO_498 (O_498,N_2958,N_2990);
and UO_499 (O_499,N_2961,N_2976);
endmodule