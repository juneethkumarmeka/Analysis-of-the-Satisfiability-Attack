module basic_2000_20000_2500_25_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_84,In_269);
xor U1 (N_1,In_1631,In_107);
or U2 (N_2,In_201,In_652);
or U3 (N_3,In_1518,In_162);
and U4 (N_4,In_987,In_1418);
and U5 (N_5,In_573,In_1360);
nor U6 (N_6,In_1299,In_1571);
and U7 (N_7,In_1099,In_1496);
xnor U8 (N_8,In_861,In_1906);
xnor U9 (N_9,In_1648,In_1313);
and U10 (N_10,In_1672,In_988);
or U11 (N_11,In_180,In_1076);
nor U12 (N_12,In_1815,In_1785);
or U13 (N_13,In_1008,In_57);
nor U14 (N_14,In_590,In_431);
nand U15 (N_15,In_1966,In_1037);
xor U16 (N_16,In_696,In_754);
nand U17 (N_17,In_1370,In_273);
and U18 (N_18,In_1034,In_1124);
nand U19 (N_19,In_1539,In_246);
nand U20 (N_20,In_879,In_902);
xnor U21 (N_21,In_1472,In_1082);
nor U22 (N_22,In_272,In_20);
and U23 (N_23,In_487,In_1187);
xnor U24 (N_24,In_1736,In_1419);
xnor U25 (N_25,In_699,In_1149);
and U26 (N_26,In_302,In_1381);
xor U27 (N_27,In_1288,In_981);
or U28 (N_28,In_460,In_1028);
or U29 (N_29,In_206,In_673);
nand U30 (N_30,In_1139,In_760);
or U31 (N_31,In_1685,In_1737);
xor U32 (N_32,In_1477,In_504);
nand U33 (N_33,In_405,In_1554);
nand U34 (N_34,In_733,In_767);
nor U35 (N_35,In_907,In_1172);
and U36 (N_36,In_948,In_1192);
and U37 (N_37,In_806,In_892);
xnor U38 (N_38,In_1503,In_224);
nor U39 (N_39,In_597,In_1030);
nor U40 (N_40,In_476,In_1461);
and U41 (N_41,In_886,In_1275);
nor U42 (N_42,In_1052,In_1733);
nor U43 (N_43,In_1445,In_922);
nand U44 (N_44,In_689,In_841);
nand U45 (N_45,In_480,In_370);
nor U46 (N_46,In_1473,In_1555);
and U47 (N_47,In_1661,In_303);
xor U48 (N_48,In_1176,In_204);
xor U49 (N_49,In_401,In_581);
or U50 (N_50,In_167,In_1905);
or U51 (N_51,In_184,In_884);
nand U52 (N_52,In_1625,In_1235);
xor U53 (N_53,In_1501,In_1043);
and U54 (N_54,In_1427,In_1975);
or U55 (N_55,In_833,In_1358);
nand U56 (N_56,In_1831,In_444);
and U57 (N_57,In_1420,In_1440);
or U58 (N_58,In_825,In_908);
nand U59 (N_59,In_514,In_1639);
nor U60 (N_60,In_1933,In_662);
and U61 (N_61,In_900,In_441);
or U62 (N_62,In_1526,In_457);
xnor U63 (N_63,In_517,In_1336);
or U64 (N_64,In_554,In_929);
or U65 (N_65,In_1810,In_51);
and U66 (N_66,In_1886,In_904);
or U67 (N_67,In_332,In_1368);
xnor U68 (N_68,In_1927,In_1502);
xnor U69 (N_69,In_678,In_1219);
xor U70 (N_70,In_89,In_1561);
and U71 (N_71,In_1786,In_464);
or U72 (N_72,In_1878,In_589);
nand U73 (N_73,In_1307,In_1829);
or U74 (N_74,In_1085,In_1750);
and U75 (N_75,In_1668,In_1464);
or U76 (N_76,In_599,In_231);
or U77 (N_77,In_940,In_1179);
and U78 (N_78,In_1867,In_1106);
nand U79 (N_79,In_1154,In_1723);
or U80 (N_80,In_1021,In_1449);
and U81 (N_81,In_1882,In_1848);
nor U82 (N_82,In_1215,In_1936);
nor U83 (N_83,In_1399,In_1392);
xnor U84 (N_84,In_782,In_1494);
or U85 (N_85,In_877,In_209);
nor U86 (N_86,In_1673,In_1078);
or U87 (N_87,In_483,In_1650);
and U88 (N_88,In_1731,In_1186);
and U89 (N_89,In_1115,In_372);
nand U90 (N_90,In_1870,In_15);
nor U91 (N_91,In_968,In_1703);
nor U92 (N_92,In_838,In_1682);
xor U93 (N_93,In_214,In_1627);
nand U94 (N_94,In_1892,In_1541);
and U95 (N_95,In_1677,In_351);
nor U96 (N_96,In_394,In_281);
xnor U97 (N_97,In_154,In_113);
xor U98 (N_98,In_1328,In_526);
nand U99 (N_99,In_1603,In_1863);
nor U100 (N_100,In_722,In_1642);
xnor U101 (N_101,In_291,In_1210);
and U102 (N_102,In_208,In_452);
or U103 (N_103,In_921,In_1083);
nand U104 (N_104,In_759,In_1263);
xor U105 (N_105,In_112,In_1132);
nor U106 (N_106,In_1610,In_1220);
nand U107 (N_107,In_449,In_1365);
or U108 (N_108,In_65,In_1908);
nand U109 (N_109,In_789,In_488);
nor U110 (N_110,In_1509,In_426);
nand U111 (N_111,In_1559,In_1155);
nor U112 (N_112,In_1321,In_1894);
nor U113 (N_113,In_1017,In_1634);
and U114 (N_114,In_1080,In_957);
or U115 (N_115,In_682,In_367);
nand U116 (N_116,In_1506,In_713);
and U117 (N_117,In_670,In_679);
xnor U118 (N_118,In_466,In_1758);
xor U119 (N_119,In_1611,In_442);
nor U120 (N_120,In_1129,In_1230);
and U121 (N_121,In_1126,In_758);
or U122 (N_122,In_1734,In_933);
xor U123 (N_123,In_334,In_583);
xor U124 (N_124,In_55,In_410);
nor U125 (N_125,In_1931,In_1589);
nand U126 (N_126,In_298,In_1973);
xnor U127 (N_127,In_508,In_1852);
and U128 (N_128,In_1040,In_999);
nor U129 (N_129,In_0,In_947);
or U130 (N_130,In_572,In_651);
xor U131 (N_131,In_1970,In_627);
xnor U132 (N_132,In_1049,In_1553);
or U133 (N_133,In_1072,In_1983);
and U134 (N_134,In_63,In_558);
or U135 (N_135,In_1264,In_537);
xor U136 (N_136,In_1893,In_1721);
nand U137 (N_137,In_1497,In_425);
nand U138 (N_138,In_501,In_605);
or U139 (N_139,In_1720,In_1962);
nand U140 (N_140,In_730,In_970);
and U141 (N_141,In_1362,In_27);
nand U142 (N_142,In_761,In_1698);
xnor U143 (N_143,In_1849,In_1422);
or U144 (N_144,In_815,In_749);
nand U145 (N_145,In_587,In_230);
xnor U146 (N_146,In_1993,In_380);
and U147 (N_147,In_18,In_1689);
nand U148 (N_148,In_1641,In_23);
nor U149 (N_149,In_1659,In_396);
nand U150 (N_150,In_976,In_1812);
xor U151 (N_151,In_1122,In_1820);
nor U152 (N_152,In_306,In_642);
nand U153 (N_153,In_832,In_1617);
or U154 (N_154,In_1879,In_1880);
nor U155 (N_155,In_915,In_700);
xnor U156 (N_156,In_997,In_1029);
or U157 (N_157,In_984,In_1408);
nand U158 (N_158,In_936,In_980);
xnor U159 (N_159,In_1955,In_862);
nand U160 (N_160,In_1782,In_683);
and U161 (N_161,In_1570,In_482);
or U162 (N_162,In_898,In_1988);
nor U163 (N_163,In_638,In_477);
xor U164 (N_164,In_336,In_608);
nand U165 (N_165,In_93,In_579);
and U166 (N_166,In_637,In_650);
or U167 (N_167,In_829,In_1699);
and U168 (N_168,In_525,In_261);
or U169 (N_169,In_555,In_601);
or U170 (N_170,In_724,In_1252);
nor U171 (N_171,In_916,In_518);
nand U172 (N_172,In_1918,In_366);
or U173 (N_173,In_328,In_1596);
or U174 (N_174,In_1079,In_326);
nand U175 (N_175,In_147,In_169);
and U176 (N_176,In_239,In_1629);
nor U177 (N_177,In_739,In_1926);
and U178 (N_178,In_562,In_316);
or U179 (N_179,In_238,In_1361);
or U180 (N_180,In_669,In_1696);
nand U181 (N_181,In_1505,In_604);
nand U182 (N_182,In_887,In_223);
and U183 (N_183,In_1110,In_1591);
nor U184 (N_184,In_116,In_645);
nand U185 (N_185,In_59,In_165);
xnor U186 (N_186,In_1267,In_1658);
nor U187 (N_187,In_1031,In_543);
nor U188 (N_188,In_1050,In_1015);
xor U189 (N_189,In_1406,In_119);
and U190 (N_190,In_1100,In_436);
or U191 (N_191,In_1854,In_743);
nand U192 (N_192,In_1002,In_568);
nand U193 (N_193,In_354,In_956);
or U194 (N_194,In_1489,In_1171);
nor U195 (N_195,In_1843,In_468);
xnor U196 (N_196,In_1003,In_268);
xnor U197 (N_197,In_1294,In_855);
xor U198 (N_198,In_1792,In_47);
nor U199 (N_199,In_346,In_923);
nor U200 (N_200,In_1719,In_828);
and U201 (N_201,In_1763,In_1910);
nand U202 (N_202,In_456,In_294);
nor U203 (N_203,In_21,In_909);
and U204 (N_204,In_1081,In_1619);
nor U205 (N_205,In_719,In_1088);
nor U206 (N_206,In_1075,In_926);
xnor U207 (N_207,In_1289,In_132);
nor U208 (N_208,In_819,In_250);
or U209 (N_209,In_786,In_614);
or U210 (N_210,In_1766,In_1114);
or U211 (N_211,In_1874,In_959);
nand U212 (N_212,In_1222,In_865);
nand U213 (N_213,In_891,In_1018);
or U214 (N_214,In_378,In_860);
or U215 (N_215,In_402,In_462);
or U216 (N_216,In_1779,In_166);
and U217 (N_217,In_76,In_1920);
xnor U218 (N_218,In_1058,In_271);
and U219 (N_219,In_258,In_1984);
and U220 (N_220,In_1208,In_86);
and U221 (N_221,In_873,In_395);
nand U222 (N_222,In_288,In_955);
nor U223 (N_223,In_1044,In_1);
or U224 (N_224,In_690,In_1396);
nand U225 (N_225,In_50,In_684);
xor U226 (N_226,In_1168,In_1806);
or U227 (N_227,In_379,In_1855);
nand U228 (N_228,In_1701,In_1051);
nor U229 (N_229,In_746,In_1146);
and U230 (N_230,In_1569,In_1976);
nand U231 (N_231,In_327,In_322);
nor U232 (N_232,In_663,In_38);
nand U233 (N_233,In_1654,In_315);
nand U234 (N_234,In_1759,In_227);
xor U235 (N_235,In_523,In_672);
nor U236 (N_236,In_1388,In_485);
and U237 (N_237,In_1287,In_992);
xor U238 (N_238,In_1460,In_878);
nand U239 (N_239,In_561,In_840);
or U240 (N_240,In_971,In_1257);
nor U241 (N_241,In_1304,In_105);
and U242 (N_242,In_1904,In_1487);
nor U243 (N_243,In_1943,In_1097);
or U244 (N_244,In_257,In_1861);
nor U245 (N_245,In_391,In_170);
and U246 (N_246,In_1528,In_1057);
or U247 (N_247,In_609,In_748);
nor U248 (N_248,In_977,In_626);
nand U249 (N_249,In_1451,In_577);
and U250 (N_250,In_1405,In_454);
xnor U251 (N_251,In_567,In_698);
xnor U252 (N_252,In_1985,In_967);
xor U253 (N_253,In_1979,In_793);
or U254 (N_254,In_91,In_376);
or U255 (N_255,In_676,In_1557);
or U256 (N_256,In_805,In_31);
and U257 (N_257,In_1194,In_1046);
xnor U258 (N_258,In_513,In_681);
nor U259 (N_259,In_983,In_1117);
nand U260 (N_260,In_1202,In_199);
and U261 (N_261,In_318,In_1990);
nand U262 (N_262,In_158,In_1315);
nand U263 (N_263,In_437,In_582);
nand U264 (N_264,In_149,In_1919);
xnor U265 (N_265,In_1417,In_499);
xnor U266 (N_266,In_197,In_944);
and U267 (N_267,In_337,In_1369);
nand U268 (N_268,In_19,In_1441);
nand U269 (N_269,In_177,In_1101);
or U270 (N_270,In_1423,In_643);
xnor U271 (N_271,In_446,In_1764);
nor U272 (N_272,In_1375,In_1415);
and U273 (N_273,In_1374,In_393);
nor U274 (N_274,In_1340,In_3);
nor U275 (N_275,In_191,In_1481);
nand U276 (N_276,In_1317,In_808);
or U277 (N_277,In_1318,In_1711);
nand U278 (N_278,In_1019,In_471);
or U279 (N_279,In_1808,In_45);
nor U280 (N_280,In_615,In_930);
and U281 (N_281,In_1712,In_335);
xor U282 (N_282,In_1679,In_1229);
nand U283 (N_283,In_1457,In_1873);
and U284 (N_284,In_675,In_1607);
nand U285 (N_285,In_935,In_1183);
and U286 (N_286,In_1327,In_639);
nand U287 (N_287,In_434,In_1372);
nand U288 (N_288,In_235,In_1322);
or U289 (N_289,In_1236,In_404);
nor U290 (N_290,In_1690,In_795);
or U291 (N_291,In_1425,In_1104);
or U292 (N_292,In_2,In_356);
or U293 (N_293,In_1379,In_686);
and U294 (N_294,In_450,In_510);
nor U295 (N_295,In_1945,In_1671);
nor U296 (N_296,In_1265,In_1549);
xnor U297 (N_297,In_1657,In_1400);
nand U298 (N_298,In_28,In_389);
xnor U299 (N_299,In_1411,In_1134);
xor U300 (N_300,In_1128,In_150);
and U301 (N_301,In_1412,In_1924);
and U302 (N_302,In_1300,In_317);
xnor U303 (N_303,In_1160,In_1092);
xor U304 (N_304,In_259,In_1162);
nand U305 (N_305,In_1453,In_931);
nand U306 (N_306,In_133,In_1952);
nand U307 (N_307,In_1038,In_175);
and U308 (N_308,In_74,In_1256);
or U309 (N_309,In_540,In_1876);
nor U310 (N_310,In_1298,In_509);
or U311 (N_311,In_1530,In_668);
nor U312 (N_312,In_240,In_1306);
nor U313 (N_313,In_479,In_1628);
or U314 (N_314,In_1013,In_274);
nand U315 (N_315,In_155,In_1799);
xnor U316 (N_316,In_804,In_11);
nor U317 (N_317,In_1067,In_818);
or U318 (N_318,In_1705,In_495);
or U319 (N_319,In_622,In_1470);
or U320 (N_320,In_106,In_1475);
xor U321 (N_321,In_1398,In_226);
and U322 (N_322,In_774,In_1995);
or U323 (N_323,In_310,In_1284);
nand U324 (N_324,In_1726,In_1821);
nor U325 (N_325,In_598,In_635);
nand U326 (N_326,In_1663,In_81);
nand U327 (N_327,In_1823,In_842);
or U328 (N_328,In_1311,In_711);
xnor U329 (N_329,In_835,In_1587);
and U330 (N_330,In_1819,In_1259);
and U331 (N_331,In_7,In_1498);
xor U332 (N_332,In_813,In_530);
nor U333 (N_333,In_1430,In_623);
xnor U334 (N_334,In_810,In_1016);
and U335 (N_335,In_996,In_10);
and U336 (N_336,In_435,In_888);
or U337 (N_337,In_1483,In_1063);
nor U338 (N_338,In_674,In_1048);
or U339 (N_339,In_866,In_1191);
nor U340 (N_340,In_422,In_16);
nor U341 (N_341,In_217,In_1546);
and U342 (N_342,In_938,In_459);
or U343 (N_343,In_817,In_1278);
nor U344 (N_344,In_110,In_1747);
and U345 (N_345,In_634,In_1404);
or U346 (N_346,In_1770,In_415);
and U347 (N_347,In_492,In_1363);
nand U348 (N_348,In_807,In_497);
or U349 (N_349,In_411,In_1865);
nand U350 (N_350,In_1950,In_1478);
xor U351 (N_351,In_802,In_831);
nand U352 (N_352,In_1514,In_1238);
nor U353 (N_353,In_1638,In_228);
and U354 (N_354,In_1350,In_176);
nand U355 (N_355,In_1666,In_848);
xnor U356 (N_356,In_1433,In_1681);
nor U357 (N_357,In_1859,In_953);
and U358 (N_358,In_952,In_853);
or U359 (N_359,In_546,In_1651);
xnor U360 (N_360,In_203,In_1573);
and U361 (N_361,In_183,In_764);
or U362 (N_362,In_1776,In_712);
or U363 (N_363,In_498,In_505);
or U364 (N_364,In_1901,In_1353);
xnor U365 (N_365,In_1377,In_1798);
xnor U366 (N_366,In_1572,In_1978);
nand U367 (N_367,In_97,In_991);
nor U368 (N_368,In_1754,In_1643);
and U369 (N_369,In_413,In_120);
and U370 (N_370,In_1324,In_44);
and U371 (N_371,In_77,In_262);
xor U372 (N_372,In_1212,In_1291);
and U373 (N_373,In_1888,In_1847);
or U374 (N_374,In_121,In_277);
nand U375 (N_375,In_507,In_1409);
and U376 (N_376,In_96,In_340);
and U377 (N_377,In_69,In_1772);
xnor U378 (N_378,In_779,In_1467);
nand U379 (N_379,In_1680,In_803);
and U380 (N_380,In_737,In_858);
nor U381 (N_381,In_1319,In_1277);
nand U382 (N_382,In_266,In_29);
nor U383 (N_383,In_32,In_1105);
or U384 (N_384,In_544,In_1954);
and U385 (N_385,In_913,In_899);
or U386 (N_386,In_548,In_1748);
nor U387 (N_387,In_213,In_30);
and U388 (N_388,In_1735,In_1568);
nand U389 (N_389,In_200,In_843);
or U390 (N_390,In_1131,In_429);
nor U391 (N_391,In_1500,In_1609);
and U392 (N_392,In_785,In_1244);
nand U393 (N_393,In_34,In_205);
or U394 (N_394,In_1329,In_1184);
nand U395 (N_395,In_1940,In_1225);
nor U396 (N_396,In_1248,In_1382);
nand U397 (N_397,In_198,In_1153);
nor U398 (N_398,In_986,In_493);
nand U399 (N_399,In_244,In_1717);
xnor U400 (N_400,In_320,In_1009);
xnor U401 (N_401,In_1836,In_1280);
nor U402 (N_402,In_1310,In_1563);
nor U403 (N_403,In_1635,In_1237);
and U404 (N_404,In_1209,In_1567);
xor U405 (N_405,In_633,In_506);
nand U406 (N_406,In_1989,In_1620);
and U407 (N_407,In_1325,In_1722);
or U408 (N_408,In_1035,In_1157);
nor U409 (N_409,In_1652,In_1190);
nand U410 (N_410,In_882,In_1709);
or U411 (N_411,In_1697,In_765);
or U412 (N_412,In_1923,In_1055);
nand U413 (N_413,In_472,In_1783);
nand U414 (N_414,In_1520,In_1728);
nor U415 (N_415,In_1448,In_1270);
nor U416 (N_416,In_219,In_1787);
nand U417 (N_417,In_791,In_657);
or U418 (N_418,In_1337,In_1755);
xor U419 (N_419,In_1507,In_1669);
nor U420 (N_420,In_195,In_1391);
or U421 (N_421,In_1108,In_894);
or U422 (N_422,In_329,In_365);
nor U423 (N_423,In_52,In_151);
nand U424 (N_424,In_1207,In_1303);
nand U425 (N_425,In_1203,In_1144);
xor U426 (N_426,In_1622,In_79);
and U427 (N_427,In_275,In_1626);
nand U428 (N_428,In_1247,In_1140);
nor U429 (N_429,In_741,In_618);
or U430 (N_430,In_1074,In_776);
xor U431 (N_431,In_1316,In_22);
nor U432 (N_432,In_1471,In_144);
xnor U433 (N_433,In_1794,In_1200);
xor U434 (N_434,In_1334,In_1960);
nand U435 (N_435,In_982,In_1997);
nand U436 (N_436,In_179,In_1274);
and U437 (N_437,In_153,In_823);
xor U438 (N_438,In_1584,In_392);
nor U439 (N_439,In_511,In_140);
or U440 (N_440,In_1109,In_243);
or U441 (N_441,In_1196,In_1581);
nor U442 (N_442,In_256,In_849);
and U443 (N_443,In_751,In_461);
xnor U444 (N_444,In_969,In_1949);
nand U445 (N_445,In_344,In_260);
nor U446 (N_446,In_1338,In_1053);
xnor U447 (N_447,In_1512,In_8);
and U448 (N_448,In_649,In_1492);
nand U449 (N_449,In_1687,In_757);
or U450 (N_450,In_560,In_1604);
or U451 (N_451,In_358,In_137);
nand U452 (N_452,In_1402,In_771);
xor U453 (N_453,In_82,In_1414);
and U454 (N_454,In_578,In_216);
nand U455 (N_455,In_1045,In_566);
xor U456 (N_456,In_419,In_338);
xor U457 (N_457,In_1862,In_1476);
xor U458 (N_458,In_347,In_1232);
xnor U459 (N_459,In_591,In_1438);
nand U460 (N_460,In_595,In_1616);
nor U461 (N_461,In_278,In_797);
nand U462 (N_462,In_439,In_896);
nand U463 (N_463,In_1323,In_769);
nand U464 (N_464,In_822,In_178);
nand U465 (N_465,In_1994,In_1371);
and U466 (N_466,In_1814,In_961);
and U467 (N_467,In_1795,In_1761);
nand U468 (N_468,In_128,In_486);
or U469 (N_469,In_58,In_1664);
and U470 (N_470,In_1828,In_94);
nand U471 (N_471,In_362,In_481);
or U472 (N_472,In_289,In_12);
nand U473 (N_473,In_1913,In_1757);
and U474 (N_474,In_1401,In_280);
nand U475 (N_475,In_171,In_1929);
xnor U476 (N_476,In_1486,In_237);
xnor U477 (N_477,In_1729,In_721);
nand U478 (N_478,In_867,In_542);
nand U479 (N_479,In_1637,In_910);
xor U480 (N_480,In_1925,In_1479);
xnor U481 (N_481,In_264,In_734);
nand U482 (N_482,In_845,In_1916);
or U483 (N_483,In_80,In_1020);
nand U484 (N_484,In_1357,In_352);
nor U485 (N_485,In_1521,In_871);
xor U486 (N_486,In_95,In_1773);
and U487 (N_487,In_1613,In_917);
and U488 (N_488,In_432,In_780);
and U489 (N_489,In_893,In_1964);
nor U490 (N_490,In_1877,In_1271);
nor U491 (N_491,In_958,In_1547);
and U492 (N_492,In_1868,In_1592);
or U493 (N_493,In_1218,In_1258);
xnor U494 (N_494,In_345,In_1426);
or U495 (N_495,In_1178,In_1732);
xor U496 (N_496,In_946,In_41);
nor U497 (N_497,In_1822,In_1495);
xnor U498 (N_498,In_569,In_1938);
xnor U499 (N_499,In_667,In_323);
nor U500 (N_500,In_254,In_220);
or U501 (N_501,In_98,In_1504);
nor U502 (N_502,In_1545,In_640);
xor U503 (N_503,In_470,In_1145);
nor U504 (N_504,In_1649,In_341);
and U505 (N_505,In_631,In_1455);
and U506 (N_506,In_368,In_705);
and U507 (N_507,In_1098,In_809);
nor U508 (N_508,In_949,In_736);
xnor U509 (N_509,In_836,In_1911);
and U510 (N_510,In_972,In_1262);
or U511 (N_511,In_1407,In_99);
xnor U512 (N_512,In_37,In_787);
or U513 (N_513,In_697,In_1840);
or U514 (N_514,In_126,In_134);
xnor U515 (N_515,In_753,In_491);
nor U516 (N_516,In_1282,In_1437);
xor U517 (N_517,In_1953,In_636);
or U518 (N_518,In_1068,In_664);
nand U519 (N_519,In_263,In_409);
xor U520 (N_520,In_1713,In_1159);
nand U521 (N_521,In_407,In_906);
nor U522 (N_522,In_556,In_1790);
or U523 (N_523,In_1835,In_54);
nor U524 (N_524,In_360,In_353);
nand U525 (N_525,In_1090,In_596);
nand U526 (N_526,In_475,In_1749);
nor U527 (N_527,In_1197,In_1393);
or U528 (N_528,In_1389,In_1292);
and U529 (N_529,In_40,In_1390);
nand U530 (N_530,In_1667,In_182);
xor U531 (N_531,In_812,In_1536);
xor U532 (N_532,In_1224,In_145);
nor U533 (N_533,In_1562,In_1005);
and U534 (N_534,In_1537,In_557);
and U535 (N_535,In_1683,In_125);
nand U536 (N_536,In_279,In_265);
xor U537 (N_537,In_1421,In_1347);
nand U538 (N_538,In_869,In_222);
and U539 (N_539,In_1775,In_1800);
nand U540 (N_540,In_308,In_387);
nand U541 (N_541,In_1725,In_1102);
and U542 (N_542,In_1832,In_1780);
or U543 (N_543,In_1897,In_1228);
or U544 (N_544,In_1066,In_453);
and U545 (N_545,In_241,In_706);
and U546 (N_546,In_752,In_1198);
and U547 (N_547,In_620,In_883);
and U548 (N_548,In_606,In_1205);
and U549 (N_549,In_1577,In_1845);
and U550 (N_550,In_1181,In_361);
or U551 (N_551,In_1261,In_159);
xor U552 (N_552,In_747,In_1301);
nor U553 (N_553,In_1857,In_720);
xnor U554 (N_554,In_1674,In_100);
nor U555 (N_555,In_603,In_321);
xor U556 (N_556,In_1130,In_123);
and U557 (N_557,In_1891,In_1670);
xnor U558 (N_558,In_1804,In_1269);
or U559 (N_559,In_1718,In_1837);
or U560 (N_560,In_927,In_1781);
and U561 (N_561,In_1791,In_1551);
nand U562 (N_562,In_325,In_1948);
nor U563 (N_563,In_989,In_1590);
xnor U564 (N_564,In_529,In_1033);
xor U565 (N_565,In_1410,In_296);
nand U566 (N_566,In_1550,In_978);
or U567 (N_567,In_654,In_1214);
or U568 (N_568,In_1656,In_1004);
nor U569 (N_569,In_695,In_594);
or U570 (N_570,In_656,In_1818);
or U571 (N_571,In_124,In_522);
xnor U572 (N_572,In_1484,In_1632);
and U573 (N_573,In_881,In_837);
and U574 (N_574,In_1469,In_1450);
nor U575 (N_575,In_192,In_928);
and U576 (N_576,In_1851,In_1351);
nor U577 (N_577,In_1290,In_1151);
or U578 (N_578,In_304,In_414);
and U579 (N_579,In_1895,In_1061);
and U580 (N_580,In_148,In_1166);
nor U581 (N_581,In_1606,In_740);
xor U582 (N_582,In_538,In_872);
xor U583 (N_583,In_727,In_357);
xnor U584 (N_584,In_796,In_5);
or U585 (N_585,In_1268,In_350);
nand U586 (N_586,In_152,In_1939);
xnor U587 (N_587,In_610,In_1169);
nand U588 (N_588,In_1113,In_1026);
and U589 (N_589,In_592,In_541);
xor U590 (N_590,In_945,In_1534);
nor U591 (N_591,In_221,In_1127);
or U592 (N_592,In_1356,In_1435);
and U593 (N_593,In_1000,In_67);
and U594 (N_594,In_202,In_1745);
or U595 (N_595,In_1452,In_1813);
and U596 (N_596,In_381,In_1346);
xnor U597 (N_597,In_1142,In_212);
and U598 (N_598,In_1056,In_1930);
nand U599 (N_599,In_440,In_1706);
nand U600 (N_600,In_247,In_1490);
xor U601 (N_601,In_1951,In_1251);
xnor U602 (N_602,In_616,In_1387);
or U603 (N_603,In_1853,In_355);
nand U604 (N_604,In_1710,In_715);
nor U605 (N_605,In_1802,In_286);
xnor U606 (N_606,In_1182,In_1850);
and U607 (N_607,In_1576,In_1646);
nor U608 (N_608,In_1245,In_966);
or U609 (N_609,In_1618,In_1286);
or U610 (N_610,In_1889,In_1141);
and U611 (N_611,In_1175,In_1330);
and U612 (N_612,In_1746,In_965);
nand U613 (N_613,In_1297,In_469);
or U614 (N_614,In_1624,In_1760);
nor U615 (N_615,In_1480,In_290);
xnor U616 (N_616,In_141,In_912);
and U617 (N_617,In_1386,In_1540);
xnor U618 (N_618,In_1858,In_644);
xnor U619 (N_619,In_1598,In_463);
or U620 (N_620,In_397,In_218);
or U621 (N_621,In_1273,In_1397);
or U622 (N_622,In_73,In_630);
nor U623 (N_623,In_742,In_942);
xor U624 (N_624,In_1091,In_1560);
nand U625 (N_625,In_847,In_1533);
or U626 (N_626,In_1087,In_408);
nor U627 (N_627,In_1675,In_1765);
xor U628 (N_628,In_1739,In_1524);
xnor U629 (N_629,In_718,In_412);
and U630 (N_630,In_1150,In_104);
and U631 (N_631,In_680,In_1295);
or U632 (N_632,In_1376,In_954);
or U633 (N_633,In_755,In_1384);
and U634 (N_634,In_852,In_284);
or U635 (N_635,In_559,In_417);
nor U636 (N_636,In_1972,In_1042);
nor U637 (N_637,In_552,In_1333);
xnor U638 (N_638,In_725,In_270);
xnor U639 (N_639,In_1069,In_1474);
nand U640 (N_640,In_821,In_1707);
xor U641 (N_641,In_1511,In_839);
nand U642 (N_642,In_775,In_918);
or U643 (N_643,In_458,In_1077);
nor U644 (N_644,In_174,In_451);
and U645 (N_645,In_313,In_163);
nand U646 (N_646,In_1914,In_297);
nor U647 (N_647,In_1296,In_1692);
xor U648 (N_648,In_1583,In_1354);
nand U649 (N_649,In_161,In_993);
nor U650 (N_650,In_295,In_824);
nand U651 (N_651,In_939,In_1986);
xor U652 (N_652,In_1702,In_1320);
or U653 (N_653,In_710,In_1665);
xor U654 (N_654,In_1768,In_1001);
nor U655 (N_655,In_1281,In_406);
xnor U656 (N_656,In_1825,In_1769);
nor U657 (N_657,In_248,In_1595);
or U658 (N_658,In_1089,In_1946);
or U659 (N_659,In_1774,In_1204);
xor U660 (N_660,In_1465,In_1633);
nor U661 (N_661,In_88,In_658);
nand U662 (N_662,In_1898,In_1444);
or U663 (N_663,In_1217,In_535);
nand U664 (N_664,In_1283,In_430);
or U665 (N_665,In_607,In_1691);
nand U666 (N_666,In_564,In_1797);
nand U667 (N_667,In_1348,In_704);
nand U668 (N_668,In_1969,In_1971);
nor U669 (N_669,In_516,In_1992);
xor U670 (N_670,In_1246,In_632);
nand U671 (N_671,In_1597,In_1974);
and U672 (N_672,In_1188,In_1645);
xor U673 (N_673,In_1532,In_1743);
nor U674 (N_674,In_1189,In_1996);
or U675 (N_675,In_1064,In_905);
and U676 (N_676,In_136,In_1838);
nor U677 (N_677,In_1956,In_473);
and U678 (N_678,In_1443,In_551);
nor U679 (N_679,In_467,In_403);
or U680 (N_680,In_373,In_484);
nor U681 (N_681,In_1788,In_399);
nand U682 (N_682,In_53,In_314);
xor U683 (N_683,In_1195,In_418);
or U684 (N_684,In_943,In_1522);
nor U685 (N_685,In_1907,In_1094);
nand U686 (N_686,In_1023,In_1999);
or U687 (N_687,In_531,In_1871);
nand U688 (N_688,In_299,In_864);
xnor U689 (N_689,In_312,In_1644);
xnor U690 (N_690,In_1442,In_951);
xor U691 (N_691,In_181,In_1887);
and U692 (N_692,In_528,In_1941);
and U693 (N_693,In_142,In_26);
xnor U694 (N_694,In_1844,In_1279);
nor U695 (N_695,In_1041,In_14);
nor U696 (N_696,In_1890,In_1987);
and U697 (N_697,In_1753,In_1250);
nand U698 (N_698,In_135,In_1957);
xor U699 (N_699,In_1944,In_1883);
or U700 (N_700,In_844,In_1488);
xnor U701 (N_701,In_889,In_641);
nand U702 (N_702,In_1688,In_1856);
and U703 (N_703,In_1588,In_1434);
nand U704 (N_704,In_1579,In_1367);
nand U705 (N_705,In_895,In_427);
xnor U706 (N_706,In_762,In_1364);
or U707 (N_707,In_39,In_790);
and U708 (N_708,In_60,In_1875);
nor U709 (N_709,In_1177,In_1778);
xnor U710 (N_710,In_48,In_820);
nand U711 (N_711,In_994,In_1896);
nor U712 (N_712,In_1615,In_490);
and U713 (N_713,In_792,In_1830);
and U714 (N_714,In_876,In_330);
nor U715 (N_715,In_1803,In_1678);
nor U716 (N_716,In_660,In_611);
nand U717 (N_717,In_735,In_1084);
or U718 (N_718,In_342,In_593);
xor U719 (N_719,In_1226,In_985);
nand U720 (N_720,In_1135,In_108);
and U721 (N_721,In_348,In_157);
and U722 (N_722,In_1921,In_1086);
or U723 (N_723,In_628,In_1714);
nand U724 (N_724,In_1025,In_1185);
or U725 (N_725,In_363,In_859);
and U726 (N_726,In_68,In_196);
nand U727 (N_727,In_694,In_588);
xnor U728 (N_728,In_1807,In_768);
and U729 (N_729,In_445,In_1039);
and U730 (N_730,In_950,In_172);
xor U731 (N_731,In_1343,In_911);
nand U732 (N_732,In_1582,In_1221);
and U733 (N_733,In_1012,In_1014);
nand U734 (N_734,In_708,In_339);
nor U735 (N_735,In_799,In_1594);
and U736 (N_736,In_576,In_1934);
nor U737 (N_737,In_647,In_1585);
xor U738 (N_738,In_1700,In_242);
nor U739 (N_739,In_811,In_1959);
nand U740 (N_740,In_43,In_400);
and U741 (N_741,In_1961,In_61);
and U742 (N_742,In_925,In_1909);
and U743 (N_743,In_309,In_773);
or U744 (N_744,In_1227,In_1133);
nor U745 (N_745,In_990,In_1612);
or U746 (N_746,In_1342,In_1762);
and U747 (N_747,In_580,In_6);
or U748 (N_748,In_1341,In_772);
nor U749 (N_749,In_750,In_1636);
or U750 (N_750,In_665,In_547);
nand U751 (N_751,In_1630,In_1811);
or U752 (N_752,In_1170,In_249);
and U753 (N_753,In_875,In_1793);
nand U754 (N_754,In_267,In_1662);
nor U755 (N_755,In_287,In_550);
or U756 (N_756,In_210,In_1614);
nor U757 (N_757,In_1394,In_186);
xor U758 (N_758,In_1416,In_1513);
nand U759 (N_759,In_1693,In_502);
xnor U760 (N_760,In_1241,In_1535);
nand U761 (N_761,In_1054,In_798);
and U762 (N_762,In_1740,In_960);
or U763 (N_763,In_1805,In_1608);
or U764 (N_764,In_744,In_1789);
nor U765 (N_765,In_655,In_1314);
or U766 (N_766,In_1869,In_35);
or U767 (N_767,In_331,In_1676);
nor U768 (N_768,In_1548,In_1147);
xnor U769 (N_769,In_1148,In_646);
xnor U770 (N_770,In_731,In_1824);
xnor U771 (N_771,In_1120,In_1796);
xor U772 (N_772,In_870,In_1958);
nand U773 (N_773,In_602,In_1073);
nand U774 (N_774,In_276,In_1538);
and U775 (N_775,In_677,In_816);
xnor U776 (N_776,In_1010,In_103);
nand U777 (N_777,In_173,In_1730);
or U778 (N_778,In_364,In_738);
or U779 (N_779,In_1199,In_1095);
or U780 (N_780,In_830,In_1302);
xor U781 (N_781,In_1446,In_500);
nor U782 (N_782,In_1517,In_117);
nor U783 (N_783,In_539,In_1756);
xnor U784 (N_784,In_146,In_1060);
or U785 (N_785,In_283,In_826);
nand U786 (N_786,In_1902,In_1482);
nor U787 (N_787,In_1982,In_1272);
nand U788 (N_788,In_24,In_1600);
nor U789 (N_789,In_532,In_653);
or U790 (N_790,In_193,In_1767);
nand U791 (N_791,In_1254,In_575);
nand U792 (N_792,In_1564,In_856);
xor U793 (N_793,In_1566,In_252);
xor U794 (N_794,In_1355,In_619);
xnor U795 (N_795,In_1738,In_25);
and U796 (N_796,In_1839,In_1704);
and U797 (N_797,In_1965,In_1111);
or U798 (N_798,In_371,In_963);
or U799 (N_799,In_1694,In_1928);
xor U800 (N_800,N_366,N_585);
xor U801 (N_801,In_1593,N_416);
nand U802 (N_802,In_1841,N_690);
xnor U803 (N_803,N_79,In_763);
or U804 (N_804,In_586,In_565);
and U805 (N_805,N_740,N_411);
nand U806 (N_806,N_19,In_1239);
and U807 (N_807,N_685,N_337);
nor U808 (N_808,In_1912,In_1493);
nand U809 (N_809,N_745,In_781);
or U810 (N_810,N_159,N_23);
nor U811 (N_811,In_709,N_28);
nand U812 (N_812,N_322,N_545);
xor U813 (N_813,N_587,In_1531);
or U814 (N_814,In_827,In_374);
or U815 (N_815,N_719,N_129);
or U816 (N_816,N_384,N_221);
and U817 (N_817,In_1036,N_437);
nand U818 (N_818,In_1331,In_512);
or U819 (N_819,N_87,In_1827);
and U820 (N_820,In_1164,In_115);
nor U821 (N_821,N_608,N_458);
or U822 (N_822,In_1981,N_573);
xor U823 (N_823,In_778,N_490);
xor U824 (N_824,In_666,In_1119);
xor U825 (N_825,N_134,N_495);
nand U826 (N_826,N_140,N_654);
and U827 (N_827,N_670,In_998);
and U828 (N_828,N_396,N_408);
or U829 (N_829,N_471,N_743);
nand U830 (N_830,N_478,N_507);
or U831 (N_831,N_709,N_570);
nand U832 (N_832,In_688,N_128);
xnor U833 (N_833,In_1233,N_504);
nor U834 (N_834,N_647,N_401);
xor U835 (N_835,In_1485,N_254);
and U836 (N_836,In_919,N_750);
xnor U837 (N_837,N_89,In_130);
xor U838 (N_838,N_687,In_1431);
and U839 (N_839,N_668,N_363);
nand U840 (N_840,N_292,N_91);
or U841 (N_841,In_1070,N_315);
nand U842 (N_842,N_84,In_448);
xnor U843 (N_843,N_300,N_656);
xnor U844 (N_844,N_432,In_1447);
nor U845 (N_845,N_11,N_447);
nand U846 (N_846,N_323,N_425);
nor U847 (N_847,N_479,In_1826);
nand U848 (N_848,N_238,N_501);
or U849 (N_849,N_207,N_113);
and U850 (N_850,N_358,N_85);
xor U851 (N_851,In_433,N_622);
or U852 (N_852,N_604,In_1640);
xnor U853 (N_853,N_409,N_399);
xnor U854 (N_854,In_1578,In_1686);
nand U855 (N_855,In_1103,In_1942);
and U856 (N_856,N_413,N_591);
nor U857 (N_857,N_46,In_600);
nand U858 (N_858,N_321,In_253);
or U859 (N_859,N_592,In_1180);
nor U860 (N_860,In_1529,In_118);
and U861 (N_861,In_1032,In_421);
nor U862 (N_862,N_593,N_405);
and U863 (N_863,N_97,In_1468);
and U864 (N_864,In_190,N_331);
or U865 (N_865,In_794,N_572);
nand U866 (N_866,N_277,N_695);
nor U867 (N_867,N_686,N_137);
xor U868 (N_868,N_158,In_4);
nor U869 (N_869,N_489,N_174);
and U870 (N_870,In_863,N_496);
nor U871 (N_871,In_1260,N_403);
or U872 (N_872,N_339,In_225);
or U873 (N_873,N_602,N_83);
and U874 (N_874,N_725,In_1107);
or U875 (N_875,N_735,In_1413);
nand U876 (N_876,In_185,N_232);
nand U877 (N_877,N_394,N_285);
xor U878 (N_878,In_1884,In_515);
or U879 (N_879,N_486,N_309);
or U880 (N_880,In_1947,In_1234);
xnor U881 (N_881,N_776,N_688);
nand U882 (N_882,In_1213,In_717);
and U883 (N_883,In_1574,N_184);
nor U884 (N_884,N_148,In_1174);
xor U885 (N_885,In_1027,In_1899);
nor U886 (N_886,N_731,N_203);
xor U887 (N_887,N_280,N_152);
or U888 (N_888,In_1935,N_259);
or U889 (N_889,In_788,N_256);
xnor U890 (N_890,N_683,In_1359);
and U891 (N_891,N_206,N_787);
and U892 (N_892,N_192,N_550);
or U893 (N_893,N_705,N_90);
nor U894 (N_894,In_390,N_646);
or U895 (N_895,N_75,In_874);
nand U896 (N_896,N_373,N_382);
or U897 (N_897,In_1047,N_156);
or U898 (N_898,N_177,N_455);
and U899 (N_899,N_675,N_620);
and U900 (N_900,N_596,N_70);
nor U901 (N_901,In_834,N_420);
nor U902 (N_902,N_442,In_1096);
nand U903 (N_903,In_1708,In_685);
nor U904 (N_904,In_1385,N_308);
nor U905 (N_905,N_389,N_214);
xnor U906 (N_906,N_338,N_393);
xor U907 (N_907,In_229,N_278);
nor U908 (N_908,In_974,In_520);
or U909 (N_909,N_475,N_674);
nand U910 (N_910,N_553,In_17);
nor U911 (N_911,N_758,In_533);
or U912 (N_912,N_552,N_22);
and U913 (N_913,In_293,In_423);
nand U914 (N_914,N_194,N_726);
or U915 (N_915,In_621,N_288);
and U916 (N_916,In_102,In_549);
xnor U917 (N_917,In_1163,N_730);
nor U918 (N_918,N_357,N_736);
nand U919 (N_919,N_387,N_370);
nor U920 (N_920,In_9,N_115);
nand U921 (N_921,N_763,N_329);
or U922 (N_922,In_1917,N_345);
nor U923 (N_923,N_698,In_1599);
nor U924 (N_924,N_768,N_204);
xor U925 (N_925,N_202,In_1022);
or U926 (N_926,In_885,N_76);
nor U927 (N_927,N_136,N_333);
xnor U928 (N_928,N_746,N_0);
nand U929 (N_929,N_293,N_580);
nand U930 (N_930,N_542,N_630);
or U931 (N_931,In_745,N_556);
nor U932 (N_932,N_616,N_583);
nor U933 (N_933,In_1380,In_245);
nand U934 (N_934,N_120,N_609);
xor U935 (N_935,N_723,In_1173);
and U936 (N_936,In_1165,N_699);
and U937 (N_937,N_727,N_142);
and U938 (N_938,In_1963,N_594);
xnor U939 (N_939,N_778,N_473);
and U940 (N_940,N_679,N_410);
or U941 (N_941,N_124,N_186);
xnor U942 (N_942,N_93,N_498);
or U943 (N_943,In_846,N_151);
and U944 (N_944,In_438,N_146);
xor U945 (N_945,N_60,N_340);
and U946 (N_946,N_100,N_689);
nor U947 (N_947,In_64,In_1695);
and U948 (N_948,In_1206,In_1454);
and U949 (N_949,N_676,In_903);
xnor U950 (N_950,In_311,N_208);
nand U951 (N_951,N_633,N_273);
nor U952 (N_952,In_570,N_290);
nor U953 (N_953,N_230,N_189);
or U954 (N_954,N_527,N_771);
nand U955 (N_955,N_62,N_381);
and U956 (N_956,In_1741,In_398);
or U957 (N_957,In_1742,N_379);
nand U958 (N_958,In_1326,N_492);
nand U959 (N_959,In_377,In_671);
nor U960 (N_960,In_131,In_1866);
xnor U961 (N_961,N_515,N_354);
and U962 (N_962,N_258,N_95);
or U963 (N_963,N_536,In_800);
nand U964 (N_964,N_66,In_897);
nor U965 (N_965,N_77,In_1922);
or U966 (N_966,N_514,N_547);
nor U967 (N_967,N_505,N_421);
nor U968 (N_968,N_170,N_781);
nor U969 (N_969,In_1161,In_251);
nand U970 (N_970,N_611,N_748);
nand U971 (N_971,N_235,In_1403);
nor U972 (N_972,N_737,N_450);
and U973 (N_973,In_1112,N_794);
xnor U974 (N_974,N_243,N_69);
xor U975 (N_975,N_786,In_1801);
xor U976 (N_976,In_92,In_857);
xnor U977 (N_977,In_307,N_320);
nand U978 (N_978,In_301,N_121);
and U979 (N_979,N_739,N_37);
nand U980 (N_980,N_301,N_313);
and U981 (N_981,In_1915,N_601);
nand U982 (N_982,In_1436,N_287);
and U983 (N_983,N_215,N_352);
and U984 (N_984,N_390,In_1784);
and U985 (N_985,N_225,N_548);
nor U986 (N_986,N_239,In_1980);
xnor U987 (N_987,N_296,N_334);
nor U988 (N_988,In_189,N_708);
and U989 (N_989,N_306,In_707);
or U990 (N_990,In_1223,N_67);
or U991 (N_991,N_532,N_132);
nor U992 (N_992,N_380,N_231);
or U993 (N_993,N_759,N_664);
or U994 (N_994,N_294,N_481);
nand U995 (N_995,In_1580,In_1366);
xnor U996 (N_996,N_133,In_70);
nor U997 (N_997,N_700,N_383);
nor U998 (N_998,In_87,N_348);
or U999 (N_999,In_1308,In_56);
nor U1000 (N_1000,N_123,In_1977);
and U1001 (N_1001,N_638,In_1872);
nand U1002 (N_1002,N_782,In_1152);
xor U1003 (N_1003,N_247,N_168);
xor U1004 (N_1004,N_512,N_251);
xnor U1005 (N_1005,N_51,N_419);
nand U1006 (N_1006,N_291,In_1515);
nor U1007 (N_1007,N_377,N_35);
nand U1008 (N_1008,N_788,In_574);
xor U1009 (N_1009,N_216,In_1459);
and U1010 (N_1010,In_1349,N_402);
nor U1011 (N_1011,N_449,N_607);
nand U1012 (N_1012,N_311,In_1352);
nor U1013 (N_1013,N_369,In_1138);
and U1014 (N_1014,N_98,In_305);
and U1015 (N_1015,N_427,In_85);
or U1016 (N_1016,N_744,N_529);
nor U1017 (N_1017,N_717,N_631);
nand U1018 (N_1018,In_1249,N_330);
nand U1019 (N_1019,N_53,In_1834);
xor U1020 (N_1020,N_164,N_653);
xnor U1021 (N_1021,N_167,In_1167);
and U1022 (N_1022,N_663,In_1062);
or U1023 (N_1023,N_58,In_1817);
and U1024 (N_1024,N_274,N_147);
nor U1025 (N_1025,N_246,N_702);
or U1026 (N_1026,N_353,N_173);
xnor U1027 (N_1027,In_1253,N_196);
or U1028 (N_1028,N_165,In_78);
and U1029 (N_1029,N_252,N_680);
nor U1030 (N_1030,N_779,N_494);
nand U1031 (N_1031,N_649,In_1285);
nand U1032 (N_1032,In_1552,N_145);
xor U1033 (N_1033,N_328,N_351);
nor U1034 (N_1034,N_734,In_194);
nand U1035 (N_1035,In_1833,In_207);
xnor U1036 (N_1036,In_1276,In_489);
nor U1037 (N_1037,N_162,N_777);
nand U1038 (N_1038,N_544,N_503);
xor U1039 (N_1039,N_307,N_343);
and U1040 (N_1040,N_344,In_519);
and U1041 (N_1041,N_29,N_88);
nor U1042 (N_1042,N_710,N_102);
or U1043 (N_1043,N_452,N_444);
and U1044 (N_1044,N_283,N_71);
xor U1045 (N_1045,In_850,In_766);
nor U1046 (N_1046,In_612,N_635);
and U1047 (N_1047,In_1543,N_562);
or U1048 (N_1048,N_523,In_1373);
xor U1049 (N_1049,N_644,N_520);
nand U1050 (N_1050,N_440,In_1216);
nor U1051 (N_1051,N_227,In_934);
nand U1052 (N_1052,In_1462,N_508);
xor U1053 (N_1053,N_559,N_86);
xor U1054 (N_1054,In_880,In_122);
nor U1055 (N_1055,N_461,In_164);
or U1056 (N_1056,N_176,In_1466);
nor U1057 (N_1057,N_546,N_267);
or U1058 (N_1058,N_623,N_433);
and U1059 (N_1059,N_448,N_80);
or U1060 (N_1060,N_613,N_24);
and U1061 (N_1061,N_456,N_561);
nand U1062 (N_1062,N_472,N_528);
nand U1063 (N_1063,N_74,In_584);
xor U1064 (N_1064,In_1932,N_226);
nand U1065 (N_1065,N_697,In_962);
or U1066 (N_1066,In_1684,N_463);
nor U1067 (N_1067,N_753,N_640);
and U1068 (N_1068,In_215,N_693);
nand U1069 (N_1069,In_1240,N_733);
xnor U1070 (N_1070,In_188,N_9);
xnor U1071 (N_1071,N_398,N_648);
nand U1072 (N_1072,N_219,N_347);
or U1073 (N_1073,N_141,N_213);
nor U1074 (N_1074,N_36,N_360);
or U1075 (N_1075,N_42,N_412);
nor U1076 (N_1076,N_538,N_241);
nand U1077 (N_1077,In_924,N_289);
or U1078 (N_1078,In_1065,N_434);
and U1079 (N_1079,In_1523,N_385);
nor U1080 (N_1080,N_276,N_109);
xnor U1081 (N_1081,N_754,N_634);
and U1082 (N_1082,In_1998,N_193);
nor U1083 (N_1083,In_233,In_416);
or U1084 (N_1084,N_435,In_211);
nor U1085 (N_1085,N_732,N_324);
and U1086 (N_1086,N_262,In_692);
nor U1087 (N_1087,N_784,N_598);
nand U1088 (N_1088,In_1305,N_138);
or U1089 (N_1089,N_169,N_582);
or U1090 (N_1090,N_480,In_494);
and U1091 (N_1091,N_107,N_564);
xor U1092 (N_1092,N_453,N_792);
nor U1093 (N_1093,N_549,In_420);
xnor U1094 (N_1094,In_1093,In_127);
nor U1095 (N_1095,N_560,N_56);
xnor U1096 (N_1096,In_1991,N_302);
or U1097 (N_1097,N_588,N_579);
nand U1098 (N_1098,In_1724,N_367);
xnor U1099 (N_1099,N_755,N_483);
nand U1100 (N_1100,N_57,In_1508);
nor U1101 (N_1101,N_765,N_704);
nand U1102 (N_1102,In_1335,N_438);
nand U1103 (N_1103,In_1575,N_395);
nand U1104 (N_1104,N_793,In_1527);
xnor U1105 (N_1105,N_658,In_973);
xnor U1106 (N_1106,N_565,N_125);
xor U1107 (N_1107,N_45,N_454);
or U1108 (N_1108,N_41,N_797);
nor U1109 (N_1109,In_1309,N_639);
or U1110 (N_1110,In_1885,In_1395);
nand U1111 (N_1111,In_1525,N_185);
nor U1112 (N_1112,In_319,N_482);
xor U1113 (N_1113,N_775,N_691);
and U1114 (N_1114,N_707,N_355);
nor U1115 (N_1115,N_242,N_332);
nor U1116 (N_1116,N_197,N_183);
nor U1117 (N_1117,N_789,N_780);
xnor U1118 (N_1118,N_43,N_400);
or U1119 (N_1119,N_163,N_678);
xnor U1120 (N_1120,In_1156,N_105);
nand U1121 (N_1121,N_44,In_777);
or U1122 (N_1122,N_672,N_364);
nor U1123 (N_1123,N_667,In_143);
or U1124 (N_1124,In_723,N_397);
xor U1125 (N_1125,In_428,N_566);
xor U1126 (N_1126,N_116,In_1653);
xnor U1127 (N_1127,N_378,N_677);
or U1128 (N_1128,In_1344,N_82);
or U1129 (N_1129,N_191,N_742);
xor U1130 (N_1130,N_713,In_1655);
and U1131 (N_1131,In_343,N_533);
and U1132 (N_1132,N_513,N_669);
nor U1133 (N_1133,In_138,N_228);
nand U1134 (N_1134,N_210,In_1011);
or U1135 (N_1135,N_711,N_275);
or U1136 (N_1136,N_144,In_1499);
nand U1137 (N_1137,N_299,N_5);
or U1138 (N_1138,N_567,N_127);
and U1139 (N_1139,N_143,In_937);
nand U1140 (N_1140,N_724,In_384);
nand U1141 (N_1141,In_324,In_465);
xnor U1142 (N_1142,N_729,In_385);
xor U1143 (N_1143,N_135,In_1339);
xor U1144 (N_1144,N_773,N_554);
nand U1145 (N_1145,In_349,N_391);
or U1146 (N_1146,N_539,N_626);
xor U1147 (N_1147,In_1864,N_614);
or U1148 (N_1148,N_209,N_618);
and U1149 (N_1149,N_359,N_8);
nand U1150 (N_1150,N_428,N_459);
xor U1151 (N_1151,N_50,N_112);
nor U1152 (N_1152,N_131,In_1900);
nor U1153 (N_1153,In_300,N_571);
nand U1154 (N_1154,N_465,N_751);
or U1155 (N_1155,In_1201,N_575);
nor U1156 (N_1156,N_154,N_468);
nor U1157 (N_1157,In_701,In_1744);
nand U1158 (N_1158,N_372,N_27);
or U1159 (N_1159,In_1211,In_139);
and U1160 (N_1160,N_237,In_729);
and U1161 (N_1161,N_52,N_619);
nand U1162 (N_1162,In_1006,N_257);
and U1163 (N_1163,N_303,N_718);
or U1164 (N_1164,N_682,N_263);
xnor U1165 (N_1165,In_571,N_470);
and U1166 (N_1166,N_64,In_1383);
xor U1167 (N_1167,N_493,N_101);
nand U1168 (N_1168,N_319,N_233);
nor U1169 (N_1169,N_282,N_474);
and U1170 (N_1170,In_1231,N_198);
nand U1171 (N_1171,In_42,N_261);
xnor U1172 (N_1172,In_1556,N_476);
or U1173 (N_1173,N_108,In_62);
xor U1174 (N_1174,N_236,N_477);
nand U1175 (N_1175,In_659,N_201);
nor U1176 (N_1176,In_1491,N_31);
nor U1177 (N_1177,N_284,N_49);
xnor U1178 (N_1178,N_783,In_1332);
or U1179 (N_1179,N_388,N_597);
and U1180 (N_1180,N_599,N_55);
nand U1181 (N_1181,N_222,In_625);
or U1182 (N_1182,In_1429,N_255);
nor U1183 (N_1183,In_1586,N_268);
nor U1184 (N_1184,N_253,In_1312);
nand U1185 (N_1185,N_568,In_1439);
nand U1186 (N_1186,N_531,N_484);
and U1187 (N_1187,In_1752,In_375);
nand U1188 (N_1188,In_629,In_424);
or U1189 (N_1189,In_496,In_1118);
xor U1190 (N_1190,N_424,In_521);
or U1191 (N_1191,In_168,N_641);
xor U1192 (N_1192,N_92,In_1660);
nand U1193 (N_1193,In_1510,In_545);
nand U1194 (N_1194,In_1123,N_770);
nand U1195 (N_1195,N_327,N_712);
or U1196 (N_1196,N_722,In_1266);
nand U1197 (N_1197,N_103,N_466);
nor U1198 (N_1198,In_1621,N_166);
nor U1199 (N_1199,In_1903,N_799);
or U1200 (N_1200,In_1458,N_318);
nor U1201 (N_1201,N_681,In_726);
xnor U1202 (N_1202,N_200,In_1243);
and U1203 (N_1203,In_648,N_32);
xor U1204 (N_1204,N_63,N_636);
xor U1205 (N_1205,N_118,N_223);
and U1206 (N_1206,In_359,N_491);
nor U1207 (N_1207,N_684,N_487);
and U1208 (N_1208,N_335,N_48);
or U1209 (N_1209,In_383,In_1601);
and U1210 (N_1210,N_160,N_637);
nand U1211 (N_1211,N_417,N_171);
nand U1212 (N_1212,In_1816,In_1623);
xor U1213 (N_1213,N_392,N_502);
nand U1214 (N_1214,N_40,N_756);
nor U1215 (N_1215,N_747,N_12);
xor U1216 (N_1216,In_702,N_436);
nand U1217 (N_1217,N_589,N_603);
xor U1218 (N_1218,N_617,N_407);
xnor U1219 (N_1219,N_346,N_790);
xor U1220 (N_1220,N_281,N_673);
nand U1221 (N_1221,In_585,In_868);
or U1222 (N_1222,N_126,N_488);
and U1223 (N_1223,N_81,N_798);
nand U1224 (N_1224,N_205,N_362);
or U1225 (N_1225,N_659,N_518);
nand U1226 (N_1226,In_1542,In_292);
and U1227 (N_1227,N_180,In_72);
nor U1228 (N_1228,N_714,In_388);
xor U1229 (N_1229,N_374,N_386);
nand U1230 (N_1230,N_612,In_784);
nand U1231 (N_1231,In_975,N_16);
xnor U1232 (N_1232,In_1809,In_1716);
nand U1233 (N_1233,N_314,N_161);
or U1234 (N_1234,N_13,In_770);
and U1235 (N_1235,N_506,N_497);
or U1236 (N_1236,N_728,N_431);
nand U1237 (N_1237,In_617,N_272);
or U1238 (N_1238,N_757,In_691);
and U1239 (N_1239,In_563,N_250);
and U1240 (N_1240,N_578,N_375);
xnor U1241 (N_1241,In_932,In_109);
and U1242 (N_1242,In_455,N_600);
nor U1243 (N_1243,N_661,N_65);
nor U1244 (N_1244,N_172,In_1059);
nand U1245 (N_1245,N_509,In_1602);
and U1246 (N_1246,N_738,N_312);
or U1247 (N_1247,N_365,N_762);
nand U1248 (N_1248,N_749,In_851);
and U1249 (N_1249,In_703,N_422);
nand U1250 (N_1250,In_624,In_979);
and U1251 (N_1251,N_694,N_2);
and U1252 (N_1252,N_245,In_1842);
nor U1253 (N_1253,In_1715,N_220);
or U1254 (N_1254,N_149,N_439);
and U1255 (N_1255,N_766,N_629);
and U1256 (N_1256,N_218,N_155);
xor U1257 (N_1257,In_1137,N_537);
nand U1258 (N_1258,N_652,N_117);
and U1259 (N_1259,N_264,N_720);
or U1260 (N_1260,N_760,N_628);
or U1261 (N_1261,N_581,In_474);
xnor U1262 (N_1262,N_651,N_34);
and U1263 (N_1263,N_150,In_524);
nand U1264 (N_1264,N_99,N_540);
or U1265 (N_1265,N_541,In_83);
and U1266 (N_1266,N_761,In_1158);
xor U1267 (N_1267,N_305,In_814);
or U1268 (N_1268,N_666,N_650);
nor U1269 (N_1269,In_1751,N_73);
or U1270 (N_1270,In_553,N_18);
nand U1271 (N_1271,N_110,N_376);
nor U1272 (N_1272,N_662,N_310);
or U1273 (N_1273,N_558,In_114);
and U1274 (N_1274,N_316,In_728);
and U1275 (N_1275,In_236,In_1544);
nor U1276 (N_1276,N_271,N_469);
xor U1277 (N_1277,N_229,N_460);
or U1278 (N_1278,N_21,In_90);
xnor U1279 (N_1279,N_187,N_785);
nor U1280 (N_1280,In_1242,In_478);
and U1281 (N_1281,N_551,In_920);
and U1282 (N_1282,N_632,N_467);
xnor U1283 (N_1283,N_6,N_10);
nor U1284 (N_1284,N_178,N_543);
and U1285 (N_1285,N_286,N_769);
xor U1286 (N_1286,N_15,N_706);
and U1287 (N_1287,N_269,N_563);
nor U1288 (N_1288,N_610,N_175);
or U1289 (N_1289,N_426,N_72);
nand U1290 (N_1290,N_721,In_1125);
nand U1291 (N_1291,N_199,In_443);
nor U1292 (N_1292,N_665,In_33);
xnor U1293 (N_1293,N_181,N_244);
or U1294 (N_1294,N_249,In_1846);
xnor U1295 (N_1295,N_68,In_527);
nor U1296 (N_1296,N_26,N_188);
nor U1297 (N_1297,N_304,N_645);
nand U1298 (N_1298,N_139,N_430);
or U1299 (N_1299,N_624,N_61);
and U1300 (N_1300,In_255,In_1605);
nand U1301 (N_1301,In_1424,N_371);
and U1302 (N_1302,In_716,N_234);
nand U1303 (N_1303,In_1378,In_187);
or U1304 (N_1304,N_764,In_71);
and U1305 (N_1305,N_510,N_157);
nand U1306 (N_1306,N_96,N_605);
xor U1307 (N_1307,In_1727,In_232);
and U1308 (N_1308,N_535,N_423);
xor U1309 (N_1309,N_522,N_445);
and U1310 (N_1310,In_156,N_240);
and U1311 (N_1311,N_534,In_661);
and U1312 (N_1312,N_574,In_66);
xnor U1313 (N_1313,In_1516,N_701);
nand U1314 (N_1314,In_1255,N_104);
xor U1315 (N_1315,In_447,In_1293);
nand U1316 (N_1316,In_13,In_1558);
xor U1317 (N_1317,N_295,N_429);
or U1318 (N_1318,In_46,N_265);
or U1319 (N_1319,N_153,In_1860);
nor U1320 (N_1320,N_182,N_555);
and U1321 (N_1321,N_270,N_195);
and U1322 (N_1322,N_606,In_783);
or U1323 (N_1323,In_382,In_282);
nand U1324 (N_1324,N_341,In_534);
nand U1325 (N_1325,In_503,In_1071);
nand U1326 (N_1326,N_526,N_342);
nand U1327 (N_1327,In_333,N_441);
xor U1328 (N_1328,N_418,In_49);
or U1329 (N_1329,In_1116,N_586);
or U1330 (N_1330,N_767,In_1428);
nand U1331 (N_1331,N_111,N_54);
nor U1332 (N_1332,In_995,N_530);
and U1333 (N_1333,N_464,N_569);
xor U1334 (N_1334,N_356,N_130);
xor U1335 (N_1335,N_516,N_317);
nand U1336 (N_1336,N_615,N_217);
nor U1337 (N_1337,In_129,N_190);
nor U1338 (N_1338,N_703,In_1456);
and U1339 (N_1339,In_854,N_326);
nand U1340 (N_1340,In_160,In_1967);
nor U1341 (N_1341,In_914,N_298);
nand U1342 (N_1342,N_457,N_774);
and U1343 (N_1343,N_715,N_25);
and U1344 (N_1344,In_801,N_38);
and U1345 (N_1345,In_369,N_655);
xnor U1346 (N_1346,In_1777,N_224);
xnor U1347 (N_1347,N_78,In_714);
nand U1348 (N_1348,N_59,N_795);
xnor U1349 (N_1349,N_349,In_1771);
nor U1350 (N_1350,In_613,N_521);
or U1351 (N_1351,N_47,In_1432);
and U1352 (N_1352,N_297,In_75);
or U1353 (N_1353,In_536,In_693);
nor U1354 (N_1354,N_642,In_1143);
or U1355 (N_1355,N_772,N_595);
xnor U1356 (N_1356,N_752,N_94);
nand U1357 (N_1357,In_1345,N_696);
and U1358 (N_1358,N_119,N_499);
xnor U1359 (N_1359,In_285,N_643);
xnor U1360 (N_1360,N_660,N_657);
nand U1361 (N_1361,N_500,In_1647);
or U1362 (N_1362,N_350,In_964);
nor U1363 (N_1363,N_627,N_406);
nor U1364 (N_1364,N_796,In_1968);
or U1365 (N_1365,In_1193,N_7);
or U1366 (N_1366,N_114,N_524);
and U1367 (N_1367,N_122,N_741);
and U1368 (N_1368,In_756,N_557);
or U1369 (N_1369,N_20,N_33);
nor U1370 (N_1370,N_625,N_1);
nand U1371 (N_1371,N_404,N_30);
and U1372 (N_1372,N_621,N_576);
nand U1373 (N_1373,N_14,N_511);
nand U1374 (N_1374,In_36,N_336);
and U1375 (N_1375,N_451,N_462);
xnor U1376 (N_1376,N_446,N_179);
and U1377 (N_1377,N_17,N_260);
nor U1378 (N_1378,N_39,In_1937);
xnor U1379 (N_1379,N_692,N_361);
and U1380 (N_1380,In_687,N_4);
or U1381 (N_1381,In_1519,In_890);
xnor U1382 (N_1382,In_1463,N_212);
nand U1383 (N_1383,In_234,N_368);
nor U1384 (N_1384,In_111,In_1024);
nor U1385 (N_1385,N_791,N_525);
xor U1386 (N_1386,In_1136,N_266);
nor U1387 (N_1387,N_485,N_443);
xor U1388 (N_1388,In_901,N_590);
nand U1389 (N_1389,In_941,In_1881);
xnor U1390 (N_1390,N_517,N_325);
nor U1391 (N_1391,N_414,In_1121);
xnor U1392 (N_1392,In_101,N_279);
nand U1393 (N_1393,N_519,N_211);
nand U1394 (N_1394,N_577,N_671);
or U1395 (N_1395,In_1007,N_248);
xnor U1396 (N_1396,N_716,N_106);
nand U1397 (N_1397,N_584,N_3);
nor U1398 (N_1398,N_415,In_1565);
xor U1399 (N_1399,In_386,In_732);
xor U1400 (N_1400,N_249,N_633);
nor U1401 (N_1401,N_4,N_576);
and U1402 (N_1402,N_290,N_616);
or U1403 (N_1403,In_75,In_1519);
nand U1404 (N_1404,In_46,N_247);
nand U1405 (N_1405,In_494,N_573);
or U1406 (N_1406,N_769,In_1339);
nand U1407 (N_1407,In_1827,N_454);
xnor U1408 (N_1408,N_455,N_105);
xor U1409 (N_1409,N_218,In_382);
nor U1410 (N_1410,In_1742,In_571);
nor U1411 (N_1411,N_322,N_307);
nand U1412 (N_1412,In_1395,N_337);
or U1413 (N_1413,N_158,In_443);
and U1414 (N_1414,In_390,N_215);
nor U1415 (N_1415,In_1801,In_1937);
nor U1416 (N_1416,N_566,In_661);
nor U1417 (N_1417,N_243,N_54);
or U1418 (N_1418,In_1152,In_1161);
nor U1419 (N_1419,N_427,N_253);
or U1420 (N_1420,In_1947,In_160);
nand U1421 (N_1421,N_500,N_612);
and U1422 (N_1422,In_574,In_49);
nand U1423 (N_1423,N_539,N_271);
nand U1424 (N_1424,In_1022,In_1527);
or U1425 (N_1425,In_709,In_1771);
and U1426 (N_1426,N_635,In_382);
nand U1427 (N_1427,N_606,N_123);
or U1428 (N_1428,N_529,In_1991);
and U1429 (N_1429,N_26,N_368);
nand U1430 (N_1430,N_430,N_648);
nor U1431 (N_1431,In_1165,In_1686);
or U1432 (N_1432,N_337,In_160);
nor U1433 (N_1433,In_1432,N_27);
xor U1434 (N_1434,N_543,N_348);
or U1435 (N_1435,N_198,In_1846);
nand U1436 (N_1436,N_180,N_582);
nor U1437 (N_1437,In_1578,N_431);
and U1438 (N_1438,N_353,N_658);
nor U1439 (N_1439,N_384,N_156);
nor U1440 (N_1440,N_562,N_647);
and U1441 (N_1441,N_726,In_687);
and U1442 (N_1442,In_465,N_91);
or U1443 (N_1443,In_553,In_138);
nor U1444 (N_1444,N_341,N_632);
nor U1445 (N_1445,N_629,In_143);
and U1446 (N_1446,N_430,N_350);
nand U1447 (N_1447,In_234,N_301);
or U1448 (N_1448,N_757,N_621);
nor U1449 (N_1449,In_1468,N_108);
xnor U1450 (N_1450,N_231,In_343);
or U1451 (N_1451,N_398,In_292);
or U1452 (N_1452,In_863,N_751);
and U1453 (N_1453,N_434,N_680);
and U1454 (N_1454,N_461,N_37);
xor U1455 (N_1455,N_319,N_560);
xor U1456 (N_1456,In_1708,N_659);
xor U1457 (N_1457,N_80,N_686);
xor U1458 (N_1458,N_617,In_111);
xor U1459 (N_1459,In_1771,In_1119);
nand U1460 (N_1460,N_482,N_44);
xor U1461 (N_1461,N_707,N_157);
or U1462 (N_1462,N_105,N_614);
nor U1463 (N_1463,In_229,In_1424);
and U1464 (N_1464,N_510,In_1211);
nand U1465 (N_1465,N_80,N_350);
nand U1466 (N_1466,N_791,N_312);
xor U1467 (N_1467,In_934,N_411);
nor U1468 (N_1468,N_391,In_1383);
xnor U1469 (N_1469,In_236,N_766);
nand U1470 (N_1470,N_768,N_244);
nand U1471 (N_1471,In_1432,N_207);
or U1472 (N_1472,N_656,In_1565);
nor U1473 (N_1473,In_1915,N_621);
or U1474 (N_1474,N_616,In_1967);
nand U1475 (N_1475,N_435,N_96);
xor U1476 (N_1476,In_1968,N_40);
xnor U1477 (N_1477,N_639,In_788);
nor U1478 (N_1478,N_388,In_1180);
nor U1479 (N_1479,N_348,In_1167);
and U1480 (N_1480,In_703,N_594);
nand U1481 (N_1481,N_745,In_1605);
or U1482 (N_1482,N_454,N_162);
or U1483 (N_1483,In_732,N_380);
nor U1484 (N_1484,N_548,N_704);
or U1485 (N_1485,In_1119,In_1024);
nand U1486 (N_1486,N_213,N_207);
nand U1487 (N_1487,In_1413,N_541);
nand U1488 (N_1488,N_544,In_685);
nor U1489 (N_1489,N_290,In_691);
xnor U1490 (N_1490,N_393,N_463);
xnor U1491 (N_1491,N_332,N_682);
nor U1492 (N_1492,In_685,N_183);
or U1493 (N_1493,N_794,N_678);
and U1494 (N_1494,In_1558,N_110);
or U1495 (N_1495,N_174,In_1458);
or U1496 (N_1496,N_470,N_743);
and U1497 (N_1497,In_534,In_1428);
nor U1498 (N_1498,In_1942,In_1784);
nand U1499 (N_1499,In_1366,N_264);
nand U1500 (N_1500,N_10,N_656);
and U1501 (N_1501,N_103,In_130);
and U1502 (N_1502,N_120,N_164);
xnor U1503 (N_1503,N_233,In_187);
nand U1504 (N_1504,In_447,N_751);
xnor U1505 (N_1505,N_293,N_38);
nor U1506 (N_1506,In_1456,N_465);
nor U1507 (N_1507,In_49,In_613);
and U1508 (N_1508,N_694,N_207);
and U1509 (N_1509,N_27,In_846);
nand U1510 (N_1510,In_1439,In_941);
nand U1511 (N_1511,N_793,N_219);
nor U1512 (N_1512,N_236,N_333);
and U1513 (N_1513,N_268,N_676);
or U1514 (N_1514,In_565,N_377);
or U1515 (N_1515,N_732,N_558);
or U1516 (N_1516,N_8,In_1556);
and U1517 (N_1517,N_7,N_619);
xor U1518 (N_1518,N_454,In_1216);
xor U1519 (N_1519,N_595,N_91);
nor U1520 (N_1520,N_26,In_1447);
and U1521 (N_1521,N_732,N_648);
xnor U1522 (N_1522,N_580,In_109);
xor U1523 (N_1523,In_1872,N_12);
and U1524 (N_1524,In_1841,N_768);
nor U1525 (N_1525,N_83,In_1007);
or U1526 (N_1526,In_1552,In_1751);
and U1527 (N_1527,In_701,In_671);
xnor U1528 (N_1528,N_80,N_26);
or U1529 (N_1529,N_329,N_546);
xnor U1530 (N_1530,N_222,N_719);
or U1531 (N_1531,In_1309,N_164);
nor U1532 (N_1532,In_111,N_4);
nor U1533 (N_1533,In_215,N_530);
xor U1534 (N_1534,In_1152,N_171);
xnor U1535 (N_1535,In_377,In_613);
nor U1536 (N_1536,N_11,N_511);
xor U1537 (N_1537,N_761,N_544);
or U1538 (N_1538,In_1602,N_56);
nor U1539 (N_1539,N_298,In_1424);
and U1540 (N_1540,N_140,N_122);
or U1541 (N_1541,N_209,N_554);
nor U1542 (N_1542,In_975,In_382);
xnor U1543 (N_1543,N_430,N_57);
and U1544 (N_1544,N_751,N_480);
nor U1545 (N_1545,N_333,N_122);
or U1546 (N_1546,N_6,In_1413);
and U1547 (N_1547,In_732,In_1942);
nor U1548 (N_1548,N_6,N_438);
xor U1549 (N_1549,N_721,N_315);
xnor U1550 (N_1550,N_320,In_416);
nand U1551 (N_1551,N_761,N_299);
nand U1552 (N_1552,N_455,N_647);
xor U1553 (N_1553,N_450,N_128);
or U1554 (N_1554,In_1164,N_799);
xnor U1555 (N_1555,N_263,N_539);
or U1556 (N_1556,N_562,N_64);
or U1557 (N_1557,N_783,In_521);
xor U1558 (N_1558,N_553,N_630);
or U1559 (N_1559,N_459,N_280);
and U1560 (N_1560,In_521,N_454);
xnor U1561 (N_1561,N_272,N_524);
or U1562 (N_1562,In_455,N_451);
and U1563 (N_1563,In_139,N_532);
and U1564 (N_1564,N_739,N_563);
xnor U1565 (N_1565,N_655,N_452);
nor U1566 (N_1566,N_61,N_749);
nand U1567 (N_1567,N_709,N_461);
nand U1568 (N_1568,N_755,N_567);
or U1569 (N_1569,N_589,In_1981);
xnor U1570 (N_1570,N_67,N_228);
nor U1571 (N_1571,In_1556,N_395);
nor U1572 (N_1572,N_238,N_313);
nor U1573 (N_1573,N_767,In_211);
xor U1574 (N_1574,N_168,In_1515);
xnor U1575 (N_1575,N_527,N_423);
nor U1576 (N_1576,N_360,N_17);
or U1577 (N_1577,In_995,N_22);
and U1578 (N_1578,In_1463,N_379);
and U1579 (N_1579,N_119,N_335);
nand U1580 (N_1580,N_294,N_325);
nand U1581 (N_1581,N_505,N_314);
and U1582 (N_1582,N_524,N_673);
and U1583 (N_1583,In_9,N_785);
nand U1584 (N_1584,N_248,N_370);
and U1585 (N_1585,N_701,In_783);
nor U1586 (N_1586,In_801,N_438);
and U1587 (N_1587,N_685,N_76);
and U1588 (N_1588,In_1305,In_42);
nand U1589 (N_1589,N_253,In_1640);
xnor U1590 (N_1590,In_102,In_1556);
and U1591 (N_1591,N_182,N_122);
xnor U1592 (N_1592,N_592,N_639);
xor U1593 (N_1593,In_188,N_667);
and U1594 (N_1594,N_393,N_487);
or U1595 (N_1595,N_595,N_54);
xnor U1596 (N_1596,In_890,N_456);
nand U1597 (N_1597,In_138,N_86);
or U1598 (N_1598,N_546,N_299);
nand U1599 (N_1599,In_1335,N_474);
nand U1600 (N_1600,N_1325,N_989);
and U1601 (N_1601,N_846,N_1391);
nor U1602 (N_1602,N_944,N_1159);
xnor U1603 (N_1603,N_1440,N_804);
or U1604 (N_1604,N_1192,N_1482);
nand U1605 (N_1605,N_887,N_878);
or U1606 (N_1606,N_986,N_1409);
and U1607 (N_1607,N_1278,N_1296);
or U1608 (N_1608,N_1102,N_1164);
nand U1609 (N_1609,N_1308,N_1042);
nand U1610 (N_1610,N_1585,N_979);
or U1611 (N_1611,N_876,N_1433);
xor U1612 (N_1612,N_906,N_1481);
nor U1613 (N_1613,N_1466,N_1485);
nor U1614 (N_1614,N_1380,N_828);
nor U1615 (N_1615,N_1024,N_1026);
nand U1616 (N_1616,N_1073,N_1108);
and U1617 (N_1617,N_961,N_1570);
or U1618 (N_1618,N_1511,N_1275);
nand U1619 (N_1619,N_1154,N_1177);
nor U1620 (N_1620,N_956,N_1175);
or U1621 (N_1621,N_1543,N_917);
nand U1622 (N_1622,N_1057,N_1513);
and U1623 (N_1623,N_1335,N_1051);
nand U1624 (N_1624,N_1349,N_931);
or U1625 (N_1625,N_1503,N_1030);
or U1626 (N_1626,N_1126,N_1002);
nor U1627 (N_1627,N_1070,N_1539);
nand U1628 (N_1628,N_1087,N_1082);
nor U1629 (N_1629,N_1427,N_1295);
and U1630 (N_1630,N_1138,N_1567);
nor U1631 (N_1631,N_992,N_1314);
or U1632 (N_1632,N_953,N_1183);
xnor U1633 (N_1633,N_1007,N_1517);
xor U1634 (N_1634,N_1495,N_1194);
nor U1635 (N_1635,N_1084,N_976);
xnor U1636 (N_1636,N_1459,N_991);
xnor U1637 (N_1637,N_1086,N_1050);
or U1638 (N_1638,N_1479,N_904);
nor U1639 (N_1639,N_845,N_1040);
and U1640 (N_1640,N_885,N_1430);
and U1641 (N_1641,N_1225,N_1301);
or U1642 (N_1642,N_945,N_1117);
xor U1643 (N_1643,N_1158,N_905);
xnor U1644 (N_1644,N_1285,N_1128);
nand U1645 (N_1645,N_823,N_1027);
nor U1646 (N_1646,N_872,N_1237);
and U1647 (N_1647,N_967,N_1003);
nor U1648 (N_1648,N_1548,N_1455);
xnor U1649 (N_1649,N_1269,N_890);
nor U1650 (N_1650,N_914,N_1208);
and U1651 (N_1651,N_1276,N_1119);
nand U1652 (N_1652,N_874,N_1371);
or U1653 (N_1653,N_1350,N_941);
or U1654 (N_1654,N_910,N_946);
nor U1655 (N_1655,N_1589,N_1254);
nand U1656 (N_1656,N_1018,N_1163);
nor U1657 (N_1657,N_1520,N_1417);
nand U1658 (N_1658,N_1207,N_1556);
nand U1659 (N_1659,N_1588,N_930);
nor U1660 (N_1660,N_1578,N_957);
nand U1661 (N_1661,N_896,N_1036);
nor U1662 (N_1662,N_1533,N_1586);
nand U1663 (N_1663,N_1025,N_1331);
or U1664 (N_1664,N_1069,N_1447);
or U1665 (N_1665,N_988,N_1354);
nor U1666 (N_1666,N_884,N_1442);
xnor U1667 (N_1667,N_1516,N_1429);
nand U1668 (N_1668,N_1133,N_1425);
xnor U1669 (N_1669,N_1483,N_1394);
nor U1670 (N_1670,N_1284,N_1351);
or U1671 (N_1671,N_1530,N_863);
and U1672 (N_1672,N_1508,N_934);
nor U1673 (N_1673,N_1205,N_1591);
nand U1674 (N_1674,N_907,N_1386);
nor U1675 (N_1675,N_812,N_1569);
nor U1676 (N_1676,N_1203,N_1410);
nand U1677 (N_1677,N_1582,N_870);
nor U1678 (N_1678,N_1487,N_857);
nand U1679 (N_1679,N_973,N_1273);
and U1680 (N_1680,N_1155,N_1151);
nor U1681 (N_1681,N_954,N_1162);
and U1682 (N_1682,N_1576,N_1390);
xor U1683 (N_1683,N_1400,N_1204);
nand U1684 (N_1684,N_1313,N_1226);
xnor U1685 (N_1685,N_1240,N_1507);
or U1686 (N_1686,N_983,N_1529);
and U1687 (N_1687,N_1232,N_1109);
xor U1688 (N_1688,N_1343,N_1063);
and U1689 (N_1689,N_1506,N_1143);
xor U1690 (N_1690,N_868,N_831);
nand U1691 (N_1691,N_1404,N_1480);
nor U1692 (N_1692,N_1004,N_958);
nand U1693 (N_1693,N_1497,N_1236);
or U1694 (N_1694,N_1422,N_1190);
or U1695 (N_1695,N_1388,N_1010);
nor U1696 (N_1696,N_1141,N_864);
or U1697 (N_1697,N_943,N_1258);
and U1698 (N_1698,N_925,N_1360);
nand U1699 (N_1699,N_1157,N_1406);
nand U1700 (N_1700,N_851,N_1235);
nand U1701 (N_1701,N_940,N_1502);
and U1702 (N_1702,N_1282,N_1596);
nor U1703 (N_1703,N_1542,N_1493);
or U1704 (N_1704,N_952,N_1393);
xnor U1705 (N_1705,N_955,N_1256);
and U1706 (N_1706,N_1423,N_877);
nor U1707 (N_1707,N_1176,N_1573);
or U1708 (N_1708,N_1131,N_1260);
nor U1709 (N_1709,N_1188,N_1228);
nor U1710 (N_1710,N_927,N_1415);
nand U1711 (N_1711,N_970,N_1242);
nor U1712 (N_1712,N_939,N_1037);
nor U1713 (N_1713,N_916,N_1230);
nor U1714 (N_1714,N_1211,N_1599);
xnor U1715 (N_1715,N_1174,N_1122);
nand U1716 (N_1716,N_1233,N_1247);
nor U1717 (N_1717,N_1463,N_996);
and U1718 (N_1718,N_922,N_1424);
and U1719 (N_1719,N_1555,N_1166);
nand U1720 (N_1720,N_1381,N_1315);
nor U1721 (N_1721,N_1562,N_1271);
xor U1722 (N_1722,N_1528,N_1035);
and U1723 (N_1723,N_817,N_1379);
xor U1724 (N_1724,N_1261,N_1241);
xnor U1725 (N_1725,N_1499,N_1475);
nand U1726 (N_1726,N_1121,N_1198);
nor U1727 (N_1727,N_1078,N_1054);
or U1728 (N_1728,N_1303,N_822);
and U1729 (N_1729,N_860,N_1098);
nand U1730 (N_1730,N_1310,N_1362);
nand U1731 (N_1731,N_1146,N_1074);
nand U1732 (N_1732,N_1344,N_835);
and U1733 (N_1733,N_1353,N_1547);
nand U1734 (N_1734,N_990,N_838);
nor U1735 (N_1735,N_1106,N_919);
nor U1736 (N_1736,N_1281,N_1199);
and U1737 (N_1737,N_1105,N_1178);
xor U1738 (N_1738,N_1514,N_1571);
nor U1739 (N_1739,N_1239,N_1246);
or U1740 (N_1740,N_1013,N_1540);
nor U1741 (N_1741,N_1093,N_1405);
xor U1742 (N_1742,N_1213,N_1292);
and U1743 (N_1743,N_901,N_848);
or U1744 (N_1744,N_1470,N_867);
or U1745 (N_1745,N_1549,N_1323);
and U1746 (N_1746,N_1557,N_1244);
or U1747 (N_1747,N_929,N_1434);
and U1748 (N_1748,N_1305,N_1012);
or U1749 (N_1749,N_994,N_993);
nor U1750 (N_1750,N_847,N_1515);
and U1751 (N_1751,N_814,N_886);
nor U1752 (N_1752,N_1420,N_1465);
nand U1753 (N_1753,N_1363,N_1496);
nand U1754 (N_1754,N_893,N_1412);
nand U1755 (N_1755,N_1243,N_1553);
nand U1756 (N_1756,N_1339,N_1094);
xnor U1757 (N_1757,N_1318,N_1577);
nor U1758 (N_1758,N_1195,N_1373);
xor U1759 (N_1759,N_1289,N_1361);
or U1760 (N_1760,N_1309,N_858);
nand U1761 (N_1761,N_1512,N_1227);
nand U1762 (N_1762,N_1060,N_869);
or U1763 (N_1763,N_1136,N_1359);
nand U1764 (N_1764,N_1152,N_1377);
and U1765 (N_1765,N_1378,N_1329);
or U1766 (N_1766,N_1510,N_1123);
and U1767 (N_1767,N_1001,N_1116);
xnor U1768 (N_1768,N_969,N_1172);
and U1769 (N_1769,N_843,N_1594);
or U1770 (N_1770,N_924,N_833);
and U1771 (N_1771,N_1565,N_1579);
nand U1772 (N_1772,N_1214,N_811);
and U1773 (N_1773,N_1398,N_1234);
nand U1774 (N_1774,N_1418,N_1118);
or U1775 (N_1775,N_1115,N_1229);
xor U1776 (N_1776,N_829,N_1357);
nand U1777 (N_1777,N_900,N_1397);
nand U1778 (N_1778,N_1376,N_1000);
or U1779 (N_1779,N_1079,N_1464);
or U1780 (N_1780,N_1491,N_1222);
nor U1781 (N_1781,N_1170,N_1469);
or U1782 (N_1782,N_1471,N_1268);
and U1783 (N_1783,N_1112,N_801);
and U1784 (N_1784,N_1330,N_1402);
and U1785 (N_1785,N_960,N_1161);
or U1786 (N_1786,N_1486,N_1392);
xnor U1787 (N_1787,N_1476,N_1169);
nor U1788 (N_1788,N_1092,N_1413);
or U1789 (N_1789,N_985,N_1532);
nor U1790 (N_1790,N_1221,N_1257);
nor U1791 (N_1791,N_1137,N_1210);
nor U1792 (N_1792,N_880,N_871);
or U1793 (N_1793,N_1428,N_816);
nand U1794 (N_1794,N_1045,N_1104);
nand U1795 (N_1795,N_807,N_1048);
or U1796 (N_1796,N_1139,N_1583);
xnor U1797 (N_1797,N_1441,N_855);
or U1798 (N_1798,N_1181,N_1089);
xor U1799 (N_1799,N_1551,N_1044);
and U1800 (N_1800,N_1168,N_808);
or U1801 (N_1801,N_959,N_1266);
or U1802 (N_1802,N_1322,N_1300);
or U1803 (N_1803,N_1262,N_1009);
nor U1804 (N_1804,N_1505,N_1135);
xor U1805 (N_1805,N_1457,N_1581);
or U1806 (N_1806,N_1191,N_1259);
or U1807 (N_1807,N_825,N_920);
xor U1808 (N_1808,N_1142,N_903);
nand U1809 (N_1809,N_1358,N_1075);
or U1810 (N_1810,N_1113,N_1103);
nand U1811 (N_1811,N_1435,N_1564);
or U1812 (N_1812,N_824,N_909);
nand U1813 (N_1813,N_923,N_1253);
and U1814 (N_1814,N_842,N_981);
or U1815 (N_1815,N_1348,N_854);
and U1816 (N_1816,N_1041,N_1531);
nor U1817 (N_1817,N_1572,N_1444);
nand U1818 (N_1818,N_1312,N_1374);
or U1819 (N_1819,N_1263,N_897);
nor U1820 (N_1820,N_1446,N_1065);
or U1821 (N_1821,N_971,N_1411);
and U1822 (N_1822,N_1382,N_911);
nand U1823 (N_1823,N_1272,N_1277);
nor U1824 (N_1824,N_1526,N_1081);
nand U1825 (N_1825,N_1458,N_1375);
xor U1826 (N_1826,N_899,N_936);
nor U1827 (N_1827,N_972,N_937);
xor U1828 (N_1828,N_1120,N_1552);
nand U1829 (N_1829,N_963,N_1460);
xnor U1830 (N_1830,N_1302,N_862);
or U1831 (N_1831,N_1453,N_1445);
nand U1832 (N_1832,N_1347,N_1316);
and U1833 (N_1833,N_1008,N_1288);
and U1834 (N_1834,N_1438,N_1150);
nand U1835 (N_1835,N_938,N_1127);
xor U1836 (N_1836,N_891,N_1341);
nand U1837 (N_1837,N_1206,N_1568);
and U1838 (N_1838,N_1280,N_1217);
and U1839 (N_1839,N_844,N_1215);
and U1840 (N_1840,N_1527,N_918);
xnor U1841 (N_1841,N_1015,N_1022);
or U1842 (N_1842,N_1299,N_1561);
nor U1843 (N_1843,N_1182,N_1202);
nand U1844 (N_1844,N_827,N_1432);
and U1845 (N_1845,N_1421,N_1283);
and U1846 (N_1846,N_1090,N_1047);
nand U1847 (N_1847,N_1148,N_1401);
xor U1848 (N_1848,N_875,N_1032);
nand U1849 (N_1849,N_1403,N_1267);
nor U1850 (N_1850,N_1574,N_1021);
and U1851 (N_1851,N_1144,N_1156);
xnor U1852 (N_1852,N_1248,N_1372);
nand U1853 (N_1853,N_1537,N_1255);
nand U1854 (N_1854,N_982,N_1028);
or U1855 (N_1855,N_881,N_942);
nor U1856 (N_1856,N_1500,N_1501);
and U1857 (N_1857,N_951,N_964);
xor U1858 (N_1858,N_865,N_1245);
xor U1859 (N_1859,N_1149,N_1212);
nand U1860 (N_1860,N_1326,N_1132);
xnor U1861 (N_1861,N_1327,N_1185);
and U1862 (N_1862,N_1130,N_902);
nor U1863 (N_1863,N_1307,N_1134);
nor U1864 (N_1864,N_1218,N_947);
nor U1865 (N_1865,N_1066,N_1153);
and U1866 (N_1866,N_1456,N_800);
xnor U1867 (N_1867,N_809,N_932);
and U1868 (N_1868,N_1100,N_1566);
or U1869 (N_1869,N_1598,N_1355);
or U1870 (N_1870,N_861,N_1319);
xor U1871 (N_1871,N_856,N_1451);
nor U1872 (N_1872,N_1597,N_1550);
nor U1873 (N_1873,N_1324,N_1370);
xor U1874 (N_1874,N_1467,N_1114);
xnor U1875 (N_1875,N_1095,N_1201);
and U1876 (N_1876,N_1472,N_818);
nand U1877 (N_1877,N_1016,N_1046);
xnor U1878 (N_1878,N_1165,N_1020);
nor U1879 (N_1879,N_1490,N_1590);
and U1880 (N_1880,N_1107,N_1193);
and U1881 (N_1881,N_1356,N_998);
and U1882 (N_1882,N_1068,N_1304);
nand U1883 (N_1883,N_1477,N_1279);
nor U1884 (N_1884,N_1538,N_873);
xor U1885 (N_1885,N_1297,N_995);
nand U1886 (N_1886,N_1448,N_813);
xnor U1887 (N_1887,N_1367,N_1039);
or U1888 (N_1888,N_1488,N_1408);
nand U1889 (N_1889,N_1333,N_1274);
and U1890 (N_1890,N_1223,N_1352);
and U1891 (N_1891,N_859,N_1005);
nor U1892 (N_1892,N_975,N_837);
or U1893 (N_1893,N_1238,N_1059);
and U1894 (N_1894,N_849,N_1336);
or U1895 (N_1895,N_1454,N_1384);
and U1896 (N_1896,N_841,N_1414);
or U1897 (N_1897,N_1088,N_1439);
nand U1898 (N_1898,N_1049,N_1593);
or U1899 (N_1899,N_1494,N_1364);
xor U1900 (N_1900,N_1224,N_1019);
and U1901 (N_1901,N_949,N_1167);
nor U1902 (N_1902,N_1265,N_1545);
or U1903 (N_1903,N_966,N_820);
or U1904 (N_1904,N_1067,N_1083);
nor U1905 (N_1905,N_1345,N_933);
xnor U1906 (N_1906,N_1473,N_826);
nor U1907 (N_1907,N_1216,N_1077);
xnor U1908 (N_1908,N_1076,N_1056);
and U1909 (N_1909,N_987,N_1575);
nor U1910 (N_1910,N_1431,N_1521);
and U1911 (N_1911,N_821,N_1160);
nor U1912 (N_1912,N_1072,N_1321);
nor U1913 (N_1913,N_965,N_1014);
nor U1914 (N_1914,N_889,N_1383);
or U1915 (N_1915,N_1320,N_1011);
xor U1916 (N_1916,N_1560,N_1559);
nor U1917 (N_1917,N_1580,N_1091);
and U1918 (N_1918,N_1209,N_1525);
nor U1919 (N_1919,N_1498,N_1450);
xor U1920 (N_1920,N_915,N_1332);
xor U1921 (N_1921,N_1536,N_908);
xor U1922 (N_1922,N_948,N_984);
and U1923 (N_1923,N_1058,N_935);
nor U1924 (N_1924,N_803,N_1298);
nand U1925 (N_1925,N_1395,N_1443);
xnor U1926 (N_1926,N_832,N_815);
xor U1927 (N_1927,N_1346,N_1171);
nand U1928 (N_1928,N_1071,N_1544);
nor U1929 (N_1929,N_1587,N_928);
and U1930 (N_1930,N_1173,N_882);
nor U1931 (N_1931,N_1061,N_1252);
or U1932 (N_1932,N_1426,N_962);
nand U1933 (N_1933,N_1437,N_1053);
and U1934 (N_1934,N_926,N_1524);
xor U1935 (N_1935,N_819,N_1184);
or U1936 (N_1936,N_1294,N_1449);
xnor U1937 (N_1937,N_1293,N_1125);
and U1938 (N_1938,N_1311,N_1522);
or U1939 (N_1939,N_1147,N_1064);
or U1940 (N_1940,N_1452,N_1196);
and U1941 (N_1941,N_834,N_1006);
nor U1942 (N_1942,N_1523,N_999);
xor U1943 (N_1943,N_1368,N_805);
xnor U1944 (N_1944,N_1029,N_1592);
nand U1945 (N_1945,N_1436,N_1110);
and U1946 (N_1946,N_892,N_913);
xnor U1947 (N_1947,N_1219,N_894);
nand U1948 (N_1948,N_1097,N_1478);
nand U1949 (N_1949,N_1340,N_850);
and U1950 (N_1950,N_1518,N_1563);
nand U1951 (N_1951,N_1220,N_980);
xor U1952 (N_1952,N_802,N_806);
nand U1953 (N_1953,N_1291,N_1369);
nand U1954 (N_1954,N_895,N_1186);
and U1955 (N_1955,N_1250,N_1558);
nor U1956 (N_1956,N_1101,N_1385);
or U1957 (N_1957,N_1334,N_1419);
nand U1958 (N_1958,N_1096,N_1145);
and U1959 (N_1959,N_1052,N_898);
nor U1960 (N_1960,N_1416,N_1554);
or U1961 (N_1961,N_1387,N_1033);
xor U1962 (N_1962,N_1342,N_1317);
or U1963 (N_1963,N_997,N_1129);
nand U1964 (N_1964,N_1038,N_1338);
nand U1965 (N_1965,N_852,N_1085);
xor U1966 (N_1966,N_1231,N_1062);
xor U1967 (N_1967,N_1189,N_866);
nand U1968 (N_1968,N_1251,N_1489);
and U1969 (N_1969,N_1462,N_839);
xor U1970 (N_1970,N_1468,N_1534);
nand U1971 (N_1971,N_1407,N_1124);
nand U1972 (N_1972,N_1541,N_968);
and U1973 (N_1973,N_1200,N_1306);
and U1974 (N_1974,N_1034,N_1474);
or U1975 (N_1975,N_1584,N_879);
nand U1976 (N_1976,N_1043,N_1509);
nor U1977 (N_1977,N_1365,N_912);
xor U1978 (N_1978,N_1519,N_883);
xnor U1979 (N_1979,N_1023,N_1595);
nand U1980 (N_1980,N_978,N_840);
and U1981 (N_1981,N_1080,N_1017);
or U1982 (N_1982,N_1504,N_950);
nor U1983 (N_1983,N_1031,N_1492);
and U1984 (N_1984,N_1389,N_1179);
or U1985 (N_1985,N_1111,N_1197);
xor U1986 (N_1986,N_921,N_1396);
xor U1987 (N_1987,N_1286,N_1180);
and U1988 (N_1988,N_836,N_1328);
xnor U1989 (N_1989,N_853,N_830);
nor U1990 (N_1990,N_1287,N_1399);
and U1991 (N_1991,N_810,N_1055);
xor U1992 (N_1992,N_888,N_1249);
and U1993 (N_1993,N_1290,N_1099);
nor U1994 (N_1994,N_1484,N_1535);
xnor U1995 (N_1995,N_1461,N_1366);
nor U1996 (N_1996,N_1337,N_1270);
xor U1997 (N_1997,N_1264,N_977);
xnor U1998 (N_1998,N_1546,N_1140);
and U1999 (N_1999,N_1187,N_974);
xnor U2000 (N_2000,N_1554,N_1390);
or U2001 (N_2001,N_1102,N_1444);
nand U2002 (N_2002,N_881,N_1485);
xor U2003 (N_2003,N_1419,N_1209);
xnor U2004 (N_2004,N_1514,N_814);
xor U2005 (N_2005,N_1430,N_1151);
xnor U2006 (N_2006,N_1170,N_1026);
xor U2007 (N_2007,N_1286,N_1484);
and U2008 (N_2008,N_946,N_1040);
xnor U2009 (N_2009,N_1581,N_857);
xnor U2010 (N_2010,N_1406,N_895);
or U2011 (N_2011,N_1270,N_1449);
xor U2012 (N_2012,N_1561,N_1588);
and U2013 (N_2013,N_1327,N_1295);
xnor U2014 (N_2014,N_1436,N_1425);
xnor U2015 (N_2015,N_1554,N_1316);
nor U2016 (N_2016,N_1161,N_1443);
xor U2017 (N_2017,N_868,N_1253);
nand U2018 (N_2018,N_1341,N_1422);
and U2019 (N_2019,N_1093,N_806);
or U2020 (N_2020,N_1018,N_849);
nand U2021 (N_2021,N_1204,N_1506);
nor U2022 (N_2022,N_1543,N_1560);
and U2023 (N_2023,N_1527,N_1222);
nand U2024 (N_2024,N_1156,N_1307);
or U2025 (N_2025,N_1218,N_1404);
nor U2026 (N_2026,N_1304,N_991);
xor U2027 (N_2027,N_1311,N_1332);
and U2028 (N_2028,N_1557,N_1482);
xnor U2029 (N_2029,N_1586,N_1094);
or U2030 (N_2030,N_1398,N_1168);
or U2031 (N_2031,N_1347,N_857);
and U2032 (N_2032,N_1392,N_1570);
nor U2033 (N_2033,N_1173,N_1204);
or U2034 (N_2034,N_1315,N_1364);
xor U2035 (N_2035,N_837,N_1215);
and U2036 (N_2036,N_1380,N_1256);
and U2037 (N_2037,N_1351,N_962);
nand U2038 (N_2038,N_1099,N_1091);
or U2039 (N_2039,N_1016,N_979);
and U2040 (N_2040,N_826,N_1527);
or U2041 (N_2041,N_1501,N_1288);
or U2042 (N_2042,N_1328,N_1542);
and U2043 (N_2043,N_1187,N_1387);
and U2044 (N_2044,N_845,N_834);
nand U2045 (N_2045,N_832,N_1124);
or U2046 (N_2046,N_1187,N_1390);
nand U2047 (N_2047,N_959,N_1212);
or U2048 (N_2048,N_1209,N_826);
nand U2049 (N_2049,N_1546,N_1211);
nor U2050 (N_2050,N_1519,N_1284);
nand U2051 (N_2051,N_1209,N_1257);
or U2052 (N_2052,N_1064,N_924);
xnor U2053 (N_2053,N_1306,N_1260);
xnor U2054 (N_2054,N_1085,N_1580);
and U2055 (N_2055,N_1092,N_955);
or U2056 (N_2056,N_1004,N_1461);
and U2057 (N_2057,N_1184,N_1246);
and U2058 (N_2058,N_1312,N_1361);
nand U2059 (N_2059,N_1197,N_1449);
nand U2060 (N_2060,N_1373,N_1338);
nand U2061 (N_2061,N_1233,N_1241);
nor U2062 (N_2062,N_944,N_862);
and U2063 (N_2063,N_1202,N_1377);
and U2064 (N_2064,N_1049,N_1062);
xnor U2065 (N_2065,N_857,N_926);
or U2066 (N_2066,N_867,N_1246);
nand U2067 (N_2067,N_1413,N_1019);
or U2068 (N_2068,N_1501,N_1362);
nor U2069 (N_2069,N_1066,N_1388);
or U2070 (N_2070,N_905,N_960);
nor U2071 (N_2071,N_1368,N_1014);
xnor U2072 (N_2072,N_1228,N_1101);
or U2073 (N_2073,N_1549,N_1050);
nor U2074 (N_2074,N_988,N_871);
nand U2075 (N_2075,N_823,N_1223);
and U2076 (N_2076,N_1574,N_1308);
nor U2077 (N_2077,N_926,N_1405);
xor U2078 (N_2078,N_1587,N_1104);
or U2079 (N_2079,N_827,N_1038);
and U2080 (N_2080,N_1321,N_1048);
nand U2081 (N_2081,N_1241,N_934);
nand U2082 (N_2082,N_1002,N_1243);
and U2083 (N_2083,N_1425,N_1261);
or U2084 (N_2084,N_933,N_1188);
nor U2085 (N_2085,N_1294,N_1380);
xor U2086 (N_2086,N_1518,N_1395);
nand U2087 (N_2087,N_968,N_1092);
nand U2088 (N_2088,N_854,N_1216);
and U2089 (N_2089,N_805,N_1015);
nor U2090 (N_2090,N_1048,N_829);
or U2091 (N_2091,N_1267,N_1284);
nand U2092 (N_2092,N_866,N_1275);
nor U2093 (N_2093,N_947,N_1030);
nor U2094 (N_2094,N_1596,N_1206);
or U2095 (N_2095,N_1356,N_1449);
nand U2096 (N_2096,N_1247,N_1169);
or U2097 (N_2097,N_1394,N_905);
nor U2098 (N_2098,N_1385,N_1112);
nand U2099 (N_2099,N_922,N_1119);
and U2100 (N_2100,N_1060,N_1040);
nand U2101 (N_2101,N_1319,N_1105);
xnor U2102 (N_2102,N_1515,N_1091);
nand U2103 (N_2103,N_1310,N_977);
nand U2104 (N_2104,N_1292,N_993);
nand U2105 (N_2105,N_1254,N_1415);
or U2106 (N_2106,N_1560,N_896);
nor U2107 (N_2107,N_1205,N_986);
and U2108 (N_2108,N_979,N_963);
and U2109 (N_2109,N_1248,N_1420);
and U2110 (N_2110,N_1123,N_1286);
nand U2111 (N_2111,N_1239,N_1359);
nand U2112 (N_2112,N_878,N_1400);
or U2113 (N_2113,N_1522,N_1350);
or U2114 (N_2114,N_1565,N_1273);
nor U2115 (N_2115,N_1521,N_1595);
nor U2116 (N_2116,N_995,N_1341);
nand U2117 (N_2117,N_964,N_910);
xnor U2118 (N_2118,N_1297,N_859);
nand U2119 (N_2119,N_1117,N_1172);
and U2120 (N_2120,N_1494,N_1195);
and U2121 (N_2121,N_1093,N_1271);
or U2122 (N_2122,N_1324,N_966);
and U2123 (N_2123,N_951,N_870);
xnor U2124 (N_2124,N_1001,N_1054);
or U2125 (N_2125,N_1109,N_1293);
and U2126 (N_2126,N_967,N_1475);
xnor U2127 (N_2127,N_1357,N_1098);
nor U2128 (N_2128,N_1194,N_921);
and U2129 (N_2129,N_1479,N_1269);
xnor U2130 (N_2130,N_1306,N_1147);
and U2131 (N_2131,N_1599,N_860);
nor U2132 (N_2132,N_1267,N_925);
xnor U2133 (N_2133,N_1523,N_1079);
nand U2134 (N_2134,N_1168,N_1204);
and U2135 (N_2135,N_1156,N_925);
and U2136 (N_2136,N_1339,N_1512);
and U2137 (N_2137,N_913,N_1189);
or U2138 (N_2138,N_1206,N_1186);
nor U2139 (N_2139,N_1402,N_1069);
nand U2140 (N_2140,N_1596,N_922);
nor U2141 (N_2141,N_1127,N_1390);
nor U2142 (N_2142,N_1264,N_840);
nor U2143 (N_2143,N_1593,N_993);
xnor U2144 (N_2144,N_874,N_1099);
nor U2145 (N_2145,N_961,N_1577);
and U2146 (N_2146,N_1196,N_1127);
nor U2147 (N_2147,N_1438,N_807);
nand U2148 (N_2148,N_1368,N_1031);
nor U2149 (N_2149,N_1477,N_1444);
nor U2150 (N_2150,N_1023,N_1050);
xor U2151 (N_2151,N_1315,N_1564);
and U2152 (N_2152,N_811,N_1074);
nand U2153 (N_2153,N_1318,N_1332);
nor U2154 (N_2154,N_1564,N_839);
nor U2155 (N_2155,N_1041,N_1187);
xor U2156 (N_2156,N_1380,N_1086);
xnor U2157 (N_2157,N_1223,N_1366);
xnor U2158 (N_2158,N_1332,N_1438);
nor U2159 (N_2159,N_1279,N_1196);
nand U2160 (N_2160,N_1129,N_969);
nor U2161 (N_2161,N_1476,N_990);
nor U2162 (N_2162,N_1154,N_1339);
and U2163 (N_2163,N_1180,N_1212);
nor U2164 (N_2164,N_1190,N_1251);
and U2165 (N_2165,N_1480,N_1252);
or U2166 (N_2166,N_1184,N_1175);
or U2167 (N_2167,N_932,N_1512);
xor U2168 (N_2168,N_1119,N_876);
xor U2169 (N_2169,N_1472,N_1170);
or U2170 (N_2170,N_1413,N_1069);
nor U2171 (N_2171,N_967,N_1120);
or U2172 (N_2172,N_1318,N_1322);
nor U2173 (N_2173,N_823,N_1106);
or U2174 (N_2174,N_1068,N_1172);
or U2175 (N_2175,N_977,N_891);
or U2176 (N_2176,N_1488,N_1543);
or U2177 (N_2177,N_1381,N_1114);
xnor U2178 (N_2178,N_1248,N_1155);
or U2179 (N_2179,N_1373,N_935);
xor U2180 (N_2180,N_862,N_1328);
or U2181 (N_2181,N_1151,N_1538);
nor U2182 (N_2182,N_881,N_1215);
nor U2183 (N_2183,N_1233,N_937);
and U2184 (N_2184,N_1076,N_1546);
xor U2185 (N_2185,N_1382,N_801);
and U2186 (N_2186,N_968,N_1314);
and U2187 (N_2187,N_1247,N_1117);
nor U2188 (N_2188,N_878,N_1431);
nand U2189 (N_2189,N_868,N_1433);
xor U2190 (N_2190,N_1076,N_826);
nor U2191 (N_2191,N_1085,N_1046);
and U2192 (N_2192,N_1092,N_1269);
nand U2193 (N_2193,N_1297,N_1323);
nand U2194 (N_2194,N_1085,N_1408);
or U2195 (N_2195,N_880,N_1079);
and U2196 (N_2196,N_1134,N_1527);
nand U2197 (N_2197,N_1179,N_945);
xnor U2198 (N_2198,N_1546,N_1529);
xor U2199 (N_2199,N_1559,N_1015);
nand U2200 (N_2200,N_1452,N_1230);
or U2201 (N_2201,N_1004,N_909);
and U2202 (N_2202,N_821,N_1509);
nor U2203 (N_2203,N_1463,N_1262);
nand U2204 (N_2204,N_981,N_1426);
xor U2205 (N_2205,N_1395,N_1097);
nand U2206 (N_2206,N_1193,N_1464);
xor U2207 (N_2207,N_1202,N_1324);
and U2208 (N_2208,N_927,N_1204);
or U2209 (N_2209,N_1083,N_1198);
xnor U2210 (N_2210,N_1243,N_973);
xor U2211 (N_2211,N_1024,N_1105);
nand U2212 (N_2212,N_956,N_1210);
nor U2213 (N_2213,N_1006,N_1216);
and U2214 (N_2214,N_1347,N_1472);
xnor U2215 (N_2215,N_891,N_1233);
or U2216 (N_2216,N_1330,N_821);
nand U2217 (N_2217,N_821,N_1599);
or U2218 (N_2218,N_1584,N_1359);
nand U2219 (N_2219,N_862,N_1436);
nand U2220 (N_2220,N_1141,N_1411);
nand U2221 (N_2221,N_977,N_845);
xnor U2222 (N_2222,N_1415,N_815);
nor U2223 (N_2223,N_1254,N_1116);
xnor U2224 (N_2224,N_965,N_1325);
xor U2225 (N_2225,N_1280,N_1178);
nand U2226 (N_2226,N_1036,N_1551);
and U2227 (N_2227,N_1177,N_1123);
nand U2228 (N_2228,N_1232,N_844);
nand U2229 (N_2229,N_1456,N_960);
and U2230 (N_2230,N_1397,N_1476);
and U2231 (N_2231,N_1401,N_904);
and U2232 (N_2232,N_1569,N_948);
and U2233 (N_2233,N_1501,N_1310);
nor U2234 (N_2234,N_1207,N_1568);
nor U2235 (N_2235,N_1428,N_1472);
nor U2236 (N_2236,N_1368,N_1581);
or U2237 (N_2237,N_1356,N_1345);
or U2238 (N_2238,N_999,N_1298);
xor U2239 (N_2239,N_1449,N_1345);
or U2240 (N_2240,N_1321,N_1550);
xnor U2241 (N_2241,N_1006,N_1198);
nand U2242 (N_2242,N_1373,N_1244);
nor U2243 (N_2243,N_1239,N_832);
xnor U2244 (N_2244,N_961,N_1054);
xnor U2245 (N_2245,N_1504,N_1185);
or U2246 (N_2246,N_1410,N_838);
xnor U2247 (N_2247,N_1364,N_1473);
and U2248 (N_2248,N_1174,N_974);
xnor U2249 (N_2249,N_933,N_1096);
nand U2250 (N_2250,N_1090,N_1495);
nand U2251 (N_2251,N_1318,N_1041);
nor U2252 (N_2252,N_951,N_818);
and U2253 (N_2253,N_1119,N_1322);
and U2254 (N_2254,N_1466,N_1431);
xor U2255 (N_2255,N_1332,N_1251);
or U2256 (N_2256,N_1556,N_1005);
nor U2257 (N_2257,N_1366,N_927);
nand U2258 (N_2258,N_1020,N_1084);
nor U2259 (N_2259,N_1210,N_910);
nand U2260 (N_2260,N_1512,N_1064);
nor U2261 (N_2261,N_1519,N_1153);
and U2262 (N_2262,N_1512,N_1351);
and U2263 (N_2263,N_1442,N_982);
xor U2264 (N_2264,N_1423,N_988);
nor U2265 (N_2265,N_1535,N_872);
xnor U2266 (N_2266,N_1598,N_1425);
xnor U2267 (N_2267,N_909,N_858);
and U2268 (N_2268,N_1487,N_932);
or U2269 (N_2269,N_801,N_1196);
and U2270 (N_2270,N_1203,N_1388);
and U2271 (N_2271,N_1008,N_1290);
nor U2272 (N_2272,N_1370,N_1250);
xnor U2273 (N_2273,N_877,N_1400);
or U2274 (N_2274,N_1512,N_1320);
nand U2275 (N_2275,N_903,N_1186);
or U2276 (N_2276,N_1115,N_1156);
and U2277 (N_2277,N_805,N_980);
or U2278 (N_2278,N_867,N_1216);
xnor U2279 (N_2279,N_1446,N_1131);
xnor U2280 (N_2280,N_1125,N_1403);
and U2281 (N_2281,N_1220,N_1173);
nand U2282 (N_2282,N_962,N_824);
or U2283 (N_2283,N_1479,N_1236);
nor U2284 (N_2284,N_1076,N_1298);
xor U2285 (N_2285,N_853,N_911);
xnor U2286 (N_2286,N_1250,N_841);
and U2287 (N_2287,N_1395,N_897);
nor U2288 (N_2288,N_1377,N_997);
nor U2289 (N_2289,N_1159,N_1081);
nand U2290 (N_2290,N_1188,N_860);
nand U2291 (N_2291,N_964,N_1273);
xor U2292 (N_2292,N_1152,N_1393);
nor U2293 (N_2293,N_978,N_831);
nand U2294 (N_2294,N_1187,N_868);
xor U2295 (N_2295,N_1128,N_1453);
or U2296 (N_2296,N_1362,N_898);
xnor U2297 (N_2297,N_1044,N_1144);
nand U2298 (N_2298,N_1409,N_1057);
nor U2299 (N_2299,N_1550,N_1186);
nand U2300 (N_2300,N_904,N_1062);
and U2301 (N_2301,N_984,N_982);
nand U2302 (N_2302,N_1285,N_1356);
and U2303 (N_2303,N_1076,N_1528);
xor U2304 (N_2304,N_1147,N_1011);
xnor U2305 (N_2305,N_1084,N_1097);
and U2306 (N_2306,N_1579,N_1064);
or U2307 (N_2307,N_1402,N_1182);
nand U2308 (N_2308,N_1540,N_1299);
xnor U2309 (N_2309,N_1117,N_1448);
xor U2310 (N_2310,N_1035,N_985);
xnor U2311 (N_2311,N_1091,N_1422);
or U2312 (N_2312,N_850,N_1258);
nor U2313 (N_2313,N_1465,N_874);
nand U2314 (N_2314,N_1510,N_1379);
nand U2315 (N_2315,N_816,N_1567);
nand U2316 (N_2316,N_1014,N_1450);
xnor U2317 (N_2317,N_1582,N_1251);
and U2318 (N_2318,N_926,N_804);
nand U2319 (N_2319,N_1004,N_1371);
nor U2320 (N_2320,N_1391,N_1361);
xor U2321 (N_2321,N_1301,N_1082);
nor U2322 (N_2322,N_936,N_839);
and U2323 (N_2323,N_1162,N_821);
or U2324 (N_2324,N_965,N_999);
nor U2325 (N_2325,N_1123,N_1209);
xor U2326 (N_2326,N_1003,N_1566);
nor U2327 (N_2327,N_1447,N_1439);
nor U2328 (N_2328,N_1425,N_1574);
or U2329 (N_2329,N_945,N_815);
nor U2330 (N_2330,N_1560,N_1506);
or U2331 (N_2331,N_1577,N_1426);
nor U2332 (N_2332,N_1563,N_859);
nor U2333 (N_2333,N_1485,N_1515);
nor U2334 (N_2334,N_1468,N_1037);
nand U2335 (N_2335,N_1231,N_1501);
and U2336 (N_2336,N_1102,N_1119);
and U2337 (N_2337,N_1474,N_1032);
and U2338 (N_2338,N_1161,N_1556);
or U2339 (N_2339,N_1590,N_1414);
nor U2340 (N_2340,N_902,N_1120);
or U2341 (N_2341,N_979,N_878);
nand U2342 (N_2342,N_1257,N_1332);
and U2343 (N_2343,N_1264,N_1111);
nand U2344 (N_2344,N_1572,N_1483);
xor U2345 (N_2345,N_1206,N_898);
or U2346 (N_2346,N_893,N_1098);
xor U2347 (N_2347,N_1329,N_878);
nand U2348 (N_2348,N_814,N_1387);
or U2349 (N_2349,N_898,N_1257);
or U2350 (N_2350,N_1076,N_1052);
and U2351 (N_2351,N_1225,N_1481);
nand U2352 (N_2352,N_974,N_965);
and U2353 (N_2353,N_1481,N_1263);
and U2354 (N_2354,N_1186,N_813);
xnor U2355 (N_2355,N_1365,N_1261);
nor U2356 (N_2356,N_871,N_1538);
nand U2357 (N_2357,N_1044,N_1530);
nor U2358 (N_2358,N_1383,N_1117);
nor U2359 (N_2359,N_1088,N_1140);
and U2360 (N_2360,N_1186,N_1459);
xnor U2361 (N_2361,N_1365,N_1075);
and U2362 (N_2362,N_1226,N_1287);
nor U2363 (N_2363,N_1412,N_1269);
xnor U2364 (N_2364,N_969,N_966);
xnor U2365 (N_2365,N_1139,N_822);
or U2366 (N_2366,N_1562,N_1061);
nor U2367 (N_2367,N_1003,N_1496);
xor U2368 (N_2368,N_1152,N_1480);
xnor U2369 (N_2369,N_1097,N_865);
xnor U2370 (N_2370,N_1330,N_1424);
nor U2371 (N_2371,N_1149,N_1349);
or U2372 (N_2372,N_1409,N_887);
nand U2373 (N_2373,N_1088,N_1326);
nor U2374 (N_2374,N_1391,N_1303);
nand U2375 (N_2375,N_1261,N_1236);
and U2376 (N_2376,N_1412,N_1452);
or U2377 (N_2377,N_1472,N_849);
nor U2378 (N_2378,N_1387,N_1467);
or U2379 (N_2379,N_1474,N_1533);
nor U2380 (N_2380,N_1420,N_1164);
or U2381 (N_2381,N_1313,N_830);
and U2382 (N_2382,N_1291,N_1120);
or U2383 (N_2383,N_1599,N_1438);
nand U2384 (N_2384,N_824,N_967);
nand U2385 (N_2385,N_1498,N_1181);
or U2386 (N_2386,N_1049,N_1326);
and U2387 (N_2387,N_845,N_940);
and U2388 (N_2388,N_1451,N_974);
nand U2389 (N_2389,N_1435,N_990);
nand U2390 (N_2390,N_1142,N_1042);
nand U2391 (N_2391,N_1308,N_875);
xor U2392 (N_2392,N_1247,N_1290);
or U2393 (N_2393,N_1481,N_1074);
nand U2394 (N_2394,N_906,N_1401);
or U2395 (N_2395,N_873,N_1067);
nor U2396 (N_2396,N_1062,N_888);
nor U2397 (N_2397,N_802,N_839);
and U2398 (N_2398,N_1095,N_1429);
and U2399 (N_2399,N_1103,N_923);
nor U2400 (N_2400,N_2399,N_1782);
or U2401 (N_2401,N_1742,N_1720);
or U2402 (N_2402,N_2028,N_2397);
nand U2403 (N_2403,N_1728,N_1979);
xor U2404 (N_2404,N_1666,N_1888);
and U2405 (N_2405,N_1625,N_1818);
or U2406 (N_2406,N_1774,N_2193);
nand U2407 (N_2407,N_1982,N_2191);
xor U2408 (N_2408,N_2051,N_1848);
nand U2409 (N_2409,N_1667,N_1948);
nand U2410 (N_2410,N_2016,N_1965);
and U2411 (N_2411,N_2012,N_1943);
xor U2412 (N_2412,N_2009,N_1622);
or U2413 (N_2413,N_2286,N_1897);
nor U2414 (N_2414,N_1709,N_1820);
nand U2415 (N_2415,N_1604,N_2253);
nand U2416 (N_2416,N_1613,N_1712);
nor U2417 (N_2417,N_1792,N_1879);
nor U2418 (N_2418,N_2331,N_2206);
or U2419 (N_2419,N_1748,N_1702);
nor U2420 (N_2420,N_1843,N_2002);
nor U2421 (N_2421,N_2186,N_1877);
nor U2422 (N_2422,N_2116,N_2061);
nor U2423 (N_2423,N_2326,N_1734);
and U2424 (N_2424,N_2379,N_1911);
nor U2425 (N_2425,N_2369,N_2315);
xor U2426 (N_2426,N_2351,N_1885);
xor U2427 (N_2427,N_1790,N_2292);
nand U2428 (N_2428,N_2144,N_2333);
and U2429 (N_2429,N_1713,N_1937);
nand U2430 (N_2430,N_1696,N_1612);
nor U2431 (N_2431,N_1851,N_1983);
and U2432 (N_2432,N_2393,N_1685);
and U2433 (N_2433,N_1862,N_1936);
nor U2434 (N_2434,N_2278,N_1619);
xor U2435 (N_2435,N_1989,N_2394);
or U2436 (N_2436,N_2324,N_2280);
xnor U2437 (N_2437,N_1947,N_2110);
or U2438 (N_2438,N_2041,N_2014);
nor U2439 (N_2439,N_1892,N_2141);
xor U2440 (N_2440,N_2355,N_1896);
nor U2441 (N_2441,N_2335,N_2045);
and U2442 (N_2442,N_1973,N_2025);
and U2443 (N_2443,N_2100,N_1976);
or U2444 (N_2444,N_1995,N_2354);
xnor U2445 (N_2445,N_2299,N_2010);
and U2446 (N_2446,N_1624,N_2107);
nor U2447 (N_2447,N_1717,N_2087);
nor U2448 (N_2448,N_2273,N_1699);
or U2449 (N_2449,N_1985,N_2063);
nand U2450 (N_2450,N_1856,N_2180);
xor U2451 (N_2451,N_1700,N_1865);
nand U2452 (N_2452,N_1932,N_1652);
and U2453 (N_2453,N_2173,N_1750);
nor U2454 (N_2454,N_1978,N_2308);
xor U2455 (N_2455,N_2079,N_2313);
nor U2456 (N_2456,N_2264,N_1769);
nor U2457 (N_2457,N_2189,N_2375);
nand U2458 (N_2458,N_1955,N_1770);
nor U2459 (N_2459,N_1736,N_2266);
nor U2460 (N_2460,N_1649,N_1646);
nor U2461 (N_2461,N_2279,N_1881);
nor U2462 (N_2462,N_2203,N_1814);
xor U2463 (N_2463,N_1807,N_2175);
xor U2464 (N_2464,N_2001,N_2139);
and U2465 (N_2465,N_2338,N_2167);
nor U2466 (N_2466,N_1678,N_1762);
xnor U2467 (N_2467,N_1775,N_1751);
xor U2468 (N_2468,N_2118,N_2162);
nand U2469 (N_2469,N_2004,N_1781);
nand U2470 (N_2470,N_2199,N_2312);
nand U2471 (N_2471,N_1930,N_2201);
and U2472 (N_2472,N_2020,N_1924);
and U2473 (N_2473,N_2074,N_2123);
or U2474 (N_2474,N_1721,N_1919);
nor U2475 (N_2475,N_2067,N_2213);
nor U2476 (N_2476,N_1795,N_1954);
and U2477 (N_2477,N_2194,N_1939);
xor U2478 (N_2478,N_2026,N_2384);
nor U2479 (N_2479,N_2361,N_2306);
and U2480 (N_2480,N_1616,N_2108);
xnor U2481 (N_2481,N_2391,N_2080);
xnor U2482 (N_2482,N_1796,N_2293);
nor U2483 (N_2483,N_2225,N_2115);
and U2484 (N_2484,N_2322,N_1971);
and U2485 (N_2485,N_1968,N_2210);
nand U2486 (N_2486,N_2353,N_1910);
or U2487 (N_2487,N_1815,N_2091);
or U2488 (N_2488,N_2284,N_1600);
nand U2489 (N_2489,N_2276,N_2196);
nor U2490 (N_2490,N_1785,N_1715);
nand U2491 (N_2491,N_2321,N_1833);
xnor U2492 (N_2492,N_2140,N_2296);
nand U2493 (N_2493,N_1768,N_2114);
or U2494 (N_2494,N_2095,N_1811);
xor U2495 (N_2495,N_2132,N_2068);
nand U2496 (N_2496,N_2054,N_2064);
and U2497 (N_2497,N_1810,N_2065);
nand U2498 (N_2498,N_1732,N_1628);
and U2499 (N_2499,N_2269,N_2272);
nand U2500 (N_2500,N_1706,N_1642);
nand U2501 (N_2501,N_2268,N_2147);
xnor U2502 (N_2502,N_1730,N_2122);
or U2503 (N_2503,N_2006,N_1964);
xor U2504 (N_2504,N_2195,N_2005);
or U2505 (N_2505,N_2137,N_1725);
and U2506 (N_2506,N_1823,N_1671);
and U2507 (N_2507,N_2257,N_2128);
or U2508 (N_2508,N_1940,N_2022);
and U2509 (N_2509,N_2138,N_1743);
or U2510 (N_2510,N_1708,N_2184);
nor U2511 (N_2511,N_1765,N_1780);
xnor U2512 (N_2512,N_1640,N_1605);
and U2513 (N_2513,N_2183,N_2161);
xor U2514 (N_2514,N_1962,N_2092);
or U2515 (N_2515,N_1857,N_2304);
nand U2516 (N_2516,N_2251,N_2145);
or U2517 (N_2517,N_1816,N_1680);
or U2518 (N_2518,N_1959,N_2356);
nand U2519 (N_2519,N_2218,N_1805);
or U2520 (N_2520,N_2370,N_2382);
nand U2521 (N_2521,N_2176,N_1934);
xnor U2522 (N_2522,N_2245,N_2236);
and U2523 (N_2523,N_1657,N_2238);
nand U2524 (N_2524,N_2047,N_2055);
and U2525 (N_2525,N_1942,N_1891);
or U2526 (N_2526,N_1786,N_1791);
xor U2527 (N_2527,N_1963,N_1872);
nor U2528 (N_2528,N_2076,N_2221);
xor U2529 (N_2529,N_2015,N_2059);
nand U2530 (N_2530,N_2385,N_2259);
and U2531 (N_2531,N_1867,N_1997);
or U2532 (N_2532,N_2301,N_1996);
nand U2533 (N_2533,N_1798,N_1858);
or U2534 (N_2534,N_2159,N_1623);
nor U2535 (N_2535,N_1890,N_1821);
and U2536 (N_2536,N_1853,N_2237);
nor U2537 (N_2537,N_1710,N_2233);
or U2538 (N_2538,N_1912,N_1784);
nand U2539 (N_2539,N_1724,N_1689);
xor U2540 (N_2540,N_2071,N_2177);
xor U2541 (N_2541,N_2377,N_2214);
nor U2542 (N_2542,N_2359,N_2152);
nor U2543 (N_2543,N_2208,N_2367);
nor U2544 (N_2544,N_2003,N_1847);
and U2545 (N_2545,N_1882,N_1922);
or U2546 (N_2546,N_1719,N_2120);
xnor U2547 (N_2547,N_2376,N_1644);
xnor U2548 (N_2548,N_2182,N_2096);
nand U2549 (N_2549,N_1634,N_1741);
or U2550 (N_2550,N_1916,N_1835);
or U2551 (N_2551,N_2142,N_1793);
or U2552 (N_2552,N_2261,N_2275);
nand U2553 (N_2553,N_1905,N_1895);
and U2554 (N_2554,N_2274,N_2277);
nand U2555 (N_2555,N_1660,N_2033);
and U2556 (N_2556,N_1904,N_2227);
xor U2557 (N_2557,N_2171,N_1999);
and U2558 (N_2558,N_2255,N_1672);
xnor U2559 (N_2559,N_2373,N_2102);
or U2560 (N_2560,N_2126,N_1906);
or U2561 (N_2561,N_1630,N_1740);
nor U2562 (N_2562,N_1880,N_2216);
nand U2563 (N_2563,N_2097,N_1834);
xor U2564 (N_2564,N_2242,N_2166);
or U2565 (N_2565,N_2066,N_2050);
xnor U2566 (N_2566,N_2042,N_2111);
nor U2567 (N_2567,N_1961,N_2371);
or U2568 (N_2568,N_2327,N_1687);
nor U2569 (N_2569,N_1803,N_1938);
or U2570 (N_2570,N_2179,N_1878);
nand U2571 (N_2571,N_1944,N_2392);
nor U2572 (N_2572,N_1866,N_1871);
and U2573 (N_2573,N_2156,N_1733);
and U2574 (N_2574,N_2256,N_1650);
or U2575 (N_2575,N_1675,N_2358);
and U2576 (N_2576,N_1998,N_1714);
or U2577 (N_2577,N_2307,N_2048);
nand U2578 (N_2578,N_2360,N_1850);
and U2579 (N_2579,N_1974,N_1674);
or U2580 (N_2580,N_1663,N_2085);
nand U2581 (N_2581,N_1773,N_2000);
or U2582 (N_2582,N_1779,N_2127);
xor U2583 (N_2583,N_1837,N_2038);
xnor U2584 (N_2584,N_2336,N_2368);
or U2585 (N_2585,N_1977,N_1928);
or U2586 (N_2586,N_1949,N_1697);
nor U2587 (N_2587,N_1681,N_2332);
or U2588 (N_2588,N_1822,N_1950);
and U2589 (N_2589,N_1711,N_2270);
nand U2590 (N_2590,N_1927,N_1960);
and U2591 (N_2591,N_1956,N_1987);
nand U2592 (N_2592,N_1984,N_1637);
and U2593 (N_2593,N_1925,N_2036);
nor U2594 (N_2594,N_1731,N_2205);
and U2595 (N_2595,N_2220,N_2084);
nand U2596 (N_2596,N_2346,N_2252);
nor U2597 (N_2597,N_1836,N_2007);
xor U2598 (N_2598,N_2239,N_2146);
and U2599 (N_2599,N_1898,N_2188);
nand U2600 (N_2600,N_2112,N_2232);
nand U2601 (N_2601,N_2058,N_1855);
and U2602 (N_2602,N_2357,N_2072);
or U2603 (N_2603,N_2034,N_2363);
nor U2604 (N_2604,N_1991,N_2297);
xnor U2605 (N_2605,N_2130,N_1698);
nor U2606 (N_2606,N_1693,N_1869);
nand U2607 (N_2607,N_2030,N_2135);
nand U2608 (N_2608,N_2150,N_1726);
xor U2609 (N_2609,N_1975,N_1718);
nand U2610 (N_2610,N_2329,N_2035);
or U2611 (N_2611,N_1966,N_2386);
nand U2612 (N_2612,N_1990,N_2300);
nor U2613 (N_2613,N_2073,N_1679);
and U2614 (N_2614,N_2083,N_1643);
nand U2615 (N_2615,N_1694,N_1844);
xor U2616 (N_2616,N_2309,N_2350);
nand U2617 (N_2617,N_1602,N_1933);
and U2618 (N_2618,N_1727,N_1929);
or U2619 (N_2619,N_2263,N_1676);
xor U2620 (N_2620,N_1661,N_2197);
and U2621 (N_2621,N_2037,N_2230);
xor U2622 (N_2622,N_2364,N_2149);
nand U2623 (N_2623,N_1677,N_2075);
nand U2624 (N_2624,N_2250,N_1772);
nand U2625 (N_2625,N_2285,N_2246);
xor U2626 (N_2626,N_1825,N_2398);
nor U2627 (N_2627,N_2302,N_1819);
nand U2628 (N_2628,N_1875,N_2247);
nand U2629 (N_2629,N_2052,N_1610);
and U2630 (N_2630,N_1611,N_1887);
nand U2631 (N_2631,N_2303,N_1870);
nor U2632 (N_2632,N_1601,N_1695);
or U2633 (N_2633,N_2226,N_1705);
or U2634 (N_2634,N_2305,N_2172);
or U2635 (N_2635,N_1900,N_1902);
and U2636 (N_2636,N_1915,N_1980);
xnor U2637 (N_2637,N_1806,N_1854);
nor U2638 (N_2638,N_2101,N_2343);
nor U2639 (N_2639,N_2125,N_1658);
and U2640 (N_2640,N_1952,N_1692);
xnor U2641 (N_2641,N_2163,N_2317);
nand U2642 (N_2642,N_1703,N_2352);
or U2643 (N_2643,N_2387,N_2170);
or U2644 (N_2644,N_1941,N_2169);
nor U2645 (N_2645,N_1737,N_2287);
or U2646 (N_2646,N_1609,N_1827);
or U2647 (N_2647,N_1860,N_1921);
xor U2648 (N_2648,N_2056,N_2154);
xor U2649 (N_2649,N_2103,N_2323);
nand U2650 (N_2650,N_1620,N_1659);
and U2651 (N_2651,N_2234,N_1704);
xnor U2652 (N_2652,N_2374,N_2209);
or U2653 (N_2653,N_1761,N_2200);
nor U2654 (N_2654,N_1809,N_1842);
nor U2655 (N_2655,N_2241,N_2019);
or U2656 (N_2656,N_2053,N_1607);
and U2657 (N_2657,N_1874,N_1606);
or U2658 (N_2658,N_2046,N_1969);
nor U2659 (N_2659,N_1886,N_2235);
xnor U2660 (N_2660,N_2345,N_1994);
xnor U2661 (N_2661,N_1846,N_1618);
nand U2662 (N_2662,N_2389,N_1813);
and U2663 (N_2663,N_1838,N_1738);
nor U2664 (N_2664,N_2143,N_1883);
nand U2665 (N_2665,N_2288,N_2198);
or U2666 (N_2666,N_2168,N_2070);
nor U2667 (N_2667,N_1764,N_1669);
nor U2668 (N_2668,N_2340,N_2094);
nor U2669 (N_2669,N_1935,N_2215);
nor U2670 (N_2670,N_2160,N_2378);
xor U2671 (N_2671,N_1760,N_1788);
xnor U2672 (N_2672,N_2204,N_2105);
nor U2673 (N_2673,N_1755,N_2258);
and U2674 (N_2674,N_1655,N_1988);
nor U2675 (N_2675,N_2119,N_1758);
nand U2676 (N_2676,N_1861,N_1729);
xnor U2677 (N_2677,N_2134,N_2082);
nand U2678 (N_2678,N_2396,N_2187);
and U2679 (N_2679,N_1763,N_1923);
and U2680 (N_2680,N_2185,N_1603);
and U2681 (N_2681,N_1907,N_1893);
nor U2682 (N_2682,N_2244,N_1639);
or U2683 (N_2683,N_2289,N_2017);
xnor U2684 (N_2684,N_2318,N_1653);
or U2685 (N_2685,N_1752,N_1831);
nor U2686 (N_2686,N_2106,N_1766);
or U2687 (N_2687,N_2254,N_1670);
or U2688 (N_2688,N_2089,N_1970);
nor U2689 (N_2689,N_1638,N_1757);
and U2690 (N_2690,N_2174,N_2310);
nand U2691 (N_2691,N_1776,N_2282);
nand U2692 (N_2692,N_2207,N_1621);
nor U2693 (N_2693,N_1662,N_2212);
nor U2694 (N_2694,N_2316,N_2380);
and U2695 (N_2695,N_2018,N_2262);
or U2696 (N_2696,N_2078,N_1756);
nor U2697 (N_2697,N_1957,N_1647);
nand U2698 (N_2698,N_1626,N_1682);
and U2699 (N_2699,N_2388,N_1852);
nor U2700 (N_2700,N_1800,N_2121);
or U2701 (N_2701,N_1868,N_2032);
and U2702 (N_2702,N_1981,N_1953);
and U2703 (N_2703,N_2151,N_1967);
xnor U2704 (N_2704,N_1914,N_2027);
xnor U2705 (N_2705,N_2011,N_1668);
and U2706 (N_2706,N_1691,N_1845);
or U2707 (N_2707,N_2098,N_2362);
nor U2708 (N_2708,N_2164,N_1747);
nor U2709 (N_2709,N_2314,N_2339);
xnor U2710 (N_2710,N_2192,N_2344);
nand U2711 (N_2711,N_2031,N_2260);
nand U2712 (N_2712,N_2311,N_1629);
xnor U2713 (N_2713,N_2320,N_2349);
nand U2714 (N_2714,N_2088,N_1759);
and U2715 (N_2715,N_1617,N_1808);
nand U2716 (N_2716,N_1794,N_1873);
nand U2717 (N_2717,N_1824,N_1946);
or U2718 (N_2718,N_1986,N_1992);
xor U2719 (N_2719,N_2148,N_2295);
nand U2720 (N_2720,N_1797,N_1722);
and U2721 (N_2721,N_1841,N_1635);
xor U2722 (N_2722,N_2181,N_2158);
or U2723 (N_2723,N_1908,N_2044);
nand U2724 (N_2724,N_2228,N_2057);
nor U2725 (N_2725,N_1802,N_1632);
xor U2726 (N_2726,N_2069,N_1631);
or U2727 (N_2727,N_1884,N_2024);
nor U2728 (N_2728,N_1839,N_2298);
nor U2729 (N_2729,N_1777,N_1665);
xor U2730 (N_2730,N_2248,N_2372);
xor U2731 (N_2731,N_2395,N_1832);
and U2732 (N_2732,N_2240,N_2021);
or U2733 (N_2733,N_1686,N_2131);
xnor U2734 (N_2734,N_1749,N_2129);
xnor U2735 (N_2735,N_2283,N_2117);
nand U2736 (N_2736,N_2290,N_1826);
and U2737 (N_2737,N_2267,N_2124);
nand U2738 (N_2738,N_1688,N_1926);
nor U2739 (N_2739,N_2243,N_1723);
and U2740 (N_2740,N_1863,N_1614);
nor U2741 (N_2741,N_1789,N_1849);
or U2742 (N_2742,N_1673,N_1917);
xor U2743 (N_2743,N_2348,N_2133);
or U2744 (N_2744,N_1608,N_1828);
nand U2745 (N_2745,N_2224,N_2366);
and U2746 (N_2746,N_2086,N_2325);
nand U2747 (N_2747,N_1615,N_2060);
or U2748 (N_2748,N_1899,N_2334);
and U2749 (N_2749,N_2249,N_1951);
xnor U2750 (N_2750,N_2330,N_1901);
and U2751 (N_2751,N_1767,N_1945);
or U2752 (N_2752,N_2223,N_1913);
xor U2753 (N_2753,N_2136,N_1739);
nor U2754 (N_2754,N_2381,N_1909);
and U2755 (N_2755,N_1746,N_1684);
xnor U2756 (N_2756,N_2342,N_1787);
and U2757 (N_2757,N_1830,N_1745);
and U2758 (N_2758,N_2231,N_1889);
nand U2759 (N_2759,N_2039,N_1920);
nand U2760 (N_2760,N_2077,N_2109);
xnor U2761 (N_2761,N_1829,N_1801);
nor U2762 (N_2762,N_2023,N_2202);
nand U2763 (N_2763,N_2040,N_2190);
and U2764 (N_2764,N_1778,N_1656);
and U2765 (N_2765,N_1648,N_2219);
and U2766 (N_2766,N_1701,N_2113);
nand U2767 (N_2767,N_2157,N_2229);
xnor U2768 (N_2768,N_1799,N_1931);
xor U2769 (N_2769,N_2211,N_1804);
xor U2770 (N_2770,N_2271,N_1707);
nor U2771 (N_2771,N_2093,N_2222);
or U2772 (N_2772,N_2043,N_1683);
xor U2773 (N_2773,N_2365,N_1654);
nor U2774 (N_2774,N_2291,N_2347);
xnor U2775 (N_2775,N_2013,N_1903);
nand U2776 (N_2776,N_1812,N_1744);
nor U2777 (N_2777,N_1753,N_2029);
xor U2778 (N_2778,N_2104,N_2319);
xor U2779 (N_2779,N_2099,N_1641);
nand U2780 (N_2780,N_1651,N_2049);
nor U2781 (N_2781,N_1876,N_1690);
xor U2782 (N_2782,N_2217,N_2294);
xor U2783 (N_2783,N_2383,N_2155);
or U2784 (N_2784,N_2341,N_2265);
and U2785 (N_2785,N_2337,N_1716);
nor U2786 (N_2786,N_1958,N_2081);
or U2787 (N_2787,N_2178,N_1754);
or U2788 (N_2788,N_1894,N_2281);
nor U2789 (N_2789,N_1636,N_1993);
and U2790 (N_2790,N_2390,N_1840);
nand U2791 (N_2791,N_1664,N_1771);
xnor U2792 (N_2792,N_1817,N_1633);
xnor U2793 (N_2793,N_1972,N_2153);
and U2794 (N_2794,N_2165,N_1735);
nand U2795 (N_2795,N_1864,N_1859);
xnor U2796 (N_2796,N_2090,N_1627);
or U2797 (N_2797,N_1645,N_1783);
nor U2798 (N_2798,N_2062,N_1918);
xnor U2799 (N_2799,N_2008,N_2328);
and U2800 (N_2800,N_2068,N_1869);
or U2801 (N_2801,N_1996,N_2339);
or U2802 (N_2802,N_2365,N_2376);
nor U2803 (N_2803,N_2034,N_1785);
xor U2804 (N_2804,N_2255,N_1985);
nand U2805 (N_2805,N_2015,N_1620);
xnor U2806 (N_2806,N_2370,N_1930);
nand U2807 (N_2807,N_1708,N_1924);
nand U2808 (N_2808,N_1910,N_2096);
and U2809 (N_2809,N_2322,N_2041);
nor U2810 (N_2810,N_2140,N_1818);
xor U2811 (N_2811,N_2033,N_1768);
nand U2812 (N_2812,N_1964,N_2178);
and U2813 (N_2813,N_1755,N_1952);
xor U2814 (N_2814,N_2384,N_2207);
or U2815 (N_2815,N_2346,N_1751);
xnor U2816 (N_2816,N_2255,N_2288);
xnor U2817 (N_2817,N_2083,N_1768);
xnor U2818 (N_2818,N_1653,N_2163);
nor U2819 (N_2819,N_1849,N_1745);
or U2820 (N_2820,N_1891,N_1634);
nor U2821 (N_2821,N_1908,N_1985);
xor U2822 (N_2822,N_1993,N_2079);
nand U2823 (N_2823,N_2265,N_2385);
or U2824 (N_2824,N_2275,N_1761);
and U2825 (N_2825,N_1861,N_2173);
xnor U2826 (N_2826,N_1821,N_1701);
xor U2827 (N_2827,N_2100,N_1752);
nand U2828 (N_2828,N_1893,N_1953);
xnor U2829 (N_2829,N_2358,N_2069);
xnor U2830 (N_2830,N_1708,N_2397);
xnor U2831 (N_2831,N_2033,N_2389);
nand U2832 (N_2832,N_2073,N_1966);
and U2833 (N_2833,N_2338,N_1958);
and U2834 (N_2834,N_2014,N_2373);
nand U2835 (N_2835,N_2302,N_1768);
xnor U2836 (N_2836,N_1920,N_2205);
xor U2837 (N_2837,N_2074,N_1740);
nand U2838 (N_2838,N_1642,N_2329);
or U2839 (N_2839,N_2086,N_1717);
nor U2840 (N_2840,N_1897,N_1952);
and U2841 (N_2841,N_2077,N_1886);
xor U2842 (N_2842,N_1783,N_2276);
xor U2843 (N_2843,N_1813,N_1966);
xor U2844 (N_2844,N_1693,N_1871);
nand U2845 (N_2845,N_2240,N_1814);
xnor U2846 (N_2846,N_2378,N_1616);
nor U2847 (N_2847,N_2002,N_2037);
nor U2848 (N_2848,N_1817,N_1959);
or U2849 (N_2849,N_2105,N_1787);
nand U2850 (N_2850,N_1621,N_2181);
nor U2851 (N_2851,N_1770,N_1649);
nand U2852 (N_2852,N_2391,N_2005);
nor U2853 (N_2853,N_1603,N_1878);
nor U2854 (N_2854,N_2226,N_1827);
or U2855 (N_2855,N_2011,N_1971);
nor U2856 (N_2856,N_1896,N_1932);
nor U2857 (N_2857,N_1720,N_2331);
and U2858 (N_2858,N_1899,N_2043);
nand U2859 (N_2859,N_2133,N_1940);
xnor U2860 (N_2860,N_1890,N_1913);
xnor U2861 (N_2861,N_1741,N_1754);
nand U2862 (N_2862,N_2307,N_2191);
nand U2863 (N_2863,N_2276,N_2237);
nor U2864 (N_2864,N_1890,N_1740);
and U2865 (N_2865,N_1706,N_1814);
nand U2866 (N_2866,N_2306,N_2079);
xnor U2867 (N_2867,N_1953,N_2233);
nor U2868 (N_2868,N_1728,N_1811);
nand U2869 (N_2869,N_1767,N_2175);
xnor U2870 (N_2870,N_2253,N_2293);
or U2871 (N_2871,N_1896,N_2019);
nor U2872 (N_2872,N_2105,N_1864);
nand U2873 (N_2873,N_1673,N_2364);
nor U2874 (N_2874,N_2135,N_1871);
xnor U2875 (N_2875,N_1934,N_1855);
xnor U2876 (N_2876,N_1926,N_1832);
and U2877 (N_2877,N_2160,N_1700);
xnor U2878 (N_2878,N_2046,N_2027);
xor U2879 (N_2879,N_2212,N_1970);
and U2880 (N_2880,N_2033,N_1602);
and U2881 (N_2881,N_2322,N_1617);
and U2882 (N_2882,N_2265,N_1860);
nor U2883 (N_2883,N_1965,N_2095);
nand U2884 (N_2884,N_2302,N_2109);
and U2885 (N_2885,N_2005,N_2240);
and U2886 (N_2886,N_2050,N_2285);
nand U2887 (N_2887,N_2012,N_2142);
or U2888 (N_2888,N_2212,N_1791);
nand U2889 (N_2889,N_1968,N_2381);
xor U2890 (N_2890,N_2003,N_1785);
xor U2891 (N_2891,N_1731,N_1965);
or U2892 (N_2892,N_1947,N_1765);
nor U2893 (N_2893,N_1729,N_2140);
xor U2894 (N_2894,N_1854,N_2012);
and U2895 (N_2895,N_1653,N_2208);
and U2896 (N_2896,N_2328,N_2254);
nor U2897 (N_2897,N_2223,N_1839);
xor U2898 (N_2898,N_1969,N_2150);
nor U2899 (N_2899,N_1917,N_1939);
nor U2900 (N_2900,N_2272,N_2071);
xor U2901 (N_2901,N_1809,N_1623);
or U2902 (N_2902,N_1884,N_2055);
nand U2903 (N_2903,N_2389,N_1860);
xor U2904 (N_2904,N_2024,N_1609);
and U2905 (N_2905,N_2151,N_2098);
and U2906 (N_2906,N_2296,N_1842);
nand U2907 (N_2907,N_2290,N_2317);
xnor U2908 (N_2908,N_1873,N_1742);
and U2909 (N_2909,N_2013,N_2007);
or U2910 (N_2910,N_2334,N_1858);
nand U2911 (N_2911,N_2024,N_1694);
nand U2912 (N_2912,N_1829,N_1950);
xnor U2913 (N_2913,N_1976,N_1773);
nand U2914 (N_2914,N_2181,N_1996);
xnor U2915 (N_2915,N_1705,N_1810);
and U2916 (N_2916,N_1740,N_2207);
nand U2917 (N_2917,N_2259,N_2292);
or U2918 (N_2918,N_1677,N_2396);
xor U2919 (N_2919,N_2389,N_2004);
nor U2920 (N_2920,N_1929,N_1687);
xor U2921 (N_2921,N_2177,N_2028);
xor U2922 (N_2922,N_2287,N_2032);
nand U2923 (N_2923,N_2125,N_2266);
nor U2924 (N_2924,N_2159,N_2328);
xor U2925 (N_2925,N_1753,N_1797);
and U2926 (N_2926,N_2208,N_2115);
nand U2927 (N_2927,N_1787,N_1661);
or U2928 (N_2928,N_2366,N_1828);
or U2929 (N_2929,N_1618,N_2273);
or U2930 (N_2930,N_1723,N_2170);
and U2931 (N_2931,N_2292,N_2089);
nor U2932 (N_2932,N_1995,N_1862);
nand U2933 (N_2933,N_2018,N_2033);
and U2934 (N_2934,N_2203,N_2244);
and U2935 (N_2935,N_1841,N_1849);
nor U2936 (N_2936,N_2324,N_2348);
nor U2937 (N_2937,N_2380,N_2183);
or U2938 (N_2938,N_1622,N_1645);
xnor U2939 (N_2939,N_1881,N_1900);
xor U2940 (N_2940,N_1639,N_2378);
nor U2941 (N_2941,N_2139,N_1617);
nand U2942 (N_2942,N_2133,N_2398);
xnor U2943 (N_2943,N_2268,N_1886);
and U2944 (N_2944,N_1848,N_2153);
or U2945 (N_2945,N_1707,N_2121);
xor U2946 (N_2946,N_1608,N_1948);
and U2947 (N_2947,N_2269,N_1625);
nand U2948 (N_2948,N_1904,N_2075);
nor U2949 (N_2949,N_2126,N_1792);
or U2950 (N_2950,N_1936,N_2238);
nand U2951 (N_2951,N_1628,N_2240);
and U2952 (N_2952,N_2096,N_2172);
nand U2953 (N_2953,N_1712,N_1687);
nand U2954 (N_2954,N_2018,N_1788);
or U2955 (N_2955,N_2216,N_2382);
nor U2956 (N_2956,N_1633,N_1741);
nor U2957 (N_2957,N_1751,N_1773);
nor U2958 (N_2958,N_1967,N_2122);
and U2959 (N_2959,N_2296,N_1616);
xor U2960 (N_2960,N_2217,N_1821);
xnor U2961 (N_2961,N_2344,N_1607);
nor U2962 (N_2962,N_2211,N_2087);
nor U2963 (N_2963,N_2228,N_2010);
and U2964 (N_2964,N_2192,N_1891);
or U2965 (N_2965,N_2025,N_1920);
nand U2966 (N_2966,N_1759,N_1981);
or U2967 (N_2967,N_2025,N_1905);
xnor U2968 (N_2968,N_1661,N_1959);
nor U2969 (N_2969,N_1829,N_2054);
and U2970 (N_2970,N_1973,N_1672);
xor U2971 (N_2971,N_1669,N_1818);
xor U2972 (N_2972,N_1631,N_2126);
xor U2973 (N_2973,N_1725,N_2264);
nand U2974 (N_2974,N_1666,N_2211);
xor U2975 (N_2975,N_1793,N_1671);
nand U2976 (N_2976,N_1986,N_1750);
or U2977 (N_2977,N_2253,N_1805);
or U2978 (N_2978,N_2123,N_1885);
and U2979 (N_2979,N_1727,N_1723);
xnor U2980 (N_2980,N_1760,N_1684);
and U2981 (N_2981,N_1779,N_2316);
nand U2982 (N_2982,N_1833,N_2154);
xnor U2983 (N_2983,N_1986,N_1803);
and U2984 (N_2984,N_1631,N_2243);
xor U2985 (N_2985,N_1927,N_1674);
nand U2986 (N_2986,N_2253,N_2121);
xor U2987 (N_2987,N_1649,N_2342);
or U2988 (N_2988,N_1686,N_1953);
xor U2989 (N_2989,N_1857,N_1736);
xnor U2990 (N_2990,N_2131,N_1902);
and U2991 (N_2991,N_2280,N_1816);
or U2992 (N_2992,N_2125,N_1888);
nand U2993 (N_2993,N_1696,N_2241);
and U2994 (N_2994,N_1718,N_2262);
nand U2995 (N_2995,N_2350,N_2192);
or U2996 (N_2996,N_2377,N_2363);
and U2997 (N_2997,N_1887,N_1908);
or U2998 (N_2998,N_1667,N_1781);
and U2999 (N_2999,N_2243,N_1860);
nand U3000 (N_3000,N_2289,N_1782);
xnor U3001 (N_3001,N_2024,N_2173);
nand U3002 (N_3002,N_1887,N_2023);
nor U3003 (N_3003,N_2175,N_1916);
and U3004 (N_3004,N_2199,N_1932);
or U3005 (N_3005,N_2009,N_2303);
or U3006 (N_3006,N_2238,N_1911);
nand U3007 (N_3007,N_1758,N_1759);
xor U3008 (N_3008,N_1645,N_2066);
or U3009 (N_3009,N_1748,N_2335);
nor U3010 (N_3010,N_2232,N_1893);
and U3011 (N_3011,N_2170,N_2092);
xor U3012 (N_3012,N_2282,N_1619);
xor U3013 (N_3013,N_1949,N_1948);
xor U3014 (N_3014,N_1980,N_1928);
xnor U3015 (N_3015,N_1958,N_1816);
xor U3016 (N_3016,N_2364,N_1988);
or U3017 (N_3017,N_2267,N_2023);
nor U3018 (N_3018,N_1823,N_1609);
or U3019 (N_3019,N_1685,N_2300);
and U3020 (N_3020,N_1650,N_2058);
xnor U3021 (N_3021,N_1651,N_2051);
nand U3022 (N_3022,N_2383,N_1861);
and U3023 (N_3023,N_1844,N_1695);
or U3024 (N_3024,N_1905,N_2065);
nor U3025 (N_3025,N_1908,N_1638);
nor U3026 (N_3026,N_2054,N_2274);
or U3027 (N_3027,N_1970,N_2072);
xor U3028 (N_3028,N_1977,N_2255);
and U3029 (N_3029,N_1665,N_2005);
nand U3030 (N_3030,N_2018,N_1826);
xor U3031 (N_3031,N_1692,N_1795);
nand U3032 (N_3032,N_2098,N_2361);
or U3033 (N_3033,N_2254,N_2307);
nor U3034 (N_3034,N_2387,N_2081);
and U3035 (N_3035,N_2228,N_2244);
xnor U3036 (N_3036,N_1886,N_1648);
nand U3037 (N_3037,N_2259,N_1983);
nand U3038 (N_3038,N_2073,N_2176);
nor U3039 (N_3039,N_2394,N_1701);
or U3040 (N_3040,N_1896,N_1653);
nand U3041 (N_3041,N_2147,N_1864);
and U3042 (N_3042,N_1703,N_2038);
xor U3043 (N_3043,N_2292,N_2140);
or U3044 (N_3044,N_1872,N_1835);
or U3045 (N_3045,N_1633,N_2310);
and U3046 (N_3046,N_2098,N_2114);
or U3047 (N_3047,N_1858,N_2093);
xor U3048 (N_3048,N_1785,N_2246);
and U3049 (N_3049,N_1824,N_1776);
nor U3050 (N_3050,N_2350,N_2050);
nand U3051 (N_3051,N_1758,N_2104);
nand U3052 (N_3052,N_1909,N_1923);
xor U3053 (N_3053,N_1986,N_2398);
nand U3054 (N_3054,N_1946,N_2102);
or U3055 (N_3055,N_1907,N_1706);
nor U3056 (N_3056,N_2039,N_1737);
or U3057 (N_3057,N_1900,N_2047);
or U3058 (N_3058,N_1656,N_1987);
xor U3059 (N_3059,N_1988,N_2143);
nand U3060 (N_3060,N_1721,N_1857);
nor U3061 (N_3061,N_1767,N_2191);
nand U3062 (N_3062,N_2277,N_1974);
nor U3063 (N_3063,N_1998,N_2063);
and U3064 (N_3064,N_1925,N_2167);
or U3065 (N_3065,N_1798,N_2261);
and U3066 (N_3066,N_1762,N_2040);
or U3067 (N_3067,N_2249,N_1730);
or U3068 (N_3068,N_2286,N_1820);
nand U3069 (N_3069,N_2243,N_2051);
and U3070 (N_3070,N_2226,N_2129);
and U3071 (N_3071,N_2149,N_2243);
nor U3072 (N_3072,N_1788,N_1804);
and U3073 (N_3073,N_1920,N_2096);
xnor U3074 (N_3074,N_2269,N_1615);
nand U3075 (N_3075,N_1888,N_2130);
xnor U3076 (N_3076,N_1873,N_2119);
nor U3077 (N_3077,N_1611,N_1815);
or U3078 (N_3078,N_1600,N_2153);
nand U3079 (N_3079,N_2355,N_1993);
or U3080 (N_3080,N_2283,N_2293);
nor U3081 (N_3081,N_2043,N_2258);
or U3082 (N_3082,N_2351,N_2193);
or U3083 (N_3083,N_1650,N_2267);
and U3084 (N_3084,N_1922,N_1849);
nor U3085 (N_3085,N_2125,N_2066);
or U3086 (N_3086,N_1959,N_2084);
nand U3087 (N_3087,N_1719,N_2073);
nand U3088 (N_3088,N_2162,N_1978);
or U3089 (N_3089,N_2186,N_2142);
and U3090 (N_3090,N_2240,N_2036);
nor U3091 (N_3091,N_2016,N_1838);
and U3092 (N_3092,N_2241,N_2032);
nand U3093 (N_3093,N_1761,N_1713);
or U3094 (N_3094,N_2303,N_1813);
nor U3095 (N_3095,N_2031,N_1990);
nand U3096 (N_3096,N_1811,N_2016);
and U3097 (N_3097,N_1782,N_2237);
or U3098 (N_3098,N_1663,N_2046);
and U3099 (N_3099,N_1652,N_2040);
nor U3100 (N_3100,N_1637,N_2141);
and U3101 (N_3101,N_1812,N_1927);
nand U3102 (N_3102,N_2223,N_1806);
or U3103 (N_3103,N_1613,N_1687);
xnor U3104 (N_3104,N_2243,N_2113);
or U3105 (N_3105,N_1866,N_2214);
and U3106 (N_3106,N_1812,N_2337);
or U3107 (N_3107,N_1723,N_1708);
xor U3108 (N_3108,N_1873,N_1733);
or U3109 (N_3109,N_1783,N_1960);
nand U3110 (N_3110,N_2137,N_1913);
and U3111 (N_3111,N_2394,N_1828);
nand U3112 (N_3112,N_2353,N_1887);
xor U3113 (N_3113,N_2388,N_1918);
xnor U3114 (N_3114,N_2314,N_1841);
xnor U3115 (N_3115,N_2373,N_2229);
and U3116 (N_3116,N_1903,N_1712);
nor U3117 (N_3117,N_2323,N_2311);
and U3118 (N_3118,N_1906,N_2294);
nor U3119 (N_3119,N_1953,N_1903);
nand U3120 (N_3120,N_2018,N_1880);
and U3121 (N_3121,N_2255,N_1912);
nor U3122 (N_3122,N_1994,N_2283);
and U3123 (N_3123,N_2189,N_1965);
or U3124 (N_3124,N_2301,N_1646);
xor U3125 (N_3125,N_1899,N_2278);
xor U3126 (N_3126,N_2196,N_2255);
or U3127 (N_3127,N_1831,N_2219);
nor U3128 (N_3128,N_2119,N_1699);
or U3129 (N_3129,N_2151,N_2103);
xor U3130 (N_3130,N_2212,N_2292);
nand U3131 (N_3131,N_1628,N_2060);
xnor U3132 (N_3132,N_2034,N_2115);
xor U3133 (N_3133,N_1629,N_1846);
and U3134 (N_3134,N_2079,N_2055);
and U3135 (N_3135,N_2396,N_1813);
nor U3136 (N_3136,N_1988,N_1950);
or U3137 (N_3137,N_1946,N_2369);
xnor U3138 (N_3138,N_2118,N_2234);
nand U3139 (N_3139,N_1794,N_2399);
or U3140 (N_3140,N_1895,N_1918);
and U3141 (N_3141,N_1706,N_2042);
or U3142 (N_3142,N_2070,N_2238);
or U3143 (N_3143,N_1755,N_1906);
nor U3144 (N_3144,N_2317,N_1701);
and U3145 (N_3145,N_2129,N_1897);
xnor U3146 (N_3146,N_1912,N_2208);
nor U3147 (N_3147,N_2157,N_2356);
or U3148 (N_3148,N_1990,N_2067);
nor U3149 (N_3149,N_2339,N_1800);
xnor U3150 (N_3150,N_2129,N_2231);
nand U3151 (N_3151,N_1662,N_1703);
nor U3152 (N_3152,N_1905,N_2066);
xor U3153 (N_3153,N_1697,N_1972);
or U3154 (N_3154,N_1971,N_1693);
or U3155 (N_3155,N_2004,N_1854);
nor U3156 (N_3156,N_2295,N_1802);
and U3157 (N_3157,N_2357,N_1607);
nand U3158 (N_3158,N_2393,N_2331);
nor U3159 (N_3159,N_2067,N_2109);
xor U3160 (N_3160,N_1776,N_1941);
nor U3161 (N_3161,N_1753,N_2033);
and U3162 (N_3162,N_2326,N_2014);
or U3163 (N_3163,N_1603,N_2091);
nor U3164 (N_3164,N_1827,N_2353);
nand U3165 (N_3165,N_2144,N_2167);
xnor U3166 (N_3166,N_2300,N_2157);
nand U3167 (N_3167,N_1860,N_1866);
or U3168 (N_3168,N_1943,N_2287);
nor U3169 (N_3169,N_2165,N_2355);
xor U3170 (N_3170,N_2008,N_1966);
nor U3171 (N_3171,N_1625,N_1991);
or U3172 (N_3172,N_1833,N_1974);
or U3173 (N_3173,N_2389,N_2306);
and U3174 (N_3174,N_1924,N_1902);
or U3175 (N_3175,N_1734,N_2190);
and U3176 (N_3176,N_2280,N_2232);
nor U3177 (N_3177,N_2266,N_1616);
xor U3178 (N_3178,N_2063,N_1629);
nor U3179 (N_3179,N_1865,N_1660);
xnor U3180 (N_3180,N_2099,N_2229);
xor U3181 (N_3181,N_2176,N_1888);
xnor U3182 (N_3182,N_2277,N_1985);
xor U3183 (N_3183,N_1875,N_2100);
and U3184 (N_3184,N_2305,N_1685);
nor U3185 (N_3185,N_2077,N_1632);
xnor U3186 (N_3186,N_1620,N_1909);
nand U3187 (N_3187,N_2124,N_1676);
xnor U3188 (N_3188,N_1623,N_2051);
nor U3189 (N_3189,N_2391,N_1913);
nand U3190 (N_3190,N_2146,N_1891);
and U3191 (N_3191,N_2152,N_2346);
nor U3192 (N_3192,N_1947,N_1633);
or U3193 (N_3193,N_2354,N_1982);
nand U3194 (N_3194,N_1938,N_1869);
nand U3195 (N_3195,N_1889,N_2308);
nor U3196 (N_3196,N_2160,N_2105);
or U3197 (N_3197,N_2024,N_1710);
xor U3198 (N_3198,N_1600,N_2117);
and U3199 (N_3199,N_2274,N_1608);
and U3200 (N_3200,N_2400,N_2645);
and U3201 (N_3201,N_2833,N_2585);
or U3202 (N_3202,N_2934,N_3022);
xnor U3203 (N_3203,N_2623,N_2790);
xnor U3204 (N_3204,N_2892,N_2868);
nand U3205 (N_3205,N_2759,N_3141);
and U3206 (N_3206,N_2574,N_2722);
nor U3207 (N_3207,N_2787,N_2888);
and U3208 (N_3208,N_2429,N_2473);
or U3209 (N_3209,N_3082,N_2606);
xor U3210 (N_3210,N_2988,N_2878);
and U3211 (N_3211,N_2747,N_2426);
or U3212 (N_3212,N_2758,N_2992);
and U3213 (N_3213,N_2660,N_2766);
nor U3214 (N_3214,N_2693,N_2717);
or U3215 (N_3215,N_2430,N_3077);
and U3216 (N_3216,N_2857,N_2972);
nor U3217 (N_3217,N_2948,N_2534);
or U3218 (N_3218,N_3063,N_3161);
and U3219 (N_3219,N_2586,N_2742);
xor U3220 (N_3220,N_2712,N_2437);
xnor U3221 (N_3221,N_2726,N_2520);
and U3222 (N_3222,N_2821,N_2450);
nor U3223 (N_3223,N_2565,N_3016);
xor U3224 (N_3224,N_2556,N_2605);
and U3225 (N_3225,N_2910,N_3159);
xor U3226 (N_3226,N_2728,N_2570);
or U3227 (N_3227,N_3126,N_2705);
nand U3228 (N_3228,N_3131,N_3052);
nor U3229 (N_3229,N_2763,N_2691);
and U3230 (N_3230,N_3195,N_2996);
xor U3231 (N_3231,N_2649,N_2692);
and U3232 (N_3232,N_2466,N_2876);
and U3233 (N_3233,N_2420,N_3080);
nor U3234 (N_3234,N_2672,N_2635);
nand U3235 (N_3235,N_2898,N_2869);
and U3236 (N_3236,N_2681,N_2659);
nor U3237 (N_3237,N_2922,N_2564);
and U3238 (N_3238,N_2666,N_3041);
and U3239 (N_3239,N_2818,N_3044);
or U3240 (N_3240,N_2637,N_2825);
nand U3241 (N_3241,N_2680,N_3054);
nor U3242 (N_3242,N_3111,N_2950);
xnor U3243 (N_3243,N_2760,N_2675);
or U3244 (N_3244,N_2983,N_3134);
and U3245 (N_3245,N_2456,N_2514);
xnor U3246 (N_3246,N_2719,N_2715);
nor U3247 (N_3247,N_2573,N_3129);
nand U3248 (N_3248,N_2735,N_2871);
nor U3249 (N_3249,N_2801,N_2986);
or U3250 (N_3250,N_3119,N_2686);
and U3251 (N_3251,N_2872,N_2751);
nor U3252 (N_3252,N_2985,N_2485);
nand U3253 (N_3253,N_3187,N_2729);
nor U3254 (N_3254,N_2723,N_3081);
xor U3255 (N_3255,N_2946,N_2633);
nor U3256 (N_3256,N_3028,N_3116);
xor U3257 (N_3257,N_2906,N_2689);
nor U3258 (N_3258,N_2832,N_3047);
or U3259 (N_3259,N_2651,N_2867);
or U3260 (N_3260,N_3132,N_2447);
xnor U3261 (N_3261,N_2549,N_2834);
and U3262 (N_3262,N_3051,N_2609);
nor U3263 (N_3263,N_2552,N_2939);
nor U3264 (N_3264,N_2600,N_2638);
nor U3265 (N_3265,N_2575,N_3033);
or U3266 (N_3266,N_2612,N_2583);
and U3267 (N_3267,N_2817,N_2930);
and U3268 (N_3268,N_3065,N_2954);
nor U3269 (N_3269,N_2924,N_2940);
and U3270 (N_3270,N_2589,N_3146);
nand U3271 (N_3271,N_3196,N_3027);
nand U3272 (N_3272,N_2483,N_3074);
nor U3273 (N_3273,N_2548,N_2537);
nor U3274 (N_3274,N_2541,N_2463);
nand U3275 (N_3275,N_3173,N_2475);
xnor U3276 (N_3276,N_2554,N_2713);
and U3277 (N_3277,N_3114,N_2653);
or U3278 (N_3278,N_2655,N_3160);
xor U3279 (N_3279,N_2776,N_3099);
xnor U3280 (N_3280,N_2404,N_2740);
nand U3281 (N_3281,N_2524,N_2797);
xor U3282 (N_3282,N_2671,N_2622);
nand U3283 (N_3283,N_2525,N_3103);
and U3284 (N_3284,N_2995,N_3130);
xnor U3285 (N_3285,N_2733,N_2720);
xnor U3286 (N_3286,N_2700,N_2603);
nor U3287 (N_3287,N_3009,N_2829);
nand U3288 (N_3288,N_2804,N_3157);
nand U3289 (N_3289,N_2506,N_3006);
nor U3290 (N_3290,N_2739,N_2464);
or U3291 (N_3291,N_3172,N_2521);
nand U3292 (N_3292,N_2936,N_3045);
and U3293 (N_3293,N_2807,N_3058);
nor U3294 (N_3294,N_3198,N_3192);
nor U3295 (N_3295,N_2941,N_3064);
and U3296 (N_3296,N_3073,N_2440);
and U3297 (N_3297,N_3088,N_2744);
and U3298 (N_3298,N_2643,N_3057);
and U3299 (N_3299,N_3112,N_2488);
xor U3300 (N_3300,N_2417,N_3068);
nor U3301 (N_3301,N_2442,N_2628);
and U3302 (N_3302,N_3003,N_2592);
and U3303 (N_3303,N_2767,N_2885);
xnor U3304 (N_3304,N_2811,N_3005);
nand U3305 (N_3305,N_2487,N_2779);
nand U3306 (N_3306,N_2793,N_3169);
xor U3307 (N_3307,N_3098,N_2916);
xor U3308 (N_3308,N_3136,N_2654);
nand U3309 (N_3309,N_2962,N_2854);
and U3310 (N_3310,N_2597,N_2462);
nor U3311 (N_3311,N_2757,N_2835);
and U3312 (N_3312,N_3153,N_2465);
nor U3313 (N_3313,N_2555,N_2993);
xnor U3314 (N_3314,N_2676,N_3007);
nand U3315 (N_3315,N_2499,N_2738);
or U3316 (N_3316,N_3024,N_2734);
xor U3317 (N_3317,N_2975,N_2864);
or U3318 (N_3318,N_2953,N_3087);
xor U3319 (N_3319,N_2652,N_2781);
nor U3320 (N_3320,N_2667,N_2877);
nor U3321 (N_3321,N_2478,N_2926);
or U3322 (N_3322,N_2874,N_3182);
xnor U3323 (N_3323,N_2594,N_2412);
and U3324 (N_3324,N_2532,N_2517);
nand U3325 (N_3325,N_2852,N_3067);
or U3326 (N_3326,N_3036,N_2849);
and U3327 (N_3327,N_3122,N_2491);
xnor U3328 (N_3328,N_2631,N_2677);
nor U3329 (N_3329,N_2476,N_2904);
nand U3330 (N_3330,N_3037,N_2610);
nor U3331 (N_3331,N_2613,N_2572);
nand U3332 (N_3332,N_2981,N_2538);
nor U3333 (N_3333,N_2933,N_2596);
or U3334 (N_3334,N_3174,N_2887);
nand U3335 (N_3335,N_2706,N_2469);
xnor U3336 (N_3336,N_3050,N_2984);
or U3337 (N_3337,N_2855,N_3092);
xnor U3338 (N_3338,N_3101,N_2566);
or U3339 (N_3339,N_3177,N_2539);
and U3340 (N_3340,N_2644,N_2579);
or U3341 (N_3341,N_2727,N_2670);
nor U3342 (N_3342,N_2918,N_2703);
nor U3343 (N_3343,N_2567,N_2461);
xnor U3344 (N_3344,N_2937,N_2516);
xnor U3345 (N_3345,N_2749,N_2694);
or U3346 (N_3346,N_2646,N_2441);
nor U3347 (N_3347,N_2805,N_2658);
nor U3348 (N_3348,N_3110,N_2544);
nor U3349 (N_3349,N_3164,N_2990);
or U3350 (N_3350,N_3042,N_3113);
and U3351 (N_3351,N_2895,N_2477);
nand U3352 (N_3352,N_3061,N_2987);
and U3353 (N_3353,N_2828,N_2782);
and U3354 (N_3354,N_3185,N_2451);
and U3355 (N_3355,N_2630,N_2518);
nor U3356 (N_3356,N_2438,N_2908);
and U3357 (N_3357,N_2826,N_3035);
xor U3358 (N_3358,N_3143,N_2557);
xnor U3359 (N_3359,N_2927,N_3102);
nor U3360 (N_3360,N_2812,N_2648);
and U3361 (N_3361,N_2474,N_2695);
and U3362 (N_3362,N_2971,N_2863);
or U3363 (N_3363,N_3125,N_3107);
or U3364 (N_3364,N_2460,N_2495);
xor U3365 (N_3365,N_2591,N_2590);
and U3366 (N_3366,N_2748,N_2650);
xor U3367 (N_3367,N_2486,N_2913);
nor U3368 (N_3368,N_2900,N_2535);
or U3369 (N_3369,N_3180,N_2772);
xnor U3370 (N_3370,N_2861,N_2974);
nor U3371 (N_3371,N_2636,N_2455);
nor U3372 (N_3372,N_2813,N_2577);
or U3373 (N_3373,N_2907,N_2550);
or U3374 (N_3374,N_2512,N_2618);
nor U3375 (N_3375,N_2611,N_2444);
xnor U3376 (N_3376,N_2837,N_2911);
nor U3377 (N_3377,N_2568,N_2866);
nand U3378 (N_3378,N_2413,N_2870);
and U3379 (N_3379,N_2640,N_2980);
and U3380 (N_3380,N_2559,N_3013);
nand U3381 (N_3381,N_2416,N_2920);
and U3382 (N_3382,N_2580,N_3014);
nand U3383 (N_3383,N_3078,N_2736);
nor U3384 (N_3384,N_3175,N_2467);
or U3385 (N_3385,N_2800,N_2741);
nand U3386 (N_3386,N_2665,N_2489);
or U3387 (N_3387,N_3086,N_3097);
and U3388 (N_3388,N_2873,N_2448);
xor U3389 (N_3389,N_2824,N_2773);
and U3390 (N_3390,N_3123,N_2593);
nand U3391 (N_3391,N_2850,N_2875);
or U3392 (N_3392,N_2732,N_3090);
xor U3393 (N_3393,N_2998,N_2553);
xor U3394 (N_3394,N_2578,N_2699);
nor U3395 (N_3395,N_2507,N_2756);
nand U3396 (N_3396,N_2602,N_2752);
or U3397 (N_3397,N_2494,N_2959);
nor U3398 (N_3398,N_2961,N_2471);
nand U3399 (N_3399,N_2890,N_2533);
xnor U3400 (N_3400,N_2862,N_2625);
nand U3401 (N_3401,N_2967,N_2561);
xnor U3402 (N_3402,N_2409,N_3190);
xnor U3403 (N_3403,N_2770,N_3001);
xor U3404 (N_3404,N_2952,N_2966);
and U3405 (N_3405,N_2696,N_2428);
xor U3406 (N_3406,N_2608,N_2725);
nor U3407 (N_3407,N_2530,N_3032);
nor U3408 (N_3408,N_3019,N_2584);
nor U3409 (N_3409,N_3193,N_3165);
and U3410 (N_3410,N_3154,N_2619);
nand U3411 (N_3411,N_2702,N_2536);
nand U3412 (N_3412,N_2769,N_2528);
nor U3413 (N_3413,N_2902,N_2601);
xor U3414 (N_3414,N_2761,N_2576);
nor U3415 (N_3415,N_2803,N_2978);
xnor U3416 (N_3416,N_2755,N_3199);
nor U3417 (N_3417,N_2951,N_2663);
nand U3418 (N_3418,N_2841,N_2802);
and U3419 (N_3419,N_2458,N_3072);
or U3420 (N_3420,N_3023,N_2815);
and U3421 (N_3421,N_2647,N_3040);
xor U3422 (N_3422,N_3115,N_2546);
and U3423 (N_3423,N_3070,N_2673);
or U3424 (N_3424,N_2819,N_2683);
xor U3425 (N_3425,N_2958,N_3138);
and U3426 (N_3426,N_3139,N_3012);
or U3427 (N_3427,N_2964,N_2662);
nand U3428 (N_3428,N_3167,N_3176);
and U3429 (N_3429,N_2810,N_2994);
nand U3430 (N_3430,N_3091,N_2624);
nor U3431 (N_3431,N_2452,N_2799);
nor U3432 (N_3432,N_2840,N_3055);
nor U3433 (N_3433,N_3002,N_2500);
nand U3434 (N_3434,N_2796,N_2709);
xor U3435 (N_3435,N_2928,N_2856);
and U3436 (N_3436,N_2604,N_2425);
nor U3437 (N_3437,N_2432,N_2410);
xnor U3438 (N_3438,N_2436,N_2515);
and U3439 (N_3439,N_2714,N_3049);
nor U3440 (N_3440,N_2408,N_2415);
or U3441 (N_3441,N_2414,N_2925);
xor U3442 (N_3442,N_2457,N_2822);
nor U3443 (N_3443,N_2919,N_2778);
or U3444 (N_3444,N_2406,N_2831);
or U3445 (N_3445,N_3004,N_2771);
nor U3446 (N_3446,N_2588,N_2587);
xor U3447 (N_3447,N_2929,N_2991);
or U3448 (N_3448,N_2785,N_2669);
nor U3449 (N_3449,N_2762,N_3017);
or U3450 (N_3450,N_2982,N_2915);
xor U3451 (N_3451,N_2629,N_2768);
and U3452 (N_3452,N_3089,N_3120);
nand U3453 (N_3453,N_2627,N_2634);
and U3454 (N_3454,N_3043,N_2879);
nand U3455 (N_3455,N_2422,N_2439);
and U3456 (N_3456,N_2405,N_3093);
or U3457 (N_3457,N_2724,N_2433);
and U3458 (N_3458,N_3194,N_2968);
and U3459 (N_3459,N_3137,N_2780);
nand U3460 (N_3460,N_2632,N_2595);
or U3461 (N_3461,N_2938,N_3178);
and U3462 (N_3462,N_2884,N_2563);
nor U3463 (N_3463,N_2979,N_3000);
nor U3464 (N_3464,N_2505,N_2522);
or U3465 (N_3465,N_2783,N_3069);
and U3466 (N_3466,N_2529,N_2523);
nor U3467 (N_3467,N_2795,N_2775);
xor U3468 (N_3468,N_2730,N_3095);
nor U3469 (N_3469,N_2955,N_3179);
or U3470 (N_3470,N_2481,N_3039);
and U3471 (N_3471,N_2679,N_2468);
or U3472 (N_3472,N_2502,N_3150);
nor U3473 (N_3473,N_2582,N_2484);
xor U3474 (N_3474,N_2731,N_2657);
nor U3475 (N_3475,N_2710,N_2571);
nor U3476 (N_3476,N_3163,N_2949);
or U3477 (N_3477,N_2905,N_2668);
nand U3478 (N_3478,N_3025,N_2791);
xor U3479 (N_3479,N_2443,N_3166);
nand U3480 (N_3480,N_2880,N_2881);
or U3481 (N_3481,N_2688,N_3171);
nand U3482 (N_3482,N_3105,N_2501);
xnor U3483 (N_3483,N_2774,N_3162);
nand U3484 (N_3484,N_2743,N_2423);
nor U3485 (N_3485,N_2899,N_2737);
nor U3486 (N_3486,N_2449,N_3083);
or U3487 (N_3487,N_2997,N_2965);
or U3488 (N_3488,N_2847,N_2656);
and U3489 (N_3489,N_2492,N_2718);
xor U3490 (N_3490,N_2914,N_3015);
or U3491 (N_3491,N_3020,N_2823);
nand U3492 (N_3492,N_3084,N_3008);
and U3493 (N_3493,N_2921,N_3076);
and U3494 (N_3494,N_2615,N_2664);
xnor U3495 (N_3495,N_3010,N_2889);
nor U3496 (N_3496,N_2792,N_2510);
and U3497 (N_3497,N_3062,N_2809);
xor U3498 (N_3498,N_2682,N_2842);
and U3499 (N_3499,N_2509,N_2956);
xnor U3500 (N_3500,N_2765,N_2542);
and U3501 (N_3501,N_3100,N_3085);
xor U3502 (N_3502,N_2617,N_3094);
nor U3503 (N_3503,N_2806,N_2816);
xnor U3504 (N_3504,N_2513,N_2424);
or U3505 (N_3505,N_2479,N_2642);
nor U3506 (N_3506,N_2434,N_2970);
nor U3507 (N_3507,N_3059,N_3029);
and U3508 (N_3508,N_2891,N_2786);
nand U3509 (N_3509,N_3152,N_3144);
nor U3510 (N_3510,N_2684,N_3140);
or U3511 (N_3511,N_2543,N_2750);
and U3512 (N_3512,N_2482,N_3183);
nand U3513 (N_3513,N_2836,N_2883);
and U3514 (N_3514,N_2599,N_2707);
nor U3515 (N_3515,N_2511,N_2581);
nand U3516 (N_3516,N_3156,N_2697);
and U3517 (N_3517,N_2957,N_3060);
nor U3518 (N_3518,N_2504,N_2493);
and U3519 (N_3519,N_2935,N_2777);
xnor U3520 (N_3520,N_3147,N_3066);
and U3521 (N_3521,N_3184,N_3079);
nand U3522 (N_3522,N_2976,N_2704);
nand U3523 (N_3523,N_2894,N_2838);
nor U3524 (N_3524,N_2496,N_2814);
or U3525 (N_3525,N_2545,N_2598);
xor U3526 (N_3526,N_2947,N_3149);
and U3527 (N_3527,N_2897,N_2435);
and U3528 (N_3528,N_3145,N_2960);
nor U3529 (N_3529,N_2746,N_2620);
nor U3530 (N_3530,N_2607,N_2882);
nand U3531 (N_3531,N_2999,N_2503);
and U3532 (N_3532,N_3075,N_3181);
or U3533 (N_3533,N_2401,N_3026);
and U3534 (N_3534,N_3046,N_2419);
nor U3535 (N_3535,N_2641,N_3121);
nor U3536 (N_3536,N_2901,N_2639);
or U3537 (N_3537,N_2969,N_3053);
nand U3538 (N_3538,N_2789,N_2745);
and U3539 (N_3539,N_2896,N_2754);
xnor U3540 (N_3540,N_2716,N_2498);
nor U3541 (N_3541,N_2708,N_3108);
nand U3542 (N_3542,N_3034,N_2808);
nor U3543 (N_3543,N_3168,N_2614);
xnor U3544 (N_3544,N_2508,N_2472);
or U3545 (N_3545,N_3186,N_2865);
or U3546 (N_3546,N_2753,N_2853);
xnor U3547 (N_3547,N_2685,N_3191);
xnor U3548 (N_3548,N_2431,N_2784);
and U3549 (N_3549,N_2973,N_2519);
or U3550 (N_3550,N_2531,N_3021);
and U3551 (N_3551,N_3133,N_2687);
nand U3552 (N_3552,N_2830,N_2912);
or U3553 (N_3553,N_3142,N_2843);
and U3554 (N_3554,N_2690,N_2944);
nand U3555 (N_3555,N_2846,N_2407);
nand U3556 (N_3556,N_2445,N_2931);
xor U3557 (N_3557,N_3128,N_2674);
or U3558 (N_3558,N_2470,N_2721);
and U3559 (N_3559,N_2858,N_2551);
nor U3560 (N_3560,N_2698,N_2701);
and U3561 (N_3561,N_3124,N_2909);
and U3562 (N_3562,N_2943,N_2923);
nor U3563 (N_3563,N_2820,N_3127);
or U3564 (N_3564,N_2569,N_2886);
and U3565 (N_3565,N_2963,N_3106);
or U3566 (N_3566,N_2798,N_3096);
and U3567 (N_3567,N_2480,N_3148);
nand U3568 (N_3568,N_2711,N_3197);
nor U3569 (N_3569,N_2989,N_2794);
xnor U3570 (N_3570,N_2459,N_2893);
xnor U3571 (N_3571,N_2411,N_2839);
nand U3572 (N_3572,N_2827,N_2526);
nand U3573 (N_3573,N_3109,N_2661);
or U3574 (N_3574,N_2945,N_2932);
or U3575 (N_3575,N_3158,N_2845);
nor U3576 (N_3576,N_2421,N_2678);
and U3577 (N_3577,N_2942,N_3104);
xnor U3578 (N_3578,N_2427,N_3188);
or U3579 (N_3579,N_3189,N_2621);
and U3580 (N_3580,N_2490,N_2977);
or U3581 (N_3581,N_2848,N_3018);
or U3582 (N_3582,N_3135,N_2562);
nor U3583 (N_3583,N_3011,N_2626);
or U3584 (N_3584,N_3038,N_2764);
nor U3585 (N_3585,N_3071,N_3030);
nor U3586 (N_3586,N_3118,N_3048);
and U3587 (N_3587,N_2917,N_3151);
xor U3588 (N_3588,N_3155,N_2844);
nand U3589 (N_3589,N_2859,N_3031);
or U3590 (N_3590,N_2454,N_2547);
xor U3591 (N_3591,N_2860,N_2616);
nand U3592 (N_3592,N_2418,N_2527);
nor U3593 (N_3593,N_2403,N_2497);
xnor U3594 (N_3594,N_2446,N_2402);
nand U3595 (N_3595,N_2788,N_3056);
nand U3596 (N_3596,N_2540,N_2558);
nor U3597 (N_3597,N_3170,N_2453);
nor U3598 (N_3598,N_2560,N_2851);
xor U3599 (N_3599,N_3117,N_2903);
nand U3600 (N_3600,N_3026,N_3072);
nor U3601 (N_3601,N_3198,N_3164);
nor U3602 (N_3602,N_2962,N_3027);
or U3603 (N_3603,N_2750,N_2866);
and U3604 (N_3604,N_2760,N_2646);
or U3605 (N_3605,N_2971,N_2734);
nor U3606 (N_3606,N_2774,N_2427);
nand U3607 (N_3607,N_3139,N_2613);
xor U3608 (N_3608,N_2754,N_2644);
xnor U3609 (N_3609,N_2912,N_3160);
and U3610 (N_3610,N_2657,N_3049);
xor U3611 (N_3611,N_2566,N_2447);
nor U3612 (N_3612,N_2549,N_2713);
xor U3613 (N_3613,N_2581,N_2579);
xnor U3614 (N_3614,N_2963,N_3194);
nand U3615 (N_3615,N_2951,N_3088);
and U3616 (N_3616,N_2776,N_3135);
and U3617 (N_3617,N_2400,N_2634);
nor U3618 (N_3618,N_2852,N_3123);
nand U3619 (N_3619,N_2784,N_2477);
xnor U3620 (N_3620,N_2833,N_3032);
and U3621 (N_3621,N_2867,N_3121);
and U3622 (N_3622,N_2677,N_2547);
nand U3623 (N_3623,N_2554,N_2664);
nand U3624 (N_3624,N_2809,N_2760);
and U3625 (N_3625,N_2574,N_2562);
xor U3626 (N_3626,N_2550,N_2957);
nand U3627 (N_3627,N_2591,N_2560);
and U3628 (N_3628,N_2502,N_2480);
and U3629 (N_3629,N_2404,N_2552);
and U3630 (N_3630,N_2786,N_3021);
nor U3631 (N_3631,N_2686,N_3052);
and U3632 (N_3632,N_2930,N_2790);
nor U3633 (N_3633,N_3066,N_2834);
nand U3634 (N_3634,N_2747,N_2512);
or U3635 (N_3635,N_2470,N_2777);
nand U3636 (N_3636,N_2657,N_2579);
nor U3637 (N_3637,N_2441,N_2881);
xor U3638 (N_3638,N_2855,N_3044);
nor U3639 (N_3639,N_2427,N_3143);
nor U3640 (N_3640,N_2557,N_2725);
or U3641 (N_3641,N_2516,N_3184);
nor U3642 (N_3642,N_2621,N_2425);
nor U3643 (N_3643,N_2509,N_2579);
or U3644 (N_3644,N_2803,N_2870);
nor U3645 (N_3645,N_2774,N_2436);
nand U3646 (N_3646,N_3114,N_2970);
and U3647 (N_3647,N_2594,N_2496);
nor U3648 (N_3648,N_2567,N_2831);
xor U3649 (N_3649,N_2561,N_2579);
nand U3650 (N_3650,N_2851,N_2639);
xor U3651 (N_3651,N_2656,N_2881);
nor U3652 (N_3652,N_2735,N_2883);
nor U3653 (N_3653,N_3195,N_3029);
nand U3654 (N_3654,N_3018,N_3041);
or U3655 (N_3655,N_2464,N_2624);
nor U3656 (N_3656,N_2810,N_3035);
nor U3657 (N_3657,N_2622,N_3053);
nand U3658 (N_3658,N_2444,N_3100);
and U3659 (N_3659,N_2632,N_3183);
or U3660 (N_3660,N_3045,N_3006);
nor U3661 (N_3661,N_2970,N_3109);
or U3662 (N_3662,N_2530,N_2492);
and U3663 (N_3663,N_2925,N_2863);
nor U3664 (N_3664,N_2681,N_2458);
or U3665 (N_3665,N_2819,N_2717);
or U3666 (N_3666,N_2922,N_2966);
xor U3667 (N_3667,N_2667,N_2497);
and U3668 (N_3668,N_2803,N_2730);
and U3669 (N_3669,N_3038,N_2422);
or U3670 (N_3670,N_2753,N_2518);
xnor U3671 (N_3671,N_2907,N_3190);
nand U3672 (N_3672,N_2654,N_2450);
or U3673 (N_3673,N_2763,N_2472);
xor U3674 (N_3674,N_3064,N_2977);
nand U3675 (N_3675,N_3172,N_3183);
xnor U3676 (N_3676,N_3057,N_2479);
nand U3677 (N_3677,N_2621,N_2507);
or U3678 (N_3678,N_2597,N_2898);
xor U3679 (N_3679,N_2829,N_2962);
nor U3680 (N_3680,N_3142,N_2967);
or U3681 (N_3681,N_2507,N_2510);
xnor U3682 (N_3682,N_3157,N_3089);
or U3683 (N_3683,N_2847,N_2519);
or U3684 (N_3684,N_2845,N_3077);
and U3685 (N_3685,N_3012,N_2511);
xnor U3686 (N_3686,N_3175,N_2628);
xor U3687 (N_3687,N_3154,N_3137);
nor U3688 (N_3688,N_2725,N_2666);
xnor U3689 (N_3689,N_3117,N_3193);
xnor U3690 (N_3690,N_2841,N_2551);
xnor U3691 (N_3691,N_3016,N_2793);
or U3692 (N_3692,N_2947,N_2411);
nand U3693 (N_3693,N_2432,N_2541);
xnor U3694 (N_3694,N_2882,N_2877);
and U3695 (N_3695,N_3005,N_2463);
nand U3696 (N_3696,N_2877,N_2975);
nand U3697 (N_3697,N_3059,N_3061);
and U3698 (N_3698,N_2572,N_2468);
nand U3699 (N_3699,N_2922,N_2403);
or U3700 (N_3700,N_3100,N_3071);
or U3701 (N_3701,N_2829,N_2875);
xor U3702 (N_3702,N_2449,N_3153);
nand U3703 (N_3703,N_3115,N_2792);
nand U3704 (N_3704,N_2827,N_3114);
nor U3705 (N_3705,N_2513,N_2407);
and U3706 (N_3706,N_3005,N_2563);
nand U3707 (N_3707,N_2744,N_2557);
xnor U3708 (N_3708,N_2997,N_3048);
or U3709 (N_3709,N_3041,N_2815);
nand U3710 (N_3710,N_2525,N_2788);
xnor U3711 (N_3711,N_2732,N_3009);
xor U3712 (N_3712,N_2852,N_3042);
nor U3713 (N_3713,N_2795,N_2858);
and U3714 (N_3714,N_2573,N_2851);
or U3715 (N_3715,N_3098,N_2469);
nor U3716 (N_3716,N_2420,N_2747);
and U3717 (N_3717,N_2857,N_2800);
and U3718 (N_3718,N_2601,N_2768);
or U3719 (N_3719,N_3012,N_2781);
nor U3720 (N_3720,N_2599,N_2720);
nand U3721 (N_3721,N_2900,N_2977);
or U3722 (N_3722,N_2504,N_2791);
nand U3723 (N_3723,N_2401,N_2576);
and U3724 (N_3724,N_2980,N_2618);
nand U3725 (N_3725,N_3111,N_2897);
xnor U3726 (N_3726,N_3133,N_2931);
nand U3727 (N_3727,N_2513,N_2521);
or U3728 (N_3728,N_2549,N_2851);
xnor U3729 (N_3729,N_2431,N_2532);
nor U3730 (N_3730,N_2549,N_2815);
nand U3731 (N_3731,N_2415,N_2728);
nor U3732 (N_3732,N_3056,N_2721);
and U3733 (N_3733,N_2764,N_2731);
nor U3734 (N_3734,N_2884,N_2555);
or U3735 (N_3735,N_2860,N_2994);
or U3736 (N_3736,N_2991,N_2820);
or U3737 (N_3737,N_3108,N_2877);
nor U3738 (N_3738,N_3114,N_2666);
nand U3739 (N_3739,N_2496,N_2969);
nand U3740 (N_3740,N_3010,N_2535);
nand U3741 (N_3741,N_2601,N_2676);
xor U3742 (N_3742,N_2476,N_2789);
and U3743 (N_3743,N_2645,N_2786);
and U3744 (N_3744,N_2414,N_3113);
xnor U3745 (N_3745,N_2547,N_2560);
and U3746 (N_3746,N_2526,N_3149);
xnor U3747 (N_3747,N_2981,N_2996);
and U3748 (N_3748,N_2727,N_3188);
nor U3749 (N_3749,N_2616,N_3010);
xnor U3750 (N_3750,N_2902,N_2534);
and U3751 (N_3751,N_2969,N_2747);
xnor U3752 (N_3752,N_2627,N_3183);
or U3753 (N_3753,N_2881,N_2437);
xnor U3754 (N_3754,N_2872,N_2956);
nand U3755 (N_3755,N_3014,N_2446);
or U3756 (N_3756,N_2818,N_3018);
and U3757 (N_3757,N_2904,N_3043);
or U3758 (N_3758,N_2860,N_2717);
nand U3759 (N_3759,N_2694,N_2972);
and U3760 (N_3760,N_2603,N_3028);
nor U3761 (N_3761,N_3023,N_3073);
and U3762 (N_3762,N_2728,N_2798);
and U3763 (N_3763,N_2402,N_2565);
nand U3764 (N_3764,N_3051,N_2860);
nand U3765 (N_3765,N_2670,N_3015);
xor U3766 (N_3766,N_3049,N_2429);
nor U3767 (N_3767,N_2559,N_2720);
or U3768 (N_3768,N_2737,N_3037);
nor U3769 (N_3769,N_2883,N_3176);
nor U3770 (N_3770,N_2584,N_2766);
nor U3771 (N_3771,N_3081,N_3059);
xnor U3772 (N_3772,N_3115,N_2832);
and U3773 (N_3773,N_2456,N_2957);
xnor U3774 (N_3774,N_2510,N_2469);
xor U3775 (N_3775,N_2977,N_2529);
nor U3776 (N_3776,N_2592,N_2510);
or U3777 (N_3777,N_3140,N_2880);
or U3778 (N_3778,N_2529,N_2958);
nor U3779 (N_3779,N_2905,N_3106);
or U3780 (N_3780,N_2728,N_2736);
and U3781 (N_3781,N_2785,N_2499);
xnor U3782 (N_3782,N_3095,N_3142);
nand U3783 (N_3783,N_2825,N_3027);
xnor U3784 (N_3784,N_3121,N_2864);
nand U3785 (N_3785,N_2937,N_3011);
or U3786 (N_3786,N_2756,N_2938);
nand U3787 (N_3787,N_2874,N_2490);
nand U3788 (N_3788,N_2486,N_3048);
or U3789 (N_3789,N_3062,N_2855);
nand U3790 (N_3790,N_3077,N_2663);
nor U3791 (N_3791,N_2890,N_3150);
xnor U3792 (N_3792,N_2433,N_2636);
nor U3793 (N_3793,N_2937,N_2477);
or U3794 (N_3794,N_3131,N_2835);
or U3795 (N_3795,N_2994,N_2448);
or U3796 (N_3796,N_2803,N_2400);
xor U3797 (N_3797,N_3069,N_3042);
nor U3798 (N_3798,N_3023,N_3028);
nor U3799 (N_3799,N_2696,N_2754);
xnor U3800 (N_3800,N_2926,N_2513);
nor U3801 (N_3801,N_3010,N_3167);
or U3802 (N_3802,N_3189,N_3173);
nand U3803 (N_3803,N_2532,N_3156);
nor U3804 (N_3804,N_3195,N_2585);
nor U3805 (N_3805,N_2707,N_2557);
nor U3806 (N_3806,N_3072,N_2487);
nor U3807 (N_3807,N_3165,N_3142);
xor U3808 (N_3808,N_2543,N_2524);
nand U3809 (N_3809,N_2902,N_2911);
nor U3810 (N_3810,N_2405,N_2926);
xnor U3811 (N_3811,N_2433,N_2619);
nor U3812 (N_3812,N_2470,N_2844);
nor U3813 (N_3813,N_3028,N_2832);
xor U3814 (N_3814,N_3041,N_2982);
xnor U3815 (N_3815,N_2994,N_2727);
and U3816 (N_3816,N_2739,N_3072);
nor U3817 (N_3817,N_3170,N_2839);
nand U3818 (N_3818,N_2832,N_2685);
xnor U3819 (N_3819,N_2476,N_2671);
nor U3820 (N_3820,N_2963,N_2896);
and U3821 (N_3821,N_2634,N_2749);
nor U3822 (N_3822,N_2931,N_3052);
xnor U3823 (N_3823,N_2949,N_3113);
or U3824 (N_3824,N_2473,N_2793);
or U3825 (N_3825,N_2912,N_3085);
nand U3826 (N_3826,N_3197,N_2648);
nand U3827 (N_3827,N_2498,N_2808);
nor U3828 (N_3828,N_2439,N_3091);
nand U3829 (N_3829,N_2628,N_2803);
xor U3830 (N_3830,N_2708,N_2932);
and U3831 (N_3831,N_2499,N_3039);
or U3832 (N_3832,N_3109,N_2459);
and U3833 (N_3833,N_2647,N_2659);
or U3834 (N_3834,N_2718,N_2703);
nand U3835 (N_3835,N_2862,N_2827);
and U3836 (N_3836,N_2965,N_3148);
nor U3837 (N_3837,N_2405,N_2724);
nor U3838 (N_3838,N_3098,N_2677);
xnor U3839 (N_3839,N_2556,N_2606);
nand U3840 (N_3840,N_3048,N_2501);
or U3841 (N_3841,N_2894,N_3079);
and U3842 (N_3842,N_2416,N_2735);
nor U3843 (N_3843,N_2693,N_2611);
nor U3844 (N_3844,N_3163,N_3120);
xnor U3845 (N_3845,N_2729,N_2569);
and U3846 (N_3846,N_2902,N_2954);
and U3847 (N_3847,N_2526,N_2879);
or U3848 (N_3848,N_3025,N_2654);
nand U3849 (N_3849,N_2442,N_2666);
nor U3850 (N_3850,N_2930,N_2705);
and U3851 (N_3851,N_3047,N_2548);
xor U3852 (N_3852,N_2849,N_2528);
or U3853 (N_3853,N_2841,N_3044);
and U3854 (N_3854,N_3170,N_2407);
and U3855 (N_3855,N_2499,N_2545);
xor U3856 (N_3856,N_2513,N_2505);
xor U3857 (N_3857,N_2922,N_2676);
xnor U3858 (N_3858,N_3101,N_3052);
nor U3859 (N_3859,N_2487,N_2644);
nand U3860 (N_3860,N_2822,N_2800);
xor U3861 (N_3861,N_3010,N_2988);
nor U3862 (N_3862,N_2651,N_2897);
xnor U3863 (N_3863,N_2862,N_2848);
nand U3864 (N_3864,N_2770,N_3048);
and U3865 (N_3865,N_2589,N_3039);
and U3866 (N_3866,N_2711,N_2429);
xor U3867 (N_3867,N_2796,N_2747);
nor U3868 (N_3868,N_2724,N_2894);
nor U3869 (N_3869,N_2711,N_2619);
and U3870 (N_3870,N_2696,N_3177);
or U3871 (N_3871,N_2836,N_2920);
or U3872 (N_3872,N_2912,N_2661);
nand U3873 (N_3873,N_2629,N_2452);
nand U3874 (N_3874,N_2443,N_2714);
nand U3875 (N_3875,N_3125,N_2571);
xnor U3876 (N_3876,N_2898,N_2900);
xnor U3877 (N_3877,N_2750,N_3137);
nor U3878 (N_3878,N_2936,N_2994);
or U3879 (N_3879,N_2657,N_2524);
and U3880 (N_3880,N_2638,N_2493);
or U3881 (N_3881,N_2738,N_2587);
nand U3882 (N_3882,N_3138,N_3152);
xnor U3883 (N_3883,N_3110,N_2508);
and U3884 (N_3884,N_3059,N_2757);
nand U3885 (N_3885,N_2946,N_2817);
nor U3886 (N_3886,N_2963,N_2976);
nand U3887 (N_3887,N_2538,N_2520);
or U3888 (N_3888,N_2791,N_2454);
nand U3889 (N_3889,N_2844,N_2932);
and U3890 (N_3890,N_2858,N_2536);
nand U3891 (N_3891,N_3085,N_2453);
nand U3892 (N_3892,N_2934,N_2828);
nor U3893 (N_3893,N_3159,N_2876);
xor U3894 (N_3894,N_3127,N_2708);
nor U3895 (N_3895,N_2941,N_3191);
nand U3896 (N_3896,N_2705,N_2714);
nand U3897 (N_3897,N_2475,N_2711);
nor U3898 (N_3898,N_2910,N_3104);
and U3899 (N_3899,N_3186,N_2417);
xor U3900 (N_3900,N_3017,N_3072);
and U3901 (N_3901,N_3022,N_2548);
nand U3902 (N_3902,N_3169,N_2508);
nand U3903 (N_3903,N_2499,N_2627);
nand U3904 (N_3904,N_2924,N_2758);
nand U3905 (N_3905,N_2950,N_3043);
xnor U3906 (N_3906,N_2681,N_2743);
xor U3907 (N_3907,N_2526,N_2784);
xnor U3908 (N_3908,N_2656,N_2591);
xor U3909 (N_3909,N_2946,N_3022);
and U3910 (N_3910,N_2730,N_2900);
or U3911 (N_3911,N_3033,N_2975);
nor U3912 (N_3912,N_2659,N_2670);
nand U3913 (N_3913,N_2704,N_2734);
and U3914 (N_3914,N_2697,N_3166);
nor U3915 (N_3915,N_3012,N_2430);
xor U3916 (N_3916,N_2903,N_2730);
xor U3917 (N_3917,N_2637,N_3163);
nand U3918 (N_3918,N_2629,N_3056);
nand U3919 (N_3919,N_2517,N_2470);
xnor U3920 (N_3920,N_2779,N_2874);
and U3921 (N_3921,N_3122,N_2990);
and U3922 (N_3922,N_2516,N_2862);
nor U3923 (N_3923,N_2840,N_3034);
or U3924 (N_3924,N_2857,N_3067);
or U3925 (N_3925,N_2909,N_2945);
nand U3926 (N_3926,N_3178,N_3092);
or U3927 (N_3927,N_2744,N_2841);
nand U3928 (N_3928,N_2996,N_2974);
nor U3929 (N_3929,N_2935,N_2528);
nor U3930 (N_3930,N_2732,N_2716);
or U3931 (N_3931,N_2827,N_2789);
nor U3932 (N_3932,N_2908,N_2748);
xor U3933 (N_3933,N_2451,N_2608);
xnor U3934 (N_3934,N_2942,N_3018);
nor U3935 (N_3935,N_2734,N_2441);
nand U3936 (N_3936,N_2464,N_2581);
nand U3937 (N_3937,N_2552,N_3028);
xor U3938 (N_3938,N_3030,N_2597);
or U3939 (N_3939,N_3191,N_3023);
or U3940 (N_3940,N_3174,N_2971);
xor U3941 (N_3941,N_2659,N_2958);
nand U3942 (N_3942,N_3083,N_2610);
or U3943 (N_3943,N_2621,N_2630);
and U3944 (N_3944,N_3035,N_3172);
nor U3945 (N_3945,N_2921,N_2800);
or U3946 (N_3946,N_2674,N_2883);
nand U3947 (N_3947,N_3091,N_2684);
nand U3948 (N_3948,N_2556,N_3118);
nor U3949 (N_3949,N_2747,N_3043);
nor U3950 (N_3950,N_2705,N_2536);
nor U3951 (N_3951,N_2545,N_2709);
nor U3952 (N_3952,N_3098,N_2696);
or U3953 (N_3953,N_2752,N_2492);
nor U3954 (N_3954,N_2510,N_2994);
or U3955 (N_3955,N_3086,N_2646);
nor U3956 (N_3956,N_2643,N_3027);
xnor U3957 (N_3957,N_2879,N_2816);
nor U3958 (N_3958,N_2846,N_3042);
and U3959 (N_3959,N_2944,N_2614);
and U3960 (N_3960,N_2532,N_2870);
nor U3961 (N_3961,N_2612,N_3180);
or U3962 (N_3962,N_3127,N_3061);
xor U3963 (N_3963,N_2689,N_3097);
and U3964 (N_3964,N_2625,N_2453);
or U3965 (N_3965,N_2540,N_2417);
nand U3966 (N_3966,N_2505,N_2636);
xor U3967 (N_3967,N_2649,N_2873);
or U3968 (N_3968,N_2668,N_2707);
xnor U3969 (N_3969,N_2746,N_3100);
or U3970 (N_3970,N_2509,N_3189);
and U3971 (N_3971,N_2694,N_2869);
nand U3972 (N_3972,N_2959,N_2401);
nor U3973 (N_3973,N_2537,N_2476);
xnor U3974 (N_3974,N_3105,N_2663);
and U3975 (N_3975,N_2910,N_2622);
nor U3976 (N_3976,N_3134,N_2907);
xor U3977 (N_3977,N_2558,N_2412);
nor U3978 (N_3978,N_2433,N_2921);
and U3979 (N_3979,N_2544,N_2969);
nor U3980 (N_3980,N_2768,N_3054);
xnor U3981 (N_3981,N_2478,N_2685);
or U3982 (N_3982,N_2928,N_3064);
nand U3983 (N_3983,N_2489,N_2803);
or U3984 (N_3984,N_2780,N_3007);
and U3985 (N_3985,N_2958,N_2774);
nor U3986 (N_3986,N_2893,N_2708);
or U3987 (N_3987,N_2999,N_2616);
nand U3988 (N_3988,N_3099,N_2445);
nor U3989 (N_3989,N_2700,N_3068);
xnor U3990 (N_3990,N_3173,N_2892);
nand U3991 (N_3991,N_2426,N_3022);
and U3992 (N_3992,N_3021,N_2558);
and U3993 (N_3993,N_3002,N_2789);
nor U3994 (N_3994,N_2706,N_2712);
xor U3995 (N_3995,N_2637,N_3073);
xor U3996 (N_3996,N_3087,N_3198);
nor U3997 (N_3997,N_2666,N_2888);
or U3998 (N_3998,N_2653,N_2733);
nand U3999 (N_3999,N_2694,N_3093);
nor U4000 (N_4000,N_3272,N_3353);
nor U4001 (N_4001,N_3385,N_3460);
and U4002 (N_4002,N_3815,N_3521);
nor U4003 (N_4003,N_3605,N_3735);
nand U4004 (N_4004,N_3564,N_3297);
nand U4005 (N_4005,N_3275,N_3550);
nor U4006 (N_4006,N_3859,N_3621);
nand U4007 (N_4007,N_3343,N_3294);
nand U4008 (N_4008,N_3260,N_3854);
nand U4009 (N_4009,N_3888,N_3963);
xor U4010 (N_4010,N_3504,N_3313);
or U4011 (N_4011,N_3763,N_3723);
or U4012 (N_4012,N_3202,N_3246);
or U4013 (N_4013,N_3996,N_3666);
nor U4014 (N_4014,N_3865,N_3507);
or U4015 (N_4015,N_3549,N_3221);
nand U4016 (N_4016,N_3845,N_3810);
or U4017 (N_4017,N_3218,N_3395);
xnor U4018 (N_4018,N_3873,N_3748);
or U4019 (N_4019,N_3753,N_3286);
nor U4020 (N_4020,N_3375,N_3230);
xor U4021 (N_4021,N_3441,N_3515);
xor U4022 (N_4022,N_3821,N_3875);
or U4023 (N_4023,N_3426,N_3442);
and U4024 (N_4024,N_3971,N_3766);
nor U4025 (N_4025,N_3247,N_3572);
nor U4026 (N_4026,N_3581,N_3643);
and U4027 (N_4027,N_3390,N_3274);
nand U4028 (N_4028,N_3224,N_3596);
and U4029 (N_4029,N_3520,N_3979);
or U4030 (N_4030,N_3849,N_3938);
nor U4031 (N_4031,N_3529,N_3619);
nand U4032 (N_4032,N_3588,N_3526);
nand U4033 (N_4033,N_3743,N_3477);
and U4034 (N_4034,N_3334,N_3661);
and U4035 (N_4035,N_3695,N_3490);
nand U4036 (N_4036,N_3256,N_3703);
nor U4037 (N_4037,N_3687,N_3316);
or U4038 (N_4038,N_3842,N_3540);
nand U4039 (N_4039,N_3911,N_3203);
nand U4040 (N_4040,N_3780,N_3946);
xor U4041 (N_4041,N_3788,N_3461);
or U4042 (N_4042,N_3265,N_3555);
or U4043 (N_4043,N_3280,N_3427);
xnor U4044 (N_4044,N_3519,N_3250);
nor U4045 (N_4045,N_3301,N_3225);
xor U4046 (N_4046,N_3929,N_3864);
and U4047 (N_4047,N_3544,N_3418);
and U4048 (N_4048,N_3463,N_3640);
nand U4049 (N_4049,N_3568,N_3925);
nand U4050 (N_4050,N_3235,N_3424);
or U4051 (N_4051,N_3921,N_3811);
and U4052 (N_4052,N_3219,N_3893);
nor U4053 (N_4053,N_3908,N_3680);
nand U4054 (N_4054,N_3593,N_3878);
nand U4055 (N_4055,N_3953,N_3567);
and U4056 (N_4056,N_3772,N_3401);
or U4057 (N_4057,N_3311,N_3384);
or U4058 (N_4058,N_3415,N_3903);
xor U4059 (N_4059,N_3691,N_3833);
xnor U4060 (N_4060,N_3437,N_3764);
and U4061 (N_4061,N_3779,N_3603);
nand U4062 (N_4062,N_3647,N_3853);
nand U4063 (N_4063,N_3454,N_3350);
or U4064 (N_4064,N_3818,N_3407);
and U4065 (N_4065,N_3587,N_3402);
or U4066 (N_4066,N_3308,N_3760);
xor U4067 (N_4067,N_3312,N_3776);
nand U4068 (N_4068,N_3917,N_3399);
nor U4069 (N_4069,N_3335,N_3293);
nor U4070 (N_4070,N_3848,N_3266);
nand U4071 (N_4071,N_3993,N_3416);
and U4072 (N_4072,N_3827,N_3667);
nand U4073 (N_4073,N_3916,N_3289);
nand U4074 (N_4074,N_3762,N_3665);
nand U4075 (N_4075,N_3969,N_3278);
nand U4076 (N_4076,N_3290,N_3943);
nand U4077 (N_4077,N_3486,N_3509);
nand U4078 (N_4078,N_3361,N_3471);
or U4079 (N_4079,N_3356,N_3267);
nor U4080 (N_4080,N_3400,N_3798);
nor U4081 (N_4081,N_3360,N_3967);
nand U4082 (N_4082,N_3420,N_3241);
nand U4083 (N_4083,N_3708,N_3998);
nor U4084 (N_4084,N_3704,N_3210);
nand U4085 (N_4085,N_3654,N_3444);
nand U4086 (N_4086,N_3448,N_3981);
or U4087 (N_4087,N_3326,N_3789);
xnor U4088 (N_4088,N_3851,N_3988);
nand U4089 (N_4089,N_3485,N_3411);
nand U4090 (N_4090,N_3434,N_3589);
and U4091 (N_4091,N_3333,N_3556);
or U4092 (N_4092,N_3626,N_3577);
or U4093 (N_4093,N_3775,N_3931);
xor U4094 (N_4094,N_3215,N_3468);
nor U4095 (N_4095,N_3862,N_3646);
nand U4096 (N_4096,N_3317,N_3736);
and U4097 (N_4097,N_3462,N_3822);
and U4098 (N_4098,N_3273,N_3877);
or U4099 (N_4099,N_3599,N_3709);
xnor U4100 (N_4100,N_3569,N_3954);
nand U4101 (N_4101,N_3984,N_3770);
and U4102 (N_4102,N_3870,N_3331);
and U4103 (N_4103,N_3627,N_3548);
nor U4104 (N_4104,N_3579,N_3522);
nor U4105 (N_4105,N_3814,N_3761);
and U4106 (N_4106,N_3670,N_3320);
nand U4107 (N_4107,N_3834,N_3406);
xor U4108 (N_4108,N_3562,N_3573);
nor U4109 (N_4109,N_3642,N_3994);
nand U4110 (N_4110,N_3480,N_3724);
xor U4111 (N_4111,N_3389,N_3804);
and U4112 (N_4112,N_3547,N_3254);
nor U4113 (N_4113,N_3980,N_3365);
nor U4114 (N_4114,N_3876,N_3754);
or U4115 (N_4115,N_3511,N_3378);
and U4116 (N_4116,N_3580,N_3481);
nand U4117 (N_4117,N_3496,N_3346);
nor U4118 (N_4118,N_3238,N_3913);
and U4119 (N_4119,N_3629,N_3970);
nand U4120 (N_4120,N_3261,N_3592);
and U4121 (N_4121,N_3965,N_3591);
nor U4122 (N_4122,N_3826,N_3679);
or U4123 (N_4123,N_3872,N_3889);
xnor U4124 (N_4124,N_3348,N_3809);
nor U4125 (N_4125,N_3910,N_3227);
nand U4126 (N_4126,N_3469,N_3950);
nor U4127 (N_4127,N_3730,N_3533);
and U4128 (N_4128,N_3684,N_3492);
nand U4129 (N_4129,N_3682,N_3303);
or U4130 (N_4130,N_3398,N_3291);
nor U4131 (N_4131,N_3371,N_3982);
xor U4132 (N_4132,N_3936,N_3553);
nand U4133 (N_4133,N_3372,N_3295);
nor U4134 (N_4134,N_3505,N_3257);
nor U4135 (N_4135,N_3675,N_3287);
nor U4136 (N_4136,N_3516,N_3885);
xnor U4137 (N_4137,N_3902,N_3719);
and U4138 (N_4138,N_3574,N_3850);
or U4139 (N_4139,N_3370,N_3551);
xnor U4140 (N_4140,N_3991,N_3276);
nand U4141 (N_4141,N_3373,N_3394);
xnor U4142 (N_4142,N_3959,N_3831);
nand U4143 (N_4143,N_3807,N_3841);
xor U4144 (N_4144,N_3242,N_3524);
or U4145 (N_4145,N_3734,N_3620);
or U4146 (N_4146,N_3676,N_3816);
or U4147 (N_4147,N_3635,N_3905);
nor U4148 (N_4148,N_3582,N_3270);
or U4149 (N_4149,N_3337,N_3302);
and U4150 (N_4150,N_3729,N_3768);
nor U4151 (N_4151,N_3881,N_3344);
or U4152 (N_4152,N_3570,N_3906);
nor U4153 (N_4153,N_3380,N_3957);
and U4154 (N_4154,N_3920,N_3721);
or U4155 (N_4155,N_3467,N_3498);
nand U4156 (N_4156,N_3922,N_3632);
or U4157 (N_4157,N_3649,N_3749);
and U4158 (N_4158,N_3229,N_3506);
nor U4159 (N_4159,N_3837,N_3939);
nor U4160 (N_4160,N_3707,N_3262);
xor U4161 (N_4161,N_3586,N_3829);
and U4162 (N_4162,N_3484,N_3694);
nor U4163 (N_4163,N_3852,N_3539);
xor U4164 (N_4164,N_3501,N_3617);
nand U4165 (N_4165,N_3607,N_3783);
and U4166 (N_4166,N_3824,N_3476);
and U4167 (N_4167,N_3631,N_3512);
or U4168 (N_4168,N_3387,N_3948);
nand U4169 (N_4169,N_3808,N_3795);
or U4170 (N_4170,N_3537,N_3423);
or U4171 (N_4171,N_3915,N_3397);
xor U4172 (N_4172,N_3801,N_3858);
nand U4173 (N_4173,N_3820,N_3895);
or U4174 (N_4174,N_3937,N_3933);
and U4175 (N_4175,N_3381,N_3497);
xor U4176 (N_4176,N_3514,N_3200);
and U4177 (N_4177,N_3493,N_3961);
xor U4178 (N_4178,N_3288,N_3248);
nand U4179 (N_4179,N_3292,N_3517);
and U4180 (N_4180,N_3536,N_3692);
or U4181 (N_4181,N_3324,N_3403);
or U4182 (N_4182,N_3792,N_3330);
or U4183 (N_4183,N_3987,N_3594);
nand U4184 (N_4184,N_3304,N_3855);
xor U4185 (N_4185,N_3787,N_3585);
nor U4186 (N_4186,N_3237,N_3616);
and U4187 (N_4187,N_3638,N_3502);
or U4188 (N_4188,N_3660,N_3992);
nand U4189 (N_4189,N_3306,N_3727);
xor U4190 (N_4190,N_3758,N_3345);
nor U4191 (N_4191,N_3636,N_3447);
nand U4192 (N_4192,N_3451,N_3894);
or U4193 (N_4193,N_3773,N_3909);
xor U4194 (N_4194,N_3802,N_3534);
nor U4195 (N_4195,N_3483,N_3258);
and U4196 (N_4196,N_3685,N_3264);
nor U4197 (N_4197,N_3769,N_3774);
and U4198 (N_4198,N_3296,N_3655);
nand U4199 (N_4199,N_3377,N_3318);
and U4200 (N_4200,N_3563,N_3470);
and U4201 (N_4201,N_3923,N_3790);
nor U4202 (N_4202,N_3733,N_3503);
and U4203 (N_4203,N_3871,N_3771);
and U4204 (N_4204,N_3722,N_3355);
or U4205 (N_4205,N_3847,N_3641);
and U4206 (N_4206,N_3212,N_3874);
nor U4207 (N_4207,N_3891,N_3673);
xnor U4208 (N_4208,N_3651,N_3609);
xnor U4209 (N_4209,N_3478,N_3216);
nand U4210 (N_4210,N_3228,N_3583);
nand U4211 (N_4211,N_3803,N_3213);
nor U4212 (N_4212,N_3243,N_3614);
nand U4213 (N_4213,N_3662,N_3781);
or U4214 (N_4214,N_3738,N_3245);
nor U4215 (N_4215,N_3999,N_3611);
nand U4216 (N_4216,N_3404,N_3363);
and U4217 (N_4217,N_3597,N_3718);
or U4218 (N_4218,N_3464,N_3846);
xnor U4219 (N_4219,N_3459,N_3784);
nor U4220 (N_4220,N_3479,N_3896);
nor U4221 (N_4221,N_3731,N_3347);
xor U4222 (N_4222,N_3639,N_3417);
nand U4223 (N_4223,N_3396,N_3452);
nor U4224 (N_4224,N_3618,N_3204);
xor U4225 (N_4225,N_3752,N_3644);
and U4226 (N_4226,N_3995,N_3249);
and U4227 (N_4227,N_3699,N_3391);
nand U4228 (N_4228,N_3453,N_3805);
or U4229 (N_4229,N_3578,N_3711);
nor U4230 (N_4230,N_3368,N_3658);
nor U4231 (N_4231,N_3986,N_3500);
and U4232 (N_4232,N_3797,N_3663);
nor U4233 (N_4233,N_3930,N_3414);
nand U4234 (N_4234,N_3645,N_3924);
and U4235 (N_4235,N_3357,N_3625);
nand U4236 (N_4236,N_3951,N_3489);
nor U4237 (N_4237,N_3732,N_3211);
nand U4238 (N_4238,N_3328,N_3282);
nor U4239 (N_4239,N_3705,N_3716);
and U4240 (N_4240,N_3366,N_3234);
nor U4241 (N_4241,N_3601,N_3739);
and U4242 (N_4242,N_3340,N_3528);
nor U4243 (N_4243,N_3975,N_3861);
nor U4244 (N_4244,N_3222,N_3972);
and U4245 (N_4245,N_3446,N_3336);
nand U4246 (N_4246,N_3890,N_3491);
or U4247 (N_4247,N_3960,N_3443);
and U4248 (N_4248,N_3465,N_3510);
and U4249 (N_4249,N_3612,N_3383);
nor U4250 (N_4250,N_3755,N_3907);
or U4251 (N_4251,N_3281,N_3825);
and U4252 (N_4252,N_3508,N_3956);
xor U4253 (N_4253,N_3392,N_3901);
nor U4254 (N_4254,N_3393,N_3990);
nand U4255 (N_4255,N_3341,N_3201);
and U4256 (N_4256,N_3836,N_3325);
xor U4257 (N_4257,N_3927,N_3918);
xor U4258 (N_4258,N_3656,N_3409);
nand U4259 (N_4259,N_3206,N_3976);
nand U4260 (N_4260,N_3677,N_3314);
or U4261 (N_4261,N_3968,N_3767);
and U4262 (N_4262,N_3610,N_3702);
or U4263 (N_4263,N_3977,N_3884);
and U4264 (N_4264,N_3436,N_3253);
and U4265 (N_4265,N_3745,N_3657);
and U4266 (N_4266,N_3900,N_3793);
nor U4267 (N_4267,N_3205,N_3985);
nand U4268 (N_4268,N_3653,N_3531);
and U4269 (N_4269,N_3623,N_3786);
nor U4270 (N_4270,N_3429,N_3765);
nor U4271 (N_4271,N_3720,N_3251);
or U4272 (N_4272,N_3239,N_3697);
nor U4273 (N_4273,N_3838,N_3935);
nand U4274 (N_4274,N_3750,N_3220);
nor U4275 (N_4275,N_3435,N_3813);
nor U4276 (N_4276,N_3934,N_3332);
xor U4277 (N_4277,N_3576,N_3904);
and U4278 (N_4278,N_3882,N_3214);
xor U4279 (N_4279,N_3558,N_3305);
and U4280 (N_4280,N_3715,N_3887);
or U4281 (N_4281,N_3650,N_3487);
or U4282 (N_4282,N_3413,N_3883);
nor U4283 (N_4283,N_3674,N_3430);
xor U4284 (N_4284,N_3299,N_3571);
nand U4285 (N_4285,N_3817,N_3867);
xnor U4286 (N_4286,N_3843,N_3352);
and U4287 (N_4287,N_3523,N_3450);
nand U4288 (N_4288,N_3457,N_3778);
nand U4289 (N_4289,N_3964,N_3879);
xor U4290 (N_4290,N_3941,N_3868);
xor U4291 (N_4291,N_3604,N_3840);
nor U4292 (N_4292,N_3756,N_3367);
xor U4293 (N_4293,N_3310,N_3997);
nor U4294 (N_4294,N_3338,N_3757);
and U4295 (N_4295,N_3590,N_3869);
nand U4296 (N_4296,N_3659,N_3899);
and U4297 (N_4297,N_3785,N_3777);
and U4298 (N_4298,N_3595,N_3438);
xor U4299 (N_4299,N_3226,N_3277);
or U4300 (N_4300,N_3458,N_3408);
or U4301 (N_4301,N_3791,N_3600);
and U4302 (N_4302,N_3207,N_3472);
and U4303 (N_4303,N_3351,N_3759);
nand U4304 (N_4304,N_3892,N_3236);
or U4305 (N_4305,N_3664,N_3339);
or U4306 (N_4306,N_3542,N_3482);
and U4307 (N_4307,N_3527,N_3681);
xnor U4308 (N_4308,N_3322,N_3839);
and U4309 (N_4309,N_3947,N_3628);
nor U4310 (N_4310,N_3962,N_3726);
xnor U4311 (N_4311,N_3958,N_3671);
or U4312 (N_4312,N_3796,N_3327);
or U4313 (N_4313,N_3952,N_3532);
nand U4314 (N_4314,N_3672,N_3240);
xor U4315 (N_4315,N_3860,N_3728);
xor U4316 (N_4316,N_3557,N_3410);
xor U4317 (N_4317,N_3433,N_3912);
nand U4318 (N_4318,N_3584,N_3321);
or U4319 (N_4319,N_3379,N_3349);
xor U4320 (N_4320,N_3751,N_3737);
or U4321 (N_4321,N_3608,N_3284);
nor U4322 (N_4322,N_3560,N_3364);
nand U4323 (N_4323,N_3835,N_3648);
nand U4324 (N_4324,N_3686,N_3622);
nor U4325 (N_4325,N_3374,N_3782);
and U4326 (N_4326,N_3513,N_3263);
nand U4327 (N_4327,N_3543,N_3388);
xor U4328 (N_4328,N_3362,N_3358);
and U4329 (N_4329,N_3419,N_3412);
xor U4330 (N_4330,N_3886,N_3812);
or U4331 (N_4331,N_3473,N_3897);
nand U4332 (N_4332,N_3208,N_3945);
and U4333 (N_4333,N_3422,N_3541);
xnor U4334 (N_4334,N_3545,N_3828);
xor U4335 (N_4335,N_3857,N_3425);
and U4336 (N_4336,N_3474,N_3940);
xnor U4337 (N_4337,N_3844,N_3710);
nand U4338 (N_4338,N_3269,N_3559);
or U4339 (N_4339,N_3279,N_3973);
nand U4340 (N_4340,N_3690,N_3285);
or U4341 (N_4341,N_3342,N_3376);
and U4342 (N_4342,N_3637,N_3717);
nand U4343 (N_4343,N_3983,N_3494);
xor U4344 (N_4344,N_3740,N_3575);
and U4345 (N_4345,N_3678,N_3499);
nor U4346 (N_4346,N_3880,N_3602);
and U4347 (N_4347,N_3823,N_3565);
nand U4348 (N_4348,N_3209,N_3488);
or U4349 (N_4349,N_3696,N_3919);
and U4350 (N_4350,N_3714,N_3255);
and U4351 (N_4351,N_3706,N_3606);
nand U4352 (N_4352,N_3217,N_3698);
or U4353 (N_4353,N_3259,N_3955);
xor U4354 (N_4354,N_3832,N_3688);
nor U4355 (N_4355,N_3354,N_3633);
xor U4356 (N_4356,N_3359,N_3538);
xnor U4357 (N_4357,N_3747,N_3725);
and U4358 (N_4358,N_3223,N_3630);
nor U4359 (N_4359,N_3926,N_3949);
and U4360 (N_4360,N_3518,N_3561);
nand U4361 (N_4361,N_3307,N_3713);
or U4362 (N_4362,N_3978,N_3315);
nor U4363 (N_4363,N_3535,N_3552);
nor U4364 (N_4364,N_3283,N_3369);
or U4365 (N_4365,N_3554,N_3598);
nor U4366 (N_4366,N_3799,N_3449);
and U4367 (N_4367,N_3683,N_3914);
or U4368 (N_4368,N_3530,N_3428);
or U4369 (N_4369,N_3439,N_3455);
xor U4370 (N_4370,N_3440,N_3928);
and U4371 (N_4371,N_3244,N_3863);
or U4372 (N_4372,N_3624,N_3566);
and U4373 (N_4373,N_3830,N_3932);
xor U4374 (N_4374,N_3856,N_3319);
or U4375 (N_4375,N_3741,N_3794);
xnor U4376 (N_4376,N_3689,N_3744);
or U4377 (N_4377,N_3233,N_3456);
nor U4378 (N_4378,N_3382,N_3806);
and U4379 (N_4379,N_3309,N_3634);
nand U4380 (N_4380,N_3966,N_3974);
nand U4381 (N_4381,N_3300,N_3525);
or U4382 (N_4382,N_3898,N_3495);
and U4383 (N_4383,N_3421,N_3386);
or U4384 (N_4384,N_3746,N_3298);
nand U4385 (N_4385,N_3693,N_3232);
nand U4386 (N_4386,N_3712,N_3405);
xnor U4387 (N_4387,N_3942,N_3944);
or U4388 (N_4388,N_3445,N_3668);
nand U4389 (N_4389,N_3432,N_3615);
or U4390 (N_4390,N_3652,N_3866);
and U4391 (N_4391,N_3475,N_3701);
nand U4392 (N_4392,N_3329,N_3613);
and U4393 (N_4393,N_3800,N_3252);
and U4394 (N_4394,N_3819,N_3466);
nand U4395 (N_4395,N_3431,N_3742);
nor U4396 (N_4396,N_3323,N_3231);
or U4397 (N_4397,N_3268,N_3700);
or U4398 (N_4398,N_3989,N_3546);
nand U4399 (N_4399,N_3669,N_3271);
xor U4400 (N_4400,N_3772,N_3448);
nand U4401 (N_4401,N_3337,N_3918);
or U4402 (N_4402,N_3992,N_3438);
or U4403 (N_4403,N_3229,N_3283);
or U4404 (N_4404,N_3478,N_3676);
or U4405 (N_4405,N_3222,N_3753);
nand U4406 (N_4406,N_3469,N_3406);
or U4407 (N_4407,N_3948,N_3714);
nor U4408 (N_4408,N_3608,N_3851);
nand U4409 (N_4409,N_3958,N_3704);
and U4410 (N_4410,N_3861,N_3465);
xor U4411 (N_4411,N_3465,N_3753);
xor U4412 (N_4412,N_3694,N_3512);
and U4413 (N_4413,N_3853,N_3300);
or U4414 (N_4414,N_3505,N_3317);
xnor U4415 (N_4415,N_3495,N_3381);
xor U4416 (N_4416,N_3349,N_3747);
xor U4417 (N_4417,N_3676,N_3852);
nand U4418 (N_4418,N_3703,N_3901);
nor U4419 (N_4419,N_3292,N_3844);
or U4420 (N_4420,N_3360,N_3523);
and U4421 (N_4421,N_3938,N_3643);
xnor U4422 (N_4422,N_3945,N_3296);
xor U4423 (N_4423,N_3231,N_3414);
or U4424 (N_4424,N_3754,N_3663);
and U4425 (N_4425,N_3336,N_3813);
nand U4426 (N_4426,N_3988,N_3427);
or U4427 (N_4427,N_3718,N_3325);
and U4428 (N_4428,N_3881,N_3589);
and U4429 (N_4429,N_3541,N_3606);
nor U4430 (N_4430,N_3838,N_3405);
and U4431 (N_4431,N_3314,N_3356);
nand U4432 (N_4432,N_3421,N_3822);
nand U4433 (N_4433,N_3395,N_3758);
or U4434 (N_4434,N_3938,N_3577);
nand U4435 (N_4435,N_3933,N_3248);
xor U4436 (N_4436,N_3937,N_3265);
xnor U4437 (N_4437,N_3519,N_3814);
or U4438 (N_4438,N_3956,N_3746);
xor U4439 (N_4439,N_3450,N_3455);
or U4440 (N_4440,N_3211,N_3334);
nor U4441 (N_4441,N_3808,N_3621);
and U4442 (N_4442,N_3775,N_3883);
nand U4443 (N_4443,N_3333,N_3795);
xnor U4444 (N_4444,N_3703,N_3340);
or U4445 (N_4445,N_3791,N_3892);
or U4446 (N_4446,N_3840,N_3915);
and U4447 (N_4447,N_3787,N_3333);
and U4448 (N_4448,N_3518,N_3952);
nand U4449 (N_4449,N_3760,N_3981);
and U4450 (N_4450,N_3926,N_3811);
or U4451 (N_4451,N_3934,N_3552);
nor U4452 (N_4452,N_3847,N_3423);
xnor U4453 (N_4453,N_3737,N_3362);
xor U4454 (N_4454,N_3666,N_3617);
xnor U4455 (N_4455,N_3717,N_3550);
or U4456 (N_4456,N_3824,N_3889);
and U4457 (N_4457,N_3375,N_3568);
xor U4458 (N_4458,N_3853,N_3305);
or U4459 (N_4459,N_3234,N_3483);
and U4460 (N_4460,N_3401,N_3305);
nor U4461 (N_4461,N_3439,N_3828);
xnor U4462 (N_4462,N_3798,N_3767);
and U4463 (N_4463,N_3441,N_3503);
nor U4464 (N_4464,N_3779,N_3357);
xor U4465 (N_4465,N_3548,N_3343);
nor U4466 (N_4466,N_3592,N_3899);
and U4467 (N_4467,N_3338,N_3547);
xor U4468 (N_4468,N_3516,N_3858);
nand U4469 (N_4469,N_3542,N_3733);
or U4470 (N_4470,N_3993,N_3601);
or U4471 (N_4471,N_3773,N_3669);
xnor U4472 (N_4472,N_3425,N_3718);
or U4473 (N_4473,N_3704,N_3907);
or U4474 (N_4474,N_3406,N_3248);
and U4475 (N_4475,N_3617,N_3960);
nand U4476 (N_4476,N_3291,N_3897);
and U4477 (N_4477,N_3488,N_3256);
nand U4478 (N_4478,N_3659,N_3424);
nand U4479 (N_4479,N_3459,N_3763);
or U4480 (N_4480,N_3265,N_3491);
and U4481 (N_4481,N_3474,N_3801);
xor U4482 (N_4482,N_3252,N_3474);
nand U4483 (N_4483,N_3479,N_3834);
xnor U4484 (N_4484,N_3958,N_3353);
xnor U4485 (N_4485,N_3372,N_3307);
or U4486 (N_4486,N_3921,N_3698);
nand U4487 (N_4487,N_3367,N_3579);
or U4488 (N_4488,N_3499,N_3987);
and U4489 (N_4489,N_3416,N_3982);
or U4490 (N_4490,N_3247,N_3718);
and U4491 (N_4491,N_3759,N_3629);
xnor U4492 (N_4492,N_3786,N_3348);
xnor U4493 (N_4493,N_3797,N_3727);
xor U4494 (N_4494,N_3347,N_3922);
xor U4495 (N_4495,N_3357,N_3995);
and U4496 (N_4496,N_3513,N_3378);
xor U4497 (N_4497,N_3587,N_3575);
nor U4498 (N_4498,N_3306,N_3307);
or U4499 (N_4499,N_3440,N_3759);
nand U4500 (N_4500,N_3329,N_3555);
xnor U4501 (N_4501,N_3505,N_3227);
nor U4502 (N_4502,N_3641,N_3307);
nand U4503 (N_4503,N_3810,N_3748);
nand U4504 (N_4504,N_3818,N_3312);
or U4505 (N_4505,N_3508,N_3905);
nand U4506 (N_4506,N_3262,N_3537);
nor U4507 (N_4507,N_3217,N_3655);
nor U4508 (N_4508,N_3927,N_3362);
nor U4509 (N_4509,N_3264,N_3400);
nand U4510 (N_4510,N_3388,N_3971);
xor U4511 (N_4511,N_3547,N_3949);
xor U4512 (N_4512,N_3941,N_3957);
nor U4513 (N_4513,N_3539,N_3442);
and U4514 (N_4514,N_3292,N_3897);
and U4515 (N_4515,N_3542,N_3233);
nand U4516 (N_4516,N_3272,N_3961);
and U4517 (N_4517,N_3989,N_3484);
nand U4518 (N_4518,N_3379,N_3620);
or U4519 (N_4519,N_3842,N_3974);
nor U4520 (N_4520,N_3345,N_3431);
or U4521 (N_4521,N_3951,N_3490);
nor U4522 (N_4522,N_3529,N_3240);
nand U4523 (N_4523,N_3886,N_3331);
nor U4524 (N_4524,N_3464,N_3244);
xor U4525 (N_4525,N_3547,N_3567);
and U4526 (N_4526,N_3425,N_3841);
and U4527 (N_4527,N_3607,N_3478);
or U4528 (N_4528,N_3880,N_3610);
or U4529 (N_4529,N_3892,N_3209);
or U4530 (N_4530,N_3416,N_3949);
or U4531 (N_4531,N_3380,N_3921);
nand U4532 (N_4532,N_3937,N_3497);
xor U4533 (N_4533,N_3517,N_3684);
or U4534 (N_4534,N_3620,N_3604);
and U4535 (N_4535,N_3428,N_3386);
or U4536 (N_4536,N_3841,N_3837);
and U4537 (N_4537,N_3833,N_3372);
and U4538 (N_4538,N_3896,N_3315);
or U4539 (N_4539,N_3216,N_3504);
xnor U4540 (N_4540,N_3763,N_3886);
xnor U4541 (N_4541,N_3703,N_3255);
and U4542 (N_4542,N_3330,N_3823);
nand U4543 (N_4543,N_3459,N_3237);
and U4544 (N_4544,N_3544,N_3305);
and U4545 (N_4545,N_3283,N_3223);
nand U4546 (N_4546,N_3866,N_3715);
or U4547 (N_4547,N_3978,N_3421);
xor U4548 (N_4548,N_3504,N_3679);
xnor U4549 (N_4549,N_3928,N_3290);
or U4550 (N_4550,N_3981,N_3379);
and U4551 (N_4551,N_3847,N_3607);
or U4552 (N_4552,N_3757,N_3223);
nor U4553 (N_4553,N_3557,N_3405);
or U4554 (N_4554,N_3313,N_3591);
nand U4555 (N_4555,N_3531,N_3419);
nand U4556 (N_4556,N_3413,N_3438);
nand U4557 (N_4557,N_3363,N_3936);
nor U4558 (N_4558,N_3835,N_3554);
and U4559 (N_4559,N_3307,N_3313);
nand U4560 (N_4560,N_3968,N_3252);
nand U4561 (N_4561,N_3307,N_3341);
xor U4562 (N_4562,N_3362,N_3720);
nor U4563 (N_4563,N_3984,N_3609);
nor U4564 (N_4564,N_3317,N_3554);
nor U4565 (N_4565,N_3254,N_3770);
nand U4566 (N_4566,N_3242,N_3200);
xnor U4567 (N_4567,N_3918,N_3726);
nor U4568 (N_4568,N_3305,N_3217);
and U4569 (N_4569,N_3551,N_3564);
nand U4570 (N_4570,N_3773,N_3434);
xor U4571 (N_4571,N_3537,N_3553);
and U4572 (N_4572,N_3914,N_3921);
nor U4573 (N_4573,N_3663,N_3249);
nor U4574 (N_4574,N_3569,N_3312);
nor U4575 (N_4575,N_3345,N_3739);
xnor U4576 (N_4576,N_3285,N_3817);
or U4577 (N_4577,N_3525,N_3522);
xor U4578 (N_4578,N_3775,N_3318);
nor U4579 (N_4579,N_3397,N_3882);
nor U4580 (N_4580,N_3520,N_3539);
xnor U4581 (N_4581,N_3891,N_3374);
nor U4582 (N_4582,N_3279,N_3841);
nand U4583 (N_4583,N_3342,N_3903);
and U4584 (N_4584,N_3418,N_3509);
and U4585 (N_4585,N_3625,N_3364);
and U4586 (N_4586,N_3735,N_3390);
nor U4587 (N_4587,N_3210,N_3921);
and U4588 (N_4588,N_3746,N_3918);
nor U4589 (N_4589,N_3507,N_3397);
and U4590 (N_4590,N_3871,N_3837);
nor U4591 (N_4591,N_3310,N_3790);
and U4592 (N_4592,N_3708,N_3591);
or U4593 (N_4593,N_3893,N_3720);
and U4594 (N_4594,N_3594,N_3385);
nor U4595 (N_4595,N_3528,N_3201);
xnor U4596 (N_4596,N_3315,N_3204);
nor U4597 (N_4597,N_3830,N_3898);
nand U4598 (N_4598,N_3812,N_3361);
or U4599 (N_4599,N_3607,N_3390);
and U4600 (N_4600,N_3943,N_3239);
xnor U4601 (N_4601,N_3344,N_3932);
xor U4602 (N_4602,N_3330,N_3770);
xor U4603 (N_4603,N_3256,N_3586);
or U4604 (N_4604,N_3660,N_3895);
nand U4605 (N_4605,N_3878,N_3314);
and U4606 (N_4606,N_3509,N_3622);
nand U4607 (N_4607,N_3849,N_3688);
xnor U4608 (N_4608,N_3345,N_3246);
nor U4609 (N_4609,N_3778,N_3746);
and U4610 (N_4610,N_3710,N_3564);
nor U4611 (N_4611,N_3507,N_3711);
xnor U4612 (N_4612,N_3574,N_3554);
and U4613 (N_4613,N_3516,N_3215);
nand U4614 (N_4614,N_3321,N_3959);
and U4615 (N_4615,N_3436,N_3878);
or U4616 (N_4616,N_3589,N_3530);
nor U4617 (N_4617,N_3919,N_3537);
xnor U4618 (N_4618,N_3299,N_3368);
nand U4619 (N_4619,N_3714,N_3691);
nor U4620 (N_4620,N_3811,N_3667);
nor U4621 (N_4621,N_3245,N_3959);
xnor U4622 (N_4622,N_3574,N_3873);
nor U4623 (N_4623,N_3573,N_3567);
and U4624 (N_4624,N_3260,N_3492);
nor U4625 (N_4625,N_3904,N_3531);
nor U4626 (N_4626,N_3456,N_3701);
nand U4627 (N_4627,N_3551,N_3597);
or U4628 (N_4628,N_3619,N_3832);
or U4629 (N_4629,N_3512,N_3422);
and U4630 (N_4630,N_3819,N_3511);
xor U4631 (N_4631,N_3437,N_3560);
xor U4632 (N_4632,N_3382,N_3802);
or U4633 (N_4633,N_3665,N_3780);
xor U4634 (N_4634,N_3520,N_3402);
xor U4635 (N_4635,N_3391,N_3989);
or U4636 (N_4636,N_3551,N_3728);
xnor U4637 (N_4637,N_3564,N_3991);
or U4638 (N_4638,N_3937,N_3972);
nand U4639 (N_4639,N_3331,N_3775);
nor U4640 (N_4640,N_3547,N_3488);
xor U4641 (N_4641,N_3432,N_3400);
nand U4642 (N_4642,N_3918,N_3842);
or U4643 (N_4643,N_3712,N_3699);
and U4644 (N_4644,N_3465,N_3748);
nand U4645 (N_4645,N_3497,N_3501);
or U4646 (N_4646,N_3343,N_3512);
xor U4647 (N_4647,N_3620,N_3628);
nand U4648 (N_4648,N_3799,N_3286);
xnor U4649 (N_4649,N_3804,N_3662);
or U4650 (N_4650,N_3840,N_3650);
or U4651 (N_4651,N_3978,N_3910);
nand U4652 (N_4652,N_3354,N_3863);
and U4653 (N_4653,N_3702,N_3542);
nand U4654 (N_4654,N_3524,N_3776);
nor U4655 (N_4655,N_3553,N_3278);
and U4656 (N_4656,N_3786,N_3353);
nor U4657 (N_4657,N_3408,N_3788);
nor U4658 (N_4658,N_3569,N_3641);
or U4659 (N_4659,N_3962,N_3786);
nor U4660 (N_4660,N_3846,N_3759);
nand U4661 (N_4661,N_3653,N_3219);
nor U4662 (N_4662,N_3223,N_3440);
nand U4663 (N_4663,N_3339,N_3202);
nor U4664 (N_4664,N_3624,N_3750);
nand U4665 (N_4665,N_3540,N_3993);
or U4666 (N_4666,N_3855,N_3381);
and U4667 (N_4667,N_3920,N_3919);
nand U4668 (N_4668,N_3492,N_3298);
or U4669 (N_4669,N_3914,N_3449);
nor U4670 (N_4670,N_3938,N_3892);
xor U4671 (N_4671,N_3695,N_3550);
or U4672 (N_4672,N_3913,N_3229);
nor U4673 (N_4673,N_3751,N_3428);
xnor U4674 (N_4674,N_3280,N_3618);
nor U4675 (N_4675,N_3395,N_3270);
and U4676 (N_4676,N_3248,N_3695);
xnor U4677 (N_4677,N_3657,N_3571);
or U4678 (N_4678,N_3819,N_3330);
and U4679 (N_4679,N_3472,N_3895);
or U4680 (N_4680,N_3951,N_3674);
nand U4681 (N_4681,N_3234,N_3744);
nor U4682 (N_4682,N_3662,N_3784);
nand U4683 (N_4683,N_3200,N_3380);
nand U4684 (N_4684,N_3243,N_3709);
or U4685 (N_4685,N_3989,N_3597);
and U4686 (N_4686,N_3864,N_3416);
xnor U4687 (N_4687,N_3706,N_3809);
nand U4688 (N_4688,N_3517,N_3537);
xor U4689 (N_4689,N_3512,N_3886);
xnor U4690 (N_4690,N_3793,N_3702);
or U4691 (N_4691,N_3244,N_3352);
nand U4692 (N_4692,N_3377,N_3933);
nor U4693 (N_4693,N_3877,N_3437);
nand U4694 (N_4694,N_3513,N_3987);
and U4695 (N_4695,N_3803,N_3860);
nand U4696 (N_4696,N_3570,N_3964);
nor U4697 (N_4697,N_3202,N_3535);
xnor U4698 (N_4698,N_3319,N_3614);
or U4699 (N_4699,N_3549,N_3552);
and U4700 (N_4700,N_3727,N_3866);
xor U4701 (N_4701,N_3207,N_3960);
nor U4702 (N_4702,N_3623,N_3579);
and U4703 (N_4703,N_3995,N_3305);
nor U4704 (N_4704,N_3919,N_3425);
or U4705 (N_4705,N_3531,N_3451);
nand U4706 (N_4706,N_3905,N_3521);
or U4707 (N_4707,N_3474,N_3425);
or U4708 (N_4708,N_3970,N_3843);
nor U4709 (N_4709,N_3818,N_3823);
nor U4710 (N_4710,N_3915,N_3644);
nand U4711 (N_4711,N_3262,N_3531);
or U4712 (N_4712,N_3572,N_3451);
and U4713 (N_4713,N_3921,N_3306);
nand U4714 (N_4714,N_3907,N_3638);
or U4715 (N_4715,N_3928,N_3306);
or U4716 (N_4716,N_3381,N_3281);
and U4717 (N_4717,N_3883,N_3754);
nand U4718 (N_4718,N_3538,N_3218);
and U4719 (N_4719,N_3909,N_3846);
nand U4720 (N_4720,N_3400,N_3374);
nand U4721 (N_4721,N_3696,N_3863);
xor U4722 (N_4722,N_3513,N_3634);
and U4723 (N_4723,N_3580,N_3213);
xor U4724 (N_4724,N_3445,N_3636);
xor U4725 (N_4725,N_3392,N_3488);
nand U4726 (N_4726,N_3789,N_3818);
xnor U4727 (N_4727,N_3692,N_3668);
nand U4728 (N_4728,N_3583,N_3341);
nor U4729 (N_4729,N_3467,N_3863);
or U4730 (N_4730,N_3647,N_3736);
nand U4731 (N_4731,N_3722,N_3703);
or U4732 (N_4732,N_3637,N_3779);
and U4733 (N_4733,N_3646,N_3430);
xnor U4734 (N_4734,N_3636,N_3686);
nand U4735 (N_4735,N_3453,N_3215);
xnor U4736 (N_4736,N_3642,N_3420);
or U4737 (N_4737,N_3230,N_3663);
nor U4738 (N_4738,N_3479,N_3795);
nor U4739 (N_4739,N_3260,N_3379);
or U4740 (N_4740,N_3237,N_3663);
nand U4741 (N_4741,N_3860,N_3254);
nor U4742 (N_4742,N_3413,N_3532);
xor U4743 (N_4743,N_3782,N_3251);
and U4744 (N_4744,N_3480,N_3640);
or U4745 (N_4745,N_3633,N_3422);
nor U4746 (N_4746,N_3389,N_3745);
nand U4747 (N_4747,N_3310,N_3569);
xnor U4748 (N_4748,N_3880,N_3356);
nand U4749 (N_4749,N_3873,N_3488);
nand U4750 (N_4750,N_3256,N_3304);
and U4751 (N_4751,N_3622,N_3573);
or U4752 (N_4752,N_3411,N_3281);
nor U4753 (N_4753,N_3834,N_3922);
or U4754 (N_4754,N_3477,N_3881);
or U4755 (N_4755,N_3265,N_3916);
xor U4756 (N_4756,N_3971,N_3496);
xor U4757 (N_4757,N_3232,N_3835);
and U4758 (N_4758,N_3553,N_3979);
and U4759 (N_4759,N_3972,N_3966);
nand U4760 (N_4760,N_3829,N_3553);
nand U4761 (N_4761,N_3227,N_3794);
and U4762 (N_4762,N_3425,N_3546);
and U4763 (N_4763,N_3955,N_3865);
nor U4764 (N_4764,N_3668,N_3405);
and U4765 (N_4765,N_3270,N_3373);
or U4766 (N_4766,N_3892,N_3288);
and U4767 (N_4767,N_3436,N_3371);
or U4768 (N_4768,N_3495,N_3735);
and U4769 (N_4769,N_3632,N_3301);
and U4770 (N_4770,N_3496,N_3800);
nor U4771 (N_4771,N_3430,N_3890);
nand U4772 (N_4772,N_3730,N_3202);
xnor U4773 (N_4773,N_3802,N_3219);
or U4774 (N_4774,N_3258,N_3657);
xor U4775 (N_4775,N_3675,N_3503);
xor U4776 (N_4776,N_3785,N_3391);
or U4777 (N_4777,N_3975,N_3852);
xnor U4778 (N_4778,N_3727,N_3219);
nor U4779 (N_4779,N_3890,N_3217);
xor U4780 (N_4780,N_3318,N_3651);
xnor U4781 (N_4781,N_3821,N_3927);
xor U4782 (N_4782,N_3614,N_3502);
xnor U4783 (N_4783,N_3289,N_3654);
or U4784 (N_4784,N_3892,N_3690);
nand U4785 (N_4785,N_3824,N_3328);
nor U4786 (N_4786,N_3484,N_3977);
and U4787 (N_4787,N_3508,N_3399);
or U4788 (N_4788,N_3648,N_3321);
or U4789 (N_4789,N_3255,N_3793);
and U4790 (N_4790,N_3557,N_3584);
or U4791 (N_4791,N_3638,N_3633);
nor U4792 (N_4792,N_3382,N_3429);
nand U4793 (N_4793,N_3355,N_3970);
and U4794 (N_4794,N_3862,N_3622);
and U4795 (N_4795,N_3341,N_3323);
nand U4796 (N_4796,N_3918,N_3229);
nand U4797 (N_4797,N_3477,N_3450);
nand U4798 (N_4798,N_3330,N_3524);
xor U4799 (N_4799,N_3916,N_3980);
or U4800 (N_4800,N_4612,N_4199);
xnor U4801 (N_4801,N_4773,N_4243);
nor U4802 (N_4802,N_4033,N_4477);
nor U4803 (N_4803,N_4577,N_4781);
nor U4804 (N_4804,N_4466,N_4203);
and U4805 (N_4805,N_4427,N_4710);
nand U4806 (N_4806,N_4077,N_4788);
nand U4807 (N_4807,N_4759,N_4433);
xnor U4808 (N_4808,N_4723,N_4019);
nor U4809 (N_4809,N_4499,N_4233);
nand U4810 (N_4810,N_4753,N_4298);
or U4811 (N_4811,N_4695,N_4430);
nor U4812 (N_4812,N_4587,N_4259);
nand U4813 (N_4813,N_4217,N_4755);
and U4814 (N_4814,N_4315,N_4656);
or U4815 (N_4815,N_4646,N_4197);
and U4816 (N_4816,N_4664,N_4678);
or U4817 (N_4817,N_4729,N_4647);
nand U4818 (N_4818,N_4650,N_4031);
and U4819 (N_4819,N_4631,N_4201);
xnor U4820 (N_4820,N_4257,N_4188);
or U4821 (N_4821,N_4321,N_4114);
or U4822 (N_4822,N_4744,N_4046);
nor U4823 (N_4823,N_4281,N_4293);
and U4824 (N_4824,N_4408,N_4790);
or U4825 (N_4825,N_4275,N_4718);
or U4826 (N_4826,N_4540,N_4441);
nor U4827 (N_4827,N_4464,N_4052);
nand U4828 (N_4828,N_4276,N_4121);
and U4829 (N_4829,N_4796,N_4093);
xor U4830 (N_4830,N_4683,N_4342);
and U4831 (N_4831,N_4245,N_4359);
xnor U4832 (N_4832,N_4267,N_4367);
and U4833 (N_4833,N_4063,N_4600);
nor U4834 (N_4834,N_4331,N_4344);
nor U4835 (N_4835,N_4286,N_4487);
nand U4836 (N_4836,N_4159,N_4674);
xnor U4837 (N_4837,N_4072,N_4055);
or U4838 (N_4838,N_4546,N_4282);
and U4839 (N_4839,N_4122,N_4409);
or U4840 (N_4840,N_4137,N_4749);
nand U4841 (N_4841,N_4352,N_4307);
nor U4842 (N_4842,N_4630,N_4395);
nor U4843 (N_4843,N_4028,N_4598);
nand U4844 (N_4844,N_4016,N_4642);
nor U4845 (N_4845,N_4071,N_4009);
and U4846 (N_4846,N_4629,N_4156);
nand U4847 (N_4847,N_4239,N_4128);
or U4848 (N_4848,N_4453,N_4424);
and U4849 (N_4849,N_4020,N_4023);
nor U4850 (N_4850,N_4608,N_4509);
nand U4851 (N_4851,N_4003,N_4238);
xnor U4852 (N_4852,N_4372,N_4682);
and U4853 (N_4853,N_4732,N_4092);
nand U4854 (N_4854,N_4722,N_4295);
nor U4855 (N_4855,N_4035,N_4136);
or U4856 (N_4856,N_4076,N_4689);
and U4857 (N_4857,N_4628,N_4615);
or U4858 (N_4858,N_4731,N_4292);
nand U4859 (N_4859,N_4541,N_4780);
xor U4860 (N_4860,N_4442,N_4459);
nor U4861 (N_4861,N_4772,N_4601);
xor U4862 (N_4862,N_4445,N_4620);
xnor U4863 (N_4863,N_4090,N_4480);
xor U4864 (N_4864,N_4054,N_4719);
and U4865 (N_4865,N_4235,N_4613);
nand U4866 (N_4866,N_4524,N_4658);
xnor U4867 (N_4867,N_4701,N_4460);
xnor U4868 (N_4868,N_4747,N_4189);
xnor U4869 (N_4869,N_4446,N_4696);
xnor U4870 (N_4870,N_4703,N_4576);
and U4871 (N_4871,N_4345,N_4301);
and U4872 (N_4872,N_4638,N_4061);
or U4873 (N_4873,N_4335,N_4109);
or U4874 (N_4874,N_4145,N_4230);
or U4875 (N_4875,N_4225,N_4554);
and U4876 (N_4876,N_4380,N_4212);
xnor U4877 (N_4877,N_4505,N_4171);
or U4878 (N_4878,N_4706,N_4049);
and U4879 (N_4879,N_4165,N_4488);
nor U4880 (N_4880,N_4669,N_4462);
nor U4881 (N_4881,N_4324,N_4490);
and U4882 (N_4882,N_4566,N_4727);
nor U4883 (N_4883,N_4017,N_4178);
or U4884 (N_4884,N_4786,N_4572);
xnor U4885 (N_4885,N_4585,N_4044);
and U4886 (N_4886,N_4139,N_4338);
and U4887 (N_4887,N_4556,N_4096);
and U4888 (N_4888,N_4391,N_4024);
or U4889 (N_4889,N_4222,N_4497);
and U4890 (N_4890,N_4565,N_4758);
nand U4891 (N_4891,N_4712,N_4116);
and U4892 (N_4892,N_4508,N_4339);
and U4893 (N_4893,N_4356,N_4680);
xor U4894 (N_4894,N_4132,N_4725);
and U4895 (N_4895,N_4303,N_4370);
xnor U4896 (N_4896,N_4070,N_4036);
nand U4897 (N_4897,N_4570,N_4147);
and U4898 (N_4898,N_4495,N_4213);
nand U4899 (N_4899,N_4632,N_4143);
nand U4900 (N_4900,N_4089,N_4179);
nand U4901 (N_4901,N_4604,N_4691);
xor U4902 (N_4902,N_4580,N_4468);
xnor U4903 (N_4903,N_4368,N_4603);
and U4904 (N_4904,N_4038,N_4493);
nand U4905 (N_4905,N_4551,N_4622);
xnor U4906 (N_4906,N_4518,N_4310);
nand U4907 (N_4907,N_4062,N_4764);
or U4908 (N_4908,N_4422,N_4265);
xnor U4909 (N_4909,N_4347,N_4426);
nand U4910 (N_4910,N_4101,N_4205);
and U4911 (N_4911,N_4685,N_4249);
and U4912 (N_4912,N_4672,N_4140);
nor U4913 (N_4913,N_4154,N_4216);
or U4914 (N_4914,N_4264,N_4660);
nand U4915 (N_4915,N_4389,N_4511);
or U4916 (N_4916,N_4746,N_4714);
xnor U4917 (N_4917,N_4254,N_4045);
or U4918 (N_4918,N_4597,N_4506);
xor U4919 (N_4919,N_4482,N_4724);
nand U4920 (N_4920,N_4760,N_4256);
nor U4921 (N_4921,N_4507,N_4221);
xnor U4922 (N_4922,N_4373,N_4717);
nor U4923 (N_4923,N_4514,N_4534);
nor U4924 (N_4924,N_4381,N_4625);
nor U4925 (N_4925,N_4416,N_4590);
or U4926 (N_4926,N_4400,N_4065);
xor U4927 (N_4927,N_4793,N_4353);
and U4928 (N_4928,N_4011,N_4519);
and U4929 (N_4929,N_4473,N_4237);
and U4930 (N_4930,N_4313,N_4283);
or U4931 (N_4931,N_4255,N_4207);
nor U4932 (N_4932,N_4176,N_4361);
and U4933 (N_4933,N_4358,N_4730);
nor U4934 (N_4934,N_4053,N_4387);
nor U4935 (N_4935,N_4162,N_4716);
nand U4936 (N_4936,N_4513,N_4005);
nor U4937 (N_4937,N_4209,N_4619);
and U4938 (N_4938,N_4690,N_4439);
or U4939 (N_4939,N_4574,N_4081);
xor U4940 (N_4940,N_4336,N_4104);
xnor U4941 (N_4941,N_4571,N_4633);
and U4942 (N_4942,N_4640,N_4402);
xor U4943 (N_4943,N_4304,N_4153);
xnor U4944 (N_4944,N_4795,N_4504);
nor U4945 (N_4945,N_4227,N_4299);
xnor U4946 (N_4946,N_4302,N_4611);
or U4947 (N_4947,N_4797,N_4210);
nor U4948 (N_4948,N_4268,N_4688);
or U4949 (N_4949,N_4425,N_4787);
xor U4950 (N_4950,N_4148,N_4414);
nor U4951 (N_4951,N_4327,N_4548);
nor U4952 (N_4952,N_4393,N_4328);
and U4953 (N_4953,N_4659,N_4325);
nand U4954 (N_4954,N_4637,N_4332);
and U4955 (N_4955,N_4311,N_4700);
or U4956 (N_4956,N_4407,N_4306);
and U4957 (N_4957,N_4384,N_4419);
and U4958 (N_4958,N_4261,N_4799);
and U4959 (N_4959,N_4341,N_4467);
nand U4960 (N_4960,N_4609,N_4421);
nor U4961 (N_4961,N_4269,N_4048);
and U4962 (N_4962,N_4248,N_4056);
or U4963 (N_4963,N_4146,N_4501);
xor U4964 (N_4964,N_4666,N_4523);
and U4965 (N_4965,N_4447,N_4599);
xnor U4966 (N_4966,N_4641,N_4605);
or U4967 (N_4967,N_4349,N_4174);
and U4968 (N_4968,N_4007,N_4051);
xor U4969 (N_4969,N_4364,N_4343);
or U4970 (N_4970,N_4300,N_4115);
and U4971 (N_4971,N_4451,N_4698);
nor U4972 (N_4972,N_4596,N_4192);
and U4973 (N_4973,N_4649,N_4142);
nor U4974 (N_4974,N_4095,N_4726);
and U4975 (N_4975,N_4607,N_4757);
nand U4976 (N_4976,N_4340,N_4777);
or U4977 (N_4977,N_4280,N_4308);
nand U4978 (N_4978,N_4713,N_4151);
nand U4979 (N_4979,N_4317,N_4778);
nand U4980 (N_4980,N_4274,N_4454);
nand U4981 (N_4981,N_4774,N_4060);
and U4982 (N_4982,N_4120,N_4242);
and U4983 (N_4983,N_4091,N_4110);
or U4984 (N_4984,N_4234,N_4316);
and U4985 (N_4985,N_4521,N_4403);
nor U4986 (N_4986,N_4294,N_4030);
or U4987 (N_4987,N_4705,N_4258);
or U4988 (N_4988,N_4461,N_4652);
nand U4989 (N_4989,N_4405,N_4751);
and U4990 (N_4990,N_4512,N_4648);
or U4991 (N_4991,N_4436,N_4180);
and U4992 (N_4992,N_4043,N_4623);
xnor U4993 (N_4993,N_4643,N_4172);
or U4994 (N_4994,N_4410,N_4522);
nor U4995 (N_4995,N_4173,N_4186);
and U4996 (N_4996,N_4247,N_4510);
nand U4997 (N_4997,N_4569,N_4135);
xnor U4998 (N_4998,N_4218,N_4476);
nand U4999 (N_4999,N_4278,N_4626);
xor U5000 (N_5000,N_4157,N_4457);
nor U5001 (N_5001,N_4170,N_4677);
or U5002 (N_5002,N_4675,N_4769);
and U5003 (N_5003,N_4369,N_4699);
xnor U5004 (N_5004,N_4078,N_4579);
or U5005 (N_5005,N_4697,N_4141);
or U5006 (N_5006,N_4206,N_4333);
nand U5007 (N_5007,N_4588,N_4397);
nor U5008 (N_5008,N_4776,N_4066);
nor U5009 (N_5009,N_4635,N_4745);
nand U5010 (N_5010,N_4037,N_4232);
xor U5011 (N_5011,N_4022,N_4553);
xnor U5012 (N_5012,N_4117,N_4767);
nand U5013 (N_5013,N_4102,N_4074);
xor U5014 (N_5014,N_4709,N_4775);
and U5015 (N_5015,N_4578,N_4472);
nand U5016 (N_5016,N_4195,N_4584);
or U5017 (N_5017,N_4411,N_4443);
and U5018 (N_5018,N_4015,N_4431);
nand U5019 (N_5019,N_4485,N_4039);
xnor U5020 (N_5020,N_4515,N_4164);
and U5021 (N_5021,N_4083,N_4272);
nand U5022 (N_5022,N_4483,N_4214);
and U5023 (N_5023,N_4766,N_4193);
xnor U5024 (N_5024,N_4555,N_4069);
nor U5025 (N_5025,N_4527,N_4657);
nand U5026 (N_5026,N_4444,N_4144);
nand U5027 (N_5027,N_4099,N_4525);
or U5028 (N_5028,N_4094,N_4073);
nor U5029 (N_5029,N_4562,N_4549);
nor U5030 (N_5030,N_4768,N_4394);
or U5031 (N_5031,N_4219,N_4413);
nor U5032 (N_5032,N_4183,N_4754);
and U5033 (N_5033,N_4792,N_4463);
nand U5034 (N_5034,N_4449,N_4079);
nor U5035 (N_5035,N_4720,N_4329);
and U5036 (N_5036,N_4177,N_4624);
xnor U5037 (N_5037,N_4671,N_4517);
xor U5038 (N_5038,N_4783,N_4437);
nor U5039 (N_5039,N_4377,N_4564);
nand U5040 (N_5040,N_4531,N_4244);
and U5041 (N_5041,N_4130,N_4455);
or U5042 (N_5042,N_4415,N_4103);
nor U5043 (N_5043,N_4082,N_4251);
and U5044 (N_5044,N_4398,N_4296);
or U5045 (N_5045,N_4516,N_4004);
nor U5046 (N_5046,N_4406,N_4494);
nor U5047 (N_5047,N_4105,N_4655);
nor U5048 (N_5048,N_4175,N_4042);
nor U5049 (N_5049,N_4636,N_4289);
xor U5050 (N_5050,N_4779,N_4547);
nor U5051 (N_5051,N_4050,N_4610);
nand U5052 (N_5052,N_4673,N_4000);
and U5053 (N_5053,N_4423,N_4360);
nor U5054 (N_5054,N_4417,N_4676);
nor U5055 (N_5055,N_4595,N_4558);
nand U5056 (N_5056,N_4502,N_4404);
nand U5057 (N_5057,N_4752,N_4492);
and U5058 (N_5058,N_4435,N_4704);
nand U5059 (N_5059,N_4229,N_4450);
or U5060 (N_5060,N_4583,N_4593);
nand U5061 (N_5061,N_4080,N_4644);
or U5062 (N_5062,N_4667,N_4252);
nand U5063 (N_5063,N_4182,N_4125);
nand U5064 (N_5064,N_4215,N_4582);
nor U5065 (N_5065,N_4702,N_4594);
nor U5066 (N_5066,N_4618,N_4058);
xnor U5067 (N_5067,N_4190,N_4001);
xor U5068 (N_5068,N_4026,N_4496);
xor U5069 (N_5069,N_4277,N_4167);
nor U5070 (N_5070,N_4168,N_4385);
nand U5071 (N_5071,N_4160,N_4376);
or U5072 (N_5072,N_4651,N_4663);
and U5073 (N_5073,N_4288,N_4305);
nand U5074 (N_5074,N_4012,N_4013);
or U5075 (N_5075,N_4545,N_4412);
xor U5076 (N_5076,N_4375,N_4715);
and U5077 (N_5077,N_4085,N_4694);
and U5078 (N_5078,N_4084,N_4112);
or U5079 (N_5079,N_4040,N_4337);
xnor U5080 (N_5080,N_4390,N_4543);
or U5081 (N_5081,N_4149,N_4763);
nor U5082 (N_5082,N_4668,N_4771);
nor U5083 (N_5083,N_4432,N_4756);
or U5084 (N_5084,N_4196,N_4791);
and U5085 (N_5085,N_4616,N_4348);
nor U5086 (N_5086,N_4434,N_4319);
and U5087 (N_5087,N_4320,N_4204);
or U5088 (N_5088,N_4470,N_4191);
nand U5089 (N_5089,N_4351,N_4231);
xor U5090 (N_5090,N_4498,N_4479);
xnor U5091 (N_5091,N_4386,N_4284);
nor U5092 (N_5092,N_4575,N_4323);
and U5093 (N_5093,N_4378,N_4542);
xnor U5094 (N_5094,N_4163,N_4529);
nand U5095 (N_5095,N_4737,N_4489);
xnor U5096 (N_5096,N_4010,N_4067);
or U5097 (N_5097,N_4382,N_4246);
nand U5098 (N_5098,N_4532,N_4365);
nand U5099 (N_5099,N_4208,N_4739);
or U5100 (N_5100,N_4735,N_4187);
nand U5101 (N_5101,N_4106,N_4029);
and U5102 (N_5102,N_4263,N_4330);
nor U5103 (N_5103,N_4291,N_4322);
nor U5104 (N_5104,N_4111,N_4097);
xor U5105 (N_5105,N_4526,N_4075);
and U5106 (N_5106,N_4262,N_4138);
nand U5107 (N_5107,N_4544,N_4784);
and U5108 (N_5108,N_4032,N_4500);
nand U5109 (N_5109,N_4537,N_4059);
and U5110 (N_5110,N_4133,N_4350);
and U5111 (N_5111,N_4550,N_4270);
or U5112 (N_5112,N_4158,N_4363);
nand U5113 (N_5113,N_4484,N_4503);
xnor U5114 (N_5114,N_4670,N_4679);
or U5115 (N_5115,N_4456,N_4150);
nor U5116 (N_5116,N_4169,N_4355);
and U5117 (N_5117,N_4279,N_4686);
xnor U5118 (N_5118,N_4568,N_4220);
or U5119 (N_5119,N_4374,N_4662);
nor U5120 (N_5120,N_4458,N_4018);
or U5121 (N_5121,N_4765,N_4741);
nor U5122 (N_5122,N_4559,N_4354);
and U5123 (N_5123,N_4736,N_4692);
nor U5124 (N_5124,N_4728,N_4021);
and U5125 (N_5125,N_4557,N_4057);
or U5126 (N_5126,N_4086,N_4606);
xor U5127 (N_5127,N_4383,N_4014);
nand U5128 (N_5128,N_4334,N_4440);
xor U5129 (N_5129,N_4124,N_4491);
and U5130 (N_5130,N_4236,N_4185);
nor U5131 (N_5131,N_4474,N_4748);
or U5132 (N_5132,N_4738,N_4379);
and U5133 (N_5133,N_4762,N_4181);
and U5134 (N_5134,N_4366,N_4155);
and U5135 (N_5135,N_4734,N_4047);
nor U5136 (N_5136,N_4194,N_4100);
nor U5137 (N_5137,N_4260,N_4027);
xnor U5138 (N_5138,N_4312,N_4127);
or U5139 (N_5139,N_4761,N_4687);
xor U5140 (N_5140,N_4740,N_4708);
nand U5141 (N_5141,N_4614,N_4743);
and U5142 (N_5142,N_4253,N_4271);
nor U5143 (N_5143,N_4224,N_4538);
or U5144 (N_5144,N_4589,N_4418);
nor U5145 (N_5145,N_4429,N_4123);
nand U5146 (N_5146,N_4025,N_4008);
xnor U5147 (N_5147,N_4362,N_4126);
and U5148 (N_5148,N_4287,N_4627);
and U5149 (N_5149,N_4399,N_4707);
nor U5150 (N_5150,N_4087,N_4634);
xor U5151 (N_5151,N_4034,N_4166);
xor U5152 (N_5152,N_4733,N_4693);
nor U5153 (N_5153,N_4285,N_4346);
nor U5154 (N_5154,N_4581,N_4563);
or U5155 (N_5155,N_4586,N_4684);
and U5156 (N_5156,N_4198,N_4661);
nand U5157 (N_5157,N_4520,N_4107);
and U5158 (N_5158,N_4721,N_4420);
and U5159 (N_5159,N_4592,N_4002);
xnor U5160 (N_5160,N_4645,N_4131);
xor U5161 (N_5161,N_4223,N_4152);
nand U5162 (N_5162,N_4161,N_4118);
or U5163 (N_5163,N_4471,N_4465);
nand U5164 (N_5164,N_4535,N_4654);
and U5165 (N_5165,N_4357,N_4481);
or U5166 (N_5166,N_4770,N_4475);
nand U5167 (N_5167,N_4639,N_4200);
and U5168 (N_5168,N_4438,N_4567);
or U5169 (N_5169,N_4392,N_4241);
nor U5170 (N_5170,N_4088,N_4552);
xnor U5171 (N_5171,N_4533,N_4266);
and U5172 (N_5172,N_4396,N_4560);
nand U5173 (N_5173,N_4309,N_4113);
xnor U5174 (N_5174,N_4448,N_4064);
or U5175 (N_5175,N_4602,N_4250);
nand U5176 (N_5176,N_4108,N_4314);
nor U5177 (N_5177,N_4530,N_4665);
or U5178 (N_5178,N_4528,N_4798);
nand U5179 (N_5179,N_4068,N_4536);
xnor U5180 (N_5180,N_4539,N_4273);
and U5181 (N_5181,N_4202,N_4318);
xor U5182 (N_5182,N_4134,N_4478);
nand U5183 (N_5183,N_4388,N_4617);
nand U5184 (N_5184,N_4401,N_4785);
or U5185 (N_5185,N_4119,N_4211);
or U5186 (N_5186,N_4452,N_4184);
nor U5187 (N_5187,N_4782,N_4240);
nor U5188 (N_5188,N_4653,N_4711);
and U5189 (N_5189,N_4750,N_4226);
nor U5190 (N_5190,N_4228,N_4326);
nand U5191 (N_5191,N_4681,N_4041);
nand U5192 (N_5192,N_4006,N_4789);
or U5193 (N_5193,N_4621,N_4742);
nor U5194 (N_5194,N_4129,N_4486);
nand U5195 (N_5195,N_4290,N_4573);
nand U5196 (N_5196,N_4371,N_4469);
and U5197 (N_5197,N_4561,N_4098);
and U5198 (N_5198,N_4794,N_4297);
nor U5199 (N_5199,N_4591,N_4428);
xnor U5200 (N_5200,N_4244,N_4527);
nand U5201 (N_5201,N_4583,N_4301);
nand U5202 (N_5202,N_4429,N_4366);
nand U5203 (N_5203,N_4607,N_4736);
nand U5204 (N_5204,N_4629,N_4437);
nand U5205 (N_5205,N_4142,N_4755);
nand U5206 (N_5206,N_4780,N_4149);
and U5207 (N_5207,N_4296,N_4484);
and U5208 (N_5208,N_4563,N_4493);
and U5209 (N_5209,N_4307,N_4065);
or U5210 (N_5210,N_4445,N_4117);
or U5211 (N_5211,N_4168,N_4386);
nand U5212 (N_5212,N_4632,N_4704);
nor U5213 (N_5213,N_4509,N_4154);
xor U5214 (N_5214,N_4736,N_4427);
and U5215 (N_5215,N_4015,N_4523);
and U5216 (N_5216,N_4620,N_4077);
nor U5217 (N_5217,N_4363,N_4506);
xor U5218 (N_5218,N_4737,N_4574);
xnor U5219 (N_5219,N_4170,N_4740);
xnor U5220 (N_5220,N_4353,N_4785);
nand U5221 (N_5221,N_4078,N_4044);
nor U5222 (N_5222,N_4635,N_4333);
and U5223 (N_5223,N_4758,N_4321);
or U5224 (N_5224,N_4280,N_4448);
xnor U5225 (N_5225,N_4203,N_4147);
nand U5226 (N_5226,N_4567,N_4768);
xnor U5227 (N_5227,N_4086,N_4360);
nor U5228 (N_5228,N_4116,N_4610);
or U5229 (N_5229,N_4121,N_4538);
xnor U5230 (N_5230,N_4385,N_4026);
nand U5231 (N_5231,N_4716,N_4289);
or U5232 (N_5232,N_4736,N_4605);
nand U5233 (N_5233,N_4414,N_4486);
nand U5234 (N_5234,N_4287,N_4674);
and U5235 (N_5235,N_4600,N_4068);
and U5236 (N_5236,N_4638,N_4547);
nand U5237 (N_5237,N_4300,N_4171);
or U5238 (N_5238,N_4601,N_4133);
or U5239 (N_5239,N_4393,N_4479);
or U5240 (N_5240,N_4612,N_4269);
nor U5241 (N_5241,N_4348,N_4617);
and U5242 (N_5242,N_4197,N_4612);
xnor U5243 (N_5243,N_4790,N_4745);
xor U5244 (N_5244,N_4012,N_4655);
nand U5245 (N_5245,N_4473,N_4229);
xnor U5246 (N_5246,N_4208,N_4591);
or U5247 (N_5247,N_4620,N_4027);
or U5248 (N_5248,N_4309,N_4080);
nand U5249 (N_5249,N_4000,N_4681);
and U5250 (N_5250,N_4441,N_4569);
nor U5251 (N_5251,N_4706,N_4551);
and U5252 (N_5252,N_4700,N_4580);
nor U5253 (N_5253,N_4448,N_4309);
xor U5254 (N_5254,N_4288,N_4680);
nand U5255 (N_5255,N_4356,N_4445);
or U5256 (N_5256,N_4516,N_4177);
and U5257 (N_5257,N_4666,N_4519);
nor U5258 (N_5258,N_4294,N_4527);
nor U5259 (N_5259,N_4022,N_4251);
xor U5260 (N_5260,N_4408,N_4634);
xor U5261 (N_5261,N_4256,N_4737);
or U5262 (N_5262,N_4659,N_4448);
xnor U5263 (N_5263,N_4275,N_4721);
xor U5264 (N_5264,N_4387,N_4446);
or U5265 (N_5265,N_4161,N_4401);
xnor U5266 (N_5266,N_4298,N_4552);
nor U5267 (N_5267,N_4117,N_4579);
xor U5268 (N_5268,N_4339,N_4077);
nand U5269 (N_5269,N_4165,N_4414);
nor U5270 (N_5270,N_4283,N_4659);
or U5271 (N_5271,N_4757,N_4655);
xor U5272 (N_5272,N_4346,N_4287);
nor U5273 (N_5273,N_4381,N_4236);
xor U5274 (N_5274,N_4660,N_4612);
and U5275 (N_5275,N_4554,N_4689);
and U5276 (N_5276,N_4652,N_4163);
and U5277 (N_5277,N_4576,N_4162);
nand U5278 (N_5278,N_4149,N_4599);
xor U5279 (N_5279,N_4149,N_4499);
or U5280 (N_5280,N_4629,N_4055);
nor U5281 (N_5281,N_4004,N_4568);
nand U5282 (N_5282,N_4182,N_4052);
xnor U5283 (N_5283,N_4426,N_4624);
nor U5284 (N_5284,N_4288,N_4510);
xor U5285 (N_5285,N_4069,N_4421);
and U5286 (N_5286,N_4614,N_4134);
or U5287 (N_5287,N_4503,N_4474);
nand U5288 (N_5288,N_4271,N_4121);
xnor U5289 (N_5289,N_4145,N_4225);
nor U5290 (N_5290,N_4430,N_4405);
nand U5291 (N_5291,N_4703,N_4735);
or U5292 (N_5292,N_4755,N_4579);
and U5293 (N_5293,N_4380,N_4705);
nand U5294 (N_5294,N_4712,N_4438);
and U5295 (N_5295,N_4066,N_4643);
nand U5296 (N_5296,N_4094,N_4399);
nand U5297 (N_5297,N_4432,N_4466);
nand U5298 (N_5298,N_4207,N_4593);
nor U5299 (N_5299,N_4647,N_4181);
or U5300 (N_5300,N_4133,N_4680);
or U5301 (N_5301,N_4474,N_4338);
xnor U5302 (N_5302,N_4023,N_4722);
xnor U5303 (N_5303,N_4155,N_4195);
xor U5304 (N_5304,N_4550,N_4375);
and U5305 (N_5305,N_4015,N_4246);
nor U5306 (N_5306,N_4661,N_4344);
or U5307 (N_5307,N_4096,N_4131);
nand U5308 (N_5308,N_4627,N_4002);
nor U5309 (N_5309,N_4309,N_4546);
nand U5310 (N_5310,N_4212,N_4073);
and U5311 (N_5311,N_4629,N_4579);
xor U5312 (N_5312,N_4092,N_4045);
xnor U5313 (N_5313,N_4130,N_4302);
and U5314 (N_5314,N_4345,N_4369);
or U5315 (N_5315,N_4697,N_4076);
nor U5316 (N_5316,N_4310,N_4313);
and U5317 (N_5317,N_4433,N_4528);
nand U5318 (N_5318,N_4177,N_4473);
xnor U5319 (N_5319,N_4587,N_4289);
nand U5320 (N_5320,N_4266,N_4643);
xor U5321 (N_5321,N_4204,N_4155);
and U5322 (N_5322,N_4585,N_4277);
and U5323 (N_5323,N_4054,N_4575);
or U5324 (N_5324,N_4567,N_4719);
or U5325 (N_5325,N_4771,N_4351);
nand U5326 (N_5326,N_4023,N_4776);
or U5327 (N_5327,N_4262,N_4291);
xnor U5328 (N_5328,N_4031,N_4505);
xor U5329 (N_5329,N_4080,N_4563);
and U5330 (N_5330,N_4752,N_4370);
or U5331 (N_5331,N_4600,N_4646);
or U5332 (N_5332,N_4787,N_4709);
or U5333 (N_5333,N_4333,N_4345);
nand U5334 (N_5334,N_4727,N_4528);
nor U5335 (N_5335,N_4320,N_4149);
xor U5336 (N_5336,N_4697,N_4552);
nor U5337 (N_5337,N_4208,N_4079);
or U5338 (N_5338,N_4724,N_4546);
and U5339 (N_5339,N_4521,N_4202);
and U5340 (N_5340,N_4166,N_4086);
and U5341 (N_5341,N_4299,N_4406);
or U5342 (N_5342,N_4094,N_4498);
nand U5343 (N_5343,N_4042,N_4119);
xor U5344 (N_5344,N_4626,N_4218);
nor U5345 (N_5345,N_4173,N_4315);
and U5346 (N_5346,N_4777,N_4567);
nand U5347 (N_5347,N_4678,N_4436);
nand U5348 (N_5348,N_4799,N_4427);
and U5349 (N_5349,N_4125,N_4670);
xor U5350 (N_5350,N_4240,N_4695);
nand U5351 (N_5351,N_4235,N_4207);
and U5352 (N_5352,N_4685,N_4392);
xor U5353 (N_5353,N_4703,N_4282);
or U5354 (N_5354,N_4204,N_4705);
or U5355 (N_5355,N_4528,N_4182);
nor U5356 (N_5356,N_4605,N_4253);
xnor U5357 (N_5357,N_4283,N_4408);
nor U5358 (N_5358,N_4241,N_4299);
nor U5359 (N_5359,N_4160,N_4408);
nor U5360 (N_5360,N_4315,N_4133);
nand U5361 (N_5361,N_4021,N_4267);
xnor U5362 (N_5362,N_4383,N_4175);
xnor U5363 (N_5363,N_4635,N_4399);
xnor U5364 (N_5364,N_4611,N_4292);
nand U5365 (N_5365,N_4433,N_4319);
xnor U5366 (N_5366,N_4728,N_4179);
and U5367 (N_5367,N_4721,N_4309);
nor U5368 (N_5368,N_4495,N_4183);
nand U5369 (N_5369,N_4448,N_4469);
nand U5370 (N_5370,N_4606,N_4552);
and U5371 (N_5371,N_4402,N_4536);
nor U5372 (N_5372,N_4038,N_4736);
nand U5373 (N_5373,N_4798,N_4067);
xor U5374 (N_5374,N_4624,N_4046);
xor U5375 (N_5375,N_4017,N_4246);
xnor U5376 (N_5376,N_4284,N_4711);
nand U5377 (N_5377,N_4468,N_4150);
nor U5378 (N_5378,N_4454,N_4285);
or U5379 (N_5379,N_4767,N_4191);
nand U5380 (N_5380,N_4794,N_4155);
and U5381 (N_5381,N_4264,N_4169);
nor U5382 (N_5382,N_4082,N_4152);
xnor U5383 (N_5383,N_4537,N_4216);
and U5384 (N_5384,N_4476,N_4761);
or U5385 (N_5385,N_4553,N_4613);
nor U5386 (N_5386,N_4541,N_4752);
or U5387 (N_5387,N_4506,N_4478);
nand U5388 (N_5388,N_4400,N_4568);
nor U5389 (N_5389,N_4417,N_4419);
nor U5390 (N_5390,N_4158,N_4391);
nand U5391 (N_5391,N_4551,N_4676);
or U5392 (N_5392,N_4606,N_4061);
nor U5393 (N_5393,N_4657,N_4363);
and U5394 (N_5394,N_4396,N_4204);
and U5395 (N_5395,N_4587,N_4390);
or U5396 (N_5396,N_4103,N_4562);
and U5397 (N_5397,N_4656,N_4704);
xnor U5398 (N_5398,N_4169,N_4792);
xor U5399 (N_5399,N_4609,N_4182);
nor U5400 (N_5400,N_4770,N_4605);
xnor U5401 (N_5401,N_4782,N_4424);
or U5402 (N_5402,N_4178,N_4303);
nor U5403 (N_5403,N_4704,N_4174);
nor U5404 (N_5404,N_4757,N_4437);
nand U5405 (N_5405,N_4762,N_4132);
xor U5406 (N_5406,N_4571,N_4184);
and U5407 (N_5407,N_4371,N_4585);
nor U5408 (N_5408,N_4199,N_4057);
or U5409 (N_5409,N_4631,N_4537);
or U5410 (N_5410,N_4373,N_4464);
and U5411 (N_5411,N_4205,N_4693);
and U5412 (N_5412,N_4661,N_4338);
xor U5413 (N_5413,N_4771,N_4677);
xnor U5414 (N_5414,N_4484,N_4736);
and U5415 (N_5415,N_4126,N_4780);
and U5416 (N_5416,N_4772,N_4232);
and U5417 (N_5417,N_4264,N_4018);
or U5418 (N_5418,N_4521,N_4276);
xnor U5419 (N_5419,N_4043,N_4474);
nand U5420 (N_5420,N_4212,N_4505);
xnor U5421 (N_5421,N_4475,N_4154);
xnor U5422 (N_5422,N_4795,N_4339);
or U5423 (N_5423,N_4715,N_4017);
nand U5424 (N_5424,N_4737,N_4225);
and U5425 (N_5425,N_4467,N_4569);
or U5426 (N_5426,N_4239,N_4004);
or U5427 (N_5427,N_4325,N_4626);
or U5428 (N_5428,N_4686,N_4047);
nand U5429 (N_5429,N_4117,N_4539);
nand U5430 (N_5430,N_4179,N_4688);
and U5431 (N_5431,N_4646,N_4675);
xnor U5432 (N_5432,N_4341,N_4503);
xor U5433 (N_5433,N_4459,N_4466);
xnor U5434 (N_5434,N_4070,N_4115);
or U5435 (N_5435,N_4394,N_4570);
and U5436 (N_5436,N_4306,N_4546);
nor U5437 (N_5437,N_4466,N_4332);
or U5438 (N_5438,N_4471,N_4378);
nor U5439 (N_5439,N_4749,N_4356);
or U5440 (N_5440,N_4753,N_4226);
and U5441 (N_5441,N_4552,N_4308);
nor U5442 (N_5442,N_4240,N_4126);
or U5443 (N_5443,N_4142,N_4545);
or U5444 (N_5444,N_4744,N_4796);
and U5445 (N_5445,N_4574,N_4681);
or U5446 (N_5446,N_4637,N_4665);
xor U5447 (N_5447,N_4632,N_4506);
or U5448 (N_5448,N_4087,N_4259);
or U5449 (N_5449,N_4747,N_4350);
xor U5450 (N_5450,N_4200,N_4214);
nand U5451 (N_5451,N_4664,N_4344);
and U5452 (N_5452,N_4194,N_4168);
xor U5453 (N_5453,N_4258,N_4707);
nor U5454 (N_5454,N_4155,N_4650);
and U5455 (N_5455,N_4096,N_4670);
nand U5456 (N_5456,N_4483,N_4766);
and U5457 (N_5457,N_4009,N_4530);
nor U5458 (N_5458,N_4635,N_4726);
nand U5459 (N_5459,N_4253,N_4036);
or U5460 (N_5460,N_4246,N_4324);
and U5461 (N_5461,N_4724,N_4421);
or U5462 (N_5462,N_4791,N_4010);
and U5463 (N_5463,N_4533,N_4107);
xor U5464 (N_5464,N_4394,N_4630);
and U5465 (N_5465,N_4632,N_4695);
or U5466 (N_5466,N_4285,N_4666);
nand U5467 (N_5467,N_4362,N_4551);
or U5468 (N_5468,N_4583,N_4154);
and U5469 (N_5469,N_4696,N_4622);
xor U5470 (N_5470,N_4268,N_4382);
xor U5471 (N_5471,N_4756,N_4656);
and U5472 (N_5472,N_4247,N_4372);
nand U5473 (N_5473,N_4360,N_4519);
and U5474 (N_5474,N_4046,N_4019);
or U5475 (N_5475,N_4248,N_4065);
nor U5476 (N_5476,N_4367,N_4272);
xor U5477 (N_5477,N_4586,N_4519);
nand U5478 (N_5478,N_4769,N_4583);
and U5479 (N_5479,N_4410,N_4720);
xnor U5480 (N_5480,N_4107,N_4237);
or U5481 (N_5481,N_4260,N_4455);
xor U5482 (N_5482,N_4559,N_4501);
and U5483 (N_5483,N_4035,N_4584);
or U5484 (N_5484,N_4507,N_4298);
nor U5485 (N_5485,N_4694,N_4392);
xor U5486 (N_5486,N_4421,N_4521);
xor U5487 (N_5487,N_4346,N_4061);
and U5488 (N_5488,N_4707,N_4565);
nand U5489 (N_5489,N_4283,N_4512);
nor U5490 (N_5490,N_4644,N_4343);
xor U5491 (N_5491,N_4025,N_4790);
nand U5492 (N_5492,N_4699,N_4140);
nor U5493 (N_5493,N_4780,N_4233);
xor U5494 (N_5494,N_4199,N_4148);
nand U5495 (N_5495,N_4012,N_4600);
nand U5496 (N_5496,N_4097,N_4064);
xor U5497 (N_5497,N_4369,N_4393);
xnor U5498 (N_5498,N_4420,N_4194);
xnor U5499 (N_5499,N_4161,N_4542);
nor U5500 (N_5500,N_4445,N_4653);
xor U5501 (N_5501,N_4793,N_4695);
nand U5502 (N_5502,N_4621,N_4495);
or U5503 (N_5503,N_4561,N_4026);
nand U5504 (N_5504,N_4279,N_4289);
nand U5505 (N_5505,N_4676,N_4553);
xnor U5506 (N_5506,N_4655,N_4013);
xor U5507 (N_5507,N_4080,N_4490);
or U5508 (N_5508,N_4021,N_4147);
or U5509 (N_5509,N_4533,N_4035);
or U5510 (N_5510,N_4579,N_4672);
or U5511 (N_5511,N_4411,N_4456);
or U5512 (N_5512,N_4219,N_4131);
and U5513 (N_5513,N_4617,N_4405);
xor U5514 (N_5514,N_4170,N_4191);
nand U5515 (N_5515,N_4251,N_4721);
nand U5516 (N_5516,N_4034,N_4699);
nand U5517 (N_5517,N_4684,N_4544);
nand U5518 (N_5518,N_4475,N_4733);
or U5519 (N_5519,N_4056,N_4582);
xor U5520 (N_5520,N_4062,N_4250);
or U5521 (N_5521,N_4660,N_4005);
and U5522 (N_5522,N_4311,N_4456);
or U5523 (N_5523,N_4140,N_4650);
xor U5524 (N_5524,N_4584,N_4728);
nor U5525 (N_5525,N_4035,N_4269);
and U5526 (N_5526,N_4759,N_4773);
nor U5527 (N_5527,N_4366,N_4418);
and U5528 (N_5528,N_4423,N_4230);
nand U5529 (N_5529,N_4032,N_4472);
or U5530 (N_5530,N_4073,N_4196);
nor U5531 (N_5531,N_4799,N_4473);
nor U5532 (N_5532,N_4367,N_4193);
or U5533 (N_5533,N_4536,N_4345);
and U5534 (N_5534,N_4101,N_4144);
nand U5535 (N_5535,N_4177,N_4359);
or U5536 (N_5536,N_4485,N_4041);
xnor U5537 (N_5537,N_4496,N_4549);
or U5538 (N_5538,N_4786,N_4448);
and U5539 (N_5539,N_4509,N_4512);
xor U5540 (N_5540,N_4137,N_4625);
xnor U5541 (N_5541,N_4408,N_4137);
or U5542 (N_5542,N_4098,N_4369);
or U5543 (N_5543,N_4103,N_4586);
nand U5544 (N_5544,N_4232,N_4392);
or U5545 (N_5545,N_4271,N_4745);
xor U5546 (N_5546,N_4616,N_4648);
xor U5547 (N_5547,N_4517,N_4159);
and U5548 (N_5548,N_4155,N_4331);
nand U5549 (N_5549,N_4764,N_4028);
xor U5550 (N_5550,N_4723,N_4447);
nand U5551 (N_5551,N_4665,N_4243);
nand U5552 (N_5552,N_4258,N_4324);
or U5553 (N_5553,N_4352,N_4764);
nor U5554 (N_5554,N_4444,N_4193);
nor U5555 (N_5555,N_4312,N_4064);
and U5556 (N_5556,N_4775,N_4604);
xnor U5557 (N_5557,N_4311,N_4531);
nor U5558 (N_5558,N_4403,N_4603);
nand U5559 (N_5559,N_4219,N_4682);
or U5560 (N_5560,N_4041,N_4547);
or U5561 (N_5561,N_4695,N_4188);
nor U5562 (N_5562,N_4415,N_4569);
xnor U5563 (N_5563,N_4364,N_4502);
xor U5564 (N_5564,N_4192,N_4029);
nor U5565 (N_5565,N_4139,N_4733);
nor U5566 (N_5566,N_4520,N_4606);
nor U5567 (N_5567,N_4093,N_4495);
xor U5568 (N_5568,N_4357,N_4713);
nor U5569 (N_5569,N_4559,N_4633);
nand U5570 (N_5570,N_4428,N_4232);
or U5571 (N_5571,N_4399,N_4781);
xnor U5572 (N_5572,N_4781,N_4149);
or U5573 (N_5573,N_4164,N_4174);
or U5574 (N_5574,N_4530,N_4798);
or U5575 (N_5575,N_4076,N_4100);
and U5576 (N_5576,N_4785,N_4307);
and U5577 (N_5577,N_4385,N_4720);
nand U5578 (N_5578,N_4419,N_4281);
xor U5579 (N_5579,N_4497,N_4505);
nand U5580 (N_5580,N_4545,N_4727);
nand U5581 (N_5581,N_4044,N_4143);
and U5582 (N_5582,N_4270,N_4595);
nor U5583 (N_5583,N_4599,N_4647);
or U5584 (N_5584,N_4282,N_4403);
nor U5585 (N_5585,N_4010,N_4672);
or U5586 (N_5586,N_4679,N_4348);
or U5587 (N_5587,N_4680,N_4703);
nor U5588 (N_5588,N_4328,N_4542);
nand U5589 (N_5589,N_4577,N_4180);
and U5590 (N_5590,N_4125,N_4612);
and U5591 (N_5591,N_4089,N_4231);
and U5592 (N_5592,N_4539,N_4058);
and U5593 (N_5593,N_4417,N_4527);
xnor U5594 (N_5594,N_4220,N_4463);
or U5595 (N_5595,N_4121,N_4359);
nand U5596 (N_5596,N_4773,N_4449);
and U5597 (N_5597,N_4102,N_4158);
and U5598 (N_5598,N_4478,N_4388);
or U5599 (N_5599,N_4549,N_4322);
or U5600 (N_5600,N_4870,N_5561);
nand U5601 (N_5601,N_5428,N_4891);
xnor U5602 (N_5602,N_4855,N_5360);
nor U5603 (N_5603,N_4850,N_5212);
nor U5604 (N_5604,N_5300,N_5149);
xnor U5605 (N_5605,N_5227,N_5399);
nand U5606 (N_5606,N_5412,N_5543);
or U5607 (N_5607,N_5186,N_5295);
and U5608 (N_5608,N_4848,N_5043);
nand U5609 (N_5609,N_5336,N_5488);
nor U5610 (N_5610,N_5196,N_5278);
xor U5611 (N_5611,N_5550,N_4814);
xnor U5612 (N_5612,N_5093,N_5234);
nor U5613 (N_5613,N_5144,N_4902);
nand U5614 (N_5614,N_4963,N_5071);
and U5615 (N_5615,N_5297,N_4898);
nor U5616 (N_5616,N_5502,N_4880);
nand U5617 (N_5617,N_5587,N_5537);
and U5618 (N_5618,N_4923,N_4985);
or U5619 (N_5619,N_5563,N_5010);
nor U5620 (N_5620,N_5568,N_5358);
nor U5621 (N_5621,N_5530,N_5244);
nand U5622 (N_5622,N_5275,N_5433);
and U5623 (N_5623,N_4852,N_5231);
xnor U5624 (N_5624,N_5283,N_5210);
nor U5625 (N_5625,N_5396,N_5238);
nand U5626 (N_5626,N_5299,N_5486);
or U5627 (N_5627,N_4926,N_5450);
nor U5628 (N_5628,N_5110,N_4817);
nand U5629 (N_5629,N_4900,N_5407);
nand U5630 (N_5630,N_5138,N_5484);
xor U5631 (N_5631,N_5007,N_5024);
nor U5632 (N_5632,N_5245,N_5103);
nor U5633 (N_5633,N_5585,N_4876);
nor U5634 (N_5634,N_5558,N_4966);
nand U5635 (N_5635,N_5174,N_5386);
xor U5636 (N_5636,N_5239,N_5286);
and U5637 (N_5637,N_4980,N_5124);
xor U5638 (N_5638,N_4962,N_5025);
nor U5639 (N_5639,N_5437,N_5122);
or U5640 (N_5640,N_4942,N_5288);
nand U5641 (N_5641,N_5084,N_5081);
nor U5642 (N_5642,N_5107,N_5158);
xor U5643 (N_5643,N_5083,N_5355);
or U5644 (N_5644,N_5116,N_5304);
or U5645 (N_5645,N_5390,N_4928);
xnor U5646 (N_5646,N_4911,N_5415);
nor U5647 (N_5647,N_4912,N_5513);
and U5648 (N_5648,N_5435,N_5385);
xor U5649 (N_5649,N_4973,N_5205);
or U5650 (N_5650,N_4836,N_5020);
nand U5651 (N_5651,N_5152,N_5564);
nor U5652 (N_5652,N_5487,N_5254);
nand U5653 (N_5653,N_5303,N_4976);
nor U5654 (N_5654,N_5281,N_5137);
nor U5655 (N_5655,N_5596,N_5185);
nor U5656 (N_5656,N_4968,N_5426);
and U5657 (N_5657,N_5177,N_5459);
xor U5658 (N_5658,N_5542,N_5371);
xnor U5659 (N_5659,N_5246,N_5593);
xor U5660 (N_5660,N_5482,N_4935);
nor U5661 (N_5661,N_4945,N_5023);
nand U5662 (N_5662,N_5269,N_5001);
or U5663 (N_5663,N_5148,N_5074);
or U5664 (N_5664,N_5580,N_4934);
nand U5665 (N_5665,N_5452,N_5471);
xnor U5666 (N_5666,N_5445,N_5141);
nor U5667 (N_5667,N_5125,N_5349);
xor U5668 (N_5668,N_5361,N_5500);
xnor U5669 (N_5669,N_5576,N_4864);
nor U5670 (N_5670,N_5479,N_5508);
nor U5671 (N_5671,N_4938,N_5095);
xor U5672 (N_5672,N_4987,N_4967);
nor U5673 (N_5673,N_4932,N_5492);
and U5674 (N_5674,N_5540,N_4809);
nor U5675 (N_5675,N_5345,N_5485);
xnor U5676 (N_5676,N_4916,N_5251);
nand U5677 (N_5677,N_5014,N_5217);
xor U5678 (N_5678,N_5541,N_5153);
xor U5679 (N_5679,N_4933,N_5397);
nand U5680 (N_5680,N_5041,N_5092);
nor U5681 (N_5681,N_4847,N_5357);
nor U5682 (N_5682,N_5599,N_4894);
nor U5683 (N_5683,N_5421,N_5378);
xor U5684 (N_5684,N_5526,N_5105);
nor U5685 (N_5685,N_5581,N_5455);
xnor U5686 (N_5686,N_5190,N_5442);
nor U5687 (N_5687,N_5392,N_5277);
nand U5688 (N_5688,N_5062,N_5061);
nand U5689 (N_5689,N_5424,N_5533);
xor U5690 (N_5690,N_5047,N_4803);
and U5691 (N_5691,N_5070,N_5341);
xnor U5692 (N_5692,N_5404,N_5598);
or U5693 (N_5693,N_5100,N_5156);
and U5694 (N_5694,N_5069,N_5194);
nor U5695 (N_5695,N_5272,N_5091);
and U5696 (N_5696,N_4965,N_5334);
nand U5697 (N_5697,N_4979,N_5298);
xor U5698 (N_5698,N_5539,N_4883);
xor U5699 (N_5699,N_5060,N_5466);
and U5700 (N_5700,N_5005,N_5344);
or U5701 (N_5701,N_5225,N_5570);
nand U5702 (N_5702,N_5119,N_5055);
xnor U5703 (N_5703,N_5520,N_5409);
and U5704 (N_5704,N_5208,N_4820);
nand U5705 (N_5705,N_4990,N_5490);
and U5706 (N_5706,N_5551,N_5094);
or U5707 (N_5707,N_5028,N_5525);
xor U5708 (N_5708,N_5139,N_5270);
or U5709 (N_5709,N_5160,N_4800);
or U5710 (N_5710,N_4819,N_5247);
xor U5711 (N_5711,N_5253,N_5521);
nor U5712 (N_5712,N_4995,N_4869);
nor U5713 (N_5713,N_4878,N_4867);
and U5714 (N_5714,N_5219,N_5590);
xor U5715 (N_5715,N_5380,N_5516);
or U5716 (N_5716,N_5274,N_5154);
or U5717 (N_5717,N_5207,N_4879);
or U5718 (N_5718,N_5181,N_5519);
and U5719 (N_5719,N_5040,N_5259);
nand U5720 (N_5720,N_5309,N_5438);
xnor U5721 (N_5721,N_4948,N_5058);
nand U5722 (N_5722,N_5117,N_5209);
or U5723 (N_5723,N_4984,N_5066);
or U5724 (N_5724,N_5322,N_5106);
nor U5725 (N_5725,N_5584,N_5577);
nor U5726 (N_5726,N_5464,N_5574);
nor U5727 (N_5727,N_5008,N_5536);
and U5728 (N_5728,N_5036,N_5302);
nor U5729 (N_5729,N_5211,N_5104);
or U5730 (N_5730,N_5328,N_5401);
nand U5731 (N_5731,N_5501,N_5050);
and U5732 (N_5732,N_4840,N_4931);
and U5733 (N_5733,N_5446,N_5178);
or U5734 (N_5734,N_5556,N_5032);
xnor U5735 (N_5735,N_5402,N_4947);
xnor U5736 (N_5736,N_4949,N_5215);
xor U5737 (N_5737,N_5367,N_5579);
and U5738 (N_5738,N_5268,N_4802);
xnor U5739 (N_5739,N_5495,N_5534);
or U5740 (N_5740,N_5132,N_5049);
and U5741 (N_5741,N_5381,N_4854);
nor U5742 (N_5742,N_4944,N_5097);
nor U5743 (N_5743,N_5226,N_5423);
nand U5744 (N_5744,N_4868,N_5547);
nor U5745 (N_5745,N_5056,N_5059);
and U5746 (N_5746,N_5594,N_5221);
and U5747 (N_5747,N_4858,N_5368);
and U5748 (N_5748,N_5434,N_4826);
nor U5749 (N_5749,N_5481,N_4881);
nor U5750 (N_5750,N_5443,N_5123);
nand U5751 (N_5751,N_4953,N_5170);
or U5752 (N_5752,N_4837,N_4896);
and U5753 (N_5753,N_5553,N_5376);
nor U5754 (N_5754,N_5507,N_5366);
or U5755 (N_5755,N_4815,N_4919);
and U5756 (N_5756,N_5037,N_5391);
and U5757 (N_5757,N_5477,N_5108);
nor U5758 (N_5758,N_4908,N_5162);
or U5759 (N_5759,N_5009,N_5469);
xor U5760 (N_5760,N_5048,N_4839);
xor U5761 (N_5761,N_5191,N_4853);
xor U5762 (N_5762,N_5291,N_5276);
xnor U5763 (N_5763,N_5389,N_5133);
or U5764 (N_5764,N_5483,N_4961);
xor U5765 (N_5765,N_5565,N_5359);
nand U5766 (N_5766,N_5496,N_5235);
or U5767 (N_5767,N_5175,N_5535);
nor U5768 (N_5768,N_5311,N_4970);
or U5769 (N_5769,N_5354,N_5240);
nand U5770 (N_5770,N_5575,N_5347);
or U5771 (N_5771,N_5130,N_5339);
nand U5772 (N_5772,N_4807,N_5578);
or U5773 (N_5773,N_4917,N_5128);
and U5774 (N_5774,N_4921,N_5489);
nor U5775 (N_5775,N_5063,N_5476);
and U5776 (N_5776,N_5363,N_5332);
xnor U5777 (N_5777,N_4981,N_5429);
nor U5778 (N_5778,N_5290,N_5072);
nand U5779 (N_5779,N_5427,N_4895);
or U5780 (N_5780,N_5155,N_4986);
nand U5781 (N_5781,N_5287,N_5078);
nand U5782 (N_5782,N_5314,N_5377);
xnor U5783 (N_5783,N_5499,N_5224);
nor U5784 (N_5784,N_4846,N_5187);
xnor U5785 (N_5785,N_4808,N_5467);
xnor U5786 (N_5786,N_5046,N_5086);
nand U5787 (N_5787,N_5447,N_4831);
and U5788 (N_5788,N_5528,N_5098);
xor U5789 (N_5789,N_5035,N_4842);
xnor U5790 (N_5790,N_4920,N_5414);
and U5791 (N_5791,N_4982,N_4838);
nand U5792 (N_5792,N_4857,N_5329);
or U5793 (N_5793,N_5305,N_4994);
nor U5794 (N_5794,N_5171,N_5375);
and U5795 (N_5795,N_5370,N_5146);
and U5796 (N_5796,N_4887,N_5263);
and U5797 (N_5797,N_5232,N_5260);
and U5798 (N_5798,N_4884,N_4950);
nand U5799 (N_5799,N_5372,N_5431);
or U5800 (N_5800,N_5456,N_4951);
nand U5801 (N_5801,N_5549,N_5324);
nand U5802 (N_5802,N_4977,N_5505);
and U5803 (N_5803,N_5085,N_4863);
and U5804 (N_5804,N_5134,N_5356);
nor U5805 (N_5805,N_5261,N_5282);
or U5806 (N_5806,N_5463,N_5013);
and U5807 (N_5807,N_5465,N_4877);
nor U5808 (N_5808,N_5201,N_5015);
nor U5809 (N_5809,N_5557,N_5420);
xor U5810 (N_5810,N_5088,N_4806);
nand U5811 (N_5811,N_5182,N_5292);
nand U5812 (N_5812,N_5257,N_5019);
and U5813 (N_5813,N_5111,N_5338);
xor U5814 (N_5814,N_5068,N_5545);
and U5815 (N_5815,N_5364,N_5184);
nand U5816 (N_5816,N_5457,N_5462);
or U5817 (N_5817,N_5112,N_5441);
nand U5818 (N_5818,N_5242,N_5192);
nand U5819 (N_5819,N_4983,N_5284);
nand U5820 (N_5820,N_5589,N_5218);
nand U5821 (N_5821,N_5315,N_5419);
xor U5822 (N_5822,N_4882,N_4909);
nor U5823 (N_5823,N_5096,N_5374);
or U5824 (N_5824,N_5422,N_5440);
or U5825 (N_5825,N_5538,N_4943);
or U5826 (N_5826,N_5183,N_5518);
or U5827 (N_5827,N_5475,N_5460);
and U5828 (N_5828,N_5002,N_5510);
xor U5829 (N_5829,N_5101,N_4969);
nand U5830 (N_5830,N_5472,N_5038);
xor U5831 (N_5831,N_5480,N_5405);
or U5832 (N_5832,N_5161,N_5410);
or U5833 (N_5833,N_4805,N_4940);
and U5834 (N_5834,N_5418,N_4924);
nor U5835 (N_5835,N_4975,N_5362);
nor U5836 (N_5836,N_4885,N_4890);
and U5837 (N_5837,N_5403,N_5451);
and U5838 (N_5838,N_5393,N_5301);
nand U5839 (N_5839,N_5319,N_5473);
or U5840 (N_5840,N_5195,N_5400);
nand U5841 (N_5841,N_5265,N_5204);
and U5842 (N_5842,N_5216,N_4810);
xor U5843 (N_5843,N_5065,N_5279);
nand U5844 (N_5844,N_5200,N_5494);
nor U5845 (N_5845,N_5250,N_5523);
nor U5846 (N_5846,N_4874,N_4816);
nor U5847 (N_5847,N_5323,N_4835);
nor U5848 (N_5848,N_5252,N_4866);
nor U5849 (N_5849,N_4833,N_5229);
and U5850 (N_5850,N_4957,N_4865);
nor U5851 (N_5851,N_4978,N_4832);
xor U5852 (N_5852,N_5021,N_4939);
nand U5853 (N_5853,N_5089,N_5512);
xnor U5854 (N_5854,N_4906,N_4910);
xnor U5855 (N_5855,N_4812,N_5214);
or U5856 (N_5856,N_5143,N_5317);
or U5857 (N_5857,N_5033,N_5006);
nor U5858 (N_5858,N_5591,N_5454);
and U5859 (N_5859,N_5118,N_5076);
and U5860 (N_5860,N_5326,N_5053);
or U5861 (N_5861,N_4851,N_5230);
nor U5862 (N_5862,N_5388,N_5560);
and U5863 (N_5863,N_5387,N_5016);
xnor U5864 (N_5864,N_4897,N_5318);
nor U5865 (N_5865,N_5213,N_5249);
or U5866 (N_5866,N_5258,N_4998);
nor U5867 (N_5867,N_5237,N_5307);
xor U5868 (N_5868,N_5327,N_5515);
xnor U5869 (N_5869,N_4960,N_4915);
nor U5870 (N_5870,N_5202,N_5168);
nor U5871 (N_5871,N_5030,N_5289);
xnor U5872 (N_5872,N_5064,N_5504);
and U5873 (N_5873,N_5176,N_5271);
or U5874 (N_5874,N_5478,N_5312);
nand U5875 (N_5875,N_4822,N_5382);
nand U5876 (N_5876,N_4834,N_4830);
nand U5877 (N_5877,N_5498,N_5497);
nor U5878 (N_5878,N_5082,N_4997);
nand U5879 (N_5879,N_5529,N_4958);
or U5880 (N_5880,N_5057,N_5203);
and U5881 (N_5881,N_5206,N_5582);
nor U5882 (N_5882,N_4843,N_5012);
and U5883 (N_5883,N_4813,N_5562);
and U5884 (N_5884,N_5109,N_4849);
xor U5885 (N_5885,N_4823,N_4922);
or U5886 (N_5886,N_5436,N_5145);
xnor U5887 (N_5887,N_4929,N_5115);
xnor U5888 (N_5888,N_4964,N_5506);
or U5889 (N_5889,N_5342,N_4956);
xor U5890 (N_5890,N_5416,N_5430);
nor U5891 (N_5891,N_5102,N_5126);
and U5892 (N_5892,N_5042,N_5353);
xor U5893 (N_5893,N_5017,N_5503);
nor U5894 (N_5894,N_4914,N_4925);
xnor U5895 (N_5895,N_4801,N_5461);
and U5896 (N_5896,N_4872,N_5554);
nor U5897 (N_5897,N_5198,N_4892);
and U5898 (N_5898,N_5567,N_5524);
and U5899 (N_5899,N_5532,N_5011);
nand U5900 (N_5900,N_5129,N_5316);
nand U5901 (N_5901,N_5348,N_5384);
or U5902 (N_5902,N_5188,N_5280);
and U5903 (N_5903,N_5294,N_5310);
nand U5904 (N_5904,N_4989,N_4862);
and U5905 (N_5905,N_5169,N_5571);
and U5906 (N_5906,N_5468,N_5255);
and U5907 (N_5907,N_5142,N_5439);
and U5908 (N_5908,N_4993,N_5340);
nor U5909 (N_5909,N_5337,N_4907);
or U5910 (N_5910,N_5267,N_5173);
nand U5911 (N_5911,N_4893,N_5449);
nand U5912 (N_5912,N_5151,N_4991);
xnor U5913 (N_5913,N_5022,N_5079);
nand U5914 (N_5914,N_5548,N_5511);
or U5915 (N_5915,N_5003,N_5165);
nand U5916 (N_5916,N_5136,N_4845);
nand U5917 (N_5917,N_5406,N_5131);
xnor U5918 (N_5918,N_4959,N_5425);
or U5919 (N_5919,N_4818,N_5527);
nand U5920 (N_5920,N_5027,N_5262);
nand U5921 (N_5921,N_4829,N_5164);
xor U5922 (N_5922,N_5569,N_5113);
nand U5923 (N_5923,N_4860,N_5222);
xnor U5924 (N_5924,N_4904,N_5383);
or U5925 (N_5925,N_5592,N_5099);
or U5926 (N_5926,N_5248,N_5373);
xnor U5927 (N_5927,N_5597,N_4905);
xnor U5928 (N_5928,N_5331,N_5051);
and U5929 (N_5929,N_5150,N_5335);
nand U5930 (N_5930,N_5163,N_5127);
xnor U5931 (N_5931,N_5179,N_5266);
nand U5932 (N_5932,N_4901,N_4844);
nor U5933 (N_5933,N_5167,N_5413);
and U5934 (N_5934,N_5306,N_4988);
xnor U5935 (N_5935,N_5273,N_5052);
or U5936 (N_5936,N_5509,N_5199);
and U5937 (N_5937,N_5432,N_5285);
xnor U5938 (N_5938,N_4871,N_5352);
xnor U5939 (N_5939,N_4889,N_5080);
xor U5940 (N_5940,N_5448,N_5120);
nor U5941 (N_5941,N_5411,N_5350);
nand U5942 (N_5942,N_4971,N_5087);
and U5943 (N_5943,N_5140,N_5379);
nor U5944 (N_5944,N_5333,N_4899);
or U5945 (N_5945,N_4936,N_5147);
nand U5946 (N_5946,N_4828,N_5514);
xor U5947 (N_5947,N_5073,N_4903);
xnor U5948 (N_5948,N_4821,N_5583);
and U5949 (N_5949,N_4937,N_4972);
nor U5950 (N_5950,N_5453,N_4804);
nand U5951 (N_5951,N_5233,N_5296);
or U5952 (N_5952,N_4996,N_5351);
xor U5953 (N_5953,N_5365,N_5517);
xnor U5954 (N_5954,N_5018,N_5159);
or U5955 (N_5955,N_5075,N_5308);
and U5956 (N_5956,N_5031,N_5243);
and U5957 (N_5957,N_5444,N_5077);
nor U5958 (N_5958,N_5236,N_5408);
nor U5959 (N_5959,N_5458,N_5474);
or U5960 (N_5960,N_5531,N_5552);
nand U5961 (N_5961,N_4888,N_5135);
xor U5962 (N_5962,N_5264,N_5029);
nor U5963 (N_5963,N_5000,N_4930);
xnor U5964 (N_5964,N_5172,N_5321);
nand U5965 (N_5965,N_5325,N_5346);
and U5966 (N_5966,N_5223,N_5573);
xor U5967 (N_5967,N_5220,N_4954);
nor U5968 (N_5968,N_5595,N_4825);
nand U5969 (N_5969,N_5586,N_5559);
and U5970 (N_5970,N_5026,N_4941);
and U5971 (N_5971,N_5369,N_5189);
and U5972 (N_5972,N_4856,N_5034);
xor U5973 (N_5973,N_5157,N_5588);
nor U5974 (N_5974,N_4992,N_4875);
or U5975 (N_5975,N_4811,N_5544);
xor U5976 (N_5976,N_5343,N_5555);
xor U5977 (N_5977,N_5394,N_5039);
xor U5978 (N_5978,N_5330,N_5044);
and U5979 (N_5979,N_5491,N_5193);
and U5980 (N_5980,N_5241,N_4824);
xnor U5981 (N_5981,N_5546,N_4955);
or U5982 (N_5982,N_5045,N_5121);
xor U5983 (N_5983,N_4946,N_5417);
nand U5984 (N_5984,N_5493,N_5313);
nand U5985 (N_5985,N_5522,N_4861);
and U5986 (N_5986,N_5293,N_4952);
or U5987 (N_5987,N_5090,N_4999);
xor U5988 (N_5988,N_5398,N_5067);
and U5989 (N_5989,N_4859,N_5054);
nand U5990 (N_5990,N_4918,N_5256);
nand U5991 (N_5991,N_4841,N_5470);
nor U5992 (N_5992,N_5395,N_5197);
nand U5993 (N_5993,N_5114,N_4913);
nor U5994 (N_5994,N_4974,N_5566);
nand U5995 (N_5995,N_4827,N_5320);
or U5996 (N_5996,N_5180,N_5572);
and U5997 (N_5997,N_5166,N_5004);
nor U5998 (N_5998,N_5228,N_4927);
nand U5999 (N_5999,N_4873,N_4886);
nor U6000 (N_6000,N_5240,N_5556);
or U6001 (N_6001,N_5087,N_5080);
and U6002 (N_6002,N_5421,N_5592);
or U6003 (N_6003,N_4909,N_4968);
and U6004 (N_6004,N_5092,N_5251);
nand U6005 (N_6005,N_5199,N_5297);
nand U6006 (N_6006,N_5216,N_5263);
xor U6007 (N_6007,N_4951,N_5542);
xor U6008 (N_6008,N_5052,N_4894);
xor U6009 (N_6009,N_5083,N_4990);
or U6010 (N_6010,N_5515,N_5463);
or U6011 (N_6011,N_5191,N_5034);
or U6012 (N_6012,N_5026,N_5059);
or U6013 (N_6013,N_5560,N_5541);
xor U6014 (N_6014,N_5071,N_5093);
xnor U6015 (N_6015,N_5493,N_5010);
and U6016 (N_6016,N_5584,N_5448);
and U6017 (N_6017,N_5401,N_5165);
and U6018 (N_6018,N_5571,N_5186);
or U6019 (N_6019,N_5114,N_4866);
nand U6020 (N_6020,N_5414,N_5499);
or U6021 (N_6021,N_5539,N_4806);
nor U6022 (N_6022,N_5226,N_5048);
nor U6023 (N_6023,N_5053,N_4894);
or U6024 (N_6024,N_5351,N_5269);
xnor U6025 (N_6025,N_4992,N_4949);
and U6026 (N_6026,N_5342,N_5516);
nor U6027 (N_6027,N_4866,N_5294);
and U6028 (N_6028,N_4915,N_5522);
xnor U6029 (N_6029,N_5086,N_5127);
nor U6030 (N_6030,N_4970,N_4842);
xnor U6031 (N_6031,N_4865,N_4849);
nor U6032 (N_6032,N_5237,N_5109);
and U6033 (N_6033,N_5064,N_4954);
or U6034 (N_6034,N_4964,N_5313);
and U6035 (N_6035,N_4873,N_5197);
and U6036 (N_6036,N_4986,N_5298);
nand U6037 (N_6037,N_5362,N_5339);
and U6038 (N_6038,N_4816,N_5129);
nand U6039 (N_6039,N_5018,N_4895);
xnor U6040 (N_6040,N_5596,N_5059);
nor U6041 (N_6041,N_5476,N_5554);
xor U6042 (N_6042,N_4806,N_5377);
nor U6043 (N_6043,N_5075,N_5379);
xnor U6044 (N_6044,N_5571,N_5046);
and U6045 (N_6045,N_5004,N_5085);
nand U6046 (N_6046,N_4848,N_4861);
nor U6047 (N_6047,N_5494,N_5194);
nor U6048 (N_6048,N_4846,N_4955);
nor U6049 (N_6049,N_5501,N_5567);
or U6050 (N_6050,N_5409,N_5472);
and U6051 (N_6051,N_5312,N_5119);
or U6052 (N_6052,N_4861,N_5135);
nand U6053 (N_6053,N_4818,N_5104);
nand U6054 (N_6054,N_5098,N_5588);
and U6055 (N_6055,N_5574,N_5485);
nand U6056 (N_6056,N_4910,N_5309);
nand U6057 (N_6057,N_5056,N_5341);
or U6058 (N_6058,N_4940,N_5194);
and U6059 (N_6059,N_5112,N_5323);
nor U6060 (N_6060,N_5025,N_4822);
and U6061 (N_6061,N_5181,N_5539);
or U6062 (N_6062,N_4876,N_5479);
and U6063 (N_6063,N_4857,N_4846);
nand U6064 (N_6064,N_5256,N_5559);
nor U6065 (N_6065,N_4802,N_5014);
or U6066 (N_6066,N_5417,N_5584);
nor U6067 (N_6067,N_4930,N_5280);
and U6068 (N_6068,N_5271,N_5268);
nor U6069 (N_6069,N_5390,N_5017);
or U6070 (N_6070,N_4859,N_5309);
xnor U6071 (N_6071,N_5351,N_5406);
nand U6072 (N_6072,N_4880,N_5046);
or U6073 (N_6073,N_5121,N_5134);
and U6074 (N_6074,N_4991,N_5177);
nor U6075 (N_6075,N_5135,N_4900);
nor U6076 (N_6076,N_5197,N_5278);
nand U6077 (N_6077,N_5413,N_5201);
and U6078 (N_6078,N_5520,N_4951);
or U6079 (N_6079,N_5534,N_5585);
and U6080 (N_6080,N_5480,N_5237);
nand U6081 (N_6081,N_5371,N_5473);
xor U6082 (N_6082,N_5514,N_4823);
or U6083 (N_6083,N_5393,N_5097);
nand U6084 (N_6084,N_4976,N_5266);
or U6085 (N_6085,N_5077,N_5063);
and U6086 (N_6086,N_4866,N_5317);
and U6087 (N_6087,N_5306,N_5170);
xor U6088 (N_6088,N_4906,N_5250);
nor U6089 (N_6089,N_4810,N_5403);
and U6090 (N_6090,N_5459,N_5198);
nand U6091 (N_6091,N_5079,N_5020);
nor U6092 (N_6092,N_5126,N_5002);
or U6093 (N_6093,N_5468,N_5055);
nor U6094 (N_6094,N_5229,N_5293);
or U6095 (N_6095,N_4842,N_5074);
and U6096 (N_6096,N_5364,N_4966);
and U6097 (N_6097,N_5059,N_5314);
nor U6098 (N_6098,N_4840,N_5366);
nor U6099 (N_6099,N_5225,N_5023);
nand U6100 (N_6100,N_5248,N_5214);
and U6101 (N_6101,N_5511,N_5467);
nor U6102 (N_6102,N_5586,N_5308);
nor U6103 (N_6103,N_4817,N_5129);
and U6104 (N_6104,N_5095,N_5297);
nor U6105 (N_6105,N_5133,N_5277);
nor U6106 (N_6106,N_5340,N_4839);
nand U6107 (N_6107,N_5059,N_4867);
or U6108 (N_6108,N_5213,N_5559);
nor U6109 (N_6109,N_4894,N_5421);
nand U6110 (N_6110,N_5336,N_5168);
or U6111 (N_6111,N_5493,N_4962);
and U6112 (N_6112,N_5341,N_5371);
and U6113 (N_6113,N_5093,N_4944);
xnor U6114 (N_6114,N_5216,N_5422);
nand U6115 (N_6115,N_5171,N_5287);
and U6116 (N_6116,N_5449,N_5409);
or U6117 (N_6117,N_5089,N_5448);
nor U6118 (N_6118,N_4828,N_4964);
or U6119 (N_6119,N_5528,N_5003);
or U6120 (N_6120,N_4972,N_5339);
and U6121 (N_6121,N_5113,N_4957);
nor U6122 (N_6122,N_4868,N_4971);
and U6123 (N_6123,N_5499,N_5524);
or U6124 (N_6124,N_4926,N_5387);
nor U6125 (N_6125,N_5170,N_5200);
nor U6126 (N_6126,N_5208,N_5346);
nor U6127 (N_6127,N_5362,N_5172);
or U6128 (N_6128,N_5056,N_5567);
and U6129 (N_6129,N_5526,N_5018);
nand U6130 (N_6130,N_5151,N_4863);
and U6131 (N_6131,N_5223,N_4977);
nor U6132 (N_6132,N_5329,N_5086);
nor U6133 (N_6133,N_4883,N_5069);
xor U6134 (N_6134,N_4838,N_4834);
or U6135 (N_6135,N_5208,N_5398);
nor U6136 (N_6136,N_5079,N_4885);
and U6137 (N_6137,N_5334,N_5384);
and U6138 (N_6138,N_5495,N_5558);
nor U6139 (N_6139,N_5375,N_4843);
nand U6140 (N_6140,N_5395,N_5015);
and U6141 (N_6141,N_4858,N_5176);
xnor U6142 (N_6142,N_5333,N_5324);
xnor U6143 (N_6143,N_4983,N_5285);
nand U6144 (N_6144,N_5094,N_4852);
nor U6145 (N_6145,N_5279,N_4920);
nand U6146 (N_6146,N_4916,N_4851);
and U6147 (N_6147,N_4990,N_5387);
or U6148 (N_6148,N_5250,N_5004);
nor U6149 (N_6149,N_5251,N_4853);
xor U6150 (N_6150,N_4834,N_5089);
and U6151 (N_6151,N_4831,N_5339);
nor U6152 (N_6152,N_5355,N_5029);
or U6153 (N_6153,N_4892,N_4870);
nor U6154 (N_6154,N_5126,N_5170);
or U6155 (N_6155,N_5329,N_5078);
nor U6156 (N_6156,N_5410,N_5249);
xnor U6157 (N_6157,N_5563,N_5163);
or U6158 (N_6158,N_5165,N_5310);
xnor U6159 (N_6159,N_4808,N_4917);
or U6160 (N_6160,N_5252,N_5214);
nand U6161 (N_6161,N_5123,N_5257);
xnor U6162 (N_6162,N_5283,N_5493);
and U6163 (N_6163,N_5075,N_5014);
or U6164 (N_6164,N_5224,N_5231);
and U6165 (N_6165,N_5255,N_4929);
nand U6166 (N_6166,N_5574,N_5327);
nor U6167 (N_6167,N_5403,N_4893);
nor U6168 (N_6168,N_5309,N_5301);
nand U6169 (N_6169,N_4919,N_5160);
nor U6170 (N_6170,N_5482,N_5315);
nor U6171 (N_6171,N_4839,N_5117);
and U6172 (N_6172,N_5041,N_5215);
nor U6173 (N_6173,N_4970,N_5240);
and U6174 (N_6174,N_4962,N_5379);
nor U6175 (N_6175,N_4877,N_5571);
or U6176 (N_6176,N_5074,N_5077);
or U6177 (N_6177,N_5316,N_4996);
nand U6178 (N_6178,N_5163,N_5110);
or U6179 (N_6179,N_5134,N_5059);
or U6180 (N_6180,N_5436,N_5472);
nor U6181 (N_6181,N_5204,N_5312);
nor U6182 (N_6182,N_5506,N_4867);
nor U6183 (N_6183,N_5153,N_5490);
or U6184 (N_6184,N_5595,N_5561);
xnor U6185 (N_6185,N_5531,N_5071);
xnor U6186 (N_6186,N_5297,N_4838);
and U6187 (N_6187,N_5206,N_4941);
xnor U6188 (N_6188,N_5007,N_5335);
or U6189 (N_6189,N_5352,N_4889);
and U6190 (N_6190,N_5213,N_5435);
nor U6191 (N_6191,N_5088,N_5308);
xnor U6192 (N_6192,N_4845,N_4848);
and U6193 (N_6193,N_5480,N_5131);
nand U6194 (N_6194,N_5261,N_5473);
nor U6195 (N_6195,N_5252,N_5048);
nor U6196 (N_6196,N_5059,N_4988);
and U6197 (N_6197,N_5435,N_5221);
or U6198 (N_6198,N_5148,N_5173);
nand U6199 (N_6199,N_5042,N_5273);
or U6200 (N_6200,N_5196,N_5178);
and U6201 (N_6201,N_5243,N_4902);
and U6202 (N_6202,N_4995,N_5078);
nand U6203 (N_6203,N_5321,N_4813);
nor U6204 (N_6204,N_4923,N_5527);
and U6205 (N_6205,N_5488,N_4874);
and U6206 (N_6206,N_5286,N_5358);
nand U6207 (N_6207,N_5497,N_5477);
nand U6208 (N_6208,N_5221,N_5394);
and U6209 (N_6209,N_5361,N_5523);
or U6210 (N_6210,N_5402,N_5564);
xor U6211 (N_6211,N_4870,N_5293);
xor U6212 (N_6212,N_5436,N_4984);
or U6213 (N_6213,N_5170,N_5322);
or U6214 (N_6214,N_4821,N_5297);
xnor U6215 (N_6215,N_5115,N_4945);
and U6216 (N_6216,N_5038,N_5235);
xnor U6217 (N_6217,N_5413,N_4979);
xor U6218 (N_6218,N_5133,N_4946);
or U6219 (N_6219,N_5497,N_5450);
nor U6220 (N_6220,N_5127,N_5093);
xor U6221 (N_6221,N_5008,N_4969);
and U6222 (N_6222,N_5164,N_4972);
nor U6223 (N_6223,N_5402,N_4863);
xor U6224 (N_6224,N_5453,N_5150);
xnor U6225 (N_6225,N_4910,N_5110);
nor U6226 (N_6226,N_4933,N_5068);
xnor U6227 (N_6227,N_5317,N_5253);
or U6228 (N_6228,N_5127,N_5400);
nor U6229 (N_6229,N_5389,N_5039);
nor U6230 (N_6230,N_5571,N_5000);
or U6231 (N_6231,N_5061,N_4935);
nand U6232 (N_6232,N_5531,N_5028);
nor U6233 (N_6233,N_5272,N_4886);
or U6234 (N_6234,N_4806,N_5202);
xor U6235 (N_6235,N_5136,N_4923);
or U6236 (N_6236,N_5223,N_4825);
nor U6237 (N_6237,N_5035,N_5053);
nand U6238 (N_6238,N_4840,N_5499);
nand U6239 (N_6239,N_4832,N_4962);
and U6240 (N_6240,N_5187,N_5491);
nand U6241 (N_6241,N_4986,N_5007);
and U6242 (N_6242,N_4883,N_4815);
or U6243 (N_6243,N_5214,N_5363);
and U6244 (N_6244,N_5569,N_5220);
and U6245 (N_6245,N_5532,N_5423);
nand U6246 (N_6246,N_4847,N_5589);
nand U6247 (N_6247,N_5577,N_4989);
or U6248 (N_6248,N_5479,N_5428);
or U6249 (N_6249,N_5263,N_5013);
nor U6250 (N_6250,N_5067,N_5030);
and U6251 (N_6251,N_5461,N_4861);
or U6252 (N_6252,N_5570,N_4889);
and U6253 (N_6253,N_4982,N_5102);
nor U6254 (N_6254,N_4943,N_5117);
nor U6255 (N_6255,N_5450,N_4975);
and U6256 (N_6256,N_5258,N_5099);
xor U6257 (N_6257,N_4996,N_5299);
and U6258 (N_6258,N_4857,N_5549);
and U6259 (N_6259,N_4921,N_5067);
or U6260 (N_6260,N_5409,N_5565);
xnor U6261 (N_6261,N_5481,N_4925);
xnor U6262 (N_6262,N_5312,N_5038);
and U6263 (N_6263,N_5141,N_5200);
nand U6264 (N_6264,N_4877,N_5424);
or U6265 (N_6265,N_5363,N_5018);
nand U6266 (N_6266,N_5376,N_5151);
or U6267 (N_6267,N_5451,N_5166);
xnor U6268 (N_6268,N_4915,N_5209);
xnor U6269 (N_6269,N_5178,N_5409);
or U6270 (N_6270,N_5415,N_5017);
xor U6271 (N_6271,N_5341,N_5177);
nor U6272 (N_6272,N_5193,N_5127);
nor U6273 (N_6273,N_5030,N_4900);
xor U6274 (N_6274,N_5534,N_5028);
nand U6275 (N_6275,N_5035,N_5019);
or U6276 (N_6276,N_5326,N_5441);
or U6277 (N_6277,N_5555,N_5050);
nand U6278 (N_6278,N_4972,N_4950);
xnor U6279 (N_6279,N_5070,N_4903);
or U6280 (N_6280,N_5266,N_4952);
and U6281 (N_6281,N_4922,N_4878);
xnor U6282 (N_6282,N_5519,N_5309);
and U6283 (N_6283,N_4887,N_5597);
xor U6284 (N_6284,N_5238,N_5586);
xnor U6285 (N_6285,N_5586,N_5526);
nor U6286 (N_6286,N_5553,N_4939);
and U6287 (N_6287,N_5089,N_5148);
nor U6288 (N_6288,N_5349,N_5092);
and U6289 (N_6289,N_5344,N_4865);
and U6290 (N_6290,N_4990,N_5474);
nor U6291 (N_6291,N_5352,N_4973);
nor U6292 (N_6292,N_5354,N_4819);
or U6293 (N_6293,N_5372,N_5262);
xnor U6294 (N_6294,N_5135,N_5077);
or U6295 (N_6295,N_5314,N_5516);
and U6296 (N_6296,N_5545,N_5216);
nor U6297 (N_6297,N_5542,N_4822);
nor U6298 (N_6298,N_5082,N_5406);
xor U6299 (N_6299,N_4991,N_5462);
or U6300 (N_6300,N_5596,N_5093);
and U6301 (N_6301,N_5262,N_5271);
nor U6302 (N_6302,N_5403,N_5307);
nand U6303 (N_6303,N_5312,N_5025);
or U6304 (N_6304,N_5528,N_5060);
or U6305 (N_6305,N_5366,N_4947);
xnor U6306 (N_6306,N_4851,N_5146);
or U6307 (N_6307,N_4815,N_5133);
xor U6308 (N_6308,N_4847,N_5242);
xor U6309 (N_6309,N_5349,N_5509);
nor U6310 (N_6310,N_5340,N_5110);
or U6311 (N_6311,N_4881,N_5075);
or U6312 (N_6312,N_5379,N_5090);
nand U6313 (N_6313,N_4817,N_5309);
and U6314 (N_6314,N_5083,N_4905);
or U6315 (N_6315,N_5450,N_4832);
or U6316 (N_6316,N_4975,N_5255);
or U6317 (N_6317,N_5367,N_5284);
nor U6318 (N_6318,N_5238,N_5435);
xor U6319 (N_6319,N_5101,N_4988);
xnor U6320 (N_6320,N_5307,N_5502);
nand U6321 (N_6321,N_4959,N_5235);
or U6322 (N_6322,N_5391,N_5023);
xor U6323 (N_6323,N_5297,N_5456);
nor U6324 (N_6324,N_5499,N_5370);
nand U6325 (N_6325,N_5536,N_5348);
and U6326 (N_6326,N_4981,N_5150);
xnor U6327 (N_6327,N_4942,N_4934);
nor U6328 (N_6328,N_5166,N_5023);
and U6329 (N_6329,N_5522,N_5195);
xor U6330 (N_6330,N_5391,N_5503);
nand U6331 (N_6331,N_5068,N_5311);
or U6332 (N_6332,N_5384,N_4927);
xor U6333 (N_6333,N_5418,N_5106);
and U6334 (N_6334,N_5114,N_5383);
or U6335 (N_6335,N_4941,N_5160);
nor U6336 (N_6336,N_5261,N_5575);
or U6337 (N_6337,N_5095,N_5354);
xnor U6338 (N_6338,N_5472,N_5049);
or U6339 (N_6339,N_4814,N_4954);
nand U6340 (N_6340,N_4824,N_5480);
or U6341 (N_6341,N_5592,N_5280);
xor U6342 (N_6342,N_5414,N_5157);
or U6343 (N_6343,N_5096,N_5457);
and U6344 (N_6344,N_5254,N_5577);
nor U6345 (N_6345,N_4915,N_4878);
and U6346 (N_6346,N_5439,N_5444);
and U6347 (N_6347,N_5112,N_5109);
and U6348 (N_6348,N_5528,N_5426);
or U6349 (N_6349,N_5179,N_4913);
xnor U6350 (N_6350,N_5366,N_5049);
xor U6351 (N_6351,N_5154,N_4814);
nand U6352 (N_6352,N_4988,N_5187);
and U6353 (N_6353,N_5155,N_5104);
and U6354 (N_6354,N_5267,N_4806);
nand U6355 (N_6355,N_5076,N_5343);
nand U6356 (N_6356,N_5067,N_5331);
and U6357 (N_6357,N_5446,N_4987);
and U6358 (N_6358,N_5216,N_5498);
nor U6359 (N_6359,N_5165,N_4985);
or U6360 (N_6360,N_5116,N_5464);
or U6361 (N_6361,N_5306,N_5590);
nand U6362 (N_6362,N_5093,N_5477);
nor U6363 (N_6363,N_5255,N_5441);
and U6364 (N_6364,N_4928,N_4920);
nor U6365 (N_6365,N_5234,N_5089);
and U6366 (N_6366,N_5514,N_4856);
and U6367 (N_6367,N_5493,N_5174);
nand U6368 (N_6368,N_4903,N_5551);
xor U6369 (N_6369,N_4803,N_4872);
nor U6370 (N_6370,N_5576,N_5237);
nand U6371 (N_6371,N_5259,N_5218);
nor U6372 (N_6372,N_4959,N_5190);
nor U6373 (N_6373,N_4901,N_5046);
or U6374 (N_6374,N_5483,N_5577);
xor U6375 (N_6375,N_4806,N_5254);
and U6376 (N_6376,N_5456,N_5065);
or U6377 (N_6377,N_5414,N_5011);
and U6378 (N_6378,N_5297,N_4805);
or U6379 (N_6379,N_5356,N_4943);
xnor U6380 (N_6380,N_5284,N_5290);
and U6381 (N_6381,N_4898,N_5569);
or U6382 (N_6382,N_5229,N_5526);
nor U6383 (N_6383,N_5473,N_4832);
nor U6384 (N_6384,N_5091,N_5454);
nand U6385 (N_6385,N_5205,N_5587);
xor U6386 (N_6386,N_5178,N_5002);
and U6387 (N_6387,N_5558,N_4890);
xor U6388 (N_6388,N_4932,N_5182);
nor U6389 (N_6389,N_5391,N_5193);
or U6390 (N_6390,N_5483,N_5347);
or U6391 (N_6391,N_5372,N_5574);
nor U6392 (N_6392,N_4935,N_5500);
and U6393 (N_6393,N_4989,N_4926);
nor U6394 (N_6394,N_5335,N_5133);
or U6395 (N_6395,N_5327,N_5202);
nand U6396 (N_6396,N_5201,N_5149);
nand U6397 (N_6397,N_5323,N_4903);
or U6398 (N_6398,N_5168,N_5401);
nand U6399 (N_6399,N_5526,N_5388);
or U6400 (N_6400,N_5773,N_6217);
nor U6401 (N_6401,N_5900,N_6139);
nor U6402 (N_6402,N_6348,N_6282);
nor U6403 (N_6403,N_5811,N_5674);
and U6404 (N_6404,N_5887,N_5766);
nor U6405 (N_6405,N_5838,N_6198);
and U6406 (N_6406,N_5784,N_6024);
nand U6407 (N_6407,N_5851,N_6055);
nor U6408 (N_6408,N_5700,N_6357);
nor U6409 (N_6409,N_5643,N_5956);
or U6410 (N_6410,N_5721,N_5614);
nor U6411 (N_6411,N_6241,N_5878);
nand U6412 (N_6412,N_5926,N_5948);
or U6413 (N_6413,N_6371,N_5659);
nand U6414 (N_6414,N_6222,N_5911);
and U6415 (N_6415,N_5819,N_6208);
and U6416 (N_6416,N_5860,N_5769);
and U6417 (N_6417,N_5697,N_6209);
and U6418 (N_6418,N_6016,N_6324);
or U6419 (N_6419,N_6039,N_5967);
nand U6420 (N_6420,N_5994,N_6376);
or U6421 (N_6421,N_6332,N_6331);
or U6422 (N_6422,N_5861,N_5868);
or U6423 (N_6423,N_6172,N_5881);
nor U6424 (N_6424,N_6220,N_6227);
nand U6425 (N_6425,N_5915,N_5685);
nand U6426 (N_6426,N_5826,N_5934);
nand U6427 (N_6427,N_6247,N_5632);
and U6428 (N_6428,N_5693,N_6010);
nor U6429 (N_6429,N_5699,N_6078);
and U6430 (N_6430,N_5706,N_6391);
or U6431 (N_6431,N_6070,N_6344);
and U6432 (N_6432,N_6022,N_5722);
and U6433 (N_6433,N_5783,N_5607);
or U6434 (N_6434,N_6291,N_6216);
nand U6435 (N_6435,N_5741,N_6360);
or U6436 (N_6436,N_6113,N_5651);
or U6437 (N_6437,N_5715,N_5837);
nor U6438 (N_6438,N_6298,N_6012);
nand U6439 (N_6439,N_5831,N_5802);
and U6440 (N_6440,N_5758,N_6118);
nor U6441 (N_6441,N_6109,N_6119);
and U6442 (N_6442,N_6228,N_6099);
nand U6443 (N_6443,N_5919,N_6148);
and U6444 (N_6444,N_6342,N_5797);
nand U6445 (N_6445,N_6105,N_6133);
nor U6446 (N_6446,N_6037,N_5663);
and U6447 (N_6447,N_6242,N_5680);
or U6448 (N_6448,N_5692,N_6058);
nand U6449 (N_6449,N_6085,N_6128);
nand U6450 (N_6450,N_5941,N_6047);
xnor U6451 (N_6451,N_6355,N_5820);
nand U6452 (N_6452,N_6294,N_5991);
and U6453 (N_6453,N_5937,N_6062);
and U6454 (N_6454,N_5684,N_6006);
nand U6455 (N_6455,N_6056,N_6168);
nand U6456 (N_6456,N_5631,N_5818);
xor U6457 (N_6457,N_6243,N_5929);
nor U6458 (N_6458,N_5719,N_6284);
or U6459 (N_6459,N_5654,N_6397);
nand U6460 (N_6460,N_6143,N_5673);
nand U6461 (N_6461,N_6286,N_6252);
xor U6462 (N_6462,N_6175,N_6005);
nor U6463 (N_6463,N_6203,N_6102);
and U6464 (N_6464,N_6015,N_6165);
nor U6465 (N_6465,N_5622,N_6347);
and U6466 (N_6466,N_6211,N_5872);
nor U6467 (N_6467,N_5918,N_5609);
nand U6468 (N_6468,N_6383,N_5809);
and U6469 (N_6469,N_6138,N_5910);
nand U6470 (N_6470,N_6004,N_6221);
nand U6471 (N_6471,N_5730,N_6270);
and U6472 (N_6472,N_5920,N_5795);
xnor U6473 (N_6473,N_5701,N_6094);
or U6474 (N_6474,N_6303,N_6180);
nand U6475 (N_6475,N_5671,N_6275);
and U6476 (N_6476,N_5804,N_5833);
nor U6477 (N_6477,N_5738,N_5914);
nand U6478 (N_6478,N_5902,N_5862);
or U6479 (N_6479,N_5890,N_6396);
or U6480 (N_6480,N_6363,N_6301);
nand U6481 (N_6481,N_5984,N_5857);
xnor U6482 (N_6482,N_6269,N_5896);
or U6483 (N_6483,N_6368,N_5989);
or U6484 (N_6484,N_5966,N_6153);
xor U6485 (N_6485,N_5814,N_5798);
and U6486 (N_6486,N_5633,N_5964);
nor U6487 (N_6487,N_6087,N_5807);
and U6488 (N_6488,N_5664,N_5774);
nand U6489 (N_6489,N_6028,N_5959);
nand U6490 (N_6490,N_5874,N_6224);
or U6491 (N_6491,N_6213,N_6090);
nand U6492 (N_6492,N_5785,N_6356);
and U6493 (N_6493,N_5618,N_5873);
and U6494 (N_6494,N_5749,N_5679);
xnor U6495 (N_6495,N_6170,N_5825);
nor U6496 (N_6496,N_5772,N_5875);
nor U6497 (N_6497,N_6374,N_5955);
nor U6498 (N_6498,N_6382,N_6395);
or U6499 (N_6499,N_6378,N_6189);
nor U6500 (N_6500,N_6021,N_6292);
xor U6501 (N_6501,N_5880,N_6129);
xor U6502 (N_6502,N_5672,N_6364);
xor U6503 (N_6503,N_6197,N_6136);
nand U6504 (N_6504,N_5969,N_6349);
xor U6505 (N_6505,N_6163,N_6183);
nor U6506 (N_6506,N_5897,N_6326);
or U6507 (N_6507,N_6132,N_5757);
nand U6508 (N_6508,N_6256,N_5615);
and U6509 (N_6509,N_6023,N_5778);
or U6510 (N_6510,N_5626,N_6293);
nand U6511 (N_6511,N_6174,N_6315);
nor U6512 (N_6512,N_5962,N_6333);
nor U6513 (N_6513,N_5829,N_6035);
nand U6514 (N_6514,N_5817,N_6092);
or U6515 (N_6515,N_6142,N_5888);
xor U6516 (N_6516,N_6323,N_6343);
nor U6517 (N_6517,N_5950,N_5657);
nor U6518 (N_6518,N_5762,N_5999);
and U6519 (N_6519,N_6290,N_5761);
nand U6520 (N_6520,N_5763,N_6299);
nor U6521 (N_6521,N_6394,N_5736);
nand U6522 (N_6522,N_6018,N_6130);
xor U6523 (N_6523,N_5616,N_5927);
nor U6524 (N_6524,N_6025,N_5666);
nand U6525 (N_6525,N_5695,N_6073);
xnor U6526 (N_6526,N_6060,N_6111);
and U6527 (N_6527,N_5940,N_5709);
or U6528 (N_6528,N_5752,N_5648);
nand U6529 (N_6529,N_5885,N_5961);
or U6530 (N_6530,N_6193,N_6244);
nor U6531 (N_6531,N_6160,N_6246);
nor U6532 (N_6532,N_5822,N_5726);
or U6533 (N_6533,N_5960,N_6384);
xnor U6534 (N_6534,N_6151,N_5755);
nand U6535 (N_6535,N_5775,N_5863);
nand U6536 (N_6536,N_6317,N_5655);
xnor U6537 (N_6537,N_5740,N_5602);
nand U6538 (N_6538,N_6013,N_5720);
and U6539 (N_6539,N_6366,N_5690);
or U6540 (N_6540,N_5662,N_5746);
or U6541 (N_6541,N_6322,N_6135);
and U6542 (N_6542,N_6300,N_6314);
nand U6543 (N_6543,N_6386,N_6319);
nor U6544 (N_6544,N_5751,N_5904);
nor U6545 (N_6545,N_5906,N_5728);
xnor U6546 (N_6546,N_5658,N_5650);
and U6547 (N_6547,N_6184,N_6365);
or U6548 (N_6548,N_6179,N_6069);
and U6549 (N_6549,N_6036,N_5899);
nor U6550 (N_6550,N_6271,N_6181);
or U6551 (N_6551,N_5993,N_5938);
nand U6552 (N_6552,N_6166,N_6223);
xor U6553 (N_6553,N_6276,N_6178);
nor U6554 (N_6554,N_6097,N_6051);
nand U6555 (N_6555,N_6390,N_6232);
nand U6556 (N_6556,N_5976,N_6145);
nor U6557 (N_6557,N_5908,N_6158);
nand U6558 (N_6558,N_6057,N_6255);
xnor U6559 (N_6559,N_6007,N_6274);
and U6560 (N_6560,N_5889,N_5661);
xor U6561 (N_6561,N_6379,N_6345);
and U6562 (N_6562,N_6117,N_6091);
or U6563 (N_6563,N_6154,N_5744);
xnor U6564 (N_6564,N_5792,N_5641);
or U6565 (N_6565,N_6144,N_6079);
xnor U6566 (N_6566,N_6235,N_6038);
xor U6567 (N_6567,N_5852,N_6086);
xor U6568 (N_6568,N_5733,N_5942);
xor U6569 (N_6569,N_5828,N_5821);
and U6570 (N_6570,N_5882,N_5979);
or U6571 (N_6571,N_5723,N_5779);
xor U6572 (N_6572,N_6202,N_5786);
and U6573 (N_6573,N_6065,N_5714);
or U6574 (N_6574,N_5704,N_5789);
nand U6575 (N_6575,N_5869,N_5977);
and U6576 (N_6576,N_5776,N_5619);
nor U6577 (N_6577,N_6176,N_5970);
xnor U6578 (N_6578,N_5854,N_5988);
nand U6579 (N_6579,N_5803,N_5905);
or U6580 (N_6580,N_5947,N_5691);
and U6581 (N_6581,N_5639,N_6054);
xor U6582 (N_6582,N_6044,N_5806);
and U6583 (N_6583,N_6265,N_6340);
or U6584 (N_6584,N_6103,N_6104);
nand U6585 (N_6585,N_6327,N_5689);
or U6586 (N_6586,N_5865,N_6389);
nand U6587 (N_6587,N_6000,N_5844);
or U6588 (N_6588,N_5925,N_6083);
or U6589 (N_6589,N_5637,N_6393);
nor U6590 (N_6590,N_6240,N_5907);
xnor U6591 (N_6591,N_5973,N_5743);
xnor U6592 (N_6592,N_5858,N_6280);
and U6593 (N_6593,N_5933,N_5954);
or U6594 (N_6594,N_5971,N_5997);
or U6595 (N_6595,N_6249,N_5638);
nand U6596 (N_6596,N_5676,N_5670);
or U6597 (N_6597,N_6030,N_6359);
and U6598 (N_6598,N_6272,N_6146);
and U6599 (N_6599,N_6115,N_6122);
or U6600 (N_6600,N_6077,N_5866);
xnor U6601 (N_6601,N_5856,N_6302);
xor U6602 (N_6602,N_5770,N_5711);
nand U6603 (N_6603,N_6306,N_5793);
nand U6604 (N_6604,N_5739,N_5982);
xor U6605 (N_6605,N_5936,N_5600);
nand U6606 (N_6606,N_5836,N_6031);
nor U6607 (N_6607,N_6110,N_6050);
nor U6608 (N_6608,N_5879,N_6321);
nor U6609 (N_6609,N_5777,N_5805);
xnor U6610 (N_6610,N_5930,N_6120);
nand U6611 (N_6611,N_6066,N_5696);
xor U6612 (N_6612,N_5725,N_5895);
and U6613 (N_6613,N_5943,N_6096);
xor U6614 (N_6614,N_6351,N_6074);
and U6615 (N_6615,N_5644,N_6149);
and U6616 (N_6616,N_5612,N_6226);
nor U6617 (N_6617,N_6173,N_6034);
xnor U6618 (N_6618,N_6072,N_6019);
nand U6619 (N_6619,N_6212,N_5742);
or U6620 (N_6620,N_5986,N_5710);
nor U6621 (N_6621,N_5909,N_5601);
nor U6622 (N_6622,N_6352,N_6116);
and U6623 (N_6623,N_6134,N_5617);
nor U6624 (N_6624,N_6338,N_6201);
nor U6625 (N_6625,N_5951,N_5678);
nand U6626 (N_6626,N_6081,N_6215);
xor U6627 (N_6627,N_5705,N_5767);
xor U6628 (N_6628,N_5898,N_5808);
or U6629 (N_6629,N_6237,N_6353);
nand U6630 (N_6630,N_5703,N_6182);
xnor U6631 (N_6631,N_6277,N_5894);
nor U6632 (N_6632,N_6273,N_6093);
nand U6633 (N_6633,N_5974,N_5634);
or U6634 (N_6634,N_6218,N_5735);
nand U6635 (N_6635,N_6095,N_6307);
and U6636 (N_6636,N_6325,N_6191);
or U6637 (N_6637,N_5965,N_6040);
or U6638 (N_6638,N_6288,N_6289);
nor U6639 (N_6639,N_5756,N_6380);
or U6640 (N_6640,N_5669,N_6002);
xor U6641 (N_6641,N_6229,N_6046);
or U6642 (N_6642,N_5613,N_5791);
nand U6643 (N_6643,N_5698,N_6192);
xnor U6644 (N_6644,N_6346,N_6126);
nand U6645 (N_6645,N_6049,N_6084);
nand U6646 (N_6646,N_6250,N_6125);
nor U6647 (N_6647,N_5886,N_5625);
xnor U6648 (N_6648,N_5708,N_6210);
xnor U6649 (N_6649,N_6388,N_6231);
nor U6650 (N_6650,N_5635,N_5913);
and U6651 (N_6651,N_5611,N_5687);
nor U6652 (N_6652,N_6329,N_5732);
xnor U6653 (N_6653,N_5760,N_5653);
nor U6654 (N_6654,N_5668,N_6313);
nand U6655 (N_6655,N_6304,N_5975);
or U6656 (N_6656,N_6124,N_6098);
nand U6657 (N_6657,N_6205,N_5620);
xor U6658 (N_6658,N_6266,N_5652);
nand U6659 (N_6659,N_6296,N_6042);
and U6660 (N_6660,N_6233,N_5953);
xor U6661 (N_6661,N_5765,N_5848);
and U6662 (N_6662,N_6032,N_6195);
nor U6663 (N_6663,N_6358,N_6064);
nand U6664 (N_6664,N_6381,N_6337);
nand U6665 (N_6665,N_6200,N_5627);
and U6666 (N_6666,N_5630,N_6239);
and U6667 (N_6667,N_5884,N_5922);
xor U6668 (N_6668,N_5642,N_6370);
nor U6669 (N_6669,N_5623,N_6354);
xnor U6670 (N_6670,N_6279,N_6067);
nor U6671 (N_6671,N_5995,N_6372);
and U6672 (N_6672,N_5813,N_6141);
nor U6673 (N_6673,N_5771,N_6339);
or U6674 (N_6674,N_5846,N_6263);
and U6675 (N_6675,N_5605,N_5753);
nor U6676 (N_6676,N_5794,N_5647);
xor U6677 (N_6677,N_5675,N_5870);
nand U6678 (N_6678,N_5843,N_5688);
xor U6679 (N_6679,N_6234,N_5853);
or U6680 (N_6680,N_6157,N_5608);
or U6681 (N_6681,N_5629,N_6059);
and U6682 (N_6682,N_6254,N_6398);
and U6683 (N_6683,N_5864,N_5972);
and U6684 (N_6684,N_6330,N_6137);
xnor U6685 (N_6685,N_6207,N_5610);
or U6686 (N_6686,N_6335,N_5646);
nand U6687 (N_6687,N_6045,N_6107);
or U6688 (N_6688,N_6068,N_5624);
nor U6689 (N_6689,N_5801,N_5781);
nand U6690 (N_6690,N_6320,N_6162);
or U6691 (N_6691,N_6308,N_6199);
or U6692 (N_6692,N_5985,N_5747);
and U6693 (N_6693,N_5978,N_5716);
and U6694 (N_6694,N_5656,N_5963);
nand U6695 (N_6695,N_5702,N_6219);
and U6696 (N_6696,N_5901,N_6258);
nand U6697 (N_6697,N_6140,N_6262);
nand U6698 (N_6698,N_5799,N_6225);
or U6699 (N_6699,N_6147,N_6101);
nand U6700 (N_6700,N_6281,N_5754);
or U6701 (N_6701,N_5935,N_6267);
xnor U6702 (N_6702,N_5677,N_6385);
and U6703 (N_6703,N_5892,N_6186);
or U6704 (N_6704,N_6108,N_6043);
nor U6705 (N_6705,N_6399,N_6011);
xnor U6706 (N_6706,N_6114,N_6373);
nand U6707 (N_6707,N_5621,N_5945);
xnor U6708 (N_6708,N_5731,N_6251);
nand U6709 (N_6709,N_6361,N_6316);
nor U6710 (N_6710,N_6230,N_5737);
xnor U6711 (N_6711,N_6261,N_5928);
xor U6712 (N_6712,N_5812,N_6089);
and U6713 (N_6713,N_6009,N_5916);
or U6714 (N_6714,N_5847,N_6196);
xor U6715 (N_6715,N_5745,N_5796);
or U6716 (N_6716,N_5823,N_6100);
xnor U6717 (N_6717,N_5917,N_6268);
nor U6718 (N_6718,N_5727,N_6159);
nand U6719 (N_6719,N_6260,N_5724);
nor U6720 (N_6720,N_6253,N_6334);
xor U6721 (N_6721,N_6127,N_5603);
and U6722 (N_6722,N_6156,N_6369);
or U6723 (N_6723,N_5717,N_6214);
nor U6724 (N_6724,N_6312,N_6053);
xnor U6725 (N_6725,N_6106,N_6190);
nand U6726 (N_6726,N_5983,N_6367);
and U6727 (N_6727,N_5859,N_5958);
nor U6728 (N_6728,N_6029,N_5729);
nor U6729 (N_6729,N_5712,N_6052);
and U6730 (N_6730,N_6309,N_5891);
nor U6731 (N_6731,N_5944,N_6375);
and U6732 (N_6732,N_5604,N_5759);
nand U6733 (N_6733,N_6033,N_6112);
nor U6734 (N_6734,N_5946,N_6026);
or U6735 (N_6735,N_6283,N_6310);
nor U6736 (N_6736,N_5840,N_5628);
nand U6737 (N_6737,N_5924,N_6187);
nor U6738 (N_6738,N_5782,N_6063);
and U6739 (N_6739,N_6003,N_6121);
nand U6740 (N_6740,N_6167,N_6071);
xor U6741 (N_6741,N_5718,N_5665);
nand U6742 (N_6742,N_5876,N_6264);
or U6743 (N_6743,N_5734,N_5877);
or U6744 (N_6744,N_5686,N_6020);
or U6745 (N_6745,N_6171,N_6177);
and U6746 (N_6746,N_6204,N_5842);
nor U6747 (N_6747,N_5834,N_5867);
or U6748 (N_6748,N_5981,N_6238);
and U6749 (N_6749,N_5640,N_6350);
xnor U6750 (N_6750,N_6236,N_6123);
nand U6751 (N_6751,N_5903,N_5790);
nand U6752 (N_6752,N_6305,N_6075);
nand U6753 (N_6753,N_5816,N_6377);
xnor U6754 (N_6754,N_5839,N_6080);
nor U6755 (N_6755,N_5931,N_5939);
nor U6756 (N_6756,N_5824,N_6027);
xor U6757 (N_6757,N_6001,N_5992);
nand U6758 (N_6758,N_6362,N_5968);
nand U6759 (N_6759,N_5682,N_5713);
nand U6760 (N_6760,N_6061,N_5683);
xor U6761 (N_6761,N_5980,N_6008);
or U6762 (N_6762,N_5681,N_5957);
nor U6763 (N_6763,N_5827,N_6082);
and U6764 (N_6764,N_6287,N_5990);
and U6765 (N_6765,N_5694,N_6088);
nand U6766 (N_6766,N_5815,N_6259);
nor U6767 (N_6767,N_6257,N_5949);
nand U6768 (N_6768,N_6131,N_6169);
or U6769 (N_6769,N_5645,N_6188);
nand U6770 (N_6770,N_5845,N_6017);
or U6771 (N_6771,N_5912,N_5660);
xor U6772 (N_6772,N_6041,N_5841);
nor U6773 (N_6773,N_6295,N_5832);
nor U6774 (N_6774,N_6248,N_6164);
and U6775 (N_6775,N_6185,N_5996);
nand U6776 (N_6776,N_6318,N_5800);
xor U6777 (N_6777,N_6392,N_5923);
or U6778 (N_6778,N_6311,N_5883);
or U6779 (N_6779,N_5998,N_6285);
nand U6780 (N_6780,N_6297,N_5750);
nor U6781 (N_6781,N_5748,N_5788);
nand U6782 (N_6782,N_6387,N_5921);
or U6783 (N_6783,N_5667,N_5830);
nor U6784 (N_6784,N_5768,N_6076);
nor U6785 (N_6785,N_6341,N_6245);
nand U6786 (N_6786,N_5835,N_5893);
or U6787 (N_6787,N_5780,N_6194);
nor U6788 (N_6788,N_6206,N_5932);
and U6789 (N_6789,N_6150,N_5952);
xor U6790 (N_6790,N_5636,N_6152);
and U6791 (N_6791,N_5787,N_6014);
xor U6792 (N_6792,N_5606,N_5649);
nand U6793 (N_6793,N_5855,N_5871);
nand U6794 (N_6794,N_6155,N_5987);
nand U6795 (N_6795,N_5850,N_6048);
nand U6796 (N_6796,N_6328,N_6161);
and U6797 (N_6797,N_6336,N_5849);
or U6798 (N_6798,N_5810,N_5764);
nand U6799 (N_6799,N_5707,N_6278);
and U6800 (N_6800,N_5849,N_6357);
xor U6801 (N_6801,N_5718,N_6128);
xnor U6802 (N_6802,N_6213,N_5707);
or U6803 (N_6803,N_6050,N_6279);
or U6804 (N_6804,N_6157,N_6176);
and U6805 (N_6805,N_6073,N_6046);
and U6806 (N_6806,N_6362,N_5909);
or U6807 (N_6807,N_6175,N_6223);
xnor U6808 (N_6808,N_6285,N_6140);
xor U6809 (N_6809,N_5669,N_5694);
xor U6810 (N_6810,N_6384,N_6305);
and U6811 (N_6811,N_5882,N_6314);
nand U6812 (N_6812,N_6378,N_5649);
or U6813 (N_6813,N_6057,N_5685);
xnor U6814 (N_6814,N_5792,N_6298);
or U6815 (N_6815,N_5798,N_6300);
and U6816 (N_6816,N_6277,N_6145);
and U6817 (N_6817,N_5746,N_5724);
nor U6818 (N_6818,N_5704,N_5781);
nand U6819 (N_6819,N_6191,N_5849);
nand U6820 (N_6820,N_5967,N_5654);
nand U6821 (N_6821,N_5774,N_5798);
or U6822 (N_6822,N_6130,N_6071);
xnor U6823 (N_6823,N_5759,N_5986);
or U6824 (N_6824,N_5914,N_5902);
and U6825 (N_6825,N_6296,N_6279);
nand U6826 (N_6826,N_5951,N_6280);
or U6827 (N_6827,N_6316,N_5841);
or U6828 (N_6828,N_6033,N_5973);
nand U6829 (N_6829,N_5888,N_6161);
and U6830 (N_6830,N_5786,N_5600);
and U6831 (N_6831,N_6118,N_5932);
nand U6832 (N_6832,N_6357,N_5755);
xor U6833 (N_6833,N_5799,N_6166);
nand U6834 (N_6834,N_6384,N_5838);
nor U6835 (N_6835,N_5647,N_5830);
or U6836 (N_6836,N_5646,N_6342);
xor U6837 (N_6837,N_6101,N_5843);
nor U6838 (N_6838,N_6100,N_5620);
xor U6839 (N_6839,N_6378,N_6292);
nand U6840 (N_6840,N_5713,N_6142);
nand U6841 (N_6841,N_5738,N_6235);
or U6842 (N_6842,N_6357,N_6163);
nand U6843 (N_6843,N_5715,N_6106);
or U6844 (N_6844,N_6164,N_6268);
or U6845 (N_6845,N_6389,N_6095);
xnor U6846 (N_6846,N_6104,N_5799);
or U6847 (N_6847,N_5967,N_5909);
nor U6848 (N_6848,N_6164,N_6009);
and U6849 (N_6849,N_5807,N_5926);
or U6850 (N_6850,N_6074,N_6155);
or U6851 (N_6851,N_5884,N_5993);
nand U6852 (N_6852,N_5675,N_6334);
xnor U6853 (N_6853,N_5997,N_6060);
nor U6854 (N_6854,N_6069,N_5979);
nand U6855 (N_6855,N_6384,N_6078);
or U6856 (N_6856,N_6254,N_6136);
or U6857 (N_6857,N_6153,N_6131);
nand U6858 (N_6858,N_6005,N_6342);
nand U6859 (N_6859,N_6278,N_6389);
and U6860 (N_6860,N_6271,N_5747);
or U6861 (N_6861,N_6242,N_6006);
nor U6862 (N_6862,N_6373,N_5738);
xor U6863 (N_6863,N_5663,N_6339);
nand U6864 (N_6864,N_6297,N_5885);
nor U6865 (N_6865,N_6307,N_5840);
or U6866 (N_6866,N_6027,N_6081);
nand U6867 (N_6867,N_6137,N_6284);
or U6868 (N_6868,N_6011,N_5989);
nor U6869 (N_6869,N_6361,N_6347);
nand U6870 (N_6870,N_5926,N_6117);
xor U6871 (N_6871,N_5797,N_5885);
xor U6872 (N_6872,N_5705,N_6160);
or U6873 (N_6873,N_5877,N_5799);
nand U6874 (N_6874,N_5813,N_5660);
nand U6875 (N_6875,N_5704,N_6019);
nand U6876 (N_6876,N_5758,N_6004);
nor U6877 (N_6877,N_5744,N_6253);
nand U6878 (N_6878,N_5680,N_6147);
nand U6879 (N_6879,N_5619,N_6038);
or U6880 (N_6880,N_6203,N_5882);
nand U6881 (N_6881,N_5705,N_6279);
xnor U6882 (N_6882,N_6051,N_6000);
or U6883 (N_6883,N_5943,N_6142);
and U6884 (N_6884,N_5819,N_5825);
or U6885 (N_6885,N_5858,N_5673);
or U6886 (N_6886,N_6091,N_6259);
nand U6887 (N_6887,N_5651,N_6352);
and U6888 (N_6888,N_6218,N_6190);
or U6889 (N_6889,N_6079,N_5903);
nand U6890 (N_6890,N_6183,N_5967);
or U6891 (N_6891,N_6017,N_5609);
nand U6892 (N_6892,N_6241,N_6092);
xnor U6893 (N_6893,N_6306,N_6241);
xor U6894 (N_6894,N_6093,N_5788);
nor U6895 (N_6895,N_6230,N_6356);
nand U6896 (N_6896,N_6180,N_6264);
and U6897 (N_6897,N_6199,N_6219);
and U6898 (N_6898,N_6149,N_5650);
nand U6899 (N_6899,N_5603,N_6206);
xnor U6900 (N_6900,N_5887,N_5823);
or U6901 (N_6901,N_6369,N_5988);
nand U6902 (N_6902,N_5949,N_5628);
nor U6903 (N_6903,N_5654,N_5750);
nor U6904 (N_6904,N_6055,N_6281);
nor U6905 (N_6905,N_5690,N_5907);
nand U6906 (N_6906,N_6145,N_5676);
xnor U6907 (N_6907,N_5844,N_5887);
nor U6908 (N_6908,N_6361,N_5604);
xor U6909 (N_6909,N_5873,N_6139);
nor U6910 (N_6910,N_6361,N_6073);
or U6911 (N_6911,N_6157,N_5967);
nor U6912 (N_6912,N_6328,N_5610);
nand U6913 (N_6913,N_5711,N_5614);
nor U6914 (N_6914,N_5866,N_5771);
xnor U6915 (N_6915,N_6286,N_6384);
or U6916 (N_6916,N_5901,N_6010);
and U6917 (N_6917,N_6396,N_6208);
and U6918 (N_6918,N_6216,N_6082);
or U6919 (N_6919,N_5707,N_5796);
xnor U6920 (N_6920,N_5897,N_6308);
nor U6921 (N_6921,N_5817,N_6350);
nand U6922 (N_6922,N_6005,N_6274);
and U6923 (N_6923,N_5657,N_5807);
xor U6924 (N_6924,N_5838,N_6096);
nor U6925 (N_6925,N_5696,N_6335);
nor U6926 (N_6926,N_5750,N_6156);
xnor U6927 (N_6927,N_6088,N_6121);
xor U6928 (N_6928,N_6147,N_6028);
nor U6929 (N_6929,N_6114,N_6116);
and U6930 (N_6930,N_6090,N_6304);
nor U6931 (N_6931,N_5651,N_5950);
nor U6932 (N_6932,N_5637,N_5844);
and U6933 (N_6933,N_6329,N_5664);
nand U6934 (N_6934,N_6106,N_6090);
xor U6935 (N_6935,N_5823,N_6137);
and U6936 (N_6936,N_5958,N_5634);
and U6937 (N_6937,N_5740,N_5677);
and U6938 (N_6938,N_6039,N_5780);
nand U6939 (N_6939,N_5652,N_5825);
nand U6940 (N_6940,N_5640,N_5957);
nand U6941 (N_6941,N_6106,N_6265);
and U6942 (N_6942,N_6361,N_5694);
or U6943 (N_6943,N_6207,N_6074);
or U6944 (N_6944,N_6383,N_5669);
and U6945 (N_6945,N_6108,N_5842);
nor U6946 (N_6946,N_6295,N_6147);
and U6947 (N_6947,N_6023,N_6022);
xnor U6948 (N_6948,N_6040,N_5618);
and U6949 (N_6949,N_6280,N_6234);
nand U6950 (N_6950,N_5646,N_5700);
nor U6951 (N_6951,N_6398,N_5712);
or U6952 (N_6952,N_5997,N_6329);
or U6953 (N_6953,N_5994,N_6354);
nor U6954 (N_6954,N_5735,N_6150);
nor U6955 (N_6955,N_6342,N_5873);
xor U6956 (N_6956,N_5620,N_6238);
and U6957 (N_6957,N_6079,N_6173);
or U6958 (N_6958,N_6324,N_5808);
nand U6959 (N_6959,N_6337,N_5998);
nor U6960 (N_6960,N_6336,N_5832);
nand U6961 (N_6961,N_5885,N_5870);
nand U6962 (N_6962,N_5934,N_5684);
nor U6963 (N_6963,N_6247,N_5990);
nor U6964 (N_6964,N_6313,N_5890);
or U6965 (N_6965,N_6003,N_6377);
or U6966 (N_6966,N_5646,N_5733);
nor U6967 (N_6967,N_6068,N_5818);
or U6968 (N_6968,N_5772,N_6067);
or U6969 (N_6969,N_5789,N_5849);
nand U6970 (N_6970,N_5976,N_5896);
and U6971 (N_6971,N_6094,N_5909);
xnor U6972 (N_6972,N_5649,N_6002);
xor U6973 (N_6973,N_6082,N_5768);
or U6974 (N_6974,N_6130,N_6203);
or U6975 (N_6975,N_6284,N_6269);
or U6976 (N_6976,N_6344,N_5916);
or U6977 (N_6977,N_5886,N_6000);
and U6978 (N_6978,N_5825,N_6355);
xor U6979 (N_6979,N_5932,N_5745);
or U6980 (N_6980,N_5637,N_6385);
xnor U6981 (N_6981,N_5754,N_6193);
nand U6982 (N_6982,N_6164,N_6007);
and U6983 (N_6983,N_6358,N_6184);
nor U6984 (N_6984,N_6121,N_5798);
and U6985 (N_6985,N_6134,N_6173);
xor U6986 (N_6986,N_6181,N_6200);
xor U6987 (N_6987,N_6310,N_5924);
and U6988 (N_6988,N_5879,N_6295);
nand U6989 (N_6989,N_6004,N_5911);
nand U6990 (N_6990,N_6003,N_5738);
nand U6991 (N_6991,N_5681,N_6194);
nor U6992 (N_6992,N_5801,N_5681);
or U6993 (N_6993,N_6064,N_5940);
nor U6994 (N_6994,N_6050,N_6156);
xor U6995 (N_6995,N_6082,N_6255);
nand U6996 (N_6996,N_5776,N_5618);
and U6997 (N_6997,N_5724,N_6343);
and U6998 (N_6998,N_6261,N_6314);
nor U6999 (N_6999,N_5604,N_6311);
xnor U7000 (N_7000,N_6051,N_6318);
or U7001 (N_7001,N_5611,N_6140);
nand U7002 (N_7002,N_5833,N_6399);
nor U7003 (N_7003,N_5850,N_6138);
and U7004 (N_7004,N_5759,N_5893);
xor U7005 (N_7005,N_6394,N_6144);
or U7006 (N_7006,N_5817,N_6155);
or U7007 (N_7007,N_6305,N_5671);
and U7008 (N_7008,N_5982,N_6214);
and U7009 (N_7009,N_6370,N_6210);
or U7010 (N_7010,N_5771,N_5936);
nand U7011 (N_7011,N_5634,N_5661);
nand U7012 (N_7012,N_6176,N_5843);
nor U7013 (N_7013,N_6201,N_6079);
xnor U7014 (N_7014,N_5777,N_5884);
nor U7015 (N_7015,N_6387,N_6203);
or U7016 (N_7016,N_5844,N_5685);
nand U7017 (N_7017,N_5940,N_6116);
nand U7018 (N_7018,N_5822,N_6379);
nor U7019 (N_7019,N_5849,N_5954);
nor U7020 (N_7020,N_6236,N_5726);
and U7021 (N_7021,N_6297,N_6279);
xor U7022 (N_7022,N_5911,N_6142);
or U7023 (N_7023,N_6278,N_5905);
or U7024 (N_7024,N_5754,N_6352);
or U7025 (N_7025,N_5795,N_5995);
or U7026 (N_7026,N_6077,N_5921);
xor U7027 (N_7027,N_6355,N_6035);
nor U7028 (N_7028,N_6248,N_5629);
nor U7029 (N_7029,N_6237,N_6205);
or U7030 (N_7030,N_5940,N_5687);
nor U7031 (N_7031,N_5745,N_5904);
or U7032 (N_7032,N_5886,N_5742);
nor U7033 (N_7033,N_6280,N_6137);
and U7034 (N_7034,N_5914,N_5792);
and U7035 (N_7035,N_6245,N_6009);
nand U7036 (N_7036,N_5671,N_6325);
nor U7037 (N_7037,N_5921,N_6148);
xnor U7038 (N_7038,N_6010,N_5783);
nor U7039 (N_7039,N_5807,N_6060);
xnor U7040 (N_7040,N_6130,N_5837);
and U7041 (N_7041,N_5763,N_6225);
nor U7042 (N_7042,N_6344,N_5991);
nor U7043 (N_7043,N_5833,N_6217);
xnor U7044 (N_7044,N_5926,N_5636);
xor U7045 (N_7045,N_5837,N_5733);
xnor U7046 (N_7046,N_6338,N_5805);
xor U7047 (N_7047,N_6169,N_6063);
nand U7048 (N_7048,N_6149,N_5957);
nand U7049 (N_7049,N_5990,N_6201);
and U7050 (N_7050,N_6191,N_5710);
nand U7051 (N_7051,N_5838,N_6237);
and U7052 (N_7052,N_5647,N_6093);
and U7053 (N_7053,N_5808,N_5811);
nor U7054 (N_7054,N_5926,N_5729);
nor U7055 (N_7055,N_6201,N_5778);
xnor U7056 (N_7056,N_6237,N_6264);
or U7057 (N_7057,N_5646,N_5931);
nand U7058 (N_7058,N_6371,N_5951);
and U7059 (N_7059,N_5925,N_5968);
xor U7060 (N_7060,N_6283,N_5783);
or U7061 (N_7061,N_5612,N_6136);
nand U7062 (N_7062,N_5803,N_6069);
nor U7063 (N_7063,N_6205,N_5912);
nand U7064 (N_7064,N_6105,N_5640);
or U7065 (N_7065,N_6202,N_6144);
xor U7066 (N_7066,N_6355,N_6168);
nor U7067 (N_7067,N_6229,N_6378);
xor U7068 (N_7068,N_6314,N_5832);
xnor U7069 (N_7069,N_5954,N_6215);
nand U7070 (N_7070,N_6016,N_5864);
and U7071 (N_7071,N_5604,N_6262);
nand U7072 (N_7072,N_6138,N_6102);
xor U7073 (N_7073,N_6006,N_6135);
nor U7074 (N_7074,N_5759,N_6233);
xnor U7075 (N_7075,N_6222,N_5692);
or U7076 (N_7076,N_5630,N_5699);
or U7077 (N_7077,N_6029,N_6295);
or U7078 (N_7078,N_6185,N_6167);
nand U7079 (N_7079,N_6372,N_6273);
xor U7080 (N_7080,N_5809,N_5984);
or U7081 (N_7081,N_5870,N_6126);
and U7082 (N_7082,N_5978,N_6020);
nand U7083 (N_7083,N_5935,N_5680);
and U7084 (N_7084,N_6088,N_6317);
nor U7085 (N_7085,N_6021,N_6210);
nand U7086 (N_7086,N_5755,N_5721);
xor U7087 (N_7087,N_5721,N_6217);
nand U7088 (N_7088,N_5849,N_5862);
nor U7089 (N_7089,N_6253,N_5648);
or U7090 (N_7090,N_5959,N_5610);
and U7091 (N_7091,N_6275,N_5670);
nor U7092 (N_7092,N_6156,N_5843);
and U7093 (N_7093,N_6165,N_6222);
xor U7094 (N_7094,N_6388,N_5759);
nand U7095 (N_7095,N_6227,N_6356);
nor U7096 (N_7096,N_6153,N_5756);
nand U7097 (N_7097,N_5694,N_6283);
xnor U7098 (N_7098,N_6278,N_5907);
and U7099 (N_7099,N_5871,N_5654);
xnor U7100 (N_7100,N_5965,N_5801);
and U7101 (N_7101,N_5962,N_6023);
or U7102 (N_7102,N_6029,N_6181);
and U7103 (N_7103,N_6378,N_6213);
xor U7104 (N_7104,N_6141,N_5910);
xnor U7105 (N_7105,N_6125,N_5684);
or U7106 (N_7106,N_6128,N_5680);
xor U7107 (N_7107,N_5809,N_6036);
nor U7108 (N_7108,N_6267,N_6300);
and U7109 (N_7109,N_5947,N_6073);
or U7110 (N_7110,N_6078,N_6211);
or U7111 (N_7111,N_5853,N_5897);
nand U7112 (N_7112,N_5606,N_5669);
and U7113 (N_7113,N_6029,N_6172);
and U7114 (N_7114,N_5903,N_5976);
and U7115 (N_7115,N_5835,N_6290);
nor U7116 (N_7116,N_5843,N_5782);
nor U7117 (N_7117,N_5674,N_5847);
nor U7118 (N_7118,N_6080,N_6177);
and U7119 (N_7119,N_5616,N_6329);
nand U7120 (N_7120,N_6069,N_6398);
xnor U7121 (N_7121,N_6290,N_6286);
and U7122 (N_7122,N_5957,N_6029);
nand U7123 (N_7123,N_6127,N_6213);
nor U7124 (N_7124,N_5873,N_6287);
xnor U7125 (N_7125,N_6187,N_6286);
xnor U7126 (N_7126,N_5794,N_5861);
nand U7127 (N_7127,N_6161,N_6359);
and U7128 (N_7128,N_6355,N_5979);
xnor U7129 (N_7129,N_6199,N_6069);
or U7130 (N_7130,N_6394,N_5881);
or U7131 (N_7131,N_6397,N_6055);
or U7132 (N_7132,N_6025,N_6049);
xnor U7133 (N_7133,N_6168,N_5752);
and U7134 (N_7134,N_6331,N_5847);
xor U7135 (N_7135,N_5963,N_5912);
nand U7136 (N_7136,N_6003,N_5729);
or U7137 (N_7137,N_5640,N_6153);
and U7138 (N_7138,N_5785,N_5903);
or U7139 (N_7139,N_5788,N_5675);
xnor U7140 (N_7140,N_5754,N_5901);
and U7141 (N_7141,N_5724,N_6054);
xnor U7142 (N_7142,N_5845,N_5822);
nand U7143 (N_7143,N_6113,N_6057);
nand U7144 (N_7144,N_6017,N_5849);
nor U7145 (N_7145,N_6209,N_5918);
xnor U7146 (N_7146,N_6029,N_6052);
xnor U7147 (N_7147,N_6065,N_5759);
xor U7148 (N_7148,N_6317,N_6206);
nor U7149 (N_7149,N_6273,N_6293);
nand U7150 (N_7150,N_6343,N_5648);
and U7151 (N_7151,N_6267,N_6035);
nor U7152 (N_7152,N_6307,N_6230);
or U7153 (N_7153,N_6095,N_6126);
xor U7154 (N_7154,N_6083,N_5827);
xor U7155 (N_7155,N_6044,N_6388);
or U7156 (N_7156,N_6234,N_6018);
nand U7157 (N_7157,N_6178,N_6390);
or U7158 (N_7158,N_5659,N_6131);
xor U7159 (N_7159,N_5938,N_6283);
and U7160 (N_7160,N_5900,N_5656);
nor U7161 (N_7161,N_5686,N_5775);
and U7162 (N_7162,N_5901,N_6187);
nor U7163 (N_7163,N_5953,N_5834);
nand U7164 (N_7164,N_5967,N_5612);
or U7165 (N_7165,N_6046,N_5700);
nor U7166 (N_7166,N_6284,N_6114);
and U7167 (N_7167,N_5959,N_6284);
nand U7168 (N_7168,N_5711,N_6330);
xor U7169 (N_7169,N_6144,N_5760);
xor U7170 (N_7170,N_6078,N_6125);
xnor U7171 (N_7171,N_5997,N_5922);
nor U7172 (N_7172,N_6239,N_5864);
nor U7173 (N_7173,N_6018,N_6133);
xnor U7174 (N_7174,N_6120,N_5922);
nand U7175 (N_7175,N_5978,N_6315);
or U7176 (N_7176,N_5872,N_5612);
or U7177 (N_7177,N_6308,N_5652);
xor U7178 (N_7178,N_6031,N_6153);
and U7179 (N_7179,N_6099,N_5859);
and U7180 (N_7180,N_5911,N_5764);
xor U7181 (N_7181,N_6206,N_6066);
nand U7182 (N_7182,N_5759,N_6285);
xnor U7183 (N_7183,N_6273,N_6392);
or U7184 (N_7184,N_5634,N_6399);
nand U7185 (N_7185,N_5928,N_5918);
and U7186 (N_7186,N_6121,N_6137);
xnor U7187 (N_7187,N_5855,N_5926);
or U7188 (N_7188,N_5846,N_6271);
nand U7189 (N_7189,N_6302,N_6128);
nor U7190 (N_7190,N_6301,N_6134);
or U7191 (N_7191,N_5998,N_6019);
nand U7192 (N_7192,N_5769,N_5995);
nor U7193 (N_7193,N_6256,N_6301);
nand U7194 (N_7194,N_6130,N_5696);
and U7195 (N_7195,N_5715,N_6334);
xnor U7196 (N_7196,N_5804,N_6280);
or U7197 (N_7197,N_6209,N_6043);
or U7198 (N_7198,N_5686,N_6395);
and U7199 (N_7199,N_5602,N_6369);
xor U7200 (N_7200,N_6716,N_6543);
nand U7201 (N_7201,N_6905,N_6783);
xor U7202 (N_7202,N_6443,N_6625);
xor U7203 (N_7203,N_6766,N_6489);
and U7204 (N_7204,N_6646,N_6806);
nor U7205 (N_7205,N_7113,N_7094);
nor U7206 (N_7206,N_6997,N_7087);
or U7207 (N_7207,N_6577,N_6845);
nand U7208 (N_7208,N_6485,N_6718);
nand U7209 (N_7209,N_6539,N_6426);
nor U7210 (N_7210,N_7159,N_6505);
xor U7211 (N_7211,N_6675,N_7164);
xnor U7212 (N_7212,N_6690,N_6985);
or U7213 (N_7213,N_7121,N_6546);
xnor U7214 (N_7214,N_6779,N_6514);
xnor U7215 (N_7215,N_6510,N_7178);
and U7216 (N_7216,N_7131,N_6453);
and U7217 (N_7217,N_6672,N_7000);
xnor U7218 (N_7218,N_6778,N_7145);
nor U7219 (N_7219,N_6594,N_7118);
or U7220 (N_7220,N_6775,N_6428);
xor U7221 (N_7221,N_6953,N_6417);
and U7222 (N_7222,N_6970,N_6424);
xnor U7223 (N_7223,N_6527,N_6921);
nand U7224 (N_7224,N_6901,N_7122);
nor U7225 (N_7225,N_7172,N_7003);
or U7226 (N_7226,N_6759,N_6956);
or U7227 (N_7227,N_7038,N_6531);
nand U7228 (N_7228,N_7095,N_7016);
or U7229 (N_7229,N_6658,N_7082);
and U7230 (N_7230,N_6801,N_6883);
nand U7231 (N_7231,N_6873,N_6869);
and U7232 (N_7232,N_6562,N_6425);
or U7233 (N_7233,N_7054,N_6586);
and U7234 (N_7234,N_6526,N_7144);
nand U7235 (N_7235,N_6669,N_6751);
xor U7236 (N_7236,N_7179,N_7032);
nand U7237 (N_7237,N_7052,N_6976);
or U7238 (N_7238,N_7173,N_7149);
nand U7239 (N_7239,N_6939,N_6748);
and U7240 (N_7240,N_6421,N_6573);
xor U7241 (N_7241,N_6731,N_6628);
and U7242 (N_7242,N_6830,N_6816);
xor U7243 (N_7243,N_6856,N_6871);
or U7244 (N_7244,N_6853,N_6467);
nand U7245 (N_7245,N_6535,N_6482);
xnor U7246 (N_7246,N_7056,N_6663);
and U7247 (N_7247,N_6945,N_6671);
xnor U7248 (N_7248,N_7012,N_6805);
nand U7249 (N_7249,N_6844,N_7063);
and U7250 (N_7250,N_7152,N_6497);
nor U7251 (N_7251,N_6875,N_6699);
or U7252 (N_7252,N_6475,N_6578);
and U7253 (N_7253,N_7034,N_6773);
xnor U7254 (N_7254,N_7059,N_6714);
nand U7255 (N_7255,N_6787,N_6710);
or U7256 (N_7256,N_6832,N_6405);
or U7257 (N_7257,N_7141,N_6804);
and U7258 (N_7258,N_6764,N_7187);
or U7259 (N_7259,N_6612,N_6996);
nand U7260 (N_7260,N_6715,N_7027);
nand U7261 (N_7261,N_6544,N_6992);
or U7262 (N_7262,N_6471,N_6430);
nor U7263 (N_7263,N_7018,N_6684);
and U7264 (N_7264,N_6490,N_6944);
and U7265 (N_7265,N_6645,N_6673);
and U7266 (N_7266,N_6767,N_6983);
xor U7267 (N_7267,N_6906,N_6942);
nor U7268 (N_7268,N_6720,N_6643);
or U7269 (N_7269,N_7183,N_6982);
nor U7270 (N_7270,N_6460,N_6558);
nand U7271 (N_7271,N_6441,N_6818);
or U7272 (N_7272,N_6429,N_6717);
or U7273 (N_7273,N_6449,N_6677);
and U7274 (N_7274,N_6642,N_6977);
or U7275 (N_7275,N_6567,N_7073);
nor U7276 (N_7276,N_6528,N_6928);
or U7277 (N_7277,N_7083,N_6974);
nand U7278 (N_7278,N_6632,N_7142);
and U7279 (N_7279,N_6948,N_6436);
xor U7280 (N_7280,N_6515,N_6876);
nor U7281 (N_7281,N_6518,N_6617);
nor U7282 (N_7282,N_6525,N_6738);
and U7283 (N_7283,N_6861,N_6817);
and U7284 (N_7284,N_7108,N_7136);
nand U7285 (N_7285,N_6437,N_6680);
xnor U7286 (N_7286,N_6501,N_6404);
nor U7287 (N_7287,N_7065,N_6620);
nand U7288 (N_7288,N_6704,N_6828);
nor U7289 (N_7289,N_6402,N_7076);
nand U7290 (N_7290,N_6938,N_7162);
and U7291 (N_7291,N_6469,N_7060);
nand U7292 (N_7292,N_6761,N_6534);
nor U7293 (N_7293,N_6739,N_6994);
nand U7294 (N_7294,N_6752,N_6512);
or U7295 (N_7295,N_6866,N_6803);
nor U7296 (N_7296,N_7096,N_6458);
and U7297 (N_7297,N_6819,N_7024);
and U7298 (N_7298,N_6551,N_6403);
or U7299 (N_7299,N_6842,N_6622);
nand U7300 (N_7300,N_7068,N_6457);
or U7301 (N_7301,N_7110,N_7196);
and U7302 (N_7302,N_6568,N_6742);
and U7303 (N_7303,N_6653,N_6712);
xnor U7304 (N_7304,N_6656,N_6674);
and U7305 (N_7305,N_7046,N_6915);
xnor U7306 (N_7306,N_6698,N_6785);
nand U7307 (N_7307,N_6589,N_7086);
and U7308 (N_7308,N_6978,N_6445);
nand U7309 (N_7309,N_7090,N_6413);
nor U7310 (N_7310,N_6434,N_7188);
or U7311 (N_7311,N_6585,N_6823);
or U7312 (N_7312,N_6422,N_6798);
nor U7313 (N_7313,N_6611,N_7045);
nand U7314 (N_7314,N_6652,N_7098);
and U7315 (N_7315,N_6631,N_6637);
or U7316 (N_7316,N_6580,N_6750);
or U7317 (N_7317,N_7181,N_7092);
nand U7318 (N_7318,N_7015,N_7167);
or U7319 (N_7319,N_6760,N_6881);
xor U7320 (N_7320,N_7154,N_6644);
nor U7321 (N_7321,N_6919,N_6981);
or U7322 (N_7322,N_6725,N_6754);
nand U7323 (N_7323,N_6918,N_6857);
xor U7324 (N_7324,N_6797,N_6610);
xnor U7325 (N_7325,N_6519,N_6452);
xor U7326 (N_7326,N_6560,N_7064);
nor U7327 (N_7327,N_7040,N_7158);
or U7328 (N_7328,N_6814,N_6864);
nor U7329 (N_7329,N_6734,N_6912);
nand U7330 (N_7330,N_6630,N_6802);
xor U7331 (N_7331,N_6492,N_6709);
xnor U7332 (N_7332,N_6930,N_6683);
or U7333 (N_7333,N_6486,N_6595);
or U7334 (N_7334,N_7102,N_6681);
or U7335 (N_7335,N_6462,N_6911);
nand U7336 (N_7336,N_6917,N_7171);
xor U7337 (N_7337,N_6986,N_6697);
nor U7338 (N_7338,N_7100,N_6850);
nor U7339 (N_7339,N_6608,N_6524);
nor U7340 (N_7340,N_6520,N_7042);
xor U7341 (N_7341,N_6557,N_6896);
nor U7342 (N_7342,N_6964,N_6762);
xnor U7343 (N_7343,N_6989,N_6827);
or U7344 (N_7344,N_7085,N_6676);
nor U7345 (N_7345,N_7017,N_7127);
xnor U7346 (N_7346,N_6648,N_6572);
or U7347 (N_7347,N_6757,N_6416);
nor U7348 (N_7348,N_6553,N_7191);
nor U7349 (N_7349,N_6592,N_6950);
nor U7350 (N_7350,N_7157,N_6987);
nor U7351 (N_7351,N_7067,N_6897);
xor U7352 (N_7352,N_6926,N_6793);
nand U7353 (N_7353,N_7123,N_6859);
and U7354 (N_7354,N_6809,N_6604);
nor U7355 (N_7355,N_6455,N_6473);
nor U7356 (N_7356,N_6400,N_6640);
nor U7357 (N_7357,N_7057,N_6726);
or U7358 (N_7358,N_6493,N_6420);
xnor U7359 (N_7359,N_6517,N_7013);
nand U7360 (N_7360,N_6679,N_6846);
nand U7361 (N_7361,N_6633,N_7104);
or U7362 (N_7362,N_6599,N_6504);
nor U7363 (N_7363,N_7061,N_6907);
or U7364 (N_7364,N_6598,N_6641);
nor U7365 (N_7365,N_7097,N_6448);
nor U7366 (N_7366,N_6965,N_6872);
nor U7367 (N_7367,N_6729,N_6962);
or U7368 (N_7368,N_6581,N_6583);
or U7369 (N_7369,N_6979,N_6470);
and U7370 (N_7370,N_6721,N_6786);
or U7371 (N_7371,N_7043,N_6914);
and U7372 (N_7372,N_6561,N_6536);
nand U7373 (N_7373,N_6678,N_7020);
nand U7374 (N_7374,N_7036,N_7126);
or U7375 (N_7375,N_7014,N_6909);
or U7376 (N_7376,N_6496,N_7069);
nor U7377 (N_7377,N_7033,N_6870);
and U7378 (N_7378,N_6506,N_6865);
and U7379 (N_7379,N_6913,N_6967);
and U7380 (N_7380,N_6836,N_6899);
and U7381 (N_7381,N_6502,N_6831);
or U7382 (N_7382,N_7037,N_7066);
or U7383 (N_7383,N_7190,N_6481);
nor U7384 (N_7384,N_6508,N_7074);
nor U7385 (N_7385,N_7197,N_7072);
xor U7386 (N_7386,N_7137,N_6666);
nor U7387 (N_7387,N_6664,N_6660);
and U7388 (N_7388,N_6591,N_6858);
nor U7389 (N_7389,N_6924,N_6807);
or U7390 (N_7390,N_6532,N_6874);
xnor U7391 (N_7391,N_6667,N_6614);
nor U7392 (N_7392,N_6559,N_6487);
and U7393 (N_7393,N_6529,N_7019);
and U7394 (N_7394,N_6887,N_7195);
and U7395 (N_7395,N_7089,N_6756);
nand U7396 (N_7396,N_6541,N_6693);
nand U7397 (N_7397,N_6713,N_6796);
xor U7398 (N_7398,N_7161,N_6916);
xor U7399 (N_7399,N_6971,N_6743);
nand U7400 (N_7400,N_6615,N_7175);
and U7401 (N_7401,N_7115,N_6431);
nand U7402 (N_7402,N_7120,N_6900);
xnor U7403 (N_7403,N_6961,N_6507);
nor U7404 (N_7404,N_6877,N_6988);
xor U7405 (N_7405,N_6951,N_7160);
nor U7406 (N_7406,N_6477,N_7135);
or U7407 (N_7407,N_6447,N_6503);
xnor U7408 (N_7408,N_6740,N_6730);
nand U7409 (N_7409,N_7078,N_7101);
and U7410 (N_7410,N_6545,N_7114);
nand U7411 (N_7411,N_6999,N_6638);
or U7412 (N_7412,N_6835,N_7130);
nand U7413 (N_7413,N_6940,N_6694);
nand U7414 (N_7414,N_6542,N_6547);
nor U7415 (N_7415,N_6937,N_6451);
and U7416 (N_7416,N_7049,N_7143);
xnor U7417 (N_7417,N_6483,N_6623);
nor U7418 (N_7418,N_7198,N_6960);
or U7419 (N_7419,N_7129,N_6461);
or U7420 (N_7420,N_7001,N_6929);
xor U7421 (N_7421,N_7047,N_6849);
nor U7422 (N_7422,N_7091,N_6575);
and U7423 (N_7423,N_6571,N_6923);
or U7424 (N_7424,N_6934,N_7151);
or U7425 (N_7425,N_6727,N_6601);
or U7426 (N_7426,N_6891,N_7163);
xnor U7427 (N_7427,N_7008,N_6892);
nand U7428 (N_7428,N_6456,N_7062);
xor U7429 (N_7429,N_6440,N_6843);
or U7430 (N_7430,N_6975,N_6401);
xnor U7431 (N_7431,N_6593,N_6885);
nor U7432 (N_7432,N_6949,N_6834);
nor U7433 (N_7433,N_6587,N_6574);
xnor U7434 (N_7434,N_6657,N_6895);
nor U7435 (N_7435,N_7041,N_6621);
or U7436 (N_7436,N_6626,N_6549);
nor U7437 (N_7437,N_6670,N_6995);
nand U7438 (N_7438,N_7168,N_7147);
xor U7439 (N_7439,N_7165,N_6813);
or U7440 (N_7440,N_6703,N_7155);
and U7441 (N_7441,N_7088,N_6812);
nor U7442 (N_7442,N_6701,N_7093);
nor U7443 (N_7443,N_7006,N_7174);
nor U7444 (N_7444,N_6635,N_6776);
xnor U7445 (N_7445,N_6569,N_6479);
nor U7446 (N_7446,N_6605,N_7119);
nand U7447 (N_7447,N_7176,N_6735);
and U7448 (N_7448,N_6946,N_7011);
xor U7449 (N_7449,N_6533,N_6419);
xnor U7450 (N_7450,N_7186,N_7080);
xor U7451 (N_7451,N_6616,N_6565);
xor U7452 (N_7452,N_6838,N_6476);
xor U7453 (N_7453,N_7146,N_6548);
nor U7454 (N_7454,N_6882,N_6516);
xor U7455 (N_7455,N_6688,N_6736);
nor U7456 (N_7456,N_6732,N_7051);
or U7457 (N_7457,N_6855,N_6499);
xor U7458 (N_7458,N_7193,N_6465);
or U7459 (N_7459,N_7075,N_6815);
xnor U7460 (N_7460,N_6498,N_6687);
xnor U7461 (N_7461,N_7025,N_7081);
nor U7462 (N_7462,N_6662,N_6841);
nand U7463 (N_7463,N_6665,N_6579);
nand U7464 (N_7464,N_6613,N_6491);
or U7465 (N_7465,N_7048,N_6609);
xor U7466 (N_7466,N_6749,N_6737);
and U7467 (N_7467,N_6792,N_6890);
or U7468 (N_7468,N_6603,N_6692);
nand U7469 (N_7469,N_6442,N_6837);
nor U7470 (N_7470,N_6466,N_6878);
nor U7471 (N_7471,N_6418,N_7148);
xor U7472 (N_7472,N_6538,N_7079);
or U7473 (N_7473,N_6863,N_7133);
xnor U7474 (N_7474,N_7004,N_6438);
and U7475 (N_7475,N_7134,N_7031);
nor U7476 (N_7476,N_6600,N_6782);
nand U7477 (N_7477,N_6826,N_6728);
nand U7478 (N_7478,N_7170,N_6522);
xor U7479 (N_7479,N_6523,N_6556);
xnor U7480 (N_7480,N_7166,N_6634);
nor U7481 (N_7481,N_6854,N_7107);
and U7482 (N_7482,N_6597,N_6880);
nand U7483 (N_7483,N_6839,N_6920);
and U7484 (N_7484,N_6468,N_6860);
and U7485 (N_7485,N_6848,N_6500);
or U7486 (N_7486,N_7153,N_6444);
and U7487 (N_7487,N_7002,N_7005);
and U7488 (N_7488,N_7055,N_7194);
and U7489 (N_7489,N_6686,N_6790);
and U7490 (N_7490,N_6765,N_6791);
nand U7491 (N_7491,N_6636,N_6990);
nor U7492 (N_7492,N_7192,N_7124);
and U7493 (N_7493,N_6771,N_6446);
or U7494 (N_7494,N_6947,N_7071);
and U7495 (N_7495,N_6847,N_6898);
and U7496 (N_7496,N_6435,N_6833);
nor U7497 (N_7497,N_6474,N_6570);
xor U7498 (N_7498,N_6800,N_6763);
nand U7499 (N_7499,N_6563,N_7010);
and U7500 (N_7500,N_7180,N_6566);
and U7501 (N_7501,N_7199,N_6596);
nand U7502 (N_7502,N_7139,N_6682);
nand U7503 (N_7503,N_6794,N_6602);
nor U7504 (N_7504,N_6454,N_6941);
nand U7505 (N_7505,N_7169,N_6706);
xnor U7506 (N_7506,N_6409,N_6903);
xnor U7507 (N_7507,N_7030,N_6509);
and U7508 (N_7508,N_6744,N_6550);
nand U7509 (N_7509,N_7105,N_7044);
nor U7510 (N_7510,N_6980,N_6588);
nand U7511 (N_7511,N_7111,N_7021);
nor U7512 (N_7512,N_6707,N_7117);
nand U7513 (N_7513,N_7184,N_6745);
nand U7514 (N_7514,N_6927,N_6627);
and U7515 (N_7515,N_6411,N_6954);
nand U7516 (N_7516,N_6606,N_6450);
nor U7517 (N_7517,N_6552,N_6868);
nand U7518 (N_7518,N_7182,N_6689);
and U7519 (N_7519,N_6691,N_7099);
or U7520 (N_7520,N_6410,N_6655);
or U7521 (N_7521,N_6769,N_6511);
nand U7522 (N_7522,N_6433,N_6576);
xor U7523 (N_7523,N_7009,N_7050);
nand U7524 (N_7524,N_6908,N_6795);
xor U7525 (N_7525,N_6590,N_7026);
or U7526 (N_7526,N_7189,N_7185);
and U7527 (N_7527,N_6943,N_6423);
and U7528 (N_7528,N_6415,N_6733);
nand U7529 (N_7529,N_7156,N_6781);
nand U7530 (N_7530,N_6607,N_6910);
or U7531 (N_7531,N_7070,N_6582);
nor U7532 (N_7532,N_6825,N_6822);
or U7533 (N_7533,N_6893,N_7035);
or U7534 (N_7534,N_6659,N_6955);
xnor U7535 (N_7535,N_6651,N_7084);
and U7536 (N_7536,N_6537,N_6478);
nand U7537 (N_7537,N_6414,N_6821);
nor U7538 (N_7538,N_6700,N_7177);
nand U7539 (N_7539,N_6894,N_6488);
xnor U7540 (N_7540,N_6711,N_6753);
nor U7541 (N_7541,N_6968,N_6747);
or U7542 (N_7542,N_7128,N_7029);
nand U7543 (N_7543,N_6768,N_6746);
nand U7544 (N_7544,N_6777,N_6406);
nor U7545 (N_7545,N_6540,N_6902);
nor U7546 (N_7546,N_6784,N_6884);
nor U7547 (N_7547,N_6494,N_6685);
nand U7548 (N_7548,N_6584,N_6799);
nand U7549 (N_7549,N_7132,N_6879);
or U7550 (N_7550,N_6811,N_6629);
or U7551 (N_7551,N_6820,N_6789);
nand U7552 (N_7552,N_6722,N_6972);
nand U7553 (N_7553,N_6513,N_7023);
xnor U7554 (N_7554,N_6998,N_7053);
nand U7555 (N_7555,N_6649,N_7077);
nand U7556 (N_7556,N_6647,N_6932);
or U7557 (N_7557,N_6772,N_6702);
or U7558 (N_7558,N_6958,N_6464);
and U7559 (N_7559,N_6886,N_6472);
or U7560 (N_7560,N_6936,N_6619);
nor U7561 (N_7561,N_6931,N_7058);
and U7562 (N_7562,N_6695,N_6639);
or U7563 (N_7563,N_6788,N_6933);
xnor U7564 (N_7564,N_6774,N_6724);
nand U7565 (N_7565,N_7125,N_7150);
nand U7566 (N_7566,N_6973,N_7109);
and U7567 (N_7567,N_6952,N_6755);
or U7568 (N_7568,N_6654,N_6829);
xor U7569 (N_7569,N_6484,N_6554);
nor U7570 (N_7570,N_6851,N_6984);
and U7571 (N_7571,N_6564,N_6758);
xor U7572 (N_7572,N_6770,N_6925);
nand U7573 (N_7573,N_6862,N_6624);
nor U7574 (N_7574,N_7039,N_6991);
nor U7575 (N_7575,N_6780,N_6852);
xnor U7576 (N_7576,N_6969,N_6661);
nand U7577 (N_7577,N_7116,N_7112);
or U7578 (N_7578,N_6889,N_6867);
or U7579 (N_7579,N_7007,N_6555);
and U7580 (N_7580,N_6463,N_6705);
nand U7581 (N_7581,N_6935,N_7138);
nand U7582 (N_7582,N_7022,N_6495);
xor U7583 (N_7583,N_6904,N_6723);
nor U7584 (N_7584,N_6810,N_6408);
xor U7585 (N_7585,N_6708,N_6840);
xnor U7586 (N_7586,N_6719,N_6993);
nand U7587 (N_7587,N_6618,N_6966);
nand U7588 (N_7588,N_6741,N_6957);
nand U7589 (N_7589,N_7028,N_6432);
xnor U7590 (N_7590,N_7106,N_6668);
nand U7591 (N_7591,N_6922,N_6439);
xor U7592 (N_7592,N_6480,N_6427);
nand U7593 (N_7593,N_6530,N_6824);
nor U7594 (N_7594,N_6459,N_6650);
or U7595 (N_7595,N_6412,N_7103);
nand U7596 (N_7596,N_6521,N_7140);
xor U7597 (N_7597,N_6959,N_6888);
nand U7598 (N_7598,N_6407,N_6696);
nor U7599 (N_7599,N_6963,N_6808);
or U7600 (N_7600,N_6960,N_6561);
or U7601 (N_7601,N_6743,N_7107);
or U7602 (N_7602,N_7141,N_6404);
xor U7603 (N_7603,N_7114,N_6981);
nand U7604 (N_7604,N_6647,N_6523);
xor U7605 (N_7605,N_6658,N_6961);
and U7606 (N_7606,N_6927,N_6450);
and U7607 (N_7607,N_7177,N_7165);
or U7608 (N_7608,N_7101,N_6563);
and U7609 (N_7609,N_7151,N_6480);
nand U7610 (N_7610,N_6614,N_7000);
nand U7611 (N_7611,N_6577,N_6890);
or U7612 (N_7612,N_6622,N_6553);
or U7613 (N_7613,N_6519,N_6874);
xor U7614 (N_7614,N_6772,N_7016);
nor U7615 (N_7615,N_6476,N_6449);
and U7616 (N_7616,N_6971,N_6744);
nor U7617 (N_7617,N_6738,N_7143);
xnor U7618 (N_7618,N_6950,N_6684);
nor U7619 (N_7619,N_6836,N_7183);
or U7620 (N_7620,N_6941,N_6717);
and U7621 (N_7621,N_6462,N_6808);
or U7622 (N_7622,N_6729,N_6890);
nor U7623 (N_7623,N_6814,N_6723);
or U7624 (N_7624,N_7043,N_7047);
nor U7625 (N_7625,N_6481,N_7151);
or U7626 (N_7626,N_6412,N_7190);
or U7627 (N_7627,N_6960,N_6856);
nor U7628 (N_7628,N_6663,N_6593);
and U7629 (N_7629,N_6791,N_6829);
and U7630 (N_7630,N_6504,N_7088);
or U7631 (N_7631,N_6716,N_6554);
and U7632 (N_7632,N_6417,N_6430);
or U7633 (N_7633,N_6487,N_6860);
and U7634 (N_7634,N_6465,N_6678);
and U7635 (N_7635,N_6525,N_6567);
and U7636 (N_7636,N_6636,N_6475);
xor U7637 (N_7637,N_6848,N_6487);
and U7638 (N_7638,N_6788,N_6968);
xor U7639 (N_7639,N_6472,N_7052);
nand U7640 (N_7640,N_6470,N_6507);
nand U7641 (N_7641,N_6632,N_6791);
and U7642 (N_7642,N_6422,N_6573);
or U7643 (N_7643,N_6630,N_7052);
xor U7644 (N_7644,N_6780,N_6713);
xnor U7645 (N_7645,N_7070,N_7099);
and U7646 (N_7646,N_7171,N_6765);
nand U7647 (N_7647,N_6904,N_6434);
and U7648 (N_7648,N_6624,N_6577);
and U7649 (N_7649,N_6558,N_7010);
and U7650 (N_7650,N_7180,N_6688);
nand U7651 (N_7651,N_6572,N_6969);
nand U7652 (N_7652,N_6622,N_6520);
nor U7653 (N_7653,N_6922,N_6624);
nor U7654 (N_7654,N_6803,N_6474);
and U7655 (N_7655,N_6821,N_7179);
nor U7656 (N_7656,N_6654,N_6808);
and U7657 (N_7657,N_6597,N_6802);
and U7658 (N_7658,N_6486,N_6514);
xor U7659 (N_7659,N_6983,N_6987);
nor U7660 (N_7660,N_6434,N_6492);
nand U7661 (N_7661,N_6475,N_7182);
xor U7662 (N_7662,N_6870,N_7186);
xor U7663 (N_7663,N_6780,N_7172);
or U7664 (N_7664,N_7154,N_6535);
nor U7665 (N_7665,N_6927,N_6501);
or U7666 (N_7666,N_6770,N_6861);
and U7667 (N_7667,N_7078,N_6604);
xnor U7668 (N_7668,N_6611,N_6408);
nor U7669 (N_7669,N_7131,N_6573);
nand U7670 (N_7670,N_7034,N_7189);
xnor U7671 (N_7671,N_6672,N_7081);
nor U7672 (N_7672,N_6468,N_6489);
xnor U7673 (N_7673,N_6566,N_7034);
xnor U7674 (N_7674,N_7088,N_6815);
xor U7675 (N_7675,N_6912,N_7155);
and U7676 (N_7676,N_6491,N_6971);
nand U7677 (N_7677,N_6406,N_7187);
nor U7678 (N_7678,N_6534,N_7082);
nand U7679 (N_7679,N_6842,N_6708);
and U7680 (N_7680,N_6476,N_6785);
nor U7681 (N_7681,N_6496,N_7104);
or U7682 (N_7682,N_6566,N_7135);
or U7683 (N_7683,N_6476,N_6555);
xnor U7684 (N_7684,N_6588,N_7127);
or U7685 (N_7685,N_7192,N_6537);
nor U7686 (N_7686,N_6479,N_6766);
nor U7687 (N_7687,N_7107,N_6642);
nand U7688 (N_7688,N_6943,N_7081);
and U7689 (N_7689,N_6939,N_7097);
nor U7690 (N_7690,N_7025,N_7108);
nor U7691 (N_7691,N_6502,N_7024);
or U7692 (N_7692,N_7110,N_6993);
or U7693 (N_7693,N_6742,N_6656);
or U7694 (N_7694,N_7022,N_6868);
nand U7695 (N_7695,N_6552,N_7073);
nand U7696 (N_7696,N_6438,N_6832);
and U7697 (N_7697,N_6939,N_6881);
nand U7698 (N_7698,N_6974,N_6494);
xor U7699 (N_7699,N_6417,N_7184);
xor U7700 (N_7700,N_7023,N_6931);
nand U7701 (N_7701,N_6761,N_6413);
nand U7702 (N_7702,N_6645,N_7099);
or U7703 (N_7703,N_6874,N_7103);
and U7704 (N_7704,N_6966,N_6840);
and U7705 (N_7705,N_6996,N_6491);
nor U7706 (N_7706,N_6569,N_6862);
xor U7707 (N_7707,N_6591,N_6954);
xnor U7708 (N_7708,N_6423,N_7052);
and U7709 (N_7709,N_6833,N_7118);
nand U7710 (N_7710,N_7091,N_6966);
or U7711 (N_7711,N_6861,N_6871);
and U7712 (N_7712,N_6806,N_7172);
or U7713 (N_7713,N_6432,N_6875);
or U7714 (N_7714,N_6961,N_7090);
nand U7715 (N_7715,N_6915,N_6848);
nor U7716 (N_7716,N_6726,N_6719);
and U7717 (N_7717,N_6517,N_6503);
nor U7718 (N_7718,N_6933,N_7014);
and U7719 (N_7719,N_6727,N_6568);
xor U7720 (N_7720,N_6456,N_6460);
nor U7721 (N_7721,N_6571,N_7183);
xor U7722 (N_7722,N_6908,N_7105);
nor U7723 (N_7723,N_6504,N_6560);
nand U7724 (N_7724,N_6716,N_6953);
nand U7725 (N_7725,N_6951,N_6468);
and U7726 (N_7726,N_6463,N_6513);
nand U7727 (N_7727,N_7078,N_6995);
xnor U7728 (N_7728,N_6531,N_6957);
xnor U7729 (N_7729,N_6943,N_7104);
xor U7730 (N_7730,N_7153,N_6507);
and U7731 (N_7731,N_6679,N_6605);
xor U7732 (N_7732,N_6914,N_6619);
xnor U7733 (N_7733,N_6776,N_6732);
nor U7734 (N_7734,N_6514,N_7004);
xnor U7735 (N_7735,N_6739,N_7195);
xor U7736 (N_7736,N_6408,N_6773);
or U7737 (N_7737,N_7044,N_6922);
xor U7738 (N_7738,N_6951,N_6775);
or U7739 (N_7739,N_7146,N_7077);
and U7740 (N_7740,N_6717,N_7063);
nor U7741 (N_7741,N_7184,N_6818);
nand U7742 (N_7742,N_6972,N_6711);
nor U7743 (N_7743,N_6568,N_6880);
xnor U7744 (N_7744,N_6830,N_6678);
nor U7745 (N_7745,N_7149,N_6921);
nand U7746 (N_7746,N_7120,N_6547);
nand U7747 (N_7747,N_7164,N_7079);
and U7748 (N_7748,N_6440,N_6625);
nand U7749 (N_7749,N_6958,N_6613);
or U7750 (N_7750,N_6915,N_6846);
xnor U7751 (N_7751,N_6522,N_7135);
nor U7752 (N_7752,N_6956,N_7026);
and U7753 (N_7753,N_6472,N_7152);
and U7754 (N_7754,N_6918,N_6735);
or U7755 (N_7755,N_7090,N_6848);
and U7756 (N_7756,N_7138,N_6507);
nor U7757 (N_7757,N_7129,N_6751);
or U7758 (N_7758,N_6609,N_6602);
nor U7759 (N_7759,N_7091,N_6609);
xor U7760 (N_7760,N_6866,N_6477);
and U7761 (N_7761,N_6628,N_6570);
or U7762 (N_7762,N_7176,N_6870);
nor U7763 (N_7763,N_6892,N_6799);
nor U7764 (N_7764,N_7142,N_6444);
nor U7765 (N_7765,N_7164,N_6861);
and U7766 (N_7766,N_6713,N_7124);
and U7767 (N_7767,N_6741,N_6642);
and U7768 (N_7768,N_6656,N_6998);
or U7769 (N_7769,N_6415,N_7012);
and U7770 (N_7770,N_6657,N_6672);
xnor U7771 (N_7771,N_6593,N_6633);
nand U7772 (N_7772,N_7143,N_6496);
xor U7773 (N_7773,N_6690,N_6824);
and U7774 (N_7774,N_6820,N_6443);
and U7775 (N_7775,N_6848,N_6687);
or U7776 (N_7776,N_7090,N_6448);
nor U7777 (N_7777,N_6550,N_7194);
nand U7778 (N_7778,N_6534,N_6448);
and U7779 (N_7779,N_7167,N_6504);
or U7780 (N_7780,N_6594,N_6788);
or U7781 (N_7781,N_6472,N_6602);
and U7782 (N_7782,N_6869,N_6900);
nand U7783 (N_7783,N_6811,N_6644);
xnor U7784 (N_7784,N_6447,N_7082);
and U7785 (N_7785,N_6624,N_6487);
and U7786 (N_7786,N_6707,N_7119);
nor U7787 (N_7787,N_6667,N_6461);
nand U7788 (N_7788,N_6945,N_6504);
or U7789 (N_7789,N_6767,N_6939);
or U7790 (N_7790,N_6764,N_6406);
and U7791 (N_7791,N_7159,N_6532);
xnor U7792 (N_7792,N_7196,N_6757);
nor U7793 (N_7793,N_6447,N_6952);
xor U7794 (N_7794,N_7038,N_6801);
and U7795 (N_7795,N_6781,N_6768);
nand U7796 (N_7796,N_7073,N_6400);
and U7797 (N_7797,N_6414,N_7188);
nand U7798 (N_7798,N_6535,N_7194);
nor U7799 (N_7799,N_7185,N_6614);
nor U7800 (N_7800,N_7130,N_6669);
nand U7801 (N_7801,N_7086,N_6953);
and U7802 (N_7802,N_6420,N_6405);
nor U7803 (N_7803,N_6626,N_7050);
and U7804 (N_7804,N_6800,N_6854);
nand U7805 (N_7805,N_6410,N_6710);
or U7806 (N_7806,N_7128,N_6421);
xor U7807 (N_7807,N_7083,N_6630);
nand U7808 (N_7808,N_6453,N_7092);
nor U7809 (N_7809,N_6488,N_6975);
nand U7810 (N_7810,N_6785,N_7152);
nor U7811 (N_7811,N_7099,N_6983);
and U7812 (N_7812,N_7111,N_6578);
nor U7813 (N_7813,N_6883,N_6987);
and U7814 (N_7814,N_6510,N_6528);
nor U7815 (N_7815,N_7195,N_7084);
nor U7816 (N_7816,N_6550,N_7134);
nor U7817 (N_7817,N_6871,N_7145);
or U7818 (N_7818,N_6472,N_7097);
xnor U7819 (N_7819,N_6791,N_6484);
and U7820 (N_7820,N_6600,N_7154);
xnor U7821 (N_7821,N_6750,N_6827);
nor U7822 (N_7822,N_6603,N_6656);
and U7823 (N_7823,N_7081,N_7162);
nor U7824 (N_7824,N_6890,N_6767);
nor U7825 (N_7825,N_6758,N_6452);
xor U7826 (N_7826,N_6947,N_7133);
and U7827 (N_7827,N_7185,N_6836);
and U7828 (N_7828,N_6955,N_7126);
nand U7829 (N_7829,N_6867,N_6495);
and U7830 (N_7830,N_6877,N_6936);
nand U7831 (N_7831,N_7017,N_6919);
or U7832 (N_7832,N_6969,N_7153);
nand U7833 (N_7833,N_6873,N_6660);
or U7834 (N_7834,N_6745,N_7175);
and U7835 (N_7835,N_6698,N_6700);
nor U7836 (N_7836,N_6826,N_6809);
nor U7837 (N_7837,N_7099,N_7196);
xor U7838 (N_7838,N_6484,N_7189);
xnor U7839 (N_7839,N_6450,N_7009);
and U7840 (N_7840,N_6437,N_7195);
nand U7841 (N_7841,N_6654,N_7024);
and U7842 (N_7842,N_6862,N_7179);
nand U7843 (N_7843,N_6656,N_7106);
and U7844 (N_7844,N_6828,N_6870);
and U7845 (N_7845,N_6859,N_7003);
and U7846 (N_7846,N_6858,N_6966);
nand U7847 (N_7847,N_6551,N_6576);
xor U7848 (N_7848,N_7192,N_6787);
nand U7849 (N_7849,N_6530,N_6897);
nor U7850 (N_7850,N_6638,N_6532);
nand U7851 (N_7851,N_7174,N_6656);
and U7852 (N_7852,N_6933,N_6900);
or U7853 (N_7853,N_6881,N_6428);
xnor U7854 (N_7854,N_6654,N_6667);
nor U7855 (N_7855,N_6577,N_6873);
xor U7856 (N_7856,N_7170,N_6437);
or U7857 (N_7857,N_7088,N_6679);
and U7858 (N_7858,N_7160,N_6715);
nor U7859 (N_7859,N_6825,N_6631);
xnor U7860 (N_7860,N_6479,N_6558);
xor U7861 (N_7861,N_6681,N_7144);
nor U7862 (N_7862,N_6858,N_6735);
nor U7863 (N_7863,N_6892,N_7148);
and U7864 (N_7864,N_7160,N_6714);
xor U7865 (N_7865,N_6765,N_7195);
and U7866 (N_7866,N_7006,N_7079);
nor U7867 (N_7867,N_6674,N_6546);
or U7868 (N_7868,N_6986,N_6991);
xnor U7869 (N_7869,N_7154,N_6638);
or U7870 (N_7870,N_6667,N_7013);
and U7871 (N_7871,N_6482,N_6413);
or U7872 (N_7872,N_6703,N_7077);
xor U7873 (N_7873,N_6401,N_6959);
or U7874 (N_7874,N_7022,N_6547);
or U7875 (N_7875,N_6533,N_6416);
xor U7876 (N_7876,N_6438,N_6922);
or U7877 (N_7877,N_7042,N_6844);
and U7878 (N_7878,N_6498,N_6575);
and U7879 (N_7879,N_6786,N_7068);
and U7880 (N_7880,N_7003,N_6657);
nand U7881 (N_7881,N_6971,N_6563);
xnor U7882 (N_7882,N_6810,N_7077);
and U7883 (N_7883,N_6533,N_6793);
nand U7884 (N_7884,N_6627,N_6765);
xor U7885 (N_7885,N_6527,N_7130);
or U7886 (N_7886,N_6746,N_6454);
nand U7887 (N_7887,N_6580,N_6789);
and U7888 (N_7888,N_6834,N_6846);
or U7889 (N_7889,N_6532,N_6905);
and U7890 (N_7890,N_7169,N_6967);
xnor U7891 (N_7891,N_6517,N_6721);
xnor U7892 (N_7892,N_6712,N_6857);
xor U7893 (N_7893,N_6544,N_6716);
nand U7894 (N_7894,N_6405,N_6838);
xor U7895 (N_7895,N_6627,N_6669);
nor U7896 (N_7896,N_6578,N_6588);
nand U7897 (N_7897,N_6849,N_7193);
nor U7898 (N_7898,N_6824,N_6817);
and U7899 (N_7899,N_7134,N_6930);
xnor U7900 (N_7900,N_6638,N_6621);
and U7901 (N_7901,N_6985,N_6605);
nor U7902 (N_7902,N_6649,N_6406);
xor U7903 (N_7903,N_6582,N_6849);
nand U7904 (N_7904,N_6955,N_6427);
xor U7905 (N_7905,N_6610,N_6444);
and U7906 (N_7906,N_6778,N_6494);
nor U7907 (N_7907,N_7039,N_7162);
nand U7908 (N_7908,N_6855,N_6965);
xnor U7909 (N_7909,N_6996,N_6546);
xnor U7910 (N_7910,N_6678,N_6687);
nor U7911 (N_7911,N_6920,N_6656);
nand U7912 (N_7912,N_7055,N_7119);
nor U7913 (N_7913,N_6478,N_6670);
or U7914 (N_7914,N_6473,N_7045);
nand U7915 (N_7915,N_6585,N_7041);
and U7916 (N_7916,N_7038,N_6890);
nor U7917 (N_7917,N_6662,N_7114);
xor U7918 (N_7918,N_6822,N_6547);
or U7919 (N_7919,N_6676,N_6620);
or U7920 (N_7920,N_6776,N_6999);
xor U7921 (N_7921,N_6441,N_7154);
and U7922 (N_7922,N_6622,N_6800);
nand U7923 (N_7923,N_6732,N_6848);
or U7924 (N_7924,N_6891,N_6803);
nor U7925 (N_7925,N_7110,N_6850);
or U7926 (N_7926,N_6770,N_6622);
and U7927 (N_7927,N_6667,N_7092);
nor U7928 (N_7928,N_7162,N_6831);
nand U7929 (N_7929,N_6708,N_6566);
xnor U7930 (N_7930,N_6809,N_6449);
nor U7931 (N_7931,N_7181,N_7172);
xor U7932 (N_7932,N_6562,N_6938);
and U7933 (N_7933,N_6588,N_6776);
nor U7934 (N_7934,N_6595,N_6411);
nand U7935 (N_7935,N_6931,N_6831);
nor U7936 (N_7936,N_6635,N_6843);
or U7937 (N_7937,N_6701,N_7125);
nand U7938 (N_7938,N_6942,N_6493);
nor U7939 (N_7939,N_6539,N_6447);
xor U7940 (N_7940,N_6492,N_6983);
and U7941 (N_7941,N_6788,N_7175);
nand U7942 (N_7942,N_6473,N_6457);
nor U7943 (N_7943,N_6444,N_6609);
nand U7944 (N_7944,N_6971,N_6965);
xor U7945 (N_7945,N_6993,N_6770);
xor U7946 (N_7946,N_6953,N_7052);
nor U7947 (N_7947,N_6481,N_6603);
and U7948 (N_7948,N_6698,N_7135);
xor U7949 (N_7949,N_6784,N_6573);
or U7950 (N_7950,N_6557,N_6892);
nor U7951 (N_7951,N_7187,N_6640);
xor U7952 (N_7952,N_6619,N_6441);
or U7953 (N_7953,N_6664,N_6454);
or U7954 (N_7954,N_6881,N_6572);
nand U7955 (N_7955,N_6753,N_6526);
nand U7956 (N_7956,N_7008,N_6434);
nand U7957 (N_7957,N_6908,N_7177);
xnor U7958 (N_7958,N_6564,N_6819);
xnor U7959 (N_7959,N_6940,N_6409);
nand U7960 (N_7960,N_6986,N_6510);
and U7961 (N_7961,N_6653,N_6478);
nor U7962 (N_7962,N_6811,N_7054);
and U7963 (N_7963,N_6513,N_6707);
and U7964 (N_7964,N_7182,N_6512);
or U7965 (N_7965,N_7035,N_6823);
and U7966 (N_7966,N_6475,N_6446);
xor U7967 (N_7967,N_6735,N_6511);
and U7968 (N_7968,N_6524,N_6807);
or U7969 (N_7969,N_7089,N_6519);
nor U7970 (N_7970,N_7181,N_7116);
or U7971 (N_7971,N_6446,N_6610);
xnor U7972 (N_7972,N_6589,N_6747);
or U7973 (N_7973,N_6608,N_6884);
nand U7974 (N_7974,N_7060,N_7088);
xnor U7975 (N_7975,N_6755,N_6635);
xnor U7976 (N_7976,N_6761,N_6478);
nor U7977 (N_7977,N_7156,N_6637);
xor U7978 (N_7978,N_6896,N_7121);
nor U7979 (N_7979,N_6824,N_7058);
nor U7980 (N_7980,N_6860,N_6608);
nand U7981 (N_7981,N_6929,N_6727);
nor U7982 (N_7982,N_6414,N_7092);
or U7983 (N_7983,N_7068,N_6909);
and U7984 (N_7984,N_6711,N_7151);
or U7985 (N_7985,N_6795,N_7179);
and U7986 (N_7986,N_6496,N_6417);
and U7987 (N_7987,N_7004,N_6492);
nand U7988 (N_7988,N_6697,N_7065);
nor U7989 (N_7989,N_6639,N_6933);
xnor U7990 (N_7990,N_6541,N_6950);
and U7991 (N_7991,N_7130,N_6497);
xor U7992 (N_7992,N_6480,N_6732);
xnor U7993 (N_7993,N_6404,N_7056);
or U7994 (N_7994,N_6663,N_6967);
and U7995 (N_7995,N_7190,N_7122);
nand U7996 (N_7996,N_7147,N_7119);
xor U7997 (N_7997,N_6595,N_6454);
and U7998 (N_7998,N_6970,N_6445);
nor U7999 (N_7999,N_7004,N_7135);
nor U8000 (N_8000,N_7525,N_7542);
nand U8001 (N_8001,N_7565,N_7363);
or U8002 (N_8002,N_7898,N_7513);
nor U8003 (N_8003,N_7949,N_7215);
or U8004 (N_8004,N_7350,N_7429);
nand U8005 (N_8005,N_7318,N_7720);
nand U8006 (N_8006,N_7664,N_7531);
xor U8007 (N_8007,N_7374,N_7909);
nor U8008 (N_8008,N_7221,N_7815);
nand U8009 (N_8009,N_7506,N_7395);
or U8010 (N_8010,N_7871,N_7792);
nand U8011 (N_8011,N_7292,N_7763);
nand U8012 (N_8012,N_7878,N_7389);
xor U8013 (N_8013,N_7281,N_7454);
or U8014 (N_8014,N_7800,N_7366);
or U8015 (N_8015,N_7876,N_7385);
and U8016 (N_8016,N_7545,N_7834);
nor U8017 (N_8017,N_7300,N_7770);
and U8018 (N_8018,N_7904,N_7338);
and U8019 (N_8019,N_7952,N_7560);
nor U8020 (N_8020,N_7201,N_7356);
nor U8021 (N_8021,N_7825,N_7370);
or U8022 (N_8022,N_7690,N_7265);
xnor U8023 (N_8023,N_7582,N_7775);
xor U8024 (N_8024,N_7637,N_7751);
nor U8025 (N_8025,N_7620,N_7269);
and U8026 (N_8026,N_7453,N_7767);
xnor U8027 (N_8027,N_7512,N_7974);
and U8028 (N_8028,N_7655,N_7990);
or U8029 (N_8029,N_7963,N_7859);
nor U8030 (N_8030,N_7968,N_7762);
xor U8031 (N_8031,N_7564,N_7252);
and U8032 (N_8032,N_7344,N_7745);
nand U8033 (N_8033,N_7554,N_7862);
xor U8034 (N_8034,N_7803,N_7346);
xor U8035 (N_8035,N_7786,N_7724);
xor U8036 (N_8036,N_7636,N_7750);
or U8037 (N_8037,N_7302,N_7879);
and U8038 (N_8038,N_7896,N_7460);
nor U8039 (N_8039,N_7839,N_7601);
nor U8040 (N_8040,N_7541,N_7520);
xor U8041 (N_8041,N_7722,N_7309);
or U8042 (N_8042,N_7758,N_7623);
nand U8043 (N_8043,N_7549,N_7508);
or U8044 (N_8044,N_7503,N_7624);
and U8045 (N_8045,N_7980,N_7977);
xnor U8046 (N_8046,N_7659,N_7957);
nor U8047 (N_8047,N_7702,N_7440);
nand U8048 (N_8048,N_7261,N_7217);
or U8049 (N_8049,N_7243,N_7646);
nor U8050 (N_8050,N_7518,N_7324);
xor U8051 (N_8051,N_7218,N_7673);
nor U8052 (N_8052,N_7475,N_7998);
xnor U8053 (N_8053,N_7547,N_7442);
xnor U8054 (N_8054,N_7894,N_7308);
nor U8055 (N_8055,N_7956,N_7789);
and U8056 (N_8056,N_7778,N_7517);
xor U8057 (N_8057,N_7443,N_7293);
xnor U8058 (N_8058,N_7357,N_7915);
nand U8059 (N_8059,N_7887,N_7959);
or U8060 (N_8060,N_7418,N_7811);
xnor U8061 (N_8061,N_7556,N_7406);
nor U8062 (N_8062,N_7474,N_7604);
xnor U8063 (N_8063,N_7480,N_7206);
nor U8064 (N_8064,N_7929,N_7703);
and U8065 (N_8065,N_7658,N_7790);
nand U8066 (N_8066,N_7203,N_7467);
xor U8067 (N_8067,N_7596,N_7849);
and U8068 (N_8068,N_7727,N_7723);
or U8069 (N_8069,N_7852,N_7299);
nor U8070 (N_8070,N_7408,N_7526);
nand U8071 (N_8071,N_7643,N_7725);
nand U8072 (N_8072,N_7536,N_7411);
or U8073 (N_8073,N_7400,N_7414);
and U8074 (N_8074,N_7897,N_7765);
and U8075 (N_8075,N_7251,N_7900);
and U8076 (N_8076,N_7472,N_7476);
or U8077 (N_8077,N_7548,N_7449);
or U8078 (N_8078,N_7899,N_7239);
nor U8079 (N_8079,N_7779,N_7228);
nand U8080 (N_8080,N_7749,N_7985);
nand U8081 (N_8081,N_7225,N_7884);
or U8082 (N_8082,N_7841,N_7569);
or U8083 (N_8083,N_7505,N_7917);
nor U8084 (N_8084,N_7836,N_7832);
xnor U8085 (N_8085,N_7907,N_7247);
nand U8086 (N_8086,N_7425,N_7736);
or U8087 (N_8087,N_7540,N_7424);
nor U8088 (N_8088,N_7921,N_7578);
xnor U8089 (N_8089,N_7369,N_7873);
or U8090 (N_8090,N_7470,N_7784);
and U8091 (N_8091,N_7423,N_7700);
or U8092 (N_8092,N_7532,N_7240);
nand U8093 (N_8093,N_7204,N_7679);
nor U8094 (N_8094,N_7372,N_7671);
nor U8095 (N_8095,N_7960,N_7431);
and U8096 (N_8096,N_7818,N_7335);
and U8097 (N_8097,N_7823,N_7375);
xor U8098 (N_8098,N_7647,N_7202);
xor U8099 (N_8099,N_7529,N_7530);
and U8100 (N_8100,N_7735,N_7412);
nand U8101 (N_8101,N_7844,N_7500);
xor U8102 (N_8102,N_7326,N_7728);
or U8103 (N_8103,N_7696,N_7714);
nor U8104 (N_8104,N_7405,N_7427);
and U8105 (N_8105,N_7208,N_7981);
xnor U8106 (N_8106,N_7359,N_7437);
nand U8107 (N_8107,N_7978,N_7616);
xnor U8108 (N_8108,N_7448,N_7331);
or U8109 (N_8109,N_7478,N_7550);
xnor U8110 (N_8110,N_7742,N_7289);
nor U8111 (N_8111,N_7450,N_7524);
or U8112 (N_8112,N_7591,N_7386);
nand U8113 (N_8113,N_7488,N_7691);
xor U8114 (N_8114,N_7877,N_7991);
and U8115 (N_8115,N_7627,N_7222);
and U8116 (N_8116,N_7730,N_7861);
or U8117 (N_8117,N_7559,N_7330);
nand U8118 (N_8118,N_7794,N_7523);
and U8119 (N_8119,N_7989,N_7870);
xnor U8120 (N_8120,N_7705,N_7321);
nand U8121 (N_8121,N_7317,N_7988);
or U8122 (N_8122,N_7787,N_7707);
and U8123 (N_8123,N_7603,N_7504);
xor U8124 (N_8124,N_7680,N_7595);
xnor U8125 (N_8125,N_7419,N_7973);
and U8126 (N_8126,N_7864,N_7965);
xnor U8127 (N_8127,N_7902,N_7972);
or U8128 (N_8128,N_7848,N_7394);
xnor U8129 (N_8129,N_7975,N_7910);
and U8130 (N_8130,N_7342,N_7842);
or U8131 (N_8131,N_7966,N_7721);
and U8132 (N_8132,N_7320,N_7782);
nor U8133 (N_8133,N_7746,N_7783);
or U8134 (N_8134,N_7580,N_7439);
or U8135 (N_8135,N_7498,N_7490);
and U8136 (N_8136,N_7235,N_7905);
nor U8137 (N_8137,N_7641,N_7349);
and U8138 (N_8138,N_7764,N_7938);
xnor U8139 (N_8139,N_7415,N_7539);
nand U8140 (N_8140,N_7417,N_7717);
and U8141 (N_8141,N_7961,N_7734);
nand U8142 (N_8142,N_7589,N_7355);
or U8143 (N_8143,N_7666,N_7364);
and U8144 (N_8144,N_7553,N_7820);
nand U8145 (N_8145,N_7420,N_7574);
or U8146 (N_8146,N_7378,N_7607);
nor U8147 (N_8147,N_7285,N_7934);
nor U8148 (N_8148,N_7477,N_7947);
nor U8149 (N_8149,N_7813,N_7528);
or U8150 (N_8150,N_7983,N_7708);
or U8151 (N_8151,N_7583,N_7796);
xnor U8152 (N_8152,N_7986,N_7935);
nand U8153 (N_8153,N_7692,N_7371);
xnor U8154 (N_8154,N_7447,N_7821);
xor U8155 (N_8155,N_7737,N_7812);
and U8156 (N_8156,N_7927,N_7459);
and U8157 (N_8157,N_7808,N_7592);
nor U8158 (N_8158,N_7576,N_7916);
xnor U8159 (N_8159,N_7209,N_7482);
xnor U8160 (N_8160,N_7455,N_7367);
and U8161 (N_8161,N_7587,N_7280);
and U8162 (N_8162,N_7855,N_7451);
and U8163 (N_8163,N_7584,N_7628);
and U8164 (N_8164,N_7510,N_7826);
nand U8165 (N_8165,N_7889,N_7801);
nor U8166 (N_8166,N_7464,N_7639);
nor U8167 (N_8167,N_7997,N_7594);
nand U8168 (N_8168,N_7245,N_7713);
and U8169 (N_8169,N_7341,N_7581);
nand U8170 (N_8170,N_7885,N_7469);
xor U8171 (N_8171,N_7617,N_7630);
nor U8172 (N_8172,N_7492,N_7279);
xnor U8173 (N_8173,N_7755,N_7631);
nand U8174 (N_8174,N_7267,N_7211);
nor U8175 (N_8175,N_7283,N_7828);
nor U8176 (N_8176,N_7567,N_7964);
nor U8177 (N_8177,N_7872,N_7835);
xnor U8178 (N_8178,N_7901,N_7798);
nor U8179 (N_8179,N_7468,N_7648);
xnor U8180 (N_8180,N_7677,N_7555);
and U8181 (N_8181,N_7345,N_7298);
nor U8182 (N_8182,N_7312,N_7716);
or U8183 (N_8183,N_7296,N_7919);
nor U8184 (N_8184,N_7231,N_7301);
xnor U8185 (N_8185,N_7230,N_7912);
nor U8186 (N_8186,N_7621,N_7942);
nand U8187 (N_8187,N_7670,N_7774);
and U8188 (N_8188,N_7939,N_7537);
nor U8189 (N_8189,N_7358,N_7996);
xor U8190 (N_8190,N_7388,N_7577);
nand U8191 (N_8191,N_7271,N_7914);
or U8192 (N_8192,N_7752,N_7333);
and U8193 (N_8193,N_7307,N_7824);
and U8194 (N_8194,N_7260,N_7436);
or U8195 (N_8195,N_7936,N_7650);
and U8196 (N_8196,N_7600,N_7651);
xnor U8197 (N_8197,N_7911,N_7390);
or U8198 (N_8198,N_7212,N_7791);
or U8199 (N_8199,N_7753,N_7501);
nor U8200 (N_8200,N_7822,N_7391);
and U8201 (N_8201,N_7586,N_7760);
nor U8202 (N_8202,N_7473,N_7274);
nor U8203 (N_8203,N_7928,N_7622);
or U8204 (N_8204,N_7984,N_7954);
xor U8205 (N_8205,N_7214,N_7731);
nand U8206 (N_8206,N_7483,N_7652);
xor U8207 (N_8207,N_7257,N_7625);
nor U8208 (N_8208,N_7270,N_7327);
nor U8209 (N_8209,N_7502,N_7404);
and U8210 (N_8210,N_7777,N_7995);
and U8211 (N_8211,N_7507,N_7881);
nand U8212 (N_8212,N_7924,N_7999);
nand U8213 (N_8213,N_7272,N_7310);
or U8214 (N_8214,N_7494,N_7612);
nor U8215 (N_8215,N_7688,N_7227);
nor U8216 (N_8216,N_7880,N_7795);
and U8217 (N_8217,N_7387,N_7804);
or U8218 (N_8218,N_7867,N_7890);
or U8219 (N_8219,N_7726,N_7223);
nand U8220 (N_8220,N_7340,N_7552);
nor U8221 (N_8221,N_7829,N_7739);
nor U8222 (N_8222,N_7718,N_7645);
nor U8223 (N_8223,N_7810,N_7273);
xnor U8224 (N_8224,N_7487,N_7433);
and U8225 (N_8225,N_7337,N_7336);
or U8226 (N_8226,N_7351,N_7781);
and U8227 (N_8227,N_7663,N_7416);
and U8228 (N_8228,N_7656,N_7869);
or U8229 (N_8229,N_7759,N_7465);
xnor U8230 (N_8230,N_7353,N_7323);
xor U8231 (N_8231,N_7496,N_7426);
nor U8232 (N_8232,N_7712,N_7729);
or U8233 (N_8233,N_7275,N_7698);
or U8234 (N_8234,N_7383,N_7410);
nor U8235 (N_8235,N_7264,N_7892);
xnor U8236 (N_8236,N_7397,N_7672);
or U8237 (N_8237,N_7238,N_7614);
and U8238 (N_8238,N_7551,N_7462);
xnor U8239 (N_8239,N_7236,N_7955);
nand U8240 (N_8240,N_7250,N_7495);
nor U8241 (N_8241,N_7807,N_7805);
nor U8242 (N_8242,N_7207,N_7930);
xnor U8243 (N_8243,N_7543,N_7237);
nor U8244 (N_8244,N_7684,N_7521);
nor U8245 (N_8245,N_7295,N_7865);
nor U8246 (N_8246,N_7976,N_7562);
or U8247 (N_8247,N_7354,N_7967);
or U8248 (N_8248,N_7969,N_7568);
and U8249 (N_8249,N_7254,N_7733);
nand U8250 (N_8250,N_7785,N_7635);
or U8251 (N_8251,N_7768,N_7944);
xor U8252 (N_8252,N_7328,N_7398);
xnor U8253 (N_8253,N_7315,N_7945);
nor U8254 (N_8254,N_7857,N_7377);
nor U8255 (N_8255,N_7788,N_7304);
nand U8256 (N_8256,N_7579,N_7799);
nor U8257 (N_8257,N_7253,N_7686);
or U8258 (N_8258,N_7706,N_7806);
and U8259 (N_8259,N_7875,N_7428);
and U8260 (N_8260,N_7863,N_7719);
nand U8261 (N_8261,N_7851,N_7435);
nand U8262 (N_8262,N_7926,N_7906);
or U8263 (N_8263,N_7937,N_7773);
xor U8264 (N_8264,N_7489,N_7516);
nor U8265 (N_8265,N_7305,N_7987);
and U8266 (N_8266,N_7886,N_7598);
xnor U8267 (N_8267,N_7827,N_7514);
xnor U8268 (N_8268,N_7258,N_7802);
xnor U8269 (N_8269,N_7544,N_7874);
or U8270 (N_8270,N_7461,N_7701);
or U8271 (N_8271,N_7845,N_7497);
xnor U8272 (N_8272,N_7840,N_7590);
xnor U8273 (N_8273,N_7399,N_7360);
nand U8274 (N_8274,N_7837,N_7754);
nor U8275 (N_8275,N_7563,N_7535);
nor U8276 (N_8276,N_7558,N_7626);
nand U8277 (N_8277,N_7678,N_7866);
and U8278 (N_8278,N_7287,N_7608);
or U8279 (N_8279,N_7226,N_7365);
nand U8280 (N_8280,N_7605,N_7421);
nor U8281 (N_8281,N_7519,N_7284);
nor U8282 (N_8282,N_7546,N_7882);
or U8283 (N_8283,N_7710,N_7573);
nand U8284 (N_8284,N_7971,N_7444);
nor U8285 (N_8285,N_7854,N_7329);
and U8286 (N_8286,N_7962,N_7611);
xor U8287 (N_8287,N_7352,N_7715);
and U8288 (N_8288,N_7649,N_7756);
and U8289 (N_8289,N_7970,N_7948);
nand U8290 (N_8290,N_7695,N_7681);
or U8291 (N_8291,N_7402,N_7610);
or U8292 (N_8292,N_7255,N_7950);
nand U8293 (N_8293,N_7561,N_7943);
xnor U8294 (N_8294,N_7286,N_7527);
or U8295 (N_8295,N_7891,N_7241);
or U8296 (N_8296,N_7657,N_7566);
xor U8297 (N_8297,N_7632,N_7994);
or U8298 (N_8298,N_7619,N_7456);
xor U8299 (N_8299,N_7484,N_7893);
nor U8300 (N_8300,N_7668,N_7888);
nand U8301 (N_8301,N_7757,N_7282);
nand U8302 (N_8302,N_7362,N_7660);
xor U8303 (N_8303,N_7422,N_7618);
xor U8304 (N_8304,N_7856,N_7325);
and U8305 (N_8305,N_7316,N_7446);
and U8306 (N_8306,N_7599,N_7846);
nand U8307 (N_8307,N_7220,N_7382);
nand U8308 (N_8308,N_7709,N_7339);
or U8309 (N_8309,N_7693,N_7920);
xor U8310 (N_8310,N_7593,N_7819);
or U8311 (N_8311,N_7993,N_7361);
nand U8312 (N_8312,N_7430,N_7638);
nor U8313 (N_8313,N_7923,N_7653);
nor U8314 (N_8314,N_7268,N_7740);
nor U8315 (N_8315,N_7306,N_7908);
nand U8316 (N_8316,N_7667,N_7953);
and U8317 (N_8317,N_7931,N_7457);
and U8318 (N_8318,N_7689,N_7249);
nor U8319 (N_8319,N_7588,N_7373);
nor U8320 (N_8320,N_7933,N_7633);
nor U8321 (N_8321,N_7244,N_7452);
or U8322 (N_8322,N_7232,N_7748);
xnor U8323 (N_8323,N_7246,N_7368);
nand U8324 (N_8324,N_7259,N_7683);
or U8325 (N_8325,N_7613,N_7860);
or U8326 (N_8326,N_7445,N_7946);
xor U8327 (N_8327,N_7343,N_7615);
or U8328 (N_8328,N_7311,N_7982);
or U8329 (N_8329,N_7675,N_7533);
nand U8330 (N_8330,N_7511,N_7644);
and U8331 (N_8331,N_7485,N_7932);
nor U8332 (N_8332,N_7704,N_7229);
or U8333 (N_8333,N_7850,N_7216);
nand U8334 (N_8334,N_7674,N_7409);
xnor U8335 (N_8335,N_7522,N_7200);
or U8336 (N_8336,N_7654,N_7413);
nor U8337 (N_8337,N_7471,N_7780);
nor U8338 (N_8338,N_7817,N_7438);
xor U8339 (N_8339,N_7699,N_7233);
xnor U8340 (N_8340,N_7381,N_7458);
and U8341 (N_8341,N_7687,N_7662);
nand U8342 (N_8342,N_7407,N_7772);
xor U8343 (N_8343,N_7843,N_7738);
nand U8344 (N_8344,N_7481,N_7314);
nor U8345 (N_8345,N_7868,N_7682);
nor U8346 (N_8346,N_7294,N_7515);
or U8347 (N_8347,N_7379,N_7297);
and U8348 (N_8348,N_7711,N_7732);
nor U8349 (N_8349,N_7769,N_7833);
xor U8350 (N_8350,N_7277,N_7266);
xor U8351 (N_8351,N_7831,N_7205);
nand U8352 (N_8352,N_7744,N_7883);
or U8353 (N_8353,N_7847,N_7376);
nand U8354 (N_8354,N_7463,N_7219);
or U8355 (N_8355,N_7838,N_7224);
nor U8356 (N_8356,N_7771,N_7303);
xor U8357 (N_8357,N_7992,N_7441);
and U8358 (N_8358,N_7491,N_7640);
or U8359 (N_8359,N_7776,N_7384);
nor U8360 (N_8360,N_7816,N_7741);
nand U8361 (N_8361,N_7572,N_7597);
nand U8362 (N_8362,N_7697,N_7669);
and U8363 (N_8363,N_7922,N_7348);
or U8364 (N_8364,N_7256,N_7747);
and U8365 (N_8365,N_7557,N_7858);
or U8366 (N_8366,N_7380,N_7940);
or U8367 (N_8367,N_7918,N_7466);
and U8368 (N_8368,N_7629,N_7634);
and U8369 (N_8369,N_7234,N_7392);
xnor U8370 (N_8370,N_7432,N_7575);
and U8371 (N_8371,N_7814,N_7534);
and U8372 (N_8372,N_7661,N_7322);
nand U8373 (N_8373,N_7913,N_7694);
xnor U8374 (N_8374,N_7895,N_7665);
nand U8375 (N_8375,N_7334,N_7830);
nor U8376 (N_8376,N_7210,N_7213);
xor U8377 (N_8377,N_7979,N_7403);
nor U8378 (N_8378,N_7606,N_7676);
or U8379 (N_8379,N_7493,N_7290);
xnor U8380 (N_8380,N_7262,N_7538);
and U8381 (N_8381,N_7479,N_7347);
or U8382 (N_8382,N_7642,N_7958);
nand U8383 (N_8383,N_7499,N_7685);
and U8384 (N_8384,N_7396,N_7288);
nor U8385 (N_8385,N_7486,N_7570);
xor U8386 (N_8386,N_7585,N_7809);
or U8387 (N_8387,N_7263,N_7925);
and U8388 (N_8388,N_7797,N_7609);
xnor U8389 (N_8389,N_7766,N_7248);
nor U8390 (N_8390,N_7276,N_7761);
and U8391 (N_8391,N_7903,N_7509);
or U8392 (N_8392,N_7571,N_7793);
nor U8393 (N_8393,N_7434,N_7602);
and U8394 (N_8394,N_7853,N_7319);
or U8395 (N_8395,N_7278,N_7951);
xnor U8396 (N_8396,N_7313,N_7743);
or U8397 (N_8397,N_7242,N_7401);
and U8398 (N_8398,N_7291,N_7941);
nand U8399 (N_8399,N_7393,N_7332);
or U8400 (N_8400,N_7605,N_7997);
or U8401 (N_8401,N_7649,N_7847);
nor U8402 (N_8402,N_7511,N_7364);
or U8403 (N_8403,N_7992,N_7835);
nor U8404 (N_8404,N_7710,N_7748);
nor U8405 (N_8405,N_7941,N_7240);
or U8406 (N_8406,N_7943,N_7764);
xnor U8407 (N_8407,N_7408,N_7531);
nor U8408 (N_8408,N_7441,N_7974);
xor U8409 (N_8409,N_7454,N_7982);
xor U8410 (N_8410,N_7516,N_7977);
or U8411 (N_8411,N_7643,N_7388);
xor U8412 (N_8412,N_7559,N_7834);
nand U8413 (N_8413,N_7505,N_7859);
and U8414 (N_8414,N_7263,N_7991);
xor U8415 (N_8415,N_7683,N_7598);
and U8416 (N_8416,N_7531,N_7303);
or U8417 (N_8417,N_7723,N_7458);
or U8418 (N_8418,N_7626,N_7201);
nand U8419 (N_8419,N_7658,N_7716);
nor U8420 (N_8420,N_7984,N_7627);
nand U8421 (N_8421,N_7405,N_7942);
or U8422 (N_8422,N_7243,N_7665);
nor U8423 (N_8423,N_7651,N_7971);
nand U8424 (N_8424,N_7759,N_7637);
nand U8425 (N_8425,N_7500,N_7830);
nand U8426 (N_8426,N_7938,N_7702);
and U8427 (N_8427,N_7838,N_7395);
nor U8428 (N_8428,N_7443,N_7789);
xnor U8429 (N_8429,N_7377,N_7489);
xnor U8430 (N_8430,N_7222,N_7290);
nor U8431 (N_8431,N_7894,N_7727);
nand U8432 (N_8432,N_7857,N_7950);
nor U8433 (N_8433,N_7215,N_7575);
xor U8434 (N_8434,N_7621,N_7474);
or U8435 (N_8435,N_7245,N_7526);
nand U8436 (N_8436,N_7577,N_7857);
nor U8437 (N_8437,N_7383,N_7683);
xor U8438 (N_8438,N_7654,N_7670);
nor U8439 (N_8439,N_7661,N_7478);
nand U8440 (N_8440,N_7765,N_7676);
or U8441 (N_8441,N_7878,N_7812);
xnor U8442 (N_8442,N_7577,N_7837);
nor U8443 (N_8443,N_7752,N_7649);
and U8444 (N_8444,N_7576,N_7563);
nor U8445 (N_8445,N_7518,N_7959);
nand U8446 (N_8446,N_7783,N_7865);
nand U8447 (N_8447,N_7282,N_7325);
xnor U8448 (N_8448,N_7693,N_7285);
xnor U8449 (N_8449,N_7549,N_7784);
or U8450 (N_8450,N_7692,N_7231);
nor U8451 (N_8451,N_7636,N_7335);
xnor U8452 (N_8452,N_7627,N_7630);
or U8453 (N_8453,N_7876,N_7406);
xor U8454 (N_8454,N_7488,N_7637);
or U8455 (N_8455,N_7556,N_7614);
or U8456 (N_8456,N_7584,N_7413);
nor U8457 (N_8457,N_7625,N_7925);
nand U8458 (N_8458,N_7830,N_7397);
and U8459 (N_8459,N_7261,N_7320);
or U8460 (N_8460,N_7816,N_7807);
nand U8461 (N_8461,N_7616,N_7664);
nand U8462 (N_8462,N_7924,N_7454);
xor U8463 (N_8463,N_7939,N_7927);
and U8464 (N_8464,N_7989,N_7625);
nand U8465 (N_8465,N_7635,N_7505);
or U8466 (N_8466,N_7579,N_7550);
and U8467 (N_8467,N_7640,N_7853);
xnor U8468 (N_8468,N_7756,N_7850);
nand U8469 (N_8469,N_7710,N_7253);
or U8470 (N_8470,N_7722,N_7282);
and U8471 (N_8471,N_7901,N_7567);
or U8472 (N_8472,N_7587,N_7596);
xor U8473 (N_8473,N_7506,N_7727);
xnor U8474 (N_8474,N_7327,N_7307);
and U8475 (N_8475,N_7665,N_7825);
nand U8476 (N_8476,N_7430,N_7431);
and U8477 (N_8477,N_7299,N_7820);
xnor U8478 (N_8478,N_7280,N_7940);
and U8479 (N_8479,N_7216,N_7241);
nand U8480 (N_8480,N_7212,N_7202);
nor U8481 (N_8481,N_7450,N_7733);
or U8482 (N_8482,N_7615,N_7654);
xnor U8483 (N_8483,N_7768,N_7398);
and U8484 (N_8484,N_7372,N_7455);
xnor U8485 (N_8485,N_7850,N_7468);
nand U8486 (N_8486,N_7885,N_7474);
and U8487 (N_8487,N_7345,N_7676);
or U8488 (N_8488,N_7579,N_7415);
nand U8489 (N_8489,N_7565,N_7304);
xor U8490 (N_8490,N_7399,N_7811);
nor U8491 (N_8491,N_7310,N_7720);
xnor U8492 (N_8492,N_7203,N_7942);
nand U8493 (N_8493,N_7339,N_7837);
xor U8494 (N_8494,N_7817,N_7274);
nand U8495 (N_8495,N_7378,N_7472);
nand U8496 (N_8496,N_7461,N_7837);
nor U8497 (N_8497,N_7528,N_7769);
xor U8498 (N_8498,N_7288,N_7309);
nand U8499 (N_8499,N_7321,N_7206);
xor U8500 (N_8500,N_7657,N_7516);
and U8501 (N_8501,N_7786,N_7481);
and U8502 (N_8502,N_7898,N_7693);
nor U8503 (N_8503,N_7391,N_7510);
nand U8504 (N_8504,N_7843,N_7204);
nor U8505 (N_8505,N_7913,N_7902);
xnor U8506 (N_8506,N_7931,N_7985);
or U8507 (N_8507,N_7722,N_7242);
nor U8508 (N_8508,N_7759,N_7760);
and U8509 (N_8509,N_7451,N_7338);
xnor U8510 (N_8510,N_7595,N_7261);
and U8511 (N_8511,N_7487,N_7443);
nand U8512 (N_8512,N_7734,N_7260);
nor U8513 (N_8513,N_7789,N_7366);
and U8514 (N_8514,N_7722,N_7627);
or U8515 (N_8515,N_7244,N_7963);
nand U8516 (N_8516,N_7350,N_7231);
nand U8517 (N_8517,N_7760,N_7821);
xnor U8518 (N_8518,N_7292,N_7696);
or U8519 (N_8519,N_7723,N_7884);
or U8520 (N_8520,N_7938,N_7262);
and U8521 (N_8521,N_7802,N_7670);
or U8522 (N_8522,N_7562,N_7566);
and U8523 (N_8523,N_7812,N_7861);
and U8524 (N_8524,N_7258,N_7443);
and U8525 (N_8525,N_7992,N_7940);
nor U8526 (N_8526,N_7481,N_7798);
and U8527 (N_8527,N_7264,N_7705);
or U8528 (N_8528,N_7227,N_7283);
or U8529 (N_8529,N_7281,N_7930);
nor U8530 (N_8530,N_7239,N_7937);
xor U8531 (N_8531,N_7366,N_7530);
and U8532 (N_8532,N_7540,N_7474);
nor U8533 (N_8533,N_7351,N_7649);
or U8534 (N_8534,N_7498,N_7628);
nand U8535 (N_8535,N_7280,N_7617);
nor U8536 (N_8536,N_7282,N_7476);
or U8537 (N_8537,N_7536,N_7367);
nand U8538 (N_8538,N_7325,N_7878);
and U8539 (N_8539,N_7214,N_7403);
nor U8540 (N_8540,N_7374,N_7309);
nand U8541 (N_8541,N_7672,N_7986);
nor U8542 (N_8542,N_7680,N_7738);
nand U8543 (N_8543,N_7919,N_7597);
nor U8544 (N_8544,N_7447,N_7338);
nor U8545 (N_8545,N_7539,N_7778);
nor U8546 (N_8546,N_7613,N_7237);
xor U8547 (N_8547,N_7408,N_7651);
nand U8548 (N_8548,N_7396,N_7394);
xnor U8549 (N_8549,N_7633,N_7858);
nand U8550 (N_8550,N_7851,N_7244);
and U8551 (N_8551,N_7820,N_7413);
nand U8552 (N_8552,N_7307,N_7865);
nor U8553 (N_8553,N_7773,N_7227);
and U8554 (N_8554,N_7963,N_7200);
or U8555 (N_8555,N_7759,N_7502);
nor U8556 (N_8556,N_7857,N_7587);
or U8557 (N_8557,N_7888,N_7891);
nor U8558 (N_8558,N_7359,N_7985);
xnor U8559 (N_8559,N_7241,N_7335);
and U8560 (N_8560,N_7216,N_7830);
nor U8561 (N_8561,N_7750,N_7965);
or U8562 (N_8562,N_7669,N_7993);
or U8563 (N_8563,N_7943,N_7570);
nand U8564 (N_8564,N_7306,N_7222);
nor U8565 (N_8565,N_7339,N_7286);
or U8566 (N_8566,N_7201,N_7860);
or U8567 (N_8567,N_7548,N_7804);
and U8568 (N_8568,N_7625,N_7982);
nor U8569 (N_8569,N_7956,N_7861);
xor U8570 (N_8570,N_7858,N_7234);
and U8571 (N_8571,N_7807,N_7956);
nor U8572 (N_8572,N_7772,N_7361);
nor U8573 (N_8573,N_7442,N_7752);
nor U8574 (N_8574,N_7416,N_7207);
or U8575 (N_8575,N_7569,N_7745);
nand U8576 (N_8576,N_7882,N_7755);
nand U8577 (N_8577,N_7834,N_7631);
xnor U8578 (N_8578,N_7658,N_7745);
xor U8579 (N_8579,N_7262,N_7678);
or U8580 (N_8580,N_7649,N_7711);
or U8581 (N_8581,N_7207,N_7985);
or U8582 (N_8582,N_7219,N_7469);
nor U8583 (N_8583,N_7418,N_7605);
or U8584 (N_8584,N_7300,N_7922);
nand U8585 (N_8585,N_7410,N_7584);
xor U8586 (N_8586,N_7439,N_7906);
nand U8587 (N_8587,N_7345,N_7794);
nor U8588 (N_8588,N_7559,N_7560);
nor U8589 (N_8589,N_7866,N_7563);
and U8590 (N_8590,N_7912,N_7591);
nor U8591 (N_8591,N_7297,N_7588);
and U8592 (N_8592,N_7979,N_7428);
nand U8593 (N_8593,N_7242,N_7628);
nand U8594 (N_8594,N_7413,N_7494);
xor U8595 (N_8595,N_7400,N_7233);
nor U8596 (N_8596,N_7389,N_7421);
and U8597 (N_8597,N_7938,N_7316);
or U8598 (N_8598,N_7595,N_7783);
or U8599 (N_8599,N_7364,N_7937);
nor U8600 (N_8600,N_7639,N_7283);
nor U8601 (N_8601,N_7875,N_7638);
nor U8602 (N_8602,N_7845,N_7320);
and U8603 (N_8603,N_7641,N_7403);
or U8604 (N_8604,N_7448,N_7830);
and U8605 (N_8605,N_7444,N_7892);
xnor U8606 (N_8606,N_7765,N_7408);
or U8607 (N_8607,N_7650,N_7542);
nand U8608 (N_8608,N_7947,N_7837);
nor U8609 (N_8609,N_7551,N_7508);
nor U8610 (N_8610,N_7499,N_7577);
or U8611 (N_8611,N_7677,N_7867);
nor U8612 (N_8612,N_7206,N_7491);
nand U8613 (N_8613,N_7666,N_7655);
nand U8614 (N_8614,N_7791,N_7844);
nor U8615 (N_8615,N_7929,N_7605);
nand U8616 (N_8616,N_7895,N_7918);
and U8617 (N_8617,N_7897,N_7872);
and U8618 (N_8618,N_7536,N_7789);
xor U8619 (N_8619,N_7642,N_7828);
nand U8620 (N_8620,N_7876,N_7376);
nor U8621 (N_8621,N_7205,N_7852);
nand U8622 (N_8622,N_7749,N_7738);
and U8623 (N_8623,N_7312,N_7288);
xnor U8624 (N_8624,N_7458,N_7619);
or U8625 (N_8625,N_7562,N_7347);
or U8626 (N_8626,N_7423,N_7362);
nor U8627 (N_8627,N_7599,N_7281);
nor U8628 (N_8628,N_7218,N_7397);
xnor U8629 (N_8629,N_7284,N_7233);
nor U8630 (N_8630,N_7594,N_7801);
or U8631 (N_8631,N_7813,N_7928);
nor U8632 (N_8632,N_7717,N_7759);
xnor U8633 (N_8633,N_7931,N_7958);
nand U8634 (N_8634,N_7766,N_7457);
nor U8635 (N_8635,N_7681,N_7953);
nor U8636 (N_8636,N_7405,N_7864);
xnor U8637 (N_8637,N_7653,N_7284);
nand U8638 (N_8638,N_7513,N_7316);
xnor U8639 (N_8639,N_7401,N_7988);
and U8640 (N_8640,N_7692,N_7241);
and U8641 (N_8641,N_7205,N_7816);
nor U8642 (N_8642,N_7744,N_7816);
nand U8643 (N_8643,N_7480,N_7940);
xor U8644 (N_8644,N_7589,N_7954);
or U8645 (N_8645,N_7965,N_7441);
nand U8646 (N_8646,N_7225,N_7412);
xnor U8647 (N_8647,N_7230,N_7992);
and U8648 (N_8648,N_7673,N_7989);
nor U8649 (N_8649,N_7460,N_7220);
xor U8650 (N_8650,N_7746,N_7256);
and U8651 (N_8651,N_7538,N_7795);
nor U8652 (N_8652,N_7377,N_7482);
or U8653 (N_8653,N_7618,N_7914);
nand U8654 (N_8654,N_7653,N_7726);
xnor U8655 (N_8655,N_7615,N_7204);
nand U8656 (N_8656,N_7796,N_7840);
and U8657 (N_8657,N_7897,N_7374);
or U8658 (N_8658,N_7880,N_7906);
xor U8659 (N_8659,N_7659,N_7483);
and U8660 (N_8660,N_7819,N_7955);
and U8661 (N_8661,N_7863,N_7241);
and U8662 (N_8662,N_7300,N_7837);
nor U8663 (N_8663,N_7526,N_7634);
and U8664 (N_8664,N_7470,N_7621);
xor U8665 (N_8665,N_7701,N_7708);
or U8666 (N_8666,N_7559,N_7457);
or U8667 (N_8667,N_7761,N_7218);
and U8668 (N_8668,N_7239,N_7598);
xor U8669 (N_8669,N_7657,N_7747);
nor U8670 (N_8670,N_7891,N_7718);
and U8671 (N_8671,N_7887,N_7553);
and U8672 (N_8672,N_7659,N_7863);
and U8673 (N_8673,N_7619,N_7621);
nand U8674 (N_8674,N_7419,N_7830);
xnor U8675 (N_8675,N_7329,N_7605);
and U8676 (N_8676,N_7320,N_7636);
xnor U8677 (N_8677,N_7407,N_7264);
nor U8678 (N_8678,N_7471,N_7536);
nand U8679 (N_8679,N_7339,N_7952);
nor U8680 (N_8680,N_7847,N_7678);
nand U8681 (N_8681,N_7476,N_7887);
xor U8682 (N_8682,N_7825,N_7982);
xnor U8683 (N_8683,N_7729,N_7424);
and U8684 (N_8684,N_7951,N_7656);
xor U8685 (N_8685,N_7243,N_7627);
xor U8686 (N_8686,N_7294,N_7372);
or U8687 (N_8687,N_7815,N_7939);
or U8688 (N_8688,N_7733,N_7942);
nor U8689 (N_8689,N_7800,N_7683);
nor U8690 (N_8690,N_7714,N_7590);
xor U8691 (N_8691,N_7749,N_7293);
and U8692 (N_8692,N_7459,N_7763);
nor U8693 (N_8693,N_7982,N_7880);
and U8694 (N_8694,N_7256,N_7366);
nor U8695 (N_8695,N_7300,N_7243);
nor U8696 (N_8696,N_7955,N_7587);
or U8697 (N_8697,N_7404,N_7773);
nand U8698 (N_8698,N_7642,N_7733);
xor U8699 (N_8699,N_7851,N_7533);
xnor U8700 (N_8700,N_7263,N_7429);
or U8701 (N_8701,N_7200,N_7491);
xnor U8702 (N_8702,N_7407,N_7643);
and U8703 (N_8703,N_7392,N_7612);
or U8704 (N_8704,N_7848,N_7790);
or U8705 (N_8705,N_7348,N_7655);
or U8706 (N_8706,N_7617,N_7744);
xor U8707 (N_8707,N_7268,N_7383);
nand U8708 (N_8708,N_7682,N_7383);
nor U8709 (N_8709,N_7491,N_7920);
nand U8710 (N_8710,N_7928,N_7716);
and U8711 (N_8711,N_7384,N_7583);
or U8712 (N_8712,N_7320,N_7905);
nand U8713 (N_8713,N_7932,N_7307);
nor U8714 (N_8714,N_7920,N_7268);
nor U8715 (N_8715,N_7306,N_7261);
nand U8716 (N_8716,N_7671,N_7888);
and U8717 (N_8717,N_7653,N_7996);
nor U8718 (N_8718,N_7339,N_7956);
and U8719 (N_8719,N_7522,N_7732);
or U8720 (N_8720,N_7921,N_7954);
or U8721 (N_8721,N_7440,N_7731);
nand U8722 (N_8722,N_7791,N_7578);
and U8723 (N_8723,N_7717,N_7414);
or U8724 (N_8724,N_7876,N_7396);
and U8725 (N_8725,N_7559,N_7443);
nand U8726 (N_8726,N_7398,N_7575);
nand U8727 (N_8727,N_7746,N_7967);
nand U8728 (N_8728,N_7886,N_7503);
nand U8729 (N_8729,N_7213,N_7666);
and U8730 (N_8730,N_7947,N_7622);
nor U8731 (N_8731,N_7665,N_7338);
and U8732 (N_8732,N_7922,N_7923);
and U8733 (N_8733,N_7752,N_7730);
or U8734 (N_8734,N_7824,N_7265);
and U8735 (N_8735,N_7854,N_7860);
nand U8736 (N_8736,N_7848,N_7996);
or U8737 (N_8737,N_7265,N_7640);
and U8738 (N_8738,N_7577,N_7426);
nor U8739 (N_8739,N_7409,N_7784);
nand U8740 (N_8740,N_7848,N_7817);
and U8741 (N_8741,N_7660,N_7593);
or U8742 (N_8742,N_7855,N_7262);
xnor U8743 (N_8743,N_7800,N_7907);
xor U8744 (N_8744,N_7774,N_7857);
or U8745 (N_8745,N_7999,N_7484);
or U8746 (N_8746,N_7517,N_7718);
nand U8747 (N_8747,N_7418,N_7407);
or U8748 (N_8748,N_7765,N_7506);
and U8749 (N_8749,N_7381,N_7460);
xnor U8750 (N_8750,N_7459,N_7218);
nor U8751 (N_8751,N_7655,N_7905);
nor U8752 (N_8752,N_7502,N_7540);
nor U8753 (N_8753,N_7806,N_7208);
and U8754 (N_8754,N_7618,N_7591);
nor U8755 (N_8755,N_7688,N_7587);
or U8756 (N_8756,N_7768,N_7891);
xor U8757 (N_8757,N_7851,N_7686);
xnor U8758 (N_8758,N_7411,N_7261);
and U8759 (N_8759,N_7799,N_7648);
or U8760 (N_8760,N_7972,N_7398);
or U8761 (N_8761,N_7608,N_7358);
nor U8762 (N_8762,N_7779,N_7717);
and U8763 (N_8763,N_7434,N_7244);
xor U8764 (N_8764,N_7928,N_7410);
and U8765 (N_8765,N_7621,N_7700);
xnor U8766 (N_8766,N_7470,N_7716);
nand U8767 (N_8767,N_7611,N_7867);
and U8768 (N_8768,N_7951,N_7925);
nor U8769 (N_8769,N_7418,N_7905);
xor U8770 (N_8770,N_7264,N_7647);
and U8771 (N_8771,N_7465,N_7951);
and U8772 (N_8772,N_7667,N_7571);
nor U8773 (N_8773,N_7474,N_7276);
or U8774 (N_8774,N_7353,N_7832);
xnor U8775 (N_8775,N_7768,N_7709);
nand U8776 (N_8776,N_7492,N_7667);
or U8777 (N_8777,N_7288,N_7501);
or U8778 (N_8778,N_7414,N_7673);
or U8779 (N_8779,N_7230,N_7592);
or U8780 (N_8780,N_7604,N_7523);
xor U8781 (N_8781,N_7321,N_7292);
nor U8782 (N_8782,N_7975,N_7703);
xor U8783 (N_8783,N_7703,N_7264);
xor U8784 (N_8784,N_7625,N_7986);
and U8785 (N_8785,N_7573,N_7511);
or U8786 (N_8786,N_7978,N_7814);
xnor U8787 (N_8787,N_7902,N_7824);
and U8788 (N_8788,N_7920,N_7629);
or U8789 (N_8789,N_7868,N_7237);
xnor U8790 (N_8790,N_7369,N_7677);
xor U8791 (N_8791,N_7582,N_7363);
and U8792 (N_8792,N_7573,N_7380);
and U8793 (N_8793,N_7735,N_7206);
nor U8794 (N_8794,N_7701,N_7662);
xor U8795 (N_8795,N_7488,N_7812);
or U8796 (N_8796,N_7832,N_7699);
and U8797 (N_8797,N_7646,N_7937);
nand U8798 (N_8798,N_7914,N_7298);
xnor U8799 (N_8799,N_7478,N_7499);
nand U8800 (N_8800,N_8202,N_8068);
and U8801 (N_8801,N_8584,N_8115);
and U8802 (N_8802,N_8407,N_8253);
nand U8803 (N_8803,N_8344,N_8363);
and U8804 (N_8804,N_8266,N_8170);
xnor U8805 (N_8805,N_8587,N_8576);
or U8806 (N_8806,N_8108,N_8753);
nand U8807 (N_8807,N_8606,N_8769);
or U8808 (N_8808,N_8163,N_8403);
xnor U8809 (N_8809,N_8348,N_8455);
xnor U8810 (N_8810,N_8744,N_8159);
nand U8811 (N_8811,N_8129,N_8719);
nand U8812 (N_8812,N_8454,N_8689);
or U8813 (N_8813,N_8405,N_8377);
nand U8814 (N_8814,N_8514,N_8140);
and U8815 (N_8815,N_8730,N_8349);
nor U8816 (N_8816,N_8201,N_8300);
xor U8817 (N_8817,N_8641,N_8620);
or U8818 (N_8818,N_8192,N_8729);
nand U8819 (N_8819,N_8207,N_8145);
xnor U8820 (N_8820,N_8604,N_8590);
and U8821 (N_8821,N_8530,N_8197);
or U8822 (N_8822,N_8570,N_8413);
nand U8823 (N_8823,N_8128,N_8257);
and U8824 (N_8824,N_8165,N_8489);
and U8825 (N_8825,N_8658,N_8143);
and U8826 (N_8826,N_8338,N_8668);
and U8827 (N_8827,N_8303,N_8011);
and U8828 (N_8828,N_8282,N_8473);
and U8829 (N_8829,N_8162,N_8182);
xnor U8830 (N_8830,N_8275,N_8085);
or U8831 (N_8831,N_8628,N_8718);
and U8832 (N_8832,N_8336,N_8123);
xnor U8833 (N_8833,N_8644,N_8397);
or U8834 (N_8834,N_8208,N_8311);
xnor U8835 (N_8835,N_8404,N_8623);
and U8836 (N_8836,N_8146,N_8660);
or U8837 (N_8837,N_8515,N_8786);
nand U8838 (N_8838,N_8597,N_8245);
or U8839 (N_8839,N_8542,N_8635);
or U8840 (N_8840,N_8087,N_8567);
nor U8841 (N_8841,N_8012,N_8083);
xor U8842 (N_8842,N_8160,N_8610);
or U8843 (N_8843,N_8575,N_8181);
nor U8844 (N_8844,N_8399,N_8588);
xnor U8845 (N_8845,N_8156,N_8410);
nor U8846 (N_8846,N_8780,N_8010);
or U8847 (N_8847,N_8713,N_8234);
or U8848 (N_8848,N_8395,N_8130);
or U8849 (N_8849,N_8464,N_8287);
xnor U8850 (N_8850,N_8703,N_8414);
xnor U8851 (N_8851,N_8033,N_8366);
xnor U8852 (N_8852,N_8390,N_8560);
nor U8853 (N_8853,N_8497,N_8273);
nand U8854 (N_8854,N_8070,N_8465);
nor U8855 (N_8855,N_8652,N_8500);
and U8856 (N_8856,N_8425,N_8158);
xor U8857 (N_8857,N_8081,N_8037);
nand U8858 (N_8858,N_8193,N_8431);
and U8859 (N_8859,N_8639,N_8712);
nor U8860 (N_8860,N_8482,N_8215);
or U8861 (N_8861,N_8750,N_8647);
xor U8862 (N_8862,N_8651,N_8428);
nand U8863 (N_8863,N_8762,N_8002);
xor U8864 (N_8864,N_8100,N_8239);
nor U8865 (N_8865,N_8286,N_8490);
nand U8866 (N_8866,N_8132,N_8634);
nand U8867 (N_8867,N_8330,N_8749);
or U8868 (N_8868,N_8320,N_8675);
and U8869 (N_8869,N_8793,N_8408);
and U8870 (N_8870,N_8378,N_8552);
nand U8871 (N_8871,N_8095,N_8035);
or U8872 (N_8872,N_8080,N_8327);
nand U8873 (N_8873,N_8737,N_8358);
nand U8874 (N_8874,N_8000,N_8781);
nor U8875 (N_8875,N_8219,N_8477);
or U8876 (N_8876,N_8723,N_8369);
nand U8877 (N_8877,N_8797,N_8732);
and U8878 (N_8878,N_8496,N_8415);
nor U8879 (N_8879,N_8633,N_8186);
or U8880 (N_8880,N_8581,N_8671);
or U8881 (N_8881,N_8400,N_8721);
or U8882 (N_8882,N_8183,N_8487);
or U8883 (N_8883,N_8701,N_8442);
nor U8884 (N_8884,N_8134,N_8558);
or U8885 (N_8885,N_8184,N_8638);
or U8886 (N_8886,N_8784,N_8393);
and U8887 (N_8887,N_8476,N_8285);
nand U8888 (N_8888,N_8195,N_8064);
nor U8889 (N_8889,N_8006,N_8645);
or U8890 (N_8890,N_8227,N_8724);
nand U8891 (N_8891,N_8507,N_8044);
or U8892 (N_8892,N_8502,N_8655);
xor U8893 (N_8893,N_8448,N_8516);
nor U8894 (N_8894,N_8328,N_8102);
and U8895 (N_8895,N_8602,N_8302);
nand U8896 (N_8896,N_8040,N_8025);
nor U8897 (N_8897,N_8682,N_8359);
and U8898 (N_8898,N_8636,N_8775);
and U8899 (N_8899,N_8392,N_8746);
nand U8900 (N_8900,N_8458,N_8056);
nor U8901 (N_8901,N_8733,N_8614);
nand U8902 (N_8902,N_8013,N_8131);
xor U8903 (N_8903,N_8173,N_8767);
xor U8904 (N_8904,N_8446,N_8007);
or U8905 (N_8905,N_8382,N_8466);
xnor U8906 (N_8906,N_8371,N_8295);
nor U8907 (N_8907,N_8662,N_8356);
nand U8908 (N_8908,N_8074,N_8423);
xnor U8909 (N_8909,N_8435,N_8650);
and U8910 (N_8910,N_8726,N_8450);
nand U8911 (N_8911,N_8376,N_8406);
nor U8912 (N_8912,N_8770,N_8761);
and U8913 (N_8913,N_8568,N_8351);
nor U8914 (N_8914,N_8149,N_8709);
xor U8915 (N_8915,N_8504,N_8562);
nand U8916 (N_8916,N_8757,N_8795);
and U8917 (N_8917,N_8688,N_8113);
and U8918 (N_8918,N_8642,N_8783);
or U8919 (N_8919,N_8079,N_8772);
nor U8920 (N_8920,N_8151,N_8596);
xor U8921 (N_8921,N_8622,N_8028);
or U8922 (N_8922,N_8362,N_8787);
nor U8923 (N_8923,N_8294,N_8608);
xor U8924 (N_8924,N_8189,N_8734);
or U8925 (N_8925,N_8307,N_8155);
or U8926 (N_8926,N_8547,N_8677);
nand U8927 (N_8927,N_8544,N_8727);
nor U8928 (N_8928,N_8523,N_8096);
xor U8929 (N_8929,N_8191,N_8290);
or U8930 (N_8930,N_8402,N_8672);
or U8931 (N_8931,N_8598,N_8763);
xor U8932 (N_8932,N_8243,N_8133);
or U8933 (N_8933,N_8698,N_8276);
xor U8934 (N_8934,N_8117,N_8251);
or U8935 (N_8935,N_8069,N_8052);
nand U8936 (N_8936,N_8077,N_8493);
xnor U8937 (N_8937,N_8053,N_8538);
nor U8938 (N_8938,N_8019,N_8443);
nand U8939 (N_8939,N_8441,N_8126);
and U8940 (N_8940,N_8518,N_8419);
nand U8941 (N_8941,N_8475,N_8764);
and U8942 (N_8942,N_8522,N_8765);
nand U8943 (N_8943,N_8714,N_8009);
nor U8944 (N_8944,N_8657,N_8034);
and U8945 (N_8945,N_8691,N_8334);
and U8946 (N_8946,N_8297,N_8339);
xnor U8947 (N_8947,N_8340,N_8078);
nor U8948 (N_8948,N_8372,N_8495);
nor U8949 (N_8949,N_8292,N_8768);
or U8950 (N_8950,N_8244,N_8664);
nor U8951 (N_8951,N_8648,N_8469);
nor U8952 (N_8952,N_8274,N_8209);
xnor U8953 (N_8953,N_8022,N_8293);
nand U8954 (N_8954,N_8778,N_8388);
nor U8955 (N_8955,N_8488,N_8663);
or U8956 (N_8956,N_8073,N_8252);
nand U8957 (N_8957,N_8699,N_8609);
xor U8958 (N_8958,N_8260,N_8016);
nand U8959 (N_8959,N_8106,N_8176);
or U8960 (N_8960,N_8799,N_8343);
nand U8961 (N_8961,N_8326,N_8157);
xnor U8962 (N_8962,N_8531,N_8433);
nor U8963 (N_8963,N_8686,N_8178);
or U8964 (N_8964,N_8629,N_8105);
and U8965 (N_8965,N_8386,N_8271);
nor U8966 (N_8966,N_8103,N_8508);
xor U8967 (N_8967,N_8312,N_8472);
nand U8968 (N_8968,N_8550,N_8017);
nor U8969 (N_8969,N_8687,N_8247);
nand U8970 (N_8970,N_8478,N_8439);
or U8971 (N_8971,N_8391,N_8137);
nand U8972 (N_8972,N_8221,N_8461);
nand U8973 (N_8973,N_8357,N_8583);
nor U8974 (N_8974,N_8429,N_8580);
nand U8975 (N_8975,N_8166,N_8259);
or U8976 (N_8976,N_8440,N_8409);
or U8977 (N_8977,N_8118,N_8537);
or U8978 (N_8978,N_8485,N_8211);
nor U8979 (N_8979,N_8084,N_8317);
and U8980 (N_8980,N_8229,N_8745);
nand U8981 (N_8981,N_8352,N_8536);
nor U8982 (N_8982,N_8373,N_8059);
and U8983 (N_8983,N_8420,N_8449);
nor U8984 (N_8984,N_8654,N_8171);
xnor U8985 (N_8985,N_8617,N_8179);
xnor U8986 (N_8986,N_8319,N_8298);
nand U8987 (N_8987,N_8527,N_8578);
and U8988 (N_8988,N_8685,N_8154);
xnor U8989 (N_8989,N_8572,N_8548);
nor U8990 (N_8990,N_8135,N_8557);
xor U8991 (N_8991,N_8444,N_8705);
and U8992 (N_8992,N_8364,N_8055);
xor U8993 (N_8993,N_8088,N_8172);
or U8994 (N_8994,N_8099,N_8418);
nand U8995 (N_8995,N_8329,N_8659);
or U8996 (N_8996,N_8272,N_8725);
nand U8997 (N_8997,N_8296,N_8754);
nand U8998 (N_8998,N_8226,N_8667);
nor U8999 (N_8999,N_8127,N_8041);
nand U9000 (N_9000,N_8177,N_8569);
and U9001 (N_9001,N_8314,N_8354);
and U9002 (N_9002,N_8457,N_8759);
xnor U9003 (N_9003,N_8785,N_8062);
xor U9004 (N_9004,N_8566,N_8223);
or U9005 (N_9005,N_8057,N_8679);
or U9006 (N_9006,N_8299,N_8014);
nand U9007 (N_9007,N_8666,N_8212);
or U9008 (N_9008,N_8445,N_8540);
xor U9009 (N_9009,N_8199,N_8249);
nor U9010 (N_9010,N_8573,N_8467);
xor U9011 (N_9011,N_8605,N_8791);
or U9012 (N_9012,N_8061,N_8438);
nand U9013 (N_9013,N_8198,N_8039);
xnor U9014 (N_9014,N_8646,N_8242);
nand U9015 (N_9015,N_8385,N_8342);
xor U9016 (N_9016,N_8152,N_8023);
and U9017 (N_9017,N_8470,N_8318);
or U9018 (N_9018,N_8690,N_8396);
and U9019 (N_9019,N_8355,N_8661);
nor U9020 (N_9020,N_8751,N_8291);
xnor U9021 (N_9021,N_8107,N_8093);
or U9022 (N_9022,N_8174,N_8111);
or U9023 (N_9023,N_8046,N_8038);
or U9024 (N_9024,N_8519,N_8365);
or U9025 (N_9025,N_8031,N_8238);
or U9026 (N_9026,N_8164,N_8036);
or U9027 (N_9027,N_8109,N_8593);
or U9028 (N_9028,N_8072,N_8559);
nor U9029 (N_9029,N_8771,N_8313);
xnor U9030 (N_9030,N_8571,N_8513);
xnor U9031 (N_9031,N_8517,N_8563);
xor U9032 (N_9032,N_8412,N_8250);
nor U9033 (N_9033,N_8486,N_8091);
nand U9034 (N_9034,N_8345,N_8112);
and U9035 (N_9035,N_8743,N_8268);
nand U9036 (N_9036,N_8119,N_8760);
xor U9037 (N_9037,N_8187,N_8777);
and U9038 (N_9038,N_8051,N_8674);
nor U9039 (N_9039,N_8389,N_8706);
nand U9040 (N_9040,N_8564,N_8310);
and U9041 (N_9041,N_8471,N_8535);
and U9042 (N_9042,N_8521,N_8416);
and U9043 (N_9043,N_8462,N_8353);
or U9044 (N_9044,N_8230,N_8381);
and U9045 (N_9045,N_8694,N_8316);
nor U9046 (N_9046,N_8168,N_8139);
or U9047 (N_9047,N_8700,N_8141);
or U9048 (N_9048,N_8032,N_8774);
and U9049 (N_9049,N_8335,N_8283);
or U9050 (N_9050,N_8256,N_8539);
or U9051 (N_9051,N_8030,N_8434);
xor U9052 (N_9052,N_8379,N_8265);
and U9053 (N_9053,N_8427,N_8175);
nor U9054 (N_9054,N_8255,N_8543);
nor U9055 (N_9055,N_8447,N_8267);
or U9056 (N_9056,N_8161,N_8185);
nand U9057 (N_9057,N_8621,N_8739);
nor U9058 (N_9058,N_8167,N_8001);
and U9059 (N_9059,N_8090,N_8015);
nand U9060 (N_9060,N_8738,N_8098);
or U9061 (N_9061,N_8360,N_8630);
and U9062 (N_9062,N_8625,N_8148);
nor U9063 (N_9063,N_8577,N_8218);
nor U9064 (N_9064,N_8480,N_8284);
xnor U9065 (N_9065,N_8341,N_8528);
xor U9066 (N_9066,N_8796,N_8600);
or U9067 (N_9067,N_8708,N_8067);
or U9068 (N_9068,N_8411,N_8254);
or U9069 (N_9069,N_8220,N_8323);
and U9070 (N_9070,N_8720,N_8479);
nand U9071 (N_9071,N_8231,N_8054);
nor U9072 (N_9072,N_8262,N_8766);
nor U9073 (N_9073,N_8616,N_8735);
or U9074 (N_9074,N_8094,N_8526);
and U9075 (N_9075,N_8144,N_8018);
nand U9076 (N_9076,N_8499,N_8370);
and U9077 (N_9077,N_8520,N_8501);
nand U9078 (N_9078,N_8716,N_8432);
nand U9079 (N_9079,N_8269,N_8387);
or U9080 (N_9080,N_8153,N_8050);
or U9081 (N_9081,N_8782,N_8075);
xnor U9082 (N_9082,N_8509,N_8024);
nand U9083 (N_9083,N_8758,N_8384);
xnor U9084 (N_9084,N_8676,N_8204);
nor U9085 (N_9085,N_8451,N_8368);
nand U9086 (N_9086,N_8715,N_8599);
and U9087 (N_9087,N_8665,N_8790);
or U9088 (N_9088,N_8756,N_8545);
xnor U9089 (N_9089,N_8346,N_8524);
and U9090 (N_9090,N_8532,N_8203);
xnor U9091 (N_9091,N_8188,N_8066);
and U9092 (N_9092,N_8607,N_8696);
nand U9093 (N_9093,N_8048,N_8142);
and U9094 (N_9094,N_8506,N_8436);
xor U9095 (N_9095,N_8643,N_8792);
xnor U9096 (N_9096,N_8322,N_8492);
nand U9097 (N_9097,N_8005,N_8277);
xnor U9098 (N_9098,N_8511,N_8683);
or U9099 (N_9099,N_8225,N_8640);
or U9100 (N_9100,N_8586,N_8213);
and U9101 (N_9101,N_8589,N_8301);
nor U9102 (N_9102,N_8460,N_8612);
nor U9103 (N_9103,N_8484,N_8280);
nand U9104 (N_9104,N_8248,N_8263);
and U9105 (N_9105,N_8337,N_8624);
or U9106 (N_9106,N_8710,N_8711);
nor U9107 (N_9107,N_8210,N_8190);
xor U9108 (N_9108,N_8742,N_8553);
and U9109 (N_9109,N_8541,N_8731);
and U9110 (N_9110,N_8430,N_8049);
or U9111 (N_9111,N_8670,N_8422);
or U9112 (N_9112,N_8678,N_8585);
or U9113 (N_9113,N_8288,N_8681);
or U9114 (N_9114,N_8684,N_8045);
and U9115 (N_9115,N_8456,N_8169);
nor U9116 (N_9116,N_8626,N_8306);
nor U9117 (N_9117,N_8082,N_8003);
nand U9118 (N_9118,N_8529,N_8374);
and U9119 (N_9119,N_8494,N_8089);
nor U9120 (N_9120,N_8021,N_8525);
nand U9121 (N_9121,N_8752,N_8261);
nor U9122 (N_9122,N_8398,N_8755);
nand U9123 (N_9123,N_8579,N_8324);
and U9124 (N_9124,N_8637,N_8121);
nor U9125 (N_9125,N_8228,N_8549);
or U9126 (N_9126,N_8788,N_8206);
and U9127 (N_9127,N_8217,N_8058);
and U9128 (N_9128,N_8264,N_8008);
xnor U9129 (N_9129,N_8063,N_8669);
or U9130 (N_9130,N_8483,N_8047);
or U9131 (N_9131,N_8196,N_8592);
or U9132 (N_9132,N_8595,N_8350);
nand U9133 (N_9133,N_8779,N_8618);
nor U9134 (N_9134,N_8534,N_8125);
nor U9135 (N_9135,N_8512,N_8114);
and U9136 (N_9136,N_8383,N_8332);
xnor U9137 (N_9137,N_8503,N_8321);
or U9138 (N_9138,N_8122,N_8594);
nand U9139 (N_9139,N_8554,N_8697);
nand U9140 (N_9140,N_8120,N_8104);
nand U9141 (N_9141,N_8693,N_8305);
or U9142 (N_9142,N_8235,N_8510);
nand U9143 (N_9143,N_8736,N_8491);
nand U9144 (N_9144,N_8424,N_8308);
and U9145 (N_9145,N_8246,N_8279);
and U9146 (N_9146,N_8498,N_8653);
or U9147 (N_9147,N_8707,N_8060);
or U9148 (N_9148,N_8020,N_8546);
and U9149 (N_9149,N_8728,N_8582);
or U9150 (N_9150,N_8237,N_8071);
and U9151 (N_9151,N_8632,N_8097);
nor U9152 (N_9152,N_8222,N_8722);
nand U9153 (N_9153,N_8794,N_8043);
nor U9154 (N_9154,N_8695,N_8333);
nand U9155 (N_9155,N_8331,N_8101);
nor U9156 (N_9156,N_8555,N_8551);
xnor U9157 (N_9157,N_8401,N_8656);
nand U9158 (N_9158,N_8673,N_8042);
nor U9159 (N_9159,N_8325,N_8026);
xor U9160 (N_9160,N_8240,N_8086);
nor U9161 (N_9161,N_8232,N_8601);
xor U9162 (N_9162,N_8027,N_8347);
or U9163 (N_9163,N_8361,N_8748);
nand U9164 (N_9164,N_8315,N_8704);
nor U9165 (N_9165,N_8281,N_8453);
xnor U9166 (N_9166,N_8004,N_8776);
or U9167 (N_9167,N_8138,N_8241);
or U9168 (N_9168,N_8110,N_8505);
and U9169 (N_9169,N_8789,N_8216);
or U9170 (N_9170,N_8613,N_8574);
nor U9171 (N_9171,N_8309,N_8065);
xnor U9172 (N_9172,N_8692,N_8417);
xnor U9173 (N_9173,N_8147,N_8741);
nor U9174 (N_9174,N_8463,N_8136);
and U9175 (N_9175,N_8615,N_8200);
nand U9176 (N_9176,N_8627,N_8533);
nand U9177 (N_9177,N_8224,N_8561);
xor U9178 (N_9178,N_8375,N_8565);
and U9179 (N_9179,N_8631,N_8740);
xnor U9180 (N_9180,N_8180,N_8233);
or U9181 (N_9181,N_8258,N_8214);
xor U9182 (N_9182,N_8304,N_8798);
nor U9183 (N_9183,N_8747,N_8421);
and U9184 (N_9184,N_8270,N_8367);
nand U9185 (N_9185,N_8426,N_8194);
nor U9186 (N_9186,N_8437,N_8076);
and U9187 (N_9187,N_8459,N_8556);
nand U9188 (N_9188,N_8649,N_8394);
or U9189 (N_9189,N_8092,N_8452);
xor U9190 (N_9190,N_8680,N_8481);
nand U9191 (N_9191,N_8603,N_8474);
nor U9192 (N_9192,N_8278,N_8611);
or U9193 (N_9193,N_8150,N_8619);
xnor U9194 (N_9194,N_8380,N_8116);
and U9195 (N_9195,N_8591,N_8029);
or U9196 (N_9196,N_8468,N_8717);
xnor U9197 (N_9197,N_8124,N_8289);
and U9198 (N_9198,N_8773,N_8702);
and U9199 (N_9199,N_8236,N_8205);
and U9200 (N_9200,N_8786,N_8305);
xor U9201 (N_9201,N_8340,N_8383);
and U9202 (N_9202,N_8284,N_8324);
nand U9203 (N_9203,N_8265,N_8198);
nor U9204 (N_9204,N_8263,N_8314);
nand U9205 (N_9205,N_8668,N_8497);
nor U9206 (N_9206,N_8248,N_8556);
and U9207 (N_9207,N_8522,N_8456);
nor U9208 (N_9208,N_8752,N_8411);
xnor U9209 (N_9209,N_8690,N_8634);
nand U9210 (N_9210,N_8457,N_8216);
nand U9211 (N_9211,N_8717,N_8745);
nor U9212 (N_9212,N_8644,N_8695);
or U9213 (N_9213,N_8769,N_8354);
nand U9214 (N_9214,N_8670,N_8550);
and U9215 (N_9215,N_8541,N_8226);
nand U9216 (N_9216,N_8537,N_8067);
nor U9217 (N_9217,N_8476,N_8007);
and U9218 (N_9218,N_8225,N_8037);
xnor U9219 (N_9219,N_8428,N_8203);
nor U9220 (N_9220,N_8689,N_8617);
nand U9221 (N_9221,N_8210,N_8605);
nor U9222 (N_9222,N_8034,N_8652);
or U9223 (N_9223,N_8610,N_8055);
nand U9224 (N_9224,N_8648,N_8310);
and U9225 (N_9225,N_8019,N_8067);
xnor U9226 (N_9226,N_8379,N_8452);
or U9227 (N_9227,N_8176,N_8126);
nor U9228 (N_9228,N_8424,N_8659);
nor U9229 (N_9229,N_8386,N_8072);
xnor U9230 (N_9230,N_8381,N_8265);
nand U9231 (N_9231,N_8311,N_8721);
or U9232 (N_9232,N_8123,N_8378);
or U9233 (N_9233,N_8139,N_8525);
or U9234 (N_9234,N_8171,N_8571);
or U9235 (N_9235,N_8525,N_8136);
nor U9236 (N_9236,N_8666,N_8667);
xnor U9237 (N_9237,N_8076,N_8054);
nor U9238 (N_9238,N_8595,N_8610);
nand U9239 (N_9239,N_8145,N_8132);
or U9240 (N_9240,N_8462,N_8436);
nor U9241 (N_9241,N_8227,N_8182);
or U9242 (N_9242,N_8248,N_8629);
or U9243 (N_9243,N_8587,N_8535);
xor U9244 (N_9244,N_8408,N_8611);
nand U9245 (N_9245,N_8582,N_8072);
xor U9246 (N_9246,N_8046,N_8034);
or U9247 (N_9247,N_8315,N_8128);
nand U9248 (N_9248,N_8551,N_8487);
and U9249 (N_9249,N_8424,N_8299);
nor U9250 (N_9250,N_8347,N_8526);
nand U9251 (N_9251,N_8109,N_8369);
nor U9252 (N_9252,N_8231,N_8629);
or U9253 (N_9253,N_8192,N_8454);
xnor U9254 (N_9254,N_8279,N_8735);
nand U9255 (N_9255,N_8614,N_8363);
nor U9256 (N_9256,N_8695,N_8110);
and U9257 (N_9257,N_8098,N_8786);
nor U9258 (N_9258,N_8088,N_8593);
nor U9259 (N_9259,N_8374,N_8393);
and U9260 (N_9260,N_8680,N_8560);
or U9261 (N_9261,N_8338,N_8361);
xor U9262 (N_9262,N_8632,N_8264);
nand U9263 (N_9263,N_8110,N_8298);
and U9264 (N_9264,N_8254,N_8394);
and U9265 (N_9265,N_8012,N_8762);
nor U9266 (N_9266,N_8498,N_8166);
nor U9267 (N_9267,N_8368,N_8277);
or U9268 (N_9268,N_8566,N_8140);
nand U9269 (N_9269,N_8197,N_8246);
nand U9270 (N_9270,N_8288,N_8767);
xnor U9271 (N_9271,N_8160,N_8716);
or U9272 (N_9272,N_8653,N_8035);
and U9273 (N_9273,N_8315,N_8214);
and U9274 (N_9274,N_8797,N_8274);
or U9275 (N_9275,N_8693,N_8740);
nand U9276 (N_9276,N_8775,N_8407);
and U9277 (N_9277,N_8509,N_8105);
nor U9278 (N_9278,N_8134,N_8711);
nand U9279 (N_9279,N_8725,N_8624);
or U9280 (N_9280,N_8764,N_8212);
and U9281 (N_9281,N_8324,N_8455);
and U9282 (N_9282,N_8642,N_8471);
xor U9283 (N_9283,N_8669,N_8600);
and U9284 (N_9284,N_8423,N_8252);
or U9285 (N_9285,N_8771,N_8770);
xnor U9286 (N_9286,N_8645,N_8475);
nor U9287 (N_9287,N_8271,N_8392);
nand U9288 (N_9288,N_8154,N_8384);
or U9289 (N_9289,N_8342,N_8475);
xor U9290 (N_9290,N_8231,N_8745);
or U9291 (N_9291,N_8583,N_8084);
nor U9292 (N_9292,N_8542,N_8353);
and U9293 (N_9293,N_8209,N_8493);
or U9294 (N_9294,N_8613,N_8026);
nand U9295 (N_9295,N_8457,N_8518);
and U9296 (N_9296,N_8338,N_8232);
nor U9297 (N_9297,N_8035,N_8043);
nand U9298 (N_9298,N_8014,N_8569);
xnor U9299 (N_9299,N_8113,N_8793);
nor U9300 (N_9300,N_8189,N_8693);
nand U9301 (N_9301,N_8631,N_8052);
nand U9302 (N_9302,N_8246,N_8352);
and U9303 (N_9303,N_8203,N_8775);
nor U9304 (N_9304,N_8406,N_8753);
or U9305 (N_9305,N_8713,N_8569);
and U9306 (N_9306,N_8516,N_8615);
nor U9307 (N_9307,N_8394,N_8003);
nand U9308 (N_9308,N_8753,N_8658);
and U9309 (N_9309,N_8141,N_8143);
or U9310 (N_9310,N_8000,N_8240);
nand U9311 (N_9311,N_8731,N_8430);
or U9312 (N_9312,N_8626,N_8410);
nor U9313 (N_9313,N_8669,N_8024);
xnor U9314 (N_9314,N_8030,N_8250);
nor U9315 (N_9315,N_8755,N_8306);
nand U9316 (N_9316,N_8731,N_8083);
nand U9317 (N_9317,N_8670,N_8223);
nand U9318 (N_9318,N_8154,N_8690);
or U9319 (N_9319,N_8277,N_8688);
nor U9320 (N_9320,N_8462,N_8252);
or U9321 (N_9321,N_8179,N_8590);
xnor U9322 (N_9322,N_8545,N_8532);
xor U9323 (N_9323,N_8245,N_8328);
nor U9324 (N_9324,N_8656,N_8625);
and U9325 (N_9325,N_8094,N_8553);
nand U9326 (N_9326,N_8329,N_8221);
and U9327 (N_9327,N_8518,N_8559);
nor U9328 (N_9328,N_8257,N_8662);
and U9329 (N_9329,N_8262,N_8269);
nor U9330 (N_9330,N_8264,N_8372);
and U9331 (N_9331,N_8074,N_8700);
xor U9332 (N_9332,N_8699,N_8433);
or U9333 (N_9333,N_8725,N_8524);
nand U9334 (N_9334,N_8641,N_8061);
and U9335 (N_9335,N_8194,N_8318);
or U9336 (N_9336,N_8621,N_8016);
xor U9337 (N_9337,N_8160,N_8256);
or U9338 (N_9338,N_8047,N_8793);
or U9339 (N_9339,N_8382,N_8517);
or U9340 (N_9340,N_8451,N_8511);
or U9341 (N_9341,N_8343,N_8200);
nor U9342 (N_9342,N_8733,N_8112);
and U9343 (N_9343,N_8312,N_8177);
xnor U9344 (N_9344,N_8641,N_8388);
nand U9345 (N_9345,N_8006,N_8288);
nand U9346 (N_9346,N_8058,N_8626);
nand U9347 (N_9347,N_8426,N_8722);
or U9348 (N_9348,N_8514,N_8486);
and U9349 (N_9349,N_8697,N_8490);
or U9350 (N_9350,N_8098,N_8159);
and U9351 (N_9351,N_8632,N_8348);
or U9352 (N_9352,N_8196,N_8194);
nand U9353 (N_9353,N_8511,N_8216);
and U9354 (N_9354,N_8668,N_8683);
and U9355 (N_9355,N_8223,N_8021);
nor U9356 (N_9356,N_8358,N_8198);
nand U9357 (N_9357,N_8430,N_8214);
and U9358 (N_9358,N_8728,N_8672);
xnor U9359 (N_9359,N_8508,N_8394);
or U9360 (N_9360,N_8251,N_8715);
or U9361 (N_9361,N_8775,N_8422);
and U9362 (N_9362,N_8262,N_8196);
xnor U9363 (N_9363,N_8381,N_8512);
nor U9364 (N_9364,N_8526,N_8427);
nand U9365 (N_9365,N_8707,N_8342);
nand U9366 (N_9366,N_8222,N_8083);
and U9367 (N_9367,N_8414,N_8721);
nor U9368 (N_9368,N_8723,N_8373);
or U9369 (N_9369,N_8352,N_8343);
nor U9370 (N_9370,N_8787,N_8022);
nor U9371 (N_9371,N_8659,N_8092);
xor U9372 (N_9372,N_8519,N_8685);
or U9373 (N_9373,N_8713,N_8454);
or U9374 (N_9374,N_8392,N_8006);
or U9375 (N_9375,N_8728,N_8124);
nor U9376 (N_9376,N_8427,N_8040);
nor U9377 (N_9377,N_8636,N_8128);
or U9378 (N_9378,N_8192,N_8484);
nand U9379 (N_9379,N_8242,N_8363);
nand U9380 (N_9380,N_8209,N_8671);
and U9381 (N_9381,N_8585,N_8264);
nand U9382 (N_9382,N_8483,N_8344);
and U9383 (N_9383,N_8732,N_8116);
nand U9384 (N_9384,N_8663,N_8446);
or U9385 (N_9385,N_8531,N_8427);
or U9386 (N_9386,N_8106,N_8419);
nand U9387 (N_9387,N_8321,N_8315);
or U9388 (N_9388,N_8767,N_8531);
or U9389 (N_9389,N_8532,N_8780);
or U9390 (N_9390,N_8407,N_8258);
and U9391 (N_9391,N_8756,N_8379);
xor U9392 (N_9392,N_8535,N_8795);
nand U9393 (N_9393,N_8773,N_8369);
and U9394 (N_9394,N_8604,N_8287);
or U9395 (N_9395,N_8468,N_8703);
nor U9396 (N_9396,N_8262,N_8251);
nand U9397 (N_9397,N_8267,N_8513);
and U9398 (N_9398,N_8214,N_8444);
nor U9399 (N_9399,N_8734,N_8394);
xor U9400 (N_9400,N_8354,N_8296);
xnor U9401 (N_9401,N_8044,N_8337);
and U9402 (N_9402,N_8485,N_8666);
xnor U9403 (N_9403,N_8618,N_8174);
nor U9404 (N_9404,N_8679,N_8105);
nor U9405 (N_9405,N_8280,N_8474);
or U9406 (N_9406,N_8241,N_8007);
or U9407 (N_9407,N_8636,N_8370);
nand U9408 (N_9408,N_8115,N_8769);
nor U9409 (N_9409,N_8396,N_8785);
and U9410 (N_9410,N_8125,N_8146);
or U9411 (N_9411,N_8039,N_8169);
xor U9412 (N_9412,N_8492,N_8464);
and U9413 (N_9413,N_8519,N_8159);
xnor U9414 (N_9414,N_8494,N_8274);
or U9415 (N_9415,N_8621,N_8235);
xor U9416 (N_9416,N_8191,N_8527);
or U9417 (N_9417,N_8518,N_8085);
or U9418 (N_9418,N_8783,N_8115);
and U9419 (N_9419,N_8648,N_8321);
nand U9420 (N_9420,N_8787,N_8329);
nand U9421 (N_9421,N_8136,N_8537);
xor U9422 (N_9422,N_8665,N_8516);
nor U9423 (N_9423,N_8120,N_8155);
or U9424 (N_9424,N_8278,N_8719);
xnor U9425 (N_9425,N_8120,N_8248);
xor U9426 (N_9426,N_8797,N_8705);
xnor U9427 (N_9427,N_8063,N_8333);
nor U9428 (N_9428,N_8399,N_8581);
xor U9429 (N_9429,N_8608,N_8515);
xor U9430 (N_9430,N_8421,N_8241);
or U9431 (N_9431,N_8270,N_8675);
nand U9432 (N_9432,N_8678,N_8752);
nand U9433 (N_9433,N_8303,N_8206);
or U9434 (N_9434,N_8655,N_8009);
and U9435 (N_9435,N_8437,N_8205);
xor U9436 (N_9436,N_8614,N_8682);
nand U9437 (N_9437,N_8258,N_8653);
and U9438 (N_9438,N_8494,N_8565);
nand U9439 (N_9439,N_8153,N_8541);
nand U9440 (N_9440,N_8175,N_8439);
and U9441 (N_9441,N_8070,N_8241);
and U9442 (N_9442,N_8770,N_8042);
and U9443 (N_9443,N_8484,N_8430);
xor U9444 (N_9444,N_8599,N_8411);
xor U9445 (N_9445,N_8327,N_8790);
or U9446 (N_9446,N_8046,N_8025);
and U9447 (N_9447,N_8111,N_8718);
nand U9448 (N_9448,N_8580,N_8404);
or U9449 (N_9449,N_8338,N_8202);
xnor U9450 (N_9450,N_8090,N_8752);
nor U9451 (N_9451,N_8262,N_8522);
xnor U9452 (N_9452,N_8419,N_8789);
nor U9453 (N_9453,N_8468,N_8245);
nand U9454 (N_9454,N_8450,N_8114);
xor U9455 (N_9455,N_8314,N_8371);
and U9456 (N_9456,N_8699,N_8706);
or U9457 (N_9457,N_8066,N_8727);
xnor U9458 (N_9458,N_8459,N_8171);
xor U9459 (N_9459,N_8137,N_8468);
nor U9460 (N_9460,N_8281,N_8390);
and U9461 (N_9461,N_8477,N_8606);
nor U9462 (N_9462,N_8214,N_8271);
or U9463 (N_9463,N_8246,N_8638);
and U9464 (N_9464,N_8280,N_8407);
and U9465 (N_9465,N_8447,N_8141);
or U9466 (N_9466,N_8070,N_8032);
nand U9467 (N_9467,N_8125,N_8504);
nand U9468 (N_9468,N_8389,N_8637);
nor U9469 (N_9469,N_8644,N_8204);
nor U9470 (N_9470,N_8709,N_8107);
nand U9471 (N_9471,N_8124,N_8650);
and U9472 (N_9472,N_8655,N_8379);
or U9473 (N_9473,N_8303,N_8669);
nand U9474 (N_9474,N_8681,N_8062);
nor U9475 (N_9475,N_8073,N_8481);
and U9476 (N_9476,N_8257,N_8536);
and U9477 (N_9477,N_8585,N_8418);
xnor U9478 (N_9478,N_8366,N_8489);
nor U9479 (N_9479,N_8067,N_8135);
nand U9480 (N_9480,N_8426,N_8798);
nor U9481 (N_9481,N_8132,N_8623);
nor U9482 (N_9482,N_8159,N_8711);
nor U9483 (N_9483,N_8176,N_8784);
or U9484 (N_9484,N_8392,N_8733);
xnor U9485 (N_9485,N_8550,N_8515);
xor U9486 (N_9486,N_8150,N_8793);
or U9487 (N_9487,N_8783,N_8192);
or U9488 (N_9488,N_8094,N_8689);
nor U9489 (N_9489,N_8098,N_8493);
xor U9490 (N_9490,N_8028,N_8091);
or U9491 (N_9491,N_8153,N_8406);
nor U9492 (N_9492,N_8428,N_8101);
nand U9493 (N_9493,N_8013,N_8587);
or U9494 (N_9494,N_8727,N_8212);
and U9495 (N_9495,N_8213,N_8419);
nand U9496 (N_9496,N_8592,N_8698);
nand U9497 (N_9497,N_8146,N_8626);
xor U9498 (N_9498,N_8283,N_8194);
and U9499 (N_9499,N_8415,N_8555);
xnor U9500 (N_9500,N_8048,N_8195);
nand U9501 (N_9501,N_8702,N_8576);
or U9502 (N_9502,N_8498,N_8675);
and U9503 (N_9503,N_8029,N_8534);
nand U9504 (N_9504,N_8646,N_8583);
and U9505 (N_9505,N_8336,N_8350);
nor U9506 (N_9506,N_8116,N_8680);
and U9507 (N_9507,N_8300,N_8374);
nor U9508 (N_9508,N_8085,N_8451);
or U9509 (N_9509,N_8232,N_8264);
or U9510 (N_9510,N_8440,N_8527);
nand U9511 (N_9511,N_8083,N_8639);
and U9512 (N_9512,N_8196,N_8471);
nand U9513 (N_9513,N_8282,N_8367);
nand U9514 (N_9514,N_8230,N_8799);
xor U9515 (N_9515,N_8123,N_8486);
and U9516 (N_9516,N_8188,N_8072);
or U9517 (N_9517,N_8348,N_8580);
or U9518 (N_9518,N_8359,N_8369);
nor U9519 (N_9519,N_8131,N_8502);
or U9520 (N_9520,N_8508,N_8795);
nor U9521 (N_9521,N_8564,N_8524);
or U9522 (N_9522,N_8254,N_8431);
or U9523 (N_9523,N_8195,N_8766);
nand U9524 (N_9524,N_8547,N_8061);
and U9525 (N_9525,N_8781,N_8798);
and U9526 (N_9526,N_8231,N_8337);
nor U9527 (N_9527,N_8278,N_8671);
nand U9528 (N_9528,N_8448,N_8477);
or U9529 (N_9529,N_8709,N_8170);
and U9530 (N_9530,N_8305,N_8133);
or U9531 (N_9531,N_8396,N_8341);
nand U9532 (N_9532,N_8101,N_8168);
nor U9533 (N_9533,N_8463,N_8411);
xor U9534 (N_9534,N_8235,N_8640);
xnor U9535 (N_9535,N_8681,N_8721);
nor U9536 (N_9536,N_8286,N_8426);
xnor U9537 (N_9537,N_8696,N_8332);
xor U9538 (N_9538,N_8395,N_8465);
nor U9539 (N_9539,N_8244,N_8659);
nand U9540 (N_9540,N_8142,N_8347);
xor U9541 (N_9541,N_8426,N_8147);
nor U9542 (N_9542,N_8641,N_8598);
nor U9543 (N_9543,N_8524,N_8077);
and U9544 (N_9544,N_8463,N_8586);
or U9545 (N_9545,N_8486,N_8769);
and U9546 (N_9546,N_8346,N_8164);
and U9547 (N_9547,N_8693,N_8327);
xnor U9548 (N_9548,N_8129,N_8522);
nor U9549 (N_9549,N_8341,N_8440);
nor U9550 (N_9550,N_8518,N_8240);
nand U9551 (N_9551,N_8232,N_8531);
and U9552 (N_9552,N_8374,N_8483);
xor U9553 (N_9553,N_8059,N_8558);
and U9554 (N_9554,N_8070,N_8739);
and U9555 (N_9555,N_8300,N_8458);
nor U9556 (N_9556,N_8444,N_8284);
xor U9557 (N_9557,N_8198,N_8400);
nor U9558 (N_9558,N_8345,N_8457);
nor U9559 (N_9559,N_8107,N_8240);
and U9560 (N_9560,N_8572,N_8379);
xnor U9561 (N_9561,N_8045,N_8332);
nand U9562 (N_9562,N_8021,N_8721);
nand U9563 (N_9563,N_8452,N_8546);
xor U9564 (N_9564,N_8538,N_8217);
xor U9565 (N_9565,N_8759,N_8118);
nor U9566 (N_9566,N_8224,N_8171);
xnor U9567 (N_9567,N_8750,N_8557);
nor U9568 (N_9568,N_8514,N_8132);
nor U9569 (N_9569,N_8588,N_8640);
xor U9570 (N_9570,N_8292,N_8761);
xnor U9571 (N_9571,N_8194,N_8337);
xnor U9572 (N_9572,N_8325,N_8076);
and U9573 (N_9573,N_8182,N_8519);
and U9574 (N_9574,N_8729,N_8701);
xor U9575 (N_9575,N_8158,N_8422);
xor U9576 (N_9576,N_8161,N_8648);
and U9577 (N_9577,N_8019,N_8266);
nand U9578 (N_9578,N_8386,N_8290);
or U9579 (N_9579,N_8602,N_8634);
nor U9580 (N_9580,N_8461,N_8390);
or U9581 (N_9581,N_8503,N_8025);
nor U9582 (N_9582,N_8579,N_8382);
or U9583 (N_9583,N_8098,N_8039);
nand U9584 (N_9584,N_8123,N_8326);
and U9585 (N_9585,N_8081,N_8397);
or U9586 (N_9586,N_8638,N_8586);
and U9587 (N_9587,N_8586,N_8147);
or U9588 (N_9588,N_8253,N_8298);
nor U9589 (N_9589,N_8342,N_8032);
nand U9590 (N_9590,N_8491,N_8681);
xnor U9591 (N_9591,N_8681,N_8203);
and U9592 (N_9592,N_8266,N_8248);
xnor U9593 (N_9593,N_8611,N_8755);
and U9594 (N_9594,N_8384,N_8389);
and U9595 (N_9595,N_8434,N_8335);
nor U9596 (N_9596,N_8698,N_8643);
nor U9597 (N_9597,N_8008,N_8401);
nand U9598 (N_9598,N_8475,N_8019);
and U9599 (N_9599,N_8365,N_8082);
nor U9600 (N_9600,N_9589,N_9582);
or U9601 (N_9601,N_9461,N_9519);
or U9602 (N_9602,N_8986,N_9206);
nand U9603 (N_9603,N_9306,N_9154);
nor U9604 (N_9604,N_9413,N_9246);
xor U9605 (N_9605,N_9277,N_9363);
xnor U9606 (N_9606,N_9553,N_9533);
and U9607 (N_9607,N_9076,N_8804);
nor U9608 (N_9608,N_8886,N_9019);
nand U9609 (N_9609,N_9479,N_9152);
xor U9610 (N_9610,N_9230,N_9010);
or U9611 (N_9611,N_9333,N_9531);
or U9612 (N_9612,N_9327,N_9437);
nand U9613 (N_9613,N_9569,N_9263);
and U9614 (N_9614,N_9298,N_9551);
nor U9615 (N_9615,N_9105,N_9383);
nand U9616 (N_9616,N_8803,N_9258);
nand U9617 (N_9617,N_9360,N_9501);
nor U9618 (N_9618,N_9460,N_9492);
xor U9619 (N_9619,N_9068,N_9332);
nand U9620 (N_9620,N_9245,N_8834);
or U9621 (N_9621,N_9336,N_8924);
nor U9622 (N_9622,N_9155,N_8955);
or U9623 (N_9623,N_9491,N_9381);
or U9624 (N_9624,N_9335,N_9186);
xnor U9625 (N_9625,N_8928,N_8968);
xor U9626 (N_9626,N_8808,N_9073);
and U9627 (N_9627,N_8809,N_9573);
nand U9628 (N_9628,N_9398,N_8855);
nor U9629 (N_9629,N_9495,N_8909);
nand U9630 (N_9630,N_9557,N_8853);
xor U9631 (N_9631,N_9188,N_9140);
xnor U9632 (N_9632,N_9564,N_9013);
and U9633 (N_9633,N_9240,N_9069);
nand U9634 (N_9634,N_9545,N_9421);
or U9635 (N_9635,N_9117,N_9474);
or U9636 (N_9636,N_9365,N_9144);
xnor U9637 (N_9637,N_9418,N_9414);
and U9638 (N_9638,N_9279,N_8841);
or U9639 (N_9639,N_9447,N_9425);
and U9640 (N_9640,N_8941,N_9256);
nand U9641 (N_9641,N_8917,N_9391);
xnor U9642 (N_9642,N_8813,N_8830);
nor U9643 (N_9643,N_9162,N_8817);
nor U9644 (N_9644,N_9172,N_9035);
and U9645 (N_9645,N_8980,N_9346);
nand U9646 (N_9646,N_9351,N_9149);
nand U9647 (N_9647,N_8812,N_9259);
xnor U9648 (N_9648,N_9348,N_9469);
nand U9649 (N_9649,N_9563,N_9176);
nor U9650 (N_9650,N_8829,N_9173);
or U9651 (N_9651,N_9185,N_9102);
or U9652 (N_9652,N_9012,N_9429);
xor U9653 (N_9653,N_8961,N_9135);
nor U9654 (N_9654,N_9020,N_8802);
and U9655 (N_9655,N_8871,N_9310);
nor U9656 (N_9656,N_9517,N_9254);
nand U9657 (N_9657,N_8800,N_8989);
nand U9658 (N_9658,N_9318,N_9093);
xnor U9659 (N_9659,N_9122,N_9187);
nor U9660 (N_9660,N_9527,N_9085);
xnor U9661 (N_9661,N_8907,N_9534);
nand U9662 (N_9662,N_8876,N_8940);
nor U9663 (N_9663,N_9544,N_9147);
nor U9664 (N_9664,N_8922,N_8805);
and U9665 (N_9665,N_9473,N_9134);
or U9666 (N_9666,N_9394,N_9316);
and U9667 (N_9667,N_9023,N_9520);
xnor U9668 (N_9668,N_9549,N_9404);
nor U9669 (N_9669,N_9378,N_9111);
and U9670 (N_9670,N_9079,N_8903);
nor U9671 (N_9671,N_8880,N_8807);
and U9672 (N_9672,N_8872,N_8934);
nand U9673 (N_9673,N_8822,N_9315);
nand U9674 (N_9674,N_9008,N_9065);
nand U9675 (N_9675,N_9281,N_9177);
or U9676 (N_9676,N_9107,N_9587);
and U9677 (N_9677,N_8947,N_9530);
or U9678 (N_9678,N_9060,N_9101);
and U9679 (N_9679,N_8927,N_9400);
nand U9680 (N_9680,N_8993,N_9294);
and U9681 (N_9681,N_9434,N_8966);
or U9682 (N_9682,N_9410,N_8981);
nand U9683 (N_9683,N_8930,N_9201);
xnor U9684 (N_9684,N_9312,N_9158);
nand U9685 (N_9685,N_9220,N_9320);
nor U9686 (N_9686,N_9537,N_9471);
nand U9687 (N_9687,N_9170,N_9067);
nand U9688 (N_9688,N_9248,N_9022);
xnor U9689 (N_9689,N_8965,N_9450);
and U9690 (N_9690,N_9299,N_9126);
xor U9691 (N_9691,N_9331,N_9499);
xnor U9692 (N_9692,N_8882,N_9132);
nor U9693 (N_9693,N_8828,N_8977);
and U9694 (N_9694,N_9130,N_9511);
and U9695 (N_9695,N_9039,N_9222);
or U9696 (N_9696,N_9243,N_9238);
or U9697 (N_9697,N_8923,N_9487);
or U9698 (N_9698,N_9124,N_9493);
xnor U9699 (N_9699,N_9242,N_8949);
nor U9700 (N_9700,N_9150,N_8982);
nor U9701 (N_9701,N_9114,N_9497);
or U9702 (N_9702,N_9225,N_9321);
xor U9703 (N_9703,N_9542,N_8908);
and U9704 (N_9704,N_9043,N_8819);
xnor U9705 (N_9705,N_9558,N_8956);
and U9706 (N_9706,N_9211,N_9146);
xnor U9707 (N_9707,N_9467,N_9007);
xnor U9708 (N_9708,N_9163,N_9326);
xor U9709 (N_9709,N_8849,N_9133);
nor U9710 (N_9710,N_9484,N_8978);
nor U9711 (N_9711,N_9000,N_8873);
nor U9712 (N_9712,N_9396,N_8942);
and U9713 (N_9713,N_9157,N_9044);
or U9714 (N_9714,N_9369,N_9156);
or U9715 (N_9715,N_9342,N_8862);
or U9716 (N_9716,N_8952,N_8999);
or U9717 (N_9717,N_8892,N_9417);
nand U9718 (N_9718,N_8996,N_9538);
nor U9719 (N_9719,N_9411,N_9016);
nor U9720 (N_9720,N_9349,N_9518);
and U9721 (N_9721,N_9585,N_9370);
and U9722 (N_9722,N_9374,N_9488);
nand U9723 (N_9723,N_9006,N_9141);
or U9724 (N_9724,N_8836,N_8905);
nor U9725 (N_9725,N_8953,N_9169);
and U9726 (N_9726,N_8843,N_8842);
or U9727 (N_9727,N_9325,N_8895);
or U9728 (N_9728,N_8902,N_8943);
or U9729 (N_9729,N_9462,N_9485);
or U9730 (N_9730,N_9232,N_9406);
nor U9731 (N_9731,N_9503,N_9208);
or U9732 (N_9732,N_9047,N_9057);
nor U9733 (N_9733,N_8840,N_9455);
xnor U9734 (N_9734,N_9030,N_9160);
xnor U9735 (N_9735,N_9388,N_9502);
nor U9736 (N_9736,N_9372,N_9449);
and U9737 (N_9737,N_9546,N_9366);
nand U9738 (N_9738,N_9489,N_8823);
nand U9739 (N_9739,N_9215,N_9061);
xor U9740 (N_9740,N_9226,N_8933);
or U9741 (N_9741,N_9109,N_8857);
nor U9742 (N_9742,N_9514,N_9203);
nor U9743 (N_9743,N_9081,N_9066);
and U9744 (N_9744,N_9344,N_9470);
nor U9745 (N_9745,N_9415,N_8850);
or U9746 (N_9746,N_8863,N_9056);
nor U9747 (N_9747,N_9078,N_9084);
nor U9748 (N_9748,N_9042,N_9422);
nand U9749 (N_9749,N_9382,N_9583);
or U9750 (N_9750,N_8814,N_8900);
nor U9751 (N_9751,N_9424,N_8833);
nand U9752 (N_9752,N_8811,N_8931);
and U9753 (N_9753,N_9265,N_9297);
or U9754 (N_9754,N_8854,N_9269);
and U9755 (N_9755,N_9392,N_9251);
nor U9756 (N_9756,N_9592,N_9459);
or U9757 (N_9757,N_9241,N_9174);
xor U9758 (N_9758,N_9548,N_9086);
nand U9759 (N_9759,N_9197,N_9011);
nor U9760 (N_9760,N_8988,N_9119);
or U9761 (N_9761,N_9302,N_9308);
and U9762 (N_9762,N_9090,N_9196);
nor U9763 (N_9763,N_9275,N_8998);
nor U9764 (N_9764,N_8869,N_9257);
or U9765 (N_9765,N_9322,N_9087);
nand U9766 (N_9766,N_9005,N_8839);
and U9767 (N_9767,N_8867,N_8979);
nor U9768 (N_9768,N_9500,N_8893);
nand U9769 (N_9769,N_9522,N_9218);
and U9770 (N_9770,N_9445,N_9034);
or U9771 (N_9771,N_9261,N_9182);
xor U9772 (N_9772,N_8910,N_8963);
or U9773 (N_9773,N_9266,N_9319);
or U9774 (N_9774,N_9041,N_9543);
nand U9775 (N_9775,N_8994,N_9062);
xor U9776 (N_9776,N_9282,N_8976);
nor U9777 (N_9777,N_9129,N_8920);
xnor U9778 (N_9778,N_9345,N_9561);
nand U9779 (N_9779,N_9362,N_9123);
and U9780 (N_9780,N_9192,N_9219);
nor U9781 (N_9781,N_9458,N_9283);
nand U9782 (N_9782,N_9376,N_9393);
and U9783 (N_9783,N_8815,N_9271);
and U9784 (N_9784,N_9287,N_9431);
nand U9785 (N_9785,N_9419,N_9390);
or U9786 (N_9786,N_9112,N_8865);
xnor U9787 (N_9787,N_9142,N_9599);
xnor U9788 (N_9788,N_9334,N_9405);
or U9789 (N_9789,N_9194,N_9356);
xnor U9790 (N_9790,N_9108,N_8847);
or U9791 (N_9791,N_9465,N_8946);
nor U9792 (N_9792,N_9032,N_9014);
and U9793 (N_9793,N_9286,N_9063);
xnor U9794 (N_9794,N_8883,N_9504);
nor U9795 (N_9795,N_9038,N_9236);
or U9796 (N_9796,N_9496,N_9466);
nand U9797 (N_9797,N_9324,N_8926);
nand U9798 (N_9798,N_9051,N_9195);
and U9799 (N_9799,N_9593,N_8974);
xnor U9800 (N_9800,N_8912,N_9436);
or U9801 (N_9801,N_9442,N_9359);
and U9802 (N_9802,N_9453,N_9053);
and U9803 (N_9803,N_9046,N_9494);
nand U9804 (N_9804,N_9480,N_8919);
xnor U9805 (N_9805,N_9200,N_9532);
nand U9806 (N_9806,N_9443,N_9024);
or U9807 (N_9807,N_9395,N_8856);
nand U9808 (N_9808,N_9357,N_9575);
or U9809 (N_9809,N_9552,N_9472);
nand U9810 (N_9810,N_9478,N_9584);
nor U9811 (N_9811,N_9205,N_9166);
and U9812 (N_9812,N_8820,N_8985);
nand U9813 (N_9813,N_9028,N_9171);
and U9814 (N_9814,N_8970,N_9054);
or U9815 (N_9815,N_9352,N_8827);
nand U9816 (N_9816,N_9403,N_9159);
and U9817 (N_9817,N_9165,N_9168);
nor U9818 (N_9818,N_9127,N_9052);
nor U9819 (N_9819,N_8935,N_9045);
nor U9820 (N_9820,N_9083,N_8983);
or U9821 (N_9821,N_9137,N_9164);
xnor U9822 (N_9822,N_9221,N_9482);
and U9823 (N_9823,N_9110,N_9244);
xnor U9824 (N_9824,N_8936,N_9379);
xor U9825 (N_9825,N_9516,N_9323);
nand U9826 (N_9826,N_9175,N_9387);
xnor U9827 (N_9827,N_9456,N_9089);
or U9828 (N_9828,N_8960,N_9037);
nand U9829 (N_9829,N_8916,N_9586);
and U9830 (N_9830,N_8860,N_8904);
and U9831 (N_9831,N_9209,N_9490);
or U9832 (N_9832,N_9399,N_9235);
xnor U9833 (N_9833,N_9512,N_9354);
xnor U9834 (N_9834,N_9339,N_8967);
or U9835 (N_9835,N_9441,N_8969);
xnor U9836 (N_9836,N_9596,N_9535);
xor U9837 (N_9837,N_9568,N_9343);
and U9838 (N_9838,N_9386,N_9289);
nand U9839 (N_9839,N_9595,N_9296);
and U9840 (N_9840,N_8868,N_9290);
or U9841 (N_9841,N_9317,N_8810);
and U9842 (N_9842,N_8997,N_9358);
and U9843 (N_9843,N_9598,N_9428);
nand U9844 (N_9844,N_9284,N_9181);
xor U9845 (N_9845,N_9247,N_9059);
and U9846 (N_9846,N_8816,N_9523);
nand U9847 (N_9847,N_9468,N_8929);
or U9848 (N_9848,N_8881,N_9204);
or U9849 (N_9849,N_9295,N_8959);
nand U9850 (N_9850,N_8896,N_9099);
or U9851 (N_9851,N_9113,N_8825);
and U9852 (N_9852,N_9092,N_9525);
nand U9853 (N_9853,N_9361,N_8937);
or U9854 (N_9854,N_9385,N_9260);
or U9855 (N_9855,N_9291,N_9590);
or U9856 (N_9856,N_9597,N_8915);
and U9857 (N_9857,N_9526,N_9179);
and U9858 (N_9858,N_8954,N_9539);
xnor U9859 (N_9859,N_9151,N_9064);
or U9860 (N_9860,N_8972,N_9444);
xnor U9861 (N_9861,N_9217,N_8887);
or U9862 (N_9862,N_8870,N_9375);
or U9863 (N_9863,N_9448,N_9216);
nor U9864 (N_9864,N_9180,N_9329);
xnor U9865 (N_9865,N_9104,N_9021);
xnor U9866 (N_9866,N_9412,N_8835);
nor U9867 (N_9867,N_9565,N_9049);
and U9868 (N_9868,N_9273,N_9353);
and U9869 (N_9869,N_9389,N_9075);
nand U9870 (N_9870,N_8925,N_9536);
nor U9871 (N_9871,N_9031,N_8991);
nand U9872 (N_9872,N_9193,N_9288);
or U9873 (N_9873,N_9148,N_8894);
nand U9874 (N_9874,N_9004,N_9074);
or U9875 (N_9875,N_8918,N_9212);
xnor U9876 (N_9876,N_9253,N_9380);
xnor U9877 (N_9877,N_8906,N_9070);
nor U9878 (N_9878,N_9566,N_9515);
or U9879 (N_9879,N_9433,N_9594);
and U9880 (N_9880,N_9371,N_9350);
and U9881 (N_9881,N_9427,N_9128);
nand U9882 (N_9882,N_8898,N_9293);
nor U9883 (N_9883,N_9178,N_9278);
nor U9884 (N_9884,N_8837,N_9311);
nand U9885 (N_9885,N_9255,N_9377);
and U9886 (N_9886,N_8866,N_9276);
xor U9887 (N_9887,N_9072,N_9285);
or U9888 (N_9888,N_8846,N_9303);
xnor U9889 (N_9889,N_9231,N_9040);
or U9890 (N_9890,N_9095,N_9314);
nor U9891 (N_9891,N_9097,N_8858);
xor U9892 (N_9892,N_9576,N_8879);
and U9893 (N_9893,N_8884,N_8897);
and U9894 (N_9894,N_9384,N_9264);
and U9895 (N_9895,N_9570,N_8848);
and U9896 (N_9896,N_8878,N_8806);
and U9897 (N_9897,N_8859,N_9483);
or U9898 (N_9898,N_9036,N_9001);
xnor U9899 (N_9899,N_9464,N_8832);
nand U9900 (N_9900,N_9588,N_9058);
nor U9901 (N_9901,N_9402,N_9125);
and U9902 (N_9902,N_9280,N_9373);
xor U9903 (N_9903,N_8888,N_9094);
or U9904 (N_9904,N_9096,N_8987);
nor U9905 (N_9905,N_9167,N_9228);
or U9906 (N_9906,N_9224,N_8864);
nand U9907 (N_9907,N_9138,N_8875);
or U9908 (N_9908,N_9183,N_9268);
or U9909 (N_9909,N_9591,N_9340);
nor U9910 (N_9910,N_9540,N_9541);
and U9911 (N_9911,N_9571,N_9432);
xnor U9912 (N_9912,N_8901,N_9025);
nor U9913 (N_9913,N_9304,N_8971);
xor U9914 (N_9914,N_9191,N_9446);
xnor U9915 (N_9915,N_9416,N_8831);
nand U9916 (N_9916,N_8995,N_8932);
nand U9917 (N_9917,N_9574,N_9420);
or U9918 (N_9918,N_8975,N_9559);
or U9919 (N_9919,N_9309,N_9524);
nand U9920 (N_9920,N_8914,N_8958);
xor U9921 (N_9921,N_9426,N_9567);
nand U9922 (N_9922,N_8990,N_9082);
nor U9923 (N_9923,N_9513,N_9015);
and U9924 (N_9924,N_8992,N_9003);
nor U9925 (N_9925,N_9161,N_9198);
and U9926 (N_9926,N_9477,N_9476);
nor U9927 (N_9927,N_9262,N_9547);
or U9928 (N_9928,N_9002,N_9026);
xor U9929 (N_9929,N_9009,N_9091);
xor U9930 (N_9930,N_8911,N_9439);
or U9931 (N_9931,N_9407,N_9213);
and U9932 (N_9932,N_8826,N_9475);
xnor U9933 (N_9933,N_8957,N_9267);
or U9934 (N_9934,N_9581,N_9550);
xor U9935 (N_9935,N_9199,N_9272);
nand U9936 (N_9936,N_9077,N_9292);
xor U9937 (N_9937,N_9307,N_9347);
nand U9938 (N_9938,N_9528,N_8818);
nor U9939 (N_9939,N_9027,N_9050);
nand U9940 (N_9940,N_9521,N_9397);
and U9941 (N_9941,N_8845,N_8944);
or U9942 (N_9942,N_9555,N_9184);
xor U9943 (N_9943,N_9202,N_9227);
or U9944 (N_9944,N_9438,N_9018);
nor U9945 (N_9945,N_8824,N_9457);
or U9946 (N_9946,N_9560,N_9145);
and U9947 (N_9947,N_8964,N_9223);
nand U9948 (N_9948,N_9017,N_8801);
and U9949 (N_9949,N_9029,N_9234);
or U9950 (N_9950,N_8821,N_8913);
and U9951 (N_9951,N_9252,N_9554);
nor U9952 (N_9952,N_9237,N_9100);
nand U9953 (N_9953,N_9507,N_8874);
nand U9954 (N_9954,N_9452,N_9409);
xor U9955 (N_9955,N_9368,N_9116);
nand U9956 (N_9956,N_9338,N_9328);
or U9957 (N_9957,N_8890,N_9423);
nand U9958 (N_9958,N_9250,N_9249);
or U9959 (N_9959,N_9098,N_9118);
or U9960 (N_9960,N_8984,N_9115);
xor U9961 (N_9961,N_9274,N_9556);
nor U9962 (N_9962,N_9033,N_9430);
or U9963 (N_9963,N_9153,N_8899);
nand U9964 (N_9964,N_9190,N_8844);
xor U9965 (N_9965,N_8938,N_9508);
nand U9966 (N_9966,N_9088,N_9454);
or U9967 (N_9967,N_8891,N_8962);
nor U9968 (N_9968,N_8889,N_9136);
xnor U9969 (N_9969,N_9498,N_9435);
nand U9970 (N_9970,N_9578,N_8851);
or U9971 (N_9971,N_9214,N_9330);
or U9972 (N_9972,N_9139,N_8973);
nand U9973 (N_9973,N_9579,N_8852);
or U9974 (N_9974,N_9055,N_8921);
nor U9975 (N_9975,N_9341,N_9120);
or U9976 (N_9976,N_9463,N_9486);
nor U9977 (N_9977,N_9239,N_9313);
nor U9978 (N_9978,N_9301,N_9131);
and U9979 (N_9979,N_9337,N_8950);
nand U9980 (N_9980,N_9080,N_8945);
nor U9981 (N_9981,N_8951,N_9481);
nand U9982 (N_9982,N_9506,N_8877);
xnor U9983 (N_9983,N_8939,N_9509);
nand U9984 (N_9984,N_9048,N_9121);
or U9985 (N_9985,N_9229,N_9562);
nand U9986 (N_9986,N_9510,N_9210);
xor U9987 (N_9987,N_9364,N_9401);
or U9988 (N_9988,N_9440,N_9103);
or U9989 (N_9989,N_9300,N_9505);
or U9990 (N_9990,N_9355,N_9071);
nor U9991 (N_9991,N_9367,N_9270);
nor U9992 (N_9992,N_9580,N_9529);
xor U9993 (N_9993,N_9143,N_9233);
nor U9994 (N_9994,N_9577,N_9451);
nand U9995 (N_9995,N_9305,N_9207);
or U9996 (N_9996,N_8838,N_8885);
or U9997 (N_9997,N_9572,N_8861);
nand U9998 (N_9998,N_9106,N_9189);
nor U9999 (N_9999,N_9408,N_8948);
and U10000 (N_10000,N_9308,N_9562);
or U10001 (N_10001,N_9407,N_9245);
nand U10002 (N_10002,N_8921,N_9521);
nand U10003 (N_10003,N_9158,N_9580);
nor U10004 (N_10004,N_9256,N_8985);
nor U10005 (N_10005,N_9254,N_9166);
or U10006 (N_10006,N_8858,N_9194);
nand U10007 (N_10007,N_9240,N_9322);
nor U10008 (N_10008,N_9353,N_9054);
xor U10009 (N_10009,N_8906,N_9186);
nand U10010 (N_10010,N_9206,N_9243);
or U10011 (N_10011,N_9055,N_9034);
or U10012 (N_10012,N_9508,N_8880);
xor U10013 (N_10013,N_9243,N_9256);
xor U10014 (N_10014,N_9171,N_8937);
nand U10015 (N_10015,N_9507,N_9248);
nor U10016 (N_10016,N_9199,N_9317);
and U10017 (N_10017,N_9350,N_9000);
nor U10018 (N_10018,N_8847,N_9574);
and U10019 (N_10019,N_8947,N_9405);
nor U10020 (N_10020,N_9063,N_9151);
nand U10021 (N_10021,N_9028,N_9137);
and U10022 (N_10022,N_8890,N_9346);
and U10023 (N_10023,N_9259,N_9204);
nand U10024 (N_10024,N_9541,N_8848);
nor U10025 (N_10025,N_9005,N_9188);
nand U10026 (N_10026,N_9366,N_9216);
xnor U10027 (N_10027,N_9328,N_9417);
and U10028 (N_10028,N_8988,N_9313);
nor U10029 (N_10029,N_8881,N_8848);
and U10030 (N_10030,N_9235,N_8876);
and U10031 (N_10031,N_9108,N_9352);
nand U10032 (N_10032,N_9106,N_9374);
or U10033 (N_10033,N_9005,N_8803);
nor U10034 (N_10034,N_8822,N_9526);
and U10035 (N_10035,N_9509,N_9137);
nor U10036 (N_10036,N_9164,N_9382);
and U10037 (N_10037,N_9212,N_9007);
or U10038 (N_10038,N_9502,N_8897);
or U10039 (N_10039,N_9391,N_9438);
nand U10040 (N_10040,N_9436,N_9141);
nand U10041 (N_10041,N_9330,N_8977);
and U10042 (N_10042,N_9170,N_9079);
nor U10043 (N_10043,N_9348,N_9122);
and U10044 (N_10044,N_9347,N_9361);
and U10045 (N_10045,N_9595,N_8992);
xnor U10046 (N_10046,N_9240,N_9436);
or U10047 (N_10047,N_9539,N_9259);
or U10048 (N_10048,N_9404,N_9197);
nand U10049 (N_10049,N_9142,N_8903);
or U10050 (N_10050,N_9080,N_9352);
xnor U10051 (N_10051,N_9013,N_8898);
or U10052 (N_10052,N_9142,N_9470);
xnor U10053 (N_10053,N_9295,N_9302);
and U10054 (N_10054,N_9539,N_9450);
xor U10055 (N_10055,N_9247,N_9149);
nor U10056 (N_10056,N_9107,N_8994);
or U10057 (N_10057,N_9032,N_9051);
xnor U10058 (N_10058,N_9463,N_8943);
or U10059 (N_10059,N_9570,N_9235);
or U10060 (N_10060,N_9316,N_9343);
and U10061 (N_10061,N_9468,N_9573);
and U10062 (N_10062,N_8828,N_9203);
nor U10063 (N_10063,N_9097,N_9557);
nand U10064 (N_10064,N_9494,N_9598);
or U10065 (N_10065,N_8865,N_9410);
xnor U10066 (N_10066,N_9508,N_9074);
or U10067 (N_10067,N_9430,N_9083);
and U10068 (N_10068,N_9148,N_9304);
or U10069 (N_10069,N_9408,N_9240);
and U10070 (N_10070,N_9381,N_9560);
xnor U10071 (N_10071,N_9077,N_9435);
and U10072 (N_10072,N_9313,N_9337);
nor U10073 (N_10073,N_9044,N_8985);
or U10074 (N_10074,N_8842,N_8900);
nor U10075 (N_10075,N_9452,N_9372);
nor U10076 (N_10076,N_9335,N_9092);
xnor U10077 (N_10077,N_9355,N_9507);
nor U10078 (N_10078,N_9010,N_9099);
nand U10079 (N_10079,N_9381,N_8921);
nor U10080 (N_10080,N_9069,N_8849);
nor U10081 (N_10081,N_9084,N_9055);
xor U10082 (N_10082,N_8920,N_9086);
nor U10083 (N_10083,N_9161,N_9394);
nor U10084 (N_10084,N_8969,N_9024);
nand U10085 (N_10085,N_8832,N_9072);
nor U10086 (N_10086,N_9536,N_8904);
and U10087 (N_10087,N_9325,N_9440);
and U10088 (N_10088,N_9488,N_9037);
and U10089 (N_10089,N_8882,N_9063);
xnor U10090 (N_10090,N_9552,N_9456);
nor U10091 (N_10091,N_9036,N_9383);
nand U10092 (N_10092,N_8953,N_9028);
nand U10093 (N_10093,N_9337,N_9392);
nand U10094 (N_10094,N_9124,N_9038);
or U10095 (N_10095,N_8968,N_9060);
nor U10096 (N_10096,N_9372,N_9116);
or U10097 (N_10097,N_8867,N_9171);
nand U10098 (N_10098,N_9284,N_9245);
nand U10099 (N_10099,N_8912,N_9456);
and U10100 (N_10100,N_8829,N_9331);
nor U10101 (N_10101,N_9284,N_9281);
and U10102 (N_10102,N_9578,N_9076);
nor U10103 (N_10103,N_9017,N_9539);
nor U10104 (N_10104,N_9039,N_8971);
and U10105 (N_10105,N_8912,N_9472);
xnor U10106 (N_10106,N_9205,N_9283);
or U10107 (N_10107,N_9135,N_8893);
or U10108 (N_10108,N_9166,N_9209);
and U10109 (N_10109,N_9570,N_9322);
nor U10110 (N_10110,N_8914,N_9358);
or U10111 (N_10111,N_8870,N_8895);
or U10112 (N_10112,N_8851,N_9469);
xnor U10113 (N_10113,N_9163,N_9298);
nor U10114 (N_10114,N_9390,N_9399);
nand U10115 (N_10115,N_8941,N_9421);
or U10116 (N_10116,N_9274,N_8929);
and U10117 (N_10117,N_9261,N_9204);
nand U10118 (N_10118,N_9014,N_8858);
nor U10119 (N_10119,N_9224,N_9126);
nor U10120 (N_10120,N_8869,N_9142);
and U10121 (N_10121,N_9564,N_9318);
xor U10122 (N_10122,N_9164,N_9522);
nor U10123 (N_10123,N_9503,N_8924);
nor U10124 (N_10124,N_9583,N_8860);
nand U10125 (N_10125,N_8840,N_9213);
or U10126 (N_10126,N_8976,N_9429);
and U10127 (N_10127,N_9264,N_9118);
and U10128 (N_10128,N_9445,N_9468);
nor U10129 (N_10129,N_9353,N_9328);
and U10130 (N_10130,N_8842,N_9199);
nor U10131 (N_10131,N_9334,N_9510);
nand U10132 (N_10132,N_9411,N_9558);
nand U10133 (N_10133,N_9556,N_9545);
xnor U10134 (N_10134,N_9416,N_9025);
xnor U10135 (N_10135,N_8996,N_9271);
nand U10136 (N_10136,N_9212,N_9018);
or U10137 (N_10137,N_9458,N_9092);
nand U10138 (N_10138,N_9492,N_9277);
xnor U10139 (N_10139,N_9102,N_9173);
nor U10140 (N_10140,N_8819,N_9064);
and U10141 (N_10141,N_9188,N_8950);
xor U10142 (N_10142,N_9467,N_9222);
and U10143 (N_10143,N_8826,N_9275);
or U10144 (N_10144,N_9163,N_9250);
xor U10145 (N_10145,N_9097,N_9284);
nor U10146 (N_10146,N_9297,N_9588);
xor U10147 (N_10147,N_9529,N_8939);
nor U10148 (N_10148,N_9524,N_9318);
or U10149 (N_10149,N_9026,N_9095);
nand U10150 (N_10150,N_9132,N_9272);
or U10151 (N_10151,N_8827,N_9298);
nor U10152 (N_10152,N_9341,N_9106);
or U10153 (N_10153,N_9245,N_9467);
nand U10154 (N_10154,N_9086,N_9027);
and U10155 (N_10155,N_9362,N_8818);
xor U10156 (N_10156,N_9486,N_9382);
xnor U10157 (N_10157,N_9196,N_9378);
nor U10158 (N_10158,N_9392,N_9076);
or U10159 (N_10159,N_8818,N_9155);
nand U10160 (N_10160,N_9335,N_9163);
nor U10161 (N_10161,N_9273,N_8883);
nand U10162 (N_10162,N_9383,N_9221);
and U10163 (N_10163,N_9081,N_9185);
or U10164 (N_10164,N_9000,N_9317);
or U10165 (N_10165,N_9269,N_9105);
nor U10166 (N_10166,N_8934,N_9441);
nand U10167 (N_10167,N_9111,N_9218);
or U10168 (N_10168,N_9463,N_9571);
nand U10169 (N_10169,N_8967,N_9120);
or U10170 (N_10170,N_8874,N_9144);
and U10171 (N_10171,N_9297,N_9548);
nand U10172 (N_10172,N_9025,N_8946);
and U10173 (N_10173,N_9481,N_9437);
xor U10174 (N_10174,N_9218,N_9470);
nand U10175 (N_10175,N_9216,N_9152);
xnor U10176 (N_10176,N_8906,N_8876);
nor U10177 (N_10177,N_8922,N_8822);
xor U10178 (N_10178,N_8951,N_9400);
nand U10179 (N_10179,N_9036,N_9509);
or U10180 (N_10180,N_9548,N_9598);
and U10181 (N_10181,N_9394,N_9510);
or U10182 (N_10182,N_9413,N_8899);
and U10183 (N_10183,N_9153,N_8818);
or U10184 (N_10184,N_9575,N_9554);
xor U10185 (N_10185,N_9533,N_9499);
and U10186 (N_10186,N_9477,N_9337);
or U10187 (N_10187,N_9445,N_9061);
or U10188 (N_10188,N_9196,N_9235);
and U10189 (N_10189,N_8834,N_8981);
nor U10190 (N_10190,N_9330,N_9303);
or U10191 (N_10191,N_9442,N_9258);
xor U10192 (N_10192,N_9257,N_9393);
and U10193 (N_10193,N_9071,N_9296);
nand U10194 (N_10194,N_9142,N_9314);
nor U10195 (N_10195,N_9216,N_9379);
or U10196 (N_10196,N_9477,N_9475);
or U10197 (N_10197,N_9130,N_8925);
and U10198 (N_10198,N_9106,N_9218);
xnor U10199 (N_10199,N_9157,N_8860);
nor U10200 (N_10200,N_8856,N_9302);
nand U10201 (N_10201,N_9498,N_8846);
xor U10202 (N_10202,N_9349,N_9220);
or U10203 (N_10203,N_9008,N_9578);
xnor U10204 (N_10204,N_8864,N_9015);
or U10205 (N_10205,N_9196,N_9178);
or U10206 (N_10206,N_9039,N_9570);
nor U10207 (N_10207,N_9558,N_9598);
nand U10208 (N_10208,N_9351,N_9171);
or U10209 (N_10209,N_8932,N_9441);
nor U10210 (N_10210,N_9438,N_9123);
or U10211 (N_10211,N_8850,N_9529);
or U10212 (N_10212,N_9486,N_8867);
nand U10213 (N_10213,N_9201,N_8875);
and U10214 (N_10214,N_9534,N_9045);
nand U10215 (N_10215,N_9155,N_8994);
or U10216 (N_10216,N_9037,N_9219);
nor U10217 (N_10217,N_9183,N_9057);
and U10218 (N_10218,N_8829,N_9024);
xnor U10219 (N_10219,N_9598,N_9173);
nand U10220 (N_10220,N_9395,N_9075);
or U10221 (N_10221,N_9563,N_9251);
and U10222 (N_10222,N_8947,N_9456);
nor U10223 (N_10223,N_9315,N_9124);
xor U10224 (N_10224,N_9298,N_8959);
and U10225 (N_10225,N_9593,N_9216);
xor U10226 (N_10226,N_9355,N_9156);
xor U10227 (N_10227,N_9211,N_8964);
and U10228 (N_10228,N_8864,N_8969);
nand U10229 (N_10229,N_9356,N_9223);
or U10230 (N_10230,N_9504,N_9457);
or U10231 (N_10231,N_9196,N_8979);
nand U10232 (N_10232,N_9138,N_9518);
or U10233 (N_10233,N_9529,N_8819);
and U10234 (N_10234,N_9101,N_9397);
nand U10235 (N_10235,N_8846,N_9132);
nor U10236 (N_10236,N_9567,N_9333);
nor U10237 (N_10237,N_8967,N_9031);
and U10238 (N_10238,N_9039,N_9057);
xor U10239 (N_10239,N_8947,N_9292);
nor U10240 (N_10240,N_9391,N_9277);
nor U10241 (N_10241,N_9127,N_9455);
or U10242 (N_10242,N_9420,N_8818);
xnor U10243 (N_10243,N_9286,N_9204);
and U10244 (N_10244,N_9256,N_9585);
or U10245 (N_10245,N_9300,N_9374);
nor U10246 (N_10246,N_9522,N_8918);
nor U10247 (N_10247,N_8814,N_9452);
nand U10248 (N_10248,N_8821,N_9361);
nand U10249 (N_10249,N_9236,N_8867);
xor U10250 (N_10250,N_8831,N_9172);
xor U10251 (N_10251,N_9561,N_9137);
nor U10252 (N_10252,N_9262,N_8908);
xnor U10253 (N_10253,N_9049,N_9076);
xor U10254 (N_10254,N_8842,N_9009);
xnor U10255 (N_10255,N_9136,N_8862);
xor U10256 (N_10256,N_9346,N_9549);
and U10257 (N_10257,N_8935,N_8917);
and U10258 (N_10258,N_9559,N_9265);
xnor U10259 (N_10259,N_9580,N_8986);
or U10260 (N_10260,N_9508,N_9144);
xor U10261 (N_10261,N_9186,N_8843);
nand U10262 (N_10262,N_8863,N_8962);
nor U10263 (N_10263,N_9357,N_9316);
and U10264 (N_10264,N_8845,N_9565);
nand U10265 (N_10265,N_9486,N_9395);
nand U10266 (N_10266,N_9396,N_8958);
nand U10267 (N_10267,N_9172,N_8810);
and U10268 (N_10268,N_9340,N_9070);
xnor U10269 (N_10269,N_9042,N_9163);
and U10270 (N_10270,N_8999,N_9465);
xor U10271 (N_10271,N_8966,N_9219);
or U10272 (N_10272,N_9288,N_9155);
and U10273 (N_10273,N_8824,N_9565);
nand U10274 (N_10274,N_9589,N_9244);
xor U10275 (N_10275,N_9018,N_8808);
and U10276 (N_10276,N_9225,N_9358);
nand U10277 (N_10277,N_9563,N_9136);
nor U10278 (N_10278,N_9219,N_9389);
or U10279 (N_10279,N_9591,N_9557);
nand U10280 (N_10280,N_9120,N_9593);
or U10281 (N_10281,N_9028,N_8919);
nor U10282 (N_10282,N_9509,N_9460);
xor U10283 (N_10283,N_9565,N_9108);
nor U10284 (N_10284,N_8850,N_8915);
or U10285 (N_10285,N_9125,N_9193);
or U10286 (N_10286,N_9426,N_9541);
nor U10287 (N_10287,N_9031,N_9035);
nor U10288 (N_10288,N_9489,N_8834);
nand U10289 (N_10289,N_9080,N_9211);
xor U10290 (N_10290,N_9520,N_8858);
nand U10291 (N_10291,N_8961,N_9302);
nand U10292 (N_10292,N_9384,N_9519);
nand U10293 (N_10293,N_8873,N_9008);
and U10294 (N_10294,N_9228,N_8930);
or U10295 (N_10295,N_9101,N_8903);
and U10296 (N_10296,N_8941,N_9118);
nand U10297 (N_10297,N_8927,N_9019);
nand U10298 (N_10298,N_9253,N_8902);
nand U10299 (N_10299,N_9309,N_9487);
or U10300 (N_10300,N_9036,N_9124);
and U10301 (N_10301,N_9193,N_9200);
or U10302 (N_10302,N_9345,N_9504);
or U10303 (N_10303,N_9260,N_9498);
xor U10304 (N_10304,N_8837,N_9053);
or U10305 (N_10305,N_9591,N_9255);
nor U10306 (N_10306,N_9342,N_9005);
and U10307 (N_10307,N_9052,N_9368);
and U10308 (N_10308,N_9519,N_8874);
and U10309 (N_10309,N_9519,N_8947);
nor U10310 (N_10310,N_9587,N_9300);
nor U10311 (N_10311,N_9584,N_9225);
or U10312 (N_10312,N_9344,N_9453);
or U10313 (N_10313,N_9105,N_9454);
and U10314 (N_10314,N_9026,N_9190);
and U10315 (N_10315,N_9253,N_9249);
xnor U10316 (N_10316,N_9487,N_9288);
xnor U10317 (N_10317,N_8913,N_9244);
and U10318 (N_10318,N_9477,N_9307);
xor U10319 (N_10319,N_9184,N_9094);
nand U10320 (N_10320,N_9370,N_9492);
and U10321 (N_10321,N_9301,N_9339);
or U10322 (N_10322,N_9414,N_9375);
or U10323 (N_10323,N_9310,N_9462);
nor U10324 (N_10324,N_8870,N_9545);
and U10325 (N_10325,N_9268,N_8855);
xnor U10326 (N_10326,N_9542,N_9585);
nor U10327 (N_10327,N_9074,N_9344);
xor U10328 (N_10328,N_9155,N_8910);
nand U10329 (N_10329,N_9590,N_9247);
or U10330 (N_10330,N_8950,N_8822);
xor U10331 (N_10331,N_9472,N_9378);
nand U10332 (N_10332,N_9019,N_9453);
nand U10333 (N_10333,N_9537,N_8918);
nor U10334 (N_10334,N_9514,N_9475);
nor U10335 (N_10335,N_9245,N_9019);
nor U10336 (N_10336,N_8860,N_9160);
and U10337 (N_10337,N_9208,N_9390);
nor U10338 (N_10338,N_9584,N_8939);
nor U10339 (N_10339,N_9403,N_9489);
xnor U10340 (N_10340,N_8986,N_9592);
nand U10341 (N_10341,N_9068,N_9438);
and U10342 (N_10342,N_8884,N_9312);
nand U10343 (N_10343,N_9341,N_9220);
xor U10344 (N_10344,N_9505,N_9024);
and U10345 (N_10345,N_9490,N_9308);
nand U10346 (N_10346,N_9255,N_8811);
nor U10347 (N_10347,N_9517,N_8891);
nor U10348 (N_10348,N_9446,N_9562);
or U10349 (N_10349,N_9552,N_9256);
xor U10350 (N_10350,N_8825,N_8879);
nor U10351 (N_10351,N_9089,N_9405);
and U10352 (N_10352,N_9524,N_9020);
and U10353 (N_10353,N_8803,N_9219);
or U10354 (N_10354,N_9263,N_9218);
xor U10355 (N_10355,N_9294,N_9228);
xnor U10356 (N_10356,N_9536,N_8801);
xnor U10357 (N_10357,N_8849,N_8977);
xor U10358 (N_10358,N_9420,N_9327);
or U10359 (N_10359,N_9218,N_9386);
and U10360 (N_10360,N_8933,N_9150);
xnor U10361 (N_10361,N_8943,N_9281);
xnor U10362 (N_10362,N_9528,N_9246);
nand U10363 (N_10363,N_8894,N_9120);
nor U10364 (N_10364,N_9250,N_9380);
nor U10365 (N_10365,N_8922,N_8963);
and U10366 (N_10366,N_9085,N_9549);
nand U10367 (N_10367,N_9185,N_9321);
and U10368 (N_10368,N_9481,N_9519);
nor U10369 (N_10369,N_8937,N_9209);
nand U10370 (N_10370,N_9039,N_9162);
nor U10371 (N_10371,N_9467,N_9451);
xor U10372 (N_10372,N_9486,N_9358);
or U10373 (N_10373,N_8839,N_9048);
and U10374 (N_10374,N_9200,N_8998);
nand U10375 (N_10375,N_8820,N_8819);
nand U10376 (N_10376,N_8874,N_9490);
nor U10377 (N_10377,N_9490,N_8950);
or U10378 (N_10378,N_9307,N_9438);
xnor U10379 (N_10379,N_8848,N_9174);
nor U10380 (N_10380,N_9327,N_8926);
or U10381 (N_10381,N_9484,N_9487);
xnor U10382 (N_10382,N_8817,N_9204);
or U10383 (N_10383,N_8862,N_9517);
nor U10384 (N_10384,N_8958,N_9530);
or U10385 (N_10385,N_9309,N_8808);
and U10386 (N_10386,N_9128,N_8910);
nand U10387 (N_10387,N_8881,N_8915);
or U10388 (N_10388,N_9508,N_9479);
and U10389 (N_10389,N_9315,N_9049);
nand U10390 (N_10390,N_9567,N_8905);
nand U10391 (N_10391,N_9355,N_8805);
xnor U10392 (N_10392,N_9426,N_9241);
or U10393 (N_10393,N_9413,N_9301);
and U10394 (N_10394,N_9110,N_9512);
nor U10395 (N_10395,N_9535,N_9159);
and U10396 (N_10396,N_9240,N_8895);
xnor U10397 (N_10397,N_9182,N_9125);
nor U10398 (N_10398,N_9590,N_9120);
or U10399 (N_10399,N_9210,N_8858);
nor U10400 (N_10400,N_9822,N_9992);
xnor U10401 (N_10401,N_10156,N_10118);
nand U10402 (N_10402,N_9856,N_10099);
xnor U10403 (N_10403,N_10271,N_9929);
or U10404 (N_10404,N_9854,N_10061);
or U10405 (N_10405,N_10382,N_10034);
nand U10406 (N_10406,N_9804,N_9741);
xor U10407 (N_10407,N_10067,N_10303);
nand U10408 (N_10408,N_10184,N_10028);
xor U10409 (N_10409,N_9794,N_10104);
nand U10410 (N_10410,N_10189,N_9987);
or U10411 (N_10411,N_10277,N_10022);
nand U10412 (N_10412,N_10254,N_9682);
or U10413 (N_10413,N_10379,N_9905);
or U10414 (N_10414,N_10332,N_9899);
xor U10415 (N_10415,N_10179,N_9893);
or U10416 (N_10416,N_9684,N_10057);
nand U10417 (N_10417,N_10210,N_9766);
and U10418 (N_10418,N_10205,N_9633);
nand U10419 (N_10419,N_9808,N_9732);
xor U10420 (N_10420,N_10053,N_9765);
xnor U10421 (N_10421,N_9832,N_10371);
nor U10422 (N_10422,N_9887,N_10339);
and U10423 (N_10423,N_9977,N_9750);
nor U10424 (N_10424,N_10321,N_10195);
xor U10425 (N_10425,N_9613,N_9703);
nor U10426 (N_10426,N_9874,N_10030);
and U10427 (N_10427,N_10134,N_9920);
and U10428 (N_10428,N_9939,N_10250);
or U10429 (N_10429,N_10161,N_9664);
xor U10430 (N_10430,N_10244,N_9890);
nand U10431 (N_10431,N_10115,N_9966);
nor U10432 (N_10432,N_10069,N_10304);
nor U10433 (N_10433,N_9911,N_10108);
nand U10434 (N_10434,N_10079,N_10336);
and U10435 (N_10435,N_9803,N_9923);
nor U10436 (N_10436,N_9877,N_9857);
xor U10437 (N_10437,N_10138,N_9967);
xnor U10438 (N_10438,N_9697,N_9937);
xor U10439 (N_10439,N_9642,N_10007);
and U10440 (N_10440,N_9875,N_10102);
and U10441 (N_10441,N_10142,N_9747);
nand U10442 (N_10442,N_9894,N_9736);
or U10443 (N_10443,N_10077,N_9756);
xor U10444 (N_10444,N_9666,N_10005);
and U10445 (N_10445,N_10261,N_9673);
xor U10446 (N_10446,N_10284,N_9849);
and U10447 (N_10447,N_10259,N_9835);
nor U10448 (N_10448,N_10206,N_9689);
and U10449 (N_10449,N_10176,N_9652);
xnor U10450 (N_10450,N_10119,N_9897);
nor U10451 (N_10451,N_9848,N_9885);
nor U10452 (N_10452,N_10380,N_10245);
xnor U10453 (N_10453,N_9882,N_9758);
or U10454 (N_10454,N_10025,N_10145);
xor U10455 (N_10455,N_9649,N_10194);
nand U10456 (N_10456,N_10268,N_10357);
or U10457 (N_10457,N_10154,N_10133);
nor U10458 (N_10458,N_10144,N_10222);
and U10459 (N_10459,N_9918,N_9783);
or U10460 (N_10460,N_9815,N_10363);
or U10461 (N_10461,N_10399,N_9843);
and U10462 (N_10462,N_10130,N_10175);
and U10463 (N_10463,N_9974,N_9944);
and U10464 (N_10464,N_10152,N_10021);
or U10465 (N_10465,N_10188,N_10225);
xnor U10466 (N_10466,N_9996,N_9910);
xor U10467 (N_10467,N_10101,N_10345);
and U10468 (N_10468,N_9692,N_9662);
or U10469 (N_10469,N_10330,N_9892);
and U10470 (N_10470,N_9779,N_9913);
nor U10471 (N_10471,N_9611,N_10314);
nor U10472 (N_10472,N_9947,N_10275);
nor U10473 (N_10473,N_10163,N_9799);
nor U10474 (N_10474,N_10049,N_9871);
or U10475 (N_10475,N_10198,N_10323);
or U10476 (N_10476,N_9813,N_10112);
and U10477 (N_10477,N_10094,N_9789);
or U10478 (N_10478,N_9809,N_9713);
or U10479 (N_10479,N_9755,N_9694);
xor U10480 (N_10480,N_9986,N_9615);
and U10481 (N_10481,N_9601,N_9771);
and U10482 (N_10482,N_9704,N_10217);
nor U10483 (N_10483,N_10389,N_9970);
nor U10484 (N_10484,N_10238,N_9745);
or U10485 (N_10485,N_9731,N_9791);
xnor U10486 (N_10486,N_9686,N_9888);
or U10487 (N_10487,N_9717,N_9961);
xnor U10488 (N_10488,N_10291,N_10174);
nand U10489 (N_10489,N_10033,N_9817);
nand U10490 (N_10490,N_10147,N_9988);
nor U10491 (N_10491,N_10209,N_9705);
or U10492 (N_10492,N_10383,N_9814);
or U10493 (N_10493,N_10372,N_10158);
and U10494 (N_10494,N_9952,N_9979);
or U10495 (N_10495,N_10249,N_9839);
nor U10496 (N_10496,N_10204,N_9626);
xor U10497 (N_10497,N_9614,N_10087);
nor U10498 (N_10498,N_9780,N_10299);
or U10499 (N_10499,N_9716,N_10137);
nor U10500 (N_10500,N_10279,N_9786);
nor U10501 (N_10501,N_10159,N_10351);
and U10502 (N_10502,N_9619,N_9735);
or U10503 (N_10503,N_10263,N_10095);
and U10504 (N_10504,N_10125,N_9776);
or U10505 (N_10505,N_10286,N_10241);
nor U10506 (N_10506,N_10050,N_9826);
xnor U10507 (N_10507,N_9990,N_10026);
nand U10508 (N_10508,N_10006,N_10121);
or U10509 (N_10509,N_10364,N_9862);
or U10510 (N_10510,N_9721,N_9927);
or U10511 (N_10511,N_9869,N_9847);
and U10512 (N_10512,N_10038,N_10126);
xor U10513 (N_10513,N_9612,N_9775);
or U10514 (N_10514,N_9678,N_10269);
nand U10515 (N_10515,N_9914,N_10221);
nand U10516 (N_10516,N_9685,N_10172);
and U10517 (N_10517,N_10207,N_10098);
nor U10518 (N_10518,N_10350,N_10103);
or U10519 (N_10519,N_10185,N_9973);
nor U10520 (N_10520,N_9650,N_10008);
or U10521 (N_10521,N_9878,N_10012);
xnor U10522 (N_10522,N_9951,N_9753);
xor U10523 (N_10523,N_9715,N_10211);
xnor U10524 (N_10524,N_9651,N_9998);
nor U10525 (N_10525,N_10000,N_10085);
xnor U10526 (N_10526,N_10362,N_10074);
nand U10527 (N_10527,N_9722,N_9930);
nand U10528 (N_10528,N_9621,N_10310);
and U10529 (N_10529,N_9940,N_10354);
nor U10530 (N_10530,N_10231,N_10242);
nor U10531 (N_10531,N_9931,N_9773);
xnor U10532 (N_10532,N_9896,N_10122);
nor U10533 (N_10533,N_9859,N_10015);
nand U10534 (N_10534,N_9883,N_10219);
nand U10535 (N_10535,N_10088,N_10208);
or U10536 (N_10536,N_9668,N_9953);
and U10537 (N_10537,N_10042,N_9846);
xor U10538 (N_10538,N_9639,N_9797);
and U10539 (N_10539,N_10212,N_9932);
and U10540 (N_10540,N_9955,N_9627);
xnor U10541 (N_10541,N_9810,N_9657);
or U10542 (N_10542,N_10044,N_9754);
xor U10543 (N_10543,N_10325,N_10100);
or U10544 (N_10544,N_10046,N_10388);
or U10545 (N_10545,N_9984,N_9618);
and U10546 (N_10546,N_9831,N_9669);
xnor U10547 (N_10547,N_9707,N_10181);
xnor U10548 (N_10548,N_10300,N_10341);
nand U10549 (N_10549,N_9793,N_9942);
or U10550 (N_10550,N_9807,N_9980);
or U10551 (N_10551,N_9768,N_10153);
xnor U10552 (N_10552,N_10218,N_10386);
or U10553 (N_10553,N_9820,N_10045);
nor U10554 (N_10554,N_10297,N_10216);
or U10555 (N_10555,N_9746,N_9683);
or U10556 (N_10556,N_10398,N_10047);
nor U10557 (N_10557,N_10131,N_9891);
nor U10558 (N_10558,N_10281,N_9687);
or U10559 (N_10559,N_9603,N_9946);
or U10560 (N_10560,N_9965,N_9935);
xor U10561 (N_10561,N_10213,N_10240);
and U10562 (N_10562,N_10369,N_10165);
or U10563 (N_10563,N_9616,N_10318);
and U10564 (N_10564,N_10397,N_9863);
nand U10565 (N_10565,N_9895,N_9976);
or U10566 (N_10566,N_9907,N_10064);
nand U10567 (N_10567,N_10252,N_10287);
nand U10568 (N_10568,N_10083,N_9838);
and U10569 (N_10569,N_10089,N_9861);
nand U10570 (N_10570,N_10150,N_9739);
nand U10571 (N_10571,N_10296,N_10019);
xnor U10572 (N_10572,N_9749,N_9926);
and U10573 (N_10573,N_9792,N_9962);
or U10574 (N_10574,N_10348,N_9969);
xnor U10575 (N_10575,N_10331,N_9880);
or U10576 (N_10576,N_10258,N_9909);
nor U10577 (N_10577,N_10171,N_9643);
or U10578 (N_10578,N_10109,N_10023);
nand U10579 (N_10579,N_10234,N_10264);
and U10580 (N_10580,N_10370,N_10017);
or U10581 (N_10581,N_10136,N_10378);
xor U10582 (N_10582,N_10352,N_9759);
nand U10583 (N_10583,N_9624,N_10197);
and U10584 (N_10584,N_10002,N_10305);
or U10585 (N_10585,N_9901,N_10235);
nor U10586 (N_10586,N_10114,N_9855);
nand U10587 (N_10587,N_9638,N_10020);
and U10588 (N_10588,N_10368,N_10313);
xnor U10589 (N_10589,N_9630,N_10190);
or U10590 (N_10590,N_9879,N_9681);
nor U10591 (N_10591,N_10322,N_10040);
and U10592 (N_10592,N_10200,N_10082);
nor U10593 (N_10593,N_9660,N_10255);
xor U10594 (N_10594,N_9900,N_10066);
and U10595 (N_10595,N_9702,N_9873);
nand U10596 (N_10596,N_10312,N_10290);
nand U10597 (N_10597,N_10366,N_9641);
xor U10598 (N_10598,N_9622,N_10186);
nor U10599 (N_10599,N_10288,N_10282);
xor U10600 (N_10600,N_10315,N_10157);
and U10601 (N_10601,N_10056,N_9665);
or U10602 (N_10602,N_10306,N_10024);
nor U10603 (N_10603,N_9729,N_9605);
or U10604 (N_10604,N_9726,N_10004);
nand U10605 (N_10605,N_9881,N_10373);
and U10606 (N_10606,N_9632,N_10319);
xnor U10607 (N_10607,N_9671,N_10349);
nor U10608 (N_10608,N_9740,N_10224);
nand U10609 (N_10609,N_10078,N_9680);
nor U10610 (N_10610,N_9975,N_9908);
xor U10611 (N_10611,N_10143,N_9928);
or U10612 (N_10612,N_10013,N_9700);
xor U10613 (N_10613,N_10276,N_9698);
or U10614 (N_10614,N_10182,N_10072);
nand U10615 (N_10615,N_9860,N_10355);
or U10616 (N_10616,N_10274,N_10301);
and U10617 (N_10617,N_9656,N_9868);
nor U10618 (N_10618,N_10298,N_10183);
and U10619 (N_10619,N_9872,N_10228);
and U10620 (N_10620,N_10317,N_9954);
xor U10621 (N_10621,N_9634,N_9654);
or U10622 (N_10622,N_10062,N_10346);
nor U10623 (N_10623,N_10324,N_9763);
nor U10624 (N_10624,N_9922,N_10251);
or U10625 (N_10625,N_10164,N_9635);
or U10626 (N_10626,N_10141,N_9798);
xor U10627 (N_10627,N_10039,N_10215);
and U10628 (N_10628,N_9950,N_10302);
xor U10629 (N_10629,N_9864,N_9915);
xnor U10630 (N_10630,N_9772,N_9600);
and U10631 (N_10631,N_10266,N_10229);
and U10632 (N_10632,N_9806,N_10036);
nand U10633 (N_10633,N_10246,N_9934);
nor U10634 (N_10634,N_10051,N_10376);
nor U10635 (N_10635,N_10337,N_9695);
nor U10636 (N_10636,N_10377,N_10365);
nor U10637 (N_10637,N_10237,N_9606);
and U10638 (N_10638,N_10168,N_10123);
or U10639 (N_10639,N_10292,N_9706);
nand U10640 (N_10640,N_10148,N_9784);
xnor U10641 (N_10641,N_10395,N_10105);
nor U10642 (N_10642,N_9711,N_10226);
nor U10643 (N_10643,N_10359,N_9658);
and U10644 (N_10644,N_9824,N_10311);
or U10645 (N_10645,N_9995,N_10361);
or U10646 (N_10646,N_10333,N_10392);
nand U10647 (N_10647,N_9821,N_9674);
nor U10648 (N_10648,N_9938,N_9767);
and U10649 (N_10649,N_9982,N_9699);
and U10650 (N_10650,N_9933,N_9949);
nor U10651 (N_10651,N_9663,N_9919);
xor U10652 (N_10652,N_9744,N_9870);
and U10653 (N_10653,N_9943,N_10054);
or U10654 (N_10654,N_10080,N_10178);
xor U10655 (N_10655,N_9675,N_9941);
and U10656 (N_10656,N_10316,N_10353);
nor U10657 (N_10657,N_10272,N_10092);
or U10658 (N_10658,N_9620,N_10041);
and U10659 (N_10659,N_9790,N_10360);
and U10660 (N_10660,N_9655,N_9964);
and U10661 (N_10661,N_9748,N_10031);
nand U10662 (N_10662,N_10139,N_9774);
nor U10663 (N_10663,N_10214,N_9866);
or U10664 (N_10664,N_10107,N_10110);
and U10665 (N_10665,N_10055,N_9963);
and U10666 (N_10666,N_10169,N_10257);
and U10667 (N_10667,N_9836,N_9972);
xor U10668 (N_10668,N_9802,N_9898);
nor U10669 (N_10669,N_9852,N_10384);
and U10670 (N_10670,N_10394,N_9644);
nor U10671 (N_10671,N_10070,N_9936);
nand U10672 (N_10672,N_9723,N_10124);
nor U10673 (N_10673,N_9743,N_10280);
nor U10674 (N_10674,N_9762,N_9924);
or U10675 (N_10675,N_9751,N_9827);
nor U10676 (N_10676,N_10071,N_9690);
xnor U10677 (N_10677,N_10199,N_9609);
nor U10678 (N_10678,N_10278,N_10018);
or U10679 (N_10679,N_9787,N_9837);
or U10680 (N_10680,N_9805,N_9728);
xor U10681 (N_10681,N_9983,N_9816);
and U10682 (N_10682,N_10106,N_10191);
or U10683 (N_10683,N_9710,N_9727);
nor U10684 (N_10684,N_10043,N_10326);
and U10685 (N_10685,N_9989,N_9948);
or U10686 (N_10686,N_10253,N_9959);
xnor U10687 (N_10687,N_10196,N_9997);
and U10688 (N_10688,N_9628,N_10073);
or U10689 (N_10689,N_10283,N_9737);
or U10690 (N_10690,N_9676,N_9916);
nand U10691 (N_10691,N_9709,N_9757);
xor U10692 (N_10692,N_9853,N_9752);
nand U10693 (N_10693,N_10170,N_9818);
and U10694 (N_10694,N_10132,N_10256);
xnor U10695 (N_10695,N_10097,N_10381);
or U10696 (N_10696,N_9667,N_9602);
nand U10697 (N_10697,N_9886,N_9812);
and U10698 (N_10698,N_10247,N_10334);
nor U10699 (N_10699,N_9917,N_10009);
nor U10700 (N_10700,N_10265,N_9801);
or U10701 (N_10701,N_9829,N_10390);
and U10702 (N_10702,N_9617,N_9708);
or U10703 (N_10703,N_10135,N_10374);
and U10704 (N_10704,N_10270,N_10032);
xnor U10705 (N_10705,N_9670,N_10236);
nand U10706 (N_10706,N_9677,N_9884);
xor U10707 (N_10707,N_10293,N_10329);
nand U10708 (N_10708,N_10010,N_9777);
xor U10709 (N_10709,N_10289,N_10308);
nand U10710 (N_10710,N_10093,N_10267);
or U10711 (N_10711,N_9828,N_10220);
and U10712 (N_10712,N_10151,N_9957);
and U10713 (N_10713,N_9844,N_10385);
nor U10714 (N_10714,N_10192,N_10187);
nand U10715 (N_10715,N_10285,N_10003);
nand U10716 (N_10716,N_10243,N_9653);
nor U10717 (N_10717,N_9921,N_10037);
and U10718 (N_10718,N_9991,N_10375);
or U10719 (N_10719,N_10052,N_9978);
xnor U10720 (N_10720,N_10091,N_10035);
xnor U10721 (N_10721,N_9925,N_9867);
xor U10722 (N_10722,N_10233,N_9714);
and U10723 (N_10723,N_10140,N_10011);
and U10724 (N_10724,N_9718,N_10180);
or U10725 (N_10725,N_9640,N_9720);
nand U10726 (N_10726,N_9858,N_9823);
nor U10727 (N_10727,N_9761,N_9819);
and U10728 (N_10728,N_10117,N_9811);
nand U10729 (N_10729,N_10120,N_10065);
and U10730 (N_10730,N_10167,N_10127);
and U10731 (N_10731,N_9696,N_9971);
xor U10732 (N_10732,N_10129,N_9834);
or U10733 (N_10733,N_9958,N_9945);
or U10734 (N_10734,N_9993,N_10162);
xor U10735 (N_10735,N_10393,N_9769);
or U10736 (N_10736,N_9785,N_9770);
nor U10737 (N_10737,N_9841,N_10166);
or U10738 (N_10738,N_10347,N_10328);
and U10739 (N_10739,N_9742,N_10248);
or U10740 (N_10740,N_10223,N_9672);
xnor U10741 (N_10741,N_10232,N_10128);
xor U10742 (N_10742,N_10340,N_10358);
and U10743 (N_10743,N_10149,N_9730);
xnor U10744 (N_10744,N_9800,N_10273);
and U10745 (N_10745,N_9840,N_9719);
nor U10746 (N_10746,N_9679,N_10260);
nand U10747 (N_10747,N_9903,N_9889);
and U10748 (N_10748,N_10387,N_10016);
and U10749 (N_10749,N_9851,N_9647);
and U10750 (N_10750,N_9912,N_9796);
xor U10751 (N_10751,N_10335,N_10396);
and U10752 (N_10752,N_9734,N_9637);
nor U10753 (N_10753,N_10081,N_9960);
nand U10754 (N_10754,N_10084,N_10059);
or U10755 (N_10755,N_10086,N_9956);
or U10756 (N_10756,N_10113,N_9830);
nor U10757 (N_10757,N_10320,N_10344);
nor U10758 (N_10758,N_9778,N_9629);
or U10759 (N_10759,N_10201,N_9648);
or U10760 (N_10760,N_9659,N_10227);
nor U10761 (N_10761,N_10193,N_10029);
and U10762 (N_10762,N_9725,N_10060);
and U10763 (N_10763,N_10202,N_10262);
nand U10764 (N_10764,N_9782,N_10342);
and U10765 (N_10765,N_10096,N_9607);
nand U10766 (N_10766,N_9902,N_9764);
xnor U10767 (N_10767,N_9781,N_10295);
xnor U10768 (N_10768,N_9733,N_9636);
nor U10769 (N_10769,N_10294,N_10014);
and U10770 (N_10770,N_10116,N_10177);
nand U10771 (N_10771,N_9985,N_9865);
nor U10772 (N_10772,N_9693,N_10063);
and U10773 (N_10773,N_9842,N_9610);
and U10774 (N_10774,N_9645,N_10160);
and U10775 (N_10775,N_10146,N_9625);
nand U10776 (N_10776,N_9661,N_9825);
or U10777 (N_10777,N_10343,N_9701);
nand U10778 (N_10778,N_9604,N_10173);
xnor U10779 (N_10779,N_9833,N_9845);
nand U10780 (N_10780,N_10309,N_9999);
nand U10781 (N_10781,N_9688,N_10239);
nor U10782 (N_10782,N_10001,N_10076);
nand U10783 (N_10783,N_10230,N_10068);
xnor U10784 (N_10784,N_10307,N_9994);
and U10785 (N_10785,N_10090,N_9904);
nor U10786 (N_10786,N_9876,N_10338);
and U10787 (N_10787,N_10155,N_10027);
or U10788 (N_10788,N_9906,N_9738);
xor U10789 (N_10789,N_10391,N_9760);
nor U10790 (N_10790,N_10111,N_9631);
xnor U10791 (N_10791,N_9981,N_10367);
nor U10792 (N_10792,N_10203,N_9724);
nor U10793 (N_10793,N_10327,N_10058);
nor U10794 (N_10794,N_10048,N_9850);
xor U10795 (N_10795,N_9691,N_9712);
nor U10796 (N_10796,N_9646,N_10075);
or U10797 (N_10797,N_9788,N_9623);
xor U10798 (N_10798,N_9795,N_10356);
and U10799 (N_10799,N_9608,N_9968);
nand U10800 (N_10800,N_9675,N_9724);
nand U10801 (N_10801,N_9952,N_9649);
xor U10802 (N_10802,N_9762,N_9740);
nand U10803 (N_10803,N_9788,N_9866);
or U10804 (N_10804,N_9862,N_9990);
xor U10805 (N_10805,N_10122,N_9653);
nor U10806 (N_10806,N_10375,N_10117);
and U10807 (N_10807,N_10230,N_10292);
or U10808 (N_10808,N_10038,N_10357);
nand U10809 (N_10809,N_10142,N_10147);
or U10810 (N_10810,N_10128,N_10310);
nor U10811 (N_10811,N_9747,N_10375);
nand U10812 (N_10812,N_9683,N_9682);
nand U10813 (N_10813,N_10343,N_9971);
nor U10814 (N_10814,N_10344,N_10290);
nand U10815 (N_10815,N_9852,N_10138);
or U10816 (N_10816,N_10290,N_10218);
xnor U10817 (N_10817,N_10362,N_10106);
nand U10818 (N_10818,N_9921,N_9852);
and U10819 (N_10819,N_9906,N_10074);
nor U10820 (N_10820,N_10206,N_9710);
xnor U10821 (N_10821,N_10221,N_10263);
nand U10822 (N_10822,N_10384,N_10054);
nand U10823 (N_10823,N_9674,N_10395);
nand U10824 (N_10824,N_10367,N_10299);
or U10825 (N_10825,N_10275,N_9643);
nand U10826 (N_10826,N_10382,N_9979);
nor U10827 (N_10827,N_10081,N_9971);
xnor U10828 (N_10828,N_9602,N_10037);
and U10829 (N_10829,N_10074,N_9709);
xnor U10830 (N_10830,N_10068,N_10246);
nor U10831 (N_10831,N_9791,N_10267);
nor U10832 (N_10832,N_10264,N_9631);
and U10833 (N_10833,N_10373,N_9775);
or U10834 (N_10834,N_9923,N_10249);
xnor U10835 (N_10835,N_9713,N_9757);
xnor U10836 (N_10836,N_9973,N_10042);
and U10837 (N_10837,N_10208,N_9949);
or U10838 (N_10838,N_9974,N_10176);
and U10839 (N_10839,N_9814,N_9688);
nor U10840 (N_10840,N_10290,N_9626);
and U10841 (N_10841,N_9934,N_10086);
nor U10842 (N_10842,N_10082,N_9769);
or U10843 (N_10843,N_9700,N_10219);
xnor U10844 (N_10844,N_10352,N_10384);
or U10845 (N_10845,N_10184,N_9760);
nand U10846 (N_10846,N_9689,N_9771);
nand U10847 (N_10847,N_10219,N_10254);
xor U10848 (N_10848,N_10205,N_10332);
and U10849 (N_10849,N_9603,N_10278);
and U10850 (N_10850,N_10179,N_10176);
nand U10851 (N_10851,N_10147,N_10378);
xnor U10852 (N_10852,N_10327,N_9900);
nand U10853 (N_10853,N_10295,N_10055);
nor U10854 (N_10854,N_10278,N_9630);
and U10855 (N_10855,N_9709,N_9867);
nor U10856 (N_10856,N_9959,N_10242);
xnor U10857 (N_10857,N_9770,N_9838);
or U10858 (N_10858,N_9786,N_10282);
nor U10859 (N_10859,N_9714,N_10273);
nor U10860 (N_10860,N_9668,N_9908);
nand U10861 (N_10861,N_10244,N_10053);
xnor U10862 (N_10862,N_10381,N_9613);
and U10863 (N_10863,N_10124,N_9692);
xor U10864 (N_10864,N_10386,N_10280);
or U10865 (N_10865,N_9805,N_10305);
nand U10866 (N_10866,N_9957,N_9605);
nand U10867 (N_10867,N_10329,N_9913);
xor U10868 (N_10868,N_10259,N_9955);
nand U10869 (N_10869,N_10365,N_9958);
and U10870 (N_10870,N_9936,N_10244);
xnor U10871 (N_10871,N_10203,N_10014);
xnor U10872 (N_10872,N_10159,N_9620);
xnor U10873 (N_10873,N_9898,N_10135);
and U10874 (N_10874,N_10038,N_10379);
nor U10875 (N_10875,N_10163,N_9833);
nand U10876 (N_10876,N_9986,N_10142);
xnor U10877 (N_10877,N_9745,N_9693);
nand U10878 (N_10878,N_10388,N_10015);
or U10879 (N_10879,N_10181,N_9629);
and U10880 (N_10880,N_10201,N_9953);
nand U10881 (N_10881,N_10169,N_9725);
nor U10882 (N_10882,N_10368,N_9649);
or U10883 (N_10883,N_9605,N_9754);
nor U10884 (N_10884,N_10345,N_10116);
or U10885 (N_10885,N_9682,N_9772);
xor U10886 (N_10886,N_10160,N_10275);
or U10887 (N_10887,N_9873,N_9851);
xor U10888 (N_10888,N_9859,N_9738);
nand U10889 (N_10889,N_10099,N_9737);
xnor U10890 (N_10890,N_9688,N_9825);
nand U10891 (N_10891,N_9698,N_9751);
or U10892 (N_10892,N_9971,N_9704);
nand U10893 (N_10893,N_10046,N_9765);
nor U10894 (N_10894,N_10112,N_10047);
and U10895 (N_10895,N_10314,N_10366);
xor U10896 (N_10896,N_9930,N_10012);
and U10897 (N_10897,N_10043,N_9974);
or U10898 (N_10898,N_10256,N_10076);
xor U10899 (N_10899,N_9607,N_9992);
xor U10900 (N_10900,N_10312,N_9711);
nand U10901 (N_10901,N_9765,N_10080);
xnor U10902 (N_10902,N_9640,N_9635);
or U10903 (N_10903,N_9811,N_10213);
or U10904 (N_10904,N_9945,N_10133);
and U10905 (N_10905,N_10299,N_9993);
or U10906 (N_10906,N_9929,N_9931);
and U10907 (N_10907,N_9994,N_9789);
nor U10908 (N_10908,N_9811,N_9819);
nor U10909 (N_10909,N_10382,N_10340);
nand U10910 (N_10910,N_10369,N_9700);
nor U10911 (N_10911,N_9678,N_10196);
and U10912 (N_10912,N_9733,N_10175);
nor U10913 (N_10913,N_10144,N_10121);
xor U10914 (N_10914,N_9938,N_9846);
and U10915 (N_10915,N_10303,N_9824);
and U10916 (N_10916,N_10309,N_9717);
nor U10917 (N_10917,N_10195,N_9635);
nand U10918 (N_10918,N_10099,N_9944);
nor U10919 (N_10919,N_10101,N_9988);
nand U10920 (N_10920,N_10228,N_10049);
and U10921 (N_10921,N_10007,N_9947);
xnor U10922 (N_10922,N_9860,N_10364);
and U10923 (N_10923,N_10020,N_9895);
or U10924 (N_10924,N_10279,N_9940);
nor U10925 (N_10925,N_10071,N_9757);
or U10926 (N_10926,N_10141,N_9921);
and U10927 (N_10927,N_10113,N_9761);
or U10928 (N_10928,N_9606,N_9973);
nand U10929 (N_10929,N_10325,N_9701);
xor U10930 (N_10930,N_9672,N_10044);
and U10931 (N_10931,N_9745,N_10263);
and U10932 (N_10932,N_10041,N_10212);
and U10933 (N_10933,N_9654,N_10097);
xnor U10934 (N_10934,N_10252,N_9927);
and U10935 (N_10935,N_9848,N_10243);
and U10936 (N_10936,N_9779,N_9994);
or U10937 (N_10937,N_10357,N_9758);
xnor U10938 (N_10938,N_9990,N_10109);
or U10939 (N_10939,N_9969,N_10117);
and U10940 (N_10940,N_10273,N_9600);
xor U10941 (N_10941,N_9704,N_10006);
and U10942 (N_10942,N_9770,N_9775);
nand U10943 (N_10943,N_10083,N_9710);
and U10944 (N_10944,N_10132,N_10389);
nand U10945 (N_10945,N_10228,N_10249);
nand U10946 (N_10946,N_9842,N_10046);
nand U10947 (N_10947,N_9925,N_9992);
xnor U10948 (N_10948,N_9616,N_9628);
nand U10949 (N_10949,N_10016,N_9654);
nor U10950 (N_10950,N_9662,N_10253);
nand U10951 (N_10951,N_9953,N_9864);
or U10952 (N_10952,N_10262,N_10042);
nor U10953 (N_10953,N_9924,N_9604);
nand U10954 (N_10954,N_9736,N_9722);
and U10955 (N_10955,N_10055,N_10111);
xnor U10956 (N_10956,N_9687,N_9886);
and U10957 (N_10957,N_9671,N_10302);
and U10958 (N_10958,N_9916,N_10155);
and U10959 (N_10959,N_9652,N_10348);
and U10960 (N_10960,N_10149,N_9919);
xor U10961 (N_10961,N_9715,N_9603);
xor U10962 (N_10962,N_10200,N_10051);
xor U10963 (N_10963,N_10047,N_9745);
nor U10964 (N_10964,N_10019,N_10063);
nand U10965 (N_10965,N_10331,N_10135);
xor U10966 (N_10966,N_10376,N_9986);
nand U10967 (N_10967,N_9677,N_9960);
nand U10968 (N_10968,N_10158,N_10181);
nor U10969 (N_10969,N_9990,N_10013);
nor U10970 (N_10970,N_9942,N_9774);
nand U10971 (N_10971,N_10039,N_10223);
nand U10972 (N_10972,N_10085,N_9647);
and U10973 (N_10973,N_10070,N_10089);
xnor U10974 (N_10974,N_9693,N_10371);
nor U10975 (N_10975,N_9994,N_10131);
or U10976 (N_10976,N_10273,N_9945);
nand U10977 (N_10977,N_10075,N_10224);
nor U10978 (N_10978,N_9615,N_9700);
and U10979 (N_10979,N_10107,N_10258);
and U10980 (N_10980,N_9811,N_10106);
and U10981 (N_10981,N_9863,N_10072);
and U10982 (N_10982,N_9747,N_9997);
or U10983 (N_10983,N_10067,N_9958);
nor U10984 (N_10984,N_9998,N_9646);
xor U10985 (N_10985,N_9778,N_10138);
nand U10986 (N_10986,N_10209,N_10343);
and U10987 (N_10987,N_10004,N_10371);
or U10988 (N_10988,N_9937,N_10308);
or U10989 (N_10989,N_9904,N_10351);
xor U10990 (N_10990,N_10371,N_10131);
nor U10991 (N_10991,N_9710,N_10236);
nand U10992 (N_10992,N_10375,N_10174);
nor U10993 (N_10993,N_9897,N_9995);
or U10994 (N_10994,N_9909,N_10045);
nor U10995 (N_10995,N_9928,N_9609);
nor U10996 (N_10996,N_10164,N_9920);
nand U10997 (N_10997,N_10278,N_10304);
nor U10998 (N_10998,N_9707,N_10060);
xor U10999 (N_10999,N_10056,N_10128);
nand U11000 (N_11000,N_9708,N_10116);
nand U11001 (N_11001,N_10238,N_10244);
xor U11002 (N_11002,N_9731,N_10221);
and U11003 (N_11003,N_9906,N_10299);
xor U11004 (N_11004,N_10125,N_10256);
or U11005 (N_11005,N_9700,N_9824);
nor U11006 (N_11006,N_10060,N_10272);
nor U11007 (N_11007,N_10148,N_10332);
or U11008 (N_11008,N_9653,N_9671);
xnor U11009 (N_11009,N_10012,N_9609);
nand U11010 (N_11010,N_9906,N_10140);
or U11011 (N_11011,N_9683,N_9677);
and U11012 (N_11012,N_9894,N_10048);
xnor U11013 (N_11013,N_10018,N_10185);
xor U11014 (N_11014,N_10239,N_9797);
xnor U11015 (N_11015,N_10297,N_9623);
and U11016 (N_11016,N_10243,N_10005);
nand U11017 (N_11017,N_10103,N_10198);
or U11018 (N_11018,N_10321,N_10389);
nand U11019 (N_11019,N_9920,N_9721);
nor U11020 (N_11020,N_10179,N_9881);
nor U11021 (N_11021,N_10019,N_9709);
nor U11022 (N_11022,N_9659,N_9703);
and U11023 (N_11023,N_10077,N_10267);
and U11024 (N_11024,N_10031,N_9756);
xnor U11025 (N_11025,N_9844,N_9649);
xor U11026 (N_11026,N_10289,N_10320);
xnor U11027 (N_11027,N_10309,N_10271);
and U11028 (N_11028,N_9673,N_10005);
nand U11029 (N_11029,N_9999,N_9979);
xor U11030 (N_11030,N_9882,N_9865);
and U11031 (N_11031,N_9847,N_9734);
nor U11032 (N_11032,N_9914,N_9922);
nor U11033 (N_11033,N_9832,N_9817);
xnor U11034 (N_11034,N_9696,N_10026);
nand U11035 (N_11035,N_9861,N_10082);
or U11036 (N_11036,N_10129,N_9924);
and U11037 (N_11037,N_9603,N_9801);
nand U11038 (N_11038,N_10097,N_10020);
xnor U11039 (N_11039,N_9943,N_9672);
nand U11040 (N_11040,N_10140,N_10213);
nand U11041 (N_11041,N_10112,N_9969);
nor U11042 (N_11042,N_10125,N_10261);
xor U11043 (N_11043,N_9993,N_9767);
nand U11044 (N_11044,N_10111,N_9627);
xor U11045 (N_11045,N_10282,N_9607);
nor U11046 (N_11046,N_10074,N_10228);
or U11047 (N_11047,N_9920,N_9869);
and U11048 (N_11048,N_10059,N_10245);
nor U11049 (N_11049,N_10178,N_9709);
nand U11050 (N_11050,N_9846,N_9887);
nor U11051 (N_11051,N_9926,N_9961);
nand U11052 (N_11052,N_10369,N_9717);
nand U11053 (N_11053,N_10091,N_10189);
nand U11054 (N_11054,N_9890,N_9736);
nor U11055 (N_11055,N_9878,N_9700);
xor U11056 (N_11056,N_10355,N_9920);
nor U11057 (N_11057,N_9950,N_9641);
xnor U11058 (N_11058,N_10347,N_9813);
or U11059 (N_11059,N_9956,N_9602);
xnor U11060 (N_11060,N_10272,N_10269);
nor U11061 (N_11061,N_9958,N_9764);
nand U11062 (N_11062,N_10183,N_9878);
or U11063 (N_11063,N_10122,N_9882);
nand U11064 (N_11064,N_9774,N_10256);
nor U11065 (N_11065,N_9894,N_9905);
nand U11066 (N_11066,N_9726,N_9817);
xnor U11067 (N_11067,N_10367,N_9994);
and U11068 (N_11068,N_9745,N_9654);
nor U11069 (N_11069,N_9714,N_10329);
nand U11070 (N_11070,N_10257,N_9996);
or U11071 (N_11071,N_10127,N_9773);
and U11072 (N_11072,N_10316,N_9905);
nand U11073 (N_11073,N_10343,N_9915);
and U11074 (N_11074,N_10335,N_9648);
and U11075 (N_11075,N_9768,N_9887);
xor U11076 (N_11076,N_9940,N_9879);
nor U11077 (N_11077,N_9869,N_9860);
or U11078 (N_11078,N_9665,N_9924);
nor U11079 (N_11079,N_9773,N_9811);
or U11080 (N_11080,N_9942,N_10317);
nand U11081 (N_11081,N_10389,N_10009);
nand U11082 (N_11082,N_9736,N_9869);
and U11083 (N_11083,N_10321,N_10055);
nor U11084 (N_11084,N_10011,N_9667);
nor U11085 (N_11085,N_9636,N_9719);
nor U11086 (N_11086,N_9640,N_10028);
xnor U11087 (N_11087,N_10039,N_10049);
or U11088 (N_11088,N_9785,N_10367);
nand U11089 (N_11089,N_9711,N_9932);
or U11090 (N_11090,N_9798,N_9607);
nand U11091 (N_11091,N_10059,N_9870);
nand U11092 (N_11092,N_9779,N_10094);
nand U11093 (N_11093,N_9749,N_10159);
and U11094 (N_11094,N_9683,N_9715);
xnor U11095 (N_11095,N_9634,N_10191);
or U11096 (N_11096,N_10131,N_10195);
nor U11097 (N_11097,N_10329,N_10350);
nand U11098 (N_11098,N_9815,N_10247);
nor U11099 (N_11099,N_10309,N_10234);
and U11100 (N_11100,N_10134,N_10124);
and U11101 (N_11101,N_9732,N_9983);
nand U11102 (N_11102,N_10337,N_10393);
nand U11103 (N_11103,N_9877,N_10268);
nand U11104 (N_11104,N_10291,N_10284);
and U11105 (N_11105,N_9681,N_9684);
nor U11106 (N_11106,N_10068,N_9868);
xor U11107 (N_11107,N_10100,N_9629);
nand U11108 (N_11108,N_9847,N_10157);
nor U11109 (N_11109,N_10295,N_10370);
or U11110 (N_11110,N_9987,N_9856);
and U11111 (N_11111,N_10167,N_10369);
nor U11112 (N_11112,N_9901,N_10178);
xnor U11113 (N_11113,N_10181,N_10379);
nand U11114 (N_11114,N_10121,N_9659);
nand U11115 (N_11115,N_9770,N_10169);
nor U11116 (N_11116,N_10283,N_10145);
nor U11117 (N_11117,N_10221,N_10026);
nor U11118 (N_11118,N_10301,N_10356);
xor U11119 (N_11119,N_10090,N_9820);
nand U11120 (N_11120,N_9949,N_9652);
or U11121 (N_11121,N_10290,N_9797);
nand U11122 (N_11122,N_10141,N_10380);
nand U11123 (N_11123,N_10134,N_9714);
nor U11124 (N_11124,N_10007,N_9788);
nor U11125 (N_11125,N_9955,N_9616);
or U11126 (N_11126,N_10166,N_9803);
or U11127 (N_11127,N_9641,N_10168);
nand U11128 (N_11128,N_9866,N_9641);
or U11129 (N_11129,N_9802,N_10339);
and U11130 (N_11130,N_10077,N_9962);
nor U11131 (N_11131,N_9899,N_10090);
and U11132 (N_11132,N_10191,N_9655);
xnor U11133 (N_11133,N_9683,N_10075);
or U11134 (N_11134,N_9681,N_9690);
or U11135 (N_11135,N_10105,N_10272);
and U11136 (N_11136,N_9942,N_10026);
and U11137 (N_11137,N_9797,N_9875);
or U11138 (N_11138,N_9601,N_10100);
xor U11139 (N_11139,N_10255,N_9678);
nand U11140 (N_11140,N_9603,N_9768);
xor U11141 (N_11141,N_9761,N_10347);
or U11142 (N_11142,N_10041,N_9724);
nor U11143 (N_11143,N_9952,N_10036);
nand U11144 (N_11144,N_9873,N_9658);
and U11145 (N_11145,N_10318,N_10088);
nand U11146 (N_11146,N_10015,N_10385);
and U11147 (N_11147,N_9753,N_10013);
nor U11148 (N_11148,N_10005,N_10343);
nand U11149 (N_11149,N_10118,N_10051);
and U11150 (N_11150,N_9768,N_9963);
xnor U11151 (N_11151,N_9652,N_9996);
or U11152 (N_11152,N_9863,N_10343);
or U11153 (N_11153,N_10080,N_10122);
xor U11154 (N_11154,N_10035,N_10246);
nand U11155 (N_11155,N_10087,N_10212);
xnor U11156 (N_11156,N_10177,N_9943);
or U11157 (N_11157,N_10248,N_10062);
or U11158 (N_11158,N_10078,N_10004);
or U11159 (N_11159,N_10021,N_9746);
or U11160 (N_11160,N_10293,N_9861);
nor U11161 (N_11161,N_10162,N_9898);
nor U11162 (N_11162,N_10172,N_9800);
xor U11163 (N_11163,N_9787,N_10184);
nand U11164 (N_11164,N_9720,N_9680);
nor U11165 (N_11165,N_10296,N_10241);
and U11166 (N_11166,N_10149,N_10154);
or U11167 (N_11167,N_10126,N_10119);
nor U11168 (N_11168,N_10357,N_10323);
xor U11169 (N_11169,N_10083,N_9811);
xor U11170 (N_11170,N_9721,N_10003);
nand U11171 (N_11171,N_9913,N_10143);
xor U11172 (N_11172,N_10259,N_9812);
xnor U11173 (N_11173,N_9651,N_9669);
and U11174 (N_11174,N_10139,N_9961);
and U11175 (N_11175,N_9857,N_9852);
or U11176 (N_11176,N_9777,N_9670);
and U11177 (N_11177,N_9809,N_9884);
nand U11178 (N_11178,N_10070,N_9748);
xnor U11179 (N_11179,N_10263,N_9623);
xnor U11180 (N_11180,N_10060,N_10062);
nor U11181 (N_11181,N_10203,N_9844);
nor U11182 (N_11182,N_10329,N_10072);
or U11183 (N_11183,N_9789,N_10264);
nand U11184 (N_11184,N_9650,N_10074);
nand U11185 (N_11185,N_9805,N_9943);
nand U11186 (N_11186,N_10339,N_9833);
and U11187 (N_11187,N_10393,N_10207);
nor U11188 (N_11188,N_10351,N_9679);
nand U11189 (N_11189,N_10226,N_9885);
or U11190 (N_11190,N_9684,N_9651);
and U11191 (N_11191,N_9859,N_9726);
xnor U11192 (N_11192,N_10020,N_9904);
and U11193 (N_11193,N_10242,N_9909);
and U11194 (N_11194,N_9990,N_9797);
nor U11195 (N_11195,N_10072,N_9874);
xnor U11196 (N_11196,N_10050,N_9814);
or U11197 (N_11197,N_9912,N_9996);
nand U11198 (N_11198,N_9602,N_9628);
nor U11199 (N_11199,N_10201,N_10321);
nor U11200 (N_11200,N_10409,N_10534);
or U11201 (N_11201,N_10817,N_10750);
or U11202 (N_11202,N_10914,N_10622);
or U11203 (N_11203,N_10828,N_11018);
nor U11204 (N_11204,N_10406,N_10710);
nand U11205 (N_11205,N_10713,N_10469);
xor U11206 (N_11206,N_11153,N_10641);
nand U11207 (N_11207,N_10642,N_10401);
or U11208 (N_11208,N_10560,N_10597);
nand U11209 (N_11209,N_10577,N_11122);
xor U11210 (N_11210,N_10716,N_10510);
or U11211 (N_11211,N_10741,N_11103);
and U11212 (N_11212,N_10978,N_10529);
nor U11213 (N_11213,N_11115,N_11031);
nand U11214 (N_11214,N_11167,N_10747);
nand U11215 (N_11215,N_10926,N_11160);
nor U11216 (N_11216,N_11157,N_11135);
xnor U11217 (N_11217,N_11041,N_10693);
xor U11218 (N_11218,N_10790,N_10943);
and U11219 (N_11219,N_10851,N_11093);
and U11220 (N_11220,N_10743,N_11178);
nand U11221 (N_11221,N_10946,N_10781);
xnor U11222 (N_11222,N_10620,N_10488);
nor U11223 (N_11223,N_10859,N_10563);
nand U11224 (N_11224,N_10508,N_11111);
and U11225 (N_11225,N_10649,N_11173);
nand U11226 (N_11226,N_10452,N_11143);
or U11227 (N_11227,N_10681,N_10553);
or U11228 (N_11228,N_10561,N_11154);
or U11229 (N_11229,N_11015,N_10400);
nand U11230 (N_11230,N_10595,N_10800);
nand U11231 (N_11231,N_11047,N_10703);
nand U11232 (N_11232,N_10673,N_10919);
nor U11233 (N_11233,N_11027,N_10503);
nand U11234 (N_11234,N_10773,N_11013);
nand U11235 (N_11235,N_10481,N_10446);
or U11236 (N_11236,N_10835,N_10516);
or U11237 (N_11237,N_10822,N_10653);
nor U11238 (N_11238,N_11089,N_10875);
and U11239 (N_11239,N_10573,N_10700);
nand U11240 (N_11240,N_10645,N_10432);
nor U11241 (N_11241,N_10833,N_11140);
xnor U11242 (N_11242,N_10928,N_10434);
xor U11243 (N_11243,N_10632,N_10769);
or U11244 (N_11244,N_11119,N_11126);
nor U11245 (N_11245,N_11005,N_10858);
nor U11246 (N_11246,N_10813,N_10427);
and U11247 (N_11247,N_10890,N_11044);
or U11248 (N_11248,N_11083,N_10715);
xnor U11249 (N_11249,N_10707,N_10625);
nand U11250 (N_11250,N_10907,N_11149);
nor U11251 (N_11251,N_10698,N_11079);
xnor U11252 (N_11252,N_11125,N_10784);
or U11253 (N_11253,N_10610,N_11051);
xor U11254 (N_11254,N_10497,N_10479);
and U11255 (N_11255,N_10518,N_10493);
nand U11256 (N_11256,N_10902,N_10783);
nand U11257 (N_11257,N_10547,N_10473);
and U11258 (N_11258,N_11170,N_10911);
xor U11259 (N_11259,N_10635,N_11068);
nand U11260 (N_11260,N_11164,N_10687);
or U11261 (N_11261,N_10419,N_10571);
nor U11262 (N_11262,N_10604,N_10442);
xor U11263 (N_11263,N_10865,N_10850);
nand U11264 (N_11264,N_10517,N_10896);
and U11265 (N_11265,N_10466,N_10557);
or U11266 (N_11266,N_10990,N_10694);
nand U11267 (N_11267,N_10970,N_11175);
or U11268 (N_11268,N_10929,N_10788);
nand U11269 (N_11269,N_10616,N_10847);
xor U11270 (N_11270,N_11075,N_10458);
nand U11271 (N_11271,N_10941,N_10798);
xnor U11272 (N_11272,N_10898,N_10974);
or U11273 (N_11273,N_10609,N_10832);
or U11274 (N_11274,N_11024,N_10861);
or U11275 (N_11275,N_11000,N_10433);
and U11276 (N_11276,N_10845,N_10735);
xor U11277 (N_11277,N_11011,N_10712);
xor U11278 (N_11278,N_11091,N_10778);
nand U11279 (N_11279,N_10532,N_10936);
and U11280 (N_11280,N_11003,N_11107);
nand U11281 (N_11281,N_10762,N_11037);
nand U11282 (N_11282,N_11069,N_10939);
xor U11283 (N_11283,N_10869,N_10995);
and U11284 (N_11284,N_11072,N_11188);
xor U11285 (N_11285,N_10966,N_10894);
nand U11286 (N_11286,N_11120,N_10696);
nand U11287 (N_11287,N_10821,N_10945);
xnor U11288 (N_11288,N_11004,N_11033);
and U11289 (N_11289,N_10721,N_10787);
or U11290 (N_11290,N_10528,N_10470);
or U11291 (N_11291,N_10507,N_10885);
nand U11292 (N_11292,N_10905,N_10566);
nor U11293 (N_11293,N_10500,N_10531);
and U11294 (N_11294,N_10872,N_11073);
or U11295 (N_11295,N_10562,N_11195);
or U11296 (N_11296,N_11062,N_11010);
nor U11297 (N_11297,N_10570,N_11029);
or U11298 (N_11298,N_10889,N_11116);
nor U11299 (N_11299,N_10659,N_11114);
and U11300 (N_11300,N_10779,N_10668);
or U11301 (N_11301,N_10949,N_10786);
xor U11302 (N_11302,N_10957,N_10471);
nor U11303 (N_11303,N_10881,N_10756);
xor U11304 (N_11304,N_10654,N_10969);
xnor U11305 (N_11305,N_10676,N_10476);
xor U11306 (N_11306,N_10864,N_10624);
nor U11307 (N_11307,N_10414,N_10979);
nand U11308 (N_11308,N_10590,N_11058);
xor U11309 (N_11309,N_11155,N_10639);
and U11310 (N_11310,N_11057,N_10634);
xor U11311 (N_11311,N_11194,N_10648);
or U11312 (N_11312,N_11189,N_10780);
xor U11313 (N_11313,N_10491,N_11141);
nand U11314 (N_11314,N_10718,N_11106);
nor U11315 (N_11315,N_11049,N_10818);
or U11316 (N_11316,N_11007,N_10520);
xnor U11317 (N_11317,N_11076,N_10582);
or U11318 (N_11318,N_11162,N_10489);
nor U11319 (N_11319,N_11132,N_11064);
nand U11320 (N_11320,N_10525,N_10922);
nor U11321 (N_11321,N_10951,N_11008);
nor U11322 (N_11322,N_10724,N_11133);
and U11323 (N_11323,N_10499,N_10965);
xnor U11324 (N_11324,N_10695,N_10448);
or U11325 (N_11325,N_10436,N_10999);
nor U11326 (N_11326,N_10884,N_10917);
nand U11327 (N_11327,N_10888,N_11046);
xor U11328 (N_11328,N_10596,N_10853);
nor U11329 (N_11329,N_10740,N_10672);
nor U11330 (N_11330,N_10440,N_10456);
or U11331 (N_11331,N_10421,N_10876);
nor U11332 (N_11332,N_10737,N_10892);
or U11333 (N_11333,N_10468,N_10554);
and U11334 (N_11334,N_10731,N_11048);
or U11335 (N_11335,N_10738,N_11165);
or U11336 (N_11336,N_11006,N_10912);
nor U11337 (N_11337,N_10660,N_11028);
xor U11338 (N_11338,N_10956,N_10599);
nor U11339 (N_11339,N_10423,N_11053);
or U11340 (N_11340,N_10906,N_11142);
or U11341 (N_11341,N_10429,N_10708);
xor U11342 (N_11342,N_10996,N_10524);
and U11343 (N_11343,N_11012,N_10574);
nor U11344 (N_11344,N_10584,N_10730);
and U11345 (N_11345,N_10823,N_11179);
xor U11346 (N_11346,N_10474,N_10486);
or U11347 (N_11347,N_10935,N_11127);
and U11348 (N_11348,N_11022,N_10492);
or U11349 (N_11349,N_10402,N_10799);
nand U11350 (N_11350,N_10829,N_10539);
nand U11351 (N_11351,N_10496,N_10689);
nand U11352 (N_11352,N_11110,N_10722);
and U11353 (N_11353,N_11025,N_10631);
and U11354 (N_11354,N_10711,N_10580);
nand U11355 (N_11355,N_11134,N_10449);
xnor U11356 (N_11356,N_11085,N_11118);
xor U11357 (N_11357,N_11105,N_10953);
xnor U11358 (N_11358,N_10411,N_10575);
or U11359 (N_11359,N_10504,N_10831);
nand U11360 (N_11360,N_11055,N_10931);
nand U11361 (N_11361,N_10751,N_11169);
or U11362 (N_11362,N_10736,N_11067);
nor U11363 (N_11363,N_10552,N_11052);
nor U11364 (N_11364,N_10565,N_10871);
or U11365 (N_11365,N_10963,N_10512);
or U11366 (N_11366,N_10544,N_10453);
and U11367 (N_11367,N_11036,N_10691);
or U11368 (N_11368,N_11161,N_11128);
nor U11369 (N_11369,N_10412,N_10472);
xor U11370 (N_11370,N_10640,N_10704);
or U11371 (N_11371,N_10482,N_10603);
nor U11372 (N_11372,N_10623,N_11176);
and U11373 (N_11373,N_10771,N_10581);
nor U11374 (N_11374,N_10729,N_10863);
nand U11375 (N_11375,N_10723,N_10830);
or U11376 (N_11376,N_10742,N_11177);
and U11377 (N_11377,N_10579,N_11123);
nor U11378 (N_11378,N_10556,N_10985);
nand U11379 (N_11379,N_10443,N_10658);
and U11380 (N_11380,N_11113,N_10701);
nand U11381 (N_11381,N_10551,N_10594);
nor U11382 (N_11382,N_11020,N_10638);
and U11383 (N_11383,N_10606,N_11183);
and U11384 (N_11384,N_10855,N_11130);
and U11385 (N_11385,N_11019,N_10948);
nor U11386 (N_11386,N_11163,N_10820);
and U11387 (N_11387,N_10526,N_10967);
xnor U11388 (N_11388,N_10805,N_10857);
xor U11389 (N_11389,N_10464,N_10643);
xor U11390 (N_11390,N_10420,N_10842);
or U11391 (N_11391,N_10921,N_10749);
and U11392 (N_11392,N_10826,N_10618);
nor U11393 (N_11393,N_10777,N_10873);
or U11394 (N_11394,N_10761,N_10686);
nand U11395 (N_11395,N_10775,N_10734);
or U11396 (N_11396,N_10515,N_10808);
nand U11397 (N_11397,N_11171,N_11146);
xnor U11398 (N_11398,N_10568,N_10717);
nor U11399 (N_11399,N_10688,N_10569);
xor U11400 (N_11400,N_10991,N_10891);
nor U11401 (N_11401,N_10883,N_10657);
and U11402 (N_11402,N_10772,N_10984);
xor U11403 (N_11403,N_10457,N_10690);
and U11404 (N_11404,N_10454,N_10522);
nand U11405 (N_11405,N_10810,N_10932);
nor U11406 (N_11406,N_10903,N_11186);
xor U11407 (N_11407,N_10587,N_11148);
and U11408 (N_11408,N_11109,N_10795);
or U11409 (N_11409,N_11065,N_10611);
nand U11410 (N_11410,N_10460,N_10844);
nand U11411 (N_11411,N_10725,N_10886);
xor U11412 (N_11412,N_10824,N_10767);
and U11413 (N_11413,N_10564,N_10843);
nor U11414 (N_11414,N_10980,N_11151);
nand U11415 (N_11415,N_10602,N_10535);
xnor U11416 (N_11416,N_10678,N_10816);
and U11417 (N_11417,N_11040,N_10997);
nor U11418 (N_11418,N_11059,N_10484);
nand U11419 (N_11419,N_10954,N_10437);
xor U11420 (N_11420,N_10477,N_10502);
nand U11421 (N_11421,N_11166,N_10684);
nand U11422 (N_11422,N_10555,N_10438);
xnor U11423 (N_11423,N_10679,N_10768);
xor U11424 (N_11424,N_11185,N_10893);
and U11425 (N_11425,N_10913,N_10920);
or U11426 (N_11426,N_11156,N_10593);
or U11427 (N_11427,N_10656,N_10900);
xnor U11428 (N_11428,N_11192,N_10463);
or U11429 (N_11429,N_10404,N_10880);
or U11430 (N_11430,N_10827,N_11074);
nand U11431 (N_11431,N_10589,N_10930);
and U11432 (N_11432,N_11112,N_10705);
nor U11433 (N_11433,N_10462,N_10619);
or U11434 (N_11434,N_10514,N_10549);
and U11435 (N_11435,N_10495,N_10938);
nor U11436 (N_11436,N_10878,N_10692);
xnor U11437 (N_11437,N_11180,N_10754);
or U11438 (N_11438,N_10545,N_10807);
and U11439 (N_11439,N_10636,N_10674);
or U11440 (N_11440,N_10647,N_10428);
and U11441 (N_11441,N_10812,N_10766);
nand U11442 (N_11442,N_10794,N_10425);
nand U11443 (N_11443,N_10699,N_11139);
nor U11444 (N_11444,N_11100,N_11095);
nor U11445 (N_11445,N_10910,N_10637);
or U11446 (N_11446,N_10802,N_10879);
nand U11447 (N_11447,N_10803,N_11066);
nor U11448 (N_11448,N_10537,N_10973);
nand U11449 (N_11449,N_11150,N_10501);
xor U11450 (N_11450,N_10441,N_11184);
nor U11451 (N_11451,N_10804,N_11082);
or U11452 (N_11452,N_11094,N_10439);
and U11453 (N_11453,N_10998,N_10901);
or U11454 (N_11454,N_11145,N_10567);
and U11455 (N_11455,N_10986,N_10664);
nand U11456 (N_11456,N_10955,N_10494);
nor U11457 (N_11457,N_10976,N_10774);
nor U11458 (N_11458,N_10940,N_10937);
or U11459 (N_11459,N_10848,N_10870);
xor U11460 (N_11460,N_11038,N_10837);
xnor U11461 (N_11461,N_11056,N_11017);
or U11462 (N_11462,N_10644,N_10895);
or U11463 (N_11463,N_10728,N_10506);
and U11464 (N_11464,N_10485,N_10416);
and U11465 (N_11465,N_11144,N_10629);
nand U11466 (N_11466,N_10413,N_10867);
nand U11467 (N_11467,N_10916,N_10801);
xor U11468 (N_11468,N_10576,N_11191);
xor U11469 (N_11469,N_10430,N_10868);
and U11470 (N_11470,N_11078,N_10670);
and U11471 (N_11471,N_10982,N_10947);
xnor U11472 (N_11472,N_11071,N_10697);
xnor U11473 (N_11473,N_11086,N_11080);
or U11474 (N_11474,N_10809,N_10548);
nor U11475 (N_11475,N_10942,N_10748);
or U11476 (N_11476,N_11035,N_10757);
xor U11477 (N_11477,N_10760,N_10753);
nand U11478 (N_11478,N_11063,N_10509);
xor U11479 (N_11479,N_10732,N_11077);
xnor U11480 (N_11480,N_10633,N_10680);
nand U11481 (N_11481,N_10445,N_10405);
and U11482 (N_11482,N_10669,N_10988);
xor U11483 (N_11483,N_10983,N_10461);
nor U11484 (N_11484,N_10483,N_10758);
or U11485 (N_11485,N_10671,N_10585);
nor U11486 (N_11486,N_10934,N_11104);
or U11487 (N_11487,N_10615,N_10498);
nor U11488 (N_11488,N_11193,N_11026);
or U11489 (N_11489,N_10646,N_10877);
and U11490 (N_11490,N_11001,N_10543);
xnor U11491 (N_11491,N_10605,N_10887);
nand U11492 (N_11492,N_10559,N_10950);
nor U11493 (N_11493,N_11138,N_10782);
or U11494 (N_11494,N_10993,N_10770);
nor U11495 (N_11495,N_10542,N_10422);
or U11496 (N_11496,N_10661,N_10763);
xnor U11497 (N_11497,N_10811,N_10550);
nand U11498 (N_11498,N_10806,N_10431);
xor U11499 (N_11499,N_10959,N_10675);
xor U11500 (N_11500,N_11060,N_10839);
or U11501 (N_11501,N_10815,N_10987);
or U11502 (N_11502,N_10752,N_10797);
nand U11503 (N_11503,N_10796,N_10612);
and U11504 (N_11504,N_10408,N_10655);
and U11505 (N_11505,N_10765,N_11061);
xnor U11506 (N_11506,N_10992,N_10666);
xnor U11507 (N_11507,N_10600,N_10511);
nor U11508 (N_11508,N_11092,N_11102);
nor U11509 (N_11509,N_10759,N_10960);
or U11510 (N_11510,N_10685,N_11172);
xnor U11511 (N_11511,N_10410,N_10709);
xnor U11512 (N_11512,N_10519,N_10899);
nand U11513 (N_11513,N_10546,N_11131);
nor U11514 (N_11514,N_11197,N_10487);
and U11515 (N_11515,N_11136,N_11129);
or U11516 (N_11516,N_11032,N_11054);
or U11517 (N_11517,N_11023,N_10836);
or U11518 (N_11518,N_10592,N_10952);
and U11519 (N_11519,N_11137,N_11152);
nand U11520 (N_11520,N_11039,N_10746);
and U11521 (N_11521,N_11034,N_11108);
xor U11522 (N_11522,N_10683,N_10825);
nor U11523 (N_11523,N_10475,N_10521);
nand U11524 (N_11524,N_10426,N_10677);
xnor U11525 (N_11525,N_10651,N_10994);
and U11526 (N_11526,N_10846,N_10793);
xnor U11527 (N_11527,N_10706,N_11187);
nor U11528 (N_11528,N_10785,N_10650);
nor U11529 (N_11529,N_11021,N_11174);
xnor U11530 (N_11530,N_10834,N_11147);
nor U11531 (N_11531,N_11030,N_10527);
or U11532 (N_11532,N_10447,N_10424);
or U11533 (N_11533,N_10925,N_11009);
nor U11534 (N_11534,N_10933,N_10923);
and U11535 (N_11535,N_10714,N_10702);
and U11536 (N_11536,N_10613,N_11016);
xor U11537 (N_11537,N_10513,N_10478);
nor U11538 (N_11538,N_10791,N_10977);
or U11539 (N_11539,N_10862,N_11101);
xnor U11540 (N_11540,N_10918,N_10776);
or U11541 (N_11541,N_10755,N_10908);
and U11542 (N_11542,N_11168,N_10860);
nand U11543 (N_11543,N_10630,N_10958);
nand U11544 (N_11544,N_11196,N_11087);
nor U11545 (N_11545,N_11096,N_10628);
or U11546 (N_11546,N_11190,N_10989);
or U11547 (N_11547,N_10558,N_10856);
or U11548 (N_11548,N_11181,N_10682);
xnor U11549 (N_11549,N_10726,N_10444);
and U11550 (N_11550,N_10621,N_11045);
nor U11551 (N_11551,N_10418,N_10854);
or U11552 (N_11552,N_10415,N_11099);
and U11553 (N_11553,N_10578,N_10403);
nand U11554 (N_11554,N_10819,N_11002);
nor U11555 (N_11555,N_10533,N_10407);
nor U11556 (N_11556,N_10459,N_11159);
and U11557 (N_11557,N_11117,N_10662);
nor U11558 (N_11558,N_11158,N_10838);
xnor U11559 (N_11559,N_10626,N_10739);
xor U11560 (N_11560,N_10792,N_10727);
xor U11561 (N_11561,N_10764,N_10451);
and U11562 (N_11562,N_10450,N_10614);
xnor U11563 (N_11563,N_10652,N_11121);
nor U11564 (N_11564,N_10627,N_10607);
nor U11565 (N_11565,N_10598,N_11070);
nor U11566 (N_11566,N_10882,N_10435);
nand U11567 (N_11567,N_10505,N_10975);
or U11568 (N_11568,N_10540,N_10490);
or U11569 (N_11569,N_10536,N_10745);
nor U11570 (N_11570,N_10572,N_10971);
and U11571 (N_11571,N_10523,N_10719);
or U11572 (N_11572,N_10733,N_10541);
nor U11573 (N_11573,N_10455,N_10530);
nand U11574 (N_11574,N_10961,N_11042);
nand U11575 (N_11575,N_10852,N_10909);
xnor U11576 (N_11576,N_10583,N_10849);
or U11577 (N_11577,N_11014,N_11088);
nor U11578 (N_11578,N_10904,N_11124);
xor U11579 (N_11579,N_11098,N_10927);
nand U11580 (N_11580,N_10814,N_11199);
xnor U11581 (N_11581,N_10840,N_10962);
xnor U11582 (N_11582,N_10964,N_10924);
nand U11583 (N_11583,N_10538,N_10968);
nor U11584 (N_11584,N_10586,N_11198);
nand U11585 (N_11585,N_10981,N_10608);
xnor U11586 (N_11586,N_10617,N_11081);
nand U11587 (N_11587,N_11043,N_10744);
nand U11588 (N_11588,N_10874,N_10897);
or U11589 (N_11589,N_11084,N_10665);
nand U11590 (N_11590,N_10417,N_10915);
xor U11591 (N_11591,N_10866,N_10588);
xor U11592 (N_11592,N_10467,N_10465);
nand U11593 (N_11593,N_10667,N_11050);
or U11594 (N_11594,N_10601,N_11182);
and U11595 (N_11595,N_10789,N_11090);
xnor U11596 (N_11596,N_10841,N_10663);
xnor U11597 (N_11597,N_10480,N_10720);
nand U11598 (N_11598,N_10944,N_10972);
xnor U11599 (N_11599,N_10591,N_11097);
nand U11600 (N_11600,N_11029,N_11058);
nand U11601 (N_11601,N_10420,N_10744);
and U11602 (N_11602,N_10577,N_10651);
xnor U11603 (N_11603,N_10408,N_10417);
nand U11604 (N_11604,N_11130,N_10545);
nor U11605 (N_11605,N_11180,N_11074);
nor U11606 (N_11606,N_11031,N_10772);
nor U11607 (N_11607,N_11152,N_10509);
and U11608 (N_11608,N_10553,N_11029);
nand U11609 (N_11609,N_10764,N_10815);
nand U11610 (N_11610,N_10732,N_10509);
or U11611 (N_11611,N_10934,N_10441);
xnor U11612 (N_11612,N_10809,N_10552);
nand U11613 (N_11613,N_10598,N_11041);
and U11614 (N_11614,N_10623,N_10734);
xnor U11615 (N_11615,N_10732,N_11093);
xnor U11616 (N_11616,N_10542,N_10851);
and U11617 (N_11617,N_11080,N_10825);
nand U11618 (N_11618,N_11019,N_10810);
xnor U11619 (N_11619,N_10710,N_10460);
nand U11620 (N_11620,N_11131,N_10413);
or U11621 (N_11621,N_10949,N_10916);
or U11622 (N_11622,N_11189,N_10860);
nor U11623 (N_11623,N_10993,N_10543);
xor U11624 (N_11624,N_10836,N_10500);
and U11625 (N_11625,N_10715,N_11180);
nor U11626 (N_11626,N_10544,N_10983);
nand U11627 (N_11627,N_10994,N_11168);
xor U11628 (N_11628,N_10895,N_10997);
nand U11629 (N_11629,N_11071,N_11118);
or U11630 (N_11630,N_11010,N_10821);
and U11631 (N_11631,N_10485,N_11150);
and U11632 (N_11632,N_10922,N_10712);
and U11633 (N_11633,N_11146,N_11095);
xor U11634 (N_11634,N_10838,N_10799);
xor U11635 (N_11635,N_10938,N_10516);
and U11636 (N_11636,N_10867,N_10683);
nand U11637 (N_11637,N_10577,N_10828);
and U11638 (N_11638,N_10916,N_10439);
nor U11639 (N_11639,N_10949,N_10852);
nor U11640 (N_11640,N_10415,N_10900);
xnor U11641 (N_11641,N_10903,N_11080);
and U11642 (N_11642,N_11084,N_10770);
and U11643 (N_11643,N_10775,N_10741);
nand U11644 (N_11644,N_10510,N_10831);
nor U11645 (N_11645,N_11140,N_10790);
nand U11646 (N_11646,N_10845,N_10771);
nand U11647 (N_11647,N_10589,N_10780);
and U11648 (N_11648,N_10462,N_10865);
nor U11649 (N_11649,N_11111,N_11049);
or U11650 (N_11650,N_10864,N_10719);
nand U11651 (N_11651,N_10575,N_11025);
or U11652 (N_11652,N_10583,N_10417);
or U11653 (N_11653,N_10713,N_10680);
or U11654 (N_11654,N_10494,N_10815);
or U11655 (N_11655,N_10730,N_10954);
nand U11656 (N_11656,N_10926,N_10746);
or U11657 (N_11657,N_10896,N_10513);
nor U11658 (N_11658,N_10490,N_11114);
nand U11659 (N_11659,N_10533,N_11002);
or U11660 (N_11660,N_10472,N_10444);
nand U11661 (N_11661,N_11094,N_10481);
xnor U11662 (N_11662,N_10553,N_10822);
and U11663 (N_11663,N_10748,N_10951);
xnor U11664 (N_11664,N_10988,N_10840);
and U11665 (N_11665,N_11000,N_11088);
xor U11666 (N_11666,N_11126,N_10528);
nand U11667 (N_11667,N_10803,N_11052);
xor U11668 (N_11668,N_10669,N_10965);
xnor U11669 (N_11669,N_10993,N_11092);
nand U11670 (N_11670,N_10786,N_10917);
and U11671 (N_11671,N_10991,N_11023);
or U11672 (N_11672,N_10636,N_10762);
nand U11673 (N_11673,N_10411,N_10993);
or U11674 (N_11674,N_10469,N_10453);
and U11675 (N_11675,N_10984,N_10478);
nor U11676 (N_11676,N_11026,N_11030);
xnor U11677 (N_11677,N_10819,N_11182);
and U11678 (N_11678,N_10834,N_10591);
xor U11679 (N_11679,N_10586,N_10917);
xnor U11680 (N_11680,N_11001,N_10561);
xnor U11681 (N_11681,N_10663,N_10859);
xor U11682 (N_11682,N_10671,N_10456);
xnor U11683 (N_11683,N_11149,N_10424);
xor U11684 (N_11684,N_10842,N_10539);
and U11685 (N_11685,N_10478,N_10824);
nand U11686 (N_11686,N_10470,N_10987);
nand U11687 (N_11687,N_10907,N_10481);
or U11688 (N_11688,N_10504,N_10995);
nor U11689 (N_11689,N_10609,N_10907);
nand U11690 (N_11690,N_10446,N_11071);
nand U11691 (N_11691,N_10875,N_11033);
or U11692 (N_11692,N_10875,N_10401);
xnor U11693 (N_11693,N_11005,N_11014);
xnor U11694 (N_11694,N_10851,N_10634);
nand U11695 (N_11695,N_11193,N_11194);
and U11696 (N_11696,N_10911,N_10859);
or U11697 (N_11697,N_10739,N_11118);
and U11698 (N_11698,N_10464,N_10795);
nand U11699 (N_11699,N_10663,N_10985);
xnor U11700 (N_11700,N_11084,N_11162);
nor U11701 (N_11701,N_11145,N_10850);
or U11702 (N_11702,N_10521,N_10825);
nand U11703 (N_11703,N_10860,N_10760);
and U11704 (N_11704,N_10415,N_10637);
and U11705 (N_11705,N_10703,N_11012);
and U11706 (N_11706,N_11087,N_10942);
nand U11707 (N_11707,N_11043,N_11134);
or U11708 (N_11708,N_10642,N_10800);
nor U11709 (N_11709,N_10751,N_10591);
nand U11710 (N_11710,N_10863,N_10601);
or U11711 (N_11711,N_10498,N_10613);
nor U11712 (N_11712,N_10950,N_11136);
or U11713 (N_11713,N_10403,N_11185);
xor U11714 (N_11714,N_11063,N_10984);
nor U11715 (N_11715,N_10861,N_11020);
and U11716 (N_11716,N_10780,N_11127);
and U11717 (N_11717,N_10676,N_10668);
xor U11718 (N_11718,N_10440,N_10969);
and U11719 (N_11719,N_11057,N_10926);
nor U11720 (N_11720,N_10620,N_10559);
and U11721 (N_11721,N_11095,N_10434);
nor U11722 (N_11722,N_10528,N_10509);
and U11723 (N_11723,N_10852,N_10858);
nand U11724 (N_11724,N_10987,N_11010);
nand U11725 (N_11725,N_10794,N_10956);
nor U11726 (N_11726,N_10877,N_11105);
and U11727 (N_11727,N_10769,N_11097);
xor U11728 (N_11728,N_10444,N_10446);
xnor U11729 (N_11729,N_10546,N_10625);
xor U11730 (N_11730,N_11005,N_10566);
or U11731 (N_11731,N_10491,N_10961);
and U11732 (N_11732,N_10757,N_10861);
nand U11733 (N_11733,N_11063,N_10956);
or U11734 (N_11734,N_10540,N_10954);
nor U11735 (N_11735,N_11085,N_11197);
and U11736 (N_11736,N_10654,N_10867);
xor U11737 (N_11737,N_10713,N_10760);
nand U11738 (N_11738,N_10765,N_11178);
xnor U11739 (N_11739,N_11177,N_10658);
xnor U11740 (N_11740,N_10443,N_11167);
xnor U11741 (N_11741,N_11177,N_11077);
xnor U11742 (N_11742,N_10600,N_10748);
nor U11743 (N_11743,N_10655,N_10712);
or U11744 (N_11744,N_10976,N_10825);
nand U11745 (N_11745,N_10955,N_10925);
or U11746 (N_11746,N_10880,N_10844);
nand U11747 (N_11747,N_10405,N_10807);
or U11748 (N_11748,N_10424,N_10975);
xnor U11749 (N_11749,N_10482,N_11154);
nand U11750 (N_11750,N_11036,N_10611);
nor U11751 (N_11751,N_10732,N_10718);
nand U11752 (N_11752,N_10574,N_10801);
or U11753 (N_11753,N_10751,N_10877);
or U11754 (N_11754,N_10979,N_10879);
nor U11755 (N_11755,N_10685,N_10494);
and U11756 (N_11756,N_11175,N_10916);
nand U11757 (N_11757,N_11130,N_11140);
xor U11758 (N_11758,N_10609,N_10768);
and U11759 (N_11759,N_10930,N_10932);
and U11760 (N_11760,N_11138,N_11175);
nand U11761 (N_11761,N_11180,N_10740);
nand U11762 (N_11762,N_10439,N_10597);
or U11763 (N_11763,N_11081,N_10846);
xnor U11764 (N_11764,N_10505,N_10864);
xor U11765 (N_11765,N_11193,N_10554);
nand U11766 (N_11766,N_11040,N_10646);
or U11767 (N_11767,N_10866,N_11174);
nand U11768 (N_11768,N_10981,N_10953);
xnor U11769 (N_11769,N_10682,N_10739);
xnor U11770 (N_11770,N_10488,N_10931);
and U11771 (N_11771,N_10424,N_10743);
nor U11772 (N_11772,N_10675,N_10945);
nand U11773 (N_11773,N_10833,N_10609);
xor U11774 (N_11774,N_11061,N_10415);
nand U11775 (N_11775,N_10565,N_10666);
nor U11776 (N_11776,N_10461,N_10785);
and U11777 (N_11777,N_10985,N_11014);
or U11778 (N_11778,N_10857,N_10433);
nor U11779 (N_11779,N_10579,N_10442);
nor U11780 (N_11780,N_11038,N_10726);
nor U11781 (N_11781,N_10855,N_11176);
xor U11782 (N_11782,N_11141,N_10416);
xor U11783 (N_11783,N_10578,N_11012);
and U11784 (N_11784,N_10722,N_10503);
xnor U11785 (N_11785,N_10965,N_10661);
or U11786 (N_11786,N_10762,N_10455);
nor U11787 (N_11787,N_10856,N_10613);
and U11788 (N_11788,N_10998,N_10541);
or U11789 (N_11789,N_10734,N_10705);
nor U11790 (N_11790,N_10462,N_10977);
and U11791 (N_11791,N_10432,N_10791);
or U11792 (N_11792,N_11052,N_10941);
or U11793 (N_11793,N_11108,N_10867);
nor U11794 (N_11794,N_11133,N_10671);
or U11795 (N_11795,N_11160,N_10813);
nand U11796 (N_11796,N_11070,N_11178);
and U11797 (N_11797,N_10570,N_11089);
xor U11798 (N_11798,N_10410,N_10485);
or U11799 (N_11799,N_10511,N_11057);
xor U11800 (N_11800,N_10578,N_10728);
or U11801 (N_11801,N_10558,N_10404);
and U11802 (N_11802,N_11089,N_10697);
nand U11803 (N_11803,N_10757,N_10908);
xor U11804 (N_11804,N_10662,N_10538);
and U11805 (N_11805,N_11082,N_11176);
and U11806 (N_11806,N_11023,N_10950);
nor U11807 (N_11807,N_10932,N_10575);
xnor U11808 (N_11808,N_10602,N_10922);
xnor U11809 (N_11809,N_10930,N_11010);
nand U11810 (N_11810,N_11018,N_10508);
nor U11811 (N_11811,N_10984,N_10579);
xnor U11812 (N_11812,N_10424,N_10663);
or U11813 (N_11813,N_10922,N_10687);
and U11814 (N_11814,N_11143,N_10763);
and U11815 (N_11815,N_10999,N_11061);
or U11816 (N_11816,N_11044,N_11131);
xnor U11817 (N_11817,N_10499,N_10808);
or U11818 (N_11818,N_10927,N_10768);
nor U11819 (N_11819,N_10791,N_10479);
or U11820 (N_11820,N_10821,N_10667);
nand U11821 (N_11821,N_10629,N_10865);
or U11822 (N_11822,N_10850,N_10888);
or U11823 (N_11823,N_11088,N_11100);
nor U11824 (N_11824,N_11065,N_10705);
or U11825 (N_11825,N_10519,N_10488);
xor U11826 (N_11826,N_10718,N_11174);
and U11827 (N_11827,N_10568,N_10999);
nand U11828 (N_11828,N_11043,N_10646);
nand U11829 (N_11829,N_10754,N_10743);
xnor U11830 (N_11830,N_10855,N_11065);
and U11831 (N_11831,N_10708,N_11103);
xnor U11832 (N_11832,N_10950,N_10464);
nand U11833 (N_11833,N_10957,N_10853);
xnor U11834 (N_11834,N_10682,N_11042);
or U11835 (N_11835,N_11176,N_10615);
xor U11836 (N_11836,N_10577,N_10503);
nand U11837 (N_11837,N_10631,N_11111);
xnor U11838 (N_11838,N_10712,N_10671);
or U11839 (N_11839,N_10427,N_10879);
and U11840 (N_11840,N_11154,N_10897);
nor U11841 (N_11841,N_10573,N_10653);
xor U11842 (N_11842,N_10603,N_10745);
nor U11843 (N_11843,N_10586,N_10844);
or U11844 (N_11844,N_10526,N_10758);
nand U11845 (N_11845,N_10511,N_10798);
nand U11846 (N_11846,N_10400,N_10988);
nand U11847 (N_11847,N_10405,N_10562);
and U11848 (N_11848,N_10412,N_10847);
nand U11849 (N_11849,N_10658,N_10700);
xor U11850 (N_11850,N_11121,N_11078);
and U11851 (N_11851,N_10995,N_10696);
xor U11852 (N_11852,N_10675,N_10876);
nor U11853 (N_11853,N_10594,N_10605);
or U11854 (N_11854,N_10978,N_10675);
xor U11855 (N_11855,N_10835,N_11121);
nor U11856 (N_11856,N_10637,N_10440);
nor U11857 (N_11857,N_11088,N_11011);
nor U11858 (N_11858,N_11054,N_11169);
nand U11859 (N_11859,N_11064,N_10659);
or U11860 (N_11860,N_10502,N_10490);
and U11861 (N_11861,N_10628,N_10581);
and U11862 (N_11862,N_10786,N_10471);
or U11863 (N_11863,N_10663,N_10632);
nor U11864 (N_11864,N_10494,N_11176);
nand U11865 (N_11865,N_10603,N_10874);
nor U11866 (N_11866,N_11112,N_10781);
nor U11867 (N_11867,N_10789,N_10911);
xor U11868 (N_11868,N_10558,N_10679);
and U11869 (N_11869,N_10896,N_10970);
and U11870 (N_11870,N_10579,N_10695);
and U11871 (N_11871,N_10999,N_10527);
and U11872 (N_11872,N_10887,N_10574);
and U11873 (N_11873,N_10979,N_10889);
and U11874 (N_11874,N_10812,N_10692);
nand U11875 (N_11875,N_10664,N_10667);
nor U11876 (N_11876,N_10843,N_10416);
or U11877 (N_11877,N_11123,N_11115);
or U11878 (N_11878,N_11161,N_10506);
and U11879 (N_11879,N_10792,N_10403);
nor U11880 (N_11880,N_10686,N_10531);
nand U11881 (N_11881,N_11019,N_10490);
xor U11882 (N_11882,N_10669,N_10865);
nor U11883 (N_11883,N_10553,N_11167);
nand U11884 (N_11884,N_11122,N_10527);
xnor U11885 (N_11885,N_11127,N_10476);
nand U11886 (N_11886,N_11016,N_10883);
nor U11887 (N_11887,N_10538,N_10574);
xnor U11888 (N_11888,N_10913,N_10424);
or U11889 (N_11889,N_11181,N_10983);
and U11890 (N_11890,N_10505,N_10511);
nand U11891 (N_11891,N_11152,N_10610);
xor U11892 (N_11892,N_11040,N_10763);
nor U11893 (N_11893,N_10683,N_10881);
and U11894 (N_11894,N_11059,N_10825);
or U11895 (N_11895,N_10533,N_10517);
and U11896 (N_11896,N_11093,N_10432);
or U11897 (N_11897,N_10611,N_10695);
or U11898 (N_11898,N_10895,N_10804);
and U11899 (N_11899,N_10626,N_10556);
or U11900 (N_11900,N_11162,N_10775);
xnor U11901 (N_11901,N_11145,N_11118);
and U11902 (N_11902,N_10588,N_10779);
xor U11903 (N_11903,N_10960,N_10427);
or U11904 (N_11904,N_10741,N_11040);
xor U11905 (N_11905,N_10704,N_10692);
or U11906 (N_11906,N_11143,N_10809);
nor U11907 (N_11907,N_10878,N_11026);
xnor U11908 (N_11908,N_11185,N_10944);
or U11909 (N_11909,N_10893,N_10440);
xor U11910 (N_11910,N_11057,N_11089);
nand U11911 (N_11911,N_10479,N_10860);
nand U11912 (N_11912,N_10489,N_11144);
nor U11913 (N_11913,N_10871,N_11028);
nand U11914 (N_11914,N_11169,N_10913);
or U11915 (N_11915,N_10691,N_10666);
and U11916 (N_11916,N_10496,N_10904);
or U11917 (N_11917,N_10434,N_10508);
xnor U11918 (N_11918,N_10747,N_10564);
nor U11919 (N_11919,N_10580,N_10909);
nand U11920 (N_11920,N_10654,N_10820);
and U11921 (N_11921,N_11167,N_11052);
xor U11922 (N_11922,N_10980,N_10580);
nand U11923 (N_11923,N_10785,N_11199);
nor U11924 (N_11924,N_11118,N_10747);
nand U11925 (N_11925,N_11040,N_10824);
and U11926 (N_11926,N_10665,N_11170);
and U11927 (N_11927,N_10656,N_11009);
or U11928 (N_11928,N_11113,N_10443);
nand U11929 (N_11929,N_10651,N_10483);
or U11930 (N_11930,N_10924,N_11046);
and U11931 (N_11931,N_10593,N_10517);
and U11932 (N_11932,N_10448,N_11129);
xnor U11933 (N_11933,N_11164,N_11123);
nand U11934 (N_11934,N_10742,N_10731);
nand U11935 (N_11935,N_11197,N_11143);
nand U11936 (N_11936,N_10867,N_10858);
nor U11937 (N_11937,N_11060,N_10761);
or U11938 (N_11938,N_10985,N_11183);
and U11939 (N_11939,N_11017,N_10658);
and U11940 (N_11940,N_10719,N_10663);
nand U11941 (N_11941,N_10790,N_11118);
xnor U11942 (N_11942,N_11198,N_10976);
xor U11943 (N_11943,N_10977,N_10505);
or U11944 (N_11944,N_10994,N_10599);
xor U11945 (N_11945,N_10818,N_10601);
nor U11946 (N_11946,N_10993,N_10966);
nor U11947 (N_11947,N_10950,N_10672);
nor U11948 (N_11948,N_10847,N_10584);
xnor U11949 (N_11949,N_11094,N_10631);
xnor U11950 (N_11950,N_10794,N_10631);
and U11951 (N_11951,N_11136,N_10541);
or U11952 (N_11952,N_10940,N_10410);
and U11953 (N_11953,N_11089,N_10586);
nor U11954 (N_11954,N_10816,N_10743);
nand U11955 (N_11955,N_11159,N_10954);
or U11956 (N_11956,N_11051,N_10981);
xnor U11957 (N_11957,N_11122,N_10879);
and U11958 (N_11958,N_11069,N_11035);
and U11959 (N_11959,N_11117,N_10621);
and U11960 (N_11960,N_10491,N_10842);
and U11961 (N_11961,N_10898,N_10523);
nand U11962 (N_11962,N_10818,N_10693);
nor U11963 (N_11963,N_10936,N_10553);
or U11964 (N_11964,N_10602,N_10657);
nor U11965 (N_11965,N_10550,N_10628);
nand U11966 (N_11966,N_10751,N_11184);
nand U11967 (N_11967,N_10673,N_10603);
nand U11968 (N_11968,N_10962,N_10861);
nor U11969 (N_11969,N_11054,N_10677);
xor U11970 (N_11970,N_10430,N_10899);
nor U11971 (N_11971,N_10847,N_11160);
or U11972 (N_11972,N_10820,N_11003);
xnor U11973 (N_11973,N_11190,N_11069);
nor U11974 (N_11974,N_11176,N_10868);
xnor U11975 (N_11975,N_10579,N_10895);
or U11976 (N_11976,N_10582,N_11111);
or U11977 (N_11977,N_10507,N_10900);
xor U11978 (N_11978,N_10863,N_11105);
and U11979 (N_11979,N_10786,N_10693);
and U11980 (N_11980,N_11042,N_10854);
nor U11981 (N_11981,N_10956,N_10900);
xnor U11982 (N_11982,N_10780,N_10427);
or U11983 (N_11983,N_10911,N_10769);
nand U11984 (N_11984,N_11023,N_10429);
xor U11985 (N_11985,N_11086,N_10712);
or U11986 (N_11986,N_10892,N_10549);
and U11987 (N_11987,N_10423,N_11032);
xor U11988 (N_11988,N_10901,N_10532);
xnor U11989 (N_11989,N_11188,N_10473);
nor U11990 (N_11990,N_10567,N_10739);
or U11991 (N_11991,N_11134,N_10764);
and U11992 (N_11992,N_10800,N_10538);
and U11993 (N_11993,N_10659,N_10492);
and U11994 (N_11994,N_10949,N_10722);
nand U11995 (N_11995,N_10685,N_10472);
or U11996 (N_11996,N_10513,N_10452);
nor U11997 (N_11997,N_10815,N_10913);
nor U11998 (N_11998,N_10948,N_10607);
xnor U11999 (N_11999,N_10709,N_10823);
nand U12000 (N_12000,N_11822,N_11551);
nor U12001 (N_12001,N_11695,N_11403);
or U12002 (N_12002,N_11397,N_11210);
or U12003 (N_12003,N_11703,N_11337);
nand U12004 (N_12004,N_11662,N_11277);
xor U12005 (N_12005,N_11728,N_11326);
and U12006 (N_12006,N_11531,N_11498);
and U12007 (N_12007,N_11992,N_11386);
nand U12008 (N_12008,N_11751,N_11730);
nand U12009 (N_12009,N_11886,N_11368);
and U12010 (N_12010,N_11311,N_11316);
and U12011 (N_12011,N_11793,N_11998);
and U12012 (N_12012,N_11877,N_11529);
nand U12013 (N_12013,N_11661,N_11660);
nand U12014 (N_12014,N_11307,N_11925);
nand U12015 (N_12015,N_11562,N_11421);
or U12016 (N_12016,N_11530,N_11799);
nand U12017 (N_12017,N_11617,N_11907);
or U12018 (N_12018,N_11821,N_11991);
xnor U12019 (N_12019,N_11605,N_11534);
xnor U12020 (N_12020,N_11521,N_11564);
or U12021 (N_12021,N_11591,N_11910);
xor U12022 (N_12022,N_11739,N_11758);
nand U12023 (N_12023,N_11801,N_11988);
or U12024 (N_12024,N_11688,N_11699);
nand U12025 (N_12025,N_11652,N_11327);
or U12026 (N_12026,N_11610,N_11207);
nand U12027 (N_12027,N_11537,N_11310);
or U12028 (N_12028,N_11686,N_11709);
xnor U12029 (N_12029,N_11441,N_11352);
nand U12030 (N_12030,N_11382,N_11852);
xnor U12031 (N_12031,N_11631,N_11510);
xnor U12032 (N_12032,N_11663,N_11724);
and U12033 (N_12033,N_11766,N_11477);
nor U12034 (N_12034,N_11355,N_11653);
nor U12035 (N_12035,N_11609,N_11476);
xnor U12036 (N_12036,N_11262,N_11524);
xnor U12037 (N_12037,N_11283,N_11772);
and U12038 (N_12038,N_11305,N_11978);
nand U12039 (N_12039,N_11559,N_11501);
nor U12040 (N_12040,N_11243,N_11571);
nor U12041 (N_12041,N_11471,N_11220);
xnor U12042 (N_12042,N_11595,N_11425);
and U12043 (N_12043,N_11712,N_11456);
xnor U12044 (N_12044,N_11224,N_11366);
nor U12045 (N_12045,N_11388,N_11820);
and U12046 (N_12046,N_11225,N_11912);
and U12047 (N_12047,N_11648,N_11721);
and U12048 (N_12048,N_11955,N_11216);
xnor U12049 (N_12049,N_11223,N_11764);
and U12050 (N_12050,N_11841,N_11768);
and U12051 (N_12051,N_11645,N_11936);
and U12052 (N_12052,N_11584,N_11463);
xor U12053 (N_12053,N_11902,N_11411);
and U12054 (N_12054,N_11752,N_11851);
xnor U12055 (N_12055,N_11965,N_11295);
xnor U12056 (N_12056,N_11757,N_11573);
xnor U12057 (N_12057,N_11457,N_11694);
nand U12058 (N_12058,N_11987,N_11585);
nand U12059 (N_12059,N_11565,N_11911);
nor U12060 (N_12060,N_11581,N_11480);
nand U12061 (N_12061,N_11373,N_11452);
and U12062 (N_12062,N_11487,N_11578);
or U12063 (N_12063,N_11726,N_11794);
nand U12064 (N_12064,N_11667,N_11825);
and U12065 (N_12065,N_11989,N_11824);
nand U12066 (N_12066,N_11299,N_11509);
and U12067 (N_12067,N_11418,N_11336);
nor U12068 (N_12068,N_11702,N_11738);
nor U12069 (N_12069,N_11906,N_11428);
xor U12070 (N_12070,N_11865,N_11209);
and U12071 (N_12071,N_11658,N_11389);
nor U12072 (N_12072,N_11974,N_11287);
or U12073 (N_12073,N_11933,N_11362);
nor U12074 (N_12074,N_11830,N_11265);
and U12075 (N_12075,N_11560,N_11218);
nand U12076 (N_12076,N_11996,N_11689);
nand U12077 (N_12077,N_11908,N_11475);
nor U12078 (N_12078,N_11878,N_11632);
and U12079 (N_12079,N_11438,N_11448);
nand U12080 (N_12080,N_11748,N_11629);
or U12081 (N_12081,N_11611,N_11928);
nor U12082 (N_12082,N_11783,N_11413);
nor U12083 (N_12083,N_11409,N_11672);
nand U12084 (N_12084,N_11599,N_11592);
and U12085 (N_12085,N_11485,N_11231);
nor U12086 (N_12086,N_11325,N_11508);
nand U12087 (N_12087,N_11575,N_11395);
or U12088 (N_12088,N_11453,N_11969);
nand U12089 (N_12089,N_11419,N_11634);
xnor U12090 (N_12090,N_11767,N_11993);
nand U12091 (N_12091,N_11788,N_11954);
xnor U12092 (N_12092,N_11696,N_11802);
nand U12093 (N_12093,N_11710,N_11889);
or U12094 (N_12094,N_11687,N_11205);
xor U12095 (N_12095,N_11486,N_11491);
nand U12096 (N_12096,N_11217,N_11249);
nand U12097 (N_12097,N_11750,N_11882);
nand U12098 (N_12098,N_11370,N_11725);
nand U12099 (N_12099,N_11246,N_11885);
nand U12100 (N_12100,N_11503,N_11619);
nor U12101 (N_12101,N_11839,N_11522);
nand U12102 (N_12102,N_11532,N_11828);
or U12103 (N_12103,N_11698,N_11950);
nor U12104 (N_12104,N_11365,N_11536);
or U12105 (N_12105,N_11895,N_11741);
nand U12106 (N_12106,N_11742,N_11898);
xor U12107 (N_12107,N_11240,N_11673);
xnor U12108 (N_12108,N_11615,N_11567);
or U12109 (N_12109,N_11313,N_11601);
and U12110 (N_12110,N_11525,N_11347);
xnor U12111 (N_12111,N_11319,N_11314);
nand U12112 (N_12112,N_11871,N_11637);
xor U12113 (N_12113,N_11659,N_11761);
and U12114 (N_12114,N_11228,N_11778);
nand U12115 (N_12115,N_11817,N_11588);
xnor U12116 (N_12116,N_11855,N_11398);
and U12117 (N_12117,N_11374,N_11780);
or U12118 (N_12118,N_11346,N_11893);
xnor U12119 (N_12119,N_11221,N_11986);
xnor U12120 (N_12120,N_11832,N_11940);
and U12121 (N_12121,N_11809,N_11250);
nor U12122 (N_12122,N_11460,N_11884);
nand U12123 (N_12123,N_11372,N_11546);
or U12124 (N_12124,N_11765,N_11704);
xnor U12125 (N_12125,N_11754,N_11396);
or U12126 (N_12126,N_11499,N_11812);
and U12127 (N_12127,N_11665,N_11717);
xnor U12128 (N_12128,N_11434,N_11932);
nand U12129 (N_12129,N_11384,N_11782);
nor U12130 (N_12130,N_11879,N_11201);
xor U12131 (N_12131,N_11269,N_11496);
or U12132 (N_12132,N_11935,N_11523);
and U12133 (N_12133,N_11539,N_11826);
nor U12134 (N_12134,N_11737,N_11789);
nor U12135 (N_12135,N_11437,N_11720);
nor U12136 (N_12136,N_11880,N_11268);
or U12137 (N_12137,N_11553,N_11713);
and U12138 (N_12138,N_11488,N_11735);
nor U12139 (N_12139,N_11756,N_11306);
or U12140 (N_12140,N_11233,N_11563);
nor U12141 (N_12141,N_11278,N_11469);
nor U12142 (N_12142,N_11492,N_11528);
nand U12143 (N_12143,N_11543,N_11414);
and U12144 (N_12144,N_11834,N_11763);
or U12145 (N_12145,N_11641,N_11494);
and U12146 (N_12146,N_11358,N_11837);
or U12147 (N_12147,N_11323,N_11813);
xnor U12148 (N_12148,N_11729,N_11308);
or U12149 (N_12149,N_11359,N_11232);
and U12150 (N_12150,N_11784,N_11569);
nor U12151 (N_12151,N_11391,N_11387);
nand U12152 (N_12152,N_11977,N_11442);
nand U12153 (N_12153,N_11867,N_11716);
nand U12154 (N_12154,N_11850,N_11612);
nor U12155 (N_12155,N_11861,N_11241);
xnor U12156 (N_12156,N_11651,N_11222);
or U12157 (N_12157,N_11429,N_11275);
xnor U12158 (N_12158,N_11415,N_11598);
nand U12159 (N_12159,N_11840,N_11961);
and U12160 (N_12160,N_11819,N_11271);
xor U12161 (N_12161,N_11806,N_11844);
nand U12162 (N_12162,N_11257,N_11876);
nor U12163 (N_12163,N_11800,N_11797);
nand U12164 (N_12164,N_11666,N_11450);
nand U12165 (N_12165,N_11506,N_11516);
xor U12166 (N_12166,N_11733,N_11743);
and U12167 (N_12167,N_11924,N_11482);
or U12168 (N_12168,N_11623,N_11859);
or U12169 (N_12169,N_11332,N_11613);
nor U12170 (N_12170,N_11557,N_11245);
and U12171 (N_12171,N_11848,N_11478);
xnor U12172 (N_12172,N_11315,N_11237);
nand U12173 (N_12173,N_11891,N_11625);
nor U12174 (N_12174,N_11502,N_11962);
nand U12175 (N_12175,N_11994,N_11943);
nand U12176 (N_12176,N_11272,N_11206);
xnor U12177 (N_12177,N_11676,N_11863);
xor U12178 (N_12178,N_11862,N_11566);
nand U12179 (N_12179,N_11357,N_11596);
and U12180 (N_12180,N_11416,N_11281);
nor U12181 (N_12181,N_11390,N_11650);
xnor U12182 (N_12182,N_11439,N_11309);
or U12183 (N_12183,N_11552,N_11402);
xnor U12184 (N_12184,N_11608,N_11540);
nand U12185 (N_12185,N_11646,N_11976);
and U12186 (N_12186,N_11883,N_11816);
nand U12187 (N_12187,N_11946,N_11378);
nor U12188 (N_12188,N_11999,N_11483);
xor U12189 (N_12189,N_11538,N_11638);
xor U12190 (N_12190,N_11706,N_11740);
xor U12191 (N_12191,N_11777,N_11443);
xor U12192 (N_12192,N_11636,N_11948);
nor U12193 (N_12193,N_11293,N_11680);
xor U12194 (N_12194,N_11776,N_11353);
xor U12195 (N_12195,N_11296,N_11270);
nand U12196 (N_12196,N_11679,N_11918);
and U12197 (N_12197,N_11845,N_11375);
or U12198 (N_12198,N_11512,N_11493);
nand U12199 (N_12199,N_11526,N_11732);
nand U12200 (N_12200,N_11236,N_11618);
nand U12201 (N_12201,N_11715,N_11258);
or U12202 (N_12202,N_11334,N_11602);
xor U12203 (N_12203,N_11484,N_11200);
xor U12204 (N_12204,N_11997,N_11410);
or U12205 (N_12205,N_11838,N_11371);
and U12206 (N_12206,N_11843,N_11723);
and U12207 (N_12207,N_11892,N_11234);
nor U12208 (N_12208,N_11670,N_11628);
nor U12209 (N_12209,N_11298,N_11980);
nand U12210 (N_12210,N_11970,N_11586);
nor U12211 (N_12211,N_11520,N_11656);
or U12212 (N_12212,N_11343,N_11280);
and U12213 (N_12213,N_11284,N_11968);
and U12214 (N_12214,N_11490,N_11771);
and U12215 (N_12215,N_11896,N_11995);
nand U12216 (N_12216,N_11407,N_11669);
and U12217 (N_12217,N_11930,N_11919);
and U12218 (N_12218,N_11677,N_11929);
nand U12219 (N_12219,N_11692,N_11517);
or U12220 (N_12220,N_11700,N_11266);
nor U12221 (N_12221,N_11481,N_11835);
xnor U12222 (N_12222,N_11412,N_11921);
and U12223 (N_12223,N_11972,N_11909);
and U12224 (N_12224,N_11630,N_11681);
nand U12225 (N_12225,N_11282,N_11582);
xnor U12226 (N_12226,N_11914,N_11810);
nand U12227 (N_12227,N_11213,N_11320);
nand U12228 (N_12228,N_11208,N_11811);
xor U12229 (N_12229,N_11519,N_11926);
nor U12230 (N_12230,N_11983,N_11626);
xnor U12231 (N_12231,N_11489,N_11408);
xnor U12232 (N_12232,N_11202,N_11708);
or U12233 (N_12233,N_11836,N_11392);
xnor U12234 (N_12234,N_11444,N_11760);
or U12235 (N_12235,N_11545,N_11682);
xnor U12236 (N_12236,N_11555,N_11734);
or U12237 (N_12237,N_11787,N_11576);
and U12238 (N_12238,N_11714,N_11736);
nor U12239 (N_12239,N_11937,N_11558);
nand U12240 (N_12240,N_11420,N_11860);
nor U12241 (N_12241,N_11939,N_11297);
and U12242 (N_12242,N_11866,N_11285);
and U12243 (N_12243,N_11430,N_11561);
nor U12244 (N_12244,N_11317,N_11356);
nor U12245 (N_12245,N_11785,N_11360);
or U12246 (N_12246,N_11577,N_11746);
xor U12247 (N_12247,N_11341,N_11973);
nand U12248 (N_12248,N_11400,N_11322);
and U12249 (N_12249,N_11773,N_11823);
nand U12250 (N_12250,N_11248,N_11711);
or U12251 (N_12251,N_11333,N_11624);
nand U12252 (N_12252,N_11255,N_11869);
or U12253 (N_12253,N_11684,N_11473);
and U12254 (N_12254,N_11344,N_11671);
nor U12255 (N_12255,N_11324,N_11547);
nor U12256 (N_12256,N_11639,N_11535);
or U12257 (N_12257,N_11881,N_11235);
xnor U12258 (N_12258,N_11905,N_11229);
or U12259 (N_12259,N_11796,N_11474);
or U12260 (N_12260,N_11781,N_11899);
nor U12261 (N_12261,N_11424,N_11513);
and U12262 (N_12262,N_11300,N_11468);
and U12263 (N_12263,N_11640,N_11915);
nor U12264 (N_12264,N_11616,N_11570);
xnor U12265 (N_12265,N_11204,N_11459);
nor U12266 (N_12266,N_11791,N_11829);
nand U12267 (N_12267,N_11417,N_11447);
nand U12268 (N_12268,N_11274,N_11288);
xnor U12269 (N_12269,N_11853,N_11927);
nand U12270 (N_12270,N_11900,N_11589);
and U12271 (N_12271,N_11505,N_11807);
nand U12272 (N_12272,N_11380,N_11244);
nor U12273 (N_12273,N_11227,N_11685);
nor U12274 (N_12274,N_11649,N_11583);
or U12275 (N_12275,N_11544,N_11590);
xnor U12276 (N_12276,N_11431,N_11574);
and U12277 (N_12277,N_11399,N_11975);
and U12278 (N_12278,N_11958,N_11887);
xor U12279 (N_12279,N_11707,N_11495);
and U12280 (N_12280,N_11267,N_11971);
and U12281 (N_12281,N_11461,N_11931);
nand U12282 (N_12282,N_11635,N_11597);
xnor U12283 (N_12283,N_11833,N_11226);
or U12284 (N_12284,N_11814,N_11302);
nand U12285 (N_12285,N_11642,N_11633);
nor U12286 (N_12286,N_11759,N_11423);
nand U12287 (N_12287,N_11620,N_11956);
nand U12288 (N_12288,N_11470,N_11913);
or U12289 (N_12289,N_11916,N_11705);
nand U12290 (N_12290,N_11697,N_11361);
or U12291 (N_12291,N_11579,N_11622);
and U12292 (N_12292,N_11500,N_11903);
xnor U12293 (N_12293,N_11643,N_11215);
nand U12294 (N_12294,N_11247,N_11875);
nor U12295 (N_12295,N_11321,N_11960);
and U12296 (N_12296,N_11379,N_11847);
and U12297 (N_12297,N_11944,N_11541);
xor U12298 (N_12298,N_11655,N_11897);
and U12299 (N_12299,N_11668,N_11345);
nor U12300 (N_12300,N_11718,N_11792);
xnor U12301 (N_12301,N_11294,N_11449);
xnor U12302 (N_12302,N_11849,N_11518);
nor U12303 (N_12303,N_11422,N_11291);
nand U12304 (N_12304,N_11259,N_11831);
or U12305 (N_12305,N_11264,N_11815);
xnor U12306 (N_12306,N_11394,N_11279);
xnor U12307 (N_12307,N_11945,N_11982);
nand U12308 (N_12308,N_11846,N_11693);
nand U12309 (N_12309,N_11230,N_11253);
or U12310 (N_12310,N_11458,N_11727);
nor U12311 (N_12311,N_11464,N_11856);
nand U12312 (N_12312,N_11339,N_11330);
or U12313 (N_12313,N_11774,N_11312);
and U12314 (N_12314,N_11239,N_11568);
or U12315 (N_12315,N_11304,N_11719);
xnor U12316 (N_12316,N_11857,N_11938);
and U12317 (N_12317,N_11864,N_11286);
and U12318 (N_12318,N_11678,N_11318);
nor U12319 (N_12319,N_11404,N_11804);
and U12320 (N_12320,N_11533,N_11479);
or U12321 (N_12321,N_11369,N_11606);
nand U12322 (N_12322,N_11260,N_11657);
xnor U12323 (N_12323,N_11901,N_11888);
and U12324 (N_12324,N_11383,N_11446);
or U12325 (N_12325,N_11979,N_11904);
nand U12326 (N_12326,N_11762,N_11769);
xor U12327 (N_12327,N_11550,N_11587);
nand U12328 (N_12328,N_11363,N_11644);
and U12329 (N_12329,N_11385,N_11290);
xnor U12330 (N_12330,N_11301,N_11462);
nand U12331 (N_12331,N_11964,N_11467);
nor U12332 (N_12332,N_11941,N_11858);
nand U12333 (N_12333,N_11572,N_11211);
or U12334 (N_12334,N_11934,N_11674);
or U12335 (N_12335,N_11947,N_11798);
nand U12336 (N_12336,N_11894,N_11614);
nor U12337 (N_12337,N_11252,N_11744);
and U12338 (N_12338,N_11349,N_11242);
nand U12339 (N_12339,N_11406,N_11753);
or U12340 (N_12340,N_11967,N_11377);
xnor U12341 (N_12341,N_11515,N_11854);
nor U12342 (N_12342,N_11920,N_11542);
and U12343 (N_12343,N_11445,N_11219);
or U12344 (N_12344,N_11342,N_11465);
xnor U12345 (N_12345,N_11440,N_11691);
and U12346 (N_12346,N_11786,N_11790);
or U12347 (N_12347,N_11393,N_11604);
xnor U12348 (N_12348,N_11451,N_11923);
and U12349 (N_12349,N_11556,N_11952);
nand U12350 (N_12350,N_11472,N_11507);
nor U12351 (N_12351,N_11335,N_11214);
or U12352 (N_12352,N_11580,N_11647);
nand U12353 (N_12353,N_11212,N_11984);
and U12354 (N_12354,N_11329,N_11607);
xor U12355 (N_12355,N_11949,N_11870);
nor U12356 (N_12356,N_11364,N_11654);
or U12357 (N_12357,N_11873,N_11548);
and U12358 (N_12358,N_11755,N_11747);
or U12359 (N_12359,N_11432,N_11354);
nand U12360 (N_12360,N_11435,N_11966);
nor U12361 (N_12361,N_11436,N_11405);
xor U12362 (N_12362,N_11263,N_11455);
xnor U12363 (N_12363,N_11367,N_11514);
and U12364 (N_12364,N_11942,N_11276);
or U12365 (N_12365,N_11593,N_11292);
and U12366 (N_12366,N_11401,N_11527);
xor U12367 (N_12367,N_11985,N_11981);
xnor U12368 (N_12368,N_11251,N_11795);
and U12369 (N_12369,N_11600,N_11959);
or U12370 (N_12370,N_11427,N_11261);
xor U12371 (N_12371,N_11808,N_11348);
xnor U12372 (N_12372,N_11731,N_11957);
nor U12373 (N_12373,N_11504,N_11722);
nor U12374 (N_12374,N_11627,N_11426);
nand U12375 (N_12375,N_11842,N_11331);
nand U12376 (N_12376,N_11701,N_11818);
and U12377 (N_12377,N_11664,N_11683);
nand U12378 (N_12378,N_11803,N_11775);
xor U12379 (N_12379,N_11690,N_11745);
xnor U12380 (N_12380,N_11328,N_11963);
and U12381 (N_12381,N_11953,N_11594);
nor U12382 (N_12382,N_11497,N_11238);
and U12383 (N_12383,N_11827,N_11922);
xnor U12384 (N_12384,N_11433,N_11350);
nor U12385 (N_12385,N_11872,N_11951);
nand U12386 (N_12386,N_11805,N_11675);
and U12387 (N_12387,N_11303,N_11749);
or U12388 (N_12388,N_11549,N_11273);
xnor U12389 (N_12389,N_11603,N_11254);
or U12390 (N_12390,N_11381,N_11289);
xnor U12391 (N_12391,N_11466,N_11770);
nand U12392 (N_12392,N_11376,N_11890);
or U12393 (N_12393,N_11351,N_11990);
and U12394 (N_12394,N_11340,N_11917);
nor U12395 (N_12395,N_11554,N_11874);
xnor U12396 (N_12396,N_11779,N_11511);
or U12397 (N_12397,N_11868,N_11338);
and U12398 (N_12398,N_11454,N_11256);
nor U12399 (N_12399,N_11621,N_11203);
or U12400 (N_12400,N_11493,N_11225);
nand U12401 (N_12401,N_11367,N_11684);
and U12402 (N_12402,N_11418,N_11868);
nor U12403 (N_12403,N_11694,N_11664);
nand U12404 (N_12404,N_11321,N_11218);
or U12405 (N_12405,N_11885,N_11408);
or U12406 (N_12406,N_11889,N_11886);
xnor U12407 (N_12407,N_11791,N_11735);
or U12408 (N_12408,N_11895,N_11663);
nand U12409 (N_12409,N_11267,N_11213);
or U12410 (N_12410,N_11859,N_11955);
and U12411 (N_12411,N_11232,N_11955);
xor U12412 (N_12412,N_11336,N_11265);
and U12413 (N_12413,N_11642,N_11891);
nor U12414 (N_12414,N_11432,N_11716);
and U12415 (N_12415,N_11892,N_11927);
xnor U12416 (N_12416,N_11932,N_11821);
nor U12417 (N_12417,N_11543,N_11729);
and U12418 (N_12418,N_11644,N_11621);
or U12419 (N_12419,N_11712,N_11774);
nand U12420 (N_12420,N_11231,N_11736);
nand U12421 (N_12421,N_11666,N_11240);
nand U12422 (N_12422,N_11891,N_11757);
nor U12423 (N_12423,N_11276,N_11301);
nand U12424 (N_12424,N_11369,N_11465);
or U12425 (N_12425,N_11367,N_11528);
nor U12426 (N_12426,N_11387,N_11638);
or U12427 (N_12427,N_11943,N_11844);
xor U12428 (N_12428,N_11605,N_11862);
nand U12429 (N_12429,N_11620,N_11320);
xor U12430 (N_12430,N_11657,N_11697);
nand U12431 (N_12431,N_11990,N_11387);
and U12432 (N_12432,N_11567,N_11854);
or U12433 (N_12433,N_11373,N_11909);
nor U12434 (N_12434,N_11423,N_11319);
nor U12435 (N_12435,N_11230,N_11418);
or U12436 (N_12436,N_11341,N_11527);
nor U12437 (N_12437,N_11646,N_11947);
and U12438 (N_12438,N_11532,N_11400);
nand U12439 (N_12439,N_11725,N_11695);
nand U12440 (N_12440,N_11781,N_11723);
xor U12441 (N_12441,N_11243,N_11839);
and U12442 (N_12442,N_11309,N_11441);
xor U12443 (N_12443,N_11725,N_11971);
or U12444 (N_12444,N_11421,N_11949);
or U12445 (N_12445,N_11554,N_11883);
or U12446 (N_12446,N_11647,N_11492);
and U12447 (N_12447,N_11851,N_11607);
and U12448 (N_12448,N_11476,N_11343);
nor U12449 (N_12449,N_11935,N_11637);
and U12450 (N_12450,N_11263,N_11570);
xnor U12451 (N_12451,N_11599,N_11818);
or U12452 (N_12452,N_11799,N_11309);
nand U12453 (N_12453,N_11728,N_11717);
nand U12454 (N_12454,N_11229,N_11916);
or U12455 (N_12455,N_11713,N_11368);
nor U12456 (N_12456,N_11456,N_11400);
or U12457 (N_12457,N_11821,N_11691);
and U12458 (N_12458,N_11723,N_11969);
xnor U12459 (N_12459,N_11436,N_11309);
and U12460 (N_12460,N_11974,N_11690);
or U12461 (N_12461,N_11389,N_11759);
nor U12462 (N_12462,N_11535,N_11691);
or U12463 (N_12463,N_11654,N_11535);
nor U12464 (N_12464,N_11922,N_11416);
and U12465 (N_12465,N_11920,N_11948);
nor U12466 (N_12466,N_11397,N_11759);
xor U12467 (N_12467,N_11316,N_11277);
nand U12468 (N_12468,N_11854,N_11261);
and U12469 (N_12469,N_11371,N_11641);
or U12470 (N_12470,N_11939,N_11346);
or U12471 (N_12471,N_11518,N_11333);
or U12472 (N_12472,N_11583,N_11775);
or U12473 (N_12473,N_11593,N_11868);
and U12474 (N_12474,N_11509,N_11692);
or U12475 (N_12475,N_11555,N_11665);
nor U12476 (N_12476,N_11281,N_11407);
and U12477 (N_12477,N_11696,N_11941);
nor U12478 (N_12478,N_11438,N_11725);
and U12479 (N_12479,N_11414,N_11421);
nor U12480 (N_12480,N_11590,N_11295);
or U12481 (N_12481,N_11414,N_11651);
and U12482 (N_12482,N_11674,N_11517);
or U12483 (N_12483,N_11208,N_11789);
and U12484 (N_12484,N_11291,N_11660);
and U12485 (N_12485,N_11938,N_11988);
nor U12486 (N_12486,N_11438,N_11496);
nand U12487 (N_12487,N_11668,N_11250);
nand U12488 (N_12488,N_11535,N_11735);
xnor U12489 (N_12489,N_11810,N_11948);
or U12490 (N_12490,N_11397,N_11858);
nand U12491 (N_12491,N_11621,N_11875);
xnor U12492 (N_12492,N_11647,N_11499);
nor U12493 (N_12493,N_11477,N_11335);
nor U12494 (N_12494,N_11845,N_11228);
nand U12495 (N_12495,N_11416,N_11489);
nor U12496 (N_12496,N_11965,N_11637);
and U12497 (N_12497,N_11309,N_11325);
xor U12498 (N_12498,N_11701,N_11269);
and U12499 (N_12499,N_11412,N_11914);
or U12500 (N_12500,N_11745,N_11473);
nand U12501 (N_12501,N_11948,N_11491);
nor U12502 (N_12502,N_11866,N_11557);
and U12503 (N_12503,N_11823,N_11859);
nand U12504 (N_12504,N_11751,N_11363);
and U12505 (N_12505,N_11869,N_11726);
xnor U12506 (N_12506,N_11759,N_11889);
nor U12507 (N_12507,N_11214,N_11709);
nand U12508 (N_12508,N_11886,N_11474);
nand U12509 (N_12509,N_11487,N_11515);
or U12510 (N_12510,N_11255,N_11460);
or U12511 (N_12511,N_11924,N_11895);
nor U12512 (N_12512,N_11425,N_11981);
and U12513 (N_12513,N_11514,N_11458);
and U12514 (N_12514,N_11470,N_11330);
or U12515 (N_12515,N_11404,N_11889);
nor U12516 (N_12516,N_11585,N_11373);
xor U12517 (N_12517,N_11243,N_11206);
nand U12518 (N_12518,N_11813,N_11584);
nand U12519 (N_12519,N_11796,N_11833);
nor U12520 (N_12520,N_11617,N_11478);
xor U12521 (N_12521,N_11235,N_11460);
xor U12522 (N_12522,N_11387,N_11261);
or U12523 (N_12523,N_11705,N_11425);
nand U12524 (N_12524,N_11510,N_11227);
nand U12525 (N_12525,N_11623,N_11945);
and U12526 (N_12526,N_11764,N_11970);
or U12527 (N_12527,N_11661,N_11700);
nand U12528 (N_12528,N_11342,N_11513);
or U12529 (N_12529,N_11277,N_11566);
and U12530 (N_12530,N_11246,N_11770);
nand U12531 (N_12531,N_11729,N_11451);
nand U12532 (N_12532,N_11805,N_11379);
and U12533 (N_12533,N_11250,N_11772);
xnor U12534 (N_12534,N_11686,N_11921);
nor U12535 (N_12535,N_11841,N_11937);
nand U12536 (N_12536,N_11417,N_11340);
nand U12537 (N_12537,N_11493,N_11337);
nor U12538 (N_12538,N_11669,N_11322);
xor U12539 (N_12539,N_11771,N_11799);
nor U12540 (N_12540,N_11459,N_11702);
nand U12541 (N_12541,N_11587,N_11722);
and U12542 (N_12542,N_11278,N_11432);
nand U12543 (N_12543,N_11930,N_11317);
xnor U12544 (N_12544,N_11836,N_11884);
or U12545 (N_12545,N_11786,N_11884);
and U12546 (N_12546,N_11732,N_11485);
and U12547 (N_12547,N_11345,N_11932);
or U12548 (N_12548,N_11794,N_11743);
xor U12549 (N_12549,N_11955,N_11241);
and U12550 (N_12550,N_11295,N_11362);
nand U12551 (N_12551,N_11319,N_11299);
xnor U12552 (N_12552,N_11933,N_11713);
nor U12553 (N_12553,N_11288,N_11597);
nand U12554 (N_12554,N_11234,N_11784);
nor U12555 (N_12555,N_11649,N_11694);
or U12556 (N_12556,N_11220,N_11934);
nand U12557 (N_12557,N_11514,N_11379);
nor U12558 (N_12558,N_11535,N_11624);
and U12559 (N_12559,N_11411,N_11384);
and U12560 (N_12560,N_11297,N_11277);
nand U12561 (N_12561,N_11252,N_11702);
nand U12562 (N_12562,N_11702,N_11387);
or U12563 (N_12563,N_11258,N_11596);
or U12564 (N_12564,N_11554,N_11256);
nand U12565 (N_12565,N_11912,N_11790);
nor U12566 (N_12566,N_11905,N_11601);
nand U12567 (N_12567,N_11786,N_11958);
or U12568 (N_12568,N_11308,N_11995);
nand U12569 (N_12569,N_11339,N_11836);
nor U12570 (N_12570,N_11838,N_11503);
nor U12571 (N_12571,N_11403,N_11460);
nor U12572 (N_12572,N_11662,N_11394);
nand U12573 (N_12573,N_11906,N_11464);
xor U12574 (N_12574,N_11813,N_11840);
nor U12575 (N_12575,N_11409,N_11726);
and U12576 (N_12576,N_11371,N_11853);
nor U12577 (N_12577,N_11484,N_11356);
and U12578 (N_12578,N_11364,N_11333);
or U12579 (N_12579,N_11432,N_11979);
xor U12580 (N_12580,N_11892,N_11553);
or U12581 (N_12581,N_11595,N_11283);
xor U12582 (N_12582,N_11550,N_11325);
nand U12583 (N_12583,N_11423,N_11830);
and U12584 (N_12584,N_11318,N_11537);
nor U12585 (N_12585,N_11801,N_11726);
nand U12586 (N_12586,N_11239,N_11309);
and U12587 (N_12587,N_11742,N_11690);
xor U12588 (N_12588,N_11445,N_11907);
nor U12589 (N_12589,N_11973,N_11509);
nor U12590 (N_12590,N_11975,N_11976);
nand U12591 (N_12591,N_11394,N_11443);
nand U12592 (N_12592,N_11755,N_11298);
and U12593 (N_12593,N_11267,N_11765);
nor U12594 (N_12594,N_11280,N_11928);
or U12595 (N_12595,N_11803,N_11945);
nand U12596 (N_12596,N_11807,N_11753);
or U12597 (N_12597,N_11243,N_11663);
nor U12598 (N_12598,N_11374,N_11821);
xnor U12599 (N_12599,N_11426,N_11644);
or U12600 (N_12600,N_11351,N_11939);
or U12601 (N_12601,N_11571,N_11754);
and U12602 (N_12602,N_11704,N_11514);
or U12603 (N_12603,N_11353,N_11320);
or U12604 (N_12604,N_11381,N_11205);
or U12605 (N_12605,N_11554,N_11700);
or U12606 (N_12606,N_11333,N_11525);
nand U12607 (N_12607,N_11761,N_11479);
nor U12608 (N_12608,N_11931,N_11555);
nand U12609 (N_12609,N_11879,N_11410);
xnor U12610 (N_12610,N_11856,N_11387);
nor U12611 (N_12611,N_11889,N_11269);
nor U12612 (N_12612,N_11444,N_11800);
nor U12613 (N_12613,N_11794,N_11405);
nand U12614 (N_12614,N_11338,N_11515);
xor U12615 (N_12615,N_11893,N_11969);
nor U12616 (N_12616,N_11554,N_11870);
or U12617 (N_12617,N_11952,N_11674);
and U12618 (N_12618,N_11489,N_11413);
nor U12619 (N_12619,N_11306,N_11945);
xor U12620 (N_12620,N_11317,N_11762);
xor U12621 (N_12621,N_11952,N_11935);
nand U12622 (N_12622,N_11965,N_11595);
or U12623 (N_12623,N_11667,N_11834);
or U12624 (N_12624,N_11243,N_11360);
nand U12625 (N_12625,N_11357,N_11462);
or U12626 (N_12626,N_11955,N_11205);
or U12627 (N_12627,N_11266,N_11827);
nor U12628 (N_12628,N_11713,N_11739);
xor U12629 (N_12629,N_11323,N_11936);
nor U12630 (N_12630,N_11713,N_11842);
or U12631 (N_12631,N_11386,N_11909);
and U12632 (N_12632,N_11730,N_11295);
or U12633 (N_12633,N_11970,N_11675);
or U12634 (N_12634,N_11812,N_11462);
or U12635 (N_12635,N_11262,N_11303);
xnor U12636 (N_12636,N_11421,N_11408);
or U12637 (N_12637,N_11793,N_11744);
xor U12638 (N_12638,N_11485,N_11539);
nand U12639 (N_12639,N_11694,N_11656);
nor U12640 (N_12640,N_11665,N_11873);
xor U12641 (N_12641,N_11222,N_11452);
nor U12642 (N_12642,N_11365,N_11541);
nand U12643 (N_12643,N_11939,N_11899);
and U12644 (N_12644,N_11859,N_11316);
nor U12645 (N_12645,N_11788,N_11948);
xnor U12646 (N_12646,N_11605,N_11884);
nand U12647 (N_12647,N_11275,N_11203);
and U12648 (N_12648,N_11856,N_11785);
nor U12649 (N_12649,N_11357,N_11535);
xnor U12650 (N_12650,N_11213,N_11657);
xnor U12651 (N_12651,N_11982,N_11515);
nor U12652 (N_12652,N_11384,N_11790);
and U12653 (N_12653,N_11993,N_11826);
and U12654 (N_12654,N_11339,N_11817);
nor U12655 (N_12655,N_11821,N_11668);
xor U12656 (N_12656,N_11664,N_11845);
or U12657 (N_12657,N_11808,N_11668);
nand U12658 (N_12658,N_11304,N_11522);
or U12659 (N_12659,N_11619,N_11762);
or U12660 (N_12660,N_11716,N_11670);
nand U12661 (N_12661,N_11562,N_11607);
or U12662 (N_12662,N_11576,N_11389);
or U12663 (N_12663,N_11775,N_11451);
nor U12664 (N_12664,N_11239,N_11509);
nor U12665 (N_12665,N_11934,N_11943);
xnor U12666 (N_12666,N_11339,N_11215);
or U12667 (N_12667,N_11560,N_11379);
nor U12668 (N_12668,N_11201,N_11247);
nand U12669 (N_12669,N_11347,N_11527);
xnor U12670 (N_12670,N_11485,N_11647);
and U12671 (N_12671,N_11475,N_11944);
nand U12672 (N_12672,N_11486,N_11867);
or U12673 (N_12673,N_11721,N_11216);
nor U12674 (N_12674,N_11364,N_11407);
nand U12675 (N_12675,N_11868,N_11200);
and U12676 (N_12676,N_11609,N_11282);
nand U12677 (N_12677,N_11633,N_11526);
and U12678 (N_12678,N_11619,N_11499);
xnor U12679 (N_12679,N_11550,N_11515);
nor U12680 (N_12680,N_11766,N_11244);
or U12681 (N_12681,N_11866,N_11502);
and U12682 (N_12682,N_11511,N_11617);
xnor U12683 (N_12683,N_11465,N_11958);
or U12684 (N_12684,N_11999,N_11222);
or U12685 (N_12685,N_11817,N_11753);
nand U12686 (N_12686,N_11789,N_11911);
or U12687 (N_12687,N_11891,N_11743);
nand U12688 (N_12688,N_11897,N_11987);
and U12689 (N_12689,N_11912,N_11914);
nor U12690 (N_12690,N_11490,N_11688);
nand U12691 (N_12691,N_11822,N_11435);
or U12692 (N_12692,N_11675,N_11410);
or U12693 (N_12693,N_11722,N_11764);
nor U12694 (N_12694,N_11936,N_11358);
xor U12695 (N_12695,N_11634,N_11288);
nor U12696 (N_12696,N_11253,N_11591);
xor U12697 (N_12697,N_11747,N_11386);
nor U12698 (N_12698,N_11238,N_11718);
or U12699 (N_12699,N_11829,N_11692);
or U12700 (N_12700,N_11587,N_11215);
nand U12701 (N_12701,N_11778,N_11466);
nand U12702 (N_12702,N_11204,N_11484);
or U12703 (N_12703,N_11698,N_11864);
xnor U12704 (N_12704,N_11786,N_11534);
and U12705 (N_12705,N_11353,N_11873);
nor U12706 (N_12706,N_11771,N_11782);
xnor U12707 (N_12707,N_11791,N_11523);
and U12708 (N_12708,N_11902,N_11680);
nor U12709 (N_12709,N_11924,N_11551);
nand U12710 (N_12710,N_11508,N_11491);
xnor U12711 (N_12711,N_11900,N_11253);
and U12712 (N_12712,N_11392,N_11523);
nand U12713 (N_12713,N_11371,N_11859);
or U12714 (N_12714,N_11917,N_11426);
xnor U12715 (N_12715,N_11863,N_11920);
nand U12716 (N_12716,N_11939,N_11431);
or U12717 (N_12717,N_11997,N_11797);
and U12718 (N_12718,N_11768,N_11231);
and U12719 (N_12719,N_11456,N_11740);
xor U12720 (N_12720,N_11506,N_11719);
and U12721 (N_12721,N_11585,N_11879);
and U12722 (N_12722,N_11484,N_11726);
and U12723 (N_12723,N_11789,N_11879);
or U12724 (N_12724,N_11413,N_11444);
nand U12725 (N_12725,N_11873,N_11490);
or U12726 (N_12726,N_11615,N_11677);
or U12727 (N_12727,N_11775,N_11393);
xor U12728 (N_12728,N_11650,N_11685);
and U12729 (N_12729,N_11465,N_11428);
and U12730 (N_12730,N_11378,N_11494);
xnor U12731 (N_12731,N_11916,N_11569);
and U12732 (N_12732,N_11634,N_11638);
nand U12733 (N_12733,N_11751,N_11220);
nand U12734 (N_12734,N_11565,N_11841);
nand U12735 (N_12735,N_11288,N_11795);
nand U12736 (N_12736,N_11690,N_11652);
and U12737 (N_12737,N_11795,N_11201);
nand U12738 (N_12738,N_11533,N_11340);
or U12739 (N_12739,N_11607,N_11910);
xnor U12740 (N_12740,N_11680,N_11223);
xor U12741 (N_12741,N_11980,N_11331);
nor U12742 (N_12742,N_11493,N_11517);
and U12743 (N_12743,N_11840,N_11705);
nand U12744 (N_12744,N_11599,N_11306);
or U12745 (N_12745,N_11931,N_11626);
and U12746 (N_12746,N_11695,N_11474);
or U12747 (N_12747,N_11488,N_11716);
nor U12748 (N_12748,N_11878,N_11286);
xnor U12749 (N_12749,N_11766,N_11409);
xnor U12750 (N_12750,N_11578,N_11732);
nor U12751 (N_12751,N_11608,N_11677);
nand U12752 (N_12752,N_11324,N_11524);
and U12753 (N_12753,N_11692,N_11395);
nand U12754 (N_12754,N_11751,N_11365);
nor U12755 (N_12755,N_11650,N_11304);
xnor U12756 (N_12756,N_11805,N_11898);
nor U12757 (N_12757,N_11633,N_11607);
or U12758 (N_12758,N_11596,N_11294);
or U12759 (N_12759,N_11979,N_11959);
or U12760 (N_12760,N_11884,N_11264);
xor U12761 (N_12761,N_11480,N_11226);
xnor U12762 (N_12762,N_11554,N_11846);
xor U12763 (N_12763,N_11369,N_11649);
nor U12764 (N_12764,N_11240,N_11258);
nand U12765 (N_12765,N_11438,N_11372);
and U12766 (N_12766,N_11760,N_11239);
nor U12767 (N_12767,N_11605,N_11477);
nand U12768 (N_12768,N_11751,N_11207);
or U12769 (N_12769,N_11586,N_11296);
xor U12770 (N_12770,N_11359,N_11827);
or U12771 (N_12771,N_11296,N_11332);
or U12772 (N_12772,N_11328,N_11799);
or U12773 (N_12773,N_11232,N_11493);
nor U12774 (N_12774,N_11728,N_11408);
nor U12775 (N_12775,N_11621,N_11453);
xnor U12776 (N_12776,N_11464,N_11986);
xnor U12777 (N_12777,N_11804,N_11334);
xor U12778 (N_12778,N_11616,N_11490);
and U12779 (N_12779,N_11652,N_11441);
or U12780 (N_12780,N_11964,N_11814);
nor U12781 (N_12781,N_11295,N_11678);
or U12782 (N_12782,N_11731,N_11241);
or U12783 (N_12783,N_11387,N_11964);
nor U12784 (N_12784,N_11653,N_11252);
nand U12785 (N_12785,N_11525,N_11385);
xnor U12786 (N_12786,N_11297,N_11881);
xnor U12787 (N_12787,N_11751,N_11952);
xor U12788 (N_12788,N_11617,N_11324);
and U12789 (N_12789,N_11717,N_11721);
xor U12790 (N_12790,N_11641,N_11446);
or U12791 (N_12791,N_11325,N_11394);
and U12792 (N_12792,N_11506,N_11383);
nor U12793 (N_12793,N_11412,N_11811);
xnor U12794 (N_12794,N_11522,N_11620);
nor U12795 (N_12795,N_11909,N_11946);
and U12796 (N_12796,N_11741,N_11230);
nor U12797 (N_12797,N_11461,N_11517);
xor U12798 (N_12798,N_11967,N_11965);
nand U12799 (N_12799,N_11503,N_11655);
xnor U12800 (N_12800,N_12182,N_12678);
and U12801 (N_12801,N_12484,N_12190);
nand U12802 (N_12802,N_12193,N_12043);
or U12803 (N_12803,N_12077,N_12107);
nand U12804 (N_12804,N_12125,N_12168);
nand U12805 (N_12805,N_12628,N_12195);
and U12806 (N_12806,N_12401,N_12615);
xor U12807 (N_12807,N_12067,N_12511);
and U12808 (N_12808,N_12082,N_12778);
nand U12809 (N_12809,N_12706,N_12200);
or U12810 (N_12810,N_12186,N_12666);
nor U12811 (N_12811,N_12428,N_12126);
or U12812 (N_12812,N_12728,N_12655);
xor U12813 (N_12813,N_12269,N_12748);
or U12814 (N_12814,N_12400,N_12243);
nand U12815 (N_12815,N_12339,N_12736);
nand U12816 (N_12816,N_12048,N_12592);
and U12817 (N_12817,N_12493,N_12371);
nand U12818 (N_12818,N_12064,N_12535);
nor U12819 (N_12819,N_12157,N_12754);
xnor U12820 (N_12820,N_12453,N_12506);
and U12821 (N_12821,N_12264,N_12324);
and U12822 (N_12822,N_12317,N_12167);
and U12823 (N_12823,N_12263,N_12362);
nor U12824 (N_12824,N_12220,N_12268);
xor U12825 (N_12825,N_12236,N_12792);
and U12826 (N_12826,N_12071,N_12201);
nor U12827 (N_12827,N_12407,N_12292);
or U12828 (N_12828,N_12481,N_12596);
nand U12829 (N_12829,N_12288,N_12011);
nand U12830 (N_12830,N_12088,N_12644);
and U12831 (N_12831,N_12047,N_12630);
nor U12832 (N_12832,N_12121,N_12299);
nand U12833 (N_12833,N_12468,N_12408);
nor U12834 (N_12834,N_12562,N_12141);
nand U12835 (N_12835,N_12440,N_12625);
xnor U12836 (N_12836,N_12597,N_12189);
nand U12837 (N_12837,N_12540,N_12146);
and U12838 (N_12838,N_12433,N_12240);
xor U12839 (N_12839,N_12498,N_12724);
or U12840 (N_12840,N_12109,N_12721);
nor U12841 (N_12841,N_12756,N_12673);
nand U12842 (N_12842,N_12301,N_12789);
nor U12843 (N_12843,N_12609,N_12427);
xnor U12844 (N_12844,N_12524,N_12402);
and U12845 (N_12845,N_12656,N_12050);
nand U12846 (N_12846,N_12346,N_12367);
or U12847 (N_12847,N_12612,N_12760);
nor U12848 (N_12848,N_12160,N_12398);
nor U12849 (N_12849,N_12436,N_12210);
nand U12850 (N_12850,N_12403,N_12465);
or U12851 (N_12851,N_12782,N_12775);
nor U12852 (N_12852,N_12030,N_12318);
nor U12853 (N_12853,N_12514,N_12587);
xor U12854 (N_12854,N_12545,N_12649);
and U12855 (N_12855,N_12671,N_12265);
xor U12856 (N_12856,N_12595,N_12418);
or U12857 (N_12857,N_12567,N_12576);
xnor U12858 (N_12858,N_12308,N_12298);
nand U12859 (N_12859,N_12610,N_12623);
nor U12860 (N_12860,N_12151,N_12221);
nor U12861 (N_12861,N_12590,N_12320);
nand U12862 (N_12862,N_12283,N_12667);
or U12863 (N_12863,N_12501,N_12178);
nor U12864 (N_12864,N_12155,N_12002);
nor U12865 (N_12865,N_12310,N_12518);
xnor U12866 (N_12866,N_12335,N_12505);
or U12867 (N_12867,N_12380,N_12207);
or U12868 (N_12868,N_12499,N_12683);
or U12869 (N_12869,N_12139,N_12185);
and U12870 (N_12870,N_12619,N_12564);
and U12871 (N_12871,N_12555,N_12049);
nor U12872 (N_12872,N_12253,N_12276);
nor U12873 (N_12873,N_12357,N_12578);
and U12874 (N_12874,N_12381,N_12785);
xnor U12875 (N_12875,N_12244,N_12277);
xnor U12876 (N_12876,N_12726,N_12053);
and U12877 (N_12877,N_12313,N_12156);
nand U12878 (N_12878,N_12070,N_12718);
nand U12879 (N_12879,N_12003,N_12289);
xor U12880 (N_12880,N_12140,N_12122);
nor U12881 (N_12881,N_12568,N_12412);
nor U12882 (N_12882,N_12532,N_12584);
or U12883 (N_12883,N_12589,N_12503);
nand U12884 (N_12884,N_12231,N_12653);
nor U12885 (N_12885,N_12553,N_12163);
xnor U12886 (N_12886,N_12282,N_12687);
xor U12887 (N_12887,N_12795,N_12411);
or U12888 (N_12888,N_12725,N_12364);
nand U12889 (N_12889,N_12627,N_12600);
nand U12890 (N_12890,N_12039,N_12127);
nor U12891 (N_12891,N_12672,N_12267);
nand U12892 (N_12892,N_12252,N_12617);
xor U12893 (N_12893,N_12327,N_12159);
nor U12894 (N_12894,N_12311,N_12439);
nor U12895 (N_12895,N_12080,N_12478);
and U12896 (N_12896,N_12150,N_12684);
xor U12897 (N_12897,N_12316,N_12363);
xnor U12898 (N_12898,N_12781,N_12799);
xnor U12899 (N_12899,N_12251,N_12108);
or U12900 (N_12900,N_12642,N_12093);
and U12901 (N_12901,N_12541,N_12255);
xor U12902 (N_12902,N_12487,N_12333);
or U12903 (N_12903,N_12148,N_12538);
nor U12904 (N_12904,N_12661,N_12431);
nand U12905 (N_12905,N_12010,N_12131);
and U12906 (N_12906,N_12312,N_12741);
nor U12907 (N_12907,N_12271,N_12384);
nor U12908 (N_12908,N_12476,N_12774);
and U12909 (N_12909,N_12771,N_12611);
nand U12910 (N_12910,N_12034,N_12780);
xnor U12911 (N_12911,N_12260,N_12104);
nor U12912 (N_12912,N_12099,N_12391);
nor U12913 (N_12913,N_12640,N_12044);
xor U12914 (N_12914,N_12051,N_12158);
and U12915 (N_12915,N_12566,N_12296);
or U12916 (N_12916,N_12266,N_12516);
nor U12917 (N_12917,N_12113,N_12732);
and U12918 (N_12918,N_12797,N_12211);
nor U12919 (N_12919,N_12450,N_12241);
xnor U12920 (N_12920,N_12658,N_12483);
nor U12921 (N_12921,N_12197,N_12467);
xor U12922 (N_12922,N_12056,N_12017);
xor U12923 (N_12923,N_12216,N_12084);
nand U12924 (N_12924,N_12621,N_12256);
nand U12925 (N_12925,N_12416,N_12054);
nand U12926 (N_12926,N_12677,N_12309);
nand U12927 (N_12927,N_12349,N_12032);
or U12928 (N_12928,N_12358,N_12062);
nand U12929 (N_12929,N_12437,N_12417);
nand U12930 (N_12930,N_12169,N_12191);
or U12931 (N_12931,N_12360,N_12482);
and U12932 (N_12932,N_12509,N_12347);
nand U12933 (N_12933,N_12081,N_12232);
xnor U12934 (N_12934,N_12174,N_12351);
or U12935 (N_12935,N_12114,N_12745);
and U12936 (N_12936,N_12546,N_12204);
xor U12937 (N_12937,N_12674,N_12635);
or U12938 (N_12938,N_12743,N_12175);
nand U12939 (N_12939,N_12652,N_12036);
and U12940 (N_12940,N_12006,N_12409);
nor U12941 (N_12941,N_12406,N_12660);
nand U12942 (N_12942,N_12199,N_12414);
nor U12943 (N_12943,N_12355,N_12634);
xor U12944 (N_12944,N_12507,N_12762);
xor U12945 (N_12945,N_12285,N_12528);
xnor U12946 (N_12946,N_12529,N_12340);
and U12947 (N_12947,N_12469,N_12770);
xor U12948 (N_12948,N_12101,N_12059);
nor U12949 (N_12949,N_12419,N_12764);
nand U12950 (N_12950,N_12449,N_12557);
and U12951 (N_12951,N_12793,N_12702);
or U12952 (N_12952,N_12435,N_12618);
nor U12953 (N_12953,N_12284,N_12208);
xnor U12954 (N_12954,N_12345,N_12224);
xnor U12955 (N_12955,N_12646,N_12593);
xor U12956 (N_12956,N_12549,N_12517);
xnor U12957 (N_12957,N_12286,N_12547);
nand U12958 (N_12958,N_12069,N_12365);
and U12959 (N_12959,N_12491,N_12377);
xnor U12960 (N_12960,N_12303,N_12544);
nor U12961 (N_12961,N_12306,N_12494);
and U12962 (N_12962,N_12462,N_12694);
or U12963 (N_12963,N_12510,N_12295);
or U12964 (N_12964,N_12124,N_12025);
xor U12965 (N_12965,N_12438,N_12133);
and U12966 (N_12966,N_12274,N_12396);
nor U12967 (N_12967,N_12472,N_12075);
nand U12968 (N_12968,N_12443,N_12234);
nor U12969 (N_12969,N_12657,N_12697);
or U12970 (N_12970,N_12300,N_12177);
and U12971 (N_12971,N_12373,N_12332);
nand U12972 (N_12972,N_12000,N_12446);
or U12973 (N_12973,N_12654,N_12165);
xnor U12974 (N_12974,N_12787,N_12639);
nand U12975 (N_12975,N_12123,N_12090);
or U12976 (N_12976,N_12226,N_12591);
nand U12977 (N_12977,N_12606,N_12713);
nor U12978 (N_12978,N_12112,N_12638);
nand U12979 (N_12979,N_12647,N_12040);
xnor U12980 (N_12980,N_12014,N_12563);
nor U12981 (N_12981,N_12457,N_12521);
and U12982 (N_12982,N_12063,N_12368);
and U12983 (N_12983,N_12096,N_12405);
and U12984 (N_12984,N_12083,N_12533);
or U12985 (N_12985,N_12137,N_12076);
and U12986 (N_12986,N_12029,N_12712);
nand U12987 (N_12987,N_12129,N_12455);
nor U12988 (N_12988,N_12213,N_12217);
and U12989 (N_12989,N_12343,N_12092);
nand U12990 (N_12990,N_12142,N_12788);
or U12991 (N_12991,N_12682,N_12777);
and U12992 (N_12992,N_12294,N_12474);
and U12993 (N_12993,N_12445,N_12570);
xor U12994 (N_12994,N_12536,N_12626);
xor U12995 (N_12995,N_12227,N_12086);
xnor U12996 (N_12996,N_12519,N_12508);
or U12997 (N_12997,N_12183,N_12170);
nor U12998 (N_12998,N_12046,N_12095);
xnor U12999 (N_12999,N_12691,N_12601);
and U13000 (N_13000,N_12105,N_12730);
nor U13001 (N_13001,N_12719,N_12376);
nor U13002 (N_13002,N_12558,N_12161);
or U13003 (N_13003,N_12530,N_12206);
nor U13004 (N_13004,N_12598,N_12272);
nand U13005 (N_13005,N_12512,N_12315);
or U13006 (N_13006,N_12219,N_12223);
xnor U13007 (N_13007,N_12280,N_12543);
and U13008 (N_13008,N_12643,N_12757);
or U13009 (N_13009,N_12722,N_12442);
xnor U13010 (N_13010,N_12033,N_12395);
or U13011 (N_13011,N_12631,N_12342);
and U13012 (N_13012,N_12242,N_12230);
nor U13013 (N_13013,N_12008,N_12111);
nand U13014 (N_13014,N_12523,N_12415);
or U13015 (N_13015,N_12192,N_12426);
xnor U13016 (N_13016,N_12314,N_12559);
nor U13017 (N_13017,N_12531,N_12581);
or U13018 (N_13018,N_12352,N_12744);
nor U13019 (N_13019,N_12004,N_12307);
and U13020 (N_13020,N_12542,N_12608);
and U13021 (N_13021,N_12599,N_12261);
nor U13022 (N_13022,N_12663,N_12703);
and U13023 (N_13023,N_12135,N_12057);
or U13024 (N_13024,N_12766,N_12012);
or U13025 (N_13025,N_12042,N_12369);
xnor U13026 (N_13026,N_12695,N_12100);
and U13027 (N_13027,N_12689,N_12385);
and U13028 (N_13028,N_12458,N_12106);
or U13029 (N_13029,N_12447,N_12676);
and U13030 (N_13030,N_12616,N_12548);
and U13031 (N_13031,N_12779,N_12413);
or U13032 (N_13032,N_12715,N_12188);
or U13033 (N_13033,N_12061,N_12334);
xor U13034 (N_13034,N_12279,N_12716);
xnor U13035 (N_13035,N_12586,N_12432);
or U13036 (N_13036,N_12700,N_12668);
or U13037 (N_13037,N_12710,N_12410);
xor U13038 (N_13038,N_12681,N_12239);
nor U13039 (N_13039,N_12143,N_12773);
nor U13040 (N_13040,N_12246,N_12551);
nand U13041 (N_13041,N_12669,N_12212);
nor U13042 (N_13042,N_12448,N_12055);
and U13043 (N_13043,N_12791,N_12180);
nor U13044 (N_13044,N_12539,N_12386);
nor U13045 (N_13045,N_12434,N_12035);
xor U13046 (N_13046,N_12670,N_12477);
nand U13047 (N_13047,N_12027,N_12389);
and U13048 (N_13048,N_12708,N_12074);
and U13049 (N_13049,N_12580,N_12602);
nor U13050 (N_13050,N_12783,N_12024);
nor U13051 (N_13051,N_12707,N_12293);
or U13052 (N_13052,N_12784,N_12534);
xnor U13053 (N_13053,N_12614,N_12605);
xor U13054 (N_13054,N_12078,N_12613);
xor U13055 (N_13055,N_12751,N_12451);
or U13056 (N_13056,N_12354,N_12379);
and U13057 (N_13057,N_12604,N_12128);
or U13058 (N_13058,N_12709,N_12392);
or U13059 (N_13059,N_12321,N_12739);
nand U13060 (N_13060,N_12425,N_12007);
nand U13061 (N_13061,N_12490,N_12701);
nand U13062 (N_13062,N_12073,N_12488);
and U13063 (N_13063,N_12734,N_12350);
nor U13064 (N_13064,N_12013,N_12790);
xnor U13065 (N_13065,N_12632,N_12504);
nor U13066 (N_13066,N_12685,N_12336);
xor U13067 (N_13067,N_12500,N_12233);
xnor U13068 (N_13068,N_12515,N_12575);
nand U13069 (N_13069,N_12444,N_12149);
nand U13070 (N_13070,N_12194,N_12620);
or U13071 (N_13071,N_12583,N_12696);
and U13072 (N_13072,N_12585,N_12005);
xnor U13073 (N_13073,N_12154,N_12486);
nand U13074 (N_13074,N_12574,N_12281);
nor U13075 (N_13075,N_12750,N_12187);
or U13076 (N_13076,N_12624,N_12456);
xnor U13077 (N_13077,N_12254,N_12738);
xor U13078 (N_13078,N_12520,N_12152);
and U13079 (N_13079,N_12423,N_12023);
nand U13080 (N_13080,N_12060,N_12495);
xnor U13081 (N_13081,N_12209,N_12037);
and U13082 (N_13082,N_12466,N_12337);
and U13083 (N_13083,N_12727,N_12594);
nor U13084 (N_13084,N_12537,N_12176);
xnor U13085 (N_13085,N_12258,N_12238);
nand U13086 (N_13086,N_12378,N_12330);
nor U13087 (N_13087,N_12513,N_12120);
or U13088 (N_13088,N_12755,N_12068);
and U13089 (N_13089,N_12147,N_12275);
and U13090 (N_13090,N_12262,N_12526);
nand U13091 (N_13091,N_12018,N_12196);
and U13092 (N_13092,N_12228,N_12387);
xnor U13093 (N_13093,N_12072,N_12353);
and U13094 (N_13094,N_12325,N_12424);
xor U13095 (N_13095,N_12162,N_12136);
nand U13096 (N_13096,N_12473,N_12375);
xor U13097 (N_13097,N_12441,N_12021);
and U13098 (N_13098,N_12102,N_12058);
nor U13099 (N_13099,N_12374,N_12015);
nand U13100 (N_13100,N_12214,N_12249);
xor U13101 (N_13101,N_12270,N_12502);
xnor U13102 (N_13102,N_12720,N_12248);
nor U13103 (N_13103,N_12001,N_12045);
nor U13104 (N_13104,N_12429,N_12164);
nand U13105 (N_13105,N_12475,N_12690);
and U13106 (N_13106,N_12341,N_12603);
xnor U13107 (N_13107,N_12420,N_12202);
and U13108 (N_13108,N_12383,N_12662);
and U13109 (N_13109,N_12166,N_12116);
nor U13110 (N_13110,N_12065,N_12372);
xor U13111 (N_13111,N_12679,N_12552);
or U13112 (N_13112,N_12648,N_12461);
xnor U13113 (N_13113,N_12382,N_12171);
nor U13114 (N_13114,N_12319,N_12329);
nand U13115 (N_13115,N_12370,N_12485);
and U13116 (N_13116,N_12776,N_12130);
or U13117 (N_13117,N_12290,N_12399);
nand U13118 (N_13118,N_12740,N_12711);
and U13119 (N_13119,N_12556,N_12698);
xor U13120 (N_13120,N_12464,N_12430);
nand U13121 (N_13121,N_12366,N_12091);
nor U13122 (N_13122,N_12422,N_12752);
or U13123 (N_13123,N_12489,N_12119);
or U13124 (N_13124,N_12134,N_12579);
or U13125 (N_13125,N_12153,N_12573);
or U13126 (N_13126,N_12322,N_12323);
nor U13127 (N_13127,N_12767,N_12637);
nor U13128 (N_13128,N_12470,N_12198);
nand U13129 (N_13129,N_12688,N_12229);
or U13130 (N_13130,N_12338,N_12247);
and U13131 (N_13131,N_12089,N_12404);
xor U13132 (N_13132,N_12344,N_12094);
and U13133 (N_13133,N_12737,N_12144);
and U13134 (N_13134,N_12041,N_12016);
and U13135 (N_13135,N_12066,N_12629);
xor U13136 (N_13136,N_12747,N_12028);
xor U13137 (N_13137,N_12560,N_12651);
nand U13138 (N_13138,N_12650,N_12571);
or U13139 (N_13139,N_12257,N_12421);
or U13140 (N_13140,N_12328,N_12723);
xnor U13141 (N_13141,N_12452,N_12692);
or U13142 (N_13142,N_12259,N_12145);
nand U13143 (N_13143,N_12356,N_12245);
and U13144 (N_13144,N_12714,N_12794);
and U13145 (N_13145,N_12772,N_12117);
nand U13146 (N_13146,N_12769,N_12471);
nand U13147 (N_13147,N_12235,N_12705);
or U13148 (N_13148,N_12291,N_12525);
nor U13149 (N_13149,N_12132,N_12582);
xnor U13150 (N_13150,N_12717,N_12704);
xnor U13151 (N_13151,N_12087,N_12636);
xnor U13152 (N_13152,N_12496,N_12098);
nor U13153 (N_13153,N_12393,N_12052);
nand U13154 (N_13154,N_12022,N_12173);
nand U13155 (N_13155,N_12020,N_12796);
nand U13156 (N_13156,N_12287,N_12765);
nor U13157 (N_13157,N_12622,N_12103);
xnor U13158 (N_13158,N_12768,N_12746);
nand U13159 (N_13159,N_12305,N_12565);
nor U13160 (N_13160,N_12572,N_12522);
xnor U13161 (N_13161,N_12735,N_12561);
or U13162 (N_13162,N_12361,N_12205);
xnor U13163 (N_13163,N_12675,N_12273);
xor U13164 (N_13164,N_12097,N_12693);
xnor U13165 (N_13165,N_12665,N_12731);
or U13166 (N_13166,N_12172,N_12215);
xnor U13167 (N_13167,N_12110,N_12218);
or U13168 (N_13168,N_12480,N_12659);
nand U13169 (N_13169,N_12250,N_12079);
xor U13170 (N_13170,N_12607,N_12645);
nor U13171 (N_13171,N_12497,N_12388);
nand U13172 (N_13172,N_12390,N_12118);
and U13173 (N_13173,N_12699,N_12569);
nor U13174 (N_13174,N_12019,N_12184);
nand U13175 (N_13175,N_12302,N_12479);
nor U13176 (N_13176,N_12459,N_12225);
or U13177 (N_13177,N_12554,N_12394);
nand U13178 (N_13178,N_12115,N_12492);
and U13179 (N_13179,N_12753,N_12729);
nand U13180 (N_13180,N_12179,N_12759);
xnor U13181 (N_13181,N_12237,N_12278);
and U13182 (N_13182,N_12085,N_12038);
xor U13183 (N_13183,N_12222,N_12550);
nand U13184 (N_13184,N_12749,N_12633);
nor U13185 (N_13185,N_12454,N_12397);
and U13186 (N_13186,N_12026,N_12348);
nand U13187 (N_13187,N_12297,N_12742);
xnor U13188 (N_13188,N_12798,N_12758);
and U13189 (N_13189,N_12680,N_12463);
nand U13190 (N_13190,N_12577,N_12359);
and U13191 (N_13191,N_12181,N_12763);
xnor U13192 (N_13192,N_12761,N_12686);
nand U13193 (N_13193,N_12031,N_12326);
or U13194 (N_13194,N_12203,N_12786);
and U13195 (N_13195,N_12527,N_12331);
nand U13196 (N_13196,N_12138,N_12009);
and U13197 (N_13197,N_12733,N_12460);
nand U13198 (N_13198,N_12641,N_12588);
xor U13199 (N_13199,N_12304,N_12664);
nand U13200 (N_13200,N_12687,N_12570);
and U13201 (N_13201,N_12487,N_12211);
xnor U13202 (N_13202,N_12161,N_12212);
nor U13203 (N_13203,N_12571,N_12451);
xnor U13204 (N_13204,N_12679,N_12030);
nand U13205 (N_13205,N_12277,N_12301);
and U13206 (N_13206,N_12798,N_12755);
or U13207 (N_13207,N_12645,N_12419);
xor U13208 (N_13208,N_12542,N_12681);
or U13209 (N_13209,N_12536,N_12347);
nand U13210 (N_13210,N_12027,N_12780);
or U13211 (N_13211,N_12783,N_12404);
nand U13212 (N_13212,N_12093,N_12189);
and U13213 (N_13213,N_12793,N_12531);
or U13214 (N_13214,N_12340,N_12297);
nor U13215 (N_13215,N_12542,N_12554);
xnor U13216 (N_13216,N_12165,N_12411);
xor U13217 (N_13217,N_12778,N_12026);
xor U13218 (N_13218,N_12661,N_12458);
and U13219 (N_13219,N_12739,N_12201);
and U13220 (N_13220,N_12694,N_12220);
nand U13221 (N_13221,N_12494,N_12244);
nor U13222 (N_13222,N_12556,N_12043);
xnor U13223 (N_13223,N_12339,N_12159);
nand U13224 (N_13224,N_12189,N_12459);
xor U13225 (N_13225,N_12493,N_12565);
and U13226 (N_13226,N_12527,N_12435);
or U13227 (N_13227,N_12223,N_12754);
xor U13228 (N_13228,N_12754,N_12731);
nand U13229 (N_13229,N_12297,N_12088);
xnor U13230 (N_13230,N_12435,N_12692);
and U13231 (N_13231,N_12373,N_12641);
and U13232 (N_13232,N_12552,N_12687);
and U13233 (N_13233,N_12533,N_12435);
nor U13234 (N_13234,N_12281,N_12066);
nor U13235 (N_13235,N_12790,N_12795);
and U13236 (N_13236,N_12029,N_12345);
nand U13237 (N_13237,N_12587,N_12002);
and U13238 (N_13238,N_12179,N_12141);
and U13239 (N_13239,N_12492,N_12131);
nor U13240 (N_13240,N_12166,N_12448);
or U13241 (N_13241,N_12313,N_12733);
xor U13242 (N_13242,N_12716,N_12740);
and U13243 (N_13243,N_12214,N_12402);
and U13244 (N_13244,N_12051,N_12652);
nor U13245 (N_13245,N_12002,N_12442);
xnor U13246 (N_13246,N_12038,N_12587);
and U13247 (N_13247,N_12142,N_12798);
xor U13248 (N_13248,N_12047,N_12117);
xor U13249 (N_13249,N_12636,N_12633);
nor U13250 (N_13250,N_12009,N_12714);
and U13251 (N_13251,N_12788,N_12198);
xor U13252 (N_13252,N_12744,N_12661);
or U13253 (N_13253,N_12131,N_12397);
xnor U13254 (N_13254,N_12379,N_12706);
or U13255 (N_13255,N_12579,N_12405);
nand U13256 (N_13256,N_12399,N_12105);
xor U13257 (N_13257,N_12760,N_12157);
nand U13258 (N_13258,N_12166,N_12131);
and U13259 (N_13259,N_12511,N_12291);
or U13260 (N_13260,N_12795,N_12076);
nand U13261 (N_13261,N_12567,N_12442);
nor U13262 (N_13262,N_12633,N_12245);
xor U13263 (N_13263,N_12502,N_12166);
or U13264 (N_13264,N_12556,N_12217);
nor U13265 (N_13265,N_12148,N_12689);
nor U13266 (N_13266,N_12242,N_12768);
nor U13267 (N_13267,N_12603,N_12465);
and U13268 (N_13268,N_12289,N_12281);
and U13269 (N_13269,N_12114,N_12390);
or U13270 (N_13270,N_12047,N_12365);
nor U13271 (N_13271,N_12198,N_12150);
or U13272 (N_13272,N_12783,N_12507);
xnor U13273 (N_13273,N_12305,N_12774);
nor U13274 (N_13274,N_12189,N_12343);
or U13275 (N_13275,N_12132,N_12534);
or U13276 (N_13276,N_12314,N_12639);
nand U13277 (N_13277,N_12734,N_12348);
nand U13278 (N_13278,N_12465,N_12195);
xor U13279 (N_13279,N_12162,N_12583);
nor U13280 (N_13280,N_12099,N_12445);
nor U13281 (N_13281,N_12525,N_12165);
or U13282 (N_13282,N_12322,N_12633);
xor U13283 (N_13283,N_12526,N_12701);
nand U13284 (N_13284,N_12352,N_12069);
and U13285 (N_13285,N_12073,N_12046);
xor U13286 (N_13286,N_12113,N_12250);
nor U13287 (N_13287,N_12098,N_12726);
and U13288 (N_13288,N_12608,N_12655);
and U13289 (N_13289,N_12286,N_12296);
nand U13290 (N_13290,N_12556,N_12595);
xor U13291 (N_13291,N_12124,N_12556);
and U13292 (N_13292,N_12536,N_12755);
and U13293 (N_13293,N_12483,N_12637);
or U13294 (N_13294,N_12164,N_12143);
or U13295 (N_13295,N_12102,N_12228);
xor U13296 (N_13296,N_12406,N_12105);
nand U13297 (N_13297,N_12497,N_12792);
and U13298 (N_13298,N_12498,N_12560);
and U13299 (N_13299,N_12269,N_12732);
or U13300 (N_13300,N_12392,N_12386);
nand U13301 (N_13301,N_12346,N_12394);
nor U13302 (N_13302,N_12757,N_12163);
xor U13303 (N_13303,N_12359,N_12719);
or U13304 (N_13304,N_12107,N_12412);
or U13305 (N_13305,N_12229,N_12334);
or U13306 (N_13306,N_12252,N_12451);
nor U13307 (N_13307,N_12611,N_12703);
nand U13308 (N_13308,N_12134,N_12262);
xor U13309 (N_13309,N_12367,N_12693);
nand U13310 (N_13310,N_12358,N_12627);
xnor U13311 (N_13311,N_12147,N_12652);
or U13312 (N_13312,N_12077,N_12452);
nor U13313 (N_13313,N_12689,N_12003);
or U13314 (N_13314,N_12204,N_12015);
nand U13315 (N_13315,N_12477,N_12734);
xnor U13316 (N_13316,N_12736,N_12582);
and U13317 (N_13317,N_12207,N_12025);
or U13318 (N_13318,N_12725,N_12559);
and U13319 (N_13319,N_12548,N_12623);
or U13320 (N_13320,N_12372,N_12028);
and U13321 (N_13321,N_12615,N_12408);
or U13322 (N_13322,N_12062,N_12539);
nor U13323 (N_13323,N_12181,N_12429);
and U13324 (N_13324,N_12681,N_12538);
xnor U13325 (N_13325,N_12537,N_12618);
or U13326 (N_13326,N_12101,N_12157);
nor U13327 (N_13327,N_12285,N_12741);
nor U13328 (N_13328,N_12655,N_12047);
nor U13329 (N_13329,N_12252,N_12542);
and U13330 (N_13330,N_12615,N_12222);
xor U13331 (N_13331,N_12418,N_12172);
or U13332 (N_13332,N_12185,N_12439);
or U13333 (N_13333,N_12675,N_12161);
nand U13334 (N_13334,N_12582,N_12622);
nand U13335 (N_13335,N_12781,N_12641);
nand U13336 (N_13336,N_12228,N_12321);
nor U13337 (N_13337,N_12172,N_12246);
nand U13338 (N_13338,N_12536,N_12588);
nor U13339 (N_13339,N_12623,N_12372);
nand U13340 (N_13340,N_12552,N_12691);
xor U13341 (N_13341,N_12698,N_12765);
nand U13342 (N_13342,N_12563,N_12562);
nand U13343 (N_13343,N_12055,N_12633);
nand U13344 (N_13344,N_12616,N_12112);
or U13345 (N_13345,N_12668,N_12509);
nor U13346 (N_13346,N_12013,N_12682);
nor U13347 (N_13347,N_12428,N_12000);
or U13348 (N_13348,N_12079,N_12105);
xnor U13349 (N_13349,N_12600,N_12377);
nand U13350 (N_13350,N_12079,N_12455);
xor U13351 (N_13351,N_12546,N_12713);
xor U13352 (N_13352,N_12377,N_12233);
nor U13353 (N_13353,N_12407,N_12754);
xor U13354 (N_13354,N_12215,N_12288);
or U13355 (N_13355,N_12443,N_12767);
and U13356 (N_13356,N_12443,N_12673);
and U13357 (N_13357,N_12336,N_12398);
or U13358 (N_13358,N_12460,N_12506);
and U13359 (N_13359,N_12623,N_12143);
or U13360 (N_13360,N_12693,N_12719);
and U13361 (N_13361,N_12490,N_12413);
or U13362 (N_13362,N_12247,N_12501);
and U13363 (N_13363,N_12425,N_12096);
or U13364 (N_13364,N_12338,N_12399);
and U13365 (N_13365,N_12376,N_12098);
nand U13366 (N_13366,N_12441,N_12523);
nor U13367 (N_13367,N_12195,N_12586);
nor U13368 (N_13368,N_12125,N_12385);
or U13369 (N_13369,N_12358,N_12530);
or U13370 (N_13370,N_12565,N_12710);
and U13371 (N_13371,N_12531,N_12248);
nor U13372 (N_13372,N_12449,N_12118);
and U13373 (N_13373,N_12044,N_12549);
nor U13374 (N_13374,N_12605,N_12241);
nand U13375 (N_13375,N_12423,N_12347);
nor U13376 (N_13376,N_12502,N_12747);
nor U13377 (N_13377,N_12428,N_12306);
and U13378 (N_13378,N_12593,N_12110);
nand U13379 (N_13379,N_12497,N_12785);
nor U13380 (N_13380,N_12604,N_12276);
nor U13381 (N_13381,N_12339,N_12025);
and U13382 (N_13382,N_12426,N_12531);
nand U13383 (N_13383,N_12168,N_12631);
or U13384 (N_13384,N_12518,N_12166);
xnor U13385 (N_13385,N_12702,N_12511);
or U13386 (N_13386,N_12318,N_12079);
nand U13387 (N_13387,N_12110,N_12323);
or U13388 (N_13388,N_12574,N_12136);
and U13389 (N_13389,N_12039,N_12134);
and U13390 (N_13390,N_12601,N_12774);
and U13391 (N_13391,N_12647,N_12177);
or U13392 (N_13392,N_12605,N_12011);
or U13393 (N_13393,N_12799,N_12342);
and U13394 (N_13394,N_12487,N_12370);
nor U13395 (N_13395,N_12029,N_12048);
and U13396 (N_13396,N_12618,N_12641);
or U13397 (N_13397,N_12794,N_12080);
xnor U13398 (N_13398,N_12673,N_12758);
xnor U13399 (N_13399,N_12063,N_12524);
or U13400 (N_13400,N_12110,N_12071);
nand U13401 (N_13401,N_12111,N_12169);
nor U13402 (N_13402,N_12637,N_12080);
xor U13403 (N_13403,N_12240,N_12317);
nor U13404 (N_13404,N_12314,N_12650);
and U13405 (N_13405,N_12791,N_12576);
xnor U13406 (N_13406,N_12036,N_12633);
nand U13407 (N_13407,N_12100,N_12195);
xnor U13408 (N_13408,N_12538,N_12074);
nor U13409 (N_13409,N_12030,N_12770);
nor U13410 (N_13410,N_12038,N_12115);
xnor U13411 (N_13411,N_12156,N_12023);
nor U13412 (N_13412,N_12142,N_12315);
xor U13413 (N_13413,N_12362,N_12201);
or U13414 (N_13414,N_12470,N_12412);
nand U13415 (N_13415,N_12079,N_12720);
xnor U13416 (N_13416,N_12610,N_12697);
nand U13417 (N_13417,N_12485,N_12274);
and U13418 (N_13418,N_12562,N_12325);
or U13419 (N_13419,N_12212,N_12035);
and U13420 (N_13420,N_12519,N_12487);
and U13421 (N_13421,N_12383,N_12477);
and U13422 (N_13422,N_12744,N_12055);
xnor U13423 (N_13423,N_12032,N_12224);
nor U13424 (N_13424,N_12604,N_12719);
nand U13425 (N_13425,N_12764,N_12533);
nor U13426 (N_13426,N_12736,N_12131);
and U13427 (N_13427,N_12512,N_12337);
and U13428 (N_13428,N_12614,N_12460);
xor U13429 (N_13429,N_12096,N_12698);
nand U13430 (N_13430,N_12753,N_12705);
xnor U13431 (N_13431,N_12317,N_12000);
and U13432 (N_13432,N_12190,N_12177);
xor U13433 (N_13433,N_12733,N_12084);
nand U13434 (N_13434,N_12775,N_12511);
nand U13435 (N_13435,N_12006,N_12310);
nor U13436 (N_13436,N_12468,N_12739);
nor U13437 (N_13437,N_12401,N_12195);
and U13438 (N_13438,N_12594,N_12067);
nand U13439 (N_13439,N_12319,N_12743);
or U13440 (N_13440,N_12315,N_12542);
nand U13441 (N_13441,N_12198,N_12458);
xor U13442 (N_13442,N_12183,N_12262);
nand U13443 (N_13443,N_12482,N_12121);
xnor U13444 (N_13444,N_12664,N_12198);
nand U13445 (N_13445,N_12786,N_12529);
xor U13446 (N_13446,N_12129,N_12689);
or U13447 (N_13447,N_12591,N_12057);
and U13448 (N_13448,N_12126,N_12705);
or U13449 (N_13449,N_12410,N_12226);
xnor U13450 (N_13450,N_12538,N_12697);
nand U13451 (N_13451,N_12015,N_12055);
xnor U13452 (N_13452,N_12569,N_12762);
and U13453 (N_13453,N_12764,N_12186);
xor U13454 (N_13454,N_12066,N_12587);
nor U13455 (N_13455,N_12662,N_12311);
xor U13456 (N_13456,N_12733,N_12335);
and U13457 (N_13457,N_12243,N_12240);
nor U13458 (N_13458,N_12121,N_12467);
and U13459 (N_13459,N_12139,N_12795);
nor U13460 (N_13460,N_12646,N_12724);
xor U13461 (N_13461,N_12182,N_12032);
and U13462 (N_13462,N_12181,N_12046);
and U13463 (N_13463,N_12753,N_12101);
and U13464 (N_13464,N_12150,N_12335);
or U13465 (N_13465,N_12257,N_12573);
or U13466 (N_13466,N_12521,N_12309);
nor U13467 (N_13467,N_12580,N_12623);
or U13468 (N_13468,N_12633,N_12671);
nor U13469 (N_13469,N_12390,N_12217);
xnor U13470 (N_13470,N_12259,N_12657);
nor U13471 (N_13471,N_12398,N_12270);
or U13472 (N_13472,N_12726,N_12238);
nand U13473 (N_13473,N_12287,N_12715);
nor U13474 (N_13474,N_12479,N_12234);
or U13475 (N_13475,N_12641,N_12210);
xor U13476 (N_13476,N_12424,N_12792);
xnor U13477 (N_13477,N_12387,N_12421);
xnor U13478 (N_13478,N_12737,N_12478);
and U13479 (N_13479,N_12436,N_12302);
xor U13480 (N_13480,N_12355,N_12167);
and U13481 (N_13481,N_12293,N_12711);
nor U13482 (N_13482,N_12104,N_12784);
or U13483 (N_13483,N_12145,N_12023);
and U13484 (N_13484,N_12216,N_12700);
nand U13485 (N_13485,N_12187,N_12071);
xor U13486 (N_13486,N_12053,N_12051);
nor U13487 (N_13487,N_12345,N_12281);
nand U13488 (N_13488,N_12560,N_12728);
and U13489 (N_13489,N_12023,N_12393);
and U13490 (N_13490,N_12439,N_12550);
nand U13491 (N_13491,N_12754,N_12208);
or U13492 (N_13492,N_12220,N_12341);
or U13493 (N_13493,N_12081,N_12086);
nor U13494 (N_13494,N_12196,N_12636);
and U13495 (N_13495,N_12614,N_12037);
and U13496 (N_13496,N_12480,N_12595);
xnor U13497 (N_13497,N_12304,N_12183);
or U13498 (N_13498,N_12760,N_12326);
nor U13499 (N_13499,N_12517,N_12065);
nand U13500 (N_13500,N_12431,N_12534);
nand U13501 (N_13501,N_12440,N_12451);
nand U13502 (N_13502,N_12604,N_12205);
nand U13503 (N_13503,N_12508,N_12045);
nand U13504 (N_13504,N_12784,N_12216);
and U13505 (N_13505,N_12161,N_12546);
nand U13506 (N_13506,N_12714,N_12617);
and U13507 (N_13507,N_12058,N_12602);
xnor U13508 (N_13508,N_12656,N_12117);
nor U13509 (N_13509,N_12466,N_12743);
or U13510 (N_13510,N_12164,N_12564);
nand U13511 (N_13511,N_12184,N_12286);
xor U13512 (N_13512,N_12642,N_12239);
nor U13513 (N_13513,N_12575,N_12435);
nand U13514 (N_13514,N_12427,N_12017);
or U13515 (N_13515,N_12212,N_12738);
xnor U13516 (N_13516,N_12178,N_12370);
nor U13517 (N_13517,N_12291,N_12146);
xnor U13518 (N_13518,N_12255,N_12199);
and U13519 (N_13519,N_12303,N_12325);
and U13520 (N_13520,N_12129,N_12739);
or U13521 (N_13521,N_12716,N_12013);
nor U13522 (N_13522,N_12598,N_12573);
and U13523 (N_13523,N_12539,N_12712);
xnor U13524 (N_13524,N_12047,N_12519);
or U13525 (N_13525,N_12440,N_12052);
nor U13526 (N_13526,N_12609,N_12721);
and U13527 (N_13527,N_12743,N_12279);
or U13528 (N_13528,N_12089,N_12518);
nand U13529 (N_13529,N_12428,N_12046);
nor U13530 (N_13530,N_12034,N_12006);
and U13531 (N_13531,N_12073,N_12479);
or U13532 (N_13532,N_12142,N_12519);
nor U13533 (N_13533,N_12030,N_12085);
and U13534 (N_13534,N_12421,N_12608);
nand U13535 (N_13535,N_12060,N_12432);
xor U13536 (N_13536,N_12622,N_12369);
and U13537 (N_13537,N_12038,N_12634);
nor U13538 (N_13538,N_12260,N_12013);
and U13539 (N_13539,N_12678,N_12416);
nor U13540 (N_13540,N_12173,N_12447);
or U13541 (N_13541,N_12615,N_12253);
and U13542 (N_13542,N_12249,N_12552);
or U13543 (N_13543,N_12270,N_12763);
xor U13544 (N_13544,N_12173,N_12654);
nand U13545 (N_13545,N_12553,N_12204);
or U13546 (N_13546,N_12255,N_12275);
and U13547 (N_13547,N_12650,N_12543);
xor U13548 (N_13548,N_12276,N_12372);
and U13549 (N_13549,N_12212,N_12469);
and U13550 (N_13550,N_12453,N_12372);
nor U13551 (N_13551,N_12604,N_12654);
nand U13552 (N_13552,N_12430,N_12199);
nor U13553 (N_13553,N_12161,N_12330);
nor U13554 (N_13554,N_12340,N_12463);
nand U13555 (N_13555,N_12451,N_12342);
xnor U13556 (N_13556,N_12661,N_12552);
xor U13557 (N_13557,N_12131,N_12657);
and U13558 (N_13558,N_12516,N_12414);
nand U13559 (N_13559,N_12457,N_12023);
and U13560 (N_13560,N_12200,N_12757);
nor U13561 (N_13561,N_12689,N_12600);
nor U13562 (N_13562,N_12050,N_12354);
and U13563 (N_13563,N_12397,N_12425);
nand U13564 (N_13564,N_12163,N_12313);
and U13565 (N_13565,N_12026,N_12090);
and U13566 (N_13566,N_12449,N_12101);
or U13567 (N_13567,N_12443,N_12536);
nor U13568 (N_13568,N_12279,N_12780);
xor U13569 (N_13569,N_12733,N_12128);
xor U13570 (N_13570,N_12572,N_12523);
and U13571 (N_13571,N_12045,N_12561);
nor U13572 (N_13572,N_12795,N_12056);
nor U13573 (N_13573,N_12786,N_12425);
or U13574 (N_13574,N_12245,N_12514);
or U13575 (N_13575,N_12454,N_12477);
xnor U13576 (N_13576,N_12224,N_12203);
nand U13577 (N_13577,N_12086,N_12063);
or U13578 (N_13578,N_12174,N_12138);
or U13579 (N_13579,N_12341,N_12090);
nand U13580 (N_13580,N_12124,N_12334);
or U13581 (N_13581,N_12529,N_12427);
and U13582 (N_13582,N_12775,N_12460);
or U13583 (N_13583,N_12551,N_12169);
nand U13584 (N_13584,N_12639,N_12245);
or U13585 (N_13585,N_12601,N_12103);
nand U13586 (N_13586,N_12563,N_12055);
nor U13587 (N_13587,N_12017,N_12333);
or U13588 (N_13588,N_12394,N_12757);
or U13589 (N_13589,N_12163,N_12784);
and U13590 (N_13590,N_12218,N_12564);
nor U13591 (N_13591,N_12451,N_12220);
or U13592 (N_13592,N_12309,N_12028);
nor U13593 (N_13593,N_12137,N_12345);
and U13594 (N_13594,N_12393,N_12725);
xnor U13595 (N_13595,N_12490,N_12690);
nand U13596 (N_13596,N_12579,N_12397);
or U13597 (N_13597,N_12423,N_12727);
nand U13598 (N_13598,N_12688,N_12064);
xor U13599 (N_13599,N_12685,N_12507);
nor U13600 (N_13600,N_13041,N_13340);
nor U13601 (N_13601,N_12877,N_13237);
and U13602 (N_13602,N_13234,N_12925);
nor U13603 (N_13603,N_12890,N_12905);
nor U13604 (N_13604,N_13258,N_13277);
xnor U13605 (N_13605,N_13485,N_12979);
nand U13606 (N_13606,N_13246,N_12878);
nand U13607 (N_13607,N_12961,N_13230);
or U13608 (N_13608,N_13442,N_13212);
nand U13609 (N_13609,N_13429,N_13040);
xnor U13610 (N_13610,N_12833,N_13425);
nor U13611 (N_13611,N_13427,N_12930);
or U13612 (N_13612,N_13083,N_13367);
nor U13613 (N_13613,N_13168,N_13399);
nand U13614 (N_13614,N_13387,N_13287);
nand U13615 (N_13615,N_13324,N_13097);
nor U13616 (N_13616,N_12949,N_13346);
nor U13617 (N_13617,N_12875,N_13444);
or U13618 (N_13618,N_13109,N_13231);
and U13619 (N_13619,N_13142,N_13268);
xnor U13620 (N_13620,N_13075,N_13486);
or U13621 (N_13621,N_12836,N_13291);
or U13622 (N_13622,N_13185,N_13457);
or U13623 (N_13623,N_13043,N_13025);
nand U13624 (N_13624,N_13133,N_13414);
and U13625 (N_13625,N_13065,N_12892);
nand U13626 (N_13626,N_13033,N_13283);
or U13627 (N_13627,N_13520,N_13100);
nand U13628 (N_13628,N_13064,N_13103);
nor U13629 (N_13629,N_13050,N_13526);
and U13630 (N_13630,N_13183,N_13319);
nor U13631 (N_13631,N_12856,N_13228);
nand U13632 (N_13632,N_12969,N_12842);
or U13633 (N_13633,N_13428,N_12813);
nor U13634 (N_13634,N_13015,N_12946);
xnor U13635 (N_13635,N_13587,N_12989);
nand U13636 (N_13636,N_13076,N_13078);
nand U13637 (N_13637,N_13260,N_13342);
nor U13638 (N_13638,N_13431,N_13470);
xor U13639 (N_13639,N_13560,N_13533);
nand U13640 (N_13640,N_12855,N_12826);
nor U13641 (N_13641,N_13372,N_13597);
or U13642 (N_13642,N_12904,N_12845);
nand U13643 (N_13643,N_13555,N_13378);
nor U13644 (N_13644,N_13509,N_13275);
xor U13645 (N_13645,N_13224,N_13336);
and U13646 (N_13646,N_13455,N_13039);
xor U13647 (N_13647,N_13038,N_13472);
nand U13648 (N_13648,N_13365,N_13305);
or U13649 (N_13649,N_13121,N_13052);
or U13650 (N_13650,N_13101,N_13205);
nand U13651 (N_13651,N_13528,N_13123);
nand U13652 (N_13652,N_13408,N_13127);
and U13653 (N_13653,N_13281,N_13148);
nor U13654 (N_13654,N_13513,N_13529);
nor U13655 (N_13655,N_12966,N_12906);
nand U13656 (N_13656,N_12848,N_13215);
nor U13657 (N_13657,N_12939,N_13047);
xor U13658 (N_13658,N_13337,N_13292);
xor U13659 (N_13659,N_13232,N_13499);
and U13660 (N_13660,N_12970,N_12997);
and U13661 (N_13661,N_13347,N_12827);
nand U13662 (N_13662,N_13280,N_12956);
or U13663 (N_13663,N_13360,N_13174);
nand U13664 (N_13664,N_13034,N_13490);
nand U13665 (N_13665,N_13373,N_13494);
or U13666 (N_13666,N_12850,N_13487);
or U13667 (N_13667,N_13248,N_13432);
or U13668 (N_13668,N_13573,N_13036);
xor U13669 (N_13669,N_13599,N_12927);
nand U13670 (N_13670,N_12994,N_13221);
nor U13671 (N_13671,N_12990,N_13053);
xnor U13672 (N_13672,N_13069,N_13539);
nand U13673 (N_13673,N_13299,N_13188);
nor U13674 (N_13674,N_12869,N_13393);
xnor U13675 (N_13675,N_12887,N_13492);
nor U13676 (N_13676,N_12811,N_13094);
nand U13677 (N_13677,N_13014,N_13176);
xnor U13678 (N_13678,N_12901,N_12810);
and U13679 (N_13679,N_13430,N_13358);
nand U13680 (N_13680,N_13072,N_12871);
nor U13681 (N_13681,N_13104,N_13112);
nand U13682 (N_13682,N_13451,N_13289);
or U13683 (N_13683,N_12942,N_12922);
and U13684 (N_13684,N_13536,N_13161);
or U13685 (N_13685,N_13130,N_13054);
xnor U13686 (N_13686,N_13261,N_13368);
nand U13687 (N_13687,N_13265,N_13453);
nor U13688 (N_13688,N_13374,N_13550);
nor U13689 (N_13689,N_13315,N_12806);
or U13690 (N_13690,N_13556,N_13583);
or U13691 (N_13691,N_13538,N_13596);
or U13692 (N_13692,N_12841,N_12908);
xnor U13693 (N_13693,N_13341,N_13318);
nor U13694 (N_13694,N_13421,N_12935);
and U13695 (N_13695,N_12807,N_12870);
or U13696 (N_13696,N_13448,N_13197);
nand U13697 (N_13697,N_12928,N_13377);
nor U13698 (N_13698,N_13056,N_13357);
and U13699 (N_13699,N_12872,N_13225);
or U13700 (N_13700,N_13266,N_13353);
xnor U13701 (N_13701,N_13102,N_13207);
or U13702 (N_13702,N_13276,N_13153);
or U13703 (N_13703,N_13196,N_13137);
xor U13704 (N_13704,N_12857,N_12972);
nand U13705 (N_13705,N_13402,N_13376);
or U13706 (N_13706,N_13384,N_13000);
and U13707 (N_13707,N_13589,N_12920);
nor U13708 (N_13708,N_13206,N_13344);
nor U13709 (N_13709,N_12852,N_12963);
and U13710 (N_13710,N_12802,N_13331);
xnor U13711 (N_13711,N_13297,N_13375);
xor U13712 (N_13712,N_13516,N_13482);
nand U13713 (N_13713,N_13214,N_12821);
or U13714 (N_13714,N_13070,N_13298);
nand U13715 (N_13715,N_12853,N_13023);
nand U13716 (N_13716,N_13138,N_12912);
nand U13717 (N_13717,N_13592,N_13439);
or U13718 (N_13718,N_13416,N_13046);
and U13719 (N_13719,N_13060,N_13479);
xor U13720 (N_13720,N_13316,N_13150);
nor U13721 (N_13721,N_12921,N_13433);
and U13722 (N_13722,N_13349,N_13390);
and U13723 (N_13723,N_12834,N_13508);
xnor U13724 (N_13724,N_13145,N_13217);
and U13725 (N_13725,N_13302,N_13585);
nor U13726 (N_13726,N_13203,N_13535);
xnor U13727 (N_13727,N_13012,N_13122);
and U13728 (N_13728,N_13343,N_13417);
and U13729 (N_13729,N_13327,N_13495);
nor U13730 (N_13730,N_13170,N_13129);
nand U13731 (N_13731,N_12999,N_13243);
nand U13732 (N_13732,N_13011,N_13581);
nand U13733 (N_13733,N_13326,N_12977);
or U13734 (N_13734,N_13156,N_13022);
and U13735 (N_13735,N_12953,N_13147);
nand U13736 (N_13736,N_13568,N_13106);
or U13737 (N_13737,N_13186,N_12940);
or U13738 (N_13738,N_13048,N_12945);
xnor U13739 (N_13739,N_13537,N_13561);
nand U13740 (N_13740,N_13334,N_12982);
nor U13741 (N_13741,N_13531,N_13348);
and U13742 (N_13742,N_13481,N_13379);
nand U13743 (N_13743,N_12893,N_13410);
nor U13744 (N_13744,N_13018,N_13249);
or U13745 (N_13745,N_12910,N_13002);
xnor U13746 (N_13746,N_13158,N_13128);
and U13747 (N_13747,N_12898,N_13279);
xnor U13748 (N_13748,N_13030,N_12816);
or U13749 (N_13749,N_13167,N_13363);
nor U13750 (N_13750,N_12941,N_12964);
nor U13751 (N_13751,N_12992,N_13504);
nand U13752 (N_13752,N_13532,N_13165);
or U13753 (N_13753,N_13339,N_12874);
or U13754 (N_13754,N_12902,N_13422);
nand U13755 (N_13755,N_13252,N_13037);
xor U13756 (N_13756,N_12815,N_13144);
nand U13757 (N_13757,N_13219,N_13413);
xnor U13758 (N_13758,N_13577,N_12808);
nand U13759 (N_13759,N_12801,N_13338);
or U13760 (N_13760,N_12860,N_12986);
xor U13761 (N_13761,N_12916,N_13572);
or U13762 (N_13762,N_13089,N_13471);
nand U13763 (N_13763,N_12803,N_13149);
and U13764 (N_13764,N_13222,N_13233);
or U13765 (N_13765,N_13044,N_13062);
nand U13766 (N_13766,N_13051,N_13440);
nor U13767 (N_13767,N_13063,N_12867);
nand U13768 (N_13768,N_12883,N_13391);
and U13769 (N_13769,N_13152,N_13461);
nor U13770 (N_13770,N_12876,N_13093);
and U13771 (N_13771,N_13105,N_13006);
nand U13772 (N_13772,N_13534,N_13310);
nor U13773 (N_13773,N_13380,N_13445);
nor U13774 (N_13774,N_13009,N_13042);
and U13775 (N_13775,N_13595,N_12829);
nand U13776 (N_13776,N_13304,N_13115);
nor U13777 (N_13777,N_13201,N_13437);
nor U13778 (N_13778,N_13517,N_13356);
xnor U13779 (N_13779,N_13333,N_12885);
xor U13780 (N_13780,N_13518,N_13108);
or U13781 (N_13781,N_12975,N_13091);
nand U13782 (N_13782,N_13524,N_13540);
or U13783 (N_13783,N_13454,N_13090);
nand U13784 (N_13784,N_13488,N_13135);
and U13785 (N_13785,N_13352,N_13139);
nand U13786 (N_13786,N_12911,N_12907);
nor U13787 (N_13787,N_13067,N_13396);
and U13788 (N_13788,N_13085,N_12955);
nand U13789 (N_13789,N_12968,N_12881);
xor U13790 (N_13790,N_13313,N_13452);
nor U13791 (N_13791,N_13370,N_13095);
nor U13792 (N_13792,N_13286,N_13371);
xor U13793 (N_13793,N_12894,N_13171);
and U13794 (N_13794,N_13111,N_13512);
or U13795 (N_13795,N_13411,N_13296);
nor U13796 (N_13796,N_13155,N_13546);
and U13797 (N_13797,N_13558,N_13335);
xor U13798 (N_13798,N_13119,N_13394);
xnor U13799 (N_13799,N_12913,N_13542);
xor U13800 (N_13800,N_13098,N_13026);
xor U13801 (N_13801,N_13480,N_12879);
xnor U13802 (N_13802,N_12996,N_13211);
xnor U13803 (N_13803,N_13501,N_13593);
nand U13804 (N_13804,N_13551,N_13590);
or U13805 (N_13805,N_13456,N_13184);
or U13806 (N_13806,N_12900,N_13541);
and U13807 (N_13807,N_12847,N_13463);
or U13808 (N_13808,N_13476,N_13013);
nand U13809 (N_13809,N_13199,N_13057);
or U13810 (N_13810,N_13388,N_13055);
nor U13811 (N_13811,N_13162,N_13146);
and U13812 (N_13812,N_13449,N_13303);
xor U13813 (N_13813,N_13191,N_12983);
and U13814 (N_13814,N_13465,N_13317);
nand U13815 (N_13815,N_13506,N_13180);
or U13816 (N_13816,N_13588,N_13245);
xnor U13817 (N_13817,N_13141,N_13255);
or U13818 (N_13818,N_13273,N_13157);
and U13819 (N_13819,N_13464,N_13125);
or U13820 (N_13820,N_12978,N_13567);
xnor U13821 (N_13821,N_13446,N_13350);
xor U13822 (N_13822,N_12882,N_12909);
and U13823 (N_13823,N_13574,N_13271);
nor U13824 (N_13824,N_13239,N_13061);
nand U13825 (N_13825,N_13311,N_13213);
nor U13826 (N_13826,N_12838,N_13359);
nor U13827 (N_13827,N_13362,N_13418);
or U13828 (N_13828,N_13256,N_13383);
nand U13829 (N_13829,N_13351,N_13322);
or U13830 (N_13830,N_13591,N_13385);
or U13831 (N_13831,N_13354,N_13016);
and U13832 (N_13832,N_13126,N_12886);
nor U13833 (N_13833,N_12903,N_12915);
xor U13834 (N_13834,N_13500,N_13309);
and U13835 (N_13835,N_12995,N_13290);
and U13836 (N_13836,N_12812,N_13515);
xor U13837 (N_13837,N_13080,N_12831);
nor U13838 (N_13838,N_13132,N_13216);
nand U13839 (N_13839,N_12957,N_13493);
nor U13840 (N_13840,N_12897,N_13272);
and U13841 (N_13841,N_13569,N_12931);
xor U13842 (N_13842,N_12817,N_13460);
and U13843 (N_13843,N_13443,N_13345);
and U13844 (N_13844,N_13522,N_12923);
or U13845 (N_13845,N_12985,N_13278);
and U13846 (N_13846,N_13552,N_12974);
and U13847 (N_13847,N_13229,N_13116);
nor U13848 (N_13848,N_13204,N_12822);
nand U13849 (N_13849,N_13307,N_13187);
nor U13850 (N_13850,N_13114,N_13441);
nand U13851 (N_13851,N_13074,N_13077);
and U13852 (N_13852,N_13004,N_12880);
xnor U13853 (N_13853,N_13008,N_12950);
xor U13854 (N_13854,N_13478,N_13092);
xnor U13855 (N_13855,N_12971,N_12828);
nand U13856 (N_13856,N_13267,N_12868);
nor U13857 (N_13857,N_12839,N_12830);
and U13858 (N_13858,N_13401,N_13328);
and U13859 (N_13859,N_13200,N_12919);
or U13860 (N_13860,N_13598,N_13284);
nor U13861 (N_13861,N_13447,N_13467);
and U13862 (N_13862,N_13330,N_12865);
nor U13863 (N_13863,N_12981,N_12973);
xnor U13864 (N_13864,N_13027,N_13295);
nor U13865 (N_13865,N_13566,N_13172);
nand U13866 (N_13866,N_12884,N_13124);
nor U13867 (N_13867,N_12889,N_12840);
xor U13868 (N_13868,N_12851,N_12846);
nor U13869 (N_13869,N_13110,N_12899);
and U13870 (N_13870,N_13325,N_13088);
or U13871 (N_13871,N_12936,N_13389);
nor U13872 (N_13872,N_13293,N_12962);
nand U13873 (N_13873,N_13525,N_13579);
nand U13874 (N_13874,N_13361,N_12987);
nand U13875 (N_13875,N_13163,N_13179);
nand U13876 (N_13876,N_12862,N_13270);
nand U13877 (N_13877,N_12858,N_13282);
nand U13878 (N_13878,N_13575,N_13355);
nor U13879 (N_13879,N_12804,N_12832);
nand U13880 (N_13880,N_13469,N_12805);
xor U13881 (N_13881,N_13079,N_13240);
or U13882 (N_13882,N_12959,N_13068);
or U13883 (N_13883,N_13007,N_13160);
nor U13884 (N_13884,N_13570,N_12814);
nand U13885 (N_13885,N_13314,N_13523);
xnor U13886 (N_13886,N_13466,N_12864);
nor U13887 (N_13887,N_13107,N_13192);
and U13888 (N_13888,N_13058,N_12896);
and U13889 (N_13889,N_13143,N_13017);
nor U13890 (N_13890,N_12809,N_13511);
nor U13891 (N_13891,N_13140,N_13423);
nand U13892 (N_13892,N_13329,N_13496);
nor U13893 (N_13893,N_13586,N_13226);
nor U13894 (N_13894,N_13510,N_13369);
nand U13895 (N_13895,N_13244,N_13241);
nand U13896 (N_13896,N_13117,N_13190);
nand U13897 (N_13897,N_12937,N_12948);
xnor U13898 (N_13898,N_13519,N_13262);
and U13899 (N_13899,N_13288,N_13300);
and U13900 (N_13900,N_13565,N_12895);
nor U13901 (N_13901,N_13426,N_13435);
and U13902 (N_13902,N_13242,N_13468);
nand U13903 (N_13903,N_13210,N_12967);
or U13904 (N_13904,N_13407,N_13491);
or U13905 (N_13905,N_13198,N_12951);
xor U13906 (N_13906,N_13045,N_13594);
or U13907 (N_13907,N_13547,N_13436);
nor U13908 (N_13908,N_13381,N_13475);
or U13909 (N_13909,N_13208,N_13505);
nor U13910 (N_13910,N_13169,N_13159);
or U13911 (N_13911,N_12861,N_13086);
nand U13912 (N_13912,N_13029,N_13154);
nor U13913 (N_13913,N_13415,N_13120);
xnor U13914 (N_13914,N_13312,N_13412);
xor U13915 (N_13915,N_13563,N_13032);
nand U13916 (N_13916,N_12944,N_13366);
xnor U13917 (N_13917,N_13497,N_12938);
xor U13918 (N_13918,N_13473,N_13301);
nor U13919 (N_13919,N_13521,N_12873);
or U13920 (N_13920,N_13306,N_12933);
nor U13921 (N_13921,N_12926,N_12932);
and U13922 (N_13922,N_13227,N_13514);
nand U13923 (N_13923,N_13251,N_12866);
xor U13924 (N_13924,N_12820,N_13582);
nor U13925 (N_13925,N_12917,N_13285);
nand U13926 (N_13926,N_13553,N_13166);
or U13927 (N_13927,N_13118,N_13175);
xor U13928 (N_13928,N_13136,N_13259);
nand U13929 (N_13929,N_13236,N_13202);
nand U13930 (N_13930,N_12914,N_13405);
nand U13931 (N_13931,N_13066,N_13571);
or U13932 (N_13932,N_13087,N_13459);
nor U13933 (N_13933,N_13164,N_13194);
xor U13934 (N_13934,N_13073,N_12965);
xor U13935 (N_13935,N_12818,N_12891);
or U13936 (N_13936,N_12947,N_13489);
nand U13937 (N_13937,N_13545,N_13576);
nand U13938 (N_13938,N_13173,N_13562);
nand U13939 (N_13939,N_13543,N_12952);
nand U13940 (N_13940,N_12980,N_13250);
nor U13941 (N_13941,N_13257,N_12934);
nor U13942 (N_13942,N_13382,N_13477);
xnor U13943 (N_13943,N_13580,N_13181);
nor U13944 (N_13944,N_13028,N_13308);
and U13945 (N_13945,N_13021,N_13005);
and U13946 (N_13946,N_13177,N_13321);
nand U13947 (N_13947,N_13409,N_13209);
xor U13948 (N_13948,N_13220,N_13134);
nor U13949 (N_13949,N_13059,N_13218);
nand U13950 (N_13950,N_12835,N_13019);
nor U13951 (N_13951,N_13530,N_13189);
or U13952 (N_13952,N_13182,N_13264);
or U13953 (N_13953,N_12960,N_13404);
and U13954 (N_13954,N_13403,N_12998);
or U13955 (N_13955,N_13195,N_13247);
nand U13956 (N_13956,N_12991,N_13458);
nor U13957 (N_13957,N_13364,N_13420);
nand U13958 (N_13958,N_12954,N_12859);
or U13959 (N_13959,N_12976,N_13484);
and U13960 (N_13960,N_13178,N_13294);
and U13961 (N_13961,N_13474,N_12843);
xor U13962 (N_13962,N_13151,N_12844);
nor U13963 (N_13963,N_13096,N_13462);
nor U13964 (N_13964,N_13554,N_13392);
or U13965 (N_13965,N_12993,N_13502);
nand U13966 (N_13966,N_12943,N_13557);
or U13967 (N_13967,N_13113,N_13564);
or U13968 (N_13968,N_13263,N_13274);
nor U13969 (N_13969,N_13527,N_12837);
or U13970 (N_13970,N_12924,N_13507);
or U13971 (N_13971,N_13084,N_12849);
and U13972 (N_13972,N_13131,N_12863);
nor U13973 (N_13973,N_13010,N_13223);
and U13974 (N_13974,N_13438,N_12918);
or U13975 (N_13975,N_13332,N_13024);
or U13976 (N_13976,N_13323,N_12819);
or U13977 (N_13977,N_12823,N_13548);
nor U13978 (N_13978,N_13020,N_12825);
and U13979 (N_13979,N_13320,N_13254);
nand U13980 (N_13980,N_13398,N_12888);
nor U13981 (N_13981,N_13406,N_12800);
and U13982 (N_13982,N_13559,N_13235);
nor U13983 (N_13983,N_13400,N_13584);
and U13984 (N_13984,N_13003,N_13578);
xor U13985 (N_13985,N_13269,N_13395);
and U13986 (N_13986,N_13434,N_13049);
nor U13987 (N_13987,N_13549,N_12929);
and U13988 (N_13988,N_13419,N_12958);
nor U13989 (N_13989,N_13031,N_13082);
xor U13990 (N_13990,N_13544,N_13193);
xor U13991 (N_13991,N_13238,N_13253);
nor U13992 (N_13992,N_12854,N_13498);
or U13993 (N_13993,N_13099,N_13081);
or U13994 (N_13994,N_13386,N_13001);
and U13995 (N_13995,N_12824,N_13035);
nor U13996 (N_13996,N_13397,N_12988);
xor U13997 (N_13997,N_13071,N_13503);
or U13998 (N_13998,N_13483,N_13450);
and U13999 (N_13999,N_13424,N_12984);
xor U14000 (N_14000,N_13240,N_13064);
nand U14001 (N_14001,N_13121,N_13013);
xnor U14002 (N_14002,N_13572,N_13471);
and U14003 (N_14003,N_13248,N_13132);
and U14004 (N_14004,N_12873,N_13534);
xnor U14005 (N_14005,N_13302,N_13366);
and U14006 (N_14006,N_12873,N_13133);
and U14007 (N_14007,N_13008,N_13057);
and U14008 (N_14008,N_12804,N_13197);
nand U14009 (N_14009,N_13472,N_12877);
nand U14010 (N_14010,N_13128,N_12832);
xor U14011 (N_14011,N_12883,N_13081);
and U14012 (N_14012,N_13516,N_13339);
and U14013 (N_14013,N_13175,N_13401);
nand U14014 (N_14014,N_13409,N_13143);
and U14015 (N_14015,N_13142,N_13460);
nor U14016 (N_14016,N_13139,N_12893);
nand U14017 (N_14017,N_12835,N_13374);
nor U14018 (N_14018,N_13157,N_13145);
nor U14019 (N_14019,N_12982,N_13553);
nor U14020 (N_14020,N_13517,N_13116);
nor U14021 (N_14021,N_13147,N_13240);
xnor U14022 (N_14022,N_13081,N_12927);
xor U14023 (N_14023,N_12980,N_13328);
nor U14024 (N_14024,N_13064,N_13579);
nor U14025 (N_14025,N_13071,N_12844);
nor U14026 (N_14026,N_12870,N_12996);
nor U14027 (N_14027,N_13434,N_13016);
nor U14028 (N_14028,N_13310,N_13112);
nand U14029 (N_14029,N_13517,N_12951);
or U14030 (N_14030,N_13528,N_12937);
nor U14031 (N_14031,N_12850,N_12817);
nand U14032 (N_14032,N_13304,N_13018);
and U14033 (N_14033,N_13458,N_13404);
nor U14034 (N_14034,N_13588,N_12884);
xnor U14035 (N_14035,N_12850,N_13053);
nand U14036 (N_14036,N_12992,N_13191);
nor U14037 (N_14037,N_13047,N_12941);
nand U14038 (N_14038,N_12877,N_12907);
xnor U14039 (N_14039,N_12801,N_13350);
and U14040 (N_14040,N_13445,N_13115);
or U14041 (N_14041,N_13274,N_12818);
nor U14042 (N_14042,N_13379,N_13156);
and U14043 (N_14043,N_13538,N_13121);
or U14044 (N_14044,N_12971,N_13138);
and U14045 (N_14045,N_13198,N_12946);
and U14046 (N_14046,N_13110,N_13454);
xnor U14047 (N_14047,N_12928,N_13042);
nor U14048 (N_14048,N_13274,N_13327);
and U14049 (N_14049,N_13126,N_12828);
or U14050 (N_14050,N_13097,N_13213);
or U14051 (N_14051,N_13502,N_13450);
nand U14052 (N_14052,N_13089,N_13569);
or U14053 (N_14053,N_13255,N_13341);
nand U14054 (N_14054,N_13178,N_13258);
xor U14055 (N_14055,N_13258,N_13031);
or U14056 (N_14056,N_13432,N_13057);
nand U14057 (N_14057,N_13439,N_13052);
nand U14058 (N_14058,N_13018,N_13594);
and U14059 (N_14059,N_13394,N_13437);
nand U14060 (N_14060,N_13464,N_12802);
nand U14061 (N_14061,N_13568,N_12979);
and U14062 (N_14062,N_12845,N_12850);
xor U14063 (N_14063,N_12885,N_13053);
xnor U14064 (N_14064,N_12985,N_13010);
nand U14065 (N_14065,N_13354,N_13267);
or U14066 (N_14066,N_13309,N_13334);
or U14067 (N_14067,N_12924,N_12986);
and U14068 (N_14068,N_13042,N_13391);
xor U14069 (N_14069,N_13032,N_13365);
and U14070 (N_14070,N_13387,N_13391);
or U14071 (N_14071,N_13124,N_13041);
nor U14072 (N_14072,N_13233,N_13002);
or U14073 (N_14073,N_13324,N_13313);
and U14074 (N_14074,N_13002,N_13288);
xor U14075 (N_14075,N_13354,N_13336);
and U14076 (N_14076,N_13109,N_13241);
nor U14077 (N_14077,N_13459,N_12936);
and U14078 (N_14078,N_13089,N_12868);
and U14079 (N_14079,N_13095,N_12903);
or U14080 (N_14080,N_12843,N_13279);
or U14081 (N_14081,N_13225,N_13451);
xor U14082 (N_14082,N_13251,N_12997);
nor U14083 (N_14083,N_13534,N_13455);
nor U14084 (N_14084,N_13000,N_13283);
xnor U14085 (N_14085,N_13385,N_13080);
nand U14086 (N_14086,N_12811,N_13128);
nand U14087 (N_14087,N_13584,N_13597);
nor U14088 (N_14088,N_13506,N_13285);
xnor U14089 (N_14089,N_12805,N_13136);
nor U14090 (N_14090,N_13550,N_13147);
nand U14091 (N_14091,N_13070,N_13069);
xnor U14092 (N_14092,N_13027,N_13418);
nor U14093 (N_14093,N_13335,N_13167);
and U14094 (N_14094,N_13397,N_13004);
nor U14095 (N_14095,N_12913,N_13265);
or U14096 (N_14096,N_13448,N_13458);
xnor U14097 (N_14097,N_13255,N_13110);
xor U14098 (N_14098,N_13415,N_13071);
nor U14099 (N_14099,N_13596,N_12972);
and U14100 (N_14100,N_13047,N_13021);
nand U14101 (N_14101,N_12969,N_12868);
nand U14102 (N_14102,N_12966,N_13339);
xor U14103 (N_14103,N_12987,N_13537);
xnor U14104 (N_14104,N_13322,N_13131);
xor U14105 (N_14105,N_12920,N_13576);
and U14106 (N_14106,N_13589,N_13120);
and U14107 (N_14107,N_13566,N_13011);
xor U14108 (N_14108,N_12812,N_13309);
nand U14109 (N_14109,N_13444,N_13270);
and U14110 (N_14110,N_13152,N_12853);
or U14111 (N_14111,N_13325,N_13427);
nand U14112 (N_14112,N_13412,N_13324);
nand U14113 (N_14113,N_13398,N_13465);
or U14114 (N_14114,N_13189,N_13163);
and U14115 (N_14115,N_13161,N_13220);
nor U14116 (N_14116,N_13009,N_13372);
nor U14117 (N_14117,N_13013,N_13431);
or U14118 (N_14118,N_12938,N_13024);
nand U14119 (N_14119,N_13543,N_13442);
or U14120 (N_14120,N_13446,N_12869);
nor U14121 (N_14121,N_12904,N_13037);
nand U14122 (N_14122,N_12995,N_12890);
or U14123 (N_14123,N_12918,N_12933);
xor U14124 (N_14124,N_13520,N_13531);
and U14125 (N_14125,N_13399,N_12827);
xnor U14126 (N_14126,N_13499,N_13581);
or U14127 (N_14127,N_13133,N_13527);
nor U14128 (N_14128,N_12953,N_12831);
nand U14129 (N_14129,N_13550,N_13494);
nor U14130 (N_14130,N_13055,N_12957);
nor U14131 (N_14131,N_13242,N_13047);
xnor U14132 (N_14132,N_13409,N_13571);
nand U14133 (N_14133,N_13190,N_13540);
xnor U14134 (N_14134,N_13344,N_12852);
xor U14135 (N_14135,N_13267,N_13190);
nor U14136 (N_14136,N_13205,N_12801);
nor U14137 (N_14137,N_13071,N_13125);
nand U14138 (N_14138,N_13352,N_13333);
and U14139 (N_14139,N_13162,N_13069);
xor U14140 (N_14140,N_13447,N_12929);
xor U14141 (N_14141,N_12964,N_13385);
xnor U14142 (N_14142,N_13437,N_12852);
xnor U14143 (N_14143,N_12966,N_13045);
or U14144 (N_14144,N_13266,N_13567);
xnor U14145 (N_14145,N_12944,N_13208);
and U14146 (N_14146,N_13191,N_13142);
nor U14147 (N_14147,N_12970,N_13472);
xnor U14148 (N_14148,N_13205,N_13228);
and U14149 (N_14149,N_12951,N_13469);
xnor U14150 (N_14150,N_12895,N_13261);
nand U14151 (N_14151,N_13484,N_13152);
nor U14152 (N_14152,N_13059,N_13586);
nor U14153 (N_14153,N_13597,N_13196);
and U14154 (N_14154,N_13211,N_13227);
and U14155 (N_14155,N_13257,N_13374);
and U14156 (N_14156,N_12871,N_13374);
or U14157 (N_14157,N_12931,N_13270);
nand U14158 (N_14158,N_12850,N_12880);
nor U14159 (N_14159,N_13276,N_13047);
or U14160 (N_14160,N_12869,N_13083);
xnor U14161 (N_14161,N_13078,N_12913);
or U14162 (N_14162,N_13308,N_13551);
nand U14163 (N_14163,N_13085,N_13248);
or U14164 (N_14164,N_13295,N_13599);
and U14165 (N_14165,N_13482,N_13588);
xor U14166 (N_14166,N_13066,N_13565);
or U14167 (N_14167,N_13202,N_13534);
nand U14168 (N_14168,N_13385,N_13310);
nand U14169 (N_14169,N_12915,N_12948);
xor U14170 (N_14170,N_13459,N_13078);
and U14171 (N_14171,N_12945,N_13274);
xnor U14172 (N_14172,N_12884,N_13202);
or U14173 (N_14173,N_13491,N_12951);
xor U14174 (N_14174,N_13353,N_13009);
nand U14175 (N_14175,N_13159,N_13114);
xnor U14176 (N_14176,N_13479,N_13356);
or U14177 (N_14177,N_13310,N_13242);
xor U14178 (N_14178,N_13247,N_13535);
and U14179 (N_14179,N_13292,N_13093);
nand U14180 (N_14180,N_13058,N_13198);
or U14181 (N_14181,N_13267,N_12888);
nor U14182 (N_14182,N_13441,N_13190);
nand U14183 (N_14183,N_12888,N_13364);
xor U14184 (N_14184,N_13248,N_13500);
nand U14185 (N_14185,N_12954,N_12893);
nand U14186 (N_14186,N_12955,N_13438);
nor U14187 (N_14187,N_12842,N_13550);
and U14188 (N_14188,N_13162,N_13260);
nand U14189 (N_14189,N_13298,N_12920);
nor U14190 (N_14190,N_13156,N_12920);
nor U14191 (N_14191,N_13395,N_12941);
and U14192 (N_14192,N_13415,N_12891);
nor U14193 (N_14193,N_13339,N_13104);
and U14194 (N_14194,N_13534,N_13053);
and U14195 (N_14195,N_12912,N_13504);
nand U14196 (N_14196,N_12859,N_12910);
or U14197 (N_14197,N_13394,N_13469);
nand U14198 (N_14198,N_13068,N_13295);
xnor U14199 (N_14199,N_12932,N_13219);
or U14200 (N_14200,N_13363,N_13452);
and U14201 (N_14201,N_13444,N_12990);
and U14202 (N_14202,N_13258,N_12833);
nand U14203 (N_14203,N_13481,N_13429);
xnor U14204 (N_14204,N_13117,N_13415);
or U14205 (N_14205,N_13127,N_13475);
xnor U14206 (N_14206,N_13346,N_13060);
nor U14207 (N_14207,N_13497,N_13214);
and U14208 (N_14208,N_12834,N_13511);
nand U14209 (N_14209,N_12993,N_13056);
xor U14210 (N_14210,N_12841,N_13529);
nor U14211 (N_14211,N_12815,N_12992);
or U14212 (N_14212,N_13237,N_13410);
or U14213 (N_14213,N_13498,N_13405);
nand U14214 (N_14214,N_13047,N_13096);
nand U14215 (N_14215,N_13082,N_12923);
nor U14216 (N_14216,N_13199,N_12952);
xor U14217 (N_14217,N_12956,N_13537);
nand U14218 (N_14218,N_12807,N_13532);
nor U14219 (N_14219,N_12918,N_12984);
or U14220 (N_14220,N_13224,N_12929);
and U14221 (N_14221,N_13184,N_13501);
or U14222 (N_14222,N_13193,N_13586);
or U14223 (N_14223,N_12941,N_13445);
xnor U14224 (N_14224,N_13338,N_13082);
and U14225 (N_14225,N_12993,N_13214);
and U14226 (N_14226,N_12937,N_13590);
or U14227 (N_14227,N_13066,N_13315);
or U14228 (N_14228,N_13443,N_12803);
nand U14229 (N_14229,N_13523,N_13133);
nor U14230 (N_14230,N_12875,N_13025);
and U14231 (N_14231,N_13350,N_12938);
nor U14232 (N_14232,N_13209,N_13312);
nand U14233 (N_14233,N_13455,N_13000);
nand U14234 (N_14234,N_13592,N_13546);
or U14235 (N_14235,N_12830,N_13127);
or U14236 (N_14236,N_13256,N_13051);
nor U14237 (N_14237,N_12826,N_13339);
xnor U14238 (N_14238,N_13345,N_12983);
or U14239 (N_14239,N_12859,N_13383);
xor U14240 (N_14240,N_13088,N_12877);
and U14241 (N_14241,N_13176,N_13068);
nand U14242 (N_14242,N_13467,N_13527);
and U14243 (N_14243,N_13053,N_13431);
nor U14244 (N_14244,N_12991,N_13170);
and U14245 (N_14245,N_13540,N_13207);
xnor U14246 (N_14246,N_13586,N_12931);
nand U14247 (N_14247,N_13591,N_12980);
xnor U14248 (N_14248,N_13407,N_13154);
and U14249 (N_14249,N_13136,N_12824);
nand U14250 (N_14250,N_13208,N_13044);
and U14251 (N_14251,N_13414,N_13275);
nand U14252 (N_14252,N_13476,N_13113);
xor U14253 (N_14253,N_13496,N_13134);
or U14254 (N_14254,N_13251,N_13443);
nor U14255 (N_14255,N_13028,N_13173);
nand U14256 (N_14256,N_13409,N_12971);
xor U14257 (N_14257,N_13122,N_13326);
and U14258 (N_14258,N_12923,N_13025);
nand U14259 (N_14259,N_13531,N_13086);
nor U14260 (N_14260,N_13078,N_13230);
or U14261 (N_14261,N_13164,N_13063);
nand U14262 (N_14262,N_13239,N_13070);
and U14263 (N_14263,N_12930,N_13516);
nand U14264 (N_14264,N_12814,N_13313);
nand U14265 (N_14265,N_12965,N_13205);
and U14266 (N_14266,N_13376,N_13541);
or U14267 (N_14267,N_13571,N_12936);
xor U14268 (N_14268,N_13572,N_13093);
nor U14269 (N_14269,N_12827,N_12891);
xor U14270 (N_14270,N_13437,N_13507);
xor U14271 (N_14271,N_12918,N_13089);
nor U14272 (N_14272,N_13042,N_13385);
or U14273 (N_14273,N_12813,N_12963);
and U14274 (N_14274,N_13500,N_12995);
nand U14275 (N_14275,N_13232,N_13106);
or U14276 (N_14276,N_13102,N_13199);
nand U14277 (N_14277,N_13515,N_13233);
nand U14278 (N_14278,N_13350,N_13004);
or U14279 (N_14279,N_12851,N_13458);
and U14280 (N_14280,N_13514,N_13281);
or U14281 (N_14281,N_13481,N_13145);
xor U14282 (N_14282,N_13310,N_13156);
nand U14283 (N_14283,N_13584,N_12945);
xnor U14284 (N_14284,N_12826,N_13397);
xor U14285 (N_14285,N_13541,N_13452);
nor U14286 (N_14286,N_12803,N_13390);
xor U14287 (N_14287,N_13195,N_13597);
and U14288 (N_14288,N_13340,N_13270);
and U14289 (N_14289,N_13022,N_13254);
or U14290 (N_14290,N_12804,N_13217);
nor U14291 (N_14291,N_13006,N_13214);
nor U14292 (N_14292,N_13592,N_13335);
xor U14293 (N_14293,N_13037,N_13391);
xor U14294 (N_14294,N_13092,N_13030);
or U14295 (N_14295,N_13449,N_13537);
nand U14296 (N_14296,N_13556,N_13551);
nor U14297 (N_14297,N_12983,N_12986);
or U14298 (N_14298,N_13158,N_13014);
nand U14299 (N_14299,N_12914,N_12854);
or U14300 (N_14300,N_13496,N_13205);
or U14301 (N_14301,N_13350,N_13032);
and U14302 (N_14302,N_12837,N_13451);
and U14303 (N_14303,N_13446,N_13001);
and U14304 (N_14304,N_13424,N_13156);
or U14305 (N_14305,N_12878,N_13500);
nor U14306 (N_14306,N_13253,N_13103);
or U14307 (N_14307,N_12889,N_12957);
nand U14308 (N_14308,N_12949,N_12958);
nor U14309 (N_14309,N_13568,N_12812);
and U14310 (N_14310,N_13156,N_13212);
nor U14311 (N_14311,N_13573,N_13541);
or U14312 (N_14312,N_13197,N_12882);
and U14313 (N_14313,N_13101,N_13586);
xor U14314 (N_14314,N_13113,N_13233);
xor U14315 (N_14315,N_13097,N_13352);
or U14316 (N_14316,N_13296,N_13373);
nor U14317 (N_14317,N_13403,N_13139);
xor U14318 (N_14318,N_13147,N_12869);
xnor U14319 (N_14319,N_13207,N_13274);
or U14320 (N_14320,N_13218,N_12845);
nand U14321 (N_14321,N_13372,N_13016);
xnor U14322 (N_14322,N_12935,N_13404);
or U14323 (N_14323,N_13102,N_12931);
or U14324 (N_14324,N_13479,N_12968);
or U14325 (N_14325,N_13191,N_13168);
nand U14326 (N_14326,N_13206,N_13064);
or U14327 (N_14327,N_13275,N_12836);
or U14328 (N_14328,N_12921,N_13003);
nand U14329 (N_14329,N_13003,N_12879);
nor U14330 (N_14330,N_13226,N_13203);
nor U14331 (N_14331,N_12962,N_13269);
nor U14332 (N_14332,N_12816,N_13578);
and U14333 (N_14333,N_13173,N_13315);
nor U14334 (N_14334,N_12992,N_12970);
xnor U14335 (N_14335,N_13324,N_13333);
or U14336 (N_14336,N_13376,N_13035);
and U14337 (N_14337,N_12834,N_13518);
nor U14338 (N_14338,N_13205,N_12925);
nand U14339 (N_14339,N_13338,N_12866);
nand U14340 (N_14340,N_13005,N_12981);
nand U14341 (N_14341,N_13323,N_13283);
xnor U14342 (N_14342,N_13569,N_13193);
or U14343 (N_14343,N_13504,N_13023);
nand U14344 (N_14344,N_13550,N_13493);
and U14345 (N_14345,N_13421,N_13084);
nor U14346 (N_14346,N_13125,N_13577);
nor U14347 (N_14347,N_13103,N_13340);
xor U14348 (N_14348,N_12920,N_13436);
nand U14349 (N_14349,N_13100,N_13088);
and U14350 (N_14350,N_13093,N_13072);
nor U14351 (N_14351,N_13020,N_13236);
and U14352 (N_14352,N_12951,N_13128);
and U14353 (N_14353,N_12874,N_12995);
nand U14354 (N_14354,N_13201,N_12938);
nand U14355 (N_14355,N_13430,N_13245);
nor U14356 (N_14356,N_13578,N_13217);
nand U14357 (N_14357,N_13164,N_13577);
and U14358 (N_14358,N_13180,N_13245);
and U14359 (N_14359,N_13327,N_12910);
xnor U14360 (N_14360,N_13551,N_12951);
nor U14361 (N_14361,N_13464,N_12926);
nor U14362 (N_14362,N_13155,N_13440);
xor U14363 (N_14363,N_13173,N_13296);
nor U14364 (N_14364,N_13149,N_13459);
nand U14365 (N_14365,N_13190,N_13001);
nand U14366 (N_14366,N_13231,N_13110);
nor U14367 (N_14367,N_13356,N_13332);
xor U14368 (N_14368,N_13105,N_13306);
nand U14369 (N_14369,N_13555,N_13338);
or U14370 (N_14370,N_13127,N_13536);
and U14371 (N_14371,N_13122,N_13469);
or U14372 (N_14372,N_12835,N_13463);
or U14373 (N_14373,N_12877,N_13220);
and U14374 (N_14374,N_13404,N_13029);
and U14375 (N_14375,N_12942,N_13163);
or U14376 (N_14376,N_13441,N_13378);
nor U14377 (N_14377,N_13121,N_13453);
nand U14378 (N_14378,N_12893,N_13112);
nand U14379 (N_14379,N_13395,N_13230);
or U14380 (N_14380,N_13164,N_13227);
nor U14381 (N_14381,N_13437,N_12876);
nor U14382 (N_14382,N_13241,N_13415);
and U14383 (N_14383,N_13515,N_13512);
nand U14384 (N_14384,N_12994,N_13568);
nand U14385 (N_14385,N_13404,N_13179);
nand U14386 (N_14386,N_13181,N_13195);
or U14387 (N_14387,N_12991,N_12987);
and U14388 (N_14388,N_12833,N_13285);
nand U14389 (N_14389,N_13254,N_13474);
xor U14390 (N_14390,N_13126,N_13255);
xnor U14391 (N_14391,N_13304,N_13584);
nand U14392 (N_14392,N_13472,N_13023);
nand U14393 (N_14393,N_13300,N_13012);
or U14394 (N_14394,N_12821,N_12833);
and U14395 (N_14395,N_13516,N_13441);
xnor U14396 (N_14396,N_13310,N_13015);
or U14397 (N_14397,N_12946,N_12824);
nand U14398 (N_14398,N_13222,N_13546);
or U14399 (N_14399,N_13410,N_13107);
or U14400 (N_14400,N_13849,N_13951);
or U14401 (N_14401,N_14289,N_14067);
nand U14402 (N_14402,N_14329,N_14114);
or U14403 (N_14403,N_14059,N_13611);
xor U14404 (N_14404,N_14383,N_13927);
xnor U14405 (N_14405,N_14180,N_14264);
nor U14406 (N_14406,N_13846,N_13601);
or U14407 (N_14407,N_13856,N_14094);
or U14408 (N_14408,N_14200,N_14163);
and U14409 (N_14409,N_13833,N_14013);
or U14410 (N_14410,N_13776,N_13817);
and U14411 (N_14411,N_14070,N_14288);
nand U14412 (N_14412,N_14224,N_13991);
and U14413 (N_14413,N_13753,N_13639);
and U14414 (N_14414,N_14285,N_14321);
nor U14415 (N_14415,N_13969,N_14023);
xor U14416 (N_14416,N_13735,N_13892);
nand U14417 (N_14417,N_14053,N_13744);
nor U14418 (N_14418,N_14294,N_14269);
xor U14419 (N_14419,N_13617,N_13809);
nor U14420 (N_14420,N_13997,N_14122);
nor U14421 (N_14421,N_13871,N_13768);
nand U14422 (N_14422,N_13815,N_13677);
nand U14423 (N_14423,N_14325,N_13836);
and U14424 (N_14424,N_14108,N_13612);
xor U14425 (N_14425,N_14092,N_14002);
or U14426 (N_14426,N_14334,N_13886);
or U14427 (N_14427,N_13908,N_14253);
xor U14428 (N_14428,N_13700,N_14054);
nor U14429 (N_14429,N_13681,N_14076);
or U14430 (N_14430,N_13780,N_13995);
and U14431 (N_14431,N_14035,N_14185);
or U14432 (N_14432,N_14365,N_13979);
nor U14433 (N_14433,N_13747,N_13878);
nand U14434 (N_14434,N_14102,N_14063);
or U14435 (N_14435,N_13936,N_14368);
or U14436 (N_14436,N_13767,N_14322);
nor U14437 (N_14437,N_13715,N_13873);
and U14438 (N_14438,N_13933,N_14215);
xnor U14439 (N_14439,N_14195,N_14256);
nand U14440 (N_14440,N_14111,N_14352);
and U14441 (N_14441,N_14207,N_13674);
and U14442 (N_14442,N_13689,N_13982);
nor U14443 (N_14443,N_14015,N_14228);
nand U14444 (N_14444,N_14326,N_13930);
nand U14445 (N_14445,N_14193,N_13801);
and U14446 (N_14446,N_14065,N_14171);
or U14447 (N_14447,N_14226,N_13786);
or U14448 (N_14448,N_14296,N_14240);
xor U14449 (N_14449,N_14081,N_14379);
nand U14450 (N_14450,N_13762,N_13778);
nor U14451 (N_14451,N_13822,N_14051);
nand U14452 (N_14452,N_14041,N_14055);
and U14453 (N_14453,N_14276,N_14258);
and U14454 (N_14454,N_13882,N_14290);
nor U14455 (N_14455,N_13692,N_13678);
nand U14456 (N_14456,N_14179,N_13726);
xor U14457 (N_14457,N_13804,N_14007);
and U14458 (N_14458,N_14223,N_14271);
and U14459 (N_14459,N_14221,N_14087);
nor U14460 (N_14460,N_13918,N_13683);
or U14461 (N_14461,N_14110,N_14214);
nor U14462 (N_14462,N_14170,N_14231);
and U14463 (N_14463,N_13665,N_13967);
nand U14464 (N_14464,N_13920,N_13769);
nand U14465 (N_14465,N_13713,N_13740);
or U14466 (N_14466,N_13895,N_13759);
nor U14467 (N_14467,N_14026,N_13999);
or U14468 (N_14468,N_13657,N_14299);
or U14469 (N_14469,N_13891,N_13784);
nand U14470 (N_14470,N_13864,N_13877);
and U14471 (N_14471,N_14206,N_14391);
nor U14472 (N_14472,N_13743,N_13990);
or U14473 (N_14473,N_13814,N_14199);
or U14474 (N_14474,N_14148,N_13904);
nand U14475 (N_14475,N_13876,N_14034);
nor U14476 (N_14476,N_14216,N_14336);
nand U14477 (N_14477,N_13663,N_13810);
nand U14478 (N_14478,N_14085,N_14115);
nor U14479 (N_14479,N_14038,N_14003);
xor U14480 (N_14480,N_14166,N_13884);
or U14481 (N_14481,N_14273,N_14242);
and U14482 (N_14482,N_13645,N_13988);
or U14483 (N_14483,N_14104,N_13727);
and U14484 (N_14484,N_14077,N_13627);
nand U14485 (N_14485,N_13604,N_14390);
xnor U14486 (N_14486,N_13844,N_13808);
or U14487 (N_14487,N_14138,N_14237);
nor U14488 (N_14488,N_13831,N_13782);
xor U14489 (N_14489,N_14394,N_14234);
and U14490 (N_14490,N_14342,N_14349);
nand U14491 (N_14491,N_13707,N_14083);
and U14492 (N_14492,N_13958,N_13641);
nor U14493 (N_14493,N_14249,N_13712);
xnor U14494 (N_14494,N_13977,N_14395);
nor U14495 (N_14495,N_14022,N_13935);
or U14496 (N_14496,N_14091,N_13772);
nand U14497 (N_14497,N_14292,N_14346);
xor U14498 (N_14498,N_14178,N_13981);
xnor U14499 (N_14499,N_14248,N_14020);
xnor U14500 (N_14500,N_13854,N_14181);
nand U14501 (N_14501,N_13925,N_13976);
nand U14502 (N_14502,N_14168,N_14392);
or U14503 (N_14503,N_13613,N_13656);
xor U14504 (N_14504,N_13757,N_13620);
xor U14505 (N_14505,N_14190,N_14366);
nor U14506 (N_14506,N_13652,N_13890);
nand U14507 (N_14507,N_13820,N_14123);
nor U14508 (N_14508,N_13842,N_13883);
nor U14509 (N_14509,N_13736,N_13899);
and U14510 (N_14510,N_14358,N_14050);
and U14511 (N_14511,N_14301,N_14265);
nand U14512 (N_14512,N_13862,N_13792);
nor U14513 (N_14513,N_13839,N_13887);
nand U14514 (N_14514,N_13848,N_14309);
and U14515 (N_14515,N_14119,N_13775);
or U14516 (N_14516,N_14130,N_14182);
and U14517 (N_14517,N_14361,N_13894);
xor U14518 (N_14518,N_14049,N_13860);
nor U14519 (N_14519,N_14158,N_13835);
xor U14520 (N_14520,N_13766,N_13975);
nand U14521 (N_14521,N_14159,N_14153);
and U14522 (N_14522,N_14313,N_13913);
nand U14523 (N_14523,N_13986,N_14354);
xor U14524 (N_14524,N_13946,N_13952);
nor U14525 (N_14525,N_13821,N_13909);
nand U14526 (N_14526,N_13688,N_14039);
or U14527 (N_14527,N_14239,N_14315);
nor U14528 (N_14528,N_14064,N_13722);
xor U14529 (N_14529,N_14335,N_14105);
nand U14530 (N_14530,N_13741,N_14371);
and U14531 (N_14531,N_13610,N_13916);
or U14532 (N_14532,N_13742,N_13607);
xor U14533 (N_14533,N_14137,N_13763);
nand U14534 (N_14534,N_13721,N_13797);
nand U14535 (N_14535,N_13915,N_13974);
nand U14536 (N_14536,N_14089,N_13755);
nand U14537 (N_14537,N_13694,N_14078);
nand U14538 (N_14538,N_13853,N_13931);
nand U14539 (N_14539,N_13666,N_14167);
xor U14540 (N_14540,N_14250,N_14251);
or U14541 (N_14541,N_13758,N_14120);
and U14542 (N_14542,N_14382,N_14061);
nor U14543 (N_14543,N_13903,N_14364);
and U14544 (N_14544,N_14100,N_14056);
nor U14545 (N_14545,N_14154,N_13675);
xor U14546 (N_14546,N_13970,N_14132);
and U14547 (N_14547,N_14337,N_14068);
or U14548 (N_14548,N_13834,N_14377);
nand U14549 (N_14549,N_13646,N_13658);
nand U14550 (N_14550,N_13926,N_14398);
and U14551 (N_14551,N_14149,N_14160);
nand U14552 (N_14552,N_14072,N_14362);
and U14553 (N_14553,N_14211,N_13880);
nand U14554 (N_14554,N_14006,N_14121);
nand U14555 (N_14555,N_14036,N_14270);
and U14556 (N_14556,N_14333,N_14118);
and U14557 (N_14557,N_13732,N_13954);
or U14558 (N_14558,N_13685,N_13964);
and U14559 (N_14559,N_13737,N_13671);
or U14560 (N_14560,N_14145,N_14261);
xnor U14561 (N_14561,N_13980,N_14323);
xor U14562 (N_14562,N_13996,N_13779);
and U14563 (N_14563,N_13643,N_13709);
nand U14564 (N_14564,N_13642,N_14071);
and U14565 (N_14565,N_13781,N_13672);
nand U14566 (N_14566,N_13923,N_14330);
nor U14567 (N_14567,N_13614,N_13774);
nand U14568 (N_14568,N_14197,N_13805);
xnor U14569 (N_14569,N_14241,N_13944);
and U14570 (N_14570,N_14175,N_13852);
or U14571 (N_14571,N_13752,N_13789);
nor U14572 (N_14572,N_14031,N_13858);
nor U14573 (N_14573,N_14266,N_14238);
nand U14574 (N_14574,N_13668,N_13959);
nand U14575 (N_14575,N_13843,N_14300);
or U14576 (N_14576,N_13696,N_13714);
nand U14577 (N_14577,N_14370,N_14345);
and U14578 (N_14578,N_14135,N_13670);
nor U14579 (N_14579,N_14033,N_13832);
xor U14580 (N_14580,N_13632,N_14052);
nor U14581 (N_14581,N_14219,N_13673);
nand U14582 (N_14582,N_14230,N_14128);
or U14583 (N_14583,N_14314,N_13690);
nor U14584 (N_14584,N_13968,N_14174);
or U14585 (N_14585,N_13987,N_13623);
or U14586 (N_14586,N_14097,N_14284);
nand U14587 (N_14587,N_13788,N_13902);
nand U14588 (N_14588,N_13807,N_14257);
or U14589 (N_14589,N_13651,N_14025);
nor U14590 (N_14590,N_13622,N_13708);
nand U14591 (N_14591,N_14140,N_14143);
xor U14592 (N_14592,N_13662,N_13813);
nand U14593 (N_14593,N_13921,N_14000);
nor U14594 (N_14594,N_14037,N_13669);
and U14595 (N_14595,N_14235,N_14027);
or U14596 (N_14596,N_14312,N_13724);
and U14597 (N_14597,N_13750,N_14247);
nor U14598 (N_14598,N_14277,N_13676);
nand U14599 (N_14599,N_14075,N_14169);
or U14600 (N_14600,N_13861,N_14090);
nand U14601 (N_14601,N_13697,N_13749);
xnor U14602 (N_14602,N_14217,N_14194);
nand U14603 (N_14603,N_14021,N_13901);
nor U14604 (N_14604,N_13719,N_14139);
or U14605 (N_14605,N_14355,N_14227);
nand U14606 (N_14606,N_13800,N_14307);
xnor U14607 (N_14607,N_14267,N_13992);
xor U14608 (N_14608,N_14287,N_13885);
nor U14609 (N_14609,N_13605,N_14032);
nor U14610 (N_14610,N_13634,N_13636);
and U14611 (N_14611,N_13870,N_13818);
and U14612 (N_14612,N_14351,N_13626);
nor U14613 (N_14613,N_13738,N_14019);
or U14614 (N_14614,N_14074,N_13660);
nor U14615 (N_14615,N_14373,N_14142);
nor U14616 (N_14616,N_14385,N_13806);
xor U14617 (N_14617,N_14369,N_13790);
nor U14618 (N_14618,N_13827,N_13771);
and U14619 (N_14619,N_14384,N_14232);
nand U14620 (N_14620,N_13838,N_13764);
or U14621 (N_14621,N_14374,N_14042);
xnor U14622 (N_14622,N_14045,N_13841);
or U14623 (N_14623,N_13637,N_13942);
or U14624 (N_14624,N_13941,N_13616);
and U14625 (N_14625,N_14209,N_14372);
xnor U14626 (N_14626,N_14381,N_13956);
and U14627 (N_14627,N_13633,N_13615);
or U14628 (N_14628,N_14012,N_14018);
or U14629 (N_14629,N_14009,N_13879);
and U14630 (N_14630,N_14306,N_14096);
xor U14631 (N_14631,N_14136,N_14192);
nand U14632 (N_14632,N_14201,N_14082);
or U14633 (N_14633,N_13939,N_14183);
nor U14634 (N_14634,N_13756,N_14344);
or U14635 (N_14635,N_14144,N_14332);
xor U14636 (N_14636,N_14397,N_14236);
xnor U14637 (N_14637,N_14010,N_14116);
xor U14638 (N_14638,N_14011,N_14103);
nand U14639 (N_14639,N_13705,N_13949);
or U14640 (N_14640,N_14260,N_13648);
and U14641 (N_14641,N_13654,N_14095);
xor U14642 (N_14642,N_14305,N_14311);
xor U14643 (N_14643,N_13938,N_13635);
and U14644 (N_14644,N_14328,N_13934);
and U14645 (N_14645,N_13600,N_14399);
nand U14646 (N_14646,N_13888,N_13691);
nor U14647 (N_14647,N_14079,N_14080);
xnor U14648 (N_14648,N_13794,N_14141);
nor U14649 (N_14649,N_14225,N_14376);
nand U14650 (N_14650,N_14255,N_14275);
and U14651 (N_14651,N_13911,N_14196);
nand U14652 (N_14652,N_13687,N_13739);
or U14653 (N_14653,N_14316,N_14014);
xnor U14654 (N_14654,N_13609,N_13754);
and U14655 (N_14655,N_13953,N_13994);
nor U14656 (N_14656,N_13961,N_14004);
and U14657 (N_14657,N_14088,N_13799);
or U14658 (N_14658,N_13816,N_14150);
nand U14659 (N_14659,N_13867,N_13630);
or U14660 (N_14660,N_13945,N_13865);
and U14661 (N_14661,N_13824,N_14319);
nor U14662 (N_14662,N_14298,N_14113);
and U14663 (N_14663,N_13826,N_14172);
nor U14664 (N_14664,N_13686,N_13914);
nor U14665 (N_14665,N_13785,N_13704);
and U14666 (N_14666,N_14069,N_13872);
nor U14667 (N_14667,N_13955,N_14151);
or U14668 (N_14668,N_13647,N_13787);
nor U14669 (N_14669,N_14155,N_14327);
nor U14670 (N_14670,N_13868,N_13893);
or U14671 (N_14671,N_13889,N_14302);
and U14672 (N_14672,N_13699,N_14099);
nand U14673 (N_14673,N_14263,N_13698);
nor U14674 (N_14674,N_14363,N_14367);
xnor U14675 (N_14675,N_14303,N_13619);
and U14676 (N_14676,N_14176,N_14338);
or U14677 (N_14677,N_13943,N_14106);
and U14678 (N_14678,N_13963,N_14131);
nor U14679 (N_14679,N_13659,N_13837);
or U14680 (N_14680,N_13940,N_14203);
and U14681 (N_14681,N_13695,N_13957);
nor U14682 (N_14682,N_13917,N_13649);
xnor U14683 (N_14683,N_14353,N_13830);
nor U14684 (N_14684,N_14339,N_13851);
xnor U14685 (N_14685,N_13984,N_13798);
nand U14686 (N_14686,N_14202,N_13973);
and U14687 (N_14687,N_13989,N_13723);
and U14688 (N_14688,N_13919,N_13728);
nor U14689 (N_14689,N_14308,N_13983);
xor U14690 (N_14690,N_13770,N_13629);
and U14691 (N_14691,N_13729,N_13857);
nand U14692 (N_14692,N_14073,N_14017);
nand U14693 (N_14693,N_13896,N_14218);
or U14694 (N_14694,N_13765,N_14243);
nand U14695 (N_14695,N_13929,N_13971);
xor U14696 (N_14696,N_13730,N_14210);
and U14697 (N_14697,N_13655,N_14272);
or U14698 (N_14698,N_14191,N_14040);
and U14699 (N_14699,N_14389,N_13828);
nor U14700 (N_14700,N_14350,N_13840);
or U14701 (N_14701,N_14246,N_14317);
and U14702 (N_14702,N_14396,N_13869);
nor U14703 (N_14703,N_13625,N_13948);
xnor U14704 (N_14704,N_13640,N_14008);
nor U14705 (N_14705,N_13875,N_14086);
or U14706 (N_14706,N_13985,N_14156);
xnor U14707 (N_14707,N_14386,N_14058);
and U14708 (N_14708,N_14204,N_13720);
or U14709 (N_14709,N_13682,N_14359);
xor U14710 (N_14710,N_13845,N_13793);
xnor U14711 (N_14711,N_14129,N_13928);
or U14712 (N_14712,N_13783,N_13679);
or U14713 (N_14713,N_13628,N_14343);
or U14714 (N_14714,N_13922,N_13998);
and U14715 (N_14715,N_13907,N_14286);
nor U14716 (N_14716,N_13900,N_14112);
and U14717 (N_14717,N_14279,N_13859);
nand U14718 (N_14718,N_14028,N_13684);
nand U14719 (N_14719,N_14274,N_13978);
xor U14720 (N_14720,N_13802,N_14233);
nor U14721 (N_14721,N_13725,N_14187);
nand U14722 (N_14722,N_14281,N_14016);
or U14723 (N_14723,N_13680,N_14262);
nand U14724 (N_14724,N_13905,N_14107);
or U14725 (N_14725,N_14387,N_13693);
nor U14726 (N_14726,N_14126,N_14318);
xnor U14727 (N_14727,N_14109,N_13602);
or U14728 (N_14728,N_13829,N_14189);
nor U14729 (N_14729,N_14084,N_14127);
nor U14730 (N_14730,N_13621,N_14268);
nand U14731 (N_14731,N_14259,N_14205);
nor U14732 (N_14732,N_14388,N_13608);
nor U14733 (N_14733,N_14331,N_13932);
and U14734 (N_14734,N_14297,N_13603);
and U14735 (N_14735,N_13703,N_14152);
nor U14736 (N_14736,N_14098,N_14291);
and U14737 (N_14737,N_13796,N_14245);
or U14738 (N_14738,N_13624,N_13897);
xnor U14739 (N_14739,N_13947,N_14252);
and U14740 (N_14740,N_13910,N_14024);
and U14741 (N_14741,N_14048,N_14117);
nand U14742 (N_14742,N_14244,N_13638);
xnor U14743 (N_14743,N_14093,N_13881);
xor U14744 (N_14744,N_13795,N_13650);
nand U14745 (N_14745,N_14188,N_13745);
and U14746 (N_14746,N_13731,N_13811);
and U14747 (N_14747,N_14046,N_13825);
nor U14748 (N_14748,N_13850,N_13803);
xor U14749 (N_14749,N_13701,N_13937);
and U14750 (N_14750,N_14161,N_14043);
xor U14751 (N_14751,N_14320,N_13718);
and U14752 (N_14752,N_14066,N_14304);
or U14753 (N_14753,N_13962,N_13950);
nand U14754 (N_14754,N_13965,N_13812);
nor U14755 (N_14755,N_14165,N_14005);
or U14756 (N_14756,N_14310,N_13898);
xor U14757 (N_14757,N_14125,N_14101);
nor U14758 (N_14758,N_13960,N_13734);
nor U14759 (N_14759,N_13618,N_13761);
xor U14760 (N_14760,N_13823,N_14124);
or U14761 (N_14761,N_14173,N_13863);
nor U14762 (N_14762,N_14212,N_14198);
nor U14763 (N_14763,N_13847,N_13710);
nor U14764 (N_14764,N_14133,N_14146);
xor U14765 (N_14765,N_14220,N_14295);
or U14766 (N_14766,N_14380,N_14375);
or U14767 (N_14767,N_14062,N_14030);
or U14768 (N_14768,N_13993,N_13773);
nand U14769 (N_14769,N_13706,N_14162);
nor U14770 (N_14770,N_13972,N_13711);
and U14771 (N_14771,N_13644,N_14360);
or U14772 (N_14772,N_13748,N_13866);
xor U14773 (N_14773,N_14280,N_13924);
xnor U14774 (N_14774,N_13631,N_14222);
xor U14775 (N_14775,N_14164,N_14341);
nor U14776 (N_14776,N_13733,N_14282);
or U14777 (N_14777,N_14157,N_14147);
or U14778 (N_14778,N_13966,N_13874);
and U14779 (N_14779,N_13912,N_14001);
and U14780 (N_14780,N_14283,N_14177);
nor U14781 (N_14781,N_14229,N_13855);
xor U14782 (N_14782,N_14029,N_13777);
and U14783 (N_14783,N_13716,N_13746);
xor U14784 (N_14784,N_13760,N_14208);
or U14785 (N_14785,N_14047,N_14184);
nand U14786 (N_14786,N_14060,N_13653);
nand U14787 (N_14787,N_13664,N_14134);
nand U14788 (N_14788,N_14393,N_14213);
and U14789 (N_14789,N_14357,N_14186);
nand U14790 (N_14790,N_14348,N_14340);
nor U14791 (N_14791,N_13791,N_13819);
and U14792 (N_14792,N_14044,N_13606);
nand U14793 (N_14793,N_13661,N_13751);
xor U14794 (N_14794,N_13906,N_13717);
xnor U14795 (N_14795,N_14293,N_14356);
and U14796 (N_14796,N_14347,N_14057);
nand U14797 (N_14797,N_14254,N_14324);
xor U14798 (N_14798,N_14278,N_13667);
nand U14799 (N_14799,N_14378,N_13702);
and U14800 (N_14800,N_13929,N_13860);
or U14801 (N_14801,N_14327,N_13925);
nor U14802 (N_14802,N_14253,N_13754);
and U14803 (N_14803,N_14313,N_13724);
xor U14804 (N_14804,N_13732,N_14179);
nand U14805 (N_14805,N_14322,N_14036);
nor U14806 (N_14806,N_13895,N_13784);
nor U14807 (N_14807,N_14287,N_14179);
and U14808 (N_14808,N_14106,N_13764);
nor U14809 (N_14809,N_14383,N_13608);
or U14810 (N_14810,N_14341,N_14159);
and U14811 (N_14811,N_13643,N_14355);
nand U14812 (N_14812,N_14307,N_14365);
or U14813 (N_14813,N_13841,N_13777);
or U14814 (N_14814,N_14389,N_14239);
xor U14815 (N_14815,N_13717,N_13757);
nor U14816 (N_14816,N_13626,N_13815);
and U14817 (N_14817,N_13661,N_13987);
xnor U14818 (N_14818,N_14329,N_13644);
and U14819 (N_14819,N_13612,N_14227);
or U14820 (N_14820,N_14355,N_13989);
xor U14821 (N_14821,N_13651,N_14077);
or U14822 (N_14822,N_13726,N_14017);
and U14823 (N_14823,N_13896,N_13889);
nand U14824 (N_14824,N_13717,N_13648);
or U14825 (N_14825,N_13820,N_13770);
nand U14826 (N_14826,N_13642,N_14353);
or U14827 (N_14827,N_13602,N_14141);
and U14828 (N_14828,N_13681,N_14361);
xnor U14829 (N_14829,N_14073,N_13872);
nand U14830 (N_14830,N_13630,N_13794);
nand U14831 (N_14831,N_13732,N_13718);
xor U14832 (N_14832,N_13616,N_14391);
and U14833 (N_14833,N_13870,N_13940);
and U14834 (N_14834,N_13727,N_13935);
nor U14835 (N_14835,N_13723,N_13649);
xnor U14836 (N_14836,N_14287,N_13929);
or U14837 (N_14837,N_14199,N_14062);
nand U14838 (N_14838,N_14078,N_13677);
and U14839 (N_14839,N_13739,N_13928);
and U14840 (N_14840,N_13783,N_13846);
nor U14841 (N_14841,N_13937,N_14082);
or U14842 (N_14842,N_13702,N_13704);
or U14843 (N_14843,N_14130,N_13983);
xor U14844 (N_14844,N_14368,N_14119);
or U14845 (N_14845,N_14095,N_14160);
xnor U14846 (N_14846,N_14276,N_13710);
nand U14847 (N_14847,N_14059,N_14273);
xor U14848 (N_14848,N_13842,N_14225);
and U14849 (N_14849,N_13654,N_13950);
xnor U14850 (N_14850,N_14248,N_14018);
nand U14851 (N_14851,N_13975,N_13778);
and U14852 (N_14852,N_14167,N_14233);
nand U14853 (N_14853,N_13747,N_13990);
xor U14854 (N_14854,N_14121,N_13851);
nand U14855 (N_14855,N_14136,N_13864);
nor U14856 (N_14856,N_14012,N_14370);
nand U14857 (N_14857,N_14354,N_14037);
nand U14858 (N_14858,N_14304,N_13928);
xor U14859 (N_14859,N_14002,N_14232);
nand U14860 (N_14860,N_14204,N_14095);
and U14861 (N_14861,N_13624,N_13934);
and U14862 (N_14862,N_14169,N_14217);
nor U14863 (N_14863,N_13896,N_13719);
xor U14864 (N_14864,N_13826,N_13935);
and U14865 (N_14865,N_13942,N_13870);
xnor U14866 (N_14866,N_13768,N_13908);
xor U14867 (N_14867,N_13796,N_14281);
or U14868 (N_14868,N_14340,N_13961);
xor U14869 (N_14869,N_13781,N_14064);
and U14870 (N_14870,N_13656,N_13899);
nor U14871 (N_14871,N_14069,N_14284);
or U14872 (N_14872,N_13777,N_13988);
and U14873 (N_14873,N_13704,N_14334);
and U14874 (N_14874,N_14165,N_14293);
nand U14875 (N_14875,N_14063,N_14284);
nand U14876 (N_14876,N_13705,N_13689);
nand U14877 (N_14877,N_14141,N_13771);
and U14878 (N_14878,N_13716,N_13672);
nand U14879 (N_14879,N_14349,N_14047);
xnor U14880 (N_14880,N_14398,N_13998);
nor U14881 (N_14881,N_13910,N_14339);
and U14882 (N_14882,N_13716,N_14045);
xnor U14883 (N_14883,N_13722,N_14156);
and U14884 (N_14884,N_13839,N_13714);
or U14885 (N_14885,N_13767,N_13601);
and U14886 (N_14886,N_13651,N_14068);
and U14887 (N_14887,N_13795,N_14008);
nor U14888 (N_14888,N_14304,N_14358);
xnor U14889 (N_14889,N_14344,N_14364);
nor U14890 (N_14890,N_14111,N_13772);
xor U14891 (N_14891,N_14310,N_14212);
or U14892 (N_14892,N_14193,N_14239);
xor U14893 (N_14893,N_14006,N_14337);
nand U14894 (N_14894,N_13812,N_14210);
nand U14895 (N_14895,N_14017,N_14066);
and U14896 (N_14896,N_14185,N_14247);
or U14897 (N_14897,N_13642,N_13802);
nand U14898 (N_14898,N_13634,N_13608);
or U14899 (N_14899,N_13729,N_13644);
or U14900 (N_14900,N_13673,N_13662);
or U14901 (N_14901,N_13691,N_13810);
xnor U14902 (N_14902,N_13915,N_13687);
and U14903 (N_14903,N_14053,N_13895);
and U14904 (N_14904,N_14286,N_14026);
nor U14905 (N_14905,N_13787,N_14335);
xor U14906 (N_14906,N_14133,N_14078);
and U14907 (N_14907,N_14096,N_13909);
or U14908 (N_14908,N_13768,N_14121);
nand U14909 (N_14909,N_13912,N_14118);
nand U14910 (N_14910,N_13925,N_14187);
nor U14911 (N_14911,N_13700,N_14319);
nand U14912 (N_14912,N_13904,N_13919);
and U14913 (N_14913,N_14247,N_13855);
nand U14914 (N_14914,N_14129,N_13611);
xor U14915 (N_14915,N_13752,N_14120);
xor U14916 (N_14916,N_14016,N_13994);
xor U14917 (N_14917,N_13740,N_13764);
xor U14918 (N_14918,N_13875,N_14083);
xor U14919 (N_14919,N_14230,N_13693);
xnor U14920 (N_14920,N_13810,N_14176);
nor U14921 (N_14921,N_14168,N_13845);
nor U14922 (N_14922,N_13692,N_13630);
nor U14923 (N_14923,N_13870,N_13832);
xnor U14924 (N_14924,N_13976,N_14049);
nand U14925 (N_14925,N_13923,N_13874);
nor U14926 (N_14926,N_13628,N_13836);
nor U14927 (N_14927,N_13832,N_14226);
and U14928 (N_14928,N_13734,N_13751);
and U14929 (N_14929,N_14139,N_13600);
nand U14930 (N_14930,N_13683,N_13863);
and U14931 (N_14931,N_14176,N_13695);
nor U14932 (N_14932,N_14011,N_13872);
nand U14933 (N_14933,N_13973,N_14072);
nor U14934 (N_14934,N_13744,N_14208);
xor U14935 (N_14935,N_14084,N_13828);
and U14936 (N_14936,N_14313,N_14231);
or U14937 (N_14937,N_14096,N_14386);
nor U14938 (N_14938,N_14132,N_14153);
or U14939 (N_14939,N_13902,N_14199);
nand U14940 (N_14940,N_14385,N_13793);
xnor U14941 (N_14941,N_14006,N_13659);
xnor U14942 (N_14942,N_13967,N_13884);
xnor U14943 (N_14943,N_14191,N_14223);
or U14944 (N_14944,N_14024,N_13823);
nor U14945 (N_14945,N_13750,N_13607);
and U14946 (N_14946,N_13926,N_13876);
nor U14947 (N_14947,N_13778,N_14387);
nor U14948 (N_14948,N_14189,N_13665);
or U14949 (N_14949,N_14208,N_14390);
nor U14950 (N_14950,N_13748,N_14391);
xor U14951 (N_14951,N_13812,N_13961);
nand U14952 (N_14952,N_14380,N_13957);
nand U14953 (N_14953,N_14289,N_13696);
nand U14954 (N_14954,N_14138,N_14329);
xor U14955 (N_14955,N_13626,N_14181);
xnor U14956 (N_14956,N_14213,N_13875);
nor U14957 (N_14957,N_14265,N_14040);
nor U14958 (N_14958,N_14243,N_13639);
xor U14959 (N_14959,N_14179,N_13811);
or U14960 (N_14960,N_13814,N_14104);
nor U14961 (N_14961,N_14376,N_14109);
nand U14962 (N_14962,N_13979,N_14162);
and U14963 (N_14963,N_13830,N_14169);
nor U14964 (N_14964,N_13943,N_14309);
nand U14965 (N_14965,N_14130,N_13949);
xnor U14966 (N_14966,N_13694,N_14029);
or U14967 (N_14967,N_14234,N_13921);
and U14968 (N_14968,N_13839,N_13840);
xor U14969 (N_14969,N_13752,N_14048);
xnor U14970 (N_14970,N_13897,N_13741);
and U14971 (N_14971,N_14281,N_13735);
nor U14972 (N_14972,N_14255,N_13768);
and U14973 (N_14973,N_13967,N_14109);
xor U14974 (N_14974,N_13677,N_14346);
nor U14975 (N_14975,N_14029,N_14221);
and U14976 (N_14976,N_14194,N_14363);
nand U14977 (N_14977,N_14163,N_14174);
nand U14978 (N_14978,N_14105,N_13899);
xor U14979 (N_14979,N_14235,N_13922);
or U14980 (N_14980,N_14321,N_14381);
or U14981 (N_14981,N_14266,N_13685);
xnor U14982 (N_14982,N_13664,N_13773);
nand U14983 (N_14983,N_14108,N_13882);
xor U14984 (N_14984,N_14288,N_13649);
and U14985 (N_14985,N_14107,N_14363);
xnor U14986 (N_14986,N_13661,N_13726);
nand U14987 (N_14987,N_14048,N_13741);
or U14988 (N_14988,N_13911,N_14072);
nor U14989 (N_14989,N_14055,N_14026);
and U14990 (N_14990,N_14313,N_14308);
xor U14991 (N_14991,N_13848,N_14011);
and U14992 (N_14992,N_13611,N_13988);
nor U14993 (N_14993,N_13743,N_14250);
nor U14994 (N_14994,N_14133,N_13714);
nand U14995 (N_14995,N_13674,N_13789);
and U14996 (N_14996,N_13911,N_14283);
xor U14997 (N_14997,N_14206,N_14147);
nand U14998 (N_14998,N_13936,N_14040);
and U14999 (N_14999,N_14337,N_13671);
nor U15000 (N_15000,N_14006,N_14270);
and U15001 (N_15001,N_13669,N_14258);
nor U15002 (N_15002,N_14266,N_14050);
nor U15003 (N_15003,N_13891,N_14300);
or U15004 (N_15004,N_14297,N_14392);
and U15005 (N_15005,N_13952,N_13901);
nor U15006 (N_15006,N_13965,N_14338);
and U15007 (N_15007,N_13813,N_14379);
xor U15008 (N_15008,N_14040,N_14207);
xnor U15009 (N_15009,N_13655,N_14332);
and U15010 (N_15010,N_14332,N_14232);
or U15011 (N_15011,N_14101,N_13840);
nor U15012 (N_15012,N_13651,N_13607);
and U15013 (N_15013,N_13817,N_14323);
or U15014 (N_15014,N_13734,N_13890);
nor U15015 (N_15015,N_14076,N_13909);
and U15016 (N_15016,N_14351,N_13854);
or U15017 (N_15017,N_13801,N_13819);
or U15018 (N_15018,N_13748,N_14172);
or U15019 (N_15019,N_14099,N_13978);
xnor U15020 (N_15020,N_13625,N_13777);
xor U15021 (N_15021,N_13922,N_14349);
or U15022 (N_15022,N_14193,N_13661);
and U15023 (N_15023,N_14021,N_13905);
nor U15024 (N_15024,N_14059,N_14025);
nand U15025 (N_15025,N_13685,N_13985);
nor U15026 (N_15026,N_13688,N_13649);
or U15027 (N_15027,N_13954,N_13679);
xor U15028 (N_15028,N_13674,N_13631);
xor U15029 (N_15029,N_13996,N_14204);
nor U15030 (N_15030,N_14114,N_13768);
and U15031 (N_15031,N_14045,N_14308);
nor U15032 (N_15032,N_13886,N_14239);
nand U15033 (N_15033,N_14128,N_13611);
and U15034 (N_15034,N_14392,N_13799);
nor U15035 (N_15035,N_14115,N_14065);
xor U15036 (N_15036,N_13735,N_13619);
nand U15037 (N_15037,N_13674,N_14227);
and U15038 (N_15038,N_13868,N_14248);
nor U15039 (N_15039,N_13929,N_14361);
and U15040 (N_15040,N_14240,N_14151);
nand U15041 (N_15041,N_13979,N_14314);
and U15042 (N_15042,N_14389,N_13666);
or U15043 (N_15043,N_14154,N_13608);
nor U15044 (N_15044,N_13780,N_14357);
xnor U15045 (N_15045,N_13825,N_14199);
nand U15046 (N_15046,N_13840,N_14269);
and U15047 (N_15047,N_14395,N_13816);
or U15048 (N_15048,N_13853,N_13666);
and U15049 (N_15049,N_13670,N_13830);
and U15050 (N_15050,N_14222,N_13728);
nor U15051 (N_15051,N_13600,N_14122);
xor U15052 (N_15052,N_14027,N_13943);
nand U15053 (N_15053,N_13744,N_13953);
nand U15054 (N_15054,N_13777,N_14195);
nand U15055 (N_15055,N_14312,N_14150);
xor U15056 (N_15056,N_13700,N_13912);
or U15057 (N_15057,N_13641,N_13687);
and U15058 (N_15058,N_13637,N_14370);
nor U15059 (N_15059,N_13659,N_13815);
and U15060 (N_15060,N_13746,N_13784);
and U15061 (N_15061,N_14374,N_13650);
nand U15062 (N_15062,N_13631,N_14082);
or U15063 (N_15063,N_14220,N_13696);
and U15064 (N_15064,N_13908,N_13866);
or U15065 (N_15065,N_13854,N_14255);
nor U15066 (N_15066,N_14293,N_14030);
nand U15067 (N_15067,N_13677,N_14399);
or U15068 (N_15068,N_14146,N_14280);
xnor U15069 (N_15069,N_14240,N_14313);
nor U15070 (N_15070,N_13775,N_13717);
or U15071 (N_15071,N_14056,N_13938);
nor U15072 (N_15072,N_13779,N_14005);
nand U15073 (N_15073,N_14040,N_13826);
nor U15074 (N_15074,N_13826,N_13925);
and U15075 (N_15075,N_14059,N_14183);
nand U15076 (N_15076,N_13748,N_13969);
and U15077 (N_15077,N_13601,N_14379);
nand U15078 (N_15078,N_14170,N_13822);
or U15079 (N_15079,N_14382,N_13950);
nor U15080 (N_15080,N_13914,N_13722);
xor U15081 (N_15081,N_14004,N_13723);
xor U15082 (N_15082,N_14044,N_14160);
and U15083 (N_15083,N_13965,N_13916);
nand U15084 (N_15084,N_14373,N_13661);
and U15085 (N_15085,N_13677,N_13870);
nand U15086 (N_15086,N_13833,N_14017);
nand U15087 (N_15087,N_14042,N_13619);
nand U15088 (N_15088,N_14153,N_14316);
nor U15089 (N_15089,N_13953,N_13977);
and U15090 (N_15090,N_13824,N_13759);
nor U15091 (N_15091,N_13638,N_13925);
nor U15092 (N_15092,N_14318,N_13861);
or U15093 (N_15093,N_13606,N_14055);
nand U15094 (N_15094,N_13909,N_13772);
nor U15095 (N_15095,N_13792,N_13807);
or U15096 (N_15096,N_14092,N_14168);
nor U15097 (N_15097,N_14387,N_13934);
nor U15098 (N_15098,N_13764,N_13634);
and U15099 (N_15099,N_14282,N_14364);
xnor U15100 (N_15100,N_14218,N_13919);
and U15101 (N_15101,N_13767,N_14064);
nand U15102 (N_15102,N_13862,N_14114);
xor U15103 (N_15103,N_13969,N_14339);
nor U15104 (N_15104,N_13933,N_13896);
nand U15105 (N_15105,N_13854,N_13888);
nor U15106 (N_15106,N_13756,N_13984);
xnor U15107 (N_15107,N_14230,N_13767);
or U15108 (N_15108,N_14041,N_14032);
or U15109 (N_15109,N_13857,N_13685);
xor U15110 (N_15110,N_13927,N_13918);
xnor U15111 (N_15111,N_13820,N_14328);
xor U15112 (N_15112,N_13875,N_13904);
nor U15113 (N_15113,N_14000,N_13695);
and U15114 (N_15114,N_13647,N_14074);
nor U15115 (N_15115,N_14003,N_14242);
or U15116 (N_15116,N_14385,N_14336);
nor U15117 (N_15117,N_13697,N_14137);
nand U15118 (N_15118,N_13724,N_13823);
and U15119 (N_15119,N_13999,N_13816);
nand U15120 (N_15120,N_14385,N_14023);
nor U15121 (N_15121,N_13876,N_14165);
and U15122 (N_15122,N_14150,N_14103);
nand U15123 (N_15123,N_14084,N_13621);
and U15124 (N_15124,N_14390,N_14294);
xor U15125 (N_15125,N_14164,N_13648);
and U15126 (N_15126,N_13713,N_13643);
and U15127 (N_15127,N_14032,N_14003);
nor U15128 (N_15128,N_14184,N_14318);
xnor U15129 (N_15129,N_13721,N_14130);
and U15130 (N_15130,N_14287,N_13654);
xnor U15131 (N_15131,N_14347,N_14112);
or U15132 (N_15132,N_13709,N_14262);
xnor U15133 (N_15133,N_13957,N_13913);
or U15134 (N_15134,N_14033,N_14044);
and U15135 (N_15135,N_14306,N_14368);
or U15136 (N_15136,N_14231,N_14394);
and U15137 (N_15137,N_14192,N_14082);
nor U15138 (N_15138,N_14250,N_13635);
or U15139 (N_15139,N_14357,N_13787);
nor U15140 (N_15140,N_13827,N_13854);
nand U15141 (N_15141,N_13965,N_13822);
xnor U15142 (N_15142,N_14226,N_13609);
nor U15143 (N_15143,N_13771,N_14312);
nor U15144 (N_15144,N_13838,N_13979);
nor U15145 (N_15145,N_13915,N_13601);
nor U15146 (N_15146,N_13818,N_14167);
nand U15147 (N_15147,N_14134,N_13685);
or U15148 (N_15148,N_13679,N_14382);
nand U15149 (N_15149,N_13690,N_13983);
nand U15150 (N_15150,N_13824,N_14120);
xnor U15151 (N_15151,N_14282,N_13688);
nand U15152 (N_15152,N_13719,N_14028);
and U15153 (N_15153,N_13922,N_13617);
and U15154 (N_15154,N_14028,N_14053);
or U15155 (N_15155,N_14251,N_13906);
xor U15156 (N_15156,N_13945,N_14082);
or U15157 (N_15157,N_13862,N_13784);
or U15158 (N_15158,N_14050,N_14034);
and U15159 (N_15159,N_14180,N_14223);
and U15160 (N_15160,N_14151,N_14152);
nor U15161 (N_15161,N_13665,N_13980);
nand U15162 (N_15162,N_14165,N_14196);
nand U15163 (N_15163,N_14324,N_14066);
and U15164 (N_15164,N_13899,N_13816);
or U15165 (N_15165,N_14274,N_14151);
nor U15166 (N_15166,N_13934,N_13815);
or U15167 (N_15167,N_13667,N_13640);
nand U15168 (N_15168,N_13949,N_13991);
and U15169 (N_15169,N_14259,N_14301);
or U15170 (N_15170,N_14156,N_13673);
nor U15171 (N_15171,N_14285,N_13831);
nand U15172 (N_15172,N_14252,N_14247);
nand U15173 (N_15173,N_13729,N_14068);
xor U15174 (N_15174,N_13885,N_13906);
xor U15175 (N_15175,N_13648,N_14288);
nand U15176 (N_15176,N_13603,N_13862);
xnor U15177 (N_15177,N_14105,N_13901);
xnor U15178 (N_15178,N_14394,N_13615);
and U15179 (N_15179,N_13950,N_14275);
xor U15180 (N_15180,N_13991,N_14275);
or U15181 (N_15181,N_13790,N_13978);
or U15182 (N_15182,N_13662,N_13604);
nand U15183 (N_15183,N_13791,N_14356);
and U15184 (N_15184,N_14044,N_13692);
xor U15185 (N_15185,N_14050,N_13932);
xor U15186 (N_15186,N_13600,N_14387);
and U15187 (N_15187,N_13659,N_13889);
nor U15188 (N_15188,N_13928,N_13858);
xor U15189 (N_15189,N_14039,N_13769);
or U15190 (N_15190,N_14090,N_13720);
and U15191 (N_15191,N_14343,N_13715);
and U15192 (N_15192,N_13622,N_14002);
and U15193 (N_15193,N_13651,N_14260);
and U15194 (N_15194,N_14328,N_14153);
nor U15195 (N_15195,N_14117,N_14347);
nand U15196 (N_15196,N_13799,N_14059);
and U15197 (N_15197,N_13912,N_13600);
xor U15198 (N_15198,N_14096,N_13841);
or U15199 (N_15199,N_13998,N_14344);
nor U15200 (N_15200,N_14760,N_14447);
nor U15201 (N_15201,N_15000,N_14860);
or U15202 (N_15202,N_15141,N_14530);
or U15203 (N_15203,N_14578,N_15088);
xor U15204 (N_15204,N_14518,N_14745);
and U15205 (N_15205,N_14569,N_14998);
xnor U15206 (N_15206,N_14925,N_14980);
or U15207 (N_15207,N_14579,N_14476);
and U15208 (N_15208,N_14611,N_14836);
or U15209 (N_15209,N_14939,N_14900);
nor U15210 (N_15210,N_14940,N_14794);
or U15211 (N_15211,N_14712,N_14759);
xnor U15212 (N_15212,N_15108,N_14955);
nand U15213 (N_15213,N_14947,N_15144);
nand U15214 (N_15214,N_14960,N_14634);
or U15215 (N_15215,N_14656,N_15169);
nand U15216 (N_15216,N_14461,N_14920);
or U15217 (N_15217,N_14607,N_14624);
xor U15218 (N_15218,N_15162,N_15197);
or U15219 (N_15219,N_15128,N_15111);
xor U15220 (N_15220,N_14978,N_14618);
or U15221 (N_15221,N_14943,N_14545);
and U15222 (N_15222,N_14442,N_14544);
and U15223 (N_15223,N_15164,N_14504);
and U15224 (N_15224,N_15065,N_14708);
and U15225 (N_15225,N_14553,N_14416);
nor U15226 (N_15226,N_14630,N_14730);
nor U15227 (N_15227,N_14912,N_14772);
xnor U15228 (N_15228,N_15199,N_14804);
or U15229 (N_15229,N_14781,N_14986);
and U15230 (N_15230,N_14625,N_14597);
or U15231 (N_15231,N_14401,N_15029);
or U15232 (N_15232,N_14741,N_15053);
nor U15233 (N_15233,N_14765,N_14902);
and U15234 (N_15234,N_14552,N_15193);
xor U15235 (N_15235,N_15043,N_14529);
xnor U15236 (N_15236,N_14633,N_14547);
nand U15237 (N_15237,N_15155,N_14665);
and U15238 (N_15238,N_15004,N_14414);
or U15239 (N_15239,N_14891,N_14973);
or U15240 (N_15240,N_15122,N_15070);
nor U15241 (N_15241,N_15003,N_14642);
or U15242 (N_15242,N_14937,N_15179);
or U15243 (N_15243,N_15194,N_14500);
or U15244 (N_15244,N_14729,N_14424);
or U15245 (N_15245,N_14427,N_14830);
nor U15246 (N_15246,N_14441,N_14647);
or U15247 (N_15247,N_14778,N_14697);
or U15248 (N_15248,N_14813,N_14617);
nor U15249 (N_15249,N_15107,N_14679);
xnor U15250 (N_15250,N_14546,N_14823);
and U15251 (N_15251,N_15061,N_15024);
nand U15252 (N_15252,N_14541,N_15113);
or U15253 (N_15253,N_14910,N_14586);
nand U15254 (N_15254,N_14692,N_15178);
and U15255 (N_15255,N_14975,N_15091);
nor U15256 (N_15256,N_14525,N_14946);
and U15257 (N_15257,N_14568,N_14532);
and U15258 (N_15258,N_15022,N_15160);
or U15259 (N_15259,N_14403,N_15075);
or U15260 (N_15260,N_14822,N_15123);
nand U15261 (N_15261,N_14785,N_14615);
and U15262 (N_15262,N_14793,N_14613);
and U15263 (N_15263,N_14911,N_15104);
and U15264 (N_15264,N_14872,N_14852);
or U15265 (N_15265,N_14649,N_15134);
and U15266 (N_15266,N_14677,N_14695);
nand U15267 (N_15267,N_14931,N_14845);
and U15268 (N_15268,N_14824,N_15039);
and U15269 (N_15269,N_14951,N_15035);
xnor U15270 (N_15270,N_14685,N_14868);
nand U15271 (N_15271,N_15168,N_14450);
and U15272 (N_15272,N_14735,N_14467);
xnor U15273 (N_15273,N_14537,N_14610);
nor U15274 (N_15274,N_14664,N_14731);
or U15275 (N_15275,N_14949,N_14643);
nor U15276 (N_15276,N_14658,N_14832);
and U15277 (N_15277,N_14918,N_14805);
or U15278 (N_15278,N_14746,N_14696);
or U15279 (N_15279,N_14770,N_14524);
nand U15280 (N_15280,N_14654,N_14669);
xnor U15281 (N_15281,N_14711,N_14989);
xnor U15282 (N_15282,N_14933,N_14465);
and U15283 (N_15283,N_15098,N_14879);
nor U15284 (N_15284,N_14536,N_14457);
nor U15285 (N_15285,N_14575,N_14802);
xor U15286 (N_15286,N_14909,N_15090);
or U15287 (N_15287,N_15149,N_14574);
or U15288 (N_15288,N_14971,N_15083);
or U15289 (N_15289,N_14969,N_14990);
xnor U15290 (N_15290,N_15177,N_14659);
nor U15291 (N_15291,N_15192,N_14957);
or U15292 (N_15292,N_15089,N_14854);
and U15293 (N_15293,N_15120,N_14528);
nor U15294 (N_15294,N_14859,N_15095);
nand U15295 (N_15295,N_14761,N_14663);
or U15296 (N_15296,N_14934,N_14959);
and U15297 (N_15297,N_15189,N_14871);
xor U15298 (N_15298,N_14809,N_14815);
nor U15299 (N_15299,N_14515,N_14748);
xnor U15300 (N_15300,N_15012,N_14812);
nor U15301 (N_15301,N_14440,N_14784);
xnor U15302 (N_15302,N_14531,N_14631);
nor U15303 (N_15303,N_14477,N_15064);
xnor U15304 (N_15304,N_14906,N_14619);
or U15305 (N_15305,N_15036,N_15048);
and U15306 (N_15306,N_14533,N_14593);
or U15307 (N_15307,N_14769,N_14870);
nand U15308 (N_15308,N_14865,N_15172);
xor U15309 (N_15309,N_14825,N_15067);
nand U15310 (N_15310,N_14407,N_14707);
or U15311 (N_15311,N_14795,N_15031);
nor U15312 (N_15312,N_15156,N_14437);
and U15313 (N_15313,N_14560,N_14601);
nor U15314 (N_15314,N_14837,N_14462);
and U15315 (N_15315,N_14932,N_14801);
nand U15316 (N_15316,N_14675,N_14688);
nor U15317 (N_15317,N_14542,N_14929);
or U15318 (N_15318,N_14594,N_14783);
nor U15319 (N_15319,N_15105,N_14522);
nand U15320 (N_15320,N_14562,N_14869);
and U15321 (N_15321,N_14520,N_15006);
nor U15322 (N_15322,N_15032,N_15114);
xnor U15323 (N_15323,N_14750,N_14896);
xnor U15324 (N_15324,N_14681,N_14629);
and U15325 (N_15325,N_15151,N_14556);
nand U15326 (N_15326,N_14673,N_14655);
nand U15327 (N_15327,N_15068,N_14724);
xnor U15328 (N_15328,N_15009,N_14779);
nor U15329 (N_15329,N_14502,N_14828);
xor U15330 (N_15330,N_14676,N_14786);
or U15331 (N_15331,N_14953,N_14543);
nand U15332 (N_15332,N_14490,N_15096);
and U15333 (N_15333,N_14637,N_14979);
xnor U15334 (N_15334,N_15126,N_15135);
nor U15335 (N_15335,N_14445,N_14876);
nor U15336 (N_15336,N_15109,N_14456);
nand U15337 (N_15337,N_14576,N_14981);
and U15338 (N_15338,N_14921,N_15087);
and U15339 (N_15339,N_14997,N_15052);
nand U15340 (N_15340,N_14814,N_15145);
or U15341 (N_15341,N_14421,N_15017);
xnor U15342 (N_15342,N_14811,N_15124);
xor U15343 (N_15343,N_15059,N_14999);
nor U15344 (N_15344,N_14604,N_14739);
and U15345 (N_15345,N_14928,N_14402);
or U15346 (N_15346,N_15174,N_14829);
or U15347 (N_15347,N_14598,N_14566);
nand U15348 (N_15348,N_14559,N_14964);
nand U15349 (N_15349,N_14917,N_14736);
xnor U15350 (N_15350,N_14468,N_15045);
xor U15351 (N_15351,N_14965,N_14513);
or U15352 (N_15352,N_14538,N_14833);
and U15353 (N_15353,N_14799,N_14874);
and U15354 (N_15354,N_14762,N_14432);
and U15355 (N_15355,N_14483,N_14700);
nor U15356 (N_15356,N_14493,N_14517);
nor U15357 (N_15357,N_14680,N_15026);
xnor U15358 (N_15358,N_15047,N_15118);
or U15359 (N_15359,N_15099,N_14444);
nand U15360 (N_15360,N_14540,N_14478);
or U15361 (N_15361,N_14961,N_15110);
or U15362 (N_15362,N_15101,N_14671);
nand U15363 (N_15363,N_14751,N_14609);
nor U15364 (N_15364,N_14743,N_14774);
nor U15365 (N_15365,N_14991,N_15137);
or U15366 (N_15366,N_14755,N_14587);
nand U15367 (N_15367,N_14993,N_14603);
nor U15368 (N_15368,N_15018,N_14843);
xor U15369 (N_15369,N_14858,N_14846);
nor U15370 (N_15370,N_14742,N_14678);
nor U15371 (N_15371,N_14409,N_15180);
xnor U15372 (N_15372,N_15069,N_14511);
or U15373 (N_15373,N_15159,N_14800);
xnor U15374 (N_15374,N_15115,N_15082);
nand U15375 (N_15375,N_14771,N_14495);
or U15376 (N_15376,N_14935,N_15196);
xor U15377 (N_15377,N_14738,N_14612);
nand U15378 (N_15378,N_14405,N_14627);
and U15379 (N_15379,N_14820,N_15183);
and U15380 (N_15380,N_14873,N_14577);
and U15381 (N_15381,N_15085,N_15028);
xor U15382 (N_15382,N_14428,N_14430);
nand U15383 (N_15383,N_14919,N_14880);
or U15384 (N_15384,N_14806,N_15157);
nand U15385 (N_15385,N_15187,N_15176);
and U15386 (N_15386,N_15019,N_14429);
xor U15387 (N_15387,N_15100,N_14435);
or U15388 (N_15388,N_14798,N_14704);
xor U15389 (N_15389,N_14535,N_14565);
or U15390 (N_15390,N_14448,N_14719);
or U15391 (N_15391,N_14420,N_14976);
nor U15392 (N_15392,N_14958,N_14411);
or U15393 (N_15393,N_14693,N_14791);
and U15394 (N_15394,N_14599,N_14582);
or U15395 (N_15395,N_14887,N_14952);
and U15396 (N_15396,N_14754,N_14740);
nand U15397 (N_15397,N_14670,N_15080);
xor U15398 (N_15398,N_14585,N_14458);
nor U15399 (N_15399,N_14718,N_14527);
nor U15400 (N_15400,N_14623,N_14727);
and U15401 (N_15401,N_15148,N_14459);
and U15402 (N_15402,N_15044,N_15121);
nand U15403 (N_15403,N_14914,N_15127);
and U15404 (N_15404,N_14423,N_15150);
or U15405 (N_15405,N_15106,N_15076);
xnor U15406 (N_15406,N_14486,N_15094);
nor U15407 (N_15407,N_15060,N_15030);
nand U15408 (N_15408,N_14916,N_15033);
nand U15409 (N_15409,N_14826,N_15190);
nor U15410 (N_15410,N_14714,N_14489);
or U15411 (N_15411,N_15186,N_15092);
or U15412 (N_15412,N_14996,N_14987);
and U15413 (N_15413,N_14581,N_14596);
or U15414 (N_15414,N_14897,N_14972);
xnor U15415 (N_15415,N_14705,N_14526);
nor U15416 (N_15416,N_14454,N_15001);
xnor U15417 (N_15417,N_14494,N_15152);
nand U15418 (N_15418,N_15042,N_14885);
and U15419 (N_15419,N_14963,N_14992);
or U15420 (N_15420,N_15158,N_14737);
and U15421 (N_15421,N_14954,N_14641);
xor U15422 (N_15422,N_14877,N_14867);
nand U15423 (N_15423,N_14410,N_14744);
nor U15424 (N_15424,N_14519,N_14600);
xnor U15425 (N_15425,N_15049,N_15037);
nand U15426 (N_15426,N_14451,N_14471);
or U15427 (N_15427,N_14936,N_14482);
and U15428 (N_15428,N_14775,N_14505);
and U15429 (N_15429,N_15165,N_14516);
or U15430 (N_15430,N_14819,N_14506);
and U15431 (N_15431,N_14817,N_15050);
or U15432 (N_15432,N_14583,N_15055);
or U15433 (N_15433,N_14888,N_15184);
and U15434 (N_15434,N_14474,N_14691);
nor U15435 (N_15435,N_14842,N_14473);
or U15436 (N_15436,N_14966,N_15046);
and U15437 (N_15437,N_14764,N_14408);
or U15438 (N_15438,N_14684,N_14570);
or U15439 (N_15439,N_14835,N_14758);
and U15440 (N_15440,N_14622,N_15013);
or U15441 (N_15441,N_15154,N_15056);
or U15442 (N_15442,N_15102,N_14443);
or U15443 (N_15443,N_14608,N_14807);
xor U15444 (N_15444,N_15066,N_14466);
or U15445 (N_15445,N_14849,N_14595);
nor U15446 (N_15446,N_14415,N_14564);
and U15447 (N_15447,N_15171,N_14709);
or U15448 (N_15448,N_14710,N_14584);
or U15449 (N_15449,N_15079,N_14839);
nand U15450 (N_15450,N_14882,N_14484);
or U15451 (N_15451,N_14682,N_14827);
and U15452 (N_15452,N_14591,N_15027);
nand U15453 (N_15453,N_14901,N_14653);
or U15454 (N_15454,N_14571,N_15136);
and U15455 (N_15455,N_14638,N_14509);
nor U15456 (N_15456,N_14942,N_15011);
and U15457 (N_15457,N_14881,N_14790);
nor U15458 (N_15458,N_14479,N_15072);
nor U15459 (N_15459,N_14988,N_14853);
xor U15460 (N_15460,N_14554,N_14884);
or U15461 (N_15461,N_15182,N_15117);
or U15462 (N_15462,N_15051,N_14722);
and U15463 (N_15463,N_14995,N_14662);
xor U15464 (N_15464,N_14831,N_14944);
nand U15465 (N_15465,N_14922,N_14984);
or U15466 (N_15466,N_14646,N_14683);
nand U15467 (N_15467,N_15074,N_14523);
xor U15468 (N_15468,N_14561,N_14768);
and U15469 (N_15469,N_14469,N_14555);
nand U15470 (N_15470,N_14776,N_14491);
and U15471 (N_15471,N_14892,N_14485);
nor U15472 (N_15472,N_14488,N_14503);
and U15473 (N_15473,N_14548,N_14878);
or U15474 (N_15474,N_14866,N_14487);
and U15475 (N_15475,N_15023,N_15153);
and U15476 (N_15476,N_14945,N_15130);
xnor U15477 (N_15477,N_15167,N_15125);
and U15478 (N_15478,N_14657,N_14481);
nor U15479 (N_15479,N_14893,N_14418);
nor U15480 (N_15480,N_14752,N_14521);
or U15481 (N_15481,N_14507,N_14728);
or U15482 (N_15482,N_15007,N_15057);
nor U15483 (N_15483,N_15142,N_15020);
nand U15484 (N_15484,N_14498,N_14962);
xor U15485 (N_15485,N_14694,N_14419);
or U15486 (N_15486,N_14956,N_14968);
or U15487 (N_15487,N_15040,N_14660);
nand U15488 (N_15488,N_14452,N_14650);
and U15489 (N_15489,N_14661,N_14780);
nor U15490 (N_15490,N_14766,N_14425);
nand U15491 (N_15491,N_14941,N_14938);
or U15492 (N_15492,N_14856,N_14904);
nand U15493 (N_15493,N_14715,N_14550);
and U15494 (N_15494,N_14816,N_14797);
or U15495 (N_15495,N_15112,N_15143);
and U15496 (N_15496,N_14589,N_15041);
and U15497 (N_15497,N_14834,N_14433);
and U15498 (N_15498,N_14557,N_15010);
or U15499 (N_15499,N_15173,N_14756);
nor U15500 (N_15500,N_14651,N_14439);
xor U15501 (N_15501,N_15063,N_14472);
and U15502 (N_15502,N_14453,N_15166);
nand U15503 (N_15503,N_14763,N_14590);
xnor U15504 (N_15504,N_15170,N_14463);
nor U15505 (N_15505,N_14687,N_14499);
nor U15506 (N_15506,N_15185,N_15181);
and U15507 (N_15507,N_15146,N_15016);
nor U15508 (N_15508,N_14767,N_14847);
or U15509 (N_15509,N_14703,N_14644);
and U15510 (N_15510,N_14787,N_15139);
nor U15511 (N_15511,N_14434,N_14850);
xor U15512 (N_15512,N_15097,N_14749);
nor U15513 (N_15513,N_14890,N_14431);
nor U15514 (N_15514,N_14757,N_14926);
or U15515 (N_15515,N_14475,N_14841);
nand U15516 (N_15516,N_14580,N_14863);
or U15517 (N_15517,N_14723,N_14782);
xnor U15518 (N_15518,N_14717,N_14905);
nor U15519 (N_15519,N_14789,N_14422);
nor U15520 (N_15520,N_14514,N_14666);
nand U15521 (N_15521,N_14496,N_15078);
xor U15522 (N_15522,N_14855,N_15021);
and U15523 (N_15523,N_14994,N_15198);
or U15524 (N_15524,N_14848,N_14777);
and U15525 (N_15525,N_14668,N_14400);
and U15526 (N_15526,N_15054,N_14977);
nand U15527 (N_15527,N_14635,N_15015);
xor U15528 (N_15528,N_14626,N_14413);
nor U15529 (N_15529,N_14792,N_14706);
nor U15530 (N_15530,N_14699,N_14567);
nand U15531 (N_15531,N_14861,N_14549);
or U15532 (N_15532,N_14773,N_14930);
nand U15533 (N_15533,N_15025,N_15005);
and U15534 (N_15534,N_14652,N_14983);
nor U15535 (N_15535,N_14788,N_15084);
and U15536 (N_15536,N_14672,N_14674);
nand U15537 (N_15537,N_14701,N_14606);
nand U15538 (N_15538,N_14464,N_15119);
nor U15539 (N_15539,N_14455,N_14702);
nor U15540 (N_15540,N_15071,N_14640);
and U15541 (N_15541,N_14903,N_14539);
nor U15542 (N_15542,N_15002,N_14558);
nor U15543 (N_15543,N_14970,N_14864);
xnor U15544 (N_15544,N_14639,N_15077);
and U15545 (N_15545,N_14851,N_14551);
xnor U15546 (N_15546,N_14886,N_15133);
and U15547 (N_15547,N_14508,N_14497);
and U15548 (N_15548,N_14690,N_15038);
xor U15549 (N_15549,N_14808,N_14720);
nand U15550 (N_15550,N_15161,N_14492);
and U15551 (N_15551,N_14436,N_14698);
nand U15552 (N_15552,N_14747,N_15062);
nor U15553 (N_15553,N_15073,N_14449);
or U15554 (N_15554,N_14632,N_15081);
or U15555 (N_15555,N_14898,N_14894);
nor U15556 (N_15556,N_15116,N_15188);
xor U15557 (N_15557,N_14426,N_15093);
or U15558 (N_15558,N_14862,N_14406);
nor U15559 (N_15559,N_14857,N_14985);
nand U15560 (N_15560,N_14534,N_14726);
xnor U15561 (N_15561,N_14667,N_14573);
or U15562 (N_15562,N_14716,N_15008);
xor U15563 (N_15563,N_14628,N_14721);
or U15564 (N_15564,N_15131,N_15034);
xor U15565 (N_15565,N_14908,N_15129);
nand U15566 (N_15566,N_14796,N_14889);
nand U15567 (N_15567,N_14645,N_14438);
or U15568 (N_15568,N_14927,N_14602);
xnor U15569 (N_15569,N_15058,N_14732);
nand U15570 (N_15570,N_14895,N_14883);
nor U15571 (N_15571,N_14924,N_14733);
nor U15572 (N_15572,N_14913,N_14592);
or U15573 (N_15573,N_14838,N_15132);
nand U15574 (N_15574,N_14713,N_14470);
nor U15575 (N_15575,N_15086,N_14982);
nor U15576 (N_15576,N_14948,N_14844);
or U15577 (N_15577,N_14648,N_14753);
nand U15578 (N_15578,N_14563,N_14907);
nand U15579 (N_15579,N_14572,N_15195);
xnor U15580 (N_15580,N_14803,N_14689);
nand U15581 (N_15581,N_15138,N_14460);
and U15582 (N_15582,N_14512,N_15163);
or U15583 (N_15583,N_14725,N_14501);
nand U15584 (N_15584,N_14950,N_15140);
or U15585 (N_15585,N_14636,N_15191);
nor U15586 (N_15586,N_14967,N_14621);
nand U15587 (N_15587,N_14899,N_14974);
and U15588 (N_15588,N_14821,N_14417);
or U15589 (N_15589,N_14620,N_14588);
and U15590 (N_15590,N_15014,N_14480);
xor U15591 (N_15591,N_14446,N_14605);
xor U15592 (N_15592,N_14818,N_14915);
xor U15593 (N_15593,N_14616,N_14686);
and U15594 (N_15594,N_15175,N_14404);
nand U15595 (N_15595,N_14510,N_15147);
nand U15596 (N_15596,N_14875,N_15103);
nor U15597 (N_15597,N_14840,N_14810);
and U15598 (N_15598,N_14734,N_14923);
nand U15599 (N_15599,N_14412,N_14614);
or U15600 (N_15600,N_15112,N_14744);
nor U15601 (N_15601,N_14970,N_14579);
nand U15602 (N_15602,N_14994,N_14574);
nand U15603 (N_15603,N_14603,N_14611);
nand U15604 (N_15604,N_15114,N_14917);
and U15605 (N_15605,N_15016,N_14848);
and U15606 (N_15606,N_14871,N_14439);
xnor U15607 (N_15607,N_14528,N_14633);
and U15608 (N_15608,N_14889,N_14500);
and U15609 (N_15609,N_15123,N_15153);
or U15610 (N_15610,N_14812,N_15092);
nand U15611 (N_15611,N_14563,N_14786);
nor U15612 (N_15612,N_14427,N_14794);
nor U15613 (N_15613,N_15099,N_14664);
or U15614 (N_15614,N_14513,N_14537);
nor U15615 (N_15615,N_14597,N_14826);
and U15616 (N_15616,N_14922,N_14958);
or U15617 (N_15617,N_14912,N_15079);
xnor U15618 (N_15618,N_14539,N_14511);
or U15619 (N_15619,N_14929,N_14497);
nor U15620 (N_15620,N_14775,N_14685);
nand U15621 (N_15621,N_14535,N_14845);
and U15622 (N_15622,N_14459,N_14541);
nand U15623 (N_15623,N_14836,N_14676);
xnor U15624 (N_15624,N_15156,N_14480);
and U15625 (N_15625,N_14822,N_14959);
nand U15626 (N_15626,N_14714,N_14402);
nor U15627 (N_15627,N_14474,N_14549);
or U15628 (N_15628,N_14422,N_14486);
xor U15629 (N_15629,N_15100,N_14538);
nand U15630 (N_15630,N_15121,N_14678);
nand U15631 (N_15631,N_14850,N_14977);
and U15632 (N_15632,N_14685,N_14964);
or U15633 (N_15633,N_14521,N_14409);
xnor U15634 (N_15634,N_14895,N_14680);
nor U15635 (N_15635,N_14674,N_15191);
nand U15636 (N_15636,N_14622,N_15021);
and U15637 (N_15637,N_14771,N_15001);
nand U15638 (N_15638,N_14958,N_14477);
nor U15639 (N_15639,N_14557,N_14643);
xor U15640 (N_15640,N_14743,N_14954);
nor U15641 (N_15641,N_14404,N_14774);
and U15642 (N_15642,N_15012,N_14774);
nand U15643 (N_15643,N_15110,N_14520);
and U15644 (N_15644,N_14636,N_14435);
and U15645 (N_15645,N_14709,N_15045);
xnor U15646 (N_15646,N_15000,N_15181);
or U15647 (N_15647,N_15198,N_14676);
xor U15648 (N_15648,N_14502,N_15134);
nand U15649 (N_15649,N_14750,N_14458);
nor U15650 (N_15650,N_14477,N_14669);
and U15651 (N_15651,N_15024,N_14849);
xnor U15652 (N_15652,N_14546,N_14576);
or U15653 (N_15653,N_15100,N_14596);
and U15654 (N_15654,N_14841,N_14627);
nand U15655 (N_15655,N_15143,N_15011);
nor U15656 (N_15656,N_14935,N_14649);
nand U15657 (N_15657,N_14495,N_15025);
xnor U15658 (N_15658,N_15018,N_14468);
and U15659 (N_15659,N_15050,N_14715);
nor U15660 (N_15660,N_14441,N_15122);
nand U15661 (N_15661,N_15167,N_14645);
nand U15662 (N_15662,N_14662,N_14428);
or U15663 (N_15663,N_14474,N_14822);
xnor U15664 (N_15664,N_14589,N_15175);
nor U15665 (N_15665,N_14772,N_15128);
nor U15666 (N_15666,N_14813,N_14779);
or U15667 (N_15667,N_14635,N_15093);
xor U15668 (N_15668,N_14753,N_15038);
and U15669 (N_15669,N_15132,N_14927);
nand U15670 (N_15670,N_14496,N_14862);
and U15671 (N_15671,N_14927,N_14543);
nor U15672 (N_15672,N_14540,N_15141);
and U15673 (N_15673,N_14864,N_14590);
nor U15674 (N_15674,N_14991,N_15100);
xor U15675 (N_15675,N_14590,N_14881);
nand U15676 (N_15676,N_15181,N_14943);
nor U15677 (N_15677,N_15130,N_14629);
and U15678 (N_15678,N_14528,N_15125);
or U15679 (N_15679,N_15001,N_14696);
nor U15680 (N_15680,N_14894,N_14798);
nand U15681 (N_15681,N_14767,N_14556);
xor U15682 (N_15682,N_14407,N_14835);
nand U15683 (N_15683,N_14500,N_14791);
nand U15684 (N_15684,N_14545,N_15133);
or U15685 (N_15685,N_15025,N_15045);
or U15686 (N_15686,N_14404,N_15172);
xor U15687 (N_15687,N_15112,N_14971);
nand U15688 (N_15688,N_14455,N_15123);
nand U15689 (N_15689,N_14582,N_15110);
and U15690 (N_15690,N_15007,N_14531);
and U15691 (N_15691,N_14710,N_15172);
or U15692 (N_15692,N_14791,N_14673);
xnor U15693 (N_15693,N_14850,N_14707);
xnor U15694 (N_15694,N_14606,N_15009);
or U15695 (N_15695,N_14656,N_14667);
nand U15696 (N_15696,N_15095,N_15051);
nand U15697 (N_15697,N_14868,N_14882);
and U15698 (N_15698,N_14483,N_14690);
xor U15699 (N_15699,N_14944,N_14618);
and U15700 (N_15700,N_15142,N_14547);
nand U15701 (N_15701,N_14664,N_14667);
nor U15702 (N_15702,N_15175,N_15006);
or U15703 (N_15703,N_14813,N_14749);
and U15704 (N_15704,N_14576,N_15175);
xnor U15705 (N_15705,N_14821,N_14401);
and U15706 (N_15706,N_14429,N_14464);
nor U15707 (N_15707,N_14818,N_14827);
and U15708 (N_15708,N_14921,N_15142);
xnor U15709 (N_15709,N_15149,N_14428);
nand U15710 (N_15710,N_14907,N_14613);
nor U15711 (N_15711,N_14490,N_14915);
or U15712 (N_15712,N_15073,N_15000);
nor U15713 (N_15713,N_14637,N_14434);
or U15714 (N_15714,N_14561,N_15160);
nand U15715 (N_15715,N_15045,N_14477);
and U15716 (N_15716,N_14491,N_14744);
xor U15717 (N_15717,N_14593,N_14866);
and U15718 (N_15718,N_14857,N_14500);
or U15719 (N_15719,N_14633,N_14890);
nand U15720 (N_15720,N_14780,N_14979);
nor U15721 (N_15721,N_14853,N_14451);
or U15722 (N_15722,N_15052,N_15113);
or U15723 (N_15723,N_15139,N_14889);
nand U15724 (N_15724,N_14416,N_14966);
and U15725 (N_15725,N_14581,N_15074);
nand U15726 (N_15726,N_15194,N_14651);
nand U15727 (N_15727,N_14551,N_14870);
nor U15728 (N_15728,N_14574,N_14438);
and U15729 (N_15729,N_14681,N_15051);
nand U15730 (N_15730,N_14587,N_15057);
or U15731 (N_15731,N_14768,N_14443);
xnor U15732 (N_15732,N_14960,N_14988);
or U15733 (N_15733,N_14453,N_14581);
xnor U15734 (N_15734,N_14980,N_14646);
nor U15735 (N_15735,N_14921,N_14947);
and U15736 (N_15736,N_14745,N_14961);
xnor U15737 (N_15737,N_14640,N_14480);
nor U15738 (N_15738,N_14943,N_14797);
nand U15739 (N_15739,N_14776,N_14573);
or U15740 (N_15740,N_14614,N_14655);
nor U15741 (N_15741,N_14487,N_14670);
nand U15742 (N_15742,N_14513,N_14596);
and U15743 (N_15743,N_14786,N_15145);
nor U15744 (N_15744,N_14701,N_14465);
or U15745 (N_15745,N_14705,N_15181);
or U15746 (N_15746,N_15043,N_14906);
nor U15747 (N_15747,N_14740,N_14739);
xor U15748 (N_15748,N_14819,N_14971);
xor U15749 (N_15749,N_15140,N_14729);
or U15750 (N_15750,N_14751,N_14450);
xnor U15751 (N_15751,N_14971,N_14766);
nor U15752 (N_15752,N_14844,N_14819);
or U15753 (N_15753,N_14779,N_15075);
xnor U15754 (N_15754,N_14618,N_14958);
nor U15755 (N_15755,N_15045,N_15132);
and U15756 (N_15756,N_14989,N_14821);
and U15757 (N_15757,N_14960,N_14970);
xor U15758 (N_15758,N_14770,N_14756);
nand U15759 (N_15759,N_14595,N_14712);
nand U15760 (N_15760,N_14559,N_14947);
nand U15761 (N_15761,N_14724,N_14637);
xor U15762 (N_15762,N_14476,N_15066);
xor U15763 (N_15763,N_14402,N_14496);
or U15764 (N_15764,N_15061,N_14980);
or U15765 (N_15765,N_15092,N_15096);
and U15766 (N_15766,N_15180,N_14700);
xor U15767 (N_15767,N_15025,N_14669);
or U15768 (N_15768,N_14719,N_14981);
or U15769 (N_15769,N_15065,N_14540);
xor U15770 (N_15770,N_14959,N_14456);
nand U15771 (N_15771,N_14641,N_15179);
xnor U15772 (N_15772,N_14743,N_15055);
or U15773 (N_15773,N_14599,N_14501);
nand U15774 (N_15774,N_14436,N_14610);
nor U15775 (N_15775,N_14493,N_14504);
nor U15776 (N_15776,N_14430,N_14993);
and U15777 (N_15777,N_14742,N_14878);
nand U15778 (N_15778,N_14985,N_14600);
and U15779 (N_15779,N_14898,N_15019);
or U15780 (N_15780,N_15052,N_14538);
or U15781 (N_15781,N_14994,N_14441);
nor U15782 (N_15782,N_14809,N_14672);
xnor U15783 (N_15783,N_14749,N_14560);
or U15784 (N_15784,N_14544,N_14738);
and U15785 (N_15785,N_14895,N_14813);
and U15786 (N_15786,N_14976,N_14961);
xnor U15787 (N_15787,N_15159,N_14502);
nor U15788 (N_15788,N_15145,N_15176);
xnor U15789 (N_15789,N_15029,N_15134);
nand U15790 (N_15790,N_14608,N_15020);
xnor U15791 (N_15791,N_14668,N_14679);
and U15792 (N_15792,N_15178,N_14610);
nor U15793 (N_15793,N_14546,N_15126);
or U15794 (N_15794,N_14806,N_15086);
or U15795 (N_15795,N_14694,N_14538);
nor U15796 (N_15796,N_14792,N_15145);
nand U15797 (N_15797,N_14612,N_14662);
nor U15798 (N_15798,N_14896,N_15041);
nand U15799 (N_15799,N_14978,N_14918);
or U15800 (N_15800,N_14803,N_15122);
or U15801 (N_15801,N_14536,N_15132);
or U15802 (N_15802,N_15088,N_14990);
nand U15803 (N_15803,N_14965,N_14684);
nor U15804 (N_15804,N_15054,N_14719);
nand U15805 (N_15805,N_14479,N_14991);
and U15806 (N_15806,N_15118,N_14891);
nand U15807 (N_15807,N_15033,N_14832);
nor U15808 (N_15808,N_14542,N_14906);
nor U15809 (N_15809,N_14882,N_14693);
xnor U15810 (N_15810,N_14630,N_14404);
or U15811 (N_15811,N_14649,N_14906);
xor U15812 (N_15812,N_14485,N_14548);
or U15813 (N_15813,N_15180,N_14883);
or U15814 (N_15814,N_14471,N_14521);
nor U15815 (N_15815,N_14579,N_14437);
or U15816 (N_15816,N_14745,N_14584);
xnor U15817 (N_15817,N_14408,N_14482);
nor U15818 (N_15818,N_14689,N_14574);
xnor U15819 (N_15819,N_14741,N_14807);
and U15820 (N_15820,N_14589,N_14973);
xnor U15821 (N_15821,N_14554,N_14400);
xor U15822 (N_15822,N_14486,N_15101);
and U15823 (N_15823,N_14747,N_14761);
and U15824 (N_15824,N_14689,N_14705);
nor U15825 (N_15825,N_14504,N_15020);
and U15826 (N_15826,N_14864,N_15101);
xnor U15827 (N_15827,N_14822,N_15044);
nand U15828 (N_15828,N_15085,N_14411);
nand U15829 (N_15829,N_15082,N_14719);
xor U15830 (N_15830,N_14574,N_15137);
xnor U15831 (N_15831,N_14504,N_14965);
nand U15832 (N_15832,N_14828,N_15168);
or U15833 (N_15833,N_14632,N_14757);
xor U15834 (N_15834,N_15128,N_14908);
or U15835 (N_15835,N_14694,N_14677);
nand U15836 (N_15836,N_14586,N_15100);
nand U15837 (N_15837,N_14752,N_15040);
xnor U15838 (N_15838,N_14612,N_14979);
or U15839 (N_15839,N_14646,N_14488);
nand U15840 (N_15840,N_14403,N_14765);
nand U15841 (N_15841,N_14670,N_15119);
and U15842 (N_15842,N_15104,N_14736);
nand U15843 (N_15843,N_14581,N_14466);
xor U15844 (N_15844,N_15047,N_15052);
or U15845 (N_15845,N_14998,N_14660);
xnor U15846 (N_15846,N_14665,N_15171);
nor U15847 (N_15847,N_14446,N_14487);
and U15848 (N_15848,N_14540,N_14433);
and U15849 (N_15849,N_15112,N_14952);
nor U15850 (N_15850,N_14576,N_14667);
nand U15851 (N_15851,N_14772,N_14478);
or U15852 (N_15852,N_14827,N_14537);
and U15853 (N_15853,N_14531,N_14651);
and U15854 (N_15854,N_14630,N_15131);
xor U15855 (N_15855,N_14505,N_14456);
xor U15856 (N_15856,N_14797,N_14867);
or U15857 (N_15857,N_14656,N_14744);
and U15858 (N_15858,N_14566,N_14558);
and U15859 (N_15859,N_15133,N_14938);
or U15860 (N_15860,N_15197,N_14903);
xnor U15861 (N_15861,N_14541,N_14521);
nor U15862 (N_15862,N_14482,N_15179);
nor U15863 (N_15863,N_14724,N_14899);
nand U15864 (N_15864,N_15140,N_14691);
or U15865 (N_15865,N_15147,N_14761);
nand U15866 (N_15866,N_15041,N_14496);
or U15867 (N_15867,N_14948,N_14851);
nand U15868 (N_15868,N_15156,N_15195);
or U15869 (N_15869,N_14454,N_14781);
and U15870 (N_15870,N_14876,N_14700);
nor U15871 (N_15871,N_14500,N_14414);
xor U15872 (N_15872,N_14547,N_14699);
and U15873 (N_15873,N_14418,N_14604);
and U15874 (N_15874,N_15139,N_14428);
nand U15875 (N_15875,N_14474,N_15043);
and U15876 (N_15876,N_15123,N_15127);
nor U15877 (N_15877,N_14674,N_14881);
nand U15878 (N_15878,N_15030,N_14761);
xnor U15879 (N_15879,N_14725,N_14953);
and U15880 (N_15880,N_14887,N_15153);
nor U15881 (N_15881,N_15049,N_14537);
or U15882 (N_15882,N_14582,N_14473);
and U15883 (N_15883,N_14911,N_15072);
nand U15884 (N_15884,N_14547,N_14766);
or U15885 (N_15885,N_14998,N_15094);
nor U15886 (N_15886,N_14719,N_14671);
or U15887 (N_15887,N_15063,N_14994);
nand U15888 (N_15888,N_14432,N_14490);
or U15889 (N_15889,N_14961,N_14620);
and U15890 (N_15890,N_15161,N_14755);
nand U15891 (N_15891,N_15012,N_15143);
xor U15892 (N_15892,N_14673,N_14959);
nand U15893 (N_15893,N_14759,N_14769);
nor U15894 (N_15894,N_14527,N_15126);
xnor U15895 (N_15895,N_15109,N_14981);
or U15896 (N_15896,N_15152,N_14649);
xor U15897 (N_15897,N_15195,N_15167);
and U15898 (N_15898,N_14560,N_15079);
xor U15899 (N_15899,N_14592,N_15163);
or U15900 (N_15900,N_15192,N_14521);
and U15901 (N_15901,N_14991,N_14754);
or U15902 (N_15902,N_14416,N_15142);
nor U15903 (N_15903,N_15031,N_14940);
nand U15904 (N_15904,N_14678,N_15178);
nand U15905 (N_15905,N_15130,N_15010);
nor U15906 (N_15906,N_14820,N_14440);
nand U15907 (N_15907,N_15173,N_15097);
nor U15908 (N_15908,N_14458,N_14546);
nand U15909 (N_15909,N_14856,N_14519);
or U15910 (N_15910,N_14971,N_14442);
nor U15911 (N_15911,N_14922,N_14698);
nand U15912 (N_15912,N_14492,N_14744);
nand U15913 (N_15913,N_14707,N_14787);
xor U15914 (N_15914,N_15163,N_14654);
nand U15915 (N_15915,N_15162,N_14573);
and U15916 (N_15916,N_14979,N_14936);
or U15917 (N_15917,N_15128,N_14704);
or U15918 (N_15918,N_14846,N_14811);
nand U15919 (N_15919,N_14755,N_14952);
xnor U15920 (N_15920,N_14551,N_14673);
or U15921 (N_15921,N_14748,N_15038);
or U15922 (N_15922,N_14806,N_15171);
nor U15923 (N_15923,N_14528,N_14746);
nor U15924 (N_15924,N_14885,N_15082);
or U15925 (N_15925,N_15102,N_14985);
xnor U15926 (N_15926,N_14556,N_14522);
or U15927 (N_15927,N_15124,N_14566);
or U15928 (N_15928,N_14829,N_14453);
nor U15929 (N_15929,N_14431,N_15112);
nand U15930 (N_15930,N_14959,N_14520);
nand U15931 (N_15931,N_15151,N_14992);
nor U15932 (N_15932,N_14669,N_14694);
xor U15933 (N_15933,N_14653,N_15031);
or U15934 (N_15934,N_15061,N_15004);
or U15935 (N_15935,N_15193,N_14478);
xnor U15936 (N_15936,N_14420,N_14964);
or U15937 (N_15937,N_14570,N_15060);
xor U15938 (N_15938,N_14547,N_14627);
nor U15939 (N_15939,N_14958,N_14661);
or U15940 (N_15940,N_14830,N_14661);
nor U15941 (N_15941,N_15166,N_14857);
and U15942 (N_15942,N_14403,N_14632);
and U15943 (N_15943,N_14954,N_15108);
nor U15944 (N_15944,N_14979,N_14824);
xor U15945 (N_15945,N_15008,N_14781);
nand U15946 (N_15946,N_14844,N_14813);
xnor U15947 (N_15947,N_14435,N_15058);
or U15948 (N_15948,N_14722,N_14904);
and U15949 (N_15949,N_14829,N_14521);
nor U15950 (N_15950,N_14413,N_14969);
or U15951 (N_15951,N_14627,N_14802);
nor U15952 (N_15952,N_14425,N_15132);
and U15953 (N_15953,N_14603,N_14881);
and U15954 (N_15954,N_14624,N_14986);
nand U15955 (N_15955,N_14728,N_14927);
and U15956 (N_15956,N_14902,N_15068);
nor U15957 (N_15957,N_14897,N_14401);
xor U15958 (N_15958,N_14465,N_15018);
xnor U15959 (N_15959,N_14999,N_15001);
and U15960 (N_15960,N_14932,N_14710);
and U15961 (N_15961,N_14418,N_14975);
nand U15962 (N_15962,N_14508,N_15165);
nand U15963 (N_15963,N_14977,N_15084);
nor U15964 (N_15964,N_14871,N_15018);
nor U15965 (N_15965,N_15064,N_14426);
xor U15966 (N_15966,N_14467,N_14807);
or U15967 (N_15967,N_14924,N_15007);
or U15968 (N_15968,N_14501,N_14932);
nor U15969 (N_15969,N_14518,N_14960);
and U15970 (N_15970,N_14440,N_15059);
xnor U15971 (N_15971,N_14774,N_15099);
xnor U15972 (N_15972,N_14711,N_14606);
xor U15973 (N_15973,N_15089,N_15040);
xnor U15974 (N_15974,N_15017,N_15161);
and U15975 (N_15975,N_15069,N_14672);
or U15976 (N_15976,N_14743,N_14512);
xor U15977 (N_15977,N_15016,N_14783);
nor U15978 (N_15978,N_14824,N_14458);
nor U15979 (N_15979,N_14995,N_14597);
nor U15980 (N_15980,N_14404,N_14903);
and U15981 (N_15981,N_14692,N_14769);
nor U15982 (N_15982,N_14879,N_14595);
nand U15983 (N_15983,N_15076,N_14615);
nor U15984 (N_15984,N_14804,N_14671);
xnor U15985 (N_15985,N_14494,N_14401);
xor U15986 (N_15986,N_15026,N_14562);
nor U15987 (N_15987,N_14822,N_14741);
or U15988 (N_15988,N_14848,N_14435);
nor U15989 (N_15989,N_14414,N_14803);
nand U15990 (N_15990,N_14594,N_14731);
nor U15991 (N_15991,N_15116,N_14754);
nand U15992 (N_15992,N_14494,N_14701);
nand U15993 (N_15993,N_14678,N_14962);
nand U15994 (N_15994,N_14544,N_14720);
nor U15995 (N_15995,N_14672,N_15094);
xor U15996 (N_15996,N_14749,N_14641);
or U15997 (N_15997,N_14829,N_15125);
nor U15998 (N_15998,N_14678,N_14796);
nand U15999 (N_15999,N_14431,N_14481);
and U16000 (N_16000,N_15952,N_15653);
or U16001 (N_16001,N_15771,N_15574);
xnor U16002 (N_16002,N_15210,N_15793);
and U16003 (N_16003,N_15645,N_15789);
nand U16004 (N_16004,N_15742,N_15202);
or U16005 (N_16005,N_15740,N_15205);
and U16006 (N_16006,N_15635,N_15241);
or U16007 (N_16007,N_15890,N_15569);
or U16008 (N_16008,N_15478,N_15283);
or U16009 (N_16009,N_15868,N_15856);
nand U16010 (N_16010,N_15228,N_15357);
and U16011 (N_16011,N_15258,N_15200);
nor U16012 (N_16012,N_15440,N_15932);
and U16013 (N_16013,N_15593,N_15577);
nor U16014 (N_16014,N_15855,N_15927);
nor U16015 (N_16015,N_15797,N_15829);
and U16016 (N_16016,N_15989,N_15735);
xnor U16017 (N_16017,N_15947,N_15350);
nand U16018 (N_16018,N_15631,N_15758);
xor U16019 (N_16019,N_15754,N_15570);
nand U16020 (N_16020,N_15521,N_15462);
nor U16021 (N_16021,N_15415,N_15779);
xnor U16022 (N_16022,N_15416,N_15900);
nor U16023 (N_16023,N_15311,N_15482);
nand U16024 (N_16024,N_15411,N_15883);
nand U16025 (N_16025,N_15839,N_15527);
nand U16026 (N_16026,N_15825,N_15343);
or U16027 (N_16027,N_15626,N_15409);
nand U16028 (N_16028,N_15379,N_15854);
or U16029 (N_16029,N_15360,N_15365);
nor U16030 (N_16030,N_15845,N_15559);
and U16031 (N_16031,N_15792,N_15656);
nand U16032 (N_16032,N_15345,N_15991);
or U16033 (N_16033,N_15461,N_15284);
nor U16034 (N_16034,N_15293,N_15816);
or U16035 (N_16035,N_15726,N_15739);
nand U16036 (N_16036,N_15992,N_15933);
nor U16037 (N_16037,N_15451,N_15919);
or U16038 (N_16038,N_15873,N_15308);
and U16039 (N_16039,N_15606,N_15764);
and U16040 (N_16040,N_15965,N_15326);
nand U16041 (N_16041,N_15295,N_15857);
nand U16042 (N_16042,N_15806,N_15619);
xnor U16043 (N_16043,N_15353,N_15436);
and U16044 (N_16044,N_15419,N_15807);
nand U16045 (N_16045,N_15398,N_15375);
xnor U16046 (N_16046,N_15836,N_15352);
nand U16047 (N_16047,N_15494,N_15601);
nor U16048 (N_16048,N_15460,N_15324);
xnor U16049 (N_16049,N_15891,N_15782);
nand U16050 (N_16050,N_15406,N_15566);
and U16051 (N_16051,N_15784,N_15230);
or U16052 (N_16052,N_15207,N_15731);
or U16053 (N_16053,N_15564,N_15307);
xor U16054 (N_16054,N_15982,N_15979);
or U16055 (N_16055,N_15310,N_15812);
and U16056 (N_16056,N_15496,N_15376);
and U16057 (N_16057,N_15425,N_15795);
nand U16058 (N_16058,N_15568,N_15753);
or U16059 (N_16059,N_15562,N_15649);
nand U16060 (N_16060,N_15351,N_15516);
or U16061 (N_16061,N_15604,N_15214);
and U16062 (N_16062,N_15897,N_15558);
or U16063 (N_16063,N_15655,N_15430);
nand U16064 (N_16064,N_15648,N_15944);
or U16065 (N_16065,N_15776,N_15773);
nand U16066 (N_16066,N_15849,N_15305);
xnor U16067 (N_16067,N_15251,N_15707);
xor U16068 (N_16068,N_15634,N_15701);
nand U16069 (N_16069,N_15341,N_15203);
nand U16070 (N_16070,N_15468,N_15372);
or U16071 (N_16071,N_15605,N_15957);
xnor U16072 (N_16072,N_15234,N_15628);
xor U16073 (N_16073,N_15522,N_15930);
nor U16074 (N_16074,N_15866,N_15774);
xor U16075 (N_16075,N_15955,N_15640);
xnor U16076 (N_16076,N_15909,N_15389);
nor U16077 (N_16077,N_15863,N_15526);
xnor U16078 (N_16078,N_15444,N_15543);
or U16079 (N_16079,N_15831,N_15449);
nand U16080 (N_16080,N_15560,N_15722);
nor U16081 (N_16081,N_15368,N_15412);
xnor U16082 (N_16082,N_15745,N_15408);
nand U16083 (N_16083,N_15996,N_15373);
xor U16084 (N_16084,N_15281,N_15708);
xnor U16085 (N_16085,N_15322,N_15498);
nor U16086 (N_16086,N_15392,N_15622);
xnor U16087 (N_16087,N_15715,N_15396);
nor U16088 (N_16088,N_15312,N_15859);
xnor U16089 (N_16089,N_15910,N_15928);
or U16090 (N_16090,N_15956,N_15611);
nand U16091 (N_16091,N_15269,N_15475);
and U16092 (N_16092,N_15388,N_15509);
nor U16093 (N_16093,N_15934,N_15778);
nor U16094 (N_16094,N_15867,N_15366);
nand U16095 (N_16095,N_15524,N_15877);
xor U16096 (N_16096,N_15862,N_15476);
nand U16097 (N_16097,N_15751,N_15621);
or U16098 (N_16098,N_15297,N_15765);
and U16099 (N_16099,N_15805,N_15688);
nand U16100 (N_16100,N_15960,N_15507);
nand U16101 (N_16101,N_15684,N_15788);
nand U16102 (N_16102,N_15329,N_15222);
nor U16103 (N_16103,N_15644,N_15404);
and U16104 (N_16104,N_15809,N_15441);
nand U16105 (N_16105,N_15698,N_15964);
nand U16106 (N_16106,N_15733,N_15837);
or U16107 (N_16107,N_15447,N_15950);
xnor U16108 (N_16108,N_15282,N_15827);
xor U16109 (N_16109,N_15629,N_15268);
or U16110 (N_16110,N_15467,N_15658);
nand U16111 (N_16111,N_15869,N_15725);
nor U16112 (N_16112,N_15880,N_15889);
and U16113 (N_16113,N_15572,N_15850);
nor U16114 (N_16114,N_15591,N_15670);
or U16115 (N_16115,N_15671,N_15563);
nand U16116 (N_16116,N_15995,N_15663);
and U16117 (N_16117,N_15987,N_15908);
or U16118 (N_16118,N_15677,N_15508);
nor U16119 (N_16119,N_15465,N_15453);
xnor U16120 (N_16120,N_15901,N_15780);
and U16121 (N_16121,N_15719,N_15413);
nand U16122 (N_16122,N_15612,N_15975);
nor U16123 (N_16123,N_15358,N_15935);
nor U16124 (N_16124,N_15215,N_15720);
or U16125 (N_16125,N_15800,N_15401);
and U16126 (N_16126,N_15362,N_15700);
nand U16127 (N_16127,N_15811,N_15598);
or U16128 (N_16128,N_15843,N_15844);
nor U16129 (N_16129,N_15973,N_15246);
xnor U16130 (N_16130,N_15749,N_15617);
and U16131 (N_16131,N_15875,N_15355);
and U16132 (N_16132,N_15669,N_15840);
nor U16133 (N_16133,N_15942,N_15969);
xnor U16134 (N_16134,N_15233,N_15954);
xnor U16135 (N_16135,N_15405,N_15301);
and U16136 (N_16136,N_15492,N_15378);
xnor U16137 (N_16137,N_15948,N_15431);
xnor U16138 (N_16138,N_15266,N_15256);
nor U16139 (N_16139,N_15990,N_15984);
nand U16140 (N_16140,N_15518,N_15680);
xnor U16141 (N_16141,N_15294,N_15832);
xor U16142 (N_16142,N_15292,N_15999);
and U16143 (N_16143,N_15924,N_15819);
nor U16144 (N_16144,N_15822,N_15298);
or U16145 (N_16145,N_15512,N_15446);
or U16146 (N_16146,N_15918,N_15519);
xnor U16147 (N_16147,N_15813,N_15732);
and U16148 (N_16148,N_15319,N_15466);
or U16149 (N_16149,N_15586,N_15403);
and U16150 (N_16150,N_15278,N_15736);
nor U16151 (N_16151,N_15250,N_15483);
and U16152 (N_16152,N_15511,N_15445);
nand U16153 (N_16153,N_15766,N_15510);
and U16154 (N_16154,N_15993,N_15639);
or U16155 (N_16155,N_15291,N_15998);
or U16156 (N_16156,N_15255,N_15699);
nand U16157 (N_16157,N_15347,N_15280);
nand U16158 (N_16158,N_15390,N_15463);
nand U16159 (N_16159,N_15479,N_15226);
xnor U16160 (N_16160,N_15450,N_15978);
nand U16161 (N_16161,N_15717,N_15770);
or U16162 (N_16162,N_15874,N_15435);
and U16163 (N_16163,N_15363,N_15976);
and U16164 (N_16164,N_15642,N_15876);
xor U16165 (N_16165,N_15879,N_15470);
nand U16166 (N_16166,N_15905,N_15369);
and U16167 (N_16167,N_15480,N_15321);
xor U16168 (N_16168,N_15588,N_15781);
nor U16169 (N_16169,N_15206,N_15530);
or U16170 (N_16170,N_15513,N_15439);
nor U16171 (N_16171,N_15683,N_15387);
or U16172 (N_16172,N_15240,N_15276);
and U16173 (N_16173,N_15824,N_15608);
or U16174 (N_16174,N_15499,N_15916);
or U16175 (N_16175,N_15296,N_15534);
and U16176 (N_16176,N_15437,N_15971);
nand U16177 (N_16177,N_15555,N_15624);
nand U16178 (N_16178,N_15791,N_15647);
or U16179 (N_16179,N_15917,N_15469);
and U16180 (N_16180,N_15665,N_15864);
and U16181 (N_16181,N_15761,N_15473);
xor U16182 (N_16182,N_15625,N_15356);
and U16183 (N_16183,N_15912,N_15615);
or U16184 (N_16184,N_15898,N_15994);
xor U16185 (N_16185,N_15676,N_15861);
nand U16186 (N_16186,N_15838,N_15364);
nand U16187 (N_16187,N_15486,N_15865);
xnor U16188 (N_16188,N_15249,N_15209);
nor U16189 (N_16189,N_15385,N_15841);
or U16190 (N_16190,N_15424,N_15886);
nand U16191 (N_16191,N_15495,N_15595);
nand U16192 (N_16192,N_15659,N_15941);
nor U16193 (N_16193,N_15231,N_15277);
nand U16194 (N_16194,N_15211,N_15888);
xor U16195 (N_16195,N_15237,N_15983);
nor U16196 (N_16196,N_15737,N_15515);
and U16197 (N_16197,N_15454,N_15506);
or U16198 (N_16198,N_15804,N_15734);
and U16199 (N_16199,N_15554,N_15940);
nand U16200 (N_16200,N_15536,N_15968);
xor U16201 (N_16201,N_15528,N_15661);
xor U16202 (N_16202,N_15275,N_15452);
nand U16203 (N_16203,N_15216,N_15455);
nor U16204 (N_16204,N_15585,N_15252);
or U16205 (N_16205,N_15420,N_15287);
nand U16206 (N_16206,N_15433,N_15920);
xor U16207 (N_16207,N_15911,N_15582);
or U16208 (N_16208,N_15485,N_15896);
and U16209 (N_16209,N_15235,N_15744);
nand U16210 (N_16210,N_15961,N_15710);
nand U16211 (N_16211,N_15820,N_15504);
or U16212 (N_16212,N_15223,N_15946);
nand U16213 (N_16213,N_15520,N_15525);
xor U16214 (N_16214,N_15418,N_15730);
or U16215 (N_16215,N_15422,N_15963);
xnor U16216 (N_16216,N_15220,N_15828);
and U16217 (N_16217,N_15686,N_15977);
xor U16218 (N_16218,N_15381,N_15673);
xor U16219 (N_16219,N_15623,N_15336);
or U16220 (N_16220,N_15833,N_15383);
xnor U16221 (N_16221,N_15456,N_15721);
nor U16222 (N_16222,N_15464,N_15714);
or U16223 (N_16223,N_15974,N_15288);
nor U16224 (N_16224,N_15929,N_15887);
nor U16225 (N_16225,N_15892,N_15633);
nand U16226 (N_16226,N_15627,N_15318);
nand U16227 (N_16227,N_15386,N_15253);
or U16228 (N_16228,N_15583,N_15741);
or U16229 (N_16229,N_15902,N_15922);
xnor U16230 (N_16230,N_15335,N_15858);
xnor U16231 (N_16231,N_15236,N_15748);
and U16232 (N_16232,N_15692,N_15218);
or U16233 (N_16233,N_15772,N_15229);
nand U16234 (N_16234,N_15344,N_15402);
xnor U16235 (N_16235,N_15762,N_15501);
and U16236 (N_16236,N_15613,N_15641);
or U16237 (N_16237,N_15219,N_15632);
nor U16238 (N_16238,N_15325,N_15662);
nand U16239 (N_16239,N_15395,N_15986);
nor U16240 (N_16240,N_15471,N_15337);
xnor U16241 (N_16241,N_15915,N_15729);
and U16242 (N_16242,N_15505,N_15798);
and U16243 (N_16243,N_15967,N_15636);
and U16244 (N_16244,N_15279,N_15327);
and U16245 (N_16245,N_15339,N_15417);
or U16246 (N_16246,N_15666,N_15548);
and U16247 (N_16247,N_15760,N_15893);
and U16248 (N_16248,N_15904,N_15382);
xor U16249 (N_16249,N_15539,N_15303);
nor U16250 (N_16250,N_15738,N_15302);
and U16251 (N_16251,N_15472,N_15340);
xor U16252 (N_16252,N_15263,N_15238);
nor U16253 (N_16253,N_15367,N_15227);
nand U16254 (N_16254,N_15575,N_15985);
or U16255 (N_16255,N_15607,N_15980);
xnor U16256 (N_16256,N_15550,N_15571);
xor U16257 (N_16257,N_15429,N_15217);
and U16258 (N_16258,N_15926,N_15428);
and U16259 (N_16259,N_15851,N_15407);
nand U16260 (N_16260,N_15848,N_15300);
xor U16261 (N_16261,N_15533,N_15652);
nand U16262 (N_16262,N_15556,N_15675);
nor U16263 (N_16263,N_15618,N_15306);
and U16264 (N_16264,N_15602,N_15697);
or U16265 (N_16265,N_15399,N_15690);
nor U16266 (N_16266,N_15664,N_15245);
xor U16267 (N_16267,N_15815,N_15860);
nand U16268 (N_16268,N_15212,N_15966);
nand U16269 (N_16269,N_15384,N_15576);
and U16270 (N_16270,N_15338,N_15224);
xor U16271 (N_16271,N_15884,N_15532);
and U16272 (N_16272,N_15592,N_15657);
nand U16273 (N_16273,N_15668,N_15535);
nor U16274 (N_16274,N_15921,N_15332);
or U16275 (N_16275,N_15903,N_15342);
or U16276 (N_16276,N_15201,N_15981);
nor U16277 (N_16277,N_15557,N_15544);
and U16278 (N_16278,N_15654,N_15316);
xnor U16279 (N_16279,N_15242,N_15442);
and U16280 (N_16280,N_15400,N_15561);
nor U16281 (N_16281,N_15313,N_15620);
nor U16282 (N_16282,N_15552,N_15746);
and U16283 (N_16283,N_15796,N_15247);
or U16284 (N_16284,N_15580,N_15538);
nand U16285 (N_16285,N_15274,N_15354);
xnor U16286 (N_16286,N_15551,N_15490);
nand U16287 (N_16287,N_15438,N_15531);
and U16288 (N_16288,N_15882,N_15775);
xor U16289 (N_16289,N_15938,N_15204);
or U16290 (N_16290,N_15899,N_15785);
xor U16291 (N_16291,N_15759,N_15945);
nand U16292 (N_16292,N_15881,N_15799);
nand U16293 (N_16293,N_15630,N_15315);
nor U16294 (N_16294,N_15728,N_15410);
and U16295 (N_16295,N_15810,N_15594);
and U16296 (N_16296,N_15427,N_15801);
xor U16297 (N_16297,N_15380,N_15702);
xnor U16298 (N_16298,N_15239,N_15988);
nor U16299 (N_16299,N_15747,N_15549);
nand U16300 (N_16300,N_15743,N_15553);
and U16301 (N_16301,N_15691,N_15757);
xnor U16302 (N_16302,N_15584,N_15484);
or U16303 (N_16303,N_15763,N_15711);
or U16304 (N_16304,N_15646,N_15299);
or U16305 (N_16305,N_15448,N_15213);
xor U16306 (N_16306,N_15872,N_15481);
and U16307 (N_16307,N_15545,N_15755);
or U16308 (N_16308,N_15286,N_15264);
and U16309 (N_16309,N_15225,N_15870);
nor U16310 (N_16310,N_15913,N_15232);
nor U16311 (N_16311,N_15808,N_15579);
xnor U16312 (N_16312,N_15959,N_15477);
or U16313 (N_16313,N_15638,N_15529);
nor U16314 (N_16314,N_15871,N_15939);
and U16315 (N_16315,N_15500,N_15457);
and U16316 (N_16316,N_15346,N_15434);
nor U16317 (N_16317,N_15958,N_15273);
nand U16318 (N_16318,N_15589,N_15578);
xor U16319 (N_16319,N_15547,N_15257);
nand U16320 (N_16320,N_15567,N_15503);
nand U16321 (N_16321,N_15374,N_15330);
or U16322 (N_16322,N_15260,N_15709);
or U16323 (N_16323,N_15943,N_15678);
or U16324 (N_16324,N_15681,N_15923);
nand U16325 (N_16325,N_15846,N_15493);
xor U16326 (N_16326,N_15818,N_15514);
or U16327 (N_16327,N_15637,N_15794);
nand U16328 (N_16328,N_15320,N_15672);
and U16329 (N_16329,N_15706,N_15650);
and U16330 (N_16330,N_15581,N_15423);
and U16331 (N_16331,N_15750,N_15331);
nand U16332 (N_16332,N_15285,N_15651);
xnor U16333 (N_16333,N_15685,N_15289);
xor U16334 (N_16334,N_15459,N_15616);
or U16335 (N_16335,N_15970,N_15596);
or U16336 (N_16336,N_15272,N_15487);
xnor U16337 (N_16337,N_15361,N_15823);
and U16338 (N_16338,N_15716,N_15769);
nor U16339 (N_16339,N_15667,N_15783);
nand U16340 (N_16340,N_15371,N_15502);
and U16341 (N_16341,N_15704,N_15936);
xnor U16342 (N_16342,N_15397,N_15600);
or U16343 (N_16343,N_15705,N_15643);
xnor U16344 (N_16344,N_15696,N_15718);
and U16345 (N_16345,N_15852,N_15540);
nand U16346 (N_16346,N_15682,N_15370);
and U16347 (N_16347,N_15674,N_15565);
and U16348 (N_16348,N_15694,N_15814);
nor U16349 (N_16349,N_15393,N_15787);
nor U16350 (N_16350,N_15573,N_15541);
xnor U16351 (N_16351,N_15972,N_15907);
or U16352 (N_16352,N_15727,N_15817);
or U16353 (N_16353,N_15270,N_15786);
xor U16354 (N_16354,N_15951,N_15842);
and U16355 (N_16355,N_15895,N_15885);
nand U16356 (N_16356,N_15333,N_15914);
nand U16357 (N_16357,N_15489,N_15997);
nor U16358 (N_16358,N_15309,N_15304);
nor U16359 (N_16359,N_15474,N_15208);
and U16360 (N_16360,N_15262,N_15949);
or U16361 (N_16361,N_15713,N_15853);
and U16362 (N_16362,N_15348,N_15687);
and U16363 (N_16363,N_15894,N_15610);
or U16364 (N_16364,N_15328,N_15497);
and U16365 (N_16365,N_15752,N_15432);
xnor U16366 (N_16366,N_15394,N_15314);
nor U16367 (N_16367,N_15254,N_15414);
or U16368 (N_16368,N_15517,N_15826);
nand U16369 (N_16369,N_15803,N_15359);
and U16370 (N_16370,N_15614,N_15834);
and U16371 (N_16371,N_15878,N_15821);
nor U16372 (N_16372,N_15847,N_15660);
nor U16373 (N_16373,N_15790,N_15458);
or U16374 (N_16374,N_15777,N_15377);
nand U16375 (N_16375,N_15723,N_15259);
nand U16376 (N_16376,N_15597,N_15937);
nor U16377 (N_16377,N_15599,N_15590);
xor U16378 (N_16378,N_15609,N_15523);
nor U16379 (N_16379,N_15689,N_15603);
xor U16380 (N_16380,N_15962,N_15835);
nand U16381 (N_16381,N_15421,N_15693);
nor U16382 (N_16382,N_15724,N_15906);
or U16383 (N_16383,N_15243,N_15349);
xnor U16384 (N_16384,N_15443,N_15767);
and U16385 (N_16385,N_15830,N_15703);
and U16386 (N_16386,N_15244,N_15221);
or U16387 (N_16387,N_15265,N_15802);
nor U16388 (N_16388,N_15391,N_15587);
nand U16389 (N_16389,N_15695,N_15768);
nor U16390 (N_16390,N_15334,N_15271);
xor U16391 (N_16391,N_15756,N_15679);
xnor U16392 (N_16392,N_15267,N_15931);
nor U16393 (N_16393,N_15290,N_15261);
and U16394 (N_16394,N_15317,N_15248);
and U16395 (N_16395,N_15491,N_15426);
xnor U16396 (N_16396,N_15953,N_15712);
xnor U16397 (N_16397,N_15488,N_15925);
nor U16398 (N_16398,N_15542,N_15323);
xnor U16399 (N_16399,N_15537,N_15546);
and U16400 (N_16400,N_15544,N_15415);
nand U16401 (N_16401,N_15990,N_15361);
xnor U16402 (N_16402,N_15832,N_15960);
and U16403 (N_16403,N_15742,N_15908);
xnor U16404 (N_16404,N_15811,N_15391);
nor U16405 (N_16405,N_15239,N_15309);
nand U16406 (N_16406,N_15910,N_15946);
xnor U16407 (N_16407,N_15664,N_15901);
xor U16408 (N_16408,N_15560,N_15922);
or U16409 (N_16409,N_15460,N_15601);
and U16410 (N_16410,N_15246,N_15554);
nor U16411 (N_16411,N_15559,N_15669);
and U16412 (N_16412,N_15935,N_15307);
or U16413 (N_16413,N_15506,N_15550);
and U16414 (N_16414,N_15689,N_15705);
or U16415 (N_16415,N_15433,N_15666);
nor U16416 (N_16416,N_15784,N_15438);
xnor U16417 (N_16417,N_15968,N_15649);
xnor U16418 (N_16418,N_15790,N_15892);
nor U16419 (N_16419,N_15765,N_15414);
or U16420 (N_16420,N_15942,N_15391);
xor U16421 (N_16421,N_15918,N_15312);
or U16422 (N_16422,N_15334,N_15975);
xnor U16423 (N_16423,N_15244,N_15593);
or U16424 (N_16424,N_15881,N_15691);
and U16425 (N_16425,N_15965,N_15847);
and U16426 (N_16426,N_15368,N_15913);
nor U16427 (N_16427,N_15872,N_15743);
xnor U16428 (N_16428,N_15993,N_15663);
nand U16429 (N_16429,N_15878,N_15757);
and U16430 (N_16430,N_15591,N_15859);
xnor U16431 (N_16431,N_15591,N_15775);
or U16432 (N_16432,N_15769,N_15553);
nand U16433 (N_16433,N_15635,N_15760);
xnor U16434 (N_16434,N_15606,N_15849);
or U16435 (N_16435,N_15398,N_15496);
nand U16436 (N_16436,N_15388,N_15578);
and U16437 (N_16437,N_15595,N_15669);
xor U16438 (N_16438,N_15487,N_15454);
nor U16439 (N_16439,N_15393,N_15972);
nand U16440 (N_16440,N_15775,N_15513);
or U16441 (N_16441,N_15399,N_15964);
or U16442 (N_16442,N_15506,N_15465);
or U16443 (N_16443,N_15549,N_15320);
or U16444 (N_16444,N_15895,N_15689);
nor U16445 (N_16445,N_15602,N_15281);
nand U16446 (N_16446,N_15205,N_15272);
or U16447 (N_16447,N_15632,N_15255);
or U16448 (N_16448,N_15828,N_15372);
nand U16449 (N_16449,N_15320,N_15295);
and U16450 (N_16450,N_15502,N_15326);
nand U16451 (N_16451,N_15264,N_15906);
nand U16452 (N_16452,N_15507,N_15485);
or U16453 (N_16453,N_15643,N_15430);
xor U16454 (N_16454,N_15541,N_15396);
and U16455 (N_16455,N_15213,N_15895);
or U16456 (N_16456,N_15900,N_15385);
and U16457 (N_16457,N_15437,N_15481);
xnor U16458 (N_16458,N_15777,N_15586);
and U16459 (N_16459,N_15364,N_15608);
nand U16460 (N_16460,N_15646,N_15675);
or U16461 (N_16461,N_15332,N_15388);
nor U16462 (N_16462,N_15591,N_15826);
nor U16463 (N_16463,N_15948,N_15621);
or U16464 (N_16464,N_15862,N_15661);
xor U16465 (N_16465,N_15821,N_15645);
xor U16466 (N_16466,N_15864,N_15744);
nor U16467 (N_16467,N_15973,N_15729);
and U16468 (N_16468,N_15726,N_15529);
xnor U16469 (N_16469,N_15757,N_15525);
and U16470 (N_16470,N_15526,N_15674);
xor U16471 (N_16471,N_15693,N_15420);
and U16472 (N_16472,N_15888,N_15230);
nor U16473 (N_16473,N_15674,N_15890);
nand U16474 (N_16474,N_15202,N_15567);
xor U16475 (N_16475,N_15992,N_15962);
or U16476 (N_16476,N_15799,N_15266);
nand U16477 (N_16477,N_15206,N_15444);
nor U16478 (N_16478,N_15633,N_15464);
and U16479 (N_16479,N_15840,N_15838);
xor U16480 (N_16480,N_15298,N_15585);
nand U16481 (N_16481,N_15700,N_15734);
or U16482 (N_16482,N_15692,N_15402);
xor U16483 (N_16483,N_15599,N_15404);
or U16484 (N_16484,N_15549,N_15932);
and U16485 (N_16485,N_15730,N_15235);
and U16486 (N_16486,N_15891,N_15952);
and U16487 (N_16487,N_15422,N_15928);
nand U16488 (N_16488,N_15382,N_15415);
or U16489 (N_16489,N_15386,N_15463);
xor U16490 (N_16490,N_15909,N_15212);
or U16491 (N_16491,N_15329,N_15731);
xnor U16492 (N_16492,N_15898,N_15932);
or U16493 (N_16493,N_15612,N_15732);
or U16494 (N_16494,N_15349,N_15675);
xor U16495 (N_16495,N_15224,N_15807);
nor U16496 (N_16496,N_15960,N_15617);
and U16497 (N_16497,N_15225,N_15495);
nand U16498 (N_16498,N_15924,N_15506);
xnor U16499 (N_16499,N_15722,N_15729);
or U16500 (N_16500,N_15482,N_15493);
or U16501 (N_16501,N_15692,N_15542);
nand U16502 (N_16502,N_15895,N_15273);
nor U16503 (N_16503,N_15692,N_15691);
and U16504 (N_16504,N_15556,N_15249);
xnor U16505 (N_16505,N_15954,N_15377);
and U16506 (N_16506,N_15494,N_15687);
xnor U16507 (N_16507,N_15600,N_15531);
nor U16508 (N_16508,N_15315,N_15371);
and U16509 (N_16509,N_15207,N_15297);
xnor U16510 (N_16510,N_15739,N_15478);
nand U16511 (N_16511,N_15784,N_15852);
nor U16512 (N_16512,N_15969,N_15339);
xnor U16513 (N_16513,N_15494,N_15928);
nand U16514 (N_16514,N_15343,N_15747);
nand U16515 (N_16515,N_15714,N_15841);
xnor U16516 (N_16516,N_15396,N_15224);
or U16517 (N_16517,N_15290,N_15574);
and U16518 (N_16518,N_15555,N_15538);
nand U16519 (N_16519,N_15658,N_15639);
or U16520 (N_16520,N_15681,N_15333);
nor U16521 (N_16521,N_15557,N_15552);
or U16522 (N_16522,N_15750,N_15973);
nand U16523 (N_16523,N_15758,N_15476);
xor U16524 (N_16524,N_15975,N_15553);
or U16525 (N_16525,N_15803,N_15779);
or U16526 (N_16526,N_15243,N_15315);
and U16527 (N_16527,N_15962,N_15634);
and U16528 (N_16528,N_15472,N_15742);
and U16529 (N_16529,N_15959,N_15591);
nand U16530 (N_16530,N_15425,N_15630);
xor U16531 (N_16531,N_15651,N_15906);
nor U16532 (N_16532,N_15373,N_15564);
nand U16533 (N_16533,N_15604,N_15576);
xor U16534 (N_16534,N_15210,N_15761);
nand U16535 (N_16535,N_15419,N_15255);
nor U16536 (N_16536,N_15869,N_15785);
nor U16537 (N_16537,N_15408,N_15601);
and U16538 (N_16538,N_15919,N_15750);
or U16539 (N_16539,N_15372,N_15579);
nand U16540 (N_16540,N_15969,N_15376);
nand U16541 (N_16541,N_15748,N_15790);
xor U16542 (N_16542,N_15434,N_15282);
nand U16543 (N_16543,N_15525,N_15471);
or U16544 (N_16544,N_15252,N_15219);
and U16545 (N_16545,N_15515,N_15411);
nor U16546 (N_16546,N_15768,N_15803);
or U16547 (N_16547,N_15693,N_15492);
nor U16548 (N_16548,N_15416,N_15519);
nor U16549 (N_16549,N_15281,N_15709);
nand U16550 (N_16550,N_15336,N_15858);
nor U16551 (N_16551,N_15768,N_15438);
or U16552 (N_16552,N_15307,N_15364);
nand U16553 (N_16553,N_15201,N_15289);
and U16554 (N_16554,N_15583,N_15542);
or U16555 (N_16555,N_15312,N_15635);
nor U16556 (N_16556,N_15334,N_15426);
xnor U16557 (N_16557,N_15219,N_15387);
xor U16558 (N_16558,N_15807,N_15825);
or U16559 (N_16559,N_15867,N_15904);
nor U16560 (N_16560,N_15623,N_15780);
nand U16561 (N_16561,N_15640,N_15289);
or U16562 (N_16562,N_15256,N_15662);
nand U16563 (N_16563,N_15821,N_15552);
nor U16564 (N_16564,N_15262,N_15273);
xnor U16565 (N_16565,N_15537,N_15916);
xnor U16566 (N_16566,N_15876,N_15976);
xor U16567 (N_16567,N_15387,N_15641);
nor U16568 (N_16568,N_15995,N_15789);
nor U16569 (N_16569,N_15243,N_15759);
nor U16570 (N_16570,N_15906,N_15527);
nor U16571 (N_16571,N_15449,N_15561);
and U16572 (N_16572,N_15466,N_15601);
and U16573 (N_16573,N_15932,N_15264);
xor U16574 (N_16574,N_15816,N_15860);
nor U16575 (N_16575,N_15752,N_15611);
nand U16576 (N_16576,N_15860,N_15567);
or U16577 (N_16577,N_15783,N_15655);
or U16578 (N_16578,N_15500,N_15986);
nor U16579 (N_16579,N_15859,N_15648);
xnor U16580 (N_16580,N_15284,N_15356);
or U16581 (N_16581,N_15901,N_15742);
or U16582 (N_16582,N_15961,N_15829);
nor U16583 (N_16583,N_15740,N_15435);
nand U16584 (N_16584,N_15452,N_15479);
nor U16585 (N_16585,N_15658,N_15390);
nand U16586 (N_16586,N_15843,N_15244);
nand U16587 (N_16587,N_15388,N_15303);
and U16588 (N_16588,N_15555,N_15759);
or U16589 (N_16589,N_15591,N_15665);
or U16590 (N_16590,N_15909,N_15436);
and U16591 (N_16591,N_15353,N_15707);
and U16592 (N_16592,N_15429,N_15465);
and U16593 (N_16593,N_15270,N_15423);
nor U16594 (N_16594,N_15448,N_15584);
xor U16595 (N_16595,N_15990,N_15635);
nor U16596 (N_16596,N_15965,N_15752);
and U16597 (N_16597,N_15342,N_15726);
nand U16598 (N_16598,N_15338,N_15769);
and U16599 (N_16599,N_15305,N_15941);
xnor U16600 (N_16600,N_15529,N_15669);
or U16601 (N_16601,N_15541,N_15722);
xor U16602 (N_16602,N_15610,N_15427);
or U16603 (N_16603,N_15605,N_15350);
and U16604 (N_16604,N_15716,N_15633);
or U16605 (N_16605,N_15882,N_15234);
or U16606 (N_16606,N_15564,N_15998);
nand U16607 (N_16607,N_15705,N_15279);
or U16608 (N_16608,N_15821,N_15322);
and U16609 (N_16609,N_15546,N_15613);
xnor U16610 (N_16610,N_15898,N_15217);
or U16611 (N_16611,N_15935,N_15323);
xnor U16612 (N_16612,N_15462,N_15640);
xnor U16613 (N_16613,N_15948,N_15557);
and U16614 (N_16614,N_15890,N_15851);
nor U16615 (N_16615,N_15203,N_15574);
nor U16616 (N_16616,N_15344,N_15326);
xor U16617 (N_16617,N_15895,N_15457);
and U16618 (N_16618,N_15680,N_15731);
nand U16619 (N_16619,N_15291,N_15905);
and U16620 (N_16620,N_15520,N_15899);
xnor U16621 (N_16621,N_15732,N_15214);
xor U16622 (N_16622,N_15509,N_15399);
and U16623 (N_16623,N_15719,N_15490);
or U16624 (N_16624,N_15583,N_15750);
nor U16625 (N_16625,N_15299,N_15802);
nor U16626 (N_16626,N_15817,N_15546);
xor U16627 (N_16627,N_15864,N_15273);
nor U16628 (N_16628,N_15745,N_15276);
or U16629 (N_16629,N_15751,N_15859);
and U16630 (N_16630,N_15760,N_15360);
nand U16631 (N_16631,N_15271,N_15768);
nor U16632 (N_16632,N_15778,N_15556);
xnor U16633 (N_16633,N_15598,N_15851);
nand U16634 (N_16634,N_15584,N_15440);
or U16635 (N_16635,N_15350,N_15379);
nor U16636 (N_16636,N_15805,N_15957);
nor U16637 (N_16637,N_15330,N_15415);
xnor U16638 (N_16638,N_15610,N_15800);
nand U16639 (N_16639,N_15441,N_15964);
and U16640 (N_16640,N_15231,N_15627);
nand U16641 (N_16641,N_15769,N_15418);
nor U16642 (N_16642,N_15439,N_15218);
nand U16643 (N_16643,N_15782,N_15275);
and U16644 (N_16644,N_15943,N_15650);
nand U16645 (N_16645,N_15826,N_15413);
or U16646 (N_16646,N_15908,N_15306);
and U16647 (N_16647,N_15491,N_15900);
and U16648 (N_16648,N_15408,N_15356);
xnor U16649 (N_16649,N_15572,N_15919);
and U16650 (N_16650,N_15864,N_15448);
and U16651 (N_16651,N_15224,N_15542);
or U16652 (N_16652,N_15441,N_15919);
nor U16653 (N_16653,N_15252,N_15524);
xor U16654 (N_16654,N_15722,N_15201);
and U16655 (N_16655,N_15990,N_15653);
nand U16656 (N_16656,N_15389,N_15580);
nor U16657 (N_16657,N_15220,N_15532);
nor U16658 (N_16658,N_15435,N_15542);
nor U16659 (N_16659,N_15890,N_15365);
and U16660 (N_16660,N_15867,N_15900);
or U16661 (N_16661,N_15208,N_15936);
nand U16662 (N_16662,N_15746,N_15925);
or U16663 (N_16663,N_15587,N_15978);
and U16664 (N_16664,N_15705,N_15227);
or U16665 (N_16665,N_15446,N_15301);
or U16666 (N_16666,N_15659,N_15742);
xnor U16667 (N_16667,N_15508,N_15989);
and U16668 (N_16668,N_15211,N_15348);
and U16669 (N_16669,N_15910,N_15706);
or U16670 (N_16670,N_15624,N_15850);
or U16671 (N_16671,N_15546,N_15612);
nand U16672 (N_16672,N_15478,N_15952);
and U16673 (N_16673,N_15236,N_15404);
and U16674 (N_16674,N_15278,N_15568);
xnor U16675 (N_16675,N_15604,N_15988);
and U16676 (N_16676,N_15986,N_15337);
nand U16677 (N_16677,N_15263,N_15447);
nand U16678 (N_16678,N_15715,N_15595);
and U16679 (N_16679,N_15237,N_15541);
or U16680 (N_16680,N_15597,N_15715);
nand U16681 (N_16681,N_15749,N_15963);
nand U16682 (N_16682,N_15744,N_15903);
nor U16683 (N_16683,N_15307,N_15205);
or U16684 (N_16684,N_15214,N_15530);
nor U16685 (N_16685,N_15602,N_15770);
and U16686 (N_16686,N_15246,N_15994);
xor U16687 (N_16687,N_15958,N_15997);
or U16688 (N_16688,N_15256,N_15378);
nand U16689 (N_16689,N_15688,N_15606);
nand U16690 (N_16690,N_15457,N_15917);
nor U16691 (N_16691,N_15809,N_15840);
xor U16692 (N_16692,N_15395,N_15542);
xor U16693 (N_16693,N_15673,N_15711);
nor U16694 (N_16694,N_15757,N_15769);
xor U16695 (N_16695,N_15363,N_15815);
nand U16696 (N_16696,N_15259,N_15942);
nand U16697 (N_16697,N_15390,N_15571);
and U16698 (N_16698,N_15644,N_15541);
and U16699 (N_16699,N_15280,N_15230);
xnor U16700 (N_16700,N_15834,N_15497);
or U16701 (N_16701,N_15886,N_15761);
nand U16702 (N_16702,N_15656,N_15422);
or U16703 (N_16703,N_15294,N_15206);
or U16704 (N_16704,N_15542,N_15820);
or U16705 (N_16705,N_15897,N_15870);
or U16706 (N_16706,N_15606,N_15740);
or U16707 (N_16707,N_15692,N_15963);
xor U16708 (N_16708,N_15870,N_15235);
xor U16709 (N_16709,N_15819,N_15523);
or U16710 (N_16710,N_15986,N_15473);
xnor U16711 (N_16711,N_15482,N_15775);
nor U16712 (N_16712,N_15979,N_15612);
nor U16713 (N_16713,N_15733,N_15654);
nand U16714 (N_16714,N_15491,N_15303);
nand U16715 (N_16715,N_15692,N_15888);
and U16716 (N_16716,N_15258,N_15479);
nor U16717 (N_16717,N_15703,N_15542);
xnor U16718 (N_16718,N_15295,N_15865);
nor U16719 (N_16719,N_15986,N_15984);
or U16720 (N_16720,N_15283,N_15340);
or U16721 (N_16721,N_15948,N_15826);
nor U16722 (N_16722,N_15425,N_15478);
or U16723 (N_16723,N_15324,N_15567);
and U16724 (N_16724,N_15752,N_15710);
nor U16725 (N_16725,N_15977,N_15902);
nor U16726 (N_16726,N_15304,N_15834);
nand U16727 (N_16727,N_15209,N_15983);
xnor U16728 (N_16728,N_15425,N_15798);
nand U16729 (N_16729,N_15646,N_15371);
and U16730 (N_16730,N_15953,N_15322);
or U16731 (N_16731,N_15228,N_15241);
and U16732 (N_16732,N_15767,N_15782);
xnor U16733 (N_16733,N_15303,N_15926);
nand U16734 (N_16734,N_15787,N_15740);
or U16735 (N_16735,N_15317,N_15434);
and U16736 (N_16736,N_15641,N_15446);
nor U16737 (N_16737,N_15747,N_15687);
nand U16738 (N_16738,N_15841,N_15704);
nand U16739 (N_16739,N_15616,N_15752);
nand U16740 (N_16740,N_15451,N_15346);
and U16741 (N_16741,N_15423,N_15356);
xor U16742 (N_16742,N_15270,N_15610);
and U16743 (N_16743,N_15417,N_15240);
nor U16744 (N_16744,N_15564,N_15733);
nand U16745 (N_16745,N_15488,N_15594);
and U16746 (N_16746,N_15667,N_15655);
or U16747 (N_16747,N_15380,N_15837);
nand U16748 (N_16748,N_15798,N_15984);
xor U16749 (N_16749,N_15793,N_15740);
or U16750 (N_16750,N_15959,N_15374);
and U16751 (N_16751,N_15956,N_15845);
xor U16752 (N_16752,N_15933,N_15235);
or U16753 (N_16753,N_15673,N_15248);
nand U16754 (N_16754,N_15616,N_15309);
nor U16755 (N_16755,N_15657,N_15597);
nand U16756 (N_16756,N_15355,N_15577);
nor U16757 (N_16757,N_15750,N_15540);
and U16758 (N_16758,N_15966,N_15701);
or U16759 (N_16759,N_15546,N_15903);
or U16760 (N_16760,N_15444,N_15505);
and U16761 (N_16761,N_15945,N_15488);
nand U16762 (N_16762,N_15437,N_15832);
and U16763 (N_16763,N_15857,N_15585);
nor U16764 (N_16764,N_15576,N_15386);
xor U16765 (N_16765,N_15459,N_15961);
xnor U16766 (N_16766,N_15819,N_15574);
and U16767 (N_16767,N_15621,N_15296);
xnor U16768 (N_16768,N_15602,N_15679);
nand U16769 (N_16769,N_15516,N_15687);
nor U16770 (N_16770,N_15642,N_15857);
xor U16771 (N_16771,N_15597,N_15960);
nor U16772 (N_16772,N_15909,N_15253);
nor U16773 (N_16773,N_15887,N_15698);
nand U16774 (N_16774,N_15937,N_15949);
xor U16775 (N_16775,N_15368,N_15979);
nor U16776 (N_16776,N_15445,N_15977);
and U16777 (N_16777,N_15439,N_15948);
and U16778 (N_16778,N_15541,N_15329);
xnor U16779 (N_16779,N_15569,N_15754);
xor U16780 (N_16780,N_15835,N_15378);
xor U16781 (N_16781,N_15424,N_15596);
xnor U16782 (N_16782,N_15798,N_15532);
nor U16783 (N_16783,N_15890,N_15448);
nor U16784 (N_16784,N_15959,N_15232);
and U16785 (N_16785,N_15639,N_15360);
and U16786 (N_16786,N_15545,N_15670);
nand U16787 (N_16787,N_15869,N_15270);
and U16788 (N_16788,N_15785,N_15349);
or U16789 (N_16789,N_15883,N_15359);
nand U16790 (N_16790,N_15810,N_15864);
xnor U16791 (N_16791,N_15209,N_15884);
nor U16792 (N_16792,N_15693,N_15837);
nor U16793 (N_16793,N_15694,N_15395);
or U16794 (N_16794,N_15629,N_15682);
nand U16795 (N_16795,N_15582,N_15859);
and U16796 (N_16796,N_15460,N_15905);
nand U16797 (N_16797,N_15624,N_15417);
nand U16798 (N_16798,N_15803,N_15269);
xor U16799 (N_16799,N_15858,N_15701);
or U16800 (N_16800,N_16512,N_16329);
or U16801 (N_16801,N_16377,N_16130);
nor U16802 (N_16802,N_16091,N_16068);
and U16803 (N_16803,N_16281,N_16288);
xnor U16804 (N_16804,N_16396,N_16059);
and U16805 (N_16805,N_16678,N_16717);
nand U16806 (N_16806,N_16780,N_16394);
nor U16807 (N_16807,N_16437,N_16346);
nand U16808 (N_16808,N_16737,N_16378);
xnor U16809 (N_16809,N_16334,N_16296);
and U16810 (N_16810,N_16611,N_16392);
nand U16811 (N_16811,N_16553,N_16122);
nand U16812 (N_16812,N_16694,N_16172);
nor U16813 (N_16813,N_16675,N_16715);
and U16814 (N_16814,N_16150,N_16582);
xnor U16815 (N_16815,N_16085,N_16414);
nor U16816 (N_16816,N_16719,N_16411);
xor U16817 (N_16817,N_16337,N_16053);
or U16818 (N_16818,N_16786,N_16208);
and U16819 (N_16819,N_16593,N_16467);
xnor U16820 (N_16820,N_16325,N_16341);
or U16821 (N_16821,N_16503,N_16038);
or U16822 (N_16822,N_16225,N_16400);
nand U16823 (N_16823,N_16307,N_16423);
and U16824 (N_16824,N_16072,N_16375);
and U16825 (N_16825,N_16559,N_16469);
nor U16826 (N_16826,N_16481,N_16086);
nor U16827 (N_16827,N_16441,N_16420);
or U16828 (N_16828,N_16619,N_16327);
xor U16829 (N_16829,N_16209,N_16030);
xnor U16830 (N_16830,N_16162,N_16470);
xor U16831 (N_16831,N_16480,N_16501);
nand U16832 (N_16832,N_16259,N_16710);
nor U16833 (N_16833,N_16718,N_16474);
nor U16834 (N_16834,N_16711,N_16366);
nor U16835 (N_16835,N_16041,N_16065);
and U16836 (N_16836,N_16714,N_16052);
nor U16837 (N_16837,N_16768,N_16021);
xor U16838 (N_16838,N_16279,N_16753);
or U16839 (N_16839,N_16158,N_16426);
or U16840 (N_16840,N_16029,N_16596);
xor U16841 (N_16841,N_16295,N_16624);
or U16842 (N_16842,N_16246,N_16646);
nor U16843 (N_16843,N_16354,N_16569);
xnor U16844 (N_16844,N_16496,N_16459);
or U16845 (N_16845,N_16215,N_16126);
nand U16846 (N_16846,N_16700,N_16516);
or U16847 (N_16847,N_16635,N_16545);
nor U16848 (N_16848,N_16187,N_16287);
nand U16849 (N_16849,N_16724,N_16212);
nor U16850 (N_16850,N_16016,N_16144);
nand U16851 (N_16851,N_16213,N_16040);
and U16852 (N_16852,N_16620,N_16161);
xnor U16853 (N_16853,N_16004,N_16487);
xor U16854 (N_16854,N_16749,N_16704);
and U16855 (N_16855,N_16123,N_16347);
nor U16856 (N_16856,N_16494,N_16538);
nand U16857 (N_16857,N_16644,N_16358);
and U16858 (N_16858,N_16357,N_16703);
xor U16859 (N_16859,N_16743,N_16581);
xnor U16860 (N_16860,N_16433,N_16372);
nand U16861 (N_16861,N_16572,N_16522);
or U16862 (N_16862,N_16070,N_16344);
xnor U16863 (N_16863,N_16319,N_16254);
xnor U16864 (N_16864,N_16078,N_16785);
nor U16865 (N_16865,N_16774,N_16269);
nor U16866 (N_16866,N_16497,N_16034);
xnor U16867 (N_16867,N_16778,N_16701);
or U16868 (N_16868,N_16237,N_16163);
nand U16869 (N_16869,N_16333,N_16626);
nand U16870 (N_16870,N_16140,N_16506);
xnor U16871 (N_16871,N_16783,N_16728);
or U16872 (N_16872,N_16722,N_16128);
nand U16873 (N_16873,N_16322,N_16731);
or U16874 (N_16874,N_16603,N_16077);
nand U16875 (N_16875,N_16132,N_16751);
xnor U16876 (N_16876,N_16772,N_16795);
and U16877 (N_16877,N_16230,N_16349);
nand U16878 (N_16878,N_16178,N_16397);
nand U16879 (N_16879,N_16210,N_16014);
nor U16880 (N_16880,N_16134,N_16020);
or U16881 (N_16881,N_16271,N_16075);
nand U16882 (N_16882,N_16073,N_16174);
nor U16883 (N_16883,N_16159,N_16563);
xnor U16884 (N_16884,N_16777,N_16303);
nor U16885 (N_16885,N_16629,N_16504);
nand U16886 (N_16886,N_16792,N_16054);
or U16887 (N_16887,N_16641,N_16142);
and U16888 (N_16888,N_16660,N_16647);
or U16889 (N_16889,N_16788,N_16642);
or U16890 (N_16890,N_16310,N_16449);
xor U16891 (N_16891,N_16442,N_16661);
xnor U16892 (N_16892,N_16245,N_16022);
or U16893 (N_16893,N_16507,N_16168);
and U16894 (N_16894,N_16148,N_16063);
nand U16895 (N_16895,N_16185,N_16055);
or U16896 (N_16896,N_16203,N_16137);
xnor U16897 (N_16897,N_16520,N_16422);
and U16898 (N_16898,N_16233,N_16005);
and U16899 (N_16899,N_16548,N_16705);
and U16900 (N_16900,N_16676,N_16556);
and U16901 (N_16901,N_16577,N_16668);
xor U16902 (N_16902,N_16402,N_16446);
and U16903 (N_16903,N_16121,N_16336);
nand U16904 (N_16904,N_16305,N_16659);
and U16905 (N_16905,N_16109,N_16623);
xor U16906 (N_16906,N_16525,N_16748);
or U16907 (N_16907,N_16456,N_16529);
nand U16908 (N_16908,N_16193,N_16429);
xor U16909 (N_16909,N_16550,N_16064);
or U16910 (N_16910,N_16238,N_16535);
and U16911 (N_16911,N_16139,N_16765);
nor U16912 (N_16912,N_16561,N_16227);
nor U16913 (N_16913,N_16206,N_16200);
or U16914 (N_16914,N_16046,N_16766);
and U16915 (N_16915,N_16250,N_16087);
xnor U16916 (N_16916,N_16667,N_16406);
or U16917 (N_16917,N_16453,N_16152);
nor U16918 (N_16918,N_16747,N_16679);
xor U16919 (N_16919,N_16428,N_16458);
nor U16920 (N_16920,N_16186,N_16709);
or U16921 (N_16921,N_16368,N_16395);
nor U16922 (N_16922,N_16095,N_16363);
xnor U16923 (N_16923,N_16653,N_16485);
nor U16924 (N_16924,N_16427,N_16663);
or U16925 (N_16925,N_16018,N_16373);
xnor U16926 (N_16926,N_16084,N_16464);
and U16927 (N_16927,N_16094,N_16118);
or U16928 (N_16928,N_16367,N_16199);
nand U16929 (N_16929,N_16670,N_16364);
nand U16930 (N_16930,N_16528,N_16248);
and U16931 (N_16931,N_16403,N_16071);
xor U16932 (N_16932,N_16093,N_16292);
or U16933 (N_16933,N_16081,N_16628);
or U16934 (N_16934,N_16637,N_16650);
nor U16935 (N_16935,N_16686,N_16736);
xnor U16936 (N_16936,N_16472,N_16092);
nand U16937 (N_16937,N_16002,N_16697);
nand U16938 (N_16938,N_16035,N_16583);
or U16939 (N_16939,N_16011,N_16542);
nor U16940 (N_16940,N_16273,N_16147);
nor U16941 (N_16941,N_16601,N_16539);
nor U16942 (N_16942,N_16498,N_16461);
and U16943 (N_16943,N_16184,N_16712);
nand U16944 (N_16944,N_16339,N_16475);
xor U16945 (N_16945,N_16546,N_16745);
or U16946 (N_16946,N_16332,N_16299);
nand U16947 (N_16947,N_16592,N_16784);
or U16948 (N_16948,N_16798,N_16606);
xnor U16949 (N_16949,N_16567,N_16486);
or U16950 (N_16950,N_16404,N_16008);
or U16951 (N_16951,N_16746,N_16110);
or U16952 (N_16952,N_16263,N_16484);
or U16953 (N_16953,N_16666,N_16255);
nand U16954 (N_16954,N_16182,N_16460);
xnor U16955 (N_16955,N_16338,N_16096);
and U16956 (N_16956,N_16773,N_16655);
xnor U16957 (N_16957,N_16621,N_16533);
nor U16958 (N_16958,N_16465,N_16331);
xnor U16959 (N_16959,N_16541,N_16758);
nor U16960 (N_16960,N_16519,N_16074);
and U16961 (N_16961,N_16562,N_16657);
and U16962 (N_16962,N_16775,N_16220);
xor U16963 (N_16963,N_16434,N_16707);
and U16964 (N_16964,N_16380,N_16195);
or U16965 (N_16965,N_16379,N_16612);
and U16966 (N_16966,N_16025,N_16490);
nor U16967 (N_16967,N_16277,N_16170);
nand U16968 (N_16968,N_16324,N_16471);
xor U16969 (N_16969,N_16692,N_16438);
or U16970 (N_16970,N_16216,N_16116);
xor U16971 (N_16971,N_16151,N_16419);
or U16972 (N_16972,N_16610,N_16028);
or U16973 (N_16973,N_16019,N_16106);
nand U16974 (N_16974,N_16725,N_16381);
xnor U16975 (N_16975,N_16293,N_16267);
and U16976 (N_16976,N_16756,N_16547);
nor U16977 (N_16977,N_16721,N_16568);
or U16978 (N_16978,N_16444,N_16352);
nand U16979 (N_16979,N_16431,N_16107);
and U16980 (N_16980,N_16112,N_16156);
and U16981 (N_16981,N_16505,N_16523);
and U16982 (N_16982,N_16636,N_16313);
nand U16983 (N_16983,N_16634,N_16360);
and U16984 (N_16984,N_16256,N_16067);
xor U16985 (N_16985,N_16173,N_16370);
xor U16986 (N_16986,N_16418,N_16177);
or U16987 (N_16987,N_16590,N_16204);
xor U16988 (N_16988,N_16412,N_16732);
nor U16989 (N_16989,N_16359,N_16240);
xor U16990 (N_16990,N_16007,N_16197);
and U16991 (N_16991,N_16565,N_16652);
and U16992 (N_16992,N_16145,N_16039);
xor U16993 (N_16993,N_16278,N_16032);
and U16994 (N_16994,N_16179,N_16735);
xnor U16995 (N_16995,N_16149,N_16082);
or U16996 (N_16996,N_16760,N_16146);
xnor U16997 (N_16997,N_16436,N_16673);
or U16998 (N_16998,N_16708,N_16575);
nand U16999 (N_16999,N_16207,N_16167);
and U17000 (N_17000,N_16473,N_16047);
nor U17001 (N_17001,N_16483,N_16537);
and U17002 (N_17002,N_16176,N_16228);
nand U17003 (N_17003,N_16587,N_16389);
nand U17004 (N_17004,N_16251,N_16617);
xor U17005 (N_17005,N_16764,N_16514);
nand U17006 (N_17006,N_16266,N_16750);
nor U17007 (N_17007,N_16693,N_16742);
and U17008 (N_17008,N_16131,N_16776);
nand U17009 (N_17009,N_16355,N_16320);
or U17010 (N_17010,N_16413,N_16793);
xor U17011 (N_17011,N_16317,N_16574);
and U17012 (N_17012,N_16057,N_16166);
nand U17013 (N_17013,N_16042,N_16727);
xor U17014 (N_17014,N_16120,N_16017);
nand U17015 (N_17015,N_16698,N_16060);
or U17016 (N_17016,N_16045,N_16283);
nor U17017 (N_17017,N_16219,N_16103);
xnor U17018 (N_17018,N_16479,N_16353);
nand U17019 (N_17019,N_16430,N_16416);
nand U17020 (N_17020,N_16382,N_16616);
and U17021 (N_17021,N_16509,N_16124);
nand U17022 (N_17022,N_16244,N_16164);
and U17023 (N_17023,N_16189,N_16602);
xor U17024 (N_17024,N_16242,N_16231);
and U17025 (N_17025,N_16771,N_16405);
or U17026 (N_17026,N_16010,N_16720);
and U17027 (N_17027,N_16393,N_16284);
nand U17028 (N_17028,N_16340,N_16664);
nand U17029 (N_17029,N_16687,N_16543);
or U17030 (N_17030,N_16135,N_16608);
xor U17031 (N_17031,N_16440,N_16689);
nor U17032 (N_17032,N_16221,N_16089);
and U17033 (N_17033,N_16298,N_16468);
xor U17034 (N_17034,N_16114,N_16261);
or U17035 (N_17035,N_16613,N_16680);
nor U17036 (N_17036,N_16262,N_16791);
or U17037 (N_17037,N_16605,N_16730);
and U17038 (N_17038,N_16752,N_16241);
and U17039 (N_17039,N_16155,N_16448);
and U17040 (N_17040,N_16286,N_16665);
nor U17041 (N_17041,N_16560,N_16061);
xnor U17042 (N_17042,N_16729,N_16350);
nand U17043 (N_17043,N_16326,N_16477);
nor U17044 (N_17044,N_16048,N_16175);
or U17045 (N_17045,N_16276,N_16294);
nor U17046 (N_17046,N_16571,N_16734);
and U17047 (N_17047,N_16651,N_16083);
xnor U17048 (N_17048,N_16388,N_16235);
nand U17049 (N_17049,N_16493,N_16723);
nand U17050 (N_17050,N_16138,N_16374);
nand U17051 (N_17051,N_16015,N_16387);
and U17052 (N_17052,N_16180,N_16739);
and U17053 (N_17053,N_16023,N_16598);
nor U17054 (N_17054,N_16043,N_16009);
nor U17055 (N_17055,N_16579,N_16133);
nor U17056 (N_17056,N_16044,N_16125);
nor U17057 (N_17057,N_16615,N_16789);
xor U17058 (N_17058,N_16090,N_16348);
or U17059 (N_17059,N_16645,N_16508);
or U17060 (N_17060,N_16597,N_16643);
nor U17061 (N_17061,N_16631,N_16192);
nor U17062 (N_17062,N_16390,N_16463);
xnor U17063 (N_17063,N_16079,N_16417);
nand U17064 (N_17064,N_16183,N_16169);
nor U17065 (N_17065,N_16455,N_16001);
nand U17066 (N_17066,N_16584,N_16599);
nand U17067 (N_17067,N_16289,N_16051);
or U17068 (N_17068,N_16270,N_16527);
xor U17069 (N_17069,N_16099,N_16767);
nor U17070 (N_17070,N_16532,N_16343);
or U17071 (N_17071,N_16141,N_16614);
or U17072 (N_17072,N_16328,N_16462);
and U17073 (N_17073,N_16301,N_16630);
or U17074 (N_17074,N_16618,N_16511);
and U17075 (N_17075,N_16391,N_16323);
nor U17076 (N_17076,N_16117,N_16491);
nand U17077 (N_17077,N_16321,N_16551);
nor U17078 (N_17078,N_16304,N_16536);
xnor U17079 (N_17079,N_16243,N_16787);
xnor U17080 (N_17080,N_16476,N_16268);
xnor U17081 (N_17081,N_16625,N_16335);
or U17082 (N_17082,N_16101,N_16685);
and U17083 (N_17083,N_16683,N_16451);
or U17084 (N_17084,N_16681,N_16272);
nor U17085 (N_17085,N_16297,N_16309);
xor U17086 (N_17086,N_16253,N_16258);
or U17087 (N_17087,N_16654,N_16252);
nor U17088 (N_17088,N_16257,N_16585);
xnor U17089 (N_17089,N_16576,N_16198);
xnor U17090 (N_17090,N_16489,N_16282);
or U17091 (N_17091,N_16031,N_16500);
nor U17092 (N_17092,N_16695,N_16410);
or U17093 (N_17093,N_16037,N_16672);
nor U17094 (N_17094,N_16308,N_16755);
and U17095 (N_17095,N_16143,N_16564);
nor U17096 (N_17096,N_16351,N_16492);
nand U17097 (N_17097,N_16302,N_16127);
or U17098 (N_17098,N_16058,N_16696);
and U17099 (N_17099,N_16769,N_16761);
xnor U17100 (N_17100,N_16104,N_16384);
or U17101 (N_17101,N_16640,N_16690);
or U17102 (N_17102,N_16555,N_16312);
xor U17103 (N_17103,N_16478,N_16510);
nand U17104 (N_17104,N_16639,N_16076);
nor U17105 (N_17105,N_16799,N_16443);
or U17106 (N_17106,N_16781,N_16797);
and U17107 (N_17107,N_16702,N_16188);
or U17108 (N_17108,N_16757,N_16691);
or U17109 (N_17109,N_16633,N_16656);
and U17110 (N_17110,N_16111,N_16502);
or U17111 (N_17111,N_16521,N_16578);
xnor U17112 (N_17112,N_16214,N_16290);
or U17113 (N_17113,N_16201,N_16674);
nand U17114 (N_17114,N_16100,N_16540);
nand U17115 (N_17115,N_16102,N_16097);
and U17116 (N_17116,N_16196,N_16006);
nor U17117 (N_17117,N_16759,N_16154);
xor U17118 (N_17118,N_16658,N_16108);
or U17119 (N_17119,N_16779,N_16554);
or U17120 (N_17120,N_16026,N_16398);
nand U17121 (N_17121,N_16033,N_16224);
and U17122 (N_17122,N_16062,N_16080);
and U17123 (N_17123,N_16557,N_16371);
nor U17124 (N_17124,N_16306,N_16526);
xor U17125 (N_17125,N_16407,N_16222);
or U17126 (N_17126,N_16762,N_16632);
and U17127 (N_17127,N_16638,N_16447);
nor U17128 (N_17128,N_16024,N_16782);
nor U17129 (N_17129,N_16452,N_16591);
and U17130 (N_17130,N_16239,N_16518);
nor U17131 (N_17131,N_16454,N_16012);
nand U17132 (N_17132,N_16763,N_16191);
and U17133 (N_17133,N_16365,N_16249);
xnor U17134 (N_17134,N_16066,N_16027);
and U17135 (N_17135,N_16165,N_16115);
nor U17136 (N_17136,N_16457,N_16726);
xor U17137 (N_17137,N_16716,N_16265);
nand U17138 (N_17138,N_16361,N_16580);
nand U17139 (N_17139,N_16056,N_16415);
nand U17140 (N_17140,N_16205,N_16558);
nand U17141 (N_17141,N_16383,N_16649);
xor U17142 (N_17142,N_16136,N_16600);
or U17143 (N_17143,N_16594,N_16439);
nor U17144 (N_17144,N_16069,N_16260);
xor U17145 (N_17145,N_16275,N_16408);
and U17146 (N_17146,N_16671,N_16316);
or U17147 (N_17147,N_16385,N_16586);
or U17148 (N_17148,N_16300,N_16223);
and U17149 (N_17149,N_16050,N_16386);
nand U17150 (N_17150,N_16157,N_16345);
or U17151 (N_17151,N_16401,N_16291);
nor U17152 (N_17152,N_16495,N_16744);
or U17153 (N_17153,N_16699,N_16226);
and U17154 (N_17154,N_16247,N_16688);
nor U17155 (N_17155,N_16589,N_16274);
and U17156 (N_17156,N_16342,N_16648);
xnor U17157 (N_17157,N_16524,N_16677);
or U17158 (N_17158,N_16036,N_16544);
nand U17159 (N_17159,N_16662,N_16595);
or U17160 (N_17160,N_16713,N_16549);
nor U17161 (N_17161,N_16211,N_16181);
and U17162 (N_17162,N_16770,N_16217);
and U17163 (N_17163,N_16013,N_16236);
or U17164 (N_17164,N_16000,N_16733);
xnor U17165 (N_17165,N_16609,N_16566);
xnor U17166 (N_17166,N_16432,N_16488);
or U17167 (N_17167,N_16194,N_16604);
nor U17168 (N_17168,N_16513,N_16425);
xor U17169 (N_17169,N_16588,N_16315);
nand U17170 (N_17170,N_16229,N_16129);
xnor U17171 (N_17171,N_16738,N_16482);
xor U17172 (N_17172,N_16285,N_16445);
xor U17173 (N_17173,N_16552,N_16105);
or U17174 (N_17174,N_16098,N_16153);
nand U17175 (N_17175,N_16369,N_16499);
xnor U17176 (N_17176,N_16682,N_16171);
and U17177 (N_17177,N_16421,N_16088);
xnor U17178 (N_17178,N_16534,N_16627);
nor U17179 (N_17179,N_16190,N_16232);
and U17180 (N_17180,N_16466,N_16531);
or U17181 (N_17181,N_16622,N_16049);
nor U17182 (N_17182,N_16790,N_16741);
xor U17183 (N_17183,N_16706,N_16113);
and U17184 (N_17184,N_16003,N_16314);
and U17185 (N_17185,N_16794,N_16280);
nor U17186 (N_17186,N_16218,N_16435);
and U17187 (N_17187,N_16234,N_16515);
or U17188 (N_17188,N_16450,N_16740);
or U17189 (N_17189,N_16424,N_16356);
xnor U17190 (N_17190,N_16376,N_16409);
xnor U17191 (N_17191,N_16669,N_16573);
and U17192 (N_17192,N_16754,N_16160);
nand U17193 (N_17193,N_16362,N_16570);
xnor U17194 (N_17194,N_16796,N_16311);
nand U17195 (N_17195,N_16119,N_16517);
nor U17196 (N_17196,N_16330,N_16530);
xnor U17197 (N_17197,N_16202,N_16399);
or U17198 (N_17198,N_16684,N_16318);
or U17199 (N_17199,N_16264,N_16607);
xor U17200 (N_17200,N_16022,N_16426);
and U17201 (N_17201,N_16684,N_16196);
or U17202 (N_17202,N_16740,N_16000);
nor U17203 (N_17203,N_16266,N_16131);
and U17204 (N_17204,N_16245,N_16555);
or U17205 (N_17205,N_16714,N_16460);
xnor U17206 (N_17206,N_16151,N_16684);
nand U17207 (N_17207,N_16195,N_16703);
and U17208 (N_17208,N_16242,N_16373);
nand U17209 (N_17209,N_16378,N_16153);
or U17210 (N_17210,N_16146,N_16101);
nor U17211 (N_17211,N_16055,N_16732);
xnor U17212 (N_17212,N_16458,N_16173);
or U17213 (N_17213,N_16153,N_16691);
and U17214 (N_17214,N_16731,N_16380);
xor U17215 (N_17215,N_16518,N_16088);
xnor U17216 (N_17216,N_16295,N_16191);
nand U17217 (N_17217,N_16490,N_16024);
or U17218 (N_17218,N_16085,N_16350);
and U17219 (N_17219,N_16602,N_16661);
nor U17220 (N_17220,N_16291,N_16574);
xnor U17221 (N_17221,N_16214,N_16048);
or U17222 (N_17222,N_16459,N_16121);
or U17223 (N_17223,N_16417,N_16285);
and U17224 (N_17224,N_16472,N_16112);
and U17225 (N_17225,N_16304,N_16499);
nand U17226 (N_17226,N_16453,N_16454);
xnor U17227 (N_17227,N_16028,N_16645);
nand U17228 (N_17228,N_16679,N_16530);
xnor U17229 (N_17229,N_16620,N_16348);
and U17230 (N_17230,N_16212,N_16230);
nand U17231 (N_17231,N_16193,N_16172);
nand U17232 (N_17232,N_16170,N_16440);
xnor U17233 (N_17233,N_16172,N_16779);
nand U17234 (N_17234,N_16460,N_16185);
nor U17235 (N_17235,N_16339,N_16550);
nand U17236 (N_17236,N_16341,N_16367);
or U17237 (N_17237,N_16066,N_16048);
or U17238 (N_17238,N_16174,N_16371);
xor U17239 (N_17239,N_16154,N_16290);
or U17240 (N_17240,N_16277,N_16537);
and U17241 (N_17241,N_16533,N_16260);
or U17242 (N_17242,N_16288,N_16023);
and U17243 (N_17243,N_16367,N_16054);
or U17244 (N_17244,N_16479,N_16003);
nor U17245 (N_17245,N_16442,N_16604);
and U17246 (N_17246,N_16358,N_16135);
and U17247 (N_17247,N_16705,N_16331);
nand U17248 (N_17248,N_16241,N_16768);
or U17249 (N_17249,N_16605,N_16244);
or U17250 (N_17250,N_16305,N_16500);
xor U17251 (N_17251,N_16243,N_16655);
or U17252 (N_17252,N_16205,N_16193);
nand U17253 (N_17253,N_16436,N_16578);
nor U17254 (N_17254,N_16336,N_16234);
nand U17255 (N_17255,N_16503,N_16005);
xor U17256 (N_17256,N_16384,N_16200);
nand U17257 (N_17257,N_16489,N_16750);
nand U17258 (N_17258,N_16070,N_16265);
or U17259 (N_17259,N_16006,N_16210);
or U17260 (N_17260,N_16711,N_16643);
and U17261 (N_17261,N_16421,N_16444);
nand U17262 (N_17262,N_16794,N_16027);
xnor U17263 (N_17263,N_16025,N_16782);
nor U17264 (N_17264,N_16168,N_16461);
or U17265 (N_17265,N_16482,N_16287);
xor U17266 (N_17266,N_16532,N_16144);
nor U17267 (N_17267,N_16174,N_16091);
nand U17268 (N_17268,N_16635,N_16464);
xnor U17269 (N_17269,N_16658,N_16552);
nand U17270 (N_17270,N_16011,N_16792);
nand U17271 (N_17271,N_16596,N_16398);
or U17272 (N_17272,N_16465,N_16753);
xor U17273 (N_17273,N_16156,N_16148);
nor U17274 (N_17274,N_16493,N_16766);
xnor U17275 (N_17275,N_16534,N_16173);
nor U17276 (N_17276,N_16353,N_16567);
xnor U17277 (N_17277,N_16316,N_16116);
xor U17278 (N_17278,N_16765,N_16776);
and U17279 (N_17279,N_16623,N_16609);
xor U17280 (N_17280,N_16059,N_16462);
xnor U17281 (N_17281,N_16418,N_16448);
nand U17282 (N_17282,N_16728,N_16241);
xnor U17283 (N_17283,N_16036,N_16552);
xnor U17284 (N_17284,N_16267,N_16123);
nor U17285 (N_17285,N_16504,N_16125);
xor U17286 (N_17286,N_16306,N_16425);
nor U17287 (N_17287,N_16781,N_16074);
and U17288 (N_17288,N_16697,N_16470);
or U17289 (N_17289,N_16695,N_16540);
nand U17290 (N_17290,N_16487,N_16345);
xnor U17291 (N_17291,N_16542,N_16145);
nor U17292 (N_17292,N_16599,N_16062);
nand U17293 (N_17293,N_16205,N_16506);
and U17294 (N_17294,N_16766,N_16775);
and U17295 (N_17295,N_16507,N_16171);
nand U17296 (N_17296,N_16752,N_16613);
and U17297 (N_17297,N_16227,N_16378);
nor U17298 (N_17298,N_16729,N_16498);
or U17299 (N_17299,N_16299,N_16020);
and U17300 (N_17300,N_16231,N_16394);
nand U17301 (N_17301,N_16019,N_16646);
nor U17302 (N_17302,N_16485,N_16128);
xnor U17303 (N_17303,N_16638,N_16519);
xnor U17304 (N_17304,N_16345,N_16210);
or U17305 (N_17305,N_16118,N_16750);
and U17306 (N_17306,N_16565,N_16466);
and U17307 (N_17307,N_16071,N_16167);
or U17308 (N_17308,N_16686,N_16584);
and U17309 (N_17309,N_16594,N_16613);
xor U17310 (N_17310,N_16289,N_16385);
or U17311 (N_17311,N_16656,N_16126);
nor U17312 (N_17312,N_16748,N_16766);
nand U17313 (N_17313,N_16131,N_16143);
and U17314 (N_17314,N_16374,N_16334);
nor U17315 (N_17315,N_16410,N_16483);
and U17316 (N_17316,N_16688,N_16412);
nor U17317 (N_17317,N_16089,N_16741);
nor U17318 (N_17318,N_16044,N_16634);
xnor U17319 (N_17319,N_16626,N_16661);
xnor U17320 (N_17320,N_16744,N_16155);
nor U17321 (N_17321,N_16298,N_16179);
nand U17322 (N_17322,N_16532,N_16151);
nand U17323 (N_17323,N_16714,N_16202);
and U17324 (N_17324,N_16312,N_16761);
nor U17325 (N_17325,N_16217,N_16154);
nor U17326 (N_17326,N_16312,N_16585);
nand U17327 (N_17327,N_16177,N_16613);
xnor U17328 (N_17328,N_16528,N_16570);
nand U17329 (N_17329,N_16422,N_16725);
xnor U17330 (N_17330,N_16273,N_16284);
nand U17331 (N_17331,N_16130,N_16704);
nand U17332 (N_17332,N_16049,N_16072);
and U17333 (N_17333,N_16401,N_16451);
and U17334 (N_17334,N_16007,N_16349);
nor U17335 (N_17335,N_16370,N_16321);
nor U17336 (N_17336,N_16047,N_16688);
or U17337 (N_17337,N_16204,N_16018);
nor U17338 (N_17338,N_16150,N_16600);
xnor U17339 (N_17339,N_16736,N_16753);
xnor U17340 (N_17340,N_16695,N_16350);
xnor U17341 (N_17341,N_16781,N_16520);
and U17342 (N_17342,N_16354,N_16488);
or U17343 (N_17343,N_16467,N_16763);
and U17344 (N_17344,N_16183,N_16248);
nor U17345 (N_17345,N_16462,N_16256);
or U17346 (N_17346,N_16359,N_16245);
and U17347 (N_17347,N_16765,N_16663);
nand U17348 (N_17348,N_16230,N_16344);
xor U17349 (N_17349,N_16611,N_16597);
nor U17350 (N_17350,N_16189,N_16693);
or U17351 (N_17351,N_16382,N_16128);
xor U17352 (N_17352,N_16793,N_16223);
or U17353 (N_17353,N_16418,N_16790);
xnor U17354 (N_17354,N_16612,N_16667);
and U17355 (N_17355,N_16477,N_16043);
xor U17356 (N_17356,N_16669,N_16523);
xor U17357 (N_17357,N_16622,N_16353);
nor U17358 (N_17358,N_16100,N_16233);
nor U17359 (N_17359,N_16414,N_16322);
nor U17360 (N_17360,N_16521,N_16621);
nor U17361 (N_17361,N_16317,N_16131);
nor U17362 (N_17362,N_16388,N_16616);
nor U17363 (N_17363,N_16373,N_16333);
nand U17364 (N_17364,N_16155,N_16709);
and U17365 (N_17365,N_16105,N_16449);
nor U17366 (N_17366,N_16136,N_16784);
nor U17367 (N_17367,N_16194,N_16542);
or U17368 (N_17368,N_16499,N_16659);
nand U17369 (N_17369,N_16541,N_16498);
nor U17370 (N_17370,N_16507,N_16337);
xnor U17371 (N_17371,N_16211,N_16174);
nor U17372 (N_17372,N_16548,N_16210);
nand U17373 (N_17373,N_16339,N_16707);
nor U17374 (N_17374,N_16781,N_16585);
nor U17375 (N_17375,N_16294,N_16450);
nor U17376 (N_17376,N_16437,N_16461);
xor U17377 (N_17377,N_16161,N_16215);
and U17378 (N_17378,N_16223,N_16306);
and U17379 (N_17379,N_16625,N_16431);
and U17380 (N_17380,N_16602,N_16237);
or U17381 (N_17381,N_16788,N_16402);
and U17382 (N_17382,N_16790,N_16500);
xnor U17383 (N_17383,N_16331,N_16030);
and U17384 (N_17384,N_16510,N_16564);
or U17385 (N_17385,N_16717,N_16406);
and U17386 (N_17386,N_16563,N_16376);
xnor U17387 (N_17387,N_16409,N_16298);
and U17388 (N_17388,N_16638,N_16036);
or U17389 (N_17389,N_16163,N_16449);
nand U17390 (N_17390,N_16376,N_16535);
nor U17391 (N_17391,N_16268,N_16591);
nand U17392 (N_17392,N_16395,N_16686);
xnor U17393 (N_17393,N_16436,N_16050);
and U17394 (N_17394,N_16314,N_16248);
or U17395 (N_17395,N_16541,N_16638);
or U17396 (N_17396,N_16506,N_16168);
nor U17397 (N_17397,N_16797,N_16379);
xnor U17398 (N_17398,N_16142,N_16526);
nor U17399 (N_17399,N_16134,N_16759);
or U17400 (N_17400,N_16510,N_16505);
nor U17401 (N_17401,N_16619,N_16620);
nand U17402 (N_17402,N_16724,N_16316);
or U17403 (N_17403,N_16254,N_16198);
nor U17404 (N_17404,N_16306,N_16016);
and U17405 (N_17405,N_16241,N_16463);
and U17406 (N_17406,N_16317,N_16418);
nand U17407 (N_17407,N_16362,N_16131);
and U17408 (N_17408,N_16713,N_16758);
and U17409 (N_17409,N_16192,N_16357);
nor U17410 (N_17410,N_16701,N_16521);
xnor U17411 (N_17411,N_16453,N_16161);
xor U17412 (N_17412,N_16497,N_16088);
xor U17413 (N_17413,N_16019,N_16368);
and U17414 (N_17414,N_16161,N_16741);
or U17415 (N_17415,N_16788,N_16764);
nor U17416 (N_17416,N_16330,N_16305);
nand U17417 (N_17417,N_16708,N_16426);
or U17418 (N_17418,N_16086,N_16623);
nand U17419 (N_17419,N_16033,N_16436);
nand U17420 (N_17420,N_16296,N_16555);
xnor U17421 (N_17421,N_16308,N_16009);
and U17422 (N_17422,N_16216,N_16391);
nor U17423 (N_17423,N_16667,N_16724);
nand U17424 (N_17424,N_16577,N_16333);
nand U17425 (N_17425,N_16406,N_16498);
nand U17426 (N_17426,N_16392,N_16119);
nand U17427 (N_17427,N_16665,N_16102);
or U17428 (N_17428,N_16097,N_16134);
nor U17429 (N_17429,N_16735,N_16074);
or U17430 (N_17430,N_16401,N_16072);
nor U17431 (N_17431,N_16400,N_16776);
xnor U17432 (N_17432,N_16492,N_16513);
and U17433 (N_17433,N_16756,N_16317);
and U17434 (N_17434,N_16586,N_16431);
nor U17435 (N_17435,N_16626,N_16665);
nand U17436 (N_17436,N_16002,N_16141);
or U17437 (N_17437,N_16068,N_16674);
nand U17438 (N_17438,N_16467,N_16580);
nor U17439 (N_17439,N_16146,N_16757);
or U17440 (N_17440,N_16396,N_16748);
nor U17441 (N_17441,N_16523,N_16326);
nand U17442 (N_17442,N_16759,N_16213);
nor U17443 (N_17443,N_16726,N_16740);
and U17444 (N_17444,N_16244,N_16279);
and U17445 (N_17445,N_16778,N_16317);
nand U17446 (N_17446,N_16299,N_16375);
or U17447 (N_17447,N_16595,N_16398);
xor U17448 (N_17448,N_16404,N_16038);
nand U17449 (N_17449,N_16485,N_16667);
nor U17450 (N_17450,N_16542,N_16144);
nand U17451 (N_17451,N_16292,N_16759);
xnor U17452 (N_17452,N_16675,N_16311);
and U17453 (N_17453,N_16075,N_16309);
nor U17454 (N_17454,N_16321,N_16558);
and U17455 (N_17455,N_16066,N_16355);
and U17456 (N_17456,N_16626,N_16157);
nor U17457 (N_17457,N_16145,N_16694);
and U17458 (N_17458,N_16735,N_16283);
and U17459 (N_17459,N_16784,N_16297);
xnor U17460 (N_17460,N_16421,N_16471);
or U17461 (N_17461,N_16619,N_16422);
nor U17462 (N_17462,N_16471,N_16759);
or U17463 (N_17463,N_16062,N_16137);
or U17464 (N_17464,N_16584,N_16490);
nand U17465 (N_17465,N_16284,N_16498);
nor U17466 (N_17466,N_16085,N_16221);
nand U17467 (N_17467,N_16497,N_16436);
nor U17468 (N_17468,N_16377,N_16537);
xnor U17469 (N_17469,N_16410,N_16677);
nor U17470 (N_17470,N_16090,N_16346);
nand U17471 (N_17471,N_16297,N_16480);
nand U17472 (N_17472,N_16549,N_16349);
nand U17473 (N_17473,N_16001,N_16428);
and U17474 (N_17474,N_16154,N_16232);
and U17475 (N_17475,N_16091,N_16482);
nand U17476 (N_17476,N_16784,N_16390);
nor U17477 (N_17477,N_16534,N_16086);
nor U17478 (N_17478,N_16503,N_16097);
nand U17479 (N_17479,N_16725,N_16196);
or U17480 (N_17480,N_16238,N_16127);
xor U17481 (N_17481,N_16051,N_16476);
nor U17482 (N_17482,N_16689,N_16493);
xnor U17483 (N_17483,N_16559,N_16252);
nand U17484 (N_17484,N_16642,N_16394);
nor U17485 (N_17485,N_16323,N_16701);
and U17486 (N_17486,N_16096,N_16689);
nor U17487 (N_17487,N_16241,N_16344);
and U17488 (N_17488,N_16583,N_16292);
or U17489 (N_17489,N_16245,N_16069);
xor U17490 (N_17490,N_16653,N_16437);
nor U17491 (N_17491,N_16177,N_16564);
and U17492 (N_17492,N_16011,N_16020);
xor U17493 (N_17493,N_16296,N_16792);
and U17494 (N_17494,N_16230,N_16303);
and U17495 (N_17495,N_16713,N_16591);
and U17496 (N_17496,N_16756,N_16568);
or U17497 (N_17497,N_16499,N_16407);
nand U17498 (N_17498,N_16194,N_16102);
or U17499 (N_17499,N_16713,N_16176);
and U17500 (N_17500,N_16495,N_16074);
nor U17501 (N_17501,N_16690,N_16596);
nor U17502 (N_17502,N_16173,N_16222);
nor U17503 (N_17503,N_16314,N_16500);
or U17504 (N_17504,N_16550,N_16706);
nand U17505 (N_17505,N_16508,N_16130);
or U17506 (N_17506,N_16032,N_16539);
xnor U17507 (N_17507,N_16798,N_16518);
and U17508 (N_17508,N_16482,N_16251);
or U17509 (N_17509,N_16670,N_16638);
nor U17510 (N_17510,N_16273,N_16755);
or U17511 (N_17511,N_16417,N_16520);
nand U17512 (N_17512,N_16274,N_16508);
nand U17513 (N_17513,N_16239,N_16436);
xor U17514 (N_17514,N_16461,N_16100);
nor U17515 (N_17515,N_16046,N_16038);
nor U17516 (N_17516,N_16546,N_16478);
nand U17517 (N_17517,N_16190,N_16498);
xor U17518 (N_17518,N_16362,N_16464);
or U17519 (N_17519,N_16635,N_16071);
or U17520 (N_17520,N_16552,N_16643);
or U17521 (N_17521,N_16402,N_16662);
nand U17522 (N_17522,N_16497,N_16014);
xnor U17523 (N_17523,N_16338,N_16506);
nor U17524 (N_17524,N_16377,N_16558);
xor U17525 (N_17525,N_16610,N_16589);
xor U17526 (N_17526,N_16322,N_16083);
and U17527 (N_17527,N_16034,N_16639);
nor U17528 (N_17528,N_16781,N_16416);
nand U17529 (N_17529,N_16337,N_16610);
nand U17530 (N_17530,N_16314,N_16299);
nand U17531 (N_17531,N_16128,N_16517);
xnor U17532 (N_17532,N_16452,N_16517);
nor U17533 (N_17533,N_16315,N_16545);
xnor U17534 (N_17534,N_16493,N_16522);
or U17535 (N_17535,N_16533,N_16608);
or U17536 (N_17536,N_16380,N_16399);
or U17537 (N_17537,N_16648,N_16362);
or U17538 (N_17538,N_16744,N_16482);
xor U17539 (N_17539,N_16323,N_16444);
nor U17540 (N_17540,N_16357,N_16193);
nor U17541 (N_17541,N_16129,N_16243);
and U17542 (N_17542,N_16080,N_16611);
and U17543 (N_17543,N_16229,N_16598);
or U17544 (N_17544,N_16043,N_16001);
and U17545 (N_17545,N_16103,N_16400);
and U17546 (N_17546,N_16581,N_16098);
or U17547 (N_17547,N_16209,N_16124);
and U17548 (N_17548,N_16352,N_16407);
or U17549 (N_17549,N_16464,N_16779);
or U17550 (N_17550,N_16671,N_16321);
nor U17551 (N_17551,N_16584,N_16064);
xnor U17552 (N_17552,N_16556,N_16654);
and U17553 (N_17553,N_16317,N_16450);
and U17554 (N_17554,N_16340,N_16242);
nand U17555 (N_17555,N_16345,N_16545);
and U17556 (N_17556,N_16210,N_16674);
nor U17557 (N_17557,N_16050,N_16413);
nor U17558 (N_17558,N_16592,N_16382);
nand U17559 (N_17559,N_16364,N_16173);
nor U17560 (N_17560,N_16731,N_16290);
or U17561 (N_17561,N_16091,N_16268);
xor U17562 (N_17562,N_16036,N_16453);
or U17563 (N_17563,N_16354,N_16404);
or U17564 (N_17564,N_16325,N_16363);
nand U17565 (N_17565,N_16561,N_16263);
xor U17566 (N_17566,N_16446,N_16392);
and U17567 (N_17567,N_16590,N_16114);
nand U17568 (N_17568,N_16190,N_16341);
nor U17569 (N_17569,N_16252,N_16489);
nor U17570 (N_17570,N_16604,N_16483);
or U17571 (N_17571,N_16603,N_16512);
xnor U17572 (N_17572,N_16633,N_16304);
xor U17573 (N_17573,N_16774,N_16154);
and U17574 (N_17574,N_16344,N_16154);
nor U17575 (N_17575,N_16482,N_16463);
nand U17576 (N_17576,N_16359,N_16761);
xnor U17577 (N_17577,N_16738,N_16508);
xor U17578 (N_17578,N_16599,N_16381);
nor U17579 (N_17579,N_16514,N_16328);
nand U17580 (N_17580,N_16325,N_16114);
xor U17581 (N_17581,N_16757,N_16644);
nand U17582 (N_17582,N_16156,N_16036);
and U17583 (N_17583,N_16486,N_16082);
or U17584 (N_17584,N_16672,N_16074);
xnor U17585 (N_17585,N_16097,N_16180);
nand U17586 (N_17586,N_16396,N_16696);
or U17587 (N_17587,N_16572,N_16265);
nand U17588 (N_17588,N_16798,N_16624);
and U17589 (N_17589,N_16383,N_16182);
nor U17590 (N_17590,N_16627,N_16536);
or U17591 (N_17591,N_16603,N_16165);
nand U17592 (N_17592,N_16368,N_16156);
nor U17593 (N_17593,N_16139,N_16065);
nand U17594 (N_17594,N_16766,N_16617);
or U17595 (N_17595,N_16158,N_16753);
nor U17596 (N_17596,N_16326,N_16706);
or U17597 (N_17597,N_16586,N_16514);
xor U17598 (N_17598,N_16555,N_16437);
nor U17599 (N_17599,N_16484,N_16624);
nor U17600 (N_17600,N_17330,N_17599);
or U17601 (N_17601,N_17211,N_17402);
nor U17602 (N_17602,N_17391,N_17546);
nor U17603 (N_17603,N_17499,N_17334);
xor U17604 (N_17604,N_17532,N_17295);
or U17605 (N_17605,N_17501,N_17516);
nor U17606 (N_17606,N_17449,N_17368);
and U17607 (N_17607,N_16826,N_17482);
or U17608 (N_17608,N_16935,N_17387);
xnor U17609 (N_17609,N_16854,N_16967);
or U17610 (N_17610,N_17196,N_16890);
nor U17611 (N_17611,N_17404,N_17182);
and U17612 (N_17612,N_17207,N_17531);
nand U17613 (N_17613,N_17254,N_16914);
or U17614 (N_17614,N_17432,N_17091);
nand U17615 (N_17615,N_16859,N_17525);
and U17616 (N_17616,N_17517,N_16867);
xor U17617 (N_17617,N_16877,N_17587);
and U17618 (N_17618,N_17265,N_17255);
nand U17619 (N_17619,N_17022,N_17215);
xor U17620 (N_17620,N_17104,N_17421);
and U17621 (N_17621,N_17348,N_17306);
xnor U17622 (N_17622,N_17400,N_17084);
nor U17623 (N_17623,N_17377,N_16902);
or U17624 (N_17624,N_17561,N_16960);
nor U17625 (N_17625,N_17540,N_17403);
nand U17626 (N_17626,N_16883,N_17229);
or U17627 (N_17627,N_17174,N_16983);
or U17628 (N_17628,N_16884,N_17522);
nand U17629 (N_17629,N_17333,N_17293);
and U17630 (N_17630,N_17103,N_17023);
xnor U17631 (N_17631,N_17280,N_17381);
nor U17632 (N_17632,N_16855,N_17566);
xnor U17633 (N_17633,N_17050,N_17508);
nand U17634 (N_17634,N_17453,N_16905);
nand U17635 (N_17635,N_17437,N_17030);
and U17636 (N_17636,N_17000,N_16963);
nand U17637 (N_17637,N_17596,N_17063);
xor U17638 (N_17638,N_17016,N_16866);
xnor U17639 (N_17639,N_17111,N_17493);
and U17640 (N_17640,N_16993,N_16956);
nor U17641 (N_17641,N_17494,N_17485);
nor U17642 (N_17642,N_17362,N_16808);
nand U17643 (N_17643,N_17171,N_17355);
nor U17644 (N_17644,N_17331,N_16813);
or U17645 (N_17645,N_17383,N_17337);
and U17646 (N_17646,N_17052,N_17228);
nor U17647 (N_17647,N_17079,N_17169);
nor U17648 (N_17648,N_17269,N_16822);
nor U17649 (N_17649,N_17314,N_17461);
nand U17650 (N_17650,N_17071,N_17184);
xnor U17651 (N_17651,N_17267,N_16996);
nand U17652 (N_17652,N_17183,N_17148);
nor U17653 (N_17653,N_17131,N_17231);
xor U17654 (N_17654,N_17488,N_17342);
nor U17655 (N_17655,N_16838,N_17492);
and U17656 (N_17656,N_17373,N_17570);
nor U17657 (N_17657,N_17093,N_17251);
xnor U17658 (N_17658,N_17443,N_17298);
nor U17659 (N_17659,N_17080,N_16940);
nand U17660 (N_17660,N_17436,N_17445);
and U17661 (N_17661,N_17451,N_17354);
or U17662 (N_17662,N_17285,N_17475);
xor U17663 (N_17663,N_17308,N_17160);
or U17664 (N_17664,N_17555,N_17035);
xor U17665 (N_17665,N_16958,N_17536);
nand U17666 (N_17666,N_17370,N_17512);
nand U17667 (N_17667,N_17535,N_17116);
xnor U17668 (N_17668,N_17300,N_17018);
or U17669 (N_17669,N_16954,N_17081);
xor U17670 (N_17670,N_17025,N_17444);
xor U17671 (N_17671,N_17442,N_17464);
and U17672 (N_17672,N_17162,N_17122);
nor U17673 (N_17673,N_17548,N_16819);
and U17674 (N_17674,N_17441,N_16906);
or U17675 (N_17675,N_17054,N_17090);
nand U17676 (N_17676,N_17135,N_16887);
nor U17677 (N_17677,N_17019,N_17114);
nand U17678 (N_17678,N_17328,N_17112);
xnor U17679 (N_17679,N_17012,N_17191);
nand U17680 (N_17680,N_17427,N_17176);
nand U17681 (N_17681,N_17218,N_17256);
and U17682 (N_17682,N_17438,N_17219);
and U17683 (N_17683,N_17246,N_17047);
and U17684 (N_17684,N_17205,N_16942);
and U17685 (N_17685,N_17467,N_17089);
xor U17686 (N_17686,N_16959,N_16865);
nand U17687 (N_17687,N_17459,N_17353);
nand U17688 (N_17688,N_17152,N_16835);
or U17689 (N_17689,N_17010,N_17157);
xnor U17690 (N_17690,N_17545,N_17398);
and U17691 (N_17691,N_16880,N_17263);
xor U17692 (N_17692,N_17120,N_17504);
nand U17693 (N_17693,N_17552,N_17472);
and U17694 (N_17694,N_17502,N_17509);
xor U17695 (N_17695,N_17027,N_16896);
nor U17696 (N_17696,N_16961,N_17194);
xor U17697 (N_17697,N_17107,N_17544);
xnor U17698 (N_17698,N_17235,N_17189);
xnor U17699 (N_17699,N_17573,N_16840);
or U17700 (N_17700,N_17351,N_17412);
nor U17701 (N_17701,N_17560,N_17070);
and U17702 (N_17702,N_17335,N_16926);
nand U17703 (N_17703,N_17015,N_17542);
nand U17704 (N_17704,N_17514,N_17369);
or U17705 (N_17705,N_16848,N_17311);
nor U17706 (N_17706,N_17274,N_17138);
nand U17707 (N_17707,N_17455,N_17374);
and U17708 (N_17708,N_17217,N_17266);
and U17709 (N_17709,N_16917,N_17558);
or U17710 (N_17710,N_17466,N_17420);
nand U17711 (N_17711,N_16941,N_17533);
and U17712 (N_17712,N_17193,N_17230);
nor U17713 (N_17713,N_17302,N_17159);
and U17714 (N_17714,N_17271,N_17195);
xnor U17715 (N_17715,N_17320,N_17585);
or U17716 (N_17716,N_16949,N_17396);
and U17717 (N_17717,N_17134,N_17476);
and U17718 (N_17718,N_16984,N_17495);
and U17719 (N_17719,N_16804,N_17234);
or U17720 (N_17720,N_16805,N_17456);
nor U17721 (N_17721,N_17097,N_16831);
and U17722 (N_17722,N_17260,N_17580);
nor U17723 (N_17723,N_16997,N_16807);
xor U17724 (N_17724,N_16806,N_17074);
xor U17725 (N_17725,N_17500,N_17017);
nor U17726 (N_17726,N_17382,N_16853);
nand U17727 (N_17727,N_17101,N_17061);
and U17728 (N_17728,N_17393,N_16885);
or U17729 (N_17729,N_17066,N_17105);
nor U17730 (N_17730,N_17471,N_17137);
or U17731 (N_17731,N_16882,N_16825);
nand U17732 (N_17732,N_16974,N_16879);
and U17733 (N_17733,N_16888,N_17305);
or U17734 (N_17734,N_16829,N_17004);
nor U17735 (N_17735,N_17244,N_17198);
xnor U17736 (N_17736,N_16828,N_17239);
xor U17737 (N_17737,N_17237,N_17425);
nand U17738 (N_17738,N_16889,N_17575);
or U17739 (N_17739,N_17329,N_17513);
nor U17740 (N_17740,N_16876,N_17245);
or U17741 (N_17741,N_17496,N_17128);
xor U17742 (N_17742,N_17123,N_16923);
and U17743 (N_17743,N_17188,N_17262);
and U17744 (N_17744,N_16843,N_17503);
or U17745 (N_17745,N_17537,N_17474);
xor U17746 (N_17746,N_17336,N_17319);
nor U17747 (N_17747,N_17040,N_17143);
or U17748 (N_17748,N_16928,N_17339);
nand U17749 (N_17749,N_17096,N_17209);
nor U17750 (N_17750,N_16856,N_16982);
nor U17751 (N_17751,N_16952,N_16987);
nand U17752 (N_17752,N_17357,N_17149);
or U17753 (N_17753,N_17340,N_17223);
nor U17754 (N_17754,N_17416,N_17457);
and U17755 (N_17755,N_17323,N_17236);
xnor U17756 (N_17756,N_17133,N_17327);
xor U17757 (N_17757,N_16950,N_16851);
and U17758 (N_17758,N_17272,N_17042);
xnor U17759 (N_17759,N_17121,N_16936);
nand U17760 (N_17760,N_17257,N_16810);
nand U17761 (N_17761,N_17439,N_17129);
xnor U17762 (N_17762,N_16979,N_17233);
or U17763 (N_17763,N_17507,N_17011);
nand U17764 (N_17764,N_17581,N_16852);
nand U17765 (N_17765,N_17592,N_16837);
and U17766 (N_17766,N_17534,N_16820);
nand U17767 (N_17767,N_17549,N_17250);
nor U17768 (N_17768,N_17118,N_17434);
nor U17769 (N_17769,N_16850,N_17275);
xnor U17770 (N_17770,N_17059,N_17277);
or U17771 (N_17771,N_17173,N_16868);
nor U17772 (N_17772,N_17290,N_17110);
nand U17773 (N_17773,N_17530,N_17470);
and U17774 (N_17774,N_17083,N_17248);
nor U17775 (N_17775,N_17344,N_16846);
or U17776 (N_17776,N_17478,N_16869);
and U17777 (N_17777,N_17276,N_17069);
xor U17778 (N_17778,N_17591,N_17031);
and U17779 (N_17779,N_17384,N_16832);
nand U17780 (N_17780,N_17043,N_16989);
xnor U17781 (N_17781,N_16934,N_16910);
xnor U17782 (N_17782,N_16915,N_17154);
nand U17783 (N_17783,N_17589,N_17164);
nor U17784 (N_17784,N_16976,N_17547);
and U17785 (N_17785,N_17124,N_17597);
xnor U17786 (N_17786,N_17115,N_16857);
or U17787 (N_17787,N_16924,N_17395);
nand U17788 (N_17788,N_17568,N_17372);
nand U17789 (N_17789,N_16921,N_17569);
or U17790 (N_17790,N_16842,N_17565);
nand U17791 (N_17791,N_17579,N_17551);
nor U17792 (N_17792,N_17008,N_17498);
and U17793 (N_17793,N_17379,N_17058);
nor U17794 (N_17794,N_16931,N_17187);
nor U17795 (N_17795,N_17013,N_17422);
or U17796 (N_17796,N_17224,N_16815);
and U17797 (N_17797,N_17125,N_17153);
nor U17798 (N_17798,N_17521,N_16817);
nor U17799 (N_17799,N_16834,N_16980);
xnor U17800 (N_17800,N_17594,N_16891);
nor U17801 (N_17801,N_17132,N_16985);
nand U17802 (N_17802,N_16938,N_16860);
and U17803 (N_17803,N_17297,N_17009);
nor U17804 (N_17804,N_16816,N_17588);
xnor U17805 (N_17805,N_17360,N_17206);
nand U17806 (N_17806,N_16998,N_17212);
nand U17807 (N_17807,N_16920,N_16955);
xnor U17808 (N_17808,N_16863,N_16886);
nor U17809 (N_17809,N_17316,N_17158);
xor U17810 (N_17810,N_16939,N_17102);
or U17811 (N_17811,N_17086,N_17242);
nand U17812 (N_17812,N_17287,N_17034);
and U17813 (N_17813,N_16841,N_17106);
and U17814 (N_17814,N_17026,N_16830);
and U17815 (N_17815,N_17414,N_17462);
nand U17816 (N_17816,N_17192,N_17450);
nor U17817 (N_17817,N_17454,N_17307);
xnor U17818 (N_17818,N_17388,N_17527);
or U17819 (N_17819,N_17350,N_17036);
or U17820 (N_17820,N_16811,N_17163);
xor U17821 (N_17821,N_17510,N_16968);
nand U17822 (N_17822,N_17538,N_16893);
nand U17823 (N_17823,N_16870,N_16922);
or U17824 (N_17824,N_17448,N_17590);
xor U17825 (N_17825,N_17068,N_17076);
nand U17826 (N_17826,N_17473,N_17098);
nor U17827 (N_17827,N_16861,N_17289);
nor U17828 (N_17828,N_17072,N_16969);
xnor U17829 (N_17829,N_17214,N_16972);
nor U17830 (N_17830,N_16803,N_17127);
nand U17831 (N_17831,N_16849,N_17238);
nand U17832 (N_17832,N_17078,N_17279);
and U17833 (N_17833,N_17151,N_16873);
or U17834 (N_17834,N_17550,N_17428);
or U17835 (N_17835,N_17175,N_17543);
nor U17836 (N_17836,N_17346,N_16973);
xnor U17837 (N_17837,N_16981,N_17429);
nand U17838 (N_17838,N_17073,N_17301);
nand U17839 (N_17839,N_17168,N_16809);
or U17840 (N_17840,N_17186,N_17363);
and U17841 (N_17841,N_17366,N_17062);
and U17842 (N_17842,N_17584,N_17465);
xnor U17843 (N_17843,N_17576,N_17142);
nor U17844 (N_17844,N_17578,N_17430);
xnor U17845 (N_17845,N_16971,N_17447);
nand U17846 (N_17846,N_16933,N_16953);
and U17847 (N_17847,N_17556,N_17491);
nor U17848 (N_17848,N_17284,N_16944);
and U17849 (N_17849,N_17469,N_17413);
xor U17850 (N_17850,N_16839,N_17526);
nor U17851 (N_17851,N_17225,N_17264);
nor U17852 (N_17852,N_16878,N_17356);
nand U17853 (N_17853,N_17281,N_17593);
xor U17854 (N_17854,N_17166,N_17213);
xnor U17855 (N_17855,N_17216,N_17002);
xnor U17856 (N_17856,N_16992,N_17178);
xnor U17857 (N_17857,N_16948,N_17410);
nor U17858 (N_17858,N_17349,N_17147);
xnor U17859 (N_17859,N_17347,N_17199);
and U17860 (N_17860,N_16881,N_17497);
and U17861 (N_17861,N_17222,N_17001);
and U17862 (N_17862,N_17253,N_16871);
xnor U17863 (N_17863,N_17386,N_17324);
or U17864 (N_17864,N_17446,N_17270);
nand U17865 (N_17865,N_17088,N_17595);
nand U17866 (N_17866,N_16892,N_17232);
and U17867 (N_17867,N_17479,N_16945);
nand U17868 (N_17868,N_17037,N_16916);
nand U17869 (N_17869,N_17506,N_17180);
or U17870 (N_17870,N_17202,N_17486);
or U17871 (N_17871,N_16929,N_16991);
and U17872 (N_17872,N_17358,N_16918);
nand U17873 (N_17873,N_17060,N_17511);
and U17874 (N_17874,N_17338,N_17304);
nand U17875 (N_17875,N_17051,N_17144);
nand U17876 (N_17876,N_17409,N_17559);
and U17877 (N_17877,N_17039,N_17095);
or U17878 (N_17878,N_17468,N_17415);
nor U17879 (N_17879,N_17582,N_16966);
or U17880 (N_17880,N_17385,N_17577);
nor U17881 (N_17881,N_16800,N_16964);
and U17882 (N_17882,N_17371,N_16965);
nor U17883 (N_17883,N_17041,N_17487);
nand U17884 (N_17884,N_17252,N_16932);
or U17885 (N_17885,N_17433,N_16951);
nor U17886 (N_17886,N_17563,N_16927);
or U17887 (N_17887,N_16970,N_17463);
nand U17888 (N_17888,N_17156,N_17064);
or U17889 (N_17889,N_17028,N_16912);
and U17890 (N_17890,N_17136,N_17208);
nor U17891 (N_17891,N_16911,N_17249);
nor U17892 (N_17892,N_17389,N_16901);
and U17893 (N_17893,N_17099,N_17426);
xnor U17894 (N_17894,N_17583,N_16946);
xnor U17895 (N_17895,N_17553,N_16899);
xnor U17896 (N_17896,N_17049,N_17325);
and U17897 (N_17897,N_17085,N_17489);
nor U17898 (N_17898,N_17317,N_17005);
nand U17899 (N_17899,N_17318,N_17571);
nor U17900 (N_17900,N_16986,N_16827);
or U17901 (N_17901,N_17155,N_16988);
nor U17902 (N_17902,N_16845,N_17247);
nor U17903 (N_17903,N_17460,N_17378);
nor U17904 (N_17904,N_16994,N_17201);
and U17905 (N_17905,N_17100,N_17161);
and U17906 (N_17906,N_17481,N_17203);
nand U17907 (N_17907,N_17227,N_17313);
xor U17908 (N_17908,N_16904,N_17431);
nand U17909 (N_17909,N_17179,N_17087);
xnor U17910 (N_17910,N_16864,N_17299);
nor U17911 (N_17911,N_17539,N_17390);
nand U17912 (N_17912,N_16937,N_17165);
nand U17913 (N_17913,N_17519,N_17190);
nand U17914 (N_17914,N_17044,N_17480);
nand U17915 (N_17915,N_17524,N_17452);
and U17916 (N_17916,N_16812,N_16824);
xor U17917 (N_17917,N_17490,N_16862);
and U17918 (N_17918,N_17045,N_17021);
nor U17919 (N_17919,N_17020,N_17177);
and U17920 (N_17920,N_17401,N_17367);
nor U17921 (N_17921,N_17418,N_17146);
nor U17922 (N_17922,N_16957,N_16909);
xor U17923 (N_17923,N_17520,N_17528);
xor U17924 (N_17924,N_16919,N_17278);
nand U17925 (N_17925,N_17484,N_17417);
xnor U17926 (N_17926,N_17518,N_17408);
xnor U17927 (N_17927,N_17108,N_17424);
nor U17928 (N_17928,N_17140,N_16999);
or U17929 (N_17929,N_17240,N_17322);
nand U17930 (N_17930,N_16947,N_17282);
or U17931 (N_17931,N_17291,N_17523);
nor U17932 (N_17932,N_17321,N_16990);
nor U17933 (N_17933,N_17315,N_17440);
and U17934 (N_17934,N_17376,N_17567);
xnor U17935 (N_17935,N_17332,N_17014);
or U17936 (N_17936,N_17296,N_17113);
or U17937 (N_17937,N_16925,N_17032);
xnor U17938 (N_17938,N_17141,N_17483);
and U17939 (N_17939,N_17204,N_16894);
xnor U17940 (N_17940,N_17109,N_17259);
and U17941 (N_17941,N_17185,N_17399);
xnor U17942 (N_17942,N_17341,N_16875);
xnor U17943 (N_17943,N_16814,N_16821);
nor U17944 (N_17944,N_17172,N_16930);
nand U17945 (N_17945,N_16801,N_17343);
xor U17946 (N_17946,N_16844,N_17130);
nor U17947 (N_17947,N_16943,N_17094);
xor U17948 (N_17948,N_17065,N_16975);
nand U17949 (N_17949,N_17529,N_17303);
nand U17950 (N_17950,N_17411,N_16900);
or U17951 (N_17951,N_17574,N_17226);
nand U17952 (N_17952,N_17562,N_17458);
xnor U17953 (N_17953,N_17392,N_17394);
or U17954 (N_17954,N_16823,N_16898);
xnor U17955 (N_17955,N_16978,N_16858);
or U17956 (N_17956,N_16903,N_16872);
or U17957 (N_17957,N_16833,N_17024);
nand U17958 (N_17958,N_17055,N_17048);
nand U17959 (N_17959,N_17067,N_17294);
nor U17960 (N_17960,N_16907,N_16977);
and U17961 (N_17961,N_17405,N_17273);
and U17962 (N_17962,N_17380,N_17029);
and U17963 (N_17963,N_17477,N_17326);
or U17964 (N_17964,N_17352,N_17210);
or U17965 (N_17965,N_17364,N_16802);
xnor U17966 (N_17966,N_16897,N_16818);
nor U17967 (N_17967,N_17221,N_17310);
nand U17968 (N_17968,N_17359,N_17292);
nand U17969 (N_17969,N_17312,N_17309);
nor U17970 (N_17970,N_17361,N_17419);
nor U17971 (N_17971,N_17288,N_17003);
nand U17972 (N_17972,N_16847,N_17407);
xnor U17973 (N_17973,N_17139,N_17598);
nand U17974 (N_17974,N_17268,N_17119);
nand U17975 (N_17975,N_17243,N_17375);
or U17976 (N_17976,N_17586,N_17077);
and U17977 (N_17977,N_17197,N_17082);
xor U17978 (N_17978,N_17006,N_17033);
xnor U17979 (N_17979,N_17200,N_17007);
or U17980 (N_17980,N_17150,N_17170);
and U17981 (N_17981,N_17261,N_17167);
or U17982 (N_17982,N_17345,N_17557);
or U17983 (N_17983,N_17145,N_17572);
nand U17984 (N_17984,N_17397,N_17515);
or U17985 (N_17985,N_17286,N_17406);
nor U17986 (N_17986,N_17423,N_17046);
and U17987 (N_17987,N_17258,N_17075);
nor U17988 (N_17988,N_17541,N_17554);
nand U17989 (N_17989,N_17057,N_17117);
nand U17990 (N_17990,N_17053,N_16995);
nand U17991 (N_17991,N_16913,N_16874);
and U17992 (N_17992,N_17241,N_17365);
or U17993 (N_17993,N_16895,N_17220);
or U17994 (N_17994,N_17038,N_17126);
and U17995 (N_17995,N_17564,N_16836);
nor U17996 (N_17996,N_16908,N_17435);
and U17997 (N_17997,N_16962,N_17056);
nor U17998 (N_17998,N_17181,N_17505);
and U17999 (N_17999,N_17092,N_17283);
xnor U18000 (N_18000,N_17593,N_17213);
xor U18001 (N_18001,N_17194,N_16923);
nand U18002 (N_18002,N_17540,N_17066);
and U18003 (N_18003,N_17187,N_17374);
nand U18004 (N_18004,N_17342,N_17000);
nor U18005 (N_18005,N_17568,N_17330);
nor U18006 (N_18006,N_17478,N_17116);
or U18007 (N_18007,N_17050,N_17006);
xor U18008 (N_18008,N_17296,N_17203);
or U18009 (N_18009,N_17570,N_17006);
and U18010 (N_18010,N_17105,N_16925);
and U18011 (N_18011,N_17277,N_17236);
nor U18012 (N_18012,N_17033,N_16934);
or U18013 (N_18013,N_16874,N_17495);
nor U18014 (N_18014,N_16829,N_17365);
or U18015 (N_18015,N_17348,N_17178);
and U18016 (N_18016,N_16834,N_16890);
nor U18017 (N_18017,N_16851,N_17111);
xor U18018 (N_18018,N_17477,N_17535);
and U18019 (N_18019,N_17232,N_17446);
and U18020 (N_18020,N_17201,N_17485);
nand U18021 (N_18021,N_17256,N_17588);
or U18022 (N_18022,N_17228,N_17422);
nor U18023 (N_18023,N_17147,N_17064);
and U18024 (N_18024,N_17158,N_17075);
xnor U18025 (N_18025,N_16960,N_16937);
nor U18026 (N_18026,N_17327,N_16967);
or U18027 (N_18027,N_16983,N_17477);
and U18028 (N_18028,N_17347,N_17072);
nand U18029 (N_18029,N_17422,N_17264);
xnor U18030 (N_18030,N_17218,N_17026);
xnor U18031 (N_18031,N_17213,N_16997);
xnor U18032 (N_18032,N_17118,N_17581);
or U18033 (N_18033,N_16863,N_17543);
xor U18034 (N_18034,N_17207,N_17307);
xor U18035 (N_18035,N_16978,N_17230);
and U18036 (N_18036,N_17336,N_17174);
xnor U18037 (N_18037,N_17585,N_17060);
or U18038 (N_18038,N_17337,N_17308);
nand U18039 (N_18039,N_17242,N_17583);
nor U18040 (N_18040,N_16805,N_16861);
nand U18041 (N_18041,N_17299,N_16870);
xnor U18042 (N_18042,N_17344,N_16829);
nand U18043 (N_18043,N_17579,N_17563);
and U18044 (N_18044,N_17472,N_17599);
and U18045 (N_18045,N_16995,N_17489);
xor U18046 (N_18046,N_17331,N_16817);
xor U18047 (N_18047,N_17586,N_17083);
or U18048 (N_18048,N_16895,N_17345);
xor U18049 (N_18049,N_16980,N_17467);
or U18050 (N_18050,N_16912,N_17017);
and U18051 (N_18051,N_17181,N_17026);
xor U18052 (N_18052,N_16887,N_17379);
xor U18053 (N_18053,N_17217,N_17162);
xnor U18054 (N_18054,N_17536,N_17433);
or U18055 (N_18055,N_17063,N_16912);
nor U18056 (N_18056,N_17479,N_16952);
nor U18057 (N_18057,N_17146,N_17450);
nor U18058 (N_18058,N_17326,N_16911);
or U18059 (N_18059,N_17259,N_17305);
or U18060 (N_18060,N_17443,N_17503);
xor U18061 (N_18061,N_17342,N_17159);
nor U18062 (N_18062,N_17168,N_17595);
nor U18063 (N_18063,N_17409,N_17539);
xnor U18064 (N_18064,N_17354,N_17234);
nor U18065 (N_18065,N_17545,N_16903);
and U18066 (N_18066,N_17445,N_17475);
nor U18067 (N_18067,N_16974,N_17185);
nand U18068 (N_18068,N_17578,N_17496);
nor U18069 (N_18069,N_16957,N_16942);
nand U18070 (N_18070,N_17469,N_17378);
and U18071 (N_18071,N_17336,N_17441);
or U18072 (N_18072,N_17575,N_16998);
nor U18073 (N_18073,N_17150,N_17400);
and U18074 (N_18074,N_17317,N_16989);
or U18075 (N_18075,N_17061,N_17087);
nand U18076 (N_18076,N_16988,N_16892);
nor U18077 (N_18077,N_17451,N_16903);
and U18078 (N_18078,N_17577,N_16843);
nand U18079 (N_18079,N_17458,N_17354);
or U18080 (N_18080,N_17464,N_17422);
nand U18081 (N_18081,N_17213,N_16826);
and U18082 (N_18082,N_16980,N_17434);
nor U18083 (N_18083,N_17094,N_16833);
or U18084 (N_18084,N_17553,N_16853);
nand U18085 (N_18085,N_16818,N_16814);
xnor U18086 (N_18086,N_17165,N_17238);
and U18087 (N_18087,N_17063,N_17391);
or U18088 (N_18088,N_17382,N_17271);
and U18089 (N_18089,N_17020,N_17085);
and U18090 (N_18090,N_16857,N_17060);
and U18091 (N_18091,N_16865,N_17115);
nand U18092 (N_18092,N_17037,N_16984);
xnor U18093 (N_18093,N_16886,N_17190);
nand U18094 (N_18094,N_16968,N_16934);
nand U18095 (N_18095,N_17218,N_17397);
nor U18096 (N_18096,N_17474,N_16920);
nand U18097 (N_18097,N_16848,N_16920);
nor U18098 (N_18098,N_17343,N_17360);
nor U18099 (N_18099,N_16924,N_16978);
xnor U18100 (N_18100,N_17430,N_17234);
xor U18101 (N_18101,N_17575,N_17219);
xnor U18102 (N_18102,N_17273,N_17258);
and U18103 (N_18103,N_16926,N_17080);
nand U18104 (N_18104,N_17202,N_17596);
and U18105 (N_18105,N_17476,N_16882);
nand U18106 (N_18106,N_17399,N_16936);
nand U18107 (N_18107,N_17420,N_17183);
and U18108 (N_18108,N_17427,N_16857);
and U18109 (N_18109,N_17421,N_17221);
nand U18110 (N_18110,N_17109,N_17247);
or U18111 (N_18111,N_17446,N_17463);
or U18112 (N_18112,N_17324,N_17408);
and U18113 (N_18113,N_16926,N_16877);
and U18114 (N_18114,N_17434,N_17073);
xnor U18115 (N_18115,N_16815,N_17302);
or U18116 (N_18116,N_17161,N_17056);
nand U18117 (N_18117,N_17425,N_16968);
nor U18118 (N_18118,N_17162,N_16932);
nand U18119 (N_18119,N_17373,N_17351);
or U18120 (N_18120,N_16964,N_17556);
and U18121 (N_18121,N_16908,N_17184);
nor U18122 (N_18122,N_17311,N_17310);
or U18123 (N_18123,N_17352,N_16849);
nor U18124 (N_18124,N_17349,N_16880);
nor U18125 (N_18125,N_17031,N_17058);
nand U18126 (N_18126,N_17388,N_17083);
xor U18127 (N_18127,N_17322,N_17147);
nor U18128 (N_18128,N_17116,N_17208);
or U18129 (N_18129,N_16869,N_17488);
nor U18130 (N_18130,N_17179,N_17383);
xor U18131 (N_18131,N_17478,N_17105);
and U18132 (N_18132,N_17088,N_17089);
and U18133 (N_18133,N_17337,N_17164);
xor U18134 (N_18134,N_17146,N_16950);
and U18135 (N_18135,N_16900,N_16860);
nand U18136 (N_18136,N_16838,N_17317);
xor U18137 (N_18137,N_17074,N_16969);
and U18138 (N_18138,N_17270,N_16940);
and U18139 (N_18139,N_17099,N_17032);
and U18140 (N_18140,N_17109,N_17138);
nand U18141 (N_18141,N_17098,N_17122);
nand U18142 (N_18142,N_17342,N_17545);
or U18143 (N_18143,N_16944,N_17555);
and U18144 (N_18144,N_17335,N_17002);
nand U18145 (N_18145,N_17171,N_17280);
or U18146 (N_18146,N_17161,N_16827);
xnor U18147 (N_18147,N_17227,N_17112);
and U18148 (N_18148,N_17537,N_17410);
or U18149 (N_18149,N_17553,N_17417);
xor U18150 (N_18150,N_17229,N_16991);
nand U18151 (N_18151,N_17498,N_17339);
nand U18152 (N_18152,N_17390,N_17568);
nand U18153 (N_18153,N_16812,N_16895);
xnor U18154 (N_18154,N_17436,N_17389);
or U18155 (N_18155,N_17478,N_17569);
xor U18156 (N_18156,N_17594,N_17092);
xnor U18157 (N_18157,N_16861,N_17412);
nand U18158 (N_18158,N_17219,N_16950);
nand U18159 (N_18159,N_17518,N_16898);
nand U18160 (N_18160,N_17057,N_17157);
xor U18161 (N_18161,N_17477,N_17100);
or U18162 (N_18162,N_16914,N_17007);
or U18163 (N_18163,N_17361,N_17187);
and U18164 (N_18164,N_16951,N_17496);
nor U18165 (N_18165,N_17382,N_17204);
and U18166 (N_18166,N_17497,N_17106);
nor U18167 (N_18167,N_16971,N_17110);
nand U18168 (N_18168,N_17534,N_17107);
or U18169 (N_18169,N_16887,N_17052);
nand U18170 (N_18170,N_17233,N_17104);
or U18171 (N_18171,N_17158,N_16957);
xnor U18172 (N_18172,N_17410,N_17384);
nand U18173 (N_18173,N_17229,N_17177);
and U18174 (N_18174,N_17225,N_16934);
xor U18175 (N_18175,N_17044,N_17170);
nand U18176 (N_18176,N_17584,N_17437);
nor U18177 (N_18177,N_17358,N_16889);
nor U18178 (N_18178,N_17583,N_16892);
nand U18179 (N_18179,N_17093,N_17036);
nor U18180 (N_18180,N_17289,N_17192);
nand U18181 (N_18181,N_16897,N_17269);
xnor U18182 (N_18182,N_17245,N_17114);
or U18183 (N_18183,N_17084,N_17378);
and U18184 (N_18184,N_17122,N_17356);
xor U18185 (N_18185,N_17331,N_16961);
and U18186 (N_18186,N_16881,N_17507);
nand U18187 (N_18187,N_16822,N_17582);
xor U18188 (N_18188,N_16953,N_17205);
and U18189 (N_18189,N_17351,N_17152);
xnor U18190 (N_18190,N_17080,N_17599);
and U18191 (N_18191,N_16988,N_16854);
nand U18192 (N_18192,N_16851,N_17120);
nor U18193 (N_18193,N_17030,N_17365);
nand U18194 (N_18194,N_17109,N_17173);
nand U18195 (N_18195,N_16944,N_16851);
or U18196 (N_18196,N_16805,N_17443);
nor U18197 (N_18197,N_16986,N_16809);
and U18198 (N_18198,N_17286,N_17525);
xor U18199 (N_18199,N_17594,N_17325);
xor U18200 (N_18200,N_17004,N_16825);
nand U18201 (N_18201,N_17419,N_16896);
and U18202 (N_18202,N_17150,N_17452);
nor U18203 (N_18203,N_16976,N_17317);
nor U18204 (N_18204,N_17581,N_17339);
xnor U18205 (N_18205,N_17368,N_17037);
nor U18206 (N_18206,N_17006,N_16814);
xor U18207 (N_18207,N_17091,N_16837);
nor U18208 (N_18208,N_17473,N_16946);
nor U18209 (N_18209,N_17317,N_16856);
and U18210 (N_18210,N_17573,N_16989);
and U18211 (N_18211,N_17051,N_17513);
and U18212 (N_18212,N_17237,N_17491);
xor U18213 (N_18213,N_16851,N_17491);
nor U18214 (N_18214,N_17194,N_17584);
nor U18215 (N_18215,N_17197,N_17463);
nor U18216 (N_18216,N_17113,N_17024);
xor U18217 (N_18217,N_17376,N_17288);
nor U18218 (N_18218,N_17033,N_17233);
nand U18219 (N_18219,N_16940,N_16894);
and U18220 (N_18220,N_16865,N_17509);
nor U18221 (N_18221,N_17384,N_17539);
nor U18222 (N_18222,N_17422,N_17408);
or U18223 (N_18223,N_17518,N_17244);
xor U18224 (N_18224,N_17030,N_17423);
nand U18225 (N_18225,N_17396,N_17587);
nor U18226 (N_18226,N_17344,N_16967);
and U18227 (N_18227,N_17511,N_17149);
xnor U18228 (N_18228,N_17248,N_17523);
or U18229 (N_18229,N_16918,N_17211);
or U18230 (N_18230,N_17295,N_17188);
or U18231 (N_18231,N_17192,N_17037);
nor U18232 (N_18232,N_17433,N_17263);
nor U18233 (N_18233,N_16990,N_17236);
xor U18234 (N_18234,N_17387,N_17364);
nor U18235 (N_18235,N_17488,N_17487);
and U18236 (N_18236,N_17521,N_17500);
xor U18237 (N_18237,N_17431,N_17406);
or U18238 (N_18238,N_16961,N_16809);
nor U18239 (N_18239,N_17339,N_17489);
or U18240 (N_18240,N_16927,N_17559);
and U18241 (N_18241,N_17427,N_17426);
and U18242 (N_18242,N_17364,N_17527);
and U18243 (N_18243,N_16954,N_17176);
or U18244 (N_18244,N_17182,N_16940);
nor U18245 (N_18245,N_17534,N_17565);
nand U18246 (N_18246,N_17224,N_17245);
and U18247 (N_18247,N_16995,N_17299);
nor U18248 (N_18248,N_17081,N_16807);
nor U18249 (N_18249,N_17297,N_17557);
and U18250 (N_18250,N_17128,N_16909);
nor U18251 (N_18251,N_17165,N_17469);
nand U18252 (N_18252,N_17218,N_17389);
nand U18253 (N_18253,N_17384,N_17421);
and U18254 (N_18254,N_17001,N_17237);
nand U18255 (N_18255,N_17176,N_17488);
nor U18256 (N_18256,N_16897,N_17566);
nand U18257 (N_18257,N_17168,N_17180);
or U18258 (N_18258,N_17587,N_17152);
nor U18259 (N_18259,N_17058,N_17241);
nor U18260 (N_18260,N_16858,N_17136);
or U18261 (N_18261,N_17589,N_17051);
nor U18262 (N_18262,N_16961,N_17574);
or U18263 (N_18263,N_16910,N_17093);
nor U18264 (N_18264,N_17576,N_17583);
or U18265 (N_18265,N_17166,N_17087);
nand U18266 (N_18266,N_17459,N_16954);
nand U18267 (N_18267,N_17344,N_17498);
or U18268 (N_18268,N_17138,N_17040);
nor U18269 (N_18269,N_17036,N_17047);
and U18270 (N_18270,N_17285,N_17580);
nand U18271 (N_18271,N_16910,N_16804);
and U18272 (N_18272,N_17193,N_17059);
nand U18273 (N_18273,N_17149,N_16945);
xnor U18274 (N_18274,N_17207,N_17313);
nand U18275 (N_18275,N_17191,N_17490);
and U18276 (N_18276,N_17585,N_17364);
and U18277 (N_18277,N_17592,N_17444);
and U18278 (N_18278,N_17589,N_17462);
and U18279 (N_18279,N_16947,N_17233);
and U18280 (N_18280,N_17092,N_17434);
xnor U18281 (N_18281,N_17307,N_17008);
and U18282 (N_18282,N_16868,N_17251);
nand U18283 (N_18283,N_16871,N_17431);
or U18284 (N_18284,N_16921,N_16997);
nand U18285 (N_18285,N_17051,N_17274);
nor U18286 (N_18286,N_17457,N_17074);
or U18287 (N_18287,N_17589,N_17305);
and U18288 (N_18288,N_16923,N_16928);
or U18289 (N_18289,N_17390,N_17317);
and U18290 (N_18290,N_17072,N_17506);
or U18291 (N_18291,N_16924,N_17156);
nand U18292 (N_18292,N_17241,N_17469);
nor U18293 (N_18293,N_17262,N_17108);
or U18294 (N_18294,N_17548,N_17493);
nor U18295 (N_18295,N_17456,N_17291);
nor U18296 (N_18296,N_17044,N_17563);
nand U18297 (N_18297,N_17434,N_17385);
or U18298 (N_18298,N_17361,N_17234);
nor U18299 (N_18299,N_17239,N_17149);
xnor U18300 (N_18300,N_17186,N_17367);
nand U18301 (N_18301,N_16997,N_17087);
nor U18302 (N_18302,N_16811,N_17146);
nand U18303 (N_18303,N_16860,N_17145);
xor U18304 (N_18304,N_17413,N_17180);
nor U18305 (N_18305,N_17351,N_17286);
xor U18306 (N_18306,N_16990,N_17133);
or U18307 (N_18307,N_17120,N_17282);
or U18308 (N_18308,N_17220,N_17251);
nand U18309 (N_18309,N_17369,N_17144);
xor U18310 (N_18310,N_17019,N_17470);
and U18311 (N_18311,N_17068,N_16822);
nor U18312 (N_18312,N_17513,N_17379);
nand U18313 (N_18313,N_17112,N_16879);
and U18314 (N_18314,N_17256,N_17573);
nand U18315 (N_18315,N_17583,N_17086);
nor U18316 (N_18316,N_17176,N_17198);
xor U18317 (N_18317,N_17358,N_17521);
nor U18318 (N_18318,N_17483,N_17575);
nand U18319 (N_18319,N_17338,N_17589);
xor U18320 (N_18320,N_17192,N_17142);
or U18321 (N_18321,N_17557,N_16980);
or U18322 (N_18322,N_17351,N_17279);
nor U18323 (N_18323,N_17388,N_17488);
or U18324 (N_18324,N_17242,N_17422);
nand U18325 (N_18325,N_17553,N_17208);
nor U18326 (N_18326,N_17436,N_17418);
nand U18327 (N_18327,N_17262,N_17547);
and U18328 (N_18328,N_17297,N_17521);
nand U18329 (N_18329,N_17435,N_17083);
or U18330 (N_18330,N_16804,N_16813);
and U18331 (N_18331,N_17467,N_17295);
or U18332 (N_18332,N_16857,N_17380);
xnor U18333 (N_18333,N_17341,N_16960);
or U18334 (N_18334,N_17358,N_17373);
xor U18335 (N_18335,N_16862,N_16955);
nor U18336 (N_18336,N_17519,N_17222);
or U18337 (N_18337,N_17233,N_17064);
and U18338 (N_18338,N_17488,N_17011);
nand U18339 (N_18339,N_16819,N_16802);
xnor U18340 (N_18340,N_17529,N_17168);
and U18341 (N_18341,N_17064,N_17505);
xor U18342 (N_18342,N_17346,N_17261);
xnor U18343 (N_18343,N_17212,N_17081);
and U18344 (N_18344,N_17053,N_17039);
and U18345 (N_18345,N_16992,N_17269);
xor U18346 (N_18346,N_16996,N_17036);
xnor U18347 (N_18347,N_17240,N_17453);
nor U18348 (N_18348,N_16918,N_17250);
nor U18349 (N_18349,N_16827,N_17456);
or U18350 (N_18350,N_17598,N_17356);
and U18351 (N_18351,N_17129,N_16951);
and U18352 (N_18352,N_16996,N_17276);
nor U18353 (N_18353,N_17446,N_17558);
nor U18354 (N_18354,N_16987,N_17123);
and U18355 (N_18355,N_17371,N_17444);
nor U18356 (N_18356,N_17131,N_16925);
nand U18357 (N_18357,N_17493,N_17281);
nand U18358 (N_18358,N_17072,N_16949);
and U18359 (N_18359,N_17063,N_17434);
or U18360 (N_18360,N_17353,N_17095);
xnor U18361 (N_18361,N_16903,N_17495);
and U18362 (N_18362,N_17495,N_17564);
or U18363 (N_18363,N_17491,N_17363);
nand U18364 (N_18364,N_17492,N_17348);
nand U18365 (N_18365,N_16808,N_17413);
and U18366 (N_18366,N_17185,N_17523);
xnor U18367 (N_18367,N_17080,N_16803);
and U18368 (N_18368,N_17560,N_16834);
nor U18369 (N_18369,N_17342,N_17110);
nand U18370 (N_18370,N_16839,N_17028);
and U18371 (N_18371,N_16871,N_17260);
nor U18372 (N_18372,N_17527,N_16978);
nor U18373 (N_18373,N_17301,N_16805);
nor U18374 (N_18374,N_17132,N_17549);
nand U18375 (N_18375,N_16979,N_17168);
xor U18376 (N_18376,N_17111,N_17419);
and U18377 (N_18377,N_17071,N_16819);
and U18378 (N_18378,N_17107,N_16872);
xor U18379 (N_18379,N_16877,N_17267);
and U18380 (N_18380,N_16853,N_17454);
or U18381 (N_18381,N_17406,N_17370);
nand U18382 (N_18382,N_17279,N_17027);
and U18383 (N_18383,N_16962,N_17460);
and U18384 (N_18384,N_17217,N_17355);
and U18385 (N_18385,N_17096,N_17504);
xor U18386 (N_18386,N_17290,N_16883);
nand U18387 (N_18387,N_17263,N_17419);
nor U18388 (N_18388,N_17177,N_17524);
nand U18389 (N_18389,N_17008,N_17537);
and U18390 (N_18390,N_17181,N_16976);
or U18391 (N_18391,N_17241,N_16806);
nand U18392 (N_18392,N_16938,N_16886);
nor U18393 (N_18393,N_17232,N_17053);
nand U18394 (N_18394,N_16885,N_16962);
xnor U18395 (N_18395,N_17235,N_17068);
xnor U18396 (N_18396,N_17519,N_17572);
xor U18397 (N_18397,N_17162,N_16880);
or U18398 (N_18398,N_16895,N_17172);
nand U18399 (N_18399,N_17032,N_17557);
or U18400 (N_18400,N_17976,N_17824);
and U18401 (N_18401,N_18308,N_17940);
xnor U18402 (N_18402,N_17879,N_18182);
or U18403 (N_18403,N_17967,N_17860);
nand U18404 (N_18404,N_18183,N_18144);
or U18405 (N_18405,N_18022,N_17856);
nor U18406 (N_18406,N_18113,N_17882);
nand U18407 (N_18407,N_18006,N_18373);
xnor U18408 (N_18408,N_17754,N_17947);
nor U18409 (N_18409,N_17886,N_17796);
nor U18410 (N_18410,N_17659,N_18002);
nor U18411 (N_18411,N_18205,N_18389);
or U18412 (N_18412,N_18048,N_17934);
nor U18413 (N_18413,N_18289,N_18141);
and U18414 (N_18414,N_17871,N_18210);
nand U18415 (N_18415,N_18296,N_18080);
and U18416 (N_18416,N_17952,N_17630);
and U18417 (N_18417,N_18189,N_18235);
nand U18418 (N_18418,N_17609,N_18122);
nor U18419 (N_18419,N_18324,N_18281);
nand U18420 (N_18420,N_17811,N_17668);
and U18421 (N_18421,N_18150,N_17992);
nand U18422 (N_18422,N_17677,N_18225);
xor U18423 (N_18423,N_17939,N_17624);
xnor U18424 (N_18424,N_17950,N_17721);
and U18425 (N_18425,N_18360,N_17617);
or U18426 (N_18426,N_17697,N_18128);
nand U18427 (N_18427,N_17971,N_18058);
nand U18428 (N_18428,N_17828,N_17794);
nor U18429 (N_18429,N_18019,N_18218);
and U18430 (N_18430,N_18114,N_18032);
or U18431 (N_18431,N_18226,N_17623);
xor U18432 (N_18432,N_18186,N_18378);
xnor U18433 (N_18433,N_18143,N_18387);
nor U18434 (N_18434,N_17881,N_17672);
nor U18435 (N_18435,N_17854,N_18326);
xnor U18436 (N_18436,N_18224,N_18335);
and U18437 (N_18437,N_18223,N_17965);
xnor U18438 (N_18438,N_17993,N_18142);
nand U18439 (N_18439,N_17686,N_17996);
xor U18440 (N_18440,N_18012,N_18123);
nand U18441 (N_18441,N_17994,N_17942);
or U18442 (N_18442,N_18255,N_17915);
and U18443 (N_18443,N_17983,N_18076);
nor U18444 (N_18444,N_18311,N_17767);
xnor U18445 (N_18445,N_17864,N_18202);
nand U18446 (N_18446,N_17716,N_17928);
xnor U18447 (N_18447,N_18243,N_18299);
or U18448 (N_18448,N_18383,N_17859);
and U18449 (N_18449,N_17980,N_17933);
or U18450 (N_18450,N_18093,N_17891);
nand U18451 (N_18451,N_18238,N_17615);
nand U18452 (N_18452,N_18208,N_18030);
or U18453 (N_18453,N_17665,N_18027);
xor U18454 (N_18454,N_18272,N_18021);
or U18455 (N_18455,N_17726,N_17773);
xnor U18456 (N_18456,N_17830,N_18108);
xnor U18457 (N_18457,N_17969,N_18294);
or U18458 (N_18458,N_18173,N_17739);
or U18459 (N_18459,N_18391,N_18034);
and U18460 (N_18460,N_18348,N_17874);
nor U18461 (N_18461,N_17797,N_17633);
xnor U18462 (N_18462,N_18399,N_18016);
and U18463 (N_18463,N_18178,N_17628);
nand U18464 (N_18464,N_17614,N_18117);
or U18465 (N_18465,N_17781,N_17759);
or U18466 (N_18466,N_18372,N_17745);
or U18467 (N_18467,N_18295,N_17918);
or U18468 (N_18468,N_18109,N_17990);
xor U18469 (N_18469,N_17803,N_18172);
or U18470 (N_18470,N_18338,N_17731);
and U18471 (N_18471,N_17692,N_17631);
and U18472 (N_18472,N_18074,N_18351);
and U18473 (N_18473,N_17936,N_17667);
and U18474 (N_18474,N_18177,N_17722);
and U18475 (N_18475,N_18047,N_17923);
or U18476 (N_18476,N_18070,N_17715);
xor U18477 (N_18477,N_17955,N_18363);
xor U18478 (N_18478,N_18050,N_18007);
nand U18479 (N_18479,N_17911,N_17838);
nand U18480 (N_18480,N_17742,N_17889);
nand U18481 (N_18481,N_18211,N_18337);
or U18482 (N_18482,N_17857,N_17768);
or U18483 (N_18483,N_18303,N_17613);
or U18484 (N_18484,N_18133,N_18059);
xor U18485 (N_18485,N_18162,N_18236);
nor U18486 (N_18486,N_17997,N_17638);
or U18487 (N_18487,N_17680,N_18371);
nand U18488 (N_18488,N_18207,N_17899);
nand U18489 (N_18489,N_17890,N_17682);
xor U18490 (N_18490,N_17728,N_17780);
and U18491 (N_18491,N_18126,N_17836);
and U18492 (N_18492,N_17920,N_17935);
xnor U18493 (N_18493,N_18287,N_18347);
xnor U18494 (N_18494,N_18069,N_18355);
nand U18495 (N_18495,N_17937,N_17802);
xor U18496 (N_18496,N_17647,N_18332);
and U18497 (N_18497,N_18327,N_18176);
xor U18498 (N_18498,N_18161,N_18302);
nor U18499 (N_18499,N_18271,N_18103);
or U18500 (N_18500,N_18056,N_17949);
nor U18501 (N_18501,N_17661,N_18139);
nand U18502 (N_18502,N_17821,N_17953);
and U18503 (N_18503,N_18165,N_18213);
xor U18504 (N_18504,N_17966,N_17982);
nand U18505 (N_18505,N_18341,N_18036);
and U18506 (N_18506,N_18099,N_18171);
or U18507 (N_18507,N_18220,N_17823);
nor U18508 (N_18508,N_18024,N_17629);
and U18509 (N_18509,N_18000,N_18385);
or U18510 (N_18510,N_17725,N_18314);
and U18511 (N_18511,N_18333,N_18087);
nor U18512 (N_18512,N_18288,N_18100);
xor U18513 (N_18513,N_18264,N_18204);
or U18514 (N_18514,N_17730,N_17729);
or U18515 (N_18515,N_18164,N_17960);
nor U18516 (N_18516,N_17684,N_17705);
nor U18517 (N_18517,N_18045,N_18084);
and U18518 (N_18518,N_18079,N_17998);
nand U18519 (N_18519,N_17800,N_18044);
or U18520 (N_18520,N_18107,N_18278);
nand U18521 (N_18521,N_18158,N_18366);
and U18522 (N_18522,N_17626,N_17865);
or U18523 (N_18523,N_18268,N_18038);
or U18524 (N_18524,N_18274,N_17763);
nand U18525 (N_18525,N_18257,N_18248);
nand U18526 (N_18526,N_18121,N_17883);
and U18527 (N_18527,N_18230,N_17818);
or U18528 (N_18528,N_17602,N_17708);
nand U18529 (N_18529,N_18305,N_17664);
nand U18530 (N_18530,N_17776,N_18025);
or U18531 (N_18531,N_18386,N_18357);
and U18532 (N_18532,N_17775,N_17809);
xnor U18533 (N_18533,N_18199,N_17943);
and U18534 (N_18534,N_18013,N_18188);
or U18535 (N_18535,N_17779,N_18129);
or U18536 (N_18536,N_18031,N_18276);
nor U18537 (N_18537,N_17719,N_17792);
or U18538 (N_18538,N_18376,N_17625);
or U18539 (N_18539,N_17951,N_18201);
or U18540 (N_18540,N_18346,N_17627);
nor U18541 (N_18541,N_18358,N_17801);
xor U18542 (N_18542,N_18354,N_18039);
nand U18543 (N_18543,N_17975,N_18041);
nand U18544 (N_18544,N_18067,N_17734);
nor U18545 (N_18545,N_17962,N_17701);
xor U18546 (N_18546,N_18212,N_17979);
and U18547 (N_18547,N_18124,N_17681);
nor U18548 (N_18548,N_18033,N_17663);
or U18549 (N_18549,N_17877,N_18138);
or U18550 (N_18550,N_17907,N_17932);
xor U18551 (N_18551,N_17945,N_18147);
xnor U18552 (N_18552,N_18054,N_17876);
nor U18553 (N_18553,N_17704,N_18216);
nor U18554 (N_18554,N_18170,N_18060);
nand U18555 (N_18555,N_18280,N_17656);
and U18556 (N_18556,N_18018,N_17658);
xor U18557 (N_18557,N_17924,N_17812);
nand U18558 (N_18558,N_18090,N_18397);
nor U18559 (N_18559,N_17654,N_18352);
or U18560 (N_18560,N_17646,N_17756);
or U18561 (N_18561,N_17984,N_17616);
xor U18562 (N_18562,N_18095,N_17738);
and U18563 (N_18563,N_18191,N_17851);
or U18564 (N_18564,N_17909,N_17693);
xor U18565 (N_18565,N_18301,N_18388);
or U18566 (N_18566,N_18384,N_17999);
or U18567 (N_18567,N_17825,N_17892);
or U18568 (N_18568,N_18098,N_18017);
and U18569 (N_18569,N_17764,N_18259);
nor U18570 (N_18570,N_17600,N_17695);
or U18571 (N_18571,N_17846,N_17741);
nor U18572 (N_18572,N_17862,N_17671);
xnor U18573 (N_18573,N_17927,N_17735);
and U18574 (N_18574,N_17748,N_17845);
nor U18575 (N_18575,N_17698,N_17849);
nor U18576 (N_18576,N_18367,N_18159);
xor U18577 (N_18577,N_18231,N_18187);
xor U18578 (N_18578,N_17900,N_18304);
and U18579 (N_18579,N_17806,N_17904);
xor U18580 (N_18580,N_17833,N_18250);
and U18581 (N_18581,N_18342,N_18286);
or U18582 (N_18582,N_17606,N_17981);
xor U18583 (N_18583,N_18375,N_18078);
and U18584 (N_18584,N_17605,N_17973);
xnor U18585 (N_18585,N_17944,N_18392);
nor U18586 (N_18586,N_18320,N_17926);
and U18587 (N_18587,N_18269,N_17707);
nor U18588 (N_18588,N_18313,N_17829);
nand U18589 (N_18589,N_17843,N_17957);
and U18590 (N_18590,N_17898,N_18174);
or U18591 (N_18591,N_18196,N_18061);
xnor U18592 (N_18592,N_18203,N_18394);
or U18593 (N_18593,N_17699,N_18275);
nor U18594 (N_18594,N_18146,N_17618);
and U18595 (N_18595,N_17917,N_17641);
xor U18596 (N_18596,N_18256,N_18042);
or U18597 (N_18597,N_18359,N_17676);
and U18598 (N_18598,N_18277,N_17785);
or U18599 (N_18599,N_18393,N_18240);
or U18600 (N_18600,N_18244,N_17910);
nor U18601 (N_18601,N_17750,N_17740);
or U18602 (N_18602,N_17711,N_18282);
or U18603 (N_18603,N_17956,N_18077);
xnor U18604 (N_18604,N_18330,N_18344);
and U18605 (N_18605,N_18233,N_17645);
and U18606 (N_18606,N_17896,N_18309);
nand U18607 (N_18607,N_18322,N_17880);
nor U18608 (N_18608,N_17769,N_18273);
or U18609 (N_18609,N_18005,N_17713);
nor U18610 (N_18610,N_17621,N_17835);
nand U18611 (N_18611,N_17666,N_18163);
or U18612 (N_18612,N_17690,N_17687);
or U18613 (N_18613,N_18112,N_18323);
nand U18614 (N_18614,N_17778,N_18049);
xor U18615 (N_18615,N_17986,N_17964);
or U18616 (N_18616,N_18221,N_18343);
nand U18617 (N_18617,N_17925,N_17946);
or U18618 (N_18618,N_17908,N_17977);
nor U18619 (N_18619,N_18266,N_17657);
nand U18620 (N_18620,N_17814,N_17619);
or U18621 (N_18621,N_18134,N_18145);
or U18622 (N_18622,N_17612,N_17884);
nor U18623 (N_18623,N_18063,N_17790);
and U18624 (N_18624,N_18227,N_18157);
or U18625 (N_18625,N_17736,N_17815);
nor U18626 (N_18626,N_18200,N_17755);
nor U18627 (N_18627,N_17929,N_18300);
nand U18628 (N_18628,N_17985,N_18283);
nor U18629 (N_18629,N_18246,N_17991);
and U18630 (N_18630,N_17840,N_18195);
and U18631 (N_18631,N_17675,N_18239);
xor U18632 (N_18632,N_17820,N_17674);
nand U18633 (N_18633,N_17746,N_18310);
or U18634 (N_18634,N_17938,N_17844);
nor U18635 (N_18635,N_17660,N_17685);
nor U18636 (N_18636,N_18254,N_18285);
xnor U18637 (N_18637,N_17887,N_18015);
xor U18638 (N_18638,N_17611,N_18316);
xnor U18639 (N_18639,N_17709,N_17640);
nand U18640 (N_18640,N_17930,N_17968);
xor U18641 (N_18641,N_18307,N_17604);
or U18642 (N_18642,N_18390,N_17700);
or U18643 (N_18643,N_18228,N_17751);
nor U18644 (N_18644,N_17897,N_17758);
nor U18645 (N_18645,N_18334,N_18215);
xor U18646 (N_18646,N_17872,N_18105);
or U18647 (N_18647,N_17995,N_18379);
and U18648 (N_18648,N_18149,N_18085);
xor U18649 (N_18649,N_17648,N_17831);
nand U18650 (N_18650,N_17766,N_17706);
nor U18651 (N_18651,N_18198,N_18325);
and U18652 (N_18652,N_18206,N_18279);
and U18653 (N_18653,N_17744,N_17948);
nand U18654 (N_18654,N_18319,N_17772);
and U18655 (N_18655,N_17720,N_17673);
nand U18656 (N_18656,N_17718,N_18321);
xnor U18657 (N_18657,N_18040,N_18290);
nor U18658 (N_18658,N_17789,N_18037);
or U18659 (N_18659,N_17717,N_17819);
or U18660 (N_18660,N_18380,N_18014);
nor U18661 (N_18661,N_17637,N_17888);
xor U18662 (N_18662,N_18219,N_17970);
or U18663 (N_18663,N_17683,N_17732);
xor U18664 (N_18664,N_18029,N_18026);
and U18665 (N_18665,N_17757,N_17978);
nand U18666 (N_18666,N_18291,N_17901);
and U18667 (N_18667,N_18102,N_17644);
and U18668 (N_18668,N_18328,N_17662);
nand U18669 (N_18669,N_18130,N_17799);
nor U18670 (N_18670,N_18395,N_18284);
or U18671 (N_18671,N_18020,N_17762);
and U18672 (N_18672,N_18082,N_17703);
or U18673 (N_18673,N_18247,N_18398);
xnor U18674 (N_18674,N_18065,N_18092);
xor U18675 (N_18675,N_17655,N_17847);
and U18676 (N_18676,N_18356,N_17974);
and U18677 (N_18677,N_17989,N_18062);
nor U18678 (N_18678,N_17765,N_17651);
and U18679 (N_18679,N_17834,N_18369);
and U18680 (N_18680,N_18096,N_18293);
nor U18681 (N_18681,N_18222,N_18035);
nor U18682 (N_18682,N_18306,N_17808);
nor U18683 (N_18683,N_18312,N_18263);
xnor U18684 (N_18684,N_18071,N_17837);
xnor U18685 (N_18685,N_18160,N_17761);
nor U18686 (N_18686,N_18053,N_18209);
or U18687 (N_18687,N_17678,N_17842);
nand U18688 (N_18688,N_17642,N_17941);
nor U18689 (N_18689,N_18179,N_17788);
nand U18690 (N_18690,N_18349,N_17710);
nand U18691 (N_18691,N_17634,N_17774);
nand U18692 (N_18692,N_17650,N_18131);
nand U18693 (N_18693,N_18151,N_17636);
nor U18694 (N_18694,N_17777,N_17848);
or U18695 (N_18695,N_18091,N_17839);
or U18696 (N_18696,N_18088,N_17919);
nor U18697 (N_18697,N_17791,N_18115);
xor U18698 (N_18698,N_17852,N_18153);
xor U18699 (N_18699,N_18345,N_18260);
and U18700 (N_18700,N_18253,N_17902);
nor U18701 (N_18701,N_18072,N_18336);
nor U18702 (N_18702,N_18251,N_18118);
xor U18703 (N_18703,N_17893,N_17855);
and U18704 (N_18704,N_17853,N_18270);
or U18705 (N_18705,N_17620,N_17861);
xor U18706 (N_18706,N_18043,N_18192);
nor U18707 (N_18707,N_17793,N_18073);
and U18708 (N_18708,N_18119,N_17903);
nor U18709 (N_18709,N_17724,N_18097);
xnor U18710 (N_18710,N_18362,N_17639);
nand U18711 (N_18711,N_17958,N_18132);
xor U18712 (N_18712,N_18125,N_17669);
nor U18713 (N_18713,N_18258,N_17770);
nand U18714 (N_18714,N_17954,N_18234);
xor U18715 (N_18715,N_17878,N_17870);
xor U18716 (N_18716,N_18004,N_18252);
or U18717 (N_18717,N_18217,N_18136);
or U18718 (N_18718,N_17931,N_18350);
nor U18719 (N_18719,N_17813,N_17913);
and U18720 (N_18720,N_18370,N_18377);
nor U18721 (N_18721,N_17912,N_18245);
nand U18722 (N_18722,N_18368,N_17712);
or U18723 (N_18723,N_18111,N_18120);
nand U18724 (N_18724,N_17841,N_18353);
nand U18725 (N_18725,N_18180,N_17689);
xor U18726 (N_18726,N_17747,N_17694);
nor U18727 (N_18727,N_17652,N_17622);
or U18728 (N_18728,N_17691,N_17805);
nand U18729 (N_18729,N_17727,N_18382);
xnor U18730 (N_18730,N_18051,N_18169);
and U18731 (N_18731,N_17827,N_18190);
nor U18732 (N_18732,N_18167,N_17643);
nand U18733 (N_18733,N_18086,N_18028);
nand U18734 (N_18734,N_18292,N_18361);
xor U18735 (N_18735,N_17784,N_17733);
or U18736 (N_18736,N_17702,N_18237);
xnor U18737 (N_18737,N_18242,N_17914);
nand U18738 (N_18738,N_18008,N_18262);
nand U18739 (N_18739,N_17688,N_17607);
or U18740 (N_18740,N_18185,N_17608);
or U18741 (N_18741,N_18298,N_18075);
nor U18742 (N_18742,N_17749,N_18127);
or U18743 (N_18743,N_18148,N_17922);
nor U18744 (N_18744,N_17869,N_17743);
nand U18745 (N_18745,N_17868,N_18068);
or U18746 (N_18746,N_17905,N_17610);
xor U18747 (N_18747,N_18066,N_17737);
or U18748 (N_18748,N_17921,N_18331);
nor U18749 (N_18749,N_17810,N_17670);
and U18750 (N_18750,N_17972,N_18094);
nor U18751 (N_18751,N_18194,N_17850);
or U18752 (N_18752,N_18106,N_17603);
nand U18753 (N_18753,N_17961,N_18261);
nor U18754 (N_18754,N_18318,N_17867);
nor U18755 (N_18755,N_17894,N_17988);
xor U18756 (N_18756,N_18101,N_17875);
nor U18757 (N_18757,N_18267,N_17760);
nor U18758 (N_18758,N_18046,N_18381);
and U18759 (N_18759,N_18003,N_18081);
and U18760 (N_18760,N_17832,N_18317);
or U18761 (N_18761,N_17804,N_17753);
nor U18762 (N_18762,N_17826,N_18137);
and U18763 (N_18763,N_17786,N_17807);
xor U18764 (N_18764,N_18057,N_17782);
nand U18765 (N_18765,N_18340,N_17866);
nand U18766 (N_18766,N_17906,N_18232);
nor U18767 (N_18767,N_18064,N_18110);
and U18768 (N_18768,N_18168,N_17679);
and U18769 (N_18769,N_18152,N_18365);
and U18770 (N_18770,N_17873,N_18265);
nor U18771 (N_18771,N_17895,N_17817);
nand U18772 (N_18772,N_18116,N_18010);
or U18773 (N_18773,N_18052,N_17816);
nor U18774 (N_18774,N_18009,N_18214);
nor U18775 (N_18775,N_17635,N_17963);
nand U18776 (N_18776,N_18001,N_17653);
xnor U18777 (N_18777,N_18364,N_18166);
or U18778 (N_18778,N_17714,N_17798);
and U18779 (N_18779,N_17783,N_17787);
nand U18780 (N_18780,N_18396,N_17959);
or U18781 (N_18781,N_18104,N_18229);
nand U18782 (N_18782,N_18339,N_17771);
and U18783 (N_18783,N_18329,N_17863);
nand U18784 (N_18784,N_18089,N_18297);
nor U18785 (N_18785,N_17858,N_17916);
xor U18786 (N_18786,N_18156,N_17795);
or U18787 (N_18787,N_18140,N_18249);
nor U18788 (N_18788,N_18197,N_17885);
and U18789 (N_18789,N_18184,N_18241);
or U18790 (N_18790,N_18011,N_18181);
and U18791 (N_18791,N_17632,N_18155);
xnor U18792 (N_18792,N_18175,N_18083);
and U18793 (N_18793,N_17987,N_17649);
nand U18794 (N_18794,N_18055,N_18135);
nor U18795 (N_18795,N_18315,N_18374);
xnor U18796 (N_18796,N_18193,N_17601);
and U18797 (N_18797,N_17752,N_18154);
and U18798 (N_18798,N_18023,N_17696);
nor U18799 (N_18799,N_17723,N_17822);
nand U18800 (N_18800,N_18373,N_17734);
nand U18801 (N_18801,N_17660,N_17870);
nand U18802 (N_18802,N_18031,N_17831);
nor U18803 (N_18803,N_18268,N_18349);
xor U18804 (N_18804,N_17881,N_17944);
xnor U18805 (N_18805,N_17963,N_17707);
xor U18806 (N_18806,N_18350,N_17648);
and U18807 (N_18807,N_18113,N_17760);
nor U18808 (N_18808,N_18125,N_17980);
nor U18809 (N_18809,N_18148,N_18191);
and U18810 (N_18810,N_17852,N_18117);
xor U18811 (N_18811,N_18347,N_17837);
nor U18812 (N_18812,N_18385,N_18357);
and U18813 (N_18813,N_17793,N_18279);
and U18814 (N_18814,N_18029,N_17888);
and U18815 (N_18815,N_18343,N_17760);
xor U18816 (N_18816,N_17622,N_17877);
nor U18817 (N_18817,N_18016,N_18034);
and U18818 (N_18818,N_18194,N_17763);
and U18819 (N_18819,N_17770,N_18017);
nand U18820 (N_18820,N_18112,N_18154);
xnor U18821 (N_18821,N_17926,N_17879);
nand U18822 (N_18822,N_17849,N_17845);
xor U18823 (N_18823,N_18227,N_17740);
or U18824 (N_18824,N_17949,N_18105);
nor U18825 (N_18825,N_17691,N_18170);
or U18826 (N_18826,N_18269,N_18047);
or U18827 (N_18827,N_18290,N_18389);
nand U18828 (N_18828,N_17660,N_17691);
or U18829 (N_18829,N_17648,N_17652);
and U18830 (N_18830,N_18368,N_17965);
xor U18831 (N_18831,N_17768,N_18011);
and U18832 (N_18832,N_17975,N_17968);
xnor U18833 (N_18833,N_18303,N_17878);
and U18834 (N_18834,N_18341,N_17690);
nand U18835 (N_18835,N_18191,N_17996);
and U18836 (N_18836,N_17787,N_17723);
and U18837 (N_18837,N_17718,N_17603);
or U18838 (N_18838,N_18291,N_18101);
or U18839 (N_18839,N_18094,N_18000);
nor U18840 (N_18840,N_17789,N_18176);
nand U18841 (N_18841,N_17966,N_17780);
nand U18842 (N_18842,N_17850,N_18387);
or U18843 (N_18843,N_17753,N_18072);
or U18844 (N_18844,N_17785,N_18260);
nor U18845 (N_18845,N_17641,N_17797);
xnor U18846 (N_18846,N_17718,N_18087);
or U18847 (N_18847,N_18055,N_17819);
nand U18848 (N_18848,N_18232,N_17916);
nand U18849 (N_18849,N_18277,N_18202);
nand U18850 (N_18850,N_17872,N_18174);
nand U18851 (N_18851,N_18172,N_18324);
xnor U18852 (N_18852,N_18062,N_17686);
nor U18853 (N_18853,N_17791,N_18347);
or U18854 (N_18854,N_18249,N_18048);
nand U18855 (N_18855,N_18219,N_18132);
nor U18856 (N_18856,N_18394,N_18336);
xor U18857 (N_18857,N_17762,N_18377);
and U18858 (N_18858,N_17999,N_17819);
nand U18859 (N_18859,N_17761,N_17748);
or U18860 (N_18860,N_17931,N_17656);
or U18861 (N_18861,N_18016,N_18007);
xnor U18862 (N_18862,N_18326,N_17878);
or U18863 (N_18863,N_18011,N_18283);
xnor U18864 (N_18864,N_17631,N_18276);
nor U18865 (N_18865,N_18234,N_18239);
nor U18866 (N_18866,N_18361,N_17681);
nand U18867 (N_18867,N_18280,N_17735);
or U18868 (N_18868,N_18239,N_17983);
or U18869 (N_18869,N_17945,N_17879);
nor U18870 (N_18870,N_18275,N_17907);
nand U18871 (N_18871,N_17866,N_18289);
and U18872 (N_18872,N_18239,N_18236);
xnor U18873 (N_18873,N_17956,N_17790);
nor U18874 (N_18874,N_17803,N_17968);
xor U18875 (N_18875,N_18082,N_17944);
xor U18876 (N_18876,N_18084,N_17603);
or U18877 (N_18877,N_17896,N_18107);
or U18878 (N_18878,N_17732,N_18093);
or U18879 (N_18879,N_18259,N_18036);
or U18880 (N_18880,N_17949,N_18181);
nand U18881 (N_18881,N_17996,N_18087);
or U18882 (N_18882,N_18323,N_18073);
or U18883 (N_18883,N_18384,N_17718);
nor U18884 (N_18884,N_17888,N_17698);
or U18885 (N_18885,N_18122,N_18158);
xnor U18886 (N_18886,N_17602,N_17649);
nor U18887 (N_18887,N_17665,N_18320);
nand U18888 (N_18888,N_18253,N_17654);
or U18889 (N_18889,N_17814,N_18129);
xor U18890 (N_18890,N_17813,N_18108);
nand U18891 (N_18891,N_17872,N_18389);
xnor U18892 (N_18892,N_17861,N_17615);
nor U18893 (N_18893,N_18272,N_18217);
nor U18894 (N_18894,N_17726,N_17886);
and U18895 (N_18895,N_18252,N_18078);
nand U18896 (N_18896,N_17722,N_18072);
or U18897 (N_18897,N_17620,N_17657);
nand U18898 (N_18898,N_18307,N_18155);
xnor U18899 (N_18899,N_17793,N_18032);
nand U18900 (N_18900,N_18317,N_18047);
and U18901 (N_18901,N_17997,N_18281);
xnor U18902 (N_18902,N_17821,N_18120);
xor U18903 (N_18903,N_17856,N_17891);
xor U18904 (N_18904,N_17807,N_18033);
or U18905 (N_18905,N_18046,N_17874);
xor U18906 (N_18906,N_18287,N_18182);
or U18907 (N_18907,N_17955,N_18081);
nand U18908 (N_18908,N_18238,N_17735);
or U18909 (N_18909,N_18352,N_18007);
or U18910 (N_18910,N_17727,N_17661);
or U18911 (N_18911,N_17954,N_18106);
nor U18912 (N_18912,N_18132,N_17814);
and U18913 (N_18913,N_17652,N_17689);
nor U18914 (N_18914,N_18169,N_18043);
nor U18915 (N_18915,N_17900,N_18070);
nand U18916 (N_18916,N_17954,N_17986);
xor U18917 (N_18917,N_18165,N_18309);
nor U18918 (N_18918,N_17985,N_17753);
xor U18919 (N_18919,N_18163,N_18032);
or U18920 (N_18920,N_18067,N_18296);
xnor U18921 (N_18921,N_17790,N_17954);
and U18922 (N_18922,N_17756,N_17889);
nor U18923 (N_18923,N_17980,N_17808);
and U18924 (N_18924,N_18191,N_17843);
or U18925 (N_18925,N_17926,N_17890);
xnor U18926 (N_18926,N_17631,N_17909);
xor U18927 (N_18927,N_17979,N_18026);
or U18928 (N_18928,N_18298,N_17760);
and U18929 (N_18929,N_17943,N_17807);
or U18930 (N_18930,N_17742,N_17763);
nand U18931 (N_18931,N_17997,N_18350);
nor U18932 (N_18932,N_18032,N_17718);
nor U18933 (N_18933,N_18113,N_17759);
and U18934 (N_18934,N_17608,N_18346);
nand U18935 (N_18935,N_18025,N_18075);
or U18936 (N_18936,N_18349,N_17858);
nand U18937 (N_18937,N_18128,N_18214);
or U18938 (N_18938,N_18031,N_17956);
nand U18939 (N_18939,N_17918,N_17912);
nand U18940 (N_18940,N_18315,N_18085);
nor U18941 (N_18941,N_17716,N_17870);
or U18942 (N_18942,N_17890,N_17925);
or U18943 (N_18943,N_18319,N_18310);
or U18944 (N_18944,N_17614,N_17973);
or U18945 (N_18945,N_17764,N_17637);
or U18946 (N_18946,N_17692,N_18001);
and U18947 (N_18947,N_18069,N_17754);
nor U18948 (N_18948,N_17852,N_18119);
nor U18949 (N_18949,N_17748,N_18268);
nand U18950 (N_18950,N_17974,N_18336);
and U18951 (N_18951,N_17693,N_17923);
nor U18952 (N_18952,N_17964,N_18113);
and U18953 (N_18953,N_17721,N_17632);
and U18954 (N_18954,N_18301,N_18085);
xnor U18955 (N_18955,N_18030,N_18134);
or U18956 (N_18956,N_17724,N_17676);
nor U18957 (N_18957,N_18104,N_17988);
or U18958 (N_18958,N_18235,N_17673);
nand U18959 (N_18959,N_17879,N_18076);
xor U18960 (N_18960,N_17627,N_17650);
and U18961 (N_18961,N_18067,N_18096);
and U18962 (N_18962,N_18049,N_18291);
xor U18963 (N_18963,N_18024,N_17771);
or U18964 (N_18964,N_17839,N_18209);
xor U18965 (N_18965,N_18386,N_17626);
nand U18966 (N_18966,N_17805,N_17841);
nand U18967 (N_18967,N_17669,N_18144);
or U18968 (N_18968,N_17845,N_17634);
xor U18969 (N_18969,N_18155,N_17935);
nor U18970 (N_18970,N_18070,N_18071);
xnor U18971 (N_18971,N_18019,N_18062);
xnor U18972 (N_18972,N_17999,N_17967);
nand U18973 (N_18973,N_18345,N_17970);
or U18974 (N_18974,N_18146,N_17757);
or U18975 (N_18975,N_18263,N_17890);
or U18976 (N_18976,N_18255,N_18264);
or U18977 (N_18977,N_17849,N_18261);
nor U18978 (N_18978,N_18286,N_17973);
nor U18979 (N_18979,N_17893,N_17883);
xor U18980 (N_18980,N_17709,N_17662);
nor U18981 (N_18981,N_17807,N_17891);
nand U18982 (N_18982,N_18253,N_17847);
nor U18983 (N_18983,N_17621,N_18128);
and U18984 (N_18984,N_17813,N_18200);
nor U18985 (N_18985,N_17614,N_18241);
or U18986 (N_18986,N_17638,N_17659);
xnor U18987 (N_18987,N_17921,N_17721);
and U18988 (N_18988,N_17956,N_17714);
nor U18989 (N_18989,N_18113,N_18192);
nor U18990 (N_18990,N_18018,N_18298);
nand U18991 (N_18991,N_17811,N_18340);
nor U18992 (N_18992,N_18386,N_17854);
and U18993 (N_18993,N_18285,N_18169);
and U18994 (N_18994,N_17848,N_17950);
and U18995 (N_18995,N_17689,N_18350);
xnor U18996 (N_18996,N_18079,N_18372);
and U18997 (N_18997,N_17692,N_18063);
nand U18998 (N_18998,N_18260,N_17738);
nor U18999 (N_18999,N_18084,N_17875);
nand U19000 (N_19000,N_17681,N_17705);
nand U19001 (N_19001,N_17807,N_17781);
and U19002 (N_19002,N_17854,N_18064);
nand U19003 (N_19003,N_18205,N_18119);
and U19004 (N_19004,N_18354,N_18143);
and U19005 (N_19005,N_17988,N_17949);
nand U19006 (N_19006,N_17655,N_17846);
or U19007 (N_19007,N_18313,N_17704);
or U19008 (N_19008,N_18256,N_17941);
nor U19009 (N_19009,N_17806,N_18316);
xnor U19010 (N_19010,N_17781,N_17601);
xnor U19011 (N_19011,N_18194,N_17894);
or U19012 (N_19012,N_18142,N_18077);
nor U19013 (N_19013,N_18301,N_18119);
and U19014 (N_19014,N_18264,N_18061);
nor U19015 (N_19015,N_18393,N_17606);
nand U19016 (N_19016,N_17993,N_17727);
or U19017 (N_19017,N_17976,N_18165);
nand U19018 (N_19018,N_17922,N_17986);
nand U19019 (N_19019,N_18348,N_17824);
and U19020 (N_19020,N_18036,N_18000);
nand U19021 (N_19021,N_17777,N_17792);
or U19022 (N_19022,N_17979,N_18097);
or U19023 (N_19023,N_17858,N_18099);
xor U19024 (N_19024,N_18200,N_17756);
xor U19025 (N_19025,N_18358,N_17840);
nand U19026 (N_19026,N_18312,N_18052);
nand U19027 (N_19027,N_17651,N_18063);
or U19028 (N_19028,N_17624,N_18195);
nand U19029 (N_19029,N_17865,N_18248);
and U19030 (N_19030,N_17836,N_18341);
or U19031 (N_19031,N_18094,N_17720);
xor U19032 (N_19032,N_17808,N_17746);
nand U19033 (N_19033,N_18075,N_18067);
nor U19034 (N_19034,N_17912,N_17779);
nand U19035 (N_19035,N_17645,N_18091);
and U19036 (N_19036,N_17770,N_18009);
xnor U19037 (N_19037,N_17693,N_18290);
nand U19038 (N_19038,N_18105,N_18069);
nor U19039 (N_19039,N_18127,N_18004);
nor U19040 (N_19040,N_17709,N_17672);
and U19041 (N_19041,N_17932,N_17736);
nand U19042 (N_19042,N_18364,N_18298);
nand U19043 (N_19043,N_18213,N_17903);
nor U19044 (N_19044,N_18287,N_18080);
xnor U19045 (N_19045,N_17761,N_17870);
and U19046 (N_19046,N_18134,N_17764);
or U19047 (N_19047,N_18148,N_17670);
nor U19048 (N_19048,N_17882,N_17820);
and U19049 (N_19049,N_18283,N_17848);
nor U19050 (N_19050,N_18124,N_17885);
nand U19051 (N_19051,N_18311,N_18147);
xor U19052 (N_19052,N_18106,N_17632);
nor U19053 (N_19053,N_18351,N_17849);
nand U19054 (N_19054,N_18085,N_18170);
xnor U19055 (N_19055,N_17708,N_17623);
and U19056 (N_19056,N_18349,N_17731);
xnor U19057 (N_19057,N_17641,N_17722);
xnor U19058 (N_19058,N_17769,N_17734);
nor U19059 (N_19059,N_17989,N_18364);
xor U19060 (N_19060,N_18136,N_18024);
xor U19061 (N_19061,N_18199,N_18031);
nand U19062 (N_19062,N_18014,N_17887);
or U19063 (N_19063,N_18171,N_18246);
xnor U19064 (N_19064,N_17644,N_18259);
nor U19065 (N_19065,N_18163,N_18398);
and U19066 (N_19066,N_18384,N_18048);
or U19067 (N_19067,N_18011,N_18293);
or U19068 (N_19068,N_17701,N_18221);
nor U19069 (N_19069,N_17861,N_18137);
xnor U19070 (N_19070,N_18336,N_18292);
nor U19071 (N_19071,N_17910,N_17837);
nand U19072 (N_19072,N_17898,N_17737);
xor U19073 (N_19073,N_18009,N_17656);
and U19074 (N_19074,N_17949,N_17684);
nand U19075 (N_19075,N_17869,N_17749);
or U19076 (N_19076,N_17903,N_17992);
and U19077 (N_19077,N_17712,N_18138);
nand U19078 (N_19078,N_17666,N_17940);
or U19079 (N_19079,N_18221,N_18301);
nor U19080 (N_19080,N_17833,N_17832);
and U19081 (N_19081,N_17621,N_17779);
or U19082 (N_19082,N_17753,N_17873);
or U19083 (N_19083,N_17653,N_17889);
xnor U19084 (N_19084,N_17903,N_18316);
nand U19085 (N_19085,N_17959,N_18302);
xor U19086 (N_19086,N_17899,N_18019);
and U19087 (N_19087,N_17718,N_18142);
xnor U19088 (N_19088,N_18377,N_17727);
or U19089 (N_19089,N_17815,N_18383);
and U19090 (N_19090,N_17952,N_17723);
xnor U19091 (N_19091,N_18378,N_18203);
and U19092 (N_19092,N_17951,N_18296);
xor U19093 (N_19093,N_17604,N_18003);
and U19094 (N_19094,N_18052,N_17895);
or U19095 (N_19095,N_17820,N_17804);
nor U19096 (N_19096,N_17877,N_17897);
xor U19097 (N_19097,N_18282,N_18380);
nand U19098 (N_19098,N_17679,N_18380);
nor U19099 (N_19099,N_18142,N_18169);
or U19100 (N_19100,N_17943,N_17742);
xnor U19101 (N_19101,N_17865,N_18290);
and U19102 (N_19102,N_18198,N_17658);
and U19103 (N_19103,N_17749,N_17988);
nand U19104 (N_19104,N_17722,N_18180);
and U19105 (N_19105,N_18089,N_18208);
or U19106 (N_19106,N_17639,N_17645);
or U19107 (N_19107,N_18273,N_17739);
xnor U19108 (N_19108,N_18155,N_17605);
nor U19109 (N_19109,N_18352,N_18220);
nor U19110 (N_19110,N_17887,N_17942);
and U19111 (N_19111,N_18345,N_17947);
nand U19112 (N_19112,N_17822,N_18045);
xnor U19113 (N_19113,N_17608,N_17805);
and U19114 (N_19114,N_18162,N_17994);
and U19115 (N_19115,N_17964,N_18313);
nor U19116 (N_19116,N_17601,N_17862);
nand U19117 (N_19117,N_17948,N_17776);
and U19118 (N_19118,N_17661,N_18194);
and U19119 (N_19119,N_17776,N_18037);
xor U19120 (N_19120,N_17664,N_17756);
nor U19121 (N_19121,N_17826,N_18322);
xor U19122 (N_19122,N_18113,N_18253);
xor U19123 (N_19123,N_17610,N_17736);
xnor U19124 (N_19124,N_18179,N_17943);
xor U19125 (N_19125,N_17787,N_17752);
nand U19126 (N_19126,N_18063,N_17653);
or U19127 (N_19127,N_17957,N_18342);
nor U19128 (N_19128,N_17760,N_17722);
nand U19129 (N_19129,N_17816,N_18093);
and U19130 (N_19130,N_17818,N_17906);
xnor U19131 (N_19131,N_17686,N_18137);
xnor U19132 (N_19132,N_18286,N_18037);
or U19133 (N_19133,N_18106,N_17703);
nand U19134 (N_19134,N_18213,N_17886);
nand U19135 (N_19135,N_18233,N_18064);
xor U19136 (N_19136,N_18188,N_18313);
and U19137 (N_19137,N_18301,N_17834);
nor U19138 (N_19138,N_18259,N_18015);
xnor U19139 (N_19139,N_18168,N_18205);
xor U19140 (N_19140,N_18296,N_18083);
nand U19141 (N_19141,N_18039,N_17670);
or U19142 (N_19142,N_17824,N_18109);
xor U19143 (N_19143,N_18066,N_18250);
nor U19144 (N_19144,N_18389,N_17771);
nand U19145 (N_19145,N_18085,N_18357);
and U19146 (N_19146,N_18063,N_18178);
and U19147 (N_19147,N_17998,N_18290);
nand U19148 (N_19148,N_18128,N_17661);
or U19149 (N_19149,N_17743,N_18070);
nand U19150 (N_19150,N_18062,N_18133);
or U19151 (N_19151,N_18197,N_18027);
and U19152 (N_19152,N_18315,N_17794);
and U19153 (N_19153,N_18216,N_18388);
xor U19154 (N_19154,N_17767,N_18252);
xnor U19155 (N_19155,N_17946,N_17851);
xor U19156 (N_19156,N_18152,N_18225);
and U19157 (N_19157,N_18312,N_17737);
xnor U19158 (N_19158,N_18098,N_17842);
xor U19159 (N_19159,N_17728,N_18307);
xnor U19160 (N_19160,N_18366,N_17963);
nor U19161 (N_19161,N_17923,N_17893);
and U19162 (N_19162,N_18381,N_17710);
nor U19163 (N_19163,N_17791,N_17944);
or U19164 (N_19164,N_17956,N_17624);
nand U19165 (N_19165,N_18272,N_18229);
nor U19166 (N_19166,N_18374,N_17639);
and U19167 (N_19167,N_18325,N_17913);
or U19168 (N_19168,N_17888,N_18310);
nand U19169 (N_19169,N_18287,N_17939);
or U19170 (N_19170,N_17687,N_18083);
nand U19171 (N_19171,N_18018,N_18354);
nand U19172 (N_19172,N_17972,N_18281);
nand U19173 (N_19173,N_17701,N_17824);
xnor U19174 (N_19174,N_18389,N_17854);
or U19175 (N_19175,N_17969,N_17987);
and U19176 (N_19176,N_17606,N_18315);
or U19177 (N_19177,N_17680,N_17885);
or U19178 (N_19178,N_17930,N_18343);
or U19179 (N_19179,N_18368,N_17693);
nand U19180 (N_19180,N_17954,N_17976);
and U19181 (N_19181,N_18005,N_18244);
or U19182 (N_19182,N_18250,N_17779);
nor U19183 (N_19183,N_17623,N_17947);
nand U19184 (N_19184,N_17657,N_18098);
xnor U19185 (N_19185,N_18153,N_18289);
nor U19186 (N_19186,N_18118,N_17992);
nand U19187 (N_19187,N_17971,N_18318);
nor U19188 (N_19188,N_17768,N_17816);
or U19189 (N_19189,N_17747,N_17974);
nor U19190 (N_19190,N_17989,N_17774);
and U19191 (N_19191,N_17834,N_18191);
or U19192 (N_19192,N_18151,N_18205);
xor U19193 (N_19193,N_18039,N_17902);
nor U19194 (N_19194,N_17832,N_18211);
or U19195 (N_19195,N_18018,N_18164);
or U19196 (N_19196,N_18260,N_17941);
xor U19197 (N_19197,N_18028,N_17832);
nand U19198 (N_19198,N_18185,N_17949);
or U19199 (N_19199,N_17624,N_18372);
xnor U19200 (N_19200,N_18526,N_18647);
or U19201 (N_19201,N_18772,N_18921);
or U19202 (N_19202,N_18497,N_19016);
nor U19203 (N_19203,N_19037,N_18759);
nor U19204 (N_19204,N_18673,N_19099);
and U19205 (N_19205,N_19147,N_19088);
xnor U19206 (N_19206,N_18656,N_19114);
or U19207 (N_19207,N_18778,N_18803);
nand U19208 (N_19208,N_18739,N_18812);
nand U19209 (N_19209,N_19026,N_18948);
xnor U19210 (N_19210,N_19005,N_18483);
and U19211 (N_19211,N_19188,N_18512);
xor U19212 (N_19212,N_19044,N_19042);
and U19213 (N_19213,N_18462,N_19121);
nand U19214 (N_19214,N_19194,N_18563);
or U19215 (N_19215,N_18791,N_18655);
and U19216 (N_19216,N_19067,N_18498);
xor U19217 (N_19217,N_18614,N_18826);
nor U19218 (N_19218,N_18914,N_18795);
xor U19219 (N_19219,N_18797,N_18924);
xnor U19220 (N_19220,N_18560,N_18814);
xor U19221 (N_19221,N_18474,N_18600);
xnor U19222 (N_19222,N_18876,N_19109);
and U19223 (N_19223,N_18771,N_18975);
and U19224 (N_19224,N_18405,N_18748);
or U19225 (N_19225,N_19155,N_18694);
nor U19226 (N_19226,N_18952,N_18735);
nand U19227 (N_19227,N_18603,N_18670);
nor U19228 (N_19228,N_18738,N_18666);
xnor U19229 (N_19229,N_18743,N_18710);
or U19230 (N_19230,N_18685,N_18538);
or U19231 (N_19231,N_19177,N_18686);
nor U19232 (N_19232,N_18620,N_18744);
and U19233 (N_19233,N_18494,N_18572);
or U19234 (N_19234,N_18937,N_19000);
or U19235 (N_19235,N_19186,N_18981);
and U19236 (N_19236,N_18613,N_19091);
xnor U19237 (N_19237,N_18816,N_18773);
and U19238 (N_19238,N_18467,N_19185);
nand U19239 (N_19239,N_18678,N_19065);
and U19240 (N_19240,N_19152,N_18839);
xnor U19241 (N_19241,N_18630,N_18561);
xor U19242 (N_19242,N_18945,N_19009);
nand U19243 (N_19243,N_18721,N_18882);
or U19244 (N_19244,N_18903,N_18697);
nand U19245 (N_19245,N_18523,N_18754);
or U19246 (N_19246,N_18869,N_18492);
nand U19247 (N_19247,N_18861,N_18763);
xor U19248 (N_19248,N_18764,N_18409);
and U19249 (N_19249,N_18846,N_18419);
or U19250 (N_19250,N_18435,N_18477);
or U19251 (N_19251,N_18706,N_18995);
or U19252 (N_19252,N_19193,N_18808);
or U19253 (N_19253,N_18732,N_18550);
and U19254 (N_19254,N_18902,N_18544);
nand U19255 (N_19255,N_18508,N_19124);
or U19256 (N_19256,N_18499,N_19018);
and U19257 (N_19257,N_18923,N_19003);
nor U19258 (N_19258,N_18646,N_19111);
and U19259 (N_19259,N_18968,N_18459);
xor U19260 (N_19260,N_18448,N_19174);
nand U19261 (N_19261,N_19045,N_19029);
xor U19262 (N_19262,N_18810,N_18601);
xor U19263 (N_19263,N_18885,N_19068);
or U19264 (N_19264,N_19137,N_18619);
xnor U19265 (N_19265,N_19182,N_18449);
nor U19266 (N_19266,N_18677,N_18729);
nand U19267 (N_19267,N_18667,N_18622);
or U19268 (N_19268,N_19151,N_18915);
and U19269 (N_19269,N_19004,N_18974);
nor U19270 (N_19270,N_19022,N_19138);
xor U19271 (N_19271,N_19041,N_18482);
xnor U19272 (N_19272,N_18634,N_18478);
xor U19273 (N_19273,N_19096,N_19093);
nor U19274 (N_19274,N_18446,N_19136);
xor U19275 (N_19275,N_19019,N_19198);
and U19276 (N_19276,N_18931,N_18450);
nand U19277 (N_19277,N_18940,N_19132);
xor U19278 (N_19278,N_18549,N_18755);
nand U19279 (N_19279,N_18779,N_18994);
xnor U19280 (N_19280,N_18993,N_18432);
nand U19281 (N_19281,N_18798,N_18730);
nor U19282 (N_19282,N_19144,N_19184);
nor U19283 (N_19283,N_18800,N_18919);
and U19284 (N_19284,N_19113,N_18621);
or U19285 (N_19285,N_18407,N_18645);
xnor U19286 (N_19286,N_18525,N_18946);
xor U19287 (N_19287,N_19010,N_19076);
nor U19288 (N_19288,N_19130,N_19170);
xnor U19289 (N_19289,N_18842,N_19085);
nor U19290 (N_19290,N_18980,N_19049);
or U19291 (N_19291,N_18418,N_18546);
and U19292 (N_19292,N_18695,N_18972);
nor U19293 (N_19293,N_18674,N_18648);
or U19294 (N_19294,N_18425,N_18504);
and U19295 (N_19295,N_18590,N_18401);
nor U19296 (N_19296,N_18470,N_18668);
nor U19297 (N_19297,N_18671,N_18868);
and U19298 (N_19298,N_18437,N_18468);
nand U19299 (N_19299,N_18776,N_19165);
and U19300 (N_19300,N_18616,N_18997);
and U19301 (N_19301,N_18723,N_18724);
nor U19302 (N_19302,N_18751,N_18741);
nand U19303 (N_19303,N_18978,N_18818);
xor U19304 (N_19304,N_18822,N_18782);
nand U19305 (N_19305,N_18500,N_18874);
and U19306 (N_19306,N_18951,N_18586);
xor U19307 (N_19307,N_18925,N_19122);
nor U19308 (N_19308,N_18817,N_18650);
and U19309 (N_19309,N_19169,N_18917);
and U19310 (N_19310,N_18658,N_18983);
nand U19311 (N_19311,N_18899,N_19115);
or U19312 (N_19312,N_18712,N_18889);
nand U19313 (N_19313,N_18760,N_18976);
nor U19314 (N_19314,N_19142,N_18780);
nand U19315 (N_19315,N_18688,N_18594);
and U19316 (N_19316,N_19025,N_18934);
and U19317 (N_19317,N_18959,N_18495);
xnor U19318 (N_19318,N_19059,N_18665);
and U19319 (N_19319,N_18789,N_19092);
and U19320 (N_19320,N_18774,N_19064);
or U19321 (N_19321,N_18641,N_18973);
and U19322 (N_19322,N_18871,N_19048);
and U19323 (N_19323,N_18431,N_18421);
and U19324 (N_19324,N_18570,N_18749);
nand U19325 (N_19325,N_18854,N_18740);
nor U19326 (N_19326,N_19168,N_18843);
nor U19327 (N_19327,N_18815,N_18888);
nand U19328 (N_19328,N_18480,N_19158);
nand U19329 (N_19329,N_18716,N_19011);
and U19330 (N_19330,N_18958,N_18784);
or U19331 (N_19331,N_18651,N_18460);
nand U19332 (N_19332,N_18476,N_18990);
xor U19333 (N_19333,N_19102,N_19001);
or U19334 (N_19334,N_18558,N_18583);
xnor U19335 (N_19335,N_18408,N_18631);
xor U19336 (N_19336,N_18769,N_19128);
xnor U19337 (N_19337,N_18638,N_19087);
xnor U19338 (N_19338,N_18672,N_18604);
nor U19339 (N_19339,N_19154,N_18530);
nor U19340 (N_19340,N_19020,N_18865);
xor U19341 (N_19341,N_18832,N_18676);
or U19342 (N_19342,N_18747,N_18969);
or U19343 (N_19343,N_19149,N_18593);
nor U19344 (N_19344,N_19043,N_18746);
and U19345 (N_19345,N_18720,N_19118);
nand U19346 (N_19346,N_18529,N_18768);
and U19347 (N_19347,N_19021,N_18653);
xnor U19348 (N_19348,N_18971,N_18633);
nand U19349 (N_19349,N_18841,N_18553);
nor U19350 (N_19350,N_18608,N_18813);
or U19351 (N_19351,N_18592,N_19148);
xor U19352 (N_19352,N_18873,N_19069);
and U19353 (N_19353,N_18982,N_19007);
or U19354 (N_19354,N_18829,N_18750);
or U19355 (N_19355,N_18537,N_19008);
and U19356 (N_19356,N_18488,N_19028);
or U19357 (N_19357,N_18589,N_18752);
or U19358 (N_19358,N_18949,N_18424);
nor U19359 (N_19359,N_18605,N_19112);
or U19360 (N_19360,N_19103,N_18933);
nand U19361 (N_19361,N_18491,N_18867);
or U19362 (N_19362,N_18836,N_18757);
xnor U19363 (N_19363,N_19107,N_19055);
and U19364 (N_19364,N_18442,N_19108);
or U19365 (N_19365,N_18811,N_18514);
nor U19366 (N_19366,N_19033,N_18416);
and U19367 (N_19367,N_18864,N_18484);
and U19368 (N_19368,N_18506,N_19006);
nor U19369 (N_19369,N_18535,N_19176);
xnor U19370 (N_19370,N_18696,N_18853);
or U19371 (N_19371,N_18580,N_18629);
nor U19372 (N_19372,N_18742,N_18898);
and U19373 (N_19373,N_18693,N_18922);
nor U19374 (N_19374,N_18907,N_18911);
xor U19375 (N_19375,N_18420,N_18439);
xor U19376 (N_19376,N_19190,N_18939);
and U19377 (N_19377,N_18823,N_18856);
or U19378 (N_19378,N_19027,N_18910);
nor U19379 (N_19379,N_18684,N_19105);
and U19380 (N_19380,N_18935,N_18767);
and U19381 (N_19381,N_19035,N_18878);
xnor U19382 (N_19382,N_19110,N_19036);
nand U19383 (N_19383,N_18661,N_18970);
xnor U19384 (N_19384,N_18766,N_19199);
and U19385 (N_19385,N_19046,N_18705);
and U19386 (N_19386,N_18429,N_18884);
nor U19387 (N_19387,N_19153,N_18533);
nand U19388 (N_19388,N_19082,N_18516);
xor U19389 (N_19389,N_18486,N_18963);
xnor U19390 (N_19390,N_18540,N_18479);
nand U19391 (N_19391,N_18532,N_18577);
nor U19392 (N_19392,N_18555,N_18691);
and U19393 (N_19393,N_18434,N_18441);
or U19394 (N_19394,N_18745,N_18591);
and U19395 (N_19395,N_18891,N_18414);
nor U19396 (N_19396,N_18992,N_18916);
and U19397 (N_19397,N_18675,N_18574);
and U19398 (N_19398,N_18913,N_18805);
or U19399 (N_19399,N_18636,N_19157);
and U19400 (N_19400,N_18606,N_18799);
nor U19401 (N_19401,N_18860,N_19196);
nor U19402 (N_19402,N_18834,N_18412);
and U19403 (N_19403,N_18831,N_19145);
or U19404 (N_19404,N_18528,N_18639);
or U19405 (N_19405,N_18698,N_18515);
xor U19406 (N_19406,N_18900,N_18704);
and U19407 (N_19407,N_19051,N_18699);
and U19408 (N_19408,N_18761,N_18904);
and U19409 (N_19409,N_18954,N_19095);
xnor U19410 (N_19410,N_18936,N_19050);
or U19411 (N_19411,N_18490,N_18838);
or U19412 (N_19412,N_19195,N_19141);
xnor U19413 (N_19413,N_18564,N_18796);
nand U19414 (N_19414,N_18857,N_18783);
nand U19415 (N_19415,N_18472,N_18687);
nor U19416 (N_19416,N_18897,N_18955);
xor U19417 (N_19417,N_18628,N_19191);
nor U19418 (N_19418,N_19012,N_19023);
xnor U19419 (N_19419,N_18489,N_18787);
and U19420 (N_19420,N_18422,N_18680);
nand U19421 (N_19421,N_19167,N_18962);
nor U19422 (N_19422,N_18609,N_18753);
and U19423 (N_19423,N_19057,N_19075);
and U19424 (N_19424,N_19072,N_18423);
or U19425 (N_19425,N_18711,N_19139);
nand U19426 (N_19426,N_18443,N_18596);
and U19427 (N_19427,N_18562,N_19014);
nor U19428 (N_19428,N_19120,N_18402);
xnor U19429 (N_19429,N_19156,N_18519);
and U19430 (N_19430,N_18426,N_18454);
nor U19431 (N_19431,N_18611,N_18640);
xnor U19432 (N_19432,N_19143,N_18548);
or U19433 (N_19433,N_18521,N_18623);
and U19434 (N_19434,N_18906,N_18679);
nor U19435 (N_19435,N_18481,N_18453);
nor U19436 (N_19436,N_18637,N_19056);
xnor U19437 (N_19437,N_18943,N_18880);
xnor U19438 (N_19438,N_18709,N_18452);
and U19439 (N_19439,N_18850,N_18809);
xor U19440 (N_19440,N_18966,N_18518);
nand U19441 (N_19441,N_18979,N_18602);
or U19442 (N_19442,N_19015,N_19179);
nor U19443 (N_19443,N_18828,N_18451);
nand U19444 (N_19444,N_18469,N_18447);
nor U19445 (N_19445,N_18986,N_18511);
nor U19446 (N_19446,N_18581,N_18536);
nand U19447 (N_19447,N_19030,N_18625);
nand U19448 (N_19448,N_18930,N_19162);
and U19449 (N_19449,N_18430,N_18400);
or U19450 (N_19450,N_18545,N_18587);
or U19451 (N_19451,N_18728,N_18988);
nor U19452 (N_19452,N_19058,N_18657);
xnor U19453 (N_19453,N_19052,N_18835);
xnor U19454 (N_19454,N_18840,N_18758);
xnor U19455 (N_19455,N_18820,N_19024);
xor U19456 (N_19456,N_18719,N_18554);
nand U19457 (N_19457,N_18734,N_18987);
nand U19458 (N_19458,N_18894,N_19192);
nor U19459 (N_19459,N_18819,N_18410);
nor U19460 (N_19460,N_19134,N_18870);
and U19461 (N_19461,N_18493,N_19081);
xor U19462 (N_19462,N_18612,N_19171);
nand U19463 (N_19463,N_19040,N_18547);
or U19464 (N_19464,N_19104,N_18427);
nand U19465 (N_19465,N_18542,N_18985);
nor U19466 (N_19466,N_18928,N_19013);
xor U19467 (N_19467,N_18660,N_19106);
nor U19468 (N_19468,N_18713,N_18785);
xnor U19469 (N_19469,N_18617,N_18858);
or U19470 (N_19470,N_18727,N_18411);
nand U19471 (N_19471,N_19181,N_19097);
xnor U19472 (N_19472,N_19066,N_18702);
nand U19473 (N_19473,N_18643,N_18926);
nor U19474 (N_19474,N_18918,N_19071);
xnor U19475 (N_19475,N_18568,N_18844);
nand U19476 (N_19476,N_18901,N_19146);
nand U19477 (N_19477,N_18664,N_19166);
nand U19478 (N_19478,N_18440,N_18567);
nand U19479 (N_19479,N_18588,N_19180);
or U19480 (N_19480,N_18851,N_18465);
xnor U19481 (N_19481,N_18551,N_18833);
nand U19482 (N_19482,N_18455,N_18632);
or U19483 (N_19483,N_18883,N_18837);
nand U19484 (N_19484,N_18801,N_18875);
nor U19485 (N_19485,N_19129,N_18859);
nor U19486 (N_19486,N_18659,N_18920);
xnor U19487 (N_19487,N_18615,N_18406);
and U19488 (N_19488,N_18726,N_18964);
nand U19489 (N_19489,N_18534,N_18717);
nand U19490 (N_19490,N_18627,N_18559);
xnor U19491 (N_19491,N_18989,N_18556);
and U19492 (N_19492,N_19089,N_19031);
xor U19493 (N_19493,N_18765,N_18624);
nand U19494 (N_19494,N_18775,N_18788);
nand U19495 (N_19495,N_19123,N_18579);
and U19496 (N_19496,N_18733,N_18669);
nor U19497 (N_19497,N_18737,N_18501);
nand U19498 (N_19498,N_18575,N_18965);
and U19499 (N_19499,N_19101,N_18947);
xor U19500 (N_19500,N_18731,N_18862);
xor U19501 (N_19501,N_19161,N_18517);
nor U19502 (N_19502,N_18417,N_18845);
nand U19503 (N_19503,N_18886,N_18890);
or U19504 (N_19504,N_19175,N_19032);
nand U19505 (N_19505,N_18692,N_18991);
or U19506 (N_19506,N_18824,N_18663);
nand U19507 (N_19507,N_19140,N_18777);
nand U19508 (N_19508,N_18941,N_18877);
and U19509 (N_19509,N_18908,N_18942);
nand U19510 (N_19510,N_19172,N_18967);
nor U19511 (N_19511,N_18957,N_18938);
or U19512 (N_19512,N_18652,N_18566);
xor U19513 (N_19513,N_18998,N_19100);
nor U19514 (N_19514,N_19131,N_19133);
nor U19515 (N_19515,N_18444,N_18825);
nor U19516 (N_19516,N_19090,N_19038);
nor U19517 (N_19517,N_18708,N_18509);
or U19518 (N_19518,N_18682,N_18802);
nand U19519 (N_19519,N_19150,N_18582);
and U19520 (N_19520,N_19197,N_18929);
nand U19521 (N_19521,N_18807,N_19126);
xnor U19522 (N_19522,N_19116,N_18576);
or U19523 (N_19523,N_19086,N_18565);
nand U19524 (N_19524,N_18456,N_18781);
and U19525 (N_19525,N_19002,N_18806);
or U19526 (N_19526,N_19160,N_19073);
and U19527 (N_19527,N_18642,N_18895);
xor U19528 (N_19528,N_19080,N_18863);
and U19529 (N_19529,N_18707,N_18804);
xor U19530 (N_19530,N_18520,N_18403);
and U19531 (N_19531,N_18683,N_19053);
nor U19532 (N_19532,N_19039,N_18909);
nor U19533 (N_19533,N_18585,N_19187);
nor U19534 (N_19534,N_18881,N_18793);
nand U19535 (N_19535,N_19017,N_19183);
nor U19536 (N_19536,N_18736,N_18466);
xnor U19537 (N_19537,N_18458,N_18794);
nor U19538 (N_19538,N_18996,N_18541);
nor U19539 (N_19539,N_18770,N_18896);
and U19540 (N_19540,N_18662,N_18635);
xnor U19541 (N_19541,N_18756,N_18599);
nor U19542 (N_19542,N_18984,N_18510);
or U19543 (N_19543,N_18855,N_18849);
or U19544 (N_19544,N_18953,N_19189);
nor U19545 (N_19545,N_18956,N_19034);
or U19546 (N_19546,N_18433,N_19047);
and U19547 (N_19547,N_18473,N_18999);
and U19548 (N_19548,N_18531,N_18513);
and U19549 (N_19549,N_18584,N_19077);
nor U19550 (N_19550,N_19173,N_18961);
nand U19551 (N_19551,N_18852,N_18595);
xnor U19552 (N_19552,N_19060,N_18503);
nor U19553 (N_19553,N_18438,N_18475);
or U19554 (N_19554,N_19163,N_18944);
and U19555 (N_19555,N_18415,N_19078);
nand U19556 (N_19556,N_18932,N_18912);
xnor U19557 (N_19557,N_18960,N_19117);
xor U19558 (N_19558,N_18404,N_18690);
or U19559 (N_19559,N_18507,N_18413);
nor U19560 (N_19560,N_18701,N_18654);
and U19561 (N_19561,N_18610,N_19061);
nand U19562 (N_19562,N_18821,N_18887);
and U19563 (N_19563,N_18866,N_18539);
nand U19564 (N_19564,N_18703,N_18522);
nand U19565 (N_19565,N_18893,N_18607);
and U19566 (N_19566,N_18485,N_18552);
xnor U19567 (N_19567,N_18505,N_19062);
nor U19568 (N_19568,N_19119,N_19079);
nand U19569 (N_19569,N_18524,N_19164);
nand U19570 (N_19570,N_19127,N_18905);
and U19571 (N_19571,N_19135,N_18700);
nor U19572 (N_19572,N_18471,N_18714);
or U19573 (N_19573,N_18827,N_18436);
nand U19574 (N_19574,N_18718,N_18725);
and U19575 (N_19575,N_18578,N_18598);
xnor U19576 (N_19576,N_18543,N_18848);
xnor U19577 (N_19577,N_18790,N_18464);
nand U19578 (N_19578,N_19098,N_18681);
and U19579 (N_19579,N_18597,N_19074);
nor U19580 (N_19580,N_18879,N_19125);
and U19581 (N_19581,N_18569,N_18463);
nor U19582 (N_19582,N_19083,N_19094);
nor U19583 (N_19583,N_18715,N_18722);
or U19584 (N_19584,N_18496,N_18557);
xnor U19585 (N_19585,N_18892,N_19084);
xor U19586 (N_19586,N_18786,N_18927);
nand U19587 (N_19587,N_18626,N_19063);
xnor U19588 (N_19588,N_19054,N_18487);
xor U19589 (N_19589,N_19159,N_18573);
xor U19590 (N_19590,N_18977,N_18502);
nand U19591 (N_19591,N_18689,N_18445);
or U19592 (N_19592,N_18457,N_18792);
nor U19593 (N_19593,N_18762,N_18461);
nand U19594 (N_19594,N_18950,N_18830);
nand U19595 (N_19595,N_18847,N_19070);
nor U19596 (N_19596,N_18571,N_18644);
and U19597 (N_19597,N_18872,N_18428);
nor U19598 (N_19598,N_18618,N_19178);
nor U19599 (N_19599,N_18649,N_18527);
or U19600 (N_19600,N_18891,N_19011);
or U19601 (N_19601,N_18780,N_19094);
or U19602 (N_19602,N_18529,N_18862);
or U19603 (N_19603,N_18820,N_19025);
or U19604 (N_19604,N_18547,N_18713);
and U19605 (N_19605,N_19125,N_18940);
nor U19606 (N_19606,N_18919,N_18845);
xor U19607 (N_19607,N_19157,N_19064);
or U19608 (N_19608,N_18700,N_18839);
and U19609 (N_19609,N_19126,N_18806);
xor U19610 (N_19610,N_18461,N_18418);
or U19611 (N_19611,N_19079,N_19104);
nand U19612 (N_19612,N_19164,N_18409);
and U19613 (N_19613,N_18569,N_18853);
xnor U19614 (N_19614,N_18618,N_18686);
or U19615 (N_19615,N_18681,N_18980);
xor U19616 (N_19616,N_19117,N_18827);
nand U19617 (N_19617,N_18534,N_18624);
nor U19618 (N_19618,N_19093,N_18646);
and U19619 (N_19619,N_18533,N_18829);
xnor U19620 (N_19620,N_18677,N_18835);
or U19621 (N_19621,N_19158,N_19008);
nand U19622 (N_19622,N_18866,N_18761);
or U19623 (N_19623,N_19009,N_18413);
xor U19624 (N_19624,N_18574,N_18538);
or U19625 (N_19625,N_18883,N_19152);
and U19626 (N_19626,N_18847,N_18601);
and U19627 (N_19627,N_19074,N_18436);
or U19628 (N_19628,N_19182,N_18665);
or U19629 (N_19629,N_18599,N_18598);
and U19630 (N_19630,N_18510,N_18427);
nand U19631 (N_19631,N_18500,N_18917);
or U19632 (N_19632,N_19055,N_18775);
nor U19633 (N_19633,N_18765,N_18437);
xnor U19634 (N_19634,N_18612,N_18722);
nand U19635 (N_19635,N_18958,N_18957);
nor U19636 (N_19636,N_18872,N_19012);
or U19637 (N_19637,N_18844,N_19045);
xnor U19638 (N_19638,N_18535,N_19085);
nand U19639 (N_19639,N_19120,N_18872);
xnor U19640 (N_19640,N_19150,N_18598);
xor U19641 (N_19641,N_18962,N_18536);
nand U19642 (N_19642,N_19131,N_19073);
nor U19643 (N_19643,N_18534,N_18507);
or U19644 (N_19644,N_18436,N_18412);
or U19645 (N_19645,N_18928,N_19194);
nor U19646 (N_19646,N_18496,N_19088);
xor U19647 (N_19647,N_19188,N_18456);
xnor U19648 (N_19648,N_19132,N_18968);
nor U19649 (N_19649,N_18567,N_19100);
and U19650 (N_19650,N_18891,N_18907);
or U19651 (N_19651,N_19170,N_18693);
and U19652 (N_19652,N_18764,N_18924);
xor U19653 (N_19653,N_18810,N_18692);
nand U19654 (N_19654,N_18648,N_18513);
or U19655 (N_19655,N_18627,N_18793);
or U19656 (N_19656,N_18676,N_19167);
nand U19657 (N_19657,N_18939,N_18772);
nand U19658 (N_19658,N_18690,N_19178);
nand U19659 (N_19659,N_19072,N_18501);
or U19660 (N_19660,N_18467,N_18848);
and U19661 (N_19661,N_18914,N_18943);
or U19662 (N_19662,N_18833,N_18532);
xnor U19663 (N_19663,N_18951,N_18517);
or U19664 (N_19664,N_18550,N_18424);
and U19665 (N_19665,N_19015,N_18749);
or U19666 (N_19666,N_19077,N_18939);
or U19667 (N_19667,N_19187,N_18419);
nand U19668 (N_19668,N_18775,N_18535);
or U19669 (N_19669,N_18981,N_18891);
nand U19670 (N_19670,N_18753,N_18970);
nor U19671 (N_19671,N_18511,N_18748);
and U19672 (N_19672,N_19034,N_19009);
xor U19673 (N_19673,N_18866,N_18481);
xnor U19674 (N_19674,N_18970,N_18684);
nor U19675 (N_19675,N_19071,N_18737);
nand U19676 (N_19676,N_18916,N_18668);
nand U19677 (N_19677,N_18512,N_18420);
nand U19678 (N_19678,N_18850,N_18568);
xnor U19679 (N_19679,N_19107,N_18629);
nand U19680 (N_19680,N_18733,N_19064);
or U19681 (N_19681,N_19061,N_18825);
xnor U19682 (N_19682,N_18646,N_18514);
and U19683 (N_19683,N_18919,N_18690);
and U19684 (N_19684,N_19110,N_18555);
nand U19685 (N_19685,N_19014,N_18942);
or U19686 (N_19686,N_18804,N_18693);
and U19687 (N_19687,N_18851,N_18755);
and U19688 (N_19688,N_18691,N_18857);
xor U19689 (N_19689,N_18944,N_18435);
nor U19690 (N_19690,N_18525,N_18561);
nand U19691 (N_19691,N_18835,N_19000);
nand U19692 (N_19692,N_18920,N_18868);
nor U19693 (N_19693,N_18594,N_18739);
xor U19694 (N_19694,N_18769,N_18846);
nand U19695 (N_19695,N_18649,N_18868);
nand U19696 (N_19696,N_19081,N_18816);
and U19697 (N_19697,N_18424,N_18444);
or U19698 (N_19698,N_18443,N_19024);
nand U19699 (N_19699,N_18537,N_19006);
nor U19700 (N_19700,N_18659,N_18868);
nand U19701 (N_19701,N_19003,N_19179);
nor U19702 (N_19702,N_19099,N_18539);
or U19703 (N_19703,N_19076,N_18790);
xor U19704 (N_19704,N_19061,N_18743);
and U19705 (N_19705,N_18832,N_18549);
xnor U19706 (N_19706,N_19199,N_18642);
or U19707 (N_19707,N_19181,N_18521);
xor U19708 (N_19708,N_18992,N_18716);
and U19709 (N_19709,N_19005,N_18473);
nand U19710 (N_19710,N_19055,N_19000);
nand U19711 (N_19711,N_18738,N_18840);
and U19712 (N_19712,N_18726,N_18822);
nand U19713 (N_19713,N_18615,N_18596);
or U19714 (N_19714,N_18828,N_18957);
nor U19715 (N_19715,N_18485,N_18472);
xor U19716 (N_19716,N_18681,N_18423);
xnor U19717 (N_19717,N_19167,N_19127);
xnor U19718 (N_19718,N_18406,N_18874);
and U19719 (N_19719,N_18705,N_18841);
and U19720 (N_19720,N_19158,N_19118);
xor U19721 (N_19721,N_18881,N_19191);
xor U19722 (N_19722,N_18411,N_18635);
xor U19723 (N_19723,N_18577,N_18991);
nor U19724 (N_19724,N_18430,N_18643);
or U19725 (N_19725,N_18602,N_19059);
nor U19726 (N_19726,N_18988,N_18413);
or U19727 (N_19727,N_18894,N_18940);
or U19728 (N_19728,N_19012,N_18940);
or U19729 (N_19729,N_18924,N_18720);
and U19730 (N_19730,N_19033,N_18867);
and U19731 (N_19731,N_18927,N_18402);
nor U19732 (N_19732,N_18939,N_18495);
or U19733 (N_19733,N_18717,N_18657);
nor U19734 (N_19734,N_18862,N_18866);
nor U19735 (N_19735,N_18448,N_18585);
xnor U19736 (N_19736,N_18663,N_19142);
and U19737 (N_19737,N_18937,N_18756);
nor U19738 (N_19738,N_18494,N_18448);
nor U19739 (N_19739,N_18615,N_18824);
and U19740 (N_19740,N_18647,N_19080);
or U19741 (N_19741,N_18414,N_18431);
xnor U19742 (N_19742,N_18549,N_18879);
nand U19743 (N_19743,N_19124,N_18968);
or U19744 (N_19744,N_18581,N_18548);
and U19745 (N_19745,N_18438,N_19006);
nor U19746 (N_19746,N_18892,N_18951);
or U19747 (N_19747,N_18440,N_18862);
nor U19748 (N_19748,N_18562,N_19137);
and U19749 (N_19749,N_18726,N_18469);
nor U19750 (N_19750,N_18708,N_18677);
nor U19751 (N_19751,N_18639,N_18507);
xnor U19752 (N_19752,N_18458,N_18492);
or U19753 (N_19753,N_18669,N_18564);
xor U19754 (N_19754,N_18726,N_18600);
nor U19755 (N_19755,N_18774,N_18795);
xnor U19756 (N_19756,N_18642,N_19046);
nand U19757 (N_19757,N_19188,N_18994);
and U19758 (N_19758,N_19121,N_19142);
or U19759 (N_19759,N_18867,N_18949);
xnor U19760 (N_19760,N_19162,N_18729);
nand U19761 (N_19761,N_18919,N_18467);
nand U19762 (N_19762,N_18406,N_19134);
nor U19763 (N_19763,N_18567,N_18824);
nand U19764 (N_19764,N_18942,N_18856);
xnor U19765 (N_19765,N_18903,N_18642);
nor U19766 (N_19766,N_18963,N_18736);
and U19767 (N_19767,N_19178,N_18738);
or U19768 (N_19768,N_18603,N_18892);
nor U19769 (N_19769,N_18452,N_18620);
xor U19770 (N_19770,N_19033,N_19040);
or U19771 (N_19771,N_18515,N_18751);
and U19772 (N_19772,N_18910,N_18957);
xnor U19773 (N_19773,N_19121,N_18699);
nor U19774 (N_19774,N_19107,N_18879);
nand U19775 (N_19775,N_18500,N_18852);
nor U19776 (N_19776,N_19051,N_18871);
nor U19777 (N_19777,N_18711,N_18719);
nand U19778 (N_19778,N_19017,N_19039);
or U19779 (N_19779,N_18413,N_18943);
xnor U19780 (N_19780,N_18852,N_19023);
xnor U19781 (N_19781,N_18814,N_18566);
nor U19782 (N_19782,N_18846,N_18596);
and U19783 (N_19783,N_18571,N_19034);
xnor U19784 (N_19784,N_18458,N_18956);
and U19785 (N_19785,N_18584,N_18872);
nand U19786 (N_19786,N_18737,N_19091);
xor U19787 (N_19787,N_18842,N_19083);
and U19788 (N_19788,N_19101,N_18635);
and U19789 (N_19789,N_18406,N_18828);
nand U19790 (N_19790,N_18476,N_18673);
xor U19791 (N_19791,N_18774,N_18507);
and U19792 (N_19792,N_18484,N_18407);
and U19793 (N_19793,N_18815,N_19021);
or U19794 (N_19794,N_19126,N_19029);
and U19795 (N_19795,N_18854,N_18673);
or U19796 (N_19796,N_19105,N_18814);
or U19797 (N_19797,N_18838,N_18452);
or U19798 (N_19798,N_18764,N_19156);
or U19799 (N_19799,N_18830,N_18438);
and U19800 (N_19800,N_18803,N_18593);
and U19801 (N_19801,N_18563,N_19103);
nor U19802 (N_19802,N_18644,N_18823);
xor U19803 (N_19803,N_19159,N_18971);
or U19804 (N_19804,N_18955,N_18899);
and U19805 (N_19805,N_18586,N_18763);
xor U19806 (N_19806,N_18410,N_18876);
nor U19807 (N_19807,N_18832,N_19082);
and U19808 (N_19808,N_18640,N_18974);
nor U19809 (N_19809,N_18592,N_18435);
xnor U19810 (N_19810,N_18722,N_19141);
nor U19811 (N_19811,N_19048,N_18416);
nand U19812 (N_19812,N_18679,N_18655);
nor U19813 (N_19813,N_18549,N_19155);
and U19814 (N_19814,N_18683,N_18500);
xor U19815 (N_19815,N_18916,N_19180);
or U19816 (N_19816,N_18523,N_19107);
and U19817 (N_19817,N_18685,N_18530);
and U19818 (N_19818,N_19152,N_18934);
xor U19819 (N_19819,N_18896,N_18908);
or U19820 (N_19820,N_18487,N_18611);
nand U19821 (N_19821,N_18738,N_19066);
or U19822 (N_19822,N_18970,N_18701);
xnor U19823 (N_19823,N_18433,N_18538);
and U19824 (N_19824,N_19092,N_18960);
and U19825 (N_19825,N_18729,N_19019);
xnor U19826 (N_19826,N_18511,N_18915);
and U19827 (N_19827,N_18485,N_19070);
and U19828 (N_19828,N_18729,N_18425);
xnor U19829 (N_19829,N_19047,N_18674);
xnor U19830 (N_19830,N_18754,N_18781);
nor U19831 (N_19831,N_18654,N_19084);
and U19832 (N_19832,N_19157,N_18808);
xor U19833 (N_19833,N_19133,N_18769);
nor U19834 (N_19834,N_18544,N_18991);
nor U19835 (N_19835,N_19011,N_19037);
xor U19836 (N_19836,N_19089,N_19095);
and U19837 (N_19837,N_18459,N_18443);
and U19838 (N_19838,N_18707,N_18679);
xnor U19839 (N_19839,N_19075,N_18996);
nor U19840 (N_19840,N_18789,N_18734);
xnor U19841 (N_19841,N_19085,N_19168);
nor U19842 (N_19842,N_18560,N_18803);
or U19843 (N_19843,N_19180,N_18624);
nand U19844 (N_19844,N_19145,N_18618);
nand U19845 (N_19845,N_18867,N_19023);
nand U19846 (N_19846,N_18997,N_19066);
or U19847 (N_19847,N_18584,N_19059);
nand U19848 (N_19848,N_18604,N_19078);
or U19849 (N_19849,N_18752,N_18422);
nor U19850 (N_19850,N_18407,N_18803);
and U19851 (N_19851,N_18876,N_18984);
nor U19852 (N_19852,N_18893,N_18575);
nand U19853 (N_19853,N_19056,N_18506);
nand U19854 (N_19854,N_18669,N_18843);
nand U19855 (N_19855,N_18569,N_18635);
and U19856 (N_19856,N_19011,N_18439);
and U19857 (N_19857,N_18418,N_18819);
or U19858 (N_19858,N_18707,N_18755);
nand U19859 (N_19859,N_18689,N_18901);
nand U19860 (N_19860,N_18952,N_18506);
nor U19861 (N_19861,N_18708,N_18908);
nor U19862 (N_19862,N_18838,N_18668);
nand U19863 (N_19863,N_18668,N_18751);
and U19864 (N_19864,N_18954,N_19107);
nor U19865 (N_19865,N_19115,N_18741);
nand U19866 (N_19866,N_18825,N_18923);
and U19867 (N_19867,N_18972,N_19117);
nand U19868 (N_19868,N_18980,N_18783);
or U19869 (N_19869,N_18549,N_18878);
xor U19870 (N_19870,N_19028,N_18428);
nand U19871 (N_19871,N_18820,N_18913);
nor U19872 (N_19872,N_18496,N_18956);
nand U19873 (N_19873,N_18768,N_19191);
nor U19874 (N_19874,N_18526,N_19195);
and U19875 (N_19875,N_19158,N_18666);
nand U19876 (N_19876,N_18979,N_18956);
xor U19877 (N_19877,N_18768,N_19108);
nor U19878 (N_19878,N_19040,N_19006);
or U19879 (N_19879,N_18942,N_18743);
nor U19880 (N_19880,N_19034,N_18830);
or U19881 (N_19881,N_18909,N_18720);
nor U19882 (N_19882,N_18513,N_18744);
nand U19883 (N_19883,N_18480,N_18986);
nor U19884 (N_19884,N_18679,N_18891);
and U19885 (N_19885,N_18905,N_18607);
xor U19886 (N_19886,N_18604,N_18405);
or U19887 (N_19887,N_18824,N_18675);
nand U19888 (N_19888,N_18559,N_18758);
nor U19889 (N_19889,N_19110,N_18983);
nor U19890 (N_19890,N_18557,N_18717);
or U19891 (N_19891,N_19142,N_18754);
and U19892 (N_19892,N_19052,N_18475);
or U19893 (N_19893,N_19000,N_18624);
nand U19894 (N_19894,N_18811,N_18649);
nand U19895 (N_19895,N_19099,N_19126);
or U19896 (N_19896,N_18438,N_18586);
or U19897 (N_19897,N_19111,N_19103);
nand U19898 (N_19898,N_18881,N_19177);
and U19899 (N_19899,N_18969,N_19094);
nor U19900 (N_19900,N_19074,N_18892);
and U19901 (N_19901,N_18413,N_18475);
xnor U19902 (N_19902,N_18935,N_18603);
and U19903 (N_19903,N_18590,N_18850);
nor U19904 (N_19904,N_19034,N_19109);
xnor U19905 (N_19905,N_19056,N_18733);
and U19906 (N_19906,N_19152,N_18730);
or U19907 (N_19907,N_18637,N_18935);
and U19908 (N_19908,N_19002,N_19084);
nand U19909 (N_19909,N_18671,N_18846);
nand U19910 (N_19910,N_18949,N_18464);
nand U19911 (N_19911,N_18773,N_18920);
xnor U19912 (N_19912,N_18467,N_19009);
or U19913 (N_19913,N_18859,N_19195);
nand U19914 (N_19914,N_18941,N_18516);
nor U19915 (N_19915,N_18829,N_18586);
xor U19916 (N_19916,N_18479,N_18513);
or U19917 (N_19917,N_18725,N_18644);
and U19918 (N_19918,N_19142,N_18734);
or U19919 (N_19919,N_19001,N_18802);
xnor U19920 (N_19920,N_18998,N_18655);
and U19921 (N_19921,N_19134,N_19103);
nor U19922 (N_19922,N_18527,N_19151);
and U19923 (N_19923,N_18647,N_18943);
nor U19924 (N_19924,N_18607,N_18407);
or U19925 (N_19925,N_18401,N_19167);
nand U19926 (N_19926,N_18970,N_18626);
xor U19927 (N_19927,N_19100,N_19081);
xor U19928 (N_19928,N_18616,N_18740);
nor U19929 (N_19929,N_18569,N_18717);
nor U19930 (N_19930,N_18747,N_18438);
xnor U19931 (N_19931,N_18645,N_19189);
or U19932 (N_19932,N_18514,N_18527);
and U19933 (N_19933,N_19146,N_19100);
xnor U19934 (N_19934,N_19054,N_18671);
and U19935 (N_19935,N_18815,N_18800);
or U19936 (N_19936,N_19173,N_18718);
nor U19937 (N_19937,N_18959,N_18695);
nor U19938 (N_19938,N_18806,N_18653);
nor U19939 (N_19939,N_18832,N_18821);
xor U19940 (N_19940,N_19198,N_18707);
xor U19941 (N_19941,N_18468,N_18927);
or U19942 (N_19942,N_18846,N_18885);
nor U19943 (N_19943,N_18803,N_18648);
and U19944 (N_19944,N_18599,N_18859);
and U19945 (N_19945,N_18909,N_18811);
nand U19946 (N_19946,N_18715,N_18569);
nand U19947 (N_19947,N_18792,N_18728);
nand U19948 (N_19948,N_18982,N_18427);
and U19949 (N_19949,N_18979,N_19029);
nor U19950 (N_19950,N_18906,N_19165);
xnor U19951 (N_19951,N_18517,N_18565);
or U19952 (N_19952,N_18929,N_18451);
and U19953 (N_19953,N_18851,N_18893);
and U19954 (N_19954,N_18496,N_18993);
xor U19955 (N_19955,N_18585,N_18525);
and U19956 (N_19956,N_18599,N_18544);
and U19957 (N_19957,N_18600,N_18482);
nor U19958 (N_19958,N_18993,N_18789);
and U19959 (N_19959,N_18784,N_18413);
or U19960 (N_19960,N_18452,N_18582);
xnor U19961 (N_19961,N_18995,N_19107);
nand U19962 (N_19962,N_18624,N_18637);
or U19963 (N_19963,N_18719,N_19087);
xnor U19964 (N_19964,N_19022,N_19136);
nand U19965 (N_19965,N_18778,N_19015);
xnor U19966 (N_19966,N_19065,N_18702);
or U19967 (N_19967,N_18538,N_19078);
xnor U19968 (N_19968,N_18595,N_18665);
or U19969 (N_19969,N_19019,N_18578);
or U19970 (N_19970,N_18494,N_18526);
nand U19971 (N_19971,N_19079,N_18485);
xnor U19972 (N_19972,N_18440,N_19146);
nor U19973 (N_19973,N_19186,N_18409);
xor U19974 (N_19974,N_18892,N_19118);
nand U19975 (N_19975,N_19158,N_18510);
and U19976 (N_19976,N_19147,N_19097);
or U19977 (N_19977,N_18704,N_18537);
nor U19978 (N_19978,N_18852,N_19150);
and U19979 (N_19979,N_18844,N_18713);
and U19980 (N_19980,N_18710,N_18523);
and U19981 (N_19981,N_18690,N_18710);
and U19982 (N_19982,N_18960,N_18573);
and U19983 (N_19983,N_19129,N_18867);
xnor U19984 (N_19984,N_19167,N_18838);
and U19985 (N_19985,N_18758,N_18885);
and U19986 (N_19986,N_18843,N_18556);
nor U19987 (N_19987,N_18977,N_18518);
or U19988 (N_19988,N_18528,N_18824);
nor U19989 (N_19989,N_18664,N_18546);
nor U19990 (N_19990,N_19085,N_18980);
xor U19991 (N_19991,N_18617,N_18574);
or U19992 (N_19992,N_18503,N_18909);
xor U19993 (N_19993,N_19152,N_19041);
and U19994 (N_19994,N_19145,N_18853);
or U19995 (N_19995,N_18745,N_18872);
nor U19996 (N_19996,N_19132,N_19184);
and U19997 (N_19997,N_18696,N_19002);
nor U19998 (N_19998,N_18987,N_18813);
nand U19999 (N_19999,N_18498,N_18613);
xor UO_0 (O_0,N_19492,N_19800);
and UO_1 (O_1,N_19560,N_19879);
nand UO_2 (O_2,N_19975,N_19786);
nor UO_3 (O_3,N_19547,N_19710);
xor UO_4 (O_4,N_19795,N_19214);
or UO_5 (O_5,N_19806,N_19954);
or UO_6 (O_6,N_19429,N_19421);
nor UO_7 (O_7,N_19290,N_19722);
nor UO_8 (O_8,N_19815,N_19706);
or UO_9 (O_9,N_19274,N_19759);
xor UO_10 (O_10,N_19714,N_19466);
and UO_11 (O_11,N_19976,N_19251);
nand UO_12 (O_12,N_19378,N_19310);
nor UO_13 (O_13,N_19713,N_19869);
nand UO_14 (O_14,N_19774,N_19955);
or UO_15 (O_15,N_19516,N_19600);
nand UO_16 (O_16,N_19269,N_19294);
and UO_17 (O_17,N_19902,N_19249);
xor UO_18 (O_18,N_19877,N_19458);
or UO_19 (O_19,N_19788,N_19674);
xor UO_20 (O_20,N_19809,N_19834);
nand UO_21 (O_21,N_19471,N_19632);
and UO_22 (O_22,N_19842,N_19283);
and UO_23 (O_23,N_19272,N_19338);
or UO_24 (O_24,N_19969,N_19947);
and UO_25 (O_25,N_19711,N_19704);
xor UO_26 (O_26,N_19320,N_19201);
nor UO_27 (O_27,N_19904,N_19811);
nand UO_28 (O_28,N_19716,N_19397);
xnor UO_29 (O_29,N_19921,N_19868);
xnor UO_30 (O_30,N_19991,N_19675);
nor UO_31 (O_31,N_19330,N_19723);
nor UO_32 (O_32,N_19607,N_19325);
nand UO_33 (O_33,N_19495,N_19237);
and UO_34 (O_34,N_19901,N_19460);
or UO_35 (O_35,N_19974,N_19321);
or UO_36 (O_36,N_19593,N_19410);
and UO_37 (O_37,N_19494,N_19745);
or UO_38 (O_38,N_19348,N_19878);
nand UO_39 (O_39,N_19768,N_19524);
nand UO_40 (O_40,N_19731,N_19477);
nand UO_41 (O_41,N_19452,N_19840);
xor UO_42 (O_42,N_19640,N_19635);
nand UO_43 (O_43,N_19379,N_19448);
and UO_44 (O_44,N_19864,N_19951);
nand UO_45 (O_45,N_19972,N_19944);
nand UO_46 (O_46,N_19934,N_19932);
nand UO_47 (O_47,N_19693,N_19771);
nor UO_48 (O_48,N_19555,N_19718);
nand UO_49 (O_49,N_19872,N_19803);
nand UO_50 (O_50,N_19823,N_19401);
nand UO_51 (O_51,N_19918,N_19487);
and UO_52 (O_52,N_19415,N_19246);
and UO_53 (O_53,N_19211,N_19435);
nor UO_54 (O_54,N_19529,N_19456);
xor UO_55 (O_55,N_19350,N_19522);
xor UO_56 (O_56,N_19651,N_19425);
nor UO_57 (O_57,N_19437,N_19681);
and UO_58 (O_58,N_19602,N_19644);
and UO_59 (O_59,N_19490,N_19993);
nor UO_60 (O_60,N_19850,N_19266);
nand UO_61 (O_61,N_19284,N_19942);
xnor UO_62 (O_62,N_19836,N_19796);
nor UO_63 (O_63,N_19373,N_19424);
nor UO_64 (O_64,N_19568,N_19948);
xor UO_65 (O_65,N_19531,N_19468);
and UO_66 (O_66,N_19318,N_19206);
nand UO_67 (O_67,N_19536,N_19573);
xor UO_68 (O_68,N_19608,N_19717);
or UO_69 (O_69,N_19370,N_19260);
and UO_70 (O_70,N_19790,N_19368);
and UO_71 (O_71,N_19941,N_19700);
and UO_72 (O_72,N_19474,N_19676);
or UO_73 (O_73,N_19994,N_19245);
and UO_74 (O_74,N_19347,N_19381);
or UO_75 (O_75,N_19375,N_19509);
and UO_76 (O_76,N_19553,N_19792);
or UO_77 (O_77,N_19292,N_19828);
nor UO_78 (O_78,N_19805,N_19386);
xnor UO_79 (O_79,N_19989,N_19682);
xnor UO_80 (O_80,N_19787,N_19758);
xnor UO_81 (O_81,N_19311,N_19414);
xor UO_82 (O_82,N_19739,N_19626);
and UO_83 (O_83,N_19478,N_19364);
or UO_84 (O_84,N_19735,N_19256);
xor UO_85 (O_85,N_19352,N_19654);
nand UO_86 (O_86,N_19689,N_19849);
or UO_87 (O_87,N_19688,N_19286);
or UO_88 (O_88,N_19857,N_19209);
or UO_89 (O_89,N_19899,N_19239);
nand UO_90 (O_90,N_19990,N_19469);
nand UO_91 (O_91,N_19807,N_19883);
nand UO_92 (O_92,N_19562,N_19226);
nor UO_93 (O_93,N_19761,N_19252);
nor UO_94 (O_94,N_19817,N_19846);
or UO_95 (O_95,N_19876,N_19585);
nand UO_96 (O_96,N_19963,N_19845);
nor UO_97 (O_97,N_19216,N_19413);
nor UO_98 (O_98,N_19754,N_19481);
nor UO_99 (O_99,N_19746,N_19264);
nand UO_100 (O_100,N_19223,N_19724);
and UO_101 (O_101,N_19219,N_19257);
nand UO_102 (O_102,N_19627,N_19865);
and UO_103 (O_103,N_19721,N_19960);
and UO_104 (O_104,N_19971,N_19804);
xor UO_105 (O_105,N_19664,N_19848);
and UO_106 (O_106,N_19979,N_19491);
nand UO_107 (O_107,N_19326,N_19574);
xnor UO_108 (O_108,N_19314,N_19765);
and UO_109 (O_109,N_19485,N_19762);
nand UO_110 (O_110,N_19694,N_19207);
nand UO_111 (O_111,N_19785,N_19210);
nor UO_112 (O_112,N_19416,N_19299);
nor UO_113 (O_113,N_19521,N_19821);
or UO_114 (O_114,N_19406,N_19799);
xor UO_115 (O_115,N_19958,N_19659);
nand UO_116 (O_116,N_19578,N_19645);
nand UO_117 (O_117,N_19383,N_19298);
and UO_118 (O_118,N_19905,N_19978);
nor UO_119 (O_119,N_19484,N_19698);
or UO_120 (O_120,N_19512,N_19952);
nand UO_121 (O_121,N_19808,N_19451);
and UO_122 (O_122,N_19480,N_19405);
xnor UO_123 (O_123,N_19241,N_19690);
xor UO_124 (O_124,N_19819,N_19599);
xor UO_125 (O_125,N_19967,N_19550);
and UO_126 (O_126,N_19692,N_19331);
xnor UO_127 (O_127,N_19833,N_19885);
nor UO_128 (O_128,N_19319,N_19404);
nand UO_129 (O_129,N_19212,N_19891);
xnor UO_130 (O_130,N_19570,N_19623);
and UO_131 (O_131,N_19534,N_19229);
nor UO_132 (O_132,N_19440,N_19365);
and UO_133 (O_133,N_19605,N_19385);
nor UO_134 (O_134,N_19510,N_19647);
xor UO_135 (O_135,N_19295,N_19986);
xnor UO_136 (O_136,N_19747,N_19797);
and UO_137 (O_137,N_19566,N_19648);
nor UO_138 (O_138,N_19327,N_19699);
nand UO_139 (O_139,N_19956,N_19501);
xor UO_140 (O_140,N_19341,N_19767);
and UO_141 (O_141,N_19473,N_19686);
nand UO_142 (O_142,N_19613,N_19500);
nor UO_143 (O_143,N_19793,N_19650);
nor UO_144 (O_144,N_19464,N_19371);
or UO_145 (O_145,N_19679,N_19225);
nor UO_146 (O_146,N_19467,N_19893);
and UO_147 (O_147,N_19832,N_19380);
and UO_148 (O_148,N_19399,N_19741);
or UO_149 (O_149,N_19625,N_19384);
and UO_150 (O_150,N_19366,N_19263);
and UO_151 (O_151,N_19233,N_19995);
or UO_152 (O_152,N_19776,N_19489);
xnor UO_153 (O_153,N_19445,N_19393);
and UO_154 (O_154,N_19657,N_19772);
xnor UO_155 (O_155,N_19581,N_19888);
nor UO_156 (O_156,N_19459,N_19367);
nand UO_157 (O_157,N_19691,N_19996);
nand UO_158 (O_158,N_19506,N_19557);
nor UO_159 (O_159,N_19323,N_19820);
nand UO_160 (O_160,N_19454,N_19420);
xnor UO_161 (O_161,N_19461,N_19518);
nor UO_162 (O_162,N_19496,N_19400);
or UO_163 (O_163,N_19537,N_19580);
nor UO_164 (O_164,N_19436,N_19230);
or UO_165 (O_165,N_19544,N_19752);
xor UO_166 (O_166,N_19369,N_19929);
or UO_167 (O_167,N_19822,N_19356);
and UO_168 (O_168,N_19503,N_19288);
xnor UO_169 (O_169,N_19303,N_19927);
or UO_170 (O_170,N_19712,N_19535);
nor UO_171 (O_171,N_19403,N_19950);
or UO_172 (O_172,N_19488,N_19359);
and UO_173 (O_173,N_19228,N_19411);
nand UO_174 (O_174,N_19614,N_19514);
nor UO_175 (O_175,N_19422,N_19353);
nor UO_176 (O_176,N_19344,N_19910);
nor UO_177 (O_177,N_19276,N_19897);
nor UO_178 (O_178,N_19998,N_19639);
nor UO_179 (O_179,N_19619,N_19438);
and UO_180 (O_180,N_19680,N_19838);
xnor UO_181 (O_181,N_19390,N_19360);
or UO_182 (O_182,N_19753,N_19582);
or UO_183 (O_183,N_19913,N_19250);
and UO_184 (O_184,N_19248,N_19672);
xor UO_185 (O_185,N_19965,N_19882);
nand UO_186 (O_186,N_19511,N_19351);
xor UO_187 (O_187,N_19419,N_19825);
xor UO_188 (O_188,N_19577,N_19707);
xor UO_189 (O_189,N_19813,N_19982);
or UO_190 (O_190,N_19742,N_19336);
or UO_191 (O_191,N_19446,N_19668);
xnor UO_192 (O_192,N_19928,N_19592);
nor UO_193 (O_193,N_19894,N_19280);
nand UO_194 (O_194,N_19520,N_19637);
or UO_195 (O_195,N_19775,N_19935);
nor UO_196 (O_196,N_19427,N_19638);
xor UO_197 (O_197,N_19236,N_19621);
nor UO_198 (O_198,N_19434,N_19200);
and UO_199 (O_199,N_19727,N_19282);
nand UO_200 (O_200,N_19204,N_19428);
or UO_201 (O_201,N_19636,N_19423);
xnor UO_202 (O_202,N_19202,N_19609);
nand UO_203 (O_203,N_19830,N_19355);
or UO_204 (O_204,N_19695,N_19285);
or UO_205 (O_205,N_19242,N_19728);
nand UO_206 (O_206,N_19296,N_19983);
nand UO_207 (O_207,N_19527,N_19579);
or UO_208 (O_208,N_19238,N_19870);
nand UO_209 (O_209,N_19729,N_19827);
or UO_210 (O_210,N_19784,N_19392);
xnor UO_211 (O_211,N_19791,N_19541);
or UO_212 (O_212,N_19773,N_19755);
xor UO_213 (O_213,N_19685,N_19253);
and UO_214 (O_214,N_19539,N_19760);
nor UO_215 (O_215,N_19549,N_19309);
nand UO_216 (O_216,N_19778,N_19985);
xor UO_217 (O_217,N_19439,N_19814);
nand UO_218 (O_218,N_19559,N_19715);
and UO_219 (O_219,N_19205,N_19673);
nand UO_220 (O_220,N_19981,N_19662);
and UO_221 (O_221,N_19583,N_19751);
nor UO_222 (O_222,N_19757,N_19231);
nor UO_223 (O_223,N_19395,N_19855);
and UO_224 (O_224,N_19628,N_19328);
nand UO_225 (O_225,N_19919,N_19943);
and UO_226 (O_226,N_19222,N_19709);
nor UO_227 (O_227,N_19262,N_19633);
nor UO_228 (O_228,N_19930,N_19641);
and UO_229 (O_229,N_19572,N_19702);
nor UO_230 (O_230,N_19258,N_19620);
and UO_231 (O_231,N_19959,N_19208);
nand UO_232 (O_232,N_19987,N_19507);
or UO_233 (O_233,N_19970,N_19243);
or UO_234 (O_234,N_19270,N_19756);
nand UO_235 (O_235,N_19586,N_19515);
xnor UO_236 (O_236,N_19218,N_19543);
or UO_237 (O_237,N_19312,N_19701);
or UO_238 (O_238,N_19346,N_19508);
nor UO_239 (O_239,N_19844,N_19734);
nand UO_240 (O_240,N_19293,N_19660);
nand UO_241 (O_241,N_19275,N_19431);
xor UO_242 (O_242,N_19340,N_19781);
nand UO_243 (O_243,N_19780,N_19234);
nand UO_244 (O_244,N_19387,N_19629);
and UO_245 (O_245,N_19497,N_19665);
nor UO_246 (O_246,N_19801,N_19961);
nor UO_247 (O_247,N_19450,N_19271);
or UO_248 (O_248,N_19462,N_19615);
xnor UO_249 (O_249,N_19217,N_19906);
and UO_250 (O_250,N_19412,N_19343);
and UO_251 (O_251,N_19281,N_19875);
and UO_252 (O_252,N_19931,N_19442);
nor UO_253 (O_253,N_19277,N_19743);
and UO_254 (O_254,N_19576,N_19307);
xnor UO_255 (O_255,N_19337,N_19333);
and UO_256 (O_256,N_19213,N_19453);
nor UO_257 (O_257,N_19377,N_19839);
nand UO_258 (O_258,N_19601,N_19766);
nand UO_259 (O_259,N_19925,N_19584);
or UO_260 (O_260,N_19357,N_19953);
and UO_261 (O_261,N_19342,N_19279);
and UO_262 (O_262,N_19505,N_19939);
xor UO_263 (O_263,N_19733,N_19308);
xor UO_264 (O_264,N_19575,N_19265);
or UO_265 (O_265,N_19661,N_19854);
xnor UO_266 (O_266,N_19802,N_19306);
nand UO_267 (O_267,N_19376,N_19499);
and UO_268 (O_268,N_19254,N_19908);
xor UO_269 (O_269,N_19587,N_19777);
xor UO_270 (O_270,N_19523,N_19703);
or UO_271 (O_271,N_19618,N_19968);
xnor UO_272 (O_272,N_19443,N_19203);
and UO_273 (O_273,N_19977,N_19730);
nand UO_274 (O_274,N_19432,N_19949);
nand UO_275 (O_275,N_19726,N_19880);
xor UO_276 (O_276,N_19402,N_19571);
nand UO_277 (O_277,N_19598,N_19890);
nor UO_278 (O_278,N_19551,N_19548);
and UO_279 (O_279,N_19862,N_19687);
xnor UO_280 (O_280,N_19558,N_19297);
xor UO_281 (O_281,N_19671,N_19914);
xnor UO_282 (O_282,N_19565,N_19361);
nor UO_283 (O_283,N_19519,N_19389);
or UO_284 (O_284,N_19291,N_19493);
or UO_285 (O_285,N_19606,N_19988);
xnor UO_286 (O_286,N_19391,N_19569);
and UO_287 (O_287,N_19643,N_19881);
and UO_288 (O_288,N_19358,N_19737);
or UO_289 (O_289,N_19540,N_19267);
nor UO_290 (O_290,N_19938,N_19426);
nand UO_291 (O_291,N_19259,N_19289);
or UO_292 (O_292,N_19964,N_19653);
or UO_293 (O_293,N_19235,N_19398);
xor UO_294 (O_294,N_19533,N_19696);
or UO_295 (O_295,N_19907,N_19324);
nand UO_296 (O_296,N_19463,N_19447);
xor UO_297 (O_297,N_19273,N_19764);
xnor UO_298 (O_298,N_19911,N_19526);
xnor UO_299 (O_299,N_19596,N_19818);
nand UO_300 (O_300,N_19980,N_19268);
xor UO_301 (O_301,N_19433,N_19455);
xor UO_302 (O_302,N_19334,N_19634);
nand UO_303 (O_303,N_19750,N_19457);
xnor UO_304 (O_304,N_19604,N_19313);
nor UO_305 (O_305,N_19532,N_19973);
nand UO_306 (O_306,N_19232,N_19962);
nor UO_307 (O_307,N_19669,N_19740);
nand UO_308 (O_308,N_19349,N_19444);
xnor UO_309 (O_309,N_19867,N_19603);
and UO_310 (O_310,N_19597,N_19418);
nand UO_311 (O_311,N_19920,N_19486);
or UO_312 (O_312,N_19915,N_19677);
nand UO_313 (O_313,N_19957,N_19316);
nor UO_314 (O_314,N_19590,N_19382);
or UO_315 (O_315,N_19530,N_19705);
nand UO_316 (O_316,N_19831,N_19545);
nor UO_317 (O_317,N_19221,N_19912);
xnor UO_318 (O_318,N_19683,N_19903);
xnor UO_319 (O_319,N_19656,N_19999);
nor UO_320 (O_320,N_19917,N_19502);
nand UO_321 (O_321,N_19564,N_19852);
and UO_322 (O_322,N_19826,N_19517);
nor UO_323 (O_323,N_19220,N_19887);
and UO_324 (O_324,N_19305,N_19525);
nand UO_325 (O_325,N_19892,N_19616);
nor UO_326 (O_326,N_19354,N_19430);
nand UO_327 (O_327,N_19475,N_19997);
nor UO_328 (O_328,N_19898,N_19538);
and UO_329 (O_329,N_19372,N_19789);
or UO_330 (O_330,N_19317,N_19749);
nor UO_331 (O_331,N_19362,N_19984);
nand UO_332 (O_332,N_19720,N_19363);
xnor UO_333 (O_333,N_19240,N_19856);
xnor UO_334 (O_334,N_19224,N_19546);
nand UO_335 (O_335,N_19874,N_19738);
nor UO_336 (O_336,N_19816,N_19652);
and UO_337 (O_337,N_19649,N_19926);
nor UO_338 (O_338,N_19498,N_19812);
and UO_339 (O_339,N_19227,N_19417);
xnor UO_340 (O_340,N_19782,N_19923);
and UO_341 (O_341,N_19678,N_19591);
nand UO_342 (O_342,N_19895,N_19708);
and UO_343 (O_343,N_19630,N_19408);
nor UO_344 (O_344,N_19472,N_19339);
nor UO_345 (O_345,N_19829,N_19663);
or UO_346 (O_346,N_19909,N_19642);
xor UO_347 (O_347,N_19937,N_19837);
xnor UO_348 (O_348,N_19924,N_19933);
nor UO_349 (O_349,N_19824,N_19631);
or UO_350 (O_350,N_19563,N_19900);
xor UO_351 (O_351,N_19396,N_19810);
nor UO_352 (O_352,N_19302,N_19301);
nor UO_353 (O_353,N_19732,N_19287);
xor UO_354 (O_354,N_19847,N_19783);
and UO_355 (O_355,N_19769,N_19884);
or UO_356 (O_356,N_19940,N_19278);
nand UO_357 (O_357,N_19896,N_19871);
xor UO_358 (O_358,N_19247,N_19407);
xor UO_359 (O_359,N_19483,N_19851);
and UO_360 (O_360,N_19770,N_19561);
and UO_361 (O_361,N_19394,N_19779);
xor UO_362 (O_362,N_19589,N_19858);
xor UO_363 (O_363,N_19345,N_19843);
xor UO_364 (O_364,N_19992,N_19866);
nand UO_365 (O_365,N_19889,N_19859);
nand UO_366 (O_366,N_19835,N_19315);
nor UO_367 (O_367,N_19215,N_19255);
or UO_368 (O_368,N_19666,N_19610);
nand UO_369 (O_369,N_19528,N_19617);
nand UO_370 (O_370,N_19863,N_19655);
and UO_371 (O_371,N_19465,N_19595);
xor UO_372 (O_372,N_19322,N_19725);
nand UO_373 (O_373,N_19946,N_19886);
and UO_374 (O_374,N_19476,N_19513);
nor UO_375 (O_375,N_19261,N_19794);
nand UO_376 (O_376,N_19861,N_19335);
nand UO_377 (O_377,N_19853,N_19374);
and UO_378 (O_378,N_19860,N_19658);
xor UO_379 (O_379,N_19622,N_19482);
or UO_380 (O_380,N_19763,N_19684);
and UO_381 (O_381,N_19646,N_19966);
xnor UO_382 (O_382,N_19449,N_19556);
xor UO_383 (O_383,N_19922,N_19697);
and UO_384 (O_384,N_19744,N_19504);
xor UO_385 (O_385,N_19304,N_19612);
xor UO_386 (O_386,N_19542,N_19594);
nand UO_387 (O_387,N_19554,N_19945);
nor UO_388 (O_388,N_19332,N_19588);
nor UO_389 (O_389,N_19719,N_19552);
xor UO_390 (O_390,N_19329,N_19388);
nand UO_391 (O_391,N_19748,N_19441);
and UO_392 (O_392,N_19873,N_19916);
nor UO_393 (O_393,N_19409,N_19798);
xnor UO_394 (O_394,N_19841,N_19670);
nor UO_395 (O_395,N_19936,N_19736);
nand UO_396 (O_396,N_19244,N_19470);
and UO_397 (O_397,N_19611,N_19667);
and UO_398 (O_398,N_19300,N_19567);
and UO_399 (O_399,N_19624,N_19479);
or UO_400 (O_400,N_19799,N_19355);
nand UO_401 (O_401,N_19961,N_19441);
nand UO_402 (O_402,N_19494,N_19628);
and UO_403 (O_403,N_19866,N_19224);
xnor UO_404 (O_404,N_19386,N_19898);
xor UO_405 (O_405,N_19310,N_19886);
nand UO_406 (O_406,N_19518,N_19690);
xnor UO_407 (O_407,N_19766,N_19218);
nor UO_408 (O_408,N_19612,N_19241);
xor UO_409 (O_409,N_19605,N_19283);
nor UO_410 (O_410,N_19714,N_19339);
xor UO_411 (O_411,N_19614,N_19523);
and UO_412 (O_412,N_19352,N_19915);
and UO_413 (O_413,N_19325,N_19910);
or UO_414 (O_414,N_19501,N_19459);
xor UO_415 (O_415,N_19702,N_19680);
and UO_416 (O_416,N_19583,N_19235);
nand UO_417 (O_417,N_19829,N_19478);
nand UO_418 (O_418,N_19457,N_19460);
nand UO_419 (O_419,N_19224,N_19390);
xor UO_420 (O_420,N_19239,N_19290);
and UO_421 (O_421,N_19677,N_19525);
and UO_422 (O_422,N_19978,N_19789);
nand UO_423 (O_423,N_19996,N_19707);
nor UO_424 (O_424,N_19633,N_19953);
xnor UO_425 (O_425,N_19841,N_19333);
xor UO_426 (O_426,N_19760,N_19844);
xor UO_427 (O_427,N_19708,N_19494);
or UO_428 (O_428,N_19998,N_19981);
nand UO_429 (O_429,N_19209,N_19464);
or UO_430 (O_430,N_19748,N_19511);
and UO_431 (O_431,N_19614,N_19659);
and UO_432 (O_432,N_19796,N_19866);
and UO_433 (O_433,N_19419,N_19475);
and UO_434 (O_434,N_19496,N_19976);
xor UO_435 (O_435,N_19559,N_19908);
nand UO_436 (O_436,N_19423,N_19776);
nor UO_437 (O_437,N_19898,N_19394);
nand UO_438 (O_438,N_19997,N_19984);
and UO_439 (O_439,N_19698,N_19486);
xor UO_440 (O_440,N_19353,N_19472);
or UO_441 (O_441,N_19917,N_19773);
or UO_442 (O_442,N_19847,N_19951);
and UO_443 (O_443,N_19972,N_19780);
xor UO_444 (O_444,N_19349,N_19609);
or UO_445 (O_445,N_19845,N_19985);
or UO_446 (O_446,N_19309,N_19377);
nor UO_447 (O_447,N_19625,N_19987);
nor UO_448 (O_448,N_19562,N_19952);
and UO_449 (O_449,N_19946,N_19811);
and UO_450 (O_450,N_19604,N_19606);
or UO_451 (O_451,N_19454,N_19721);
nor UO_452 (O_452,N_19296,N_19776);
or UO_453 (O_453,N_19274,N_19436);
nand UO_454 (O_454,N_19798,N_19226);
and UO_455 (O_455,N_19461,N_19598);
nand UO_456 (O_456,N_19318,N_19419);
nor UO_457 (O_457,N_19871,N_19307);
xnor UO_458 (O_458,N_19643,N_19557);
xor UO_459 (O_459,N_19666,N_19335);
or UO_460 (O_460,N_19985,N_19521);
xor UO_461 (O_461,N_19285,N_19515);
and UO_462 (O_462,N_19374,N_19267);
nor UO_463 (O_463,N_19265,N_19959);
or UO_464 (O_464,N_19417,N_19679);
nand UO_465 (O_465,N_19615,N_19497);
or UO_466 (O_466,N_19629,N_19512);
or UO_467 (O_467,N_19842,N_19334);
and UO_468 (O_468,N_19606,N_19844);
or UO_469 (O_469,N_19889,N_19712);
nand UO_470 (O_470,N_19463,N_19802);
nor UO_471 (O_471,N_19523,N_19826);
or UO_472 (O_472,N_19530,N_19527);
nand UO_473 (O_473,N_19686,N_19454);
nand UO_474 (O_474,N_19530,N_19565);
xor UO_475 (O_475,N_19377,N_19863);
nor UO_476 (O_476,N_19943,N_19426);
nor UO_477 (O_477,N_19674,N_19489);
nor UO_478 (O_478,N_19619,N_19766);
or UO_479 (O_479,N_19711,N_19900);
nand UO_480 (O_480,N_19322,N_19541);
or UO_481 (O_481,N_19325,N_19455);
nand UO_482 (O_482,N_19558,N_19612);
or UO_483 (O_483,N_19979,N_19789);
and UO_484 (O_484,N_19812,N_19464);
nand UO_485 (O_485,N_19326,N_19477);
xor UO_486 (O_486,N_19945,N_19932);
and UO_487 (O_487,N_19433,N_19676);
nand UO_488 (O_488,N_19334,N_19462);
nor UO_489 (O_489,N_19743,N_19273);
xor UO_490 (O_490,N_19729,N_19890);
nand UO_491 (O_491,N_19482,N_19663);
nor UO_492 (O_492,N_19215,N_19752);
nor UO_493 (O_493,N_19448,N_19830);
nor UO_494 (O_494,N_19869,N_19376);
or UO_495 (O_495,N_19294,N_19668);
nor UO_496 (O_496,N_19559,N_19938);
nor UO_497 (O_497,N_19398,N_19361);
nor UO_498 (O_498,N_19258,N_19707);
nor UO_499 (O_499,N_19908,N_19256);
and UO_500 (O_500,N_19478,N_19220);
and UO_501 (O_501,N_19566,N_19249);
nand UO_502 (O_502,N_19900,N_19574);
or UO_503 (O_503,N_19706,N_19840);
xor UO_504 (O_504,N_19701,N_19499);
xor UO_505 (O_505,N_19718,N_19768);
xor UO_506 (O_506,N_19721,N_19213);
or UO_507 (O_507,N_19743,N_19340);
nand UO_508 (O_508,N_19942,N_19852);
nand UO_509 (O_509,N_19747,N_19992);
or UO_510 (O_510,N_19431,N_19588);
or UO_511 (O_511,N_19856,N_19619);
or UO_512 (O_512,N_19469,N_19959);
nand UO_513 (O_513,N_19859,N_19524);
nand UO_514 (O_514,N_19848,N_19533);
and UO_515 (O_515,N_19635,N_19838);
nor UO_516 (O_516,N_19438,N_19502);
xnor UO_517 (O_517,N_19870,N_19558);
xor UO_518 (O_518,N_19966,N_19624);
and UO_519 (O_519,N_19266,N_19387);
or UO_520 (O_520,N_19315,N_19323);
and UO_521 (O_521,N_19828,N_19765);
and UO_522 (O_522,N_19564,N_19559);
or UO_523 (O_523,N_19269,N_19502);
or UO_524 (O_524,N_19542,N_19925);
and UO_525 (O_525,N_19664,N_19678);
xnor UO_526 (O_526,N_19757,N_19497);
xor UO_527 (O_527,N_19739,N_19574);
xnor UO_528 (O_528,N_19529,N_19680);
nand UO_529 (O_529,N_19651,N_19501);
nand UO_530 (O_530,N_19630,N_19853);
and UO_531 (O_531,N_19303,N_19275);
xor UO_532 (O_532,N_19326,N_19573);
xor UO_533 (O_533,N_19428,N_19829);
or UO_534 (O_534,N_19677,N_19777);
or UO_535 (O_535,N_19952,N_19699);
nand UO_536 (O_536,N_19974,N_19484);
or UO_537 (O_537,N_19544,N_19330);
xor UO_538 (O_538,N_19634,N_19279);
and UO_539 (O_539,N_19246,N_19648);
xor UO_540 (O_540,N_19651,N_19421);
xor UO_541 (O_541,N_19743,N_19357);
xor UO_542 (O_542,N_19552,N_19415);
and UO_543 (O_543,N_19209,N_19815);
xnor UO_544 (O_544,N_19353,N_19486);
and UO_545 (O_545,N_19385,N_19300);
and UO_546 (O_546,N_19729,N_19517);
nor UO_547 (O_547,N_19431,N_19962);
nor UO_548 (O_548,N_19654,N_19455);
nor UO_549 (O_549,N_19416,N_19533);
or UO_550 (O_550,N_19714,N_19845);
xor UO_551 (O_551,N_19970,N_19822);
or UO_552 (O_552,N_19317,N_19720);
nand UO_553 (O_553,N_19363,N_19222);
or UO_554 (O_554,N_19221,N_19787);
and UO_555 (O_555,N_19324,N_19777);
or UO_556 (O_556,N_19950,N_19220);
and UO_557 (O_557,N_19933,N_19541);
nor UO_558 (O_558,N_19757,N_19675);
and UO_559 (O_559,N_19543,N_19288);
xor UO_560 (O_560,N_19549,N_19590);
xnor UO_561 (O_561,N_19645,N_19867);
nand UO_562 (O_562,N_19636,N_19510);
nand UO_563 (O_563,N_19421,N_19851);
and UO_564 (O_564,N_19434,N_19259);
nand UO_565 (O_565,N_19677,N_19735);
or UO_566 (O_566,N_19800,N_19844);
nor UO_567 (O_567,N_19840,N_19417);
nor UO_568 (O_568,N_19554,N_19490);
nand UO_569 (O_569,N_19587,N_19992);
and UO_570 (O_570,N_19610,N_19494);
and UO_571 (O_571,N_19993,N_19529);
nor UO_572 (O_572,N_19386,N_19452);
or UO_573 (O_573,N_19624,N_19584);
nor UO_574 (O_574,N_19820,N_19699);
xor UO_575 (O_575,N_19373,N_19295);
nand UO_576 (O_576,N_19666,N_19544);
and UO_577 (O_577,N_19573,N_19594);
xnor UO_578 (O_578,N_19789,N_19619);
nand UO_579 (O_579,N_19608,N_19471);
nand UO_580 (O_580,N_19560,N_19841);
or UO_581 (O_581,N_19946,N_19209);
nand UO_582 (O_582,N_19976,N_19340);
or UO_583 (O_583,N_19559,N_19613);
nand UO_584 (O_584,N_19408,N_19462);
nor UO_585 (O_585,N_19961,N_19489);
xnor UO_586 (O_586,N_19932,N_19698);
and UO_587 (O_587,N_19540,N_19791);
and UO_588 (O_588,N_19802,N_19410);
nand UO_589 (O_589,N_19837,N_19538);
xnor UO_590 (O_590,N_19534,N_19407);
or UO_591 (O_591,N_19256,N_19694);
nand UO_592 (O_592,N_19342,N_19775);
or UO_593 (O_593,N_19512,N_19736);
nand UO_594 (O_594,N_19884,N_19837);
nor UO_595 (O_595,N_19840,N_19988);
and UO_596 (O_596,N_19888,N_19419);
nor UO_597 (O_597,N_19763,N_19657);
and UO_598 (O_598,N_19413,N_19617);
xor UO_599 (O_599,N_19306,N_19747);
and UO_600 (O_600,N_19700,N_19589);
nor UO_601 (O_601,N_19202,N_19622);
xor UO_602 (O_602,N_19664,N_19879);
xnor UO_603 (O_603,N_19985,N_19367);
xor UO_604 (O_604,N_19509,N_19229);
nor UO_605 (O_605,N_19310,N_19587);
or UO_606 (O_606,N_19213,N_19948);
nor UO_607 (O_607,N_19375,N_19533);
xor UO_608 (O_608,N_19664,N_19302);
or UO_609 (O_609,N_19737,N_19758);
or UO_610 (O_610,N_19234,N_19714);
xnor UO_611 (O_611,N_19291,N_19831);
nor UO_612 (O_612,N_19277,N_19850);
or UO_613 (O_613,N_19733,N_19979);
nor UO_614 (O_614,N_19726,N_19488);
and UO_615 (O_615,N_19969,N_19442);
nor UO_616 (O_616,N_19570,N_19405);
or UO_617 (O_617,N_19903,N_19861);
and UO_618 (O_618,N_19591,N_19919);
nor UO_619 (O_619,N_19626,N_19214);
nor UO_620 (O_620,N_19765,N_19916);
and UO_621 (O_621,N_19855,N_19856);
nor UO_622 (O_622,N_19606,N_19778);
or UO_623 (O_623,N_19257,N_19865);
or UO_624 (O_624,N_19327,N_19263);
nand UO_625 (O_625,N_19543,N_19763);
nor UO_626 (O_626,N_19858,N_19688);
and UO_627 (O_627,N_19445,N_19825);
or UO_628 (O_628,N_19774,N_19964);
nand UO_629 (O_629,N_19671,N_19975);
and UO_630 (O_630,N_19648,N_19497);
xor UO_631 (O_631,N_19947,N_19945);
nand UO_632 (O_632,N_19205,N_19677);
nand UO_633 (O_633,N_19739,N_19526);
or UO_634 (O_634,N_19841,N_19399);
nor UO_635 (O_635,N_19904,N_19589);
and UO_636 (O_636,N_19936,N_19464);
or UO_637 (O_637,N_19329,N_19464);
and UO_638 (O_638,N_19726,N_19627);
nand UO_639 (O_639,N_19992,N_19403);
nand UO_640 (O_640,N_19620,N_19511);
nand UO_641 (O_641,N_19320,N_19343);
xor UO_642 (O_642,N_19237,N_19439);
xor UO_643 (O_643,N_19388,N_19438);
or UO_644 (O_644,N_19401,N_19209);
nor UO_645 (O_645,N_19485,N_19258);
and UO_646 (O_646,N_19714,N_19272);
xnor UO_647 (O_647,N_19990,N_19897);
and UO_648 (O_648,N_19652,N_19952);
xnor UO_649 (O_649,N_19978,N_19880);
or UO_650 (O_650,N_19789,N_19792);
nor UO_651 (O_651,N_19489,N_19405);
nor UO_652 (O_652,N_19520,N_19901);
or UO_653 (O_653,N_19376,N_19205);
xor UO_654 (O_654,N_19308,N_19809);
nor UO_655 (O_655,N_19211,N_19523);
nand UO_656 (O_656,N_19233,N_19926);
nand UO_657 (O_657,N_19794,N_19737);
nand UO_658 (O_658,N_19629,N_19227);
or UO_659 (O_659,N_19867,N_19512);
xnor UO_660 (O_660,N_19541,N_19749);
or UO_661 (O_661,N_19758,N_19521);
or UO_662 (O_662,N_19290,N_19962);
nor UO_663 (O_663,N_19433,N_19462);
nor UO_664 (O_664,N_19638,N_19667);
and UO_665 (O_665,N_19756,N_19487);
or UO_666 (O_666,N_19911,N_19978);
xnor UO_667 (O_667,N_19302,N_19689);
nor UO_668 (O_668,N_19466,N_19500);
or UO_669 (O_669,N_19302,N_19757);
or UO_670 (O_670,N_19979,N_19247);
nand UO_671 (O_671,N_19820,N_19490);
or UO_672 (O_672,N_19237,N_19420);
xor UO_673 (O_673,N_19556,N_19973);
or UO_674 (O_674,N_19849,N_19442);
or UO_675 (O_675,N_19368,N_19597);
xnor UO_676 (O_676,N_19851,N_19744);
nand UO_677 (O_677,N_19812,N_19784);
nor UO_678 (O_678,N_19749,N_19379);
xor UO_679 (O_679,N_19467,N_19551);
nand UO_680 (O_680,N_19406,N_19984);
or UO_681 (O_681,N_19783,N_19618);
xnor UO_682 (O_682,N_19636,N_19668);
xor UO_683 (O_683,N_19306,N_19783);
xnor UO_684 (O_684,N_19982,N_19313);
nor UO_685 (O_685,N_19495,N_19470);
and UO_686 (O_686,N_19689,N_19719);
or UO_687 (O_687,N_19734,N_19889);
xor UO_688 (O_688,N_19375,N_19720);
and UO_689 (O_689,N_19747,N_19705);
xnor UO_690 (O_690,N_19631,N_19505);
nand UO_691 (O_691,N_19537,N_19870);
and UO_692 (O_692,N_19754,N_19756);
or UO_693 (O_693,N_19941,N_19881);
nand UO_694 (O_694,N_19236,N_19721);
and UO_695 (O_695,N_19637,N_19652);
or UO_696 (O_696,N_19508,N_19921);
or UO_697 (O_697,N_19743,N_19383);
nor UO_698 (O_698,N_19547,N_19324);
nor UO_699 (O_699,N_19466,N_19896);
nand UO_700 (O_700,N_19673,N_19641);
nand UO_701 (O_701,N_19552,N_19240);
or UO_702 (O_702,N_19561,N_19442);
nand UO_703 (O_703,N_19864,N_19230);
xor UO_704 (O_704,N_19485,N_19203);
and UO_705 (O_705,N_19503,N_19813);
nor UO_706 (O_706,N_19917,N_19259);
nor UO_707 (O_707,N_19930,N_19337);
nor UO_708 (O_708,N_19450,N_19433);
nand UO_709 (O_709,N_19777,N_19434);
xor UO_710 (O_710,N_19348,N_19391);
nand UO_711 (O_711,N_19634,N_19830);
and UO_712 (O_712,N_19203,N_19517);
nor UO_713 (O_713,N_19295,N_19743);
nand UO_714 (O_714,N_19251,N_19997);
or UO_715 (O_715,N_19502,N_19723);
nor UO_716 (O_716,N_19779,N_19536);
nand UO_717 (O_717,N_19316,N_19512);
nor UO_718 (O_718,N_19326,N_19899);
nor UO_719 (O_719,N_19817,N_19842);
nand UO_720 (O_720,N_19542,N_19780);
xor UO_721 (O_721,N_19631,N_19314);
nor UO_722 (O_722,N_19554,N_19648);
nor UO_723 (O_723,N_19868,N_19801);
and UO_724 (O_724,N_19453,N_19482);
nand UO_725 (O_725,N_19453,N_19889);
xnor UO_726 (O_726,N_19259,N_19221);
and UO_727 (O_727,N_19632,N_19823);
or UO_728 (O_728,N_19604,N_19951);
or UO_729 (O_729,N_19347,N_19630);
xor UO_730 (O_730,N_19298,N_19873);
or UO_731 (O_731,N_19788,N_19491);
xnor UO_732 (O_732,N_19503,N_19441);
or UO_733 (O_733,N_19390,N_19278);
nor UO_734 (O_734,N_19235,N_19481);
xor UO_735 (O_735,N_19604,N_19303);
xor UO_736 (O_736,N_19656,N_19486);
and UO_737 (O_737,N_19968,N_19202);
nor UO_738 (O_738,N_19855,N_19838);
nand UO_739 (O_739,N_19234,N_19858);
nand UO_740 (O_740,N_19246,N_19932);
nand UO_741 (O_741,N_19330,N_19898);
xor UO_742 (O_742,N_19941,N_19850);
or UO_743 (O_743,N_19300,N_19856);
or UO_744 (O_744,N_19982,N_19629);
nand UO_745 (O_745,N_19759,N_19221);
or UO_746 (O_746,N_19597,N_19523);
xnor UO_747 (O_747,N_19575,N_19222);
or UO_748 (O_748,N_19687,N_19858);
and UO_749 (O_749,N_19864,N_19963);
xor UO_750 (O_750,N_19612,N_19867);
xnor UO_751 (O_751,N_19246,N_19279);
nand UO_752 (O_752,N_19305,N_19492);
nand UO_753 (O_753,N_19955,N_19780);
and UO_754 (O_754,N_19487,N_19667);
nor UO_755 (O_755,N_19350,N_19467);
nor UO_756 (O_756,N_19662,N_19466);
or UO_757 (O_757,N_19595,N_19408);
xnor UO_758 (O_758,N_19810,N_19785);
nand UO_759 (O_759,N_19660,N_19200);
or UO_760 (O_760,N_19589,N_19698);
or UO_761 (O_761,N_19591,N_19740);
nand UO_762 (O_762,N_19247,N_19850);
and UO_763 (O_763,N_19250,N_19838);
or UO_764 (O_764,N_19861,N_19997);
xor UO_765 (O_765,N_19625,N_19514);
and UO_766 (O_766,N_19857,N_19575);
xor UO_767 (O_767,N_19815,N_19861);
or UO_768 (O_768,N_19431,N_19673);
nand UO_769 (O_769,N_19472,N_19897);
and UO_770 (O_770,N_19425,N_19244);
nor UO_771 (O_771,N_19425,N_19496);
or UO_772 (O_772,N_19871,N_19351);
nor UO_773 (O_773,N_19269,N_19908);
nand UO_774 (O_774,N_19422,N_19213);
nand UO_775 (O_775,N_19519,N_19267);
or UO_776 (O_776,N_19257,N_19548);
xnor UO_777 (O_777,N_19318,N_19902);
or UO_778 (O_778,N_19651,N_19895);
and UO_779 (O_779,N_19441,N_19553);
nor UO_780 (O_780,N_19288,N_19638);
and UO_781 (O_781,N_19331,N_19744);
and UO_782 (O_782,N_19563,N_19728);
and UO_783 (O_783,N_19686,N_19737);
or UO_784 (O_784,N_19443,N_19722);
xnor UO_785 (O_785,N_19939,N_19294);
nand UO_786 (O_786,N_19606,N_19560);
and UO_787 (O_787,N_19570,N_19855);
and UO_788 (O_788,N_19906,N_19258);
nor UO_789 (O_789,N_19744,N_19329);
and UO_790 (O_790,N_19450,N_19252);
and UO_791 (O_791,N_19561,N_19443);
nor UO_792 (O_792,N_19946,N_19945);
xor UO_793 (O_793,N_19584,N_19768);
xor UO_794 (O_794,N_19332,N_19850);
or UO_795 (O_795,N_19742,N_19952);
or UO_796 (O_796,N_19498,N_19861);
xnor UO_797 (O_797,N_19954,N_19638);
or UO_798 (O_798,N_19593,N_19238);
nand UO_799 (O_799,N_19469,N_19479);
nand UO_800 (O_800,N_19565,N_19661);
nor UO_801 (O_801,N_19331,N_19992);
or UO_802 (O_802,N_19623,N_19416);
nand UO_803 (O_803,N_19335,N_19764);
and UO_804 (O_804,N_19254,N_19537);
and UO_805 (O_805,N_19545,N_19700);
nand UO_806 (O_806,N_19802,N_19787);
nand UO_807 (O_807,N_19646,N_19463);
and UO_808 (O_808,N_19292,N_19612);
nand UO_809 (O_809,N_19285,N_19900);
and UO_810 (O_810,N_19219,N_19824);
or UO_811 (O_811,N_19369,N_19463);
xor UO_812 (O_812,N_19794,N_19399);
or UO_813 (O_813,N_19502,N_19248);
and UO_814 (O_814,N_19766,N_19846);
and UO_815 (O_815,N_19495,N_19866);
or UO_816 (O_816,N_19945,N_19878);
nand UO_817 (O_817,N_19876,N_19806);
nand UO_818 (O_818,N_19387,N_19813);
nand UO_819 (O_819,N_19676,N_19324);
and UO_820 (O_820,N_19774,N_19861);
and UO_821 (O_821,N_19889,N_19336);
and UO_822 (O_822,N_19642,N_19357);
nor UO_823 (O_823,N_19294,N_19681);
nor UO_824 (O_824,N_19763,N_19267);
nor UO_825 (O_825,N_19398,N_19632);
nor UO_826 (O_826,N_19218,N_19958);
xnor UO_827 (O_827,N_19393,N_19770);
and UO_828 (O_828,N_19217,N_19350);
xor UO_829 (O_829,N_19606,N_19610);
nor UO_830 (O_830,N_19593,N_19866);
xor UO_831 (O_831,N_19710,N_19766);
nand UO_832 (O_832,N_19860,N_19557);
nor UO_833 (O_833,N_19588,N_19258);
or UO_834 (O_834,N_19261,N_19582);
xor UO_835 (O_835,N_19872,N_19383);
nand UO_836 (O_836,N_19857,N_19943);
nand UO_837 (O_837,N_19518,N_19263);
xnor UO_838 (O_838,N_19327,N_19679);
xor UO_839 (O_839,N_19683,N_19812);
nor UO_840 (O_840,N_19946,N_19314);
and UO_841 (O_841,N_19751,N_19318);
nor UO_842 (O_842,N_19353,N_19936);
nand UO_843 (O_843,N_19667,N_19493);
nand UO_844 (O_844,N_19253,N_19293);
and UO_845 (O_845,N_19537,N_19968);
or UO_846 (O_846,N_19617,N_19574);
xor UO_847 (O_847,N_19583,N_19272);
or UO_848 (O_848,N_19845,N_19534);
xnor UO_849 (O_849,N_19500,N_19789);
or UO_850 (O_850,N_19267,N_19737);
nor UO_851 (O_851,N_19621,N_19359);
nor UO_852 (O_852,N_19669,N_19968);
xor UO_853 (O_853,N_19448,N_19988);
or UO_854 (O_854,N_19432,N_19267);
xor UO_855 (O_855,N_19631,N_19372);
or UO_856 (O_856,N_19867,N_19660);
xnor UO_857 (O_857,N_19810,N_19353);
xor UO_858 (O_858,N_19520,N_19585);
or UO_859 (O_859,N_19430,N_19499);
or UO_860 (O_860,N_19941,N_19679);
and UO_861 (O_861,N_19897,N_19258);
or UO_862 (O_862,N_19578,N_19217);
xnor UO_863 (O_863,N_19618,N_19729);
xor UO_864 (O_864,N_19254,N_19732);
nand UO_865 (O_865,N_19587,N_19527);
and UO_866 (O_866,N_19542,N_19462);
or UO_867 (O_867,N_19859,N_19968);
xor UO_868 (O_868,N_19610,N_19667);
xnor UO_869 (O_869,N_19813,N_19792);
xor UO_870 (O_870,N_19586,N_19995);
xnor UO_871 (O_871,N_19204,N_19526);
nor UO_872 (O_872,N_19932,N_19241);
xor UO_873 (O_873,N_19539,N_19579);
xor UO_874 (O_874,N_19597,N_19332);
nand UO_875 (O_875,N_19649,N_19626);
xnor UO_876 (O_876,N_19753,N_19837);
nor UO_877 (O_877,N_19642,N_19212);
xor UO_878 (O_878,N_19304,N_19736);
xnor UO_879 (O_879,N_19392,N_19731);
or UO_880 (O_880,N_19853,N_19504);
and UO_881 (O_881,N_19416,N_19786);
nor UO_882 (O_882,N_19794,N_19898);
or UO_883 (O_883,N_19335,N_19891);
and UO_884 (O_884,N_19360,N_19579);
nor UO_885 (O_885,N_19909,N_19730);
and UO_886 (O_886,N_19856,N_19295);
xor UO_887 (O_887,N_19775,N_19518);
or UO_888 (O_888,N_19230,N_19297);
nor UO_889 (O_889,N_19213,N_19391);
or UO_890 (O_890,N_19361,N_19335);
or UO_891 (O_891,N_19501,N_19502);
or UO_892 (O_892,N_19920,N_19515);
xor UO_893 (O_893,N_19959,N_19358);
and UO_894 (O_894,N_19645,N_19463);
or UO_895 (O_895,N_19632,N_19680);
and UO_896 (O_896,N_19543,N_19911);
nand UO_897 (O_897,N_19527,N_19827);
or UO_898 (O_898,N_19940,N_19273);
nand UO_899 (O_899,N_19212,N_19609);
xnor UO_900 (O_900,N_19773,N_19423);
or UO_901 (O_901,N_19987,N_19869);
nor UO_902 (O_902,N_19878,N_19305);
xnor UO_903 (O_903,N_19634,N_19958);
xor UO_904 (O_904,N_19862,N_19695);
or UO_905 (O_905,N_19492,N_19286);
and UO_906 (O_906,N_19992,N_19677);
nand UO_907 (O_907,N_19840,N_19805);
or UO_908 (O_908,N_19539,N_19463);
and UO_909 (O_909,N_19491,N_19272);
or UO_910 (O_910,N_19905,N_19259);
nor UO_911 (O_911,N_19563,N_19237);
nor UO_912 (O_912,N_19690,N_19921);
nor UO_913 (O_913,N_19268,N_19535);
nand UO_914 (O_914,N_19596,N_19335);
nor UO_915 (O_915,N_19904,N_19289);
and UO_916 (O_916,N_19299,N_19497);
nor UO_917 (O_917,N_19577,N_19239);
nand UO_918 (O_918,N_19591,N_19292);
xnor UO_919 (O_919,N_19901,N_19884);
or UO_920 (O_920,N_19319,N_19911);
or UO_921 (O_921,N_19582,N_19749);
xor UO_922 (O_922,N_19794,N_19697);
nor UO_923 (O_923,N_19325,N_19790);
nand UO_924 (O_924,N_19391,N_19555);
nand UO_925 (O_925,N_19854,N_19718);
and UO_926 (O_926,N_19399,N_19720);
or UO_927 (O_927,N_19308,N_19901);
or UO_928 (O_928,N_19205,N_19980);
and UO_929 (O_929,N_19777,N_19439);
or UO_930 (O_930,N_19764,N_19813);
and UO_931 (O_931,N_19835,N_19747);
or UO_932 (O_932,N_19650,N_19918);
xor UO_933 (O_933,N_19245,N_19894);
nand UO_934 (O_934,N_19546,N_19547);
or UO_935 (O_935,N_19649,N_19204);
and UO_936 (O_936,N_19365,N_19844);
or UO_937 (O_937,N_19417,N_19411);
and UO_938 (O_938,N_19392,N_19458);
xnor UO_939 (O_939,N_19542,N_19236);
and UO_940 (O_940,N_19687,N_19217);
nor UO_941 (O_941,N_19833,N_19970);
xor UO_942 (O_942,N_19761,N_19563);
nor UO_943 (O_943,N_19573,N_19247);
and UO_944 (O_944,N_19925,N_19945);
or UO_945 (O_945,N_19653,N_19839);
nand UO_946 (O_946,N_19734,N_19504);
xnor UO_947 (O_947,N_19269,N_19434);
and UO_948 (O_948,N_19446,N_19482);
and UO_949 (O_949,N_19722,N_19237);
or UO_950 (O_950,N_19610,N_19225);
xnor UO_951 (O_951,N_19904,N_19701);
nor UO_952 (O_952,N_19314,N_19509);
and UO_953 (O_953,N_19202,N_19517);
nor UO_954 (O_954,N_19550,N_19359);
xnor UO_955 (O_955,N_19586,N_19938);
nand UO_956 (O_956,N_19778,N_19252);
nor UO_957 (O_957,N_19870,N_19756);
or UO_958 (O_958,N_19815,N_19819);
or UO_959 (O_959,N_19407,N_19774);
or UO_960 (O_960,N_19317,N_19654);
xor UO_961 (O_961,N_19497,N_19565);
nand UO_962 (O_962,N_19781,N_19299);
or UO_963 (O_963,N_19459,N_19589);
nand UO_964 (O_964,N_19884,N_19922);
nand UO_965 (O_965,N_19542,N_19600);
xnor UO_966 (O_966,N_19218,N_19367);
xnor UO_967 (O_967,N_19885,N_19579);
or UO_968 (O_968,N_19420,N_19825);
nand UO_969 (O_969,N_19344,N_19817);
xnor UO_970 (O_970,N_19675,N_19609);
xnor UO_971 (O_971,N_19785,N_19649);
and UO_972 (O_972,N_19678,N_19634);
nor UO_973 (O_973,N_19843,N_19632);
or UO_974 (O_974,N_19572,N_19631);
xor UO_975 (O_975,N_19933,N_19949);
and UO_976 (O_976,N_19617,N_19787);
nor UO_977 (O_977,N_19233,N_19824);
xor UO_978 (O_978,N_19322,N_19343);
and UO_979 (O_979,N_19897,N_19829);
xnor UO_980 (O_980,N_19838,N_19717);
nand UO_981 (O_981,N_19327,N_19902);
and UO_982 (O_982,N_19327,N_19806);
nand UO_983 (O_983,N_19493,N_19633);
and UO_984 (O_984,N_19302,N_19232);
or UO_985 (O_985,N_19258,N_19301);
xor UO_986 (O_986,N_19587,N_19905);
xnor UO_987 (O_987,N_19576,N_19553);
nand UO_988 (O_988,N_19382,N_19480);
xor UO_989 (O_989,N_19679,N_19501);
and UO_990 (O_990,N_19211,N_19743);
or UO_991 (O_991,N_19277,N_19608);
xor UO_992 (O_992,N_19246,N_19971);
or UO_993 (O_993,N_19265,N_19876);
and UO_994 (O_994,N_19931,N_19667);
and UO_995 (O_995,N_19610,N_19354);
and UO_996 (O_996,N_19355,N_19997);
or UO_997 (O_997,N_19979,N_19760);
nor UO_998 (O_998,N_19458,N_19360);
xnor UO_999 (O_999,N_19995,N_19372);
and UO_1000 (O_1000,N_19651,N_19704);
nor UO_1001 (O_1001,N_19358,N_19581);
nor UO_1002 (O_1002,N_19571,N_19415);
nand UO_1003 (O_1003,N_19278,N_19365);
nor UO_1004 (O_1004,N_19621,N_19813);
nor UO_1005 (O_1005,N_19724,N_19462);
and UO_1006 (O_1006,N_19923,N_19382);
xnor UO_1007 (O_1007,N_19718,N_19981);
nor UO_1008 (O_1008,N_19615,N_19748);
nand UO_1009 (O_1009,N_19905,N_19275);
nand UO_1010 (O_1010,N_19908,N_19941);
nand UO_1011 (O_1011,N_19591,N_19893);
or UO_1012 (O_1012,N_19951,N_19933);
or UO_1013 (O_1013,N_19385,N_19343);
nor UO_1014 (O_1014,N_19275,N_19268);
and UO_1015 (O_1015,N_19510,N_19936);
or UO_1016 (O_1016,N_19468,N_19802);
and UO_1017 (O_1017,N_19401,N_19908);
nand UO_1018 (O_1018,N_19223,N_19645);
nor UO_1019 (O_1019,N_19892,N_19347);
or UO_1020 (O_1020,N_19621,N_19273);
nand UO_1021 (O_1021,N_19648,N_19351);
or UO_1022 (O_1022,N_19673,N_19499);
or UO_1023 (O_1023,N_19376,N_19862);
and UO_1024 (O_1024,N_19610,N_19333);
nor UO_1025 (O_1025,N_19352,N_19834);
nor UO_1026 (O_1026,N_19928,N_19258);
nor UO_1027 (O_1027,N_19954,N_19939);
xor UO_1028 (O_1028,N_19416,N_19353);
or UO_1029 (O_1029,N_19871,N_19580);
nand UO_1030 (O_1030,N_19258,N_19323);
nand UO_1031 (O_1031,N_19241,N_19688);
xnor UO_1032 (O_1032,N_19609,N_19794);
nand UO_1033 (O_1033,N_19261,N_19737);
and UO_1034 (O_1034,N_19819,N_19852);
nor UO_1035 (O_1035,N_19795,N_19763);
nand UO_1036 (O_1036,N_19598,N_19294);
or UO_1037 (O_1037,N_19312,N_19874);
nor UO_1038 (O_1038,N_19999,N_19372);
and UO_1039 (O_1039,N_19323,N_19327);
nand UO_1040 (O_1040,N_19935,N_19553);
or UO_1041 (O_1041,N_19597,N_19381);
and UO_1042 (O_1042,N_19516,N_19332);
nand UO_1043 (O_1043,N_19647,N_19504);
xnor UO_1044 (O_1044,N_19323,N_19350);
xor UO_1045 (O_1045,N_19682,N_19420);
nor UO_1046 (O_1046,N_19328,N_19563);
or UO_1047 (O_1047,N_19852,N_19296);
and UO_1048 (O_1048,N_19870,N_19730);
and UO_1049 (O_1049,N_19503,N_19328);
nor UO_1050 (O_1050,N_19603,N_19406);
xor UO_1051 (O_1051,N_19543,N_19861);
nor UO_1052 (O_1052,N_19475,N_19762);
xnor UO_1053 (O_1053,N_19881,N_19207);
nand UO_1054 (O_1054,N_19446,N_19297);
xnor UO_1055 (O_1055,N_19201,N_19277);
nor UO_1056 (O_1056,N_19420,N_19210);
nand UO_1057 (O_1057,N_19566,N_19727);
nor UO_1058 (O_1058,N_19606,N_19794);
xnor UO_1059 (O_1059,N_19854,N_19393);
or UO_1060 (O_1060,N_19423,N_19583);
or UO_1061 (O_1061,N_19499,N_19285);
nor UO_1062 (O_1062,N_19601,N_19553);
nand UO_1063 (O_1063,N_19824,N_19945);
or UO_1064 (O_1064,N_19795,N_19938);
or UO_1065 (O_1065,N_19705,N_19388);
and UO_1066 (O_1066,N_19653,N_19704);
xnor UO_1067 (O_1067,N_19618,N_19857);
and UO_1068 (O_1068,N_19305,N_19760);
xor UO_1069 (O_1069,N_19916,N_19679);
and UO_1070 (O_1070,N_19752,N_19971);
xnor UO_1071 (O_1071,N_19656,N_19848);
nor UO_1072 (O_1072,N_19710,N_19673);
or UO_1073 (O_1073,N_19509,N_19203);
xor UO_1074 (O_1074,N_19770,N_19650);
and UO_1075 (O_1075,N_19898,N_19353);
nand UO_1076 (O_1076,N_19423,N_19879);
or UO_1077 (O_1077,N_19532,N_19252);
xnor UO_1078 (O_1078,N_19775,N_19315);
and UO_1079 (O_1079,N_19332,N_19557);
xnor UO_1080 (O_1080,N_19343,N_19707);
nand UO_1081 (O_1081,N_19898,N_19492);
and UO_1082 (O_1082,N_19578,N_19338);
nand UO_1083 (O_1083,N_19343,N_19839);
or UO_1084 (O_1084,N_19598,N_19460);
nor UO_1085 (O_1085,N_19392,N_19762);
or UO_1086 (O_1086,N_19881,N_19839);
or UO_1087 (O_1087,N_19881,N_19515);
xnor UO_1088 (O_1088,N_19884,N_19820);
and UO_1089 (O_1089,N_19649,N_19730);
xnor UO_1090 (O_1090,N_19904,N_19395);
nand UO_1091 (O_1091,N_19880,N_19276);
nor UO_1092 (O_1092,N_19272,N_19728);
and UO_1093 (O_1093,N_19909,N_19285);
xnor UO_1094 (O_1094,N_19247,N_19209);
xor UO_1095 (O_1095,N_19376,N_19588);
nor UO_1096 (O_1096,N_19650,N_19312);
and UO_1097 (O_1097,N_19881,N_19523);
or UO_1098 (O_1098,N_19392,N_19326);
and UO_1099 (O_1099,N_19730,N_19838);
and UO_1100 (O_1100,N_19803,N_19564);
and UO_1101 (O_1101,N_19825,N_19348);
nor UO_1102 (O_1102,N_19703,N_19234);
nor UO_1103 (O_1103,N_19803,N_19805);
or UO_1104 (O_1104,N_19222,N_19392);
nor UO_1105 (O_1105,N_19256,N_19224);
xnor UO_1106 (O_1106,N_19446,N_19983);
or UO_1107 (O_1107,N_19847,N_19639);
or UO_1108 (O_1108,N_19933,N_19707);
nor UO_1109 (O_1109,N_19764,N_19350);
nand UO_1110 (O_1110,N_19818,N_19927);
and UO_1111 (O_1111,N_19748,N_19297);
and UO_1112 (O_1112,N_19343,N_19441);
xor UO_1113 (O_1113,N_19537,N_19452);
nand UO_1114 (O_1114,N_19300,N_19648);
xnor UO_1115 (O_1115,N_19793,N_19826);
and UO_1116 (O_1116,N_19245,N_19978);
nor UO_1117 (O_1117,N_19822,N_19911);
xor UO_1118 (O_1118,N_19634,N_19494);
or UO_1119 (O_1119,N_19767,N_19908);
nand UO_1120 (O_1120,N_19241,N_19284);
or UO_1121 (O_1121,N_19561,N_19226);
nand UO_1122 (O_1122,N_19612,N_19875);
and UO_1123 (O_1123,N_19823,N_19578);
xor UO_1124 (O_1124,N_19406,N_19521);
nand UO_1125 (O_1125,N_19999,N_19929);
nand UO_1126 (O_1126,N_19297,N_19249);
and UO_1127 (O_1127,N_19537,N_19592);
nor UO_1128 (O_1128,N_19649,N_19477);
xnor UO_1129 (O_1129,N_19768,N_19252);
nand UO_1130 (O_1130,N_19872,N_19980);
xnor UO_1131 (O_1131,N_19653,N_19639);
xnor UO_1132 (O_1132,N_19712,N_19357);
and UO_1133 (O_1133,N_19978,N_19714);
nand UO_1134 (O_1134,N_19868,N_19533);
or UO_1135 (O_1135,N_19205,N_19447);
nand UO_1136 (O_1136,N_19301,N_19519);
nor UO_1137 (O_1137,N_19348,N_19708);
xnor UO_1138 (O_1138,N_19485,N_19464);
nor UO_1139 (O_1139,N_19700,N_19656);
nor UO_1140 (O_1140,N_19224,N_19845);
xor UO_1141 (O_1141,N_19770,N_19624);
nand UO_1142 (O_1142,N_19412,N_19441);
and UO_1143 (O_1143,N_19845,N_19216);
and UO_1144 (O_1144,N_19797,N_19754);
nor UO_1145 (O_1145,N_19672,N_19372);
nand UO_1146 (O_1146,N_19410,N_19942);
nand UO_1147 (O_1147,N_19959,N_19723);
nor UO_1148 (O_1148,N_19358,N_19775);
nand UO_1149 (O_1149,N_19833,N_19567);
and UO_1150 (O_1150,N_19757,N_19645);
xnor UO_1151 (O_1151,N_19849,N_19411);
nor UO_1152 (O_1152,N_19949,N_19320);
nor UO_1153 (O_1153,N_19889,N_19742);
or UO_1154 (O_1154,N_19314,N_19928);
nor UO_1155 (O_1155,N_19574,N_19747);
nand UO_1156 (O_1156,N_19625,N_19369);
and UO_1157 (O_1157,N_19811,N_19685);
and UO_1158 (O_1158,N_19997,N_19686);
and UO_1159 (O_1159,N_19258,N_19842);
and UO_1160 (O_1160,N_19289,N_19716);
nand UO_1161 (O_1161,N_19628,N_19875);
xnor UO_1162 (O_1162,N_19635,N_19893);
and UO_1163 (O_1163,N_19387,N_19299);
or UO_1164 (O_1164,N_19295,N_19821);
or UO_1165 (O_1165,N_19971,N_19941);
nor UO_1166 (O_1166,N_19916,N_19398);
xnor UO_1167 (O_1167,N_19954,N_19516);
nor UO_1168 (O_1168,N_19426,N_19574);
xnor UO_1169 (O_1169,N_19923,N_19528);
xnor UO_1170 (O_1170,N_19620,N_19427);
nor UO_1171 (O_1171,N_19335,N_19555);
nand UO_1172 (O_1172,N_19970,N_19784);
xnor UO_1173 (O_1173,N_19589,N_19401);
or UO_1174 (O_1174,N_19589,N_19249);
nand UO_1175 (O_1175,N_19417,N_19318);
nand UO_1176 (O_1176,N_19594,N_19262);
xor UO_1177 (O_1177,N_19666,N_19596);
nor UO_1178 (O_1178,N_19553,N_19861);
xnor UO_1179 (O_1179,N_19834,N_19832);
or UO_1180 (O_1180,N_19266,N_19736);
nand UO_1181 (O_1181,N_19897,N_19778);
and UO_1182 (O_1182,N_19869,N_19732);
xor UO_1183 (O_1183,N_19235,N_19217);
nand UO_1184 (O_1184,N_19525,N_19490);
nor UO_1185 (O_1185,N_19544,N_19871);
nor UO_1186 (O_1186,N_19956,N_19513);
xor UO_1187 (O_1187,N_19573,N_19227);
nand UO_1188 (O_1188,N_19647,N_19209);
or UO_1189 (O_1189,N_19574,N_19349);
nor UO_1190 (O_1190,N_19529,N_19247);
nor UO_1191 (O_1191,N_19636,N_19290);
or UO_1192 (O_1192,N_19699,N_19203);
or UO_1193 (O_1193,N_19513,N_19270);
or UO_1194 (O_1194,N_19538,N_19484);
and UO_1195 (O_1195,N_19357,N_19702);
xnor UO_1196 (O_1196,N_19916,N_19859);
or UO_1197 (O_1197,N_19770,N_19490);
or UO_1198 (O_1198,N_19841,N_19843);
nand UO_1199 (O_1199,N_19696,N_19218);
or UO_1200 (O_1200,N_19703,N_19819);
xor UO_1201 (O_1201,N_19446,N_19541);
nor UO_1202 (O_1202,N_19976,N_19761);
or UO_1203 (O_1203,N_19613,N_19296);
nor UO_1204 (O_1204,N_19995,N_19450);
nand UO_1205 (O_1205,N_19556,N_19997);
and UO_1206 (O_1206,N_19648,N_19521);
or UO_1207 (O_1207,N_19245,N_19574);
nor UO_1208 (O_1208,N_19935,N_19425);
xor UO_1209 (O_1209,N_19688,N_19696);
nor UO_1210 (O_1210,N_19393,N_19754);
and UO_1211 (O_1211,N_19853,N_19480);
nor UO_1212 (O_1212,N_19328,N_19589);
xor UO_1213 (O_1213,N_19252,N_19598);
xor UO_1214 (O_1214,N_19361,N_19205);
nor UO_1215 (O_1215,N_19596,N_19434);
xor UO_1216 (O_1216,N_19858,N_19623);
or UO_1217 (O_1217,N_19208,N_19624);
and UO_1218 (O_1218,N_19656,N_19455);
and UO_1219 (O_1219,N_19227,N_19796);
or UO_1220 (O_1220,N_19590,N_19450);
or UO_1221 (O_1221,N_19287,N_19457);
or UO_1222 (O_1222,N_19607,N_19713);
and UO_1223 (O_1223,N_19824,N_19549);
and UO_1224 (O_1224,N_19711,N_19370);
or UO_1225 (O_1225,N_19626,N_19621);
and UO_1226 (O_1226,N_19799,N_19867);
or UO_1227 (O_1227,N_19325,N_19468);
nor UO_1228 (O_1228,N_19428,N_19859);
or UO_1229 (O_1229,N_19473,N_19839);
xnor UO_1230 (O_1230,N_19980,N_19868);
nand UO_1231 (O_1231,N_19783,N_19571);
and UO_1232 (O_1232,N_19857,N_19203);
xnor UO_1233 (O_1233,N_19596,N_19653);
nand UO_1234 (O_1234,N_19530,N_19423);
nand UO_1235 (O_1235,N_19971,N_19377);
nand UO_1236 (O_1236,N_19826,N_19583);
or UO_1237 (O_1237,N_19857,N_19745);
or UO_1238 (O_1238,N_19628,N_19426);
xor UO_1239 (O_1239,N_19984,N_19323);
or UO_1240 (O_1240,N_19927,N_19409);
xor UO_1241 (O_1241,N_19263,N_19930);
or UO_1242 (O_1242,N_19500,N_19261);
nor UO_1243 (O_1243,N_19638,N_19470);
nor UO_1244 (O_1244,N_19251,N_19252);
or UO_1245 (O_1245,N_19912,N_19662);
nor UO_1246 (O_1246,N_19557,N_19690);
nor UO_1247 (O_1247,N_19773,N_19367);
or UO_1248 (O_1248,N_19959,N_19327);
or UO_1249 (O_1249,N_19409,N_19298);
xor UO_1250 (O_1250,N_19412,N_19669);
and UO_1251 (O_1251,N_19815,N_19867);
nor UO_1252 (O_1252,N_19550,N_19495);
nor UO_1253 (O_1253,N_19688,N_19605);
nand UO_1254 (O_1254,N_19457,N_19953);
or UO_1255 (O_1255,N_19622,N_19772);
nand UO_1256 (O_1256,N_19973,N_19405);
xor UO_1257 (O_1257,N_19674,N_19720);
xnor UO_1258 (O_1258,N_19529,N_19492);
nor UO_1259 (O_1259,N_19546,N_19504);
and UO_1260 (O_1260,N_19939,N_19981);
nor UO_1261 (O_1261,N_19346,N_19751);
nor UO_1262 (O_1262,N_19599,N_19717);
and UO_1263 (O_1263,N_19355,N_19739);
nand UO_1264 (O_1264,N_19860,N_19894);
nor UO_1265 (O_1265,N_19929,N_19674);
xnor UO_1266 (O_1266,N_19643,N_19566);
or UO_1267 (O_1267,N_19497,N_19984);
and UO_1268 (O_1268,N_19400,N_19873);
xnor UO_1269 (O_1269,N_19634,N_19948);
nand UO_1270 (O_1270,N_19891,N_19378);
xnor UO_1271 (O_1271,N_19337,N_19459);
or UO_1272 (O_1272,N_19672,N_19832);
nand UO_1273 (O_1273,N_19426,N_19537);
nor UO_1274 (O_1274,N_19226,N_19275);
or UO_1275 (O_1275,N_19574,N_19510);
and UO_1276 (O_1276,N_19690,N_19473);
or UO_1277 (O_1277,N_19671,N_19602);
nor UO_1278 (O_1278,N_19209,N_19896);
nand UO_1279 (O_1279,N_19515,N_19289);
and UO_1280 (O_1280,N_19872,N_19787);
xnor UO_1281 (O_1281,N_19739,N_19285);
or UO_1282 (O_1282,N_19965,N_19262);
nor UO_1283 (O_1283,N_19923,N_19515);
xor UO_1284 (O_1284,N_19980,N_19296);
xnor UO_1285 (O_1285,N_19530,N_19998);
nand UO_1286 (O_1286,N_19689,N_19817);
xnor UO_1287 (O_1287,N_19870,N_19802);
and UO_1288 (O_1288,N_19628,N_19674);
nor UO_1289 (O_1289,N_19410,N_19230);
and UO_1290 (O_1290,N_19644,N_19219);
and UO_1291 (O_1291,N_19931,N_19841);
nand UO_1292 (O_1292,N_19359,N_19255);
nand UO_1293 (O_1293,N_19663,N_19973);
or UO_1294 (O_1294,N_19470,N_19646);
or UO_1295 (O_1295,N_19240,N_19314);
nor UO_1296 (O_1296,N_19648,N_19321);
or UO_1297 (O_1297,N_19717,N_19872);
xor UO_1298 (O_1298,N_19486,N_19558);
xor UO_1299 (O_1299,N_19370,N_19892);
and UO_1300 (O_1300,N_19947,N_19857);
nor UO_1301 (O_1301,N_19376,N_19843);
or UO_1302 (O_1302,N_19401,N_19694);
and UO_1303 (O_1303,N_19654,N_19602);
nand UO_1304 (O_1304,N_19606,N_19350);
nand UO_1305 (O_1305,N_19385,N_19794);
xnor UO_1306 (O_1306,N_19904,N_19626);
xnor UO_1307 (O_1307,N_19965,N_19976);
nand UO_1308 (O_1308,N_19821,N_19591);
xor UO_1309 (O_1309,N_19450,N_19882);
or UO_1310 (O_1310,N_19967,N_19911);
and UO_1311 (O_1311,N_19231,N_19254);
nor UO_1312 (O_1312,N_19865,N_19384);
xor UO_1313 (O_1313,N_19231,N_19269);
or UO_1314 (O_1314,N_19213,N_19650);
nor UO_1315 (O_1315,N_19749,N_19969);
nor UO_1316 (O_1316,N_19809,N_19700);
nand UO_1317 (O_1317,N_19555,N_19616);
nor UO_1318 (O_1318,N_19573,N_19684);
and UO_1319 (O_1319,N_19206,N_19904);
and UO_1320 (O_1320,N_19204,N_19375);
nand UO_1321 (O_1321,N_19639,N_19597);
or UO_1322 (O_1322,N_19295,N_19240);
and UO_1323 (O_1323,N_19869,N_19683);
nor UO_1324 (O_1324,N_19846,N_19811);
or UO_1325 (O_1325,N_19815,N_19646);
or UO_1326 (O_1326,N_19408,N_19238);
nor UO_1327 (O_1327,N_19332,N_19509);
and UO_1328 (O_1328,N_19454,N_19370);
and UO_1329 (O_1329,N_19685,N_19834);
xnor UO_1330 (O_1330,N_19531,N_19255);
nor UO_1331 (O_1331,N_19386,N_19643);
nor UO_1332 (O_1332,N_19305,N_19289);
or UO_1333 (O_1333,N_19658,N_19539);
and UO_1334 (O_1334,N_19632,N_19730);
and UO_1335 (O_1335,N_19886,N_19455);
xor UO_1336 (O_1336,N_19643,N_19587);
and UO_1337 (O_1337,N_19846,N_19241);
nor UO_1338 (O_1338,N_19934,N_19881);
nand UO_1339 (O_1339,N_19846,N_19994);
and UO_1340 (O_1340,N_19761,N_19652);
or UO_1341 (O_1341,N_19295,N_19283);
nand UO_1342 (O_1342,N_19676,N_19908);
or UO_1343 (O_1343,N_19647,N_19210);
nor UO_1344 (O_1344,N_19758,N_19828);
nand UO_1345 (O_1345,N_19884,N_19776);
xnor UO_1346 (O_1346,N_19325,N_19901);
xor UO_1347 (O_1347,N_19577,N_19254);
nand UO_1348 (O_1348,N_19430,N_19940);
nand UO_1349 (O_1349,N_19880,N_19395);
and UO_1350 (O_1350,N_19563,N_19294);
xor UO_1351 (O_1351,N_19722,N_19411);
xor UO_1352 (O_1352,N_19966,N_19251);
or UO_1353 (O_1353,N_19645,N_19696);
nor UO_1354 (O_1354,N_19971,N_19702);
or UO_1355 (O_1355,N_19539,N_19428);
or UO_1356 (O_1356,N_19612,N_19744);
or UO_1357 (O_1357,N_19813,N_19322);
xor UO_1358 (O_1358,N_19619,N_19725);
nand UO_1359 (O_1359,N_19482,N_19291);
nand UO_1360 (O_1360,N_19877,N_19795);
nand UO_1361 (O_1361,N_19955,N_19247);
nand UO_1362 (O_1362,N_19965,N_19947);
and UO_1363 (O_1363,N_19800,N_19388);
nor UO_1364 (O_1364,N_19497,N_19418);
nand UO_1365 (O_1365,N_19945,N_19643);
or UO_1366 (O_1366,N_19636,N_19273);
or UO_1367 (O_1367,N_19645,N_19534);
or UO_1368 (O_1368,N_19691,N_19608);
nor UO_1369 (O_1369,N_19394,N_19479);
nor UO_1370 (O_1370,N_19327,N_19371);
or UO_1371 (O_1371,N_19382,N_19716);
or UO_1372 (O_1372,N_19473,N_19367);
or UO_1373 (O_1373,N_19447,N_19363);
or UO_1374 (O_1374,N_19866,N_19776);
and UO_1375 (O_1375,N_19652,N_19345);
nand UO_1376 (O_1376,N_19697,N_19253);
nor UO_1377 (O_1377,N_19370,N_19562);
nor UO_1378 (O_1378,N_19854,N_19351);
and UO_1379 (O_1379,N_19233,N_19336);
xnor UO_1380 (O_1380,N_19500,N_19737);
xnor UO_1381 (O_1381,N_19299,N_19201);
nand UO_1382 (O_1382,N_19526,N_19632);
nor UO_1383 (O_1383,N_19727,N_19623);
or UO_1384 (O_1384,N_19861,N_19877);
xnor UO_1385 (O_1385,N_19219,N_19698);
nor UO_1386 (O_1386,N_19833,N_19555);
or UO_1387 (O_1387,N_19819,N_19893);
or UO_1388 (O_1388,N_19599,N_19913);
nor UO_1389 (O_1389,N_19423,N_19501);
or UO_1390 (O_1390,N_19274,N_19255);
xnor UO_1391 (O_1391,N_19846,N_19843);
and UO_1392 (O_1392,N_19340,N_19557);
or UO_1393 (O_1393,N_19362,N_19381);
and UO_1394 (O_1394,N_19459,N_19877);
xnor UO_1395 (O_1395,N_19701,N_19691);
or UO_1396 (O_1396,N_19770,N_19667);
nor UO_1397 (O_1397,N_19813,N_19299);
or UO_1398 (O_1398,N_19928,N_19346);
nor UO_1399 (O_1399,N_19425,N_19516);
xor UO_1400 (O_1400,N_19945,N_19852);
and UO_1401 (O_1401,N_19821,N_19745);
or UO_1402 (O_1402,N_19648,N_19434);
xnor UO_1403 (O_1403,N_19972,N_19271);
and UO_1404 (O_1404,N_19746,N_19480);
nor UO_1405 (O_1405,N_19407,N_19938);
or UO_1406 (O_1406,N_19687,N_19534);
nand UO_1407 (O_1407,N_19207,N_19461);
xor UO_1408 (O_1408,N_19709,N_19504);
xor UO_1409 (O_1409,N_19746,N_19490);
and UO_1410 (O_1410,N_19875,N_19878);
xor UO_1411 (O_1411,N_19735,N_19657);
and UO_1412 (O_1412,N_19280,N_19994);
nand UO_1413 (O_1413,N_19273,N_19493);
and UO_1414 (O_1414,N_19873,N_19877);
or UO_1415 (O_1415,N_19548,N_19639);
xor UO_1416 (O_1416,N_19700,N_19288);
xor UO_1417 (O_1417,N_19857,N_19966);
xor UO_1418 (O_1418,N_19647,N_19215);
xnor UO_1419 (O_1419,N_19898,N_19754);
and UO_1420 (O_1420,N_19414,N_19520);
or UO_1421 (O_1421,N_19527,N_19631);
nor UO_1422 (O_1422,N_19282,N_19816);
nor UO_1423 (O_1423,N_19240,N_19695);
nand UO_1424 (O_1424,N_19772,N_19604);
nand UO_1425 (O_1425,N_19686,N_19606);
or UO_1426 (O_1426,N_19383,N_19413);
nor UO_1427 (O_1427,N_19878,N_19342);
and UO_1428 (O_1428,N_19305,N_19469);
nor UO_1429 (O_1429,N_19508,N_19784);
nor UO_1430 (O_1430,N_19788,N_19908);
and UO_1431 (O_1431,N_19510,N_19643);
nor UO_1432 (O_1432,N_19885,N_19702);
xor UO_1433 (O_1433,N_19417,N_19293);
nand UO_1434 (O_1434,N_19389,N_19594);
and UO_1435 (O_1435,N_19381,N_19543);
nand UO_1436 (O_1436,N_19303,N_19715);
xor UO_1437 (O_1437,N_19977,N_19882);
nor UO_1438 (O_1438,N_19763,N_19502);
xor UO_1439 (O_1439,N_19831,N_19839);
nor UO_1440 (O_1440,N_19757,N_19408);
and UO_1441 (O_1441,N_19784,N_19507);
or UO_1442 (O_1442,N_19231,N_19741);
nor UO_1443 (O_1443,N_19281,N_19830);
xnor UO_1444 (O_1444,N_19276,N_19893);
nor UO_1445 (O_1445,N_19226,N_19273);
and UO_1446 (O_1446,N_19746,N_19947);
xnor UO_1447 (O_1447,N_19716,N_19521);
xor UO_1448 (O_1448,N_19633,N_19726);
xnor UO_1449 (O_1449,N_19489,N_19815);
xor UO_1450 (O_1450,N_19455,N_19397);
nand UO_1451 (O_1451,N_19904,N_19637);
nand UO_1452 (O_1452,N_19910,N_19522);
nor UO_1453 (O_1453,N_19620,N_19676);
xor UO_1454 (O_1454,N_19980,N_19813);
nor UO_1455 (O_1455,N_19514,N_19484);
nor UO_1456 (O_1456,N_19628,N_19662);
nor UO_1457 (O_1457,N_19768,N_19558);
nor UO_1458 (O_1458,N_19999,N_19976);
nor UO_1459 (O_1459,N_19824,N_19512);
xor UO_1460 (O_1460,N_19440,N_19739);
nand UO_1461 (O_1461,N_19547,N_19660);
or UO_1462 (O_1462,N_19831,N_19819);
and UO_1463 (O_1463,N_19296,N_19904);
or UO_1464 (O_1464,N_19942,N_19641);
and UO_1465 (O_1465,N_19270,N_19292);
nor UO_1466 (O_1466,N_19737,N_19726);
xor UO_1467 (O_1467,N_19534,N_19465);
nand UO_1468 (O_1468,N_19492,N_19527);
and UO_1469 (O_1469,N_19500,N_19857);
nand UO_1470 (O_1470,N_19590,N_19899);
nor UO_1471 (O_1471,N_19601,N_19893);
or UO_1472 (O_1472,N_19610,N_19473);
xnor UO_1473 (O_1473,N_19971,N_19853);
nor UO_1474 (O_1474,N_19782,N_19464);
nor UO_1475 (O_1475,N_19586,N_19524);
and UO_1476 (O_1476,N_19280,N_19325);
nand UO_1477 (O_1477,N_19360,N_19471);
or UO_1478 (O_1478,N_19688,N_19757);
nor UO_1479 (O_1479,N_19924,N_19577);
nor UO_1480 (O_1480,N_19370,N_19366);
or UO_1481 (O_1481,N_19865,N_19696);
or UO_1482 (O_1482,N_19219,N_19882);
or UO_1483 (O_1483,N_19318,N_19971);
xnor UO_1484 (O_1484,N_19721,N_19607);
xor UO_1485 (O_1485,N_19297,N_19777);
and UO_1486 (O_1486,N_19711,N_19937);
and UO_1487 (O_1487,N_19564,N_19832);
or UO_1488 (O_1488,N_19536,N_19656);
nand UO_1489 (O_1489,N_19301,N_19609);
nand UO_1490 (O_1490,N_19527,N_19880);
or UO_1491 (O_1491,N_19868,N_19410);
nand UO_1492 (O_1492,N_19281,N_19908);
or UO_1493 (O_1493,N_19777,N_19999);
xor UO_1494 (O_1494,N_19417,N_19715);
xor UO_1495 (O_1495,N_19516,N_19395);
and UO_1496 (O_1496,N_19728,N_19326);
nor UO_1497 (O_1497,N_19657,N_19433);
or UO_1498 (O_1498,N_19570,N_19932);
nor UO_1499 (O_1499,N_19462,N_19554);
or UO_1500 (O_1500,N_19653,N_19739);
and UO_1501 (O_1501,N_19701,N_19339);
or UO_1502 (O_1502,N_19936,N_19431);
nand UO_1503 (O_1503,N_19995,N_19539);
nor UO_1504 (O_1504,N_19356,N_19266);
and UO_1505 (O_1505,N_19876,N_19358);
and UO_1506 (O_1506,N_19557,N_19815);
or UO_1507 (O_1507,N_19405,N_19669);
nand UO_1508 (O_1508,N_19604,N_19839);
or UO_1509 (O_1509,N_19989,N_19831);
or UO_1510 (O_1510,N_19428,N_19230);
xor UO_1511 (O_1511,N_19634,N_19671);
nand UO_1512 (O_1512,N_19607,N_19247);
and UO_1513 (O_1513,N_19996,N_19615);
nor UO_1514 (O_1514,N_19779,N_19449);
and UO_1515 (O_1515,N_19338,N_19742);
nor UO_1516 (O_1516,N_19248,N_19739);
or UO_1517 (O_1517,N_19574,N_19835);
xnor UO_1518 (O_1518,N_19331,N_19310);
nand UO_1519 (O_1519,N_19300,N_19690);
xor UO_1520 (O_1520,N_19684,N_19405);
or UO_1521 (O_1521,N_19702,N_19576);
xnor UO_1522 (O_1522,N_19780,N_19652);
xnor UO_1523 (O_1523,N_19608,N_19248);
and UO_1524 (O_1524,N_19972,N_19772);
xor UO_1525 (O_1525,N_19947,N_19534);
nor UO_1526 (O_1526,N_19464,N_19716);
or UO_1527 (O_1527,N_19367,N_19665);
nor UO_1528 (O_1528,N_19841,N_19747);
nor UO_1529 (O_1529,N_19475,N_19486);
or UO_1530 (O_1530,N_19489,N_19640);
or UO_1531 (O_1531,N_19479,N_19571);
xor UO_1532 (O_1532,N_19612,N_19644);
xor UO_1533 (O_1533,N_19351,N_19864);
or UO_1534 (O_1534,N_19619,N_19804);
nand UO_1535 (O_1535,N_19484,N_19563);
nor UO_1536 (O_1536,N_19622,N_19354);
nand UO_1537 (O_1537,N_19786,N_19594);
and UO_1538 (O_1538,N_19771,N_19875);
nor UO_1539 (O_1539,N_19895,N_19234);
and UO_1540 (O_1540,N_19987,N_19581);
and UO_1541 (O_1541,N_19853,N_19615);
nor UO_1542 (O_1542,N_19643,N_19951);
or UO_1543 (O_1543,N_19379,N_19647);
xnor UO_1544 (O_1544,N_19628,N_19958);
xor UO_1545 (O_1545,N_19332,N_19596);
or UO_1546 (O_1546,N_19578,N_19919);
nand UO_1547 (O_1547,N_19392,N_19315);
nor UO_1548 (O_1548,N_19878,N_19529);
or UO_1549 (O_1549,N_19920,N_19794);
or UO_1550 (O_1550,N_19527,N_19845);
and UO_1551 (O_1551,N_19578,N_19577);
xor UO_1552 (O_1552,N_19229,N_19916);
xor UO_1553 (O_1553,N_19370,N_19540);
nor UO_1554 (O_1554,N_19219,N_19399);
nand UO_1555 (O_1555,N_19616,N_19312);
or UO_1556 (O_1556,N_19516,N_19396);
and UO_1557 (O_1557,N_19896,N_19827);
xor UO_1558 (O_1558,N_19283,N_19998);
and UO_1559 (O_1559,N_19335,N_19633);
or UO_1560 (O_1560,N_19243,N_19977);
nand UO_1561 (O_1561,N_19213,N_19510);
xnor UO_1562 (O_1562,N_19590,N_19393);
or UO_1563 (O_1563,N_19958,N_19668);
and UO_1564 (O_1564,N_19450,N_19321);
xor UO_1565 (O_1565,N_19951,N_19222);
or UO_1566 (O_1566,N_19873,N_19337);
and UO_1567 (O_1567,N_19440,N_19677);
or UO_1568 (O_1568,N_19656,N_19593);
nor UO_1569 (O_1569,N_19515,N_19919);
nor UO_1570 (O_1570,N_19706,N_19283);
and UO_1571 (O_1571,N_19806,N_19298);
nor UO_1572 (O_1572,N_19586,N_19900);
xor UO_1573 (O_1573,N_19475,N_19501);
nor UO_1574 (O_1574,N_19954,N_19882);
nor UO_1575 (O_1575,N_19770,N_19707);
xor UO_1576 (O_1576,N_19736,N_19535);
or UO_1577 (O_1577,N_19619,N_19930);
nor UO_1578 (O_1578,N_19810,N_19980);
and UO_1579 (O_1579,N_19343,N_19914);
or UO_1580 (O_1580,N_19938,N_19798);
nand UO_1581 (O_1581,N_19728,N_19505);
nor UO_1582 (O_1582,N_19790,N_19563);
nor UO_1583 (O_1583,N_19509,N_19987);
nor UO_1584 (O_1584,N_19358,N_19593);
and UO_1585 (O_1585,N_19664,N_19896);
and UO_1586 (O_1586,N_19683,N_19347);
nor UO_1587 (O_1587,N_19398,N_19711);
nor UO_1588 (O_1588,N_19680,N_19314);
xor UO_1589 (O_1589,N_19310,N_19810);
xor UO_1590 (O_1590,N_19905,N_19544);
and UO_1591 (O_1591,N_19581,N_19783);
nor UO_1592 (O_1592,N_19511,N_19265);
nand UO_1593 (O_1593,N_19467,N_19652);
xnor UO_1594 (O_1594,N_19252,N_19828);
nand UO_1595 (O_1595,N_19396,N_19529);
or UO_1596 (O_1596,N_19960,N_19859);
xnor UO_1597 (O_1597,N_19286,N_19480);
nand UO_1598 (O_1598,N_19891,N_19383);
xor UO_1599 (O_1599,N_19843,N_19309);
or UO_1600 (O_1600,N_19242,N_19944);
xnor UO_1601 (O_1601,N_19251,N_19499);
and UO_1602 (O_1602,N_19554,N_19522);
nor UO_1603 (O_1603,N_19857,N_19461);
or UO_1604 (O_1604,N_19466,N_19242);
nor UO_1605 (O_1605,N_19739,N_19216);
nor UO_1606 (O_1606,N_19243,N_19374);
or UO_1607 (O_1607,N_19659,N_19356);
nand UO_1608 (O_1608,N_19975,N_19688);
xor UO_1609 (O_1609,N_19528,N_19426);
or UO_1610 (O_1610,N_19735,N_19393);
and UO_1611 (O_1611,N_19532,N_19328);
and UO_1612 (O_1612,N_19586,N_19324);
nor UO_1613 (O_1613,N_19950,N_19648);
and UO_1614 (O_1614,N_19825,N_19267);
xor UO_1615 (O_1615,N_19918,N_19896);
nand UO_1616 (O_1616,N_19385,N_19498);
nand UO_1617 (O_1617,N_19331,N_19874);
nand UO_1618 (O_1618,N_19679,N_19894);
nand UO_1619 (O_1619,N_19362,N_19314);
and UO_1620 (O_1620,N_19839,N_19714);
nand UO_1621 (O_1621,N_19343,N_19794);
nor UO_1622 (O_1622,N_19932,N_19689);
nand UO_1623 (O_1623,N_19963,N_19443);
or UO_1624 (O_1624,N_19656,N_19977);
nand UO_1625 (O_1625,N_19931,N_19897);
xnor UO_1626 (O_1626,N_19799,N_19607);
nand UO_1627 (O_1627,N_19901,N_19692);
nor UO_1628 (O_1628,N_19716,N_19467);
and UO_1629 (O_1629,N_19357,N_19430);
or UO_1630 (O_1630,N_19304,N_19260);
and UO_1631 (O_1631,N_19510,N_19505);
nand UO_1632 (O_1632,N_19741,N_19559);
nand UO_1633 (O_1633,N_19888,N_19754);
and UO_1634 (O_1634,N_19789,N_19370);
nor UO_1635 (O_1635,N_19827,N_19925);
and UO_1636 (O_1636,N_19547,N_19549);
and UO_1637 (O_1637,N_19946,N_19668);
xnor UO_1638 (O_1638,N_19454,N_19346);
xnor UO_1639 (O_1639,N_19253,N_19629);
and UO_1640 (O_1640,N_19784,N_19347);
nand UO_1641 (O_1641,N_19439,N_19593);
nor UO_1642 (O_1642,N_19299,N_19220);
or UO_1643 (O_1643,N_19388,N_19453);
and UO_1644 (O_1644,N_19440,N_19599);
xor UO_1645 (O_1645,N_19619,N_19845);
nor UO_1646 (O_1646,N_19406,N_19269);
or UO_1647 (O_1647,N_19211,N_19621);
xnor UO_1648 (O_1648,N_19721,N_19858);
nand UO_1649 (O_1649,N_19559,N_19301);
and UO_1650 (O_1650,N_19468,N_19834);
nand UO_1651 (O_1651,N_19955,N_19649);
nand UO_1652 (O_1652,N_19708,N_19519);
nor UO_1653 (O_1653,N_19958,N_19687);
and UO_1654 (O_1654,N_19468,N_19738);
nor UO_1655 (O_1655,N_19574,N_19457);
and UO_1656 (O_1656,N_19782,N_19330);
nor UO_1657 (O_1657,N_19614,N_19769);
nand UO_1658 (O_1658,N_19251,N_19898);
nand UO_1659 (O_1659,N_19919,N_19202);
and UO_1660 (O_1660,N_19428,N_19596);
and UO_1661 (O_1661,N_19602,N_19897);
and UO_1662 (O_1662,N_19273,N_19556);
nor UO_1663 (O_1663,N_19981,N_19205);
and UO_1664 (O_1664,N_19382,N_19570);
xor UO_1665 (O_1665,N_19223,N_19663);
xor UO_1666 (O_1666,N_19462,N_19513);
or UO_1667 (O_1667,N_19350,N_19250);
and UO_1668 (O_1668,N_19376,N_19512);
or UO_1669 (O_1669,N_19633,N_19500);
or UO_1670 (O_1670,N_19970,N_19519);
nor UO_1671 (O_1671,N_19725,N_19617);
or UO_1672 (O_1672,N_19536,N_19422);
or UO_1673 (O_1673,N_19360,N_19903);
nand UO_1674 (O_1674,N_19495,N_19303);
nor UO_1675 (O_1675,N_19357,N_19557);
and UO_1676 (O_1676,N_19996,N_19329);
nor UO_1677 (O_1677,N_19378,N_19824);
or UO_1678 (O_1678,N_19608,N_19388);
or UO_1679 (O_1679,N_19723,N_19674);
nand UO_1680 (O_1680,N_19491,N_19725);
nor UO_1681 (O_1681,N_19760,N_19284);
nor UO_1682 (O_1682,N_19981,N_19298);
xnor UO_1683 (O_1683,N_19718,N_19669);
and UO_1684 (O_1684,N_19817,N_19801);
or UO_1685 (O_1685,N_19657,N_19434);
and UO_1686 (O_1686,N_19894,N_19346);
and UO_1687 (O_1687,N_19932,N_19794);
and UO_1688 (O_1688,N_19825,N_19699);
xor UO_1689 (O_1689,N_19813,N_19525);
or UO_1690 (O_1690,N_19451,N_19449);
nor UO_1691 (O_1691,N_19618,N_19829);
and UO_1692 (O_1692,N_19272,N_19367);
xnor UO_1693 (O_1693,N_19293,N_19576);
nand UO_1694 (O_1694,N_19349,N_19597);
or UO_1695 (O_1695,N_19617,N_19272);
xnor UO_1696 (O_1696,N_19817,N_19657);
xor UO_1697 (O_1697,N_19375,N_19398);
and UO_1698 (O_1698,N_19640,N_19221);
or UO_1699 (O_1699,N_19239,N_19379);
xor UO_1700 (O_1700,N_19422,N_19534);
xor UO_1701 (O_1701,N_19282,N_19601);
nor UO_1702 (O_1702,N_19843,N_19935);
xnor UO_1703 (O_1703,N_19967,N_19274);
or UO_1704 (O_1704,N_19441,N_19625);
and UO_1705 (O_1705,N_19468,N_19402);
nand UO_1706 (O_1706,N_19698,N_19858);
xor UO_1707 (O_1707,N_19724,N_19276);
xor UO_1708 (O_1708,N_19933,N_19415);
or UO_1709 (O_1709,N_19287,N_19267);
nand UO_1710 (O_1710,N_19214,N_19860);
xnor UO_1711 (O_1711,N_19707,N_19871);
nor UO_1712 (O_1712,N_19207,N_19427);
xor UO_1713 (O_1713,N_19330,N_19589);
or UO_1714 (O_1714,N_19475,N_19920);
xor UO_1715 (O_1715,N_19741,N_19461);
and UO_1716 (O_1716,N_19501,N_19276);
or UO_1717 (O_1717,N_19281,N_19907);
nand UO_1718 (O_1718,N_19420,N_19643);
or UO_1719 (O_1719,N_19937,N_19386);
nor UO_1720 (O_1720,N_19466,N_19393);
nor UO_1721 (O_1721,N_19387,N_19377);
nand UO_1722 (O_1722,N_19336,N_19894);
and UO_1723 (O_1723,N_19766,N_19579);
or UO_1724 (O_1724,N_19386,N_19426);
or UO_1725 (O_1725,N_19980,N_19827);
xnor UO_1726 (O_1726,N_19214,N_19623);
nor UO_1727 (O_1727,N_19506,N_19912);
nand UO_1728 (O_1728,N_19432,N_19956);
nand UO_1729 (O_1729,N_19611,N_19769);
nor UO_1730 (O_1730,N_19936,N_19596);
and UO_1731 (O_1731,N_19215,N_19517);
nand UO_1732 (O_1732,N_19447,N_19863);
or UO_1733 (O_1733,N_19705,N_19258);
nand UO_1734 (O_1734,N_19341,N_19988);
and UO_1735 (O_1735,N_19973,N_19587);
and UO_1736 (O_1736,N_19624,N_19487);
xnor UO_1737 (O_1737,N_19495,N_19789);
nor UO_1738 (O_1738,N_19252,N_19808);
xor UO_1739 (O_1739,N_19944,N_19370);
and UO_1740 (O_1740,N_19483,N_19329);
or UO_1741 (O_1741,N_19710,N_19746);
or UO_1742 (O_1742,N_19777,N_19419);
nand UO_1743 (O_1743,N_19620,N_19854);
xnor UO_1744 (O_1744,N_19531,N_19772);
nor UO_1745 (O_1745,N_19442,N_19835);
or UO_1746 (O_1746,N_19731,N_19583);
nand UO_1747 (O_1747,N_19289,N_19511);
nor UO_1748 (O_1748,N_19909,N_19337);
nor UO_1749 (O_1749,N_19607,N_19326);
nor UO_1750 (O_1750,N_19429,N_19685);
or UO_1751 (O_1751,N_19988,N_19274);
nand UO_1752 (O_1752,N_19986,N_19795);
or UO_1753 (O_1753,N_19799,N_19828);
nor UO_1754 (O_1754,N_19686,N_19451);
nand UO_1755 (O_1755,N_19251,N_19301);
or UO_1756 (O_1756,N_19224,N_19741);
nor UO_1757 (O_1757,N_19819,N_19704);
and UO_1758 (O_1758,N_19452,N_19449);
nor UO_1759 (O_1759,N_19413,N_19745);
and UO_1760 (O_1760,N_19566,N_19695);
nor UO_1761 (O_1761,N_19762,N_19866);
and UO_1762 (O_1762,N_19403,N_19705);
or UO_1763 (O_1763,N_19611,N_19760);
and UO_1764 (O_1764,N_19492,N_19389);
and UO_1765 (O_1765,N_19812,N_19269);
xnor UO_1766 (O_1766,N_19947,N_19926);
and UO_1767 (O_1767,N_19972,N_19982);
and UO_1768 (O_1768,N_19951,N_19915);
or UO_1769 (O_1769,N_19547,N_19706);
nor UO_1770 (O_1770,N_19628,N_19417);
nor UO_1771 (O_1771,N_19219,N_19314);
and UO_1772 (O_1772,N_19516,N_19882);
or UO_1773 (O_1773,N_19809,N_19869);
or UO_1774 (O_1774,N_19958,N_19257);
xor UO_1775 (O_1775,N_19678,N_19504);
nand UO_1776 (O_1776,N_19439,N_19644);
xor UO_1777 (O_1777,N_19347,N_19656);
and UO_1778 (O_1778,N_19689,N_19406);
xor UO_1779 (O_1779,N_19746,N_19628);
nor UO_1780 (O_1780,N_19633,N_19971);
and UO_1781 (O_1781,N_19311,N_19650);
xor UO_1782 (O_1782,N_19737,N_19530);
nand UO_1783 (O_1783,N_19427,N_19407);
nor UO_1784 (O_1784,N_19672,N_19524);
nor UO_1785 (O_1785,N_19370,N_19756);
nor UO_1786 (O_1786,N_19608,N_19445);
and UO_1787 (O_1787,N_19815,N_19772);
nand UO_1788 (O_1788,N_19693,N_19729);
and UO_1789 (O_1789,N_19482,N_19243);
nand UO_1790 (O_1790,N_19490,N_19590);
nand UO_1791 (O_1791,N_19845,N_19822);
nand UO_1792 (O_1792,N_19248,N_19473);
nand UO_1793 (O_1793,N_19208,N_19771);
nand UO_1794 (O_1794,N_19329,N_19240);
or UO_1795 (O_1795,N_19517,N_19688);
nand UO_1796 (O_1796,N_19461,N_19421);
nand UO_1797 (O_1797,N_19769,N_19939);
and UO_1798 (O_1798,N_19467,N_19302);
nand UO_1799 (O_1799,N_19703,N_19709);
xnor UO_1800 (O_1800,N_19969,N_19554);
and UO_1801 (O_1801,N_19331,N_19619);
or UO_1802 (O_1802,N_19269,N_19259);
xor UO_1803 (O_1803,N_19853,N_19816);
xnor UO_1804 (O_1804,N_19845,N_19404);
or UO_1805 (O_1805,N_19856,N_19261);
or UO_1806 (O_1806,N_19278,N_19615);
and UO_1807 (O_1807,N_19337,N_19987);
xor UO_1808 (O_1808,N_19464,N_19578);
xnor UO_1809 (O_1809,N_19307,N_19328);
xnor UO_1810 (O_1810,N_19735,N_19717);
and UO_1811 (O_1811,N_19318,N_19700);
xnor UO_1812 (O_1812,N_19388,N_19508);
nor UO_1813 (O_1813,N_19332,N_19820);
nand UO_1814 (O_1814,N_19970,N_19915);
xor UO_1815 (O_1815,N_19430,N_19696);
nand UO_1816 (O_1816,N_19285,N_19745);
nand UO_1817 (O_1817,N_19844,N_19591);
xnor UO_1818 (O_1818,N_19412,N_19208);
and UO_1819 (O_1819,N_19980,N_19852);
nand UO_1820 (O_1820,N_19492,N_19746);
and UO_1821 (O_1821,N_19882,N_19622);
xnor UO_1822 (O_1822,N_19511,N_19728);
nand UO_1823 (O_1823,N_19992,N_19451);
nor UO_1824 (O_1824,N_19518,N_19646);
nand UO_1825 (O_1825,N_19683,N_19878);
and UO_1826 (O_1826,N_19247,N_19579);
nand UO_1827 (O_1827,N_19407,N_19786);
or UO_1828 (O_1828,N_19935,N_19431);
or UO_1829 (O_1829,N_19619,N_19329);
nand UO_1830 (O_1830,N_19301,N_19675);
nand UO_1831 (O_1831,N_19232,N_19661);
or UO_1832 (O_1832,N_19561,N_19597);
nor UO_1833 (O_1833,N_19718,N_19621);
or UO_1834 (O_1834,N_19883,N_19508);
xor UO_1835 (O_1835,N_19528,N_19496);
nand UO_1836 (O_1836,N_19334,N_19243);
nor UO_1837 (O_1837,N_19475,N_19363);
nand UO_1838 (O_1838,N_19434,N_19904);
nor UO_1839 (O_1839,N_19490,N_19964);
or UO_1840 (O_1840,N_19780,N_19977);
and UO_1841 (O_1841,N_19289,N_19842);
nor UO_1842 (O_1842,N_19782,N_19944);
and UO_1843 (O_1843,N_19522,N_19945);
nand UO_1844 (O_1844,N_19349,N_19456);
nor UO_1845 (O_1845,N_19457,N_19565);
nand UO_1846 (O_1846,N_19637,N_19852);
nor UO_1847 (O_1847,N_19874,N_19688);
xnor UO_1848 (O_1848,N_19257,N_19636);
nor UO_1849 (O_1849,N_19611,N_19320);
xor UO_1850 (O_1850,N_19948,N_19907);
nand UO_1851 (O_1851,N_19272,N_19686);
nor UO_1852 (O_1852,N_19881,N_19642);
or UO_1853 (O_1853,N_19813,N_19647);
nand UO_1854 (O_1854,N_19905,N_19423);
nand UO_1855 (O_1855,N_19890,N_19421);
xor UO_1856 (O_1856,N_19605,N_19917);
nor UO_1857 (O_1857,N_19587,N_19354);
nand UO_1858 (O_1858,N_19247,N_19936);
nor UO_1859 (O_1859,N_19692,N_19303);
nand UO_1860 (O_1860,N_19875,N_19600);
nor UO_1861 (O_1861,N_19385,N_19213);
xnor UO_1862 (O_1862,N_19556,N_19334);
xnor UO_1863 (O_1863,N_19651,N_19233);
or UO_1864 (O_1864,N_19526,N_19374);
or UO_1865 (O_1865,N_19394,N_19271);
or UO_1866 (O_1866,N_19556,N_19776);
nor UO_1867 (O_1867,N_19467,N_19503);
nand UO_1868 (O_1868,N_19677,N_19473);
or UO_1869 (O_1869,N_19966,N_19566);
nor UO_1870 (O_1870,N_19617,N_19662);
xor UO_1871 (O_1871,N_19402,N_19481);
xor UO_1872 (O_1872,N_19802,N_19670);
nor UO_1873 (O_1873,N_19222,N_19804);
xnor UO_1874 (O_1874,N_19826,N_19474);
xor UO_1875 (O_1875,N_19356,N_19608);
xor UO_1876 (O_1876,N_19917,N_19508);
nor UO_1877 (O_1877,N_19561,N_19575);
nand UO_1878 (O_1878,N_19905,N_19644);
nor UO_1879 (O_1879,N_19608,N_19906);
nand UO_1880 (O_1880,N_19489,N_19336);
and UO_1881 (O_1881,N_19509,N_19972);
nand UO_1882 (O_1882,N_19202,N_19236);
or UO_1883 (O_1883,N_19827,N_19848);
nand UO_1884 (O_1884,N_19372,N_19964);
and UO_1885 (O_1885,N_19737,N_19805);
or UO_1886 (O_1886,N_19528,N_19473);
nor UO_1887 (O_1887,N_19847,N_19711);
or UO_1888 (O_1888,N_19764,N_19640);
xnor UO_1889 (O_1889,N_19672,N_19455);
nand UO_1890 (O_1890,N_19559,N_19536);
nand UO_1891 (O_1891,N_19577,N_19597);
or UO_1892 (O_1892,N_19732,N_19529);
nor UO_1893 (O_1893,N_19292,N_19479);
nand UO_1894 (O_1894,N_19649,N_19368);
or UO_1895 (O_1895,N_19535,N_19585);
or UO_1896 (O_1896,N_19266,N_19485);
xor UO_1897 (O_1897,N_19640,N_19829);
and UO_1898 (O_1898,N_19540,N_19538);
nor UO_1899 (O_1899,N_19643,N_19283);
or UO_1900 (O_1900,N_19838,N_19826);
and UO_1901 (O_1901,N_19709,N_19997);
or UO_1902 (O_1902,N_19759,N_19254);
or UO_1903 (O_1903,N_19290,N_19279);
nand UO_1904 (O_1904,N_19314,N_19718);
xnor UO_1905 (O_1905,N_19725,N_19574);
and UO_1906 (O_1906,N_19685,N_19616);
or UO_1907 (O_1907,N_19542,N_19771);
or UO_1908 (O_1908,N_19548,N_19877);
nor UO_1909 (O_1909,N_19497,N_19544);
nor UO_1910 (O_1910,N_19793,N_19238);
nand UO_1911 (O_1911,N_19388,N_19981);
xor UO_1912 (O_1912,N_19434,N_19969);
or UO_1913 (O_1913,N_19725,N_19605);
nor UO_1914 (O_1914,N_19287,N_19782);
and UO_1915 (O_1915,N_19757,N_19921);
xor UO_1916 (O_1916,N_19575,N_19385);
xnor UO_1917 (O_1917,N_19826,N_19228);
nand UO_1918 (O_1918,N_19272,N_19793);
and UO_1919 (O_1919,N_19342,N_19821);
xor UO_1920 (O_1920,N_19304,N_19322);
nor UO_1921 (O_1921,N_19595,N_19714);
and UO_1922 (O_1922,N_19614,N_19396);
nand UO_1923 (O_1923,N_19222,N_19461);
nor UO_1924 (O_1924,N_19697,N_19260);
and UO_1925 (O_1925,N_19889,N_19989);
or UO_1926 (O_1926,N_19983,N_19836);
and UO_1927 (O_1927,N_19551,N_19398);
xnor UO_1928 (O_1928,N_19469,N_19787);
and UO_1929 (O_1929,N_19707,N_19815);
and UO_1930 (O_1930,N_19541,N_19690);
and UO_1931 (O_1931,N_19942,N_19204);
nor UO_1932 (O_1932,N_19892,N_19601);
nor UO_1933 (O_1933,N_19236,N_19239);
or UO_1934 (O_1934,N_19798,N_19635);
nand UO_1935 (O_1935,N_19655,N_19371);
or UO_1936 (O_1936,N_19792,N_19961);
xor UO_1937 (O_1937,N_19362,N_19338);
nand UO_1938 (O_1938,N_19335,N_19411);
nand UO_1939 (O_1939,N_19822,N_19794);
xnor UO_1940 (O_1940,N_19539,N_19315);
and UO_1941 (O_1941,N_19700,N_19476);
and UO_1942 (O_1942,N_19776,N_19459);
nor UO_1943 (O_1943,N_19810,N_19493);
xor UO_1944 (O_1944,N_19228,N_19750);
nor UO_1945 (O_1945,N_19774,N_19609);
xnor UO_1946 (O_1946,N_19894,N_19214);
xnor UO_1947 (O_1947,N_19505,N_19746);
nor UO_1948 (O_1948,N_19978,N_19602);
and UO_1949 (O_1949,N_19490,N_19859);
or UO_1950 (O_1950,N_19487,N_19414);
or UO_1951 (O_1951,N_19203,N_19516);
nor UO_1952 (O_1952,N_19830,N_19724);
xnor UO_1953 (O_1953,N_19633,N_19306);
and UO_1954 (O_1954,N_19253,N_19490);
xnor UO_1955 (O_1955,N_19822,N_19290);
nand UO_1956 (O_1956,N_19403,N_19318);
and UO_1957 (O_1957,N_19529,N_19840);
or UO_1958 (O_1958,N_19420,N_19264);
nor UO_1959 (O_1959,N_19737,N_19674);
nor UO_1960 (O_1960,N_19367,N_19881);
nand UO_1961 (O_1961,N_19857,N_19954);
nand UO_1962 (O_1962,N_19637,N_19939);
and UO_1963 (O_1963,N_19338,N_19469);
xor UO_1964 (O_1964,N_19942,N_19934);
nand UO_1965 (O_1965,N_19881,N_19611);
nand UO_1966 (O_1966,N_19427,N_19909);
nand UO_1967 (O_1967,N_19694,N_19250);
or UO_1968 (O_1968,N_19968,N_19781);
and UO_1969 (O_1969,N_19551,N_19545);
and UO_1970 (O_1970,N_19319,N_19625);
and UO_1971 (O_1971,N_19571,N_19850);
nor UO_1972 (O_1972,N_19260,N_19411);
and UO_1973 (O_1973,N_19619,N_19209);
nand UO_1974 (O_1974,N_19702,N_19209);
nand UO_1975 (O_1975,N_19587,N_19646);
nor UO_1976 (O_1976,N_19404,N_19611);
and UO_1977 (O_1977,N_19638,N_19880);
or UO_1978 (O_1978,N_19242,N_19642);
nand UO_1979 (O_1979,N_19807,N_19665);
and UO_1980 (O_1980,N_19845,N_19915);
nand UO_1981 (O_1981,N_19787,N_19421);
nor UO_1982 (O_1982,N_19379,N_19548);
xor UO_1983 (O_1983,N_19611,N_19274);
xnor UO_1984 (O_1984,N_19275,N_19602);
xnor UO_1985 (O_1985,N_19429,N_19727);
or UO_1986 (O_1986,N_19380,N_19851);
and UO_1987 (O_1987,N_19257,N_19810);
and UO_1988 (O_1988,N_19553,N_19988);
xnor UO_1989 (O_1989,N_19252,N_19702);
nor UO_1990 (O_1990,N_19699,N_19930);
nand UO_1991 (O_1991,N_19604,N_19543);
xor UO_1992 (O_1992,N_19454,N_19623);
or UO_1993 (O_1993,N_19740,N_19411);
nor UO_1994 (O_1994,N_19593,N_19999);
or UO_1995 (O_1995,N_19993,N_19378);
nand UO_1996 (O_1996,N_19474,N_19278);
xor UO_1997 (O_1997,N_19949,N_19622);
and UO_1998 (O_1998,N_19591,N_19697);
or UO_1999 (O_1999,N_19204,N_19625);
nand UO_2000 (O_2000,N_19219,N_19618);
nand UO_2001 (O_2001,N_19700,N_19304);
nand UO_2002 (O_2002,N_19695,N_19751);
nor UO_2003 (O_2003,N_19637,N_19310);
nor UO_2004 (O_2004,N_19882,N_19528);
or UO_2005 (O_2005,N_19382,N_19837);
and UO_2006 (O_2006,N_19853,N_19741);
nor UO_2007 (O_2007,N_19747,N_19280);
and UO_2008 (O_2008,N_19385,N_19557);
or UO_2009 (O_2009,N_19326,N_19517);
or UO_2010 (O_2010,N_19246,N_19339);
and UO_2011 (O_2011,N_19574,N_19603);
nand UO_2012 (O_2012,N_19231,N_19220);
or UO_2013 (O_2013,N_19974,N_19658);
nand UO_2014 (O_2014,N_19751,N_19332);
xnor UO_2015 (O_2015,N_19848,N_19262);
and UO_2016 (O_2016,N_19259,N_19297);
and UO_2017 (O_2017,N_19543,N_19672);
and UO_2018 (O_2018,N_19375,N_19593);
nor UO_2019 (O_2019,N_19936,N_19228);
xor UO_2020 (O_2020,N_19595,N_19593);
and UO_2021 (O_2021,N_19692,N_19738);
nor UO_2022 (O_2022,N_19311,N_19721);
and UO_2023 (O_2023,N_19889,N_19386);
and UO_2024 (O_2024,N_19938,N_19733);
and UO_2025 (O_2025,N_19460,N_19968);
nand UO_2026 (O_2026,N_19718,N_19220);
xnor UO_2027 (O_2027,N_19952,N_19968);
and UO_2028 (O_2028,N_19272,N_19518);
nand UO_2029 (O_2029,N_19387,N_19546);
xor UO_2030 (O_2030,N_19391,N_19999);
or UO_2031 (O_2031,N_19214,N_19974);
nand UO_2032 (O_2032,N_19810,N_19873);
nor UO_2033 (O_2033,N_19256,N_19933);
and UO_2034 (O_2034,N_19290,N_19344);
nand UO_2035 (O_2035,N_19884,N_19934);
or UO_2036 (O_2036,N_19943,N_19461);
xor UO_2037 (O_2037,N_19398,N_19311);
nand UO_2038 (O_2038,N_19833,N_19587);
and UO_2039 (O_2039,N_19579,N_19850);
or UO_2040 (O_2040,N_19368,N_19932);
xor UO_2041 (O_2041,N_19798,N_19631);
or UO_2042 (O_2042,N_19704,N_19734);
nor UO_2043 (O_2043,N_19852,N_19450);
nor UO_2044 (O_2044,N_19240,N_19428);
nand UO_2045 (O_2045,N_19426,N_19271);
xor UO_2046 (O_2046,N_19856,N_19664);
nand UO_2047 (O_2047,N_19276,N_19352);
nand UO_2048 (O_2048,N_19741,N_19770);
and UO_2049 (O_2049,N_19865,N_19285);
or UO_2050 (O_2050,N_19879,N_19480);
and UO_2051 (O_2051,N_19827,N_19748);
and UO_2052 (O_2052,N_19540,N_19606);
or UO_2053 (O_2053,N_19686,N_19450);
xnor UO_2054 (O_2054,N_19323,N_19214);
nand UO_2055 (O_2055,N_19875,N_19283);
or UO_2056 (O_2056,N_19742,N_19680);
xor UO_2057 (O_2057,N_19288,N_19688);
and UO_2058 (O_2058,N_19980,N_19564);
xnor UO_2059 (O_2059,N_19815,N_19507);
nor UO_2060 (O_2060,N_19284,N_19560);
or UO_2061 (O_2061,N_19739,N_19742);
or UO_2062 (O_2062,N_19997,N_19956);
xor UO_2063 (O_2063,N_19990,N_19649);
and UO_2064 (O_2064,N_19842,N_19807);
and UO_2065 (O_2065,N_19523,N_19712);
xor UO_2066 (O_2066,N_19473,N_19830);
nor UO_2067 (O_2067,N_19375,N_19340);
and UO_2068 (O_2068,N_19849,N_19528);
and UO_2069 (O_2069,N_19905,N_19692);
nand UO_2070 (O_2070,N_19480,N_19718);
xnor UO_2071 (O_2071,N_19333,N_19987);
xor UO_2072 (O_2072,N_19217,N_19470);
and UO_2073 (O_2073,N_19885,N_19529);
xnor UO_2074 (O_2074,N_19448,N_19320);
or UO_2075 (O_2075,N_19282,N_19233);
or UO_2076 (O_2076,N_19510,N_19751);
and UO_2077 (O_2077,N_19213,N_19430);
or UO_2078 (O_2078,N_19642,N_19432);
and UO_2079 (O_2079,N_19640,N_19306);
nand UO_2080 (O_2080,N_19488,N_19596);
or UO_2081 (O_2081,N_19874,N_19539);
nand UO_2082 (O_2082,N_19293,N_19447);
and UO_2083 (O_2083,N_19935,N_19930);
or UO_2084 (O_2084,N_19746,N_19281);
or UO_2085 (O_2085,N_19809,N_19989);
or UO_2086 (O_2086,N_19447,N_19789);
and UO_2087 (O_2087,N_19387,N_19993);
or UO_2088 (O_2088,N_19842,N_19878);
or UO_2089 (O_2089,N_19388,N_19847);
or UO_2090 (O_2090,N_19596,N_19894);
nor UO_2091 (O_2091,N_19583,N_19747);
nor UO_2092 (O_2092,N_19806,N_19715);
and UO_2093 (O_2093,N_19622,N_19587);
nand UO_2094 (O_2094,N_19636,N_19265);
nor UO_2095 (O_2095,N_19506,N_19952);
nand UO_2096 (O_2096,N_19498,N_19494);
nor UO_2097 (O_2097,N_19986,N_19757);
or UO_2098 (O_2098,N_19754,N_19616);
and UO_2099 (O_2099,N_19960,N_19546);
nor UO_2100 (O_2100,N_19442,N_19609);
or UO_2101 (O_2101,N_19733,N_19627);
or UO_2102 (O_2102,N_19791,N_19415);
or UO_2103 (O_2103,N_19595,N_19601);
nor UO_2104 (O_2104,N_19224,N_19465);
xnor UO_2105 (O_2105,N_19269,N_19889);
and UO_2106 (O_2106,N_19823,N_19706);
and UO_2107 (O_2107,N_19472,N_19497);
and UO_2108 (O_2108,N_19622,N_19808);
nor UO_2109 (O_2109,N_19213,N_19740);
and UO_2110 (O_2110,N_19867,N_19849);
nand UO_2111 (O_2111,N_19347,N_19732);
and UO_2112 (O_2112,N_19996,N_19986);
xor UO_2113 (O_2113,N_19821,N_19695);
nor UO_2114 (O_2114,N_19882,N_19649);
nor UO_2115 (O_2115,N_19846,N_19924);
or UO_2116 (O_2116,N_19530,N_19402);
nand UO_2117 (O_2117,N_19964,N_19460);
xor UO_2118 (O_2118,N_19472,N_19297);
xnor UO_2119 (O_2119,N_19763,N_19236);
nor UO_2120 (O_2120,N_19952,N_19801);
or UO_2121 (O_2121,N_19327,N_19367);
xnor UO_2122 (O_2122,N_19313,N_19422);
or UO_2123 (O_2123,N_19906,N_19712);
and UO_2124 (O_2124,N_19621,N_19644);
or UO_2125 (O_2125,N_19839,N_19403);
nand UO_2126 (O_2126,N_19739,N_19814);
or UO_2127 (O_2127,N_19396,N_19663);
or UO_2128 (O_2128,N_19261,N_19226);
and UO_2129 (O_2129,N_19662,N_19489);
xor UO_2130 (O_2130,N_19896,N_19317);
nor UO_2131 (O_2131,N_19231,N_19379);
or UO_2132 (O_2132,N_19324,N_19862);
nor UO_2133 (O_2133,N_19290,N_19389);
and UO_2134 (O_2134,N_19892,N_19541);
xor UO_2135 (O_2135,N_19510,N_19274);
nor UO_2136 (O_2136,N_19618,N_19545);
nor UO_2137 (O_2137,N_19649,N_19893);
nor UO_2138 (O_2138,N_19296,N_19417);
nor UO_2139 (O_2139,N_19509,N_19329);
and UO_2140 (O_2140,N_19722,N_19967);
nor UO_2141 (O_2141,N_19524,N_19428);
and UO_2142 (O_2142,N_19869,N_19254);
or UO_2143 (O_2143,N_19930,N_19311);
xnor UO_2144 (O_2144,N_19631,N_19931);
nor UO_2145 (O_2145,N_19689,N_19942);
xor UO_2146 (O_2146,N_19788,N_19459);
nand UO_2147 (O_2147,N_19922,N_19815);
nand UO_2148 (O_2148,N_19682,N_19973);
xor UO_2149 (O_2149,N_19845,N_19290);
nand UO_2150 (O_2150,N_19641,N_19809);
and UO_2151 (O_2151,N_19240,N_19739);
nand UO_2152 (O_2152,N_19731,N_19635);
nand UO_2153 (O_2153,N_19845,N_19784);
nand UO_2154 (O_2154,N_19322,N_19975);
or UO_2155 (O_2155,N_19554,N_19976);
xnor UO_2156 (O_2156,N_19800,N_19231);
xnor UO_2157 (O_2157,N_19990,N_19965);
nand UO_2158 (O_2158,N_19571,N_19986);
or UO_2159 (O_2159,N_19608,N_19833);
and UO_2160 (O_2160,N_19951,N_19661);
xnor UO_2161 (O_2161,N_19721,N_19564);
or UO_2162 (O_2162,N_19332,N_19762);
nor UO_2163 (O_2163,N_19735,N_19998);
and UO_2164 (O_2164,N_19577,N_19521);
nor UO_2165 (O_2165,N_19863,N_19309);
xor UO_2166 (O_2166,N_19371,N_19835);
and UO_2167 (O_2167,N_19406,N_19224);
or UO_2168 (O_2168,N_19935,N_19217);
nor UO_2169 (O_2169,N_19737,N_19488);
nor UO_2170 (O_2170,N_19461,N_19804);
nand UO_2171 (O_2171,N_19664,N_19333);
nand UO_2172 (O_2172,N_19774,N_19527);
and UO_2173 (O_2173,N_19333,N_19513);
or UO_2174 (O_2174,N_19310,N_19247);
and UO_2175 (O_2175,N_19831,N_19562);
or UO_2176 (O_2176,N_19793,N_19678);
nand UO_2177 (O_2177,N_19745,N_19799);
or UO_2178 (O_2178,N_19868,N_19231);
nor UO_2179 (O_2179,N_19879,N_19857);
nor UO_2180 (O_2180,N_19959,N_19917);
nor UO_2181 (O_2181,N_19896,N_19681);
xnor UO_2182 (O_2182,N_19354,N_19519);
nand UO_2183 (O_2183,N_19788,N_19582);
or UO_2184 (O_2184,N_19660,N_19910);
nor UO_2185 (O_2185,N_19440,N_19526);
or UO_2186 (O_2186,N_19797,N_19539);
xnor UO_2187 (O_2187,N_19921,N_19245);
and UO_2188 (O_2188,N_19475,N_19554);
or UO_2189 (O_2189,N_19519,N_19900);
nor UO_2190 (O_2190,N_19327,N_19919);
or UO_2191 (O_2191,N_19973,N_19853);
or UO_2192 (O_2192,N_19228,N_19398);
xor UO_2193 (O_2193,N_19298,N_19740);
nor UO_2194 (O_2194,N_19902,N_19304);
nor UO_2195 (O_2195,N_19634,N_19867);
nand UO_2196 (O_2196,N_19743,N_19836);
nand UO_2197 (O_2197,N_19623,N_19673);
xor UO_2198 (O_2198,N_19223,N_19643);
nor UO_2199 (O_2199,N_19447,N_19544);
and UO_2200 (O_2200,N_19217,N_19279);
or UO_2201 (O_2201,N_19613,N_19548);
nand UO_2202 (O_2202,N_19963,N_19822);
xor UO_2203 (O_2203,N_19779,N_19992);
nand UO_2204 (O_2204,N_19401,N_19319);
nand UO_2205 (O_2205,N_19809,N_19379);
xor UO_2206 (O_2206,N_19589,N_19871);
xor UO_2207 (O_2207,N_19305,N_19847);
xnor UO_2208 (O_2208,N_19616,N_19205);
nand UO_2209 (O_2209,N_19670,N_19755);
nor UO_2210 (O_2210,N_19560,N_19890);
and UO_2211 (O_2211,N_19873,N_19638);
xnor UO_2212 (O_2212,N_19664,N_19352);
nor UO_2213 (O_2213,N_19639,N_19692);
and UO_2214 (O_2214,N_19693,N_19948);
and UO_2215 (O_2215,N_19213,N_19524);
or UO_2216 (O_2216,N_19905,N_19205);
xor UO_2217 (O_2217,N_19612,N_19274);
xnor UO_2218 (O_2218,N_19669,N_19860);
nor UO_2219 (O_2219,N_19649,N_19551);
xor UO_2220 (O_2220,N_19500,N_19481);
and UO_2221 (O_2221,N_19651,N_19678);
xor UO_2222 (O_2222,N_19642,N_19643);
nor UO_2223 (O_2223,N_19459,N_19898);
xnor UO_2224 (O_2224,N_19546,N_19416);
nor UO_2225 (O_2225,N_19497,N_19827);
xnor UO_2226 (O_2226,N_19428,N_19588);
nor UO_2227 (O_2227,N_19689,N_19883);
xor UO_2228 (O_2228,N_19303,N_19404);
and UO_2229 (O_2229,N_19358,N_19383);
and UO_2230 (O_2230,N_19207,N_19446);
nand UO_2231 (O_2231,N_19272,N_19457);
and UO_2232 (O_2232,N_19512,N_19387);
nand UO_2233 (O_2233,N_19797,N_19630);
xor UO_2234 (O_2234,N_19206,N_19437);
or UO_2235 (O_2235,N_19540,N_19582);
xor UO_2236 (O_2236,N_19205,N_19240);
nand UO_2237 (O_2237,N_19947,N_19717);
nor UO_2238 (O_2238,N_19417,N_19754);
xor UO_2239 (O_2239,N_19971,N_19674);
nand UO_2240 (O_2240,N_19349,N_19491);
and UO_2241 (O_2241,N_19333,N_19489);
nor UO_2242 (O_2242,N_19994,N_19817);
xnor UO_2243 (O_2243,N_19604,N_19617);
and UO_2244 (O_2244,N_19385,N_19257);
or UO_2245 (O_2245,N_19216,N_19261);
nor UO_2246 (O_2246,N_19973,N_19415);
or UO_2247 (O_2247,N_19692,N_19994);
nand UO_2248 (O_2248,N_19426,N_19473);
xnor UO_2249 (O_2249,N_19587,N_19364);
or UO_2250 (O_2250,N_19915,N_19515);
or UO_2251 (O_2251,N_19854,N_19295);
nand UO_2252 (O_2252,N_19232,N_19638);
nand UO_2253 (O_2253,N_19510,N_19462);
nand UO_2254 (O_2254,N_19837,N_19907);
nand UO_2255 (O_2255,N_19510,N_19432);
and UO_2256 (O_2256,N_19810,N_19398);
nor UO_2257 (O_2257,N_19931,N_19733);
nand UO_2258 (O_2258,N_19402,N_19252);
nor UO_2259 (O_2259,N_19336,N_19999);
nand UO_2260 (O_2260,N_19545,N_19342);
or UO_2261 (O_2261,N_19399,N_19238);
or UO_2262 (O_2262,N_19785,N_19274);
and UO_2263 (O_2263,N_19512,N_19671);
or UO_2264 (O_2264,N_19390,N_19306);
or UO_2265 (O_2265,N_19469,N_19328);
nand UO_2266 (O_2266,N_19499,N_19940);
nand UO_2267 (O_2267,N_19957,N_19579);
nand UO_2268 (O_2268,N_19437,N_19985);
xor UO_2269 (O_2269,N_19761,N_19667);
nor UO_2270 (O_2270,N_19206,N_19429);
or UO_2271 (O_2271,N_19524,N_19764);
xor UO_2272 (O_2272,N_19745,N_19789);
nand UO_2273 (O_2273,N_19836,N_19329);
and UO_2274 (O_2274,N_19634,N_19230);
and UO_2275 (O_2275,N_19878,N_19915);
nor UO_2276 (O_2276,N_19819,N_19242);
or UO_2277 (O_2277,N_19277,N_19512);
and UO_2278 (O_2278,N_19764,N_19511);
and UO_2279 (O_2279,N_19292,N_19556);
xnor UO_2280 (O_2280,N_19492,N_19985);
and UO_2281 (O_2281,N_19490,N_19666);
xnor UO_2282 (O_2282,N_19683,N_19590);
or UO_2283 (O_2283,N_19439,N_19737);
xnor UO_2284 (O_2284,N_19466,N_19791);
or UO_2285 (O_2285,N_19813,N_19614);
or UO_2286 (O_2286,N_19298,N_19271);
nor UO_2287 (O_2287,N_19244,N_19757);
or UO_2288 (O_2288,N_19814,N_19422);
nand UO_2289 (O_2289,N_19782,N_19631);
xor UO_2290 (O_2290,N_19935,N_19300);
xnor UO_2291 (O_2291,N_19400,N_19417);
nor UO_2292 (O_2292,N_19502,N_19522);
or UO_2293 (O_2293,N_19648,N_19700);
nor UO_2294 (O_2294,N_19973,N_19410);
and UO_2295 (O_2295,N_19705,N_19625);
xor UO_2296 (O_2296,N_19574,N_19810);
and UO_2297 (O_2297,N_19609,N_19389);
or UO_2298 (O_2298,N_19988,N_19780);
or UO_2299 (O_2299,N_19310,N_19589);
and UO_2300 (O_2300,N_19653,N_19598);
or UO_2301 (O_2301,N_19236,N_19654);
xor UO_2302 (O_2302,N_19847,N_19997);
xor UO_2303 (O_2303,N_19983,N_19596);
nor UO_2304 (O_2304,N_19367,N_19268);
xor UO_2305 (O_2305,N_19687,N_19578);
nor UO_2306 (O_2306,N_19979,N_19265);
nand UO_2307 (O_2307,N_19251,N_19285);
and UO_2308 (O_2308,N_19305,N_19660);
nand UO_2309 (O_2309,N_19539,N_19777);
nor UO_2310 (O_2310,N_19877,N_19493);
nand UO_2311 (O_2311,N_19315,N_19959);
nor UO_2312 (O_2312,N_19643,N_19292);
xor UO_2313 (O_2313,N_19238,N_19389);
nand UO_2314 (O_2314,N_19690,N_19422);
and UO_2315 (O_2315,N_19659,N_19540);
nand UO_2316 (O_2316,N_19649,N_19238);
nor UO_2317 (O_2317,N_19299,N_19256);
and UO_2318 (O_2318,N_19430,N_19663);
xor UO_2319 (O_2319,N_19963,N_19546);
or UO_2320 (O_2320,N_19416,N_19934);
xnor UO_2321 (O_2321,N_19833,N_19637);
nor UO_2322 (O_2322,N_19642,N_19744);
nor UO_2323 (O_2323,N_19419,N_19588);
xor UO_2324 (O_2324,N_19563,N_19862);
nand UO_2325 (O_2325,N_19300,N_19998);
xor UO_2326 (O_2326,N_19304,N_19352);
nand UO_2327 (O_2327,N_19974,N_19439);
nor UO_2328 (O_2328,N_19270,N_19299);
and UO_2329 (O_2329,N_19927,N_19500);
nor UO_2330 (O_2330,N_19504,N_19883);
or UO_2331 (O_2331,N_19781,N_19489);
nand UO_2332 (O_2332,N_19419,N_19558);
nand UO_2333 (O_2333,N_19908,N_19546);
or UO_2334 (O_2334,N_19717,N_19581);
nand UO_2335 (O_2335,N_19899,N_19688);
nor UO_2336 (O_2336,N_19907,N_19733);
and UO_2337 (O_2337,N_19412,N_19674);
or UO_2338 (O_2338,N_19363,N_19907);
nor UO_2339 (O_2339,N_19693,N_19774);
nor UO_2340 (O_2340,N_19374,N_19964);
and UO_2341 (O_2341,N_19663,N_19776);
nand UO_2342 (O_2342,N_19795,N_19343);
nand UO_2343 (O_2343,N_19480,N_19827);
xnor UO_2344 (O_2344,N_19321,N_19268);
and UO_2345 (O_2345,N_19770,N_19743);
and UO_2346 (O_2346,N_19336,N_19962);
nand UO_2347 (O_2347,N_19314,N_19301);
and UO_2348 (O_2348,N_19322,N_19943);
and UO_2349 (O_2349,N_19540,N_19306);
nor UO_2350 (O_2350,N_19810,N_19774);
nor UO_2351 (O_2351,N_19264,N_19830);
and UO_2352 (O_2352,N_19407,N_19658);
or UO_2353 (O_2353,N_19634,N_19236);
or UO_2354 (O_2354,N_19311,N_19542);
or UO_2355 (O_2355,N_19418,N_19836);
nor UO_2356 (O_2356,N_19837,N_19952);
or UO_2357 (O_2357,N_19679,N_19877);
xnor UO_2358 (O_2358,N_19545,N_19895);
or UO_2359 (O_2359,N_19406,N_19236);
nor UO_2360 (O_2360,N_19887,N_19410);
xnor UO_2361 (O_2361,N_19988,N_19222);
xnor UO_2362 (O_2362,N_19458,N_19327);
and UO_2363 (O_2363,N_19406,N_19206);
nor UO_2364 (O_2364,N_19984,N_19977);
nand UO_2365 (O_2365,N_19255,N_19798);
nor UO_2366 (O_2366,N_19454,N_19497);
xor UO_2367 (O_2367,N_19958,N_19334);
nand UO_2368 (O_2368,N_19767,N_19373);
and UO_2369 (O_2369,N_19845,N_19724);
or UO_2370 (O_2370,N_19611,N_19489);
nor UO_2371 (O_2371,N_19864,N_19787);
nor UO_2372 (O_2372,N_19953,N_19360);
nor UO_2373 (O_2373,N_19772,N_19745);
nor UO_2374 (O_2374,N_19366,N_19458);
xnor UO_2375 (O_2375,N_19308,N_19626);
and UO_2376 (O_2376,N_19782,N_19558);
or UO_2377 (O_2377,N_19577,N_19344);
or UO_2378 (O_2378,N_19871,N_19536);
or UO_2379 (O_2379,N_19914,N_19287);
xor UO_2380 (O_2380,N_19289,N_19447);
nor UO_2381 (O_2381,N_19692,N_19679);
nand UO_2382 (O_2382,N_19862,N_19208);
or UO_2383 (O_2383,N_19578,N_19359);
xor UO_2384 (O_2384,N_19729,N_19295);
nor UO_2385 (O_2385,N_19613,N_19579);
xor UO_2386 (O_2386,N_19790,N_19209);
xnor UO_2387 (O_2387,N_19686,N_19751);
or UO_2388 (O_2388,N_19930,N_19941);
nor UO_2389 (O_2389,N_19342,N_19990);
and UO_2390 (O_2390,N_19654,N_19847);
and UO_2391 (O_2391,N_19520,N_19371);
or UO_2392 (O_2392,N_19374,N_19976);
nand UO_2393 (O_2393,N_19524,N_19886);
and UO_2394 (O_2394,N_19959,N_19736);
or UO_2395 (O_2395,N_19535,N_19282);
xnor UO_2396 (O_2396,N_19735,N_19411);
xnor UO_2397 (O_2397,N_19772,N_19790);
nor UO_2398 (O_2398,N_19271,N_19669);
xor UO_2399 (O_2399,N_19881,N_19908);
or UO_2400 (O_2400,N_19583,N_19909);
nor UO_2401 (O_2401,N_19697,N_19487);
nand UO_2402 (O_2402,N_19575,N_19864);
nand UO_2403 (O_2403,N_19334,N_19747);
nor UO_2404 (O_2404,N_19463,N_19640);
nor UO_2405 (O_2405,N_19595,N_19838);
and UO_2406 (O_2406,N_19457,N_19692);
xor UO_2407 (O_2407,N_19794,N_19427);
or UO_2408 (O_2408,N_19373,N_19471);
and UO_2409 (O_2409,N_19382,N_19751);
or UO_2410 (O_2410,N_19420,N_19442);
and UO_2411 (O_2411,N_19423,N_19951);
nor UO_2412 (O_2412,N_19894,N_19749);
and UO_2413 (O_2413,N_19359,N_19528);
xnor UO_2414 (O_2414,N_19509,N_19627);
nand UO_2415 (O_2415,N_19866,N_19672);
nand UO_2416 (O_2416,N_19639,N_19691);
and UO_2417 (O_2417,N_19472,N_19730);
and UO_2418 (O_2418,N_19532,N_19201);
or UO_2419 (O_2419,N_19325,N_19807);
xnor UO_2420 (O_2420,N_19309,N_19303);
xor UO_2421 (O_2421,N_19935,N_19856);
xor UO_2422 (O_2422,N_19562,N_19880);
xor UO_2423 (O_2423,N_19913,N_19434);
nor UO_2424 (O_2424,N_19895,N_19729);
and UO_2425 (O_2425,N_19667,N_19811);
and UO_2426 (O_2426,N_19276,N_19621);
xor UO_2427 (O_2427,N_19660,N_19846);
xnor UO_2428 (O_2428,N_19595,N_19227);
xor UO_2429 (O_2429,N_19992,N_19673);
xor UO_2430 (O_2430,N_19681,N_19526);
or UO_2431 (O_2431,N_19883,N_19428);
nor UO_2432 (O_2432,N_19358,N_19460);
xnor UO_2433 (O_2433,N_19618,N_19925);
nand UO_2434 (O_2434,N_19905,N_19537);
and UO_2435 (O_2435,N_19808,N_19296);
or UO_2436 (O_2436,N_19638,N_19353);
nor UO_2437 (O_2437,N_19735,N_19353);
nand UO_2438 (O_2438,N_19949,N_19486);
nor UO_2439 (O_2439,N_19392,N_19244);
xnor UO_2440 (O_2440,N_19930,N_19515);
nand UO_2441 (O_2441,N_19677,N_19602);
and UO_2442 (O_2442,N_19262,N_19705);
nand UO_2443 (O_2443,N_19643,N_19664);
nor UO_2444 (O_2444,N_19658,N_19273);
nand UO_2445 (O_2445,N_19872,N_19676);
xor UO_2446 (O_2446,N_19666,N_19618);
and UO_2447 (O_2447,N_19873,N_19519);
and UO_2448 (O_2448,N_19323,N_19213);
nand UO_2449 (O_2449,N_19603,N_19499);
nand UO_2450 (O_2450,N_19481,N_19833);
or UO_2451 (O_2451,N_19738,N_19269);
xnor UO_2452 (O_2452,N_19941,N_19782);
nor UO_2453 (O_2453,N_19223,N_19462);
xor UO_2454 (O_2454,N_19468,N_19559);
nor UO_2455 (O_2455,N_19437,N_19459);
nor UO_2456 (O_2456,N_19810,N_19309);
xor UO_2457 (O_2457,N_19298,N_19213);
or UO_2458 (O_2458,N_19605,N_19284);
nor UO_2459 (O_2459,N_19639,N_19803);
or UO_2460 (O_2460,N_19254,N_19666);
xor UO_2461 (O_2461,N_19959,N_19758);
and UO_2462 (O_2462,N_19286,N_19760);
xnor UO_2463 (O_2463,N_19380,N_19704);
or UO_2464 (O_2464,N_19293,N_19456);
and UO_2465 (O_2465,N_19674,N_19797);
xor UO_2466 (O_2466,N_19764,N_19774);
xor UO_2467 (O_2467,N_19793,N_19534);
or UO_2468 (O_2468,N_19545,N_19297);
and UO_2469 (O_2469,N_19819,N_19234);
nor UO_2470 (O_2470,N_19844,N_19669);
nand UO_2471 (O_2471,N_19942,N_19904);
nand UO_2472 (O_2472,N_19229,N_19826);
and UO_2473 (O_2473,N_19889,N_19383);
nor UO_2474 (O_2474,N_19417,N_19926);
xnor UO_2475 (O_2475,N_19744,N_19758);
or UO_2476 (O_2476,N_19689,N_19402);
or UO_2477 (O_2477,N_19751,N_19512);
nand UO_2478 (O_2478,N_19698,N_19297);
xnor UO_2479 (O_2479,N_19312,N_19991);
xnor UO_2480 (O_2480,N_19325,N_19740);
nand UO_2481 (O_2481,N_19753,N_19846);
nor UO_2482 (O_2482,N_19864,N_19959);
and UO_2483 (O_2483,N_19719,N_19267);
xnor UO_2484 (O_2484,N_19612,N_19698);
and UO_2485 (O_2485,N_19515,N_19849);
nor UO_2486 (O_2486,N_19301,N_19927);
or UO_2487 (O_2487,N_19453,N_19888);
or UO_2488 (O_2488,N_19372,N_19791);
or UO_2489 (O_2489,N_19742,N_19615);
or UO_2490 (O_2490,N_19605,N_19487);
and UO_2491 (O_2491,N_19686,N_19656);
or UO_2492 (O_2492,N_19927,N_19205);
nand UO_2493 (O_2493,N_19878,N_19356);
or UO_2494 (O_2494,N_19622,N_19269);
and UO_2495 (O_2495,N_19988,N_19824);
xnor UO_2496 (O_2496,N_19841,N_19993);
nand UO_2497 (O_2497,N_19645,N_19904);
xor UO_2498 (O_2498,N_19455,N_19565);
or UO_2499 (O_2499,N_19305,N_19860);
endmodule