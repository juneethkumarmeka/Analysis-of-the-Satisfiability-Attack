module basic_1000_10000_1500_5_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_311,In_143);
nor U1 (N_1,In_275,In_90);
nand U2 (N_2,In_641,In_11);
or U3 (N_3,In_262,In_452);
nand U4 (N_4,In_764,In_729);
or U5 (N_5,In_328,In_897);
nand U6 (N_6,In_617,In_356);
nor U7 (N_7,In_360,In_125);
and U8 (N_8,In_997,In_248);
and U9 (N_9,In_964,In_765);
and U10 (N_10,In_166,In_514);
nor U11 (N_11,In_760,In_198);
nor U12 (N_12,In_483,In_538);
xor U13 (N_13,In_464,In_367);
and U14 (N_14,In_106,In_379);
and U15 (N_15,In_861,In_722);
and U16 (N_16,In_841,In_324);
nand U17 (N_17,In_104,In_305);
or U18 (N_18,In_644,In_107);
or U19 (N_19,In_96,In_698);
and U20 (N_20,In_315,In_974);
nor U21 (N_21,In_346,In_185);
or U22 (N_22,In_286,In_419);
and U23 (N_23,In_3,In_173);
and U24 (N_24,In_884,In_591);
and U25 (N_25,In_774,In_694);
and U26 (N_26,In_444,In_905);
xor U27 (N_27,In_755,In_81);
or U28 (N_28,In_562,In_622);
or U29 (N_29,In_500,In_706);
or U30 (N_30,In_188,In_416);
nor U31 (N_31,In_880,In_256);
nor U32 (N_32,In_522,In_136);
nand U33 (N_33,In_231,In_0);
and U34 (N_34,In_121,In_737);
nand U35 (N_35,In_882,In_909);
and U36 (N_36,In_517,In_68);
and U37 (N_37,In_948,In_359);
or U38 (N_38,In_469,In_254);
nor U39 (N_39,In_624,In_886);
nand U40 (N_40,In_128,In_17);
nand U41 (N_41,In_684,In_314);
or U42 (N_42,In_648,In_21);
nor U43 (N_43,In_708,In_931);
or U44 (N_44,In_885,In_508);
or U45 (N_45,In_425,In_131);
or U46 (N_46,In_609,In_775);
nor U47 (N_47,In_352,In_281);
nor U48 (N_48,In_656,In_435);
and U49 (N_49,In_977,In_811);
and U50 (N_50,In_716,In_134);
nand U51 (N_51,In_900,In_815);
nand U52 (N_52,In_25,In_879);
nor U53 (N_53,In_747,In_97);
nor U54 (N_54,In_877,In_678);
nor U55 (N_55,In_37,In_441);
and U56 (N_56,In_368,In_671);
and U57 (N_57,In_232,In_692);
nor U58 (N_58,In_200,In_849);
or U59 (N_59,In_734,In_763);
nand U60 (N_60,In_126,In_992);
nand U61 (N_61,In_544,In_851);
and U62 (N_62,In_753,In_109);
nand U63 (N_63,In_345,In_280);
xor U64 (N_64,In_957,In_318);
or U65 (N_65,In_389,In_610);
nand U66 (N_66,In_975,In_146);
nor U67 (N_67,In_285,In_902);
or U68 (N_68,In_525,In_284);
nor U69 (N_69,In_654,In_291);
nor U70 (N_70,In_904,In_825);
nand U71 (N_71,In_250,In_92);
or U72 (N_72,In_963,In_294);
or U73 (N_73,In_767,In_414);
nand U74 (N_74,In_167,In_968);
nand U75 (N_75,In_741,In_383);
nor U76 (N_76,In_601,In_862);
nand U77 (N_77,In_224,In_647);
and U78 (N_78,In_307,In_502);
nand U79 (N_79,In_940,In_989);
and U80 (N_80,In_440,In_703);
and U81 (N_81,In_41,In_803);
nor U82 (N_82,In_182,In_130);
nor U83 (N_83,In_1,In_55);
and U84 (N_84,In_939,In_377);
nor U85 (N_85,In_530,In_553);
or U86 (N_86,In_789,In_349);
and U87 (N_87,In_567,In_987);
and U88 (N_88,In_829,In_986);
and U89 (N_89,In_43,In_251);
nor U90 (N_90,In_407,In_757);
or U91 (N_91,In_269,In_523);
nand U92 (N_92,In_924,In_691);
nand U93 (N_93,In_598,In_18);
and U94 (N_94,In_582,In_667);
nor U95 (N_95,In_702,In_421);
nand U96 (N_96,In_898,In_922);
nor U97 (N_97,In_463,In_268);
nand U98 (N_98,In_621,In_32);
and U99 (N_99,In_586,In_850);
or U100 (N_100,In_181,In_216);
or U101 (N_101,In_215,In_101);
xnor U102 (N_102,In_645,In_679);
nor U103 (N_103,In_661,In_381);
or U104 (N_104,In_50,In_405);
nor U105 (N_105,In_744,In_242);
nor U106 (N_106,In_959,In_670);
or U107 (N_107,In_20,In_347);
nand U108 (N_108,In_29,In_852);
or U109 (N_109,In_631,In_329);
nor U110 (N_110,In_921,In_265);
nor U111 (N_111,In_933,In_701);
or U112 (N_112,In_739,In_245);
or U113 (N_113,In_48,In_298);
nand U114 (N_114,In_154,In_344);
and U115 (N_115,In_990,In_267);
nand U116 (N_116,In_149,In_445);
nor U117 (N_117,In_846,In_552);
and U118 (N_118,In_855,In_260);
nor U119 (N_119,In_161,In_779);
nand U120 (N_120,In_496,In_548);
nand U121 (N_121,In_599,In_838);
nor U122 (N_122,In_300,In_579);
xor U123 (N_123,In_778,In_836);
or U124 (N_124,In_791,In_459);
nand U125 (N_125,In_370,In_30);
nor U126 (N_126,In_369,In_222);
and U127 (N_127,In_949,In_273);
xor U128 (N_128,In_63,In_685);
or U129 (N_129,In_816,In_881);
or U130 (N_130,In_213,In_390);
nor U131 (N_131,In_235,In_287);
nand U132 (N_132,In_587,In_279);
and U133 (N_133,In_341,In_124);
and U134 (N_134,In_353,In_745);
and U135 (N_135,In_145,In_354);
xnor U136 (N_136,In_82,In_72);
nand U137 (N_137,In_332,In_288);
or U138 (N_138,In_944,In_433);
nand U139 (N_139,In_114,In_664);
and U140 (N_140,In_613,In_427);
or U141 (N_141,In_833,In_434);
or U142 (N_142,In_961,In_535);
and U143 (N_143,In_906,In_313);
or U144 (N_144,In_488,In_302);
nor U145 (N_145,In_704,In_208);
and U146 (N_146,In_118,In_66);
nand U147 (N_147,In_74,In_214);
nor U148 (N_148,In_770,In_929);
nand U149 (N_149,In_603,In_272);
or U150 (N_150,In_516,In_777);
xnor U151 (N_151,In_142,In_657);
nor U152 (N_152,In_958,In_558);
nor U153 (N_153,In_925,In_863);
nor U154 (N_154,In_804,In_955);
or U155 (N_155,In_785,In_627);
nor U156 (N_156,In_823,In_282);
nor U157 (N_157,In_511,In_355);
nor U158 (N_158,In_477,In_27);
nor U159 (N_159,In_67,In_781);
nand U160 (N_160,In_720,In_953);
and U161 (N_161,In_388,In_391);
or U162 (N_162,In_330,In_636);
nand U163 (N_163,In_787,In_759);
nand U164 (N_164,In_301,In_809);
nand U165 (N_165,In_162,In_653);
nand U166 (N_166,In_362,In_962);
xnor U167 (N_167,In_930,In_643);
nor U168 (N_168,In_190,In_283);
nor U169 (N_169,In_218,In_799);
xor U170 (N_170,In_192,In_828);
xor U171 (N_171,In_699,In_910);
nand U172 (N_172,In_139,In_151);
nand U173 (N_173,In_526,In_270);
xor U174 (N_174,In_675,In_874);
nor U175 (N_175,In_420,In_818);
or U176 (N_176,In_883,In_77);
nand U177 (N_177,In_144,In_481);
xor U178 (N_178,In_731,In_545);
nand U179 (N_179,In_709,In_70);
and U180 (N_180,In_174,In_163);
nand U181 (N_181,In_732,In_650);
nor U182 (N_182,In_61,In_674);
xor U183 (N_183,In_864,In_527);
xnor U184 (N_184,In_506,In_334);
nor U185 (N_185,In_339,In_768);
and U186 (N_186,In_533,In_393);
and U187 (N_187,In_386,In_663);
nand U188 (N_188,In_927,In_689);
nor U189 (N_189,In_292,In_264);
nor U190 (N_190,In_687,In_396);
nand U191 (N_191,In_394,In_220);
and U192 (N_192,In_229,In_872);
or U193 (N_193,In_539,In_476);
nand U194 (N_194,In_537,In_659);
or U195 (N_195,In_19,In_91);
or U196 (N_196,In_711,In_518);
nand U197 (N_197,In_998,In_385);
and U198 (N_198,In_39,In_310);
nand U199 (N_199,In_683,In_333);
and U200 (N_200,In_697,In_395);
or U201 (N_201,In_261,In_404);
nand U202 (N_202,In_856,In_903);
or U203 (N_203,In_531,In_98);
nand U204 (N_204,In_71,In_503);
and U205 (N_205,In_750,In_596);
nor U206 (N_206,In_164,In_680);
nand U207 (N_207,In_542,In_295);
nor U208 (N_208,In_171,In_465);
and U209 (N_209,In_569,In_723);
nand U210 (N_210,In_871,In_597);
nor U211 (N_211,In_802,In_954);
xnor U212 (N_212,In_9,In_608);
nand U213 (N_213,In_263,In_618);
or U214 (N_214,In_822,In_917);
xnor U215 (N_215,In_640,In_868);
nor U216 (N_216,In_150,In_202);
and U217 (N_217,In_195,In_210);
and U218 (N_218,In_387,In_102);
nor U219 (N_219,In_797,In_918);
and U220 (N_220,In_493,In_935);
nand U221 (N_221,In_632,In_588);
or U222 (N_222,In_448,In_782);
or U223 (N_223,In_730,In_411);
nor U224 (N_224,In_110,In_480);
nor U225 (N_225,In_946,In_155);
or U226 (N_226,In_695,In_572);
xnor U227 (N_227,In_672,In_570);
or U228 (N_228,In_176,In_637);
or U229 (N_229,In_605,In_956);
nor U230 (N_230,In_365,In_783);
or U231 (N_231,In_297,In_616);
or U232 (N_232,In_13,In_60);
or U233 (N_233,In_913,In_400);
and U234 (N_234,In_62,In_983);
xnor U235 (N_235,In_509,In_374);
and U236 (N_236,In_230,In_304);
or U237 (N_237,In_893,In_510);
and U238 (N_238,In_186,In_555);
and U239 (N_239,In_380,In_338);
and U240 (N_240,In_619,In_358);
nor U241 (N_241,In_688,In_331);
xor U242 (N_242,In_715,In_247);
and U243 (N_243,In_923,In_132);
nor U244 (N_244,In_988,In_57);
xor U245 (N_245,In_157,In_119);
nor U246 (N_246,In_458,In_65);
nor U247 (N_247,In_187,In_498);
nand U248 (N_248,In_470,In_981);
and U249 (N_249,In_950,In_141);
nand U250 (N_250,In_583,In_576);
nand U251 (N_251,In_436,In_446);
or U252 (N_252,In_515,In_169);
xnor U253 (N_253,In_914,In_221);
or U254 (N_254,In_575,In_225);
nand U255 (N_255,In_726,In_205);
nor U256 (N_256,In_889,In_201);
nand U257 (N_257,In_348,In_912);
or U258 (N_258,In_842,In_375);
nand U259 (N_259,In_258,In_8);
xnor U260 (N_260,In_994,In_122);
nor U261 (N_261,In_865,In_489);
or U262 (N_262,In_473,In_630);
nand U263 (N_263,In_494,In_499);
or U264 (N_264,In_372,In_505);
nor U265 (N_265,In_762,In_528);
xor U266 (N_266,In_554,In_456);
nor U267 (N_267,In_309,In_54);
nand U268 (N_268,In_581,In_159);
or U269 (N_269,In_742,In_993);
nor U270 (N_270,In_660,In_108);
xnor U271 (N_271,In_795,In_28);
and U272 (N_272,In_415,In_308);
and U273 (N_273,In_651,In_978);
nand U274 (N_274,In_976,In_79);
xnor U275 (N_275,In_487,In_551);
and U276 (N_276,In_233,In_123);
nor U277 (N_277,In_86,In_180);
nor U278 (N_278,In_42,In_758);
nand U279 (N_279,In_397,In_491);
xor U280 (N_280,In_87,In_669);
xnor U281 (N_281,In_826,In_289);
nand U282 (N_282,In_46,In_867);
and U283 (N_283,In_869,In_177);
and U284 (N_284,In_769,In_454);
nor U285 (N_285,In_343,In_735);
nor U286 (N_286,In_662,In_100);
and U287 (N_287,In_271,In_501);
nor U288 (N_288,In_634,In_830);
nor U289 (N_289,In_580,In_253);
xnor U290 (N_290,In_129,In_746);
nor U291 (N_291,In_814,In_932);
or U292 (N_292,In_686,In_529);
and U293 (N_293,In_320,In_969);
and U294 (N_294,In_590,In_47);
nand U295 (N_295,In_761,In_724);
or U296 (N_296,In_147,In_999);
nand U297 (N_297,In_199,In_784);
nor U298 (N_298,In_890,In_813);
nand U299 (N_299,In_403,In_942);
or U300 (N_300,In_408,In_547);
nor U301 (N_301,In_478,In_629);
nor U302 (N_302,In_15,In_728);
nand U303 (N_303,In_943,In_409);
and U304 (N_304,In_626,In_497);
or U305 (N_305,In_357,In_342);
or U306 (N_306,In_252,In_431);
nand U307 (N_307,In_519,In_73);
nand U308 (N_308,In_22,In_455);
nor U309 (N_309,In_95,In_982);
nor U310 (N_310,In_371,In_524);
and U311 (N_311,In_602,In_960);
and U312 (N_312,In_749,In_193);
or U313 (N_313,In_540,In_873);
or U314 (N_314,In_69,In_751);
nand U315 (N_315,In_277,In_772);
nand U316 (N_316,In_594,In_457);
xnor U317 (N_317,In_592,In_36);
or U318 (N_318,In_490,In_549);
nor U319 (N_319,In_668,In_59);
and U320 (N_320,In_475,In_866);
xnor U321 (N_321,In_76,In_839);
and U322 (N_322,In_392,In_449);
or U323 (N_323,In_156,In_895);
and U324 (N_324,In_340,In_725);
nor U325 (N_325,In_844,In_351);
nand U326 (N_326,In_399,In_936);
nor U327 (N_327,In_85,In_585);
and U328 (N_328,In_740,In_89);
nand U329 (N_329,In_401,In_612);
xnor U330 (N_330,In_424,In_361);
nor U331 (N_331,In_807,In_6);
xnor U332 (N_332,In_713,In_543);
xor U333 (N_333,In_607,In_557);
nor U334 (N_334,In_299,In_696);
and U335 (N_335,In_259,In_94);
nand U336 (N_336,In_113,In_211);
or U337 (N_337,In_373,In_565);
or U338 (N_338,In_952,In_4);
nor U339 (N_339,In_207,In_165);
nor U340 (N_340,In_550,In_12);
or U341 (N_341,In_771,In_103);
nand U342 (N_342,In_450,In_615);
and U343 (N_343,In_817,In_705);
or U344 (N_344,In_26,In_135);
and U345 (N_345,In_120,In_241);
nand U346 (N_346,In_422,In_203);
nand U347 (N_347,In_428,In_158);
or U348 (N_348,In_707,In_137);
and U349 (N_349,In_366,In_901);
xnor U350 (N_350,In_209,In_296);
or U351 (N_351,In_563,In_160);
and U352 (N_352,In_337,In_875);
and U353 (N_353,In_788,In_183);
or U354 (N_354,In_584,In_316);
xnor U355 (N_355,In_564,In_655);
nor U356 (N_356,In_153,In_801);
nand U357 (N_357,In_832,In_593);
nand U358 (N_358,In_835,In_33);
xnor U359 (N_359,In_467,In_363);
or U360 (N_360,In_892,In_513);
and U361 (N_361,In_93,In_278);
or U362 (N_362,In_853,In_541);
nor U363 (N_363,In_571,In_561);
and U364 (N_364,In_38,In_532);
xnor U365 (N_365,In_733,In_168);
nand U366 (N_366,In_718,In_468);
and U367 (N_367,In_894,In_14);
and U368 (N_368,In_611,In_717);
nand U369 (N_369,In_521,In_520);
nor U370 (N_370,In_335,In_888);
and U371 (N_371,In_620,In_152);
or U372 (N_372,In_53,In_824);
nand U373 (N_373,In_238,In_236);
nand U374 (N_374,In_577,In_682);
and U375 (N_375,In_870,In_443);
xor U376 (N_376,In_748,In_951);
xnor U377 (N_377,In_10,In_984);
nor U378 (N_378,In_430,In_973);
nor U379 (N_379,In_719,In_5);
xnor U380 (N_380,In_736,In_980);
or U381 (N_381,In_255,In_451);
nor U382 (N_382,In_827,In_796);
and U383 (N_383,In_907,In_402);
nand U384 (N_384,In_878,In_138);
and U385 (N_385,In_854,In_479);
nand U386 (N_386,In_376,In_274);
and U387 (N_387,In_721,In_820);
xnor U388 (N_388,In_325,In_116);
or U389 (N_389,In_752,In_507);
nand U390 (N_390,In_321,In_859);
and U391 (N_391,In_382,In_223);
nor U392 (N_392,In_23,In_574);
or U393 (N_393,In_996,In_447);
nor U394 (N_394,In_559,In_536);
xor U395 (N_395,In_712,In_84);
or U396 (N_396,In_217,In_112);
and U397 (N_397,In_58,In_423);
and U398 (N_398,In_681,In_714);
xnor U399 (N_399,In_56,In_410);
xnor U400 (N_400,In_972,In_945);
or U401 (N_401,In_437,In_673);
or U402 (N_402,In_111,In_776);
xnor U403 (N_403,In_676,In_896);
and U404 (N_404,In_319,In_64);
nor U405 (N_405,In_237,In_226);
nand U406 (N_406,In_908,In_947);
nor U407 (N_407,In_115,In_504);
and U408 (N_408,In_495,In_556);
or U409 (N_409,In_600,In_7);
and U410 (N_410,In_44,In_633);
nand U411 (N_411,In_858,In_244);
xor U412 (N_412,In_418,In_196);
or U413 (N_413,In_170,In_738);
or U414 (N_414,In_840,In_995);
nor U415 (N_415,In_398,In_303);
or U416 (N_416,In_614,In_234);
or U417 (N_417,In_486,In_812);
nor U418 (N_418,In_665,In_638);
nor U419 (N_419,In_628,In_926);
or U420 (N_420,In_140,In_336);
nor U421 (N_421,In_249,In_798);
nor U422 (N_422,In_189,In_184);
nand U423 (N_423,In_899,In_911);
nor U424 (N_424,In_228,In_792);
or U425 (N_425,In_327,In_790);
nand U426 (N_426,In_240,In_805);
xnor U427 (N_427,In_642,In_276);
or U428 (N_428,In_646,In_652);
nor U429 (N_429,In_179,In_40);
or U430 (N_430,In_442,In_364);
nor U431 (N_431,In_49,In_293);
nand U432 (N_432,In_306,In_413);
and U433 (N_433,In_589,In_172);
or U434 (N_434,In_378,In_246);
xor U435 (N_435,In_710,In_384);
xor U436 (N_436,In_985,In_312);
nor U437 (N_437,In_800,In_406);
nor U438 (N_438,In_78,In_290);
xor U439 (N_439,In_970,In_677);
nor U440 (N_440,In_604,In_821);
nand U441 (N_441,In_492,In_916);
or U442 (N_442,In_52,In_639);
or U443 (N_443,In_915,In_808);
xnor U444 (N_444,In_16,In_474);
or U445 (N_445,In_239,In_560);
nor U446 (N_446,In_266,In_834);
nand U447 (N_447,In_460,In_810);
nand U448 (N_448,In_928,In_243);
nor U449 (N_449,In_831,In_595);
or U450 (N_450,In_690,In_649);
or U451 (N_451,In_566,In_578);
nand U452 (N_452,In_31,In_573);
and U453 (N_453,In_991,In_979);
nor U454 (N_454,In_461,In_432);
nand U455 (N_455,In_227,In_472);
xor U456 (N_456,In_848,In_219);
or U457 (N_457,In_99,In_453);
or U458 (N_458,In_965,In_204);
nor U459 (N_459,In_773,In_105);
xnor U460 (N_460,In_756,In_485);
and U461 (N_461,In_466,In_780);
or U462 (N_462,In_133,In_786);
and U463 (N_463,In_257,In_766);
xor U464 (N_464,In_2,In_806);
nand U465 (N_465,In_794,In_971);
nand U466 (N_466,In_666,In_45);
nor U467 (N_467,In_793,In_471);
xnor U468 (N_468,In_819,In_568);
and U469 (N_469,In_484,In_887);
nor U470 (N_470,In_857,In_920);
nand U471 (N_471,In_512,In_919);
nand U472 (N_472,In_727,In_941);
nand U473 (N_473,In_412,In_837);
or U474 (N_474,In_658,In_326);
nand U475 (N_475,In_178,In_606);
or U476 (N_476,In_194,In_117);
and U477 (N_477,In_876,In_482);
and U478 (N_478,In_350,In_426);
or U479 (N_479,In_743,In_625);
nand U480 (N_480,In_546,In_323);
and U481 (N_481,In_212,In_937);
nand U482 (N_482,In_317,In_148);
and U483 (N_483,In_206,In_623);
nor U484 (N_484,In_75,In_35);
or U485 (N_485,In_80,In_934);
xnor U486 (N_486,In_845,In_462);
nand U487 (N_487,In_175,In_127);
nor U488 (N_488,In_24,In_197);
nand U489 (N_489,In_88,In_322);
nor U490 (N_490,In_417,In_51);
and U491 (N_491,In_429,In_438);
and U492 (N_492,In_191,In_700);
nand U493 (N_493,In_83,In_635);
or U494 (N_494,In_754,In_966);
or U495 (N_495,In_439,In_967);
or U496 (N_496,In_891,In_938);
nand U497 (N_497,In_693,In_534);
and U498 (N_498,In_860,In_34);
or U499 (N_499,In_843,In_847);
and U500 (N_500,In_870,In_778);
nand U501 (N_501,In_856,In_419);
or U502 (N_502,In_584,In_475);
nand U503 (N_503,In_707,In_677);
or U504 (N_504,In_62,In_605);
and U505 (N_505,In_136,In_639);
nand U506 (N_506,In_220,In_827);
or U507 (N_507,In_702,In_460);
and U508 (N_508,In_530,In_286);
nor U509 (N_509,In_191,In_885);
xor U510 (N_510,In_19,In_389);
nor U511 (N_511,In_649,In_309);
and U512 (N_512,In_906,In_810);
and U513 (N_513,In_891,In_261);
nor U514 (N_514,In_367,In_270);
nand U515 (N_515,In_603,In_828);
nand U516 (N_516,In_347,In_699);
nand U517 (N_517,In_409,In_682);
nor U518 (N_518,In_27,In_252);
nand U519 (N_519,In_360,In_807);
or U520 (N_520,In_494,In_83);
nor U521 (N_521,In_793,In_581);
nor U522 (N_522,In_748,In_105);
nor U523 (N_523,In_860,In_598);
nor U524 (N_524,In_580,In_286);
or U525 (N_525,In_279,In_948);
nand U526 (N_526,In_636,In_19);
or U527 (N_527,In_775,In_770);
or U528 (N_528,In_394,In_173);
and U529 (N_529,In_95,In_298);
or U530 (N_530,In_122,In_773);
nor U531 (N_531,In_539,In_569);
or U532 (N_532,In_840,In_357);
nand U533 (N_533,In_821,In_214);
or U534 (N_534,In_514,In_55);
nor U535 (N_535,In_194,In_601);
or U536 (N_536,In_171,In_141);
or U537 (N_537,In_859,In_702);
and U538 (N_538,In_527,In_809);
or U539 (N_539,In_853,In_889);
xor U540 (N_540,In_831,In_661);
or U541 (N_541,In_139,In_315);
and U542 (N_542,In_774,In_176);
and U543 (N_543,In_857,In_136);
nor U544 (N_544,In_960,In_699);
and U545 (N_545,In_840,In_495);
nor U546 (N_546,In_185,In_64);
nor U547 (N_547,In_381,In_710);
or U548 (N_548,In_932,In_380);
or U549 (N_549,In_919,In_336);
or U550 (N_550,In_731,In_617);
and U551 (N_551,In_671,In_224);
nor U552 (N_552,In_281,In_773);
nor U553 (N_553,In_736,In_60);
nor U554 (N_554,In_335,In_989);
nand U555 (N_555,In_364,In_188);
nor U556 (N_556,In_756,In_730);
or U557 (N_557,In_857,In_655);
and U558 (N_558,In_753,In_920);
nor U559 (N_559,In_605,In_250);
nand U560 (N_560,In_638,In_184);
and U561 (N_561,In_887,In_917);
nor U562 (N_562,In_214,In_491);
and U563 (N_563,In_886,In_518);
and U564 (N_564,In_198,In_451);
or U565 (N_565,In_441,In_260);
and U566 (N_566,In_105,In_486);
nand U567 (N_567,In_779,In_329);
xnor U568 (N_568,In_442,In_473);
xor U569 (N_569,In_146,In_253);
nand U570 (N_570,In_86,In_783);
nor U571 (N_571,In_233,In_692);
nand U572 (N_572,In_938,In_352);
and U573 (N_573,In_212,In_834);
and U574 (N_574,In_334,In_137);
nor U575 (N_575,In_683,In_589);
nand U576 (N_576,In_317,In_327);
nor U577 (N_577,In_192,In_193);
nand U578 (N_578,In_191,In_675);
nor U579 (N_579,In_724,In_686);
nand U580 (N_580,In_679,In_993);
and U581 (N_581,In_15,In_235);
nor U582 (N_582,In_438,In_248);
and U583 (N_583,In_73,In_981);
and U584 (N_584,In_808,In_378);
and U585 (N_585,In_46,In_940);
or U586 (N_586,In_866,In_454);
and U587 (N_587,In_893,In_536);
or U588 (N_588,In_15,In_685);
nor U589 (N_589,In_870,In_240);
and U590 (N_590,In_507,In_714);
nor U591 (N_591,In_428,In_725);
or U592 (N_592,In_754,In_864);
nand U593 (N_593,In_940,In_132);
or U594 (N_594,In_781,In_860);
and U595 (N_595,In_20,In_667);
nor U596 (N_596,In_626,In_111);
or U597 (N_597,In_279,In_578);
nor U598 (N_598,In_858,In_383);
nor U599 (N_599,In_438,In_3);
nor U600 (N_600,In_602,In_567);
and U601 (N_601,In_197,In_130);
nor U602 (N_602,In_685,In_178);
xnor U603 (N_603,In_503,In_216);
nand U604 (N_604,In_433,In_637);
or U605 (N_605,In_26,In_996);
or U606 (N_606,In_204,In_129);
xnor U607 (N_607,In_227,In_336);
nor U608 (N_608,In_873,In_257);
and U609 (N_609,In_313,In_563);
nand U610 (N_610,In_236,In_924);
or U611 (N_611,In_186,In_447);
nor U612 (N_612,In_238,In_539);
nor U613 (N_613,In_273,In_466);
xnor U614 (N_614,In_179,In_183);
or U615 (N_615,In_16,In_591);
and U616 (N_616,In_840,In_326);
nand U617 (N_617,In_571,In_388);
or U618 (N_618,In_253,In_12);
or U619 (N_619,In_816,In_567);
and U620 (N_620,In_304,In_326);
or U621 (N_621,In_37,In_516);
or U622 (N_622,In_590,In_485);
and U623 (N_623,In_846,In_980);
or U624 (N_624,In_453,In_674);
nor U625 (N_625,In_366,In_807);
nor U626 (N_626,In_923,In_449);
nor U627 (N_627,In_620,In_402);
or U628 (N_628,In_441,In_666);
or U629 (N_629,In_482,In_175);
or U630 (N_630,In_291,In_315);
nor U631 (N_631,In_742,In_424);
nand U632 (N_632,In_899,In_509);
nand U633 (N_633,In_856,In_919);
nor U634 (N_634,In_210,In_726);
or U635 (N_635,In_201,In_987);
or U636 (N_636,In_630,In_839);
xnor U637 (N_637,In_176,In_405);
xor U638 (N_638,In_848,In_525);
nor U639 (N_639,In_228,In_50);
nand U640 (N_640,In_876,In_667);
nand U641 (N_641,In_805,In_789);
and U642 (N_642,In_688,In_316);
or U643 (N_643,In_381,In_122);
and U644 (N_644,In_919,In_370);
and U645 (N_645,In_974,In_429);
and U646 (N_646,In_310,In_644);
nor U647 (N_647,In_661,In_194);
nand U648 (N_648,In_225,In_679);
or U649 (N_649,In_333,In_290);
xnor U650 (N_650,In_641,In_832);
and U651 (N_651,In_898,In_671);
nand U652 (N_652,In_17,In_28);
nand U653 (N_653,In_830,In_685);
nor U654 (N_654,In_649,In_560);
or U655 (N_655,In_567,In_725);
nor U656 (N_656,In_283,In_135);
and U657 (N_657,In_837,In_819);
nor U658 (N_658,In_332,In_194);
nor U659 (N_659,In_365,In_908);
xnor U660 (N_660,In_475,In_78);
nand U661 (N_661,In_9,In_135);
and U662 (N_662,In_485,In_15);
nand U663 (N_663,In_318,In_394);
or U664 (N_664,In_442,In_994);
nor U665 (N_665,In_517,In_624);
xor U666 (N_666,In_188,In_166);
and U667 (N_667,In_912,In_746);
nand U668 (N_668,In_480,In_412);
nor U669 (N_669,In_70,In_536);
and U670 (N_670,In_918,In_867);
or U671 (N_671,In_882,In_462);
xor U672 (N_672,In_699,In_834);
and U673 (N_673,In_772,In_577);
xor U674 (N_674,In_262,In_386);
nand U675 (N_675,In_425,In_205);
xor U676 (N_676,In_994,In_569);
and U677 (N_677,In_203,In_59);
nand U678 (N_678,In_326,In_818);
or U679 (N_679,In_804,In_533);
or U680 (N_680,In_28,In_461);
or U681 (N_681,In_804,In_6);
nor U682 (N_682,In_342,In_728);
nand U683 (N_683,In_701,In_190);
and U684 (N_684,In_95,In_543);
nand U685 (N_685,In_239,In_679);
and U686 (N_686,In_903,In_655);
or U687 (N_687,In_747,In_36);
xor U688 (N_688,In_969,In_786);
and U689 (N_689,In_717,In_902);
nor U690 (N_690,In_21,In_93);
nor U691 (N_691,In_451,In_539);
nand U692 (N_692,In_711,In_869);
nor U693 (N_693,In_225,In_598);
nand U694 (N_694,In_276,In_428);
and U695 (N_695,In_670,In_572);
or U696 (N_696,In_983,In_961);
or U697 (N_697,In_610,In_849);
and U698 (N_698,In_920,In_803);
and U699 (N_699,In_169,In_246);
or U700 (N_700,In_707,In_918);
and U701 (N_701,In_908,In_194);
or U702 (N_702,In_884,In_463);
or U703 (N_703,In_520,In_750);
nand U704 (N_704,In_561,In_768);
or U705 (N_705,In_607,In_975);
nor U706 (N_706,In_79,In_293);
nand U707 (N_707,In_161,In_641);
xor U708 (N_708,In_314,In_350);
and U709 (N_709,In_460,In_929);
nor U710 (N_710,In_297,In_887);
and U711 (N_711,In_875,In_595);
nor U712 (N_712,In_544,In_386);
and U713 (N_713,In_102,In_858);
or U714 (N_714,In_468,In_862);
xnor U715 (N_715,In_490,In_79);
nand U716 (N_716,In_705,In_949);
nand U717 (N_717,In_713,In_569);
or U718 (N_718,In_14,In_588);
nor U719 (N_719,In_540,In_203);
nor U720 (N_720,In_783,In_44);
and U721 (N_721,In_392,In_998);
and U722 (N_722,In_920,In_979);
nand U723 (N_723,In_387,In_706);
nand U724 (N_724,In_970,In_387);
nand U725 (N_725,In_848,In_838);
and U726 (N_726,In_683,In_568);
or U727 (N_727,In_6,In_611);
nand U728 (N_728,In_355,In_13);
and U729 (N_729,In_327,In_188);
nor U730 (N_730,In_621,In_657);
nand U731 (N_731,In_481,In_311);
or U732 (N_732,In_118,In_93);
and U733 (N_733,In_94,In_666);
nand U734 (N_734,In_971,In_628);
or U735 (N_735,In_8,In_598);
or U736 (N_736,In_165,In_940);
xnor U737 (N_737,In_859,In_940);
nor U738 (N_738,In_429,In_38);
nor U739 (N_739,In_67,In_383);
nand U740 (N_740,In_922,In_730);
nand U741 (N_741,In_424,In_930);
nand U742 (N_742,In_262,In_247);
nand U743 (N_743,In_920,In_884);
nor U744 (N_744,In_487,In_987);
nand U745 (N_745,In_333,In_776);
nand U746 (N_746,In_617,In_106);
or U747 (N_747,In_281,In_471);
nor U748 (N_748,In_281,In_326);
nor U749 (N_749,In_231,In_153);
nor U750 (N_750,In_131,In_776);
xor U751 (N_751,In_413,In_794);
nor U752 (N_752,In_397,In_166);
or U753 (N_753,In_305,In_576);
and U754 (N_754,In_565,In_179);
and U755 (N_755,In_71,In_944);
nand U756 (N_756,In_417,In_26);
or U757 (N_757,In_873,In_67);
nand U758 (N_758,In_439,In_281);
and U759 (N_759,In_925,In_985);
and U760 (N_760,In_85,In_169);
nand U761 (N_761,In_546,In_135);
nand U762 (N_762,In_541,In_459);
xor U763 (N_763,In_531,In_813);
or U764 (N_764,In_884,In_356);
and U765 (N_765,In_749,In_725);
nand U766 (N_766,In_225,In_319);
and U767 (N_767,In_767,In_294);
and U768 (N_768,In_493,In_319);
or U769 (N_769,In_609,In_293);
or U770 (N_770,In_492,In_481);
or U771 (N_771,In_789,In_604);
and U772 (N_772,In_991,In_675);
xor U773 (N_773,In_180,In_299);
xnor U774 (N_774,In_179,In_106);
nand U775 (N_775,In_639,In_409);
xnor U776 (N_776,In_536,In_164);
xnor U777 (N_777,In_458,In_592);
nor U778 (N_778,In_237,In_50);
or U779 (N_779,In_634,In_730);
and U780 (N_780,In_560,In_181);
nand U781 (N_781,In_515,In_426);
nand U782 (N_782,In_524,In_669);
nand U783 (N_783,In_490,In_623);
and U784 (N_784,In_818,In_136);
xor U785 (N_785,In_63,In_615);
or U786 (N_786,In_922,In_657);
or U787 (N_787,In_844,In_586);
or U788 (N_788,In_15,In_86);
nand U789 (N_789,In_702,In_365);
and U790 (N_790,In_173,In_748);
nand U791 (N_791,In_616,In_935);
or U792 (N_792,In_735,In_553);
or U793 (N_793,In_657,In_233);
and U794 (N_794,In_170,In_84);
xnor U795 (N_795,In_846,In_785);
and U796 (N_796,In_513,In_343);
nor U797 (N_797,In_778,In_907);
nor U798 (N_798,In_542,In_112);
nor U799 (N_799,In_767,In_306);
nand U800 (N_800,In_938,In_561);
and U801 (N_801,In_277,In_754);
or U802 (N_802,In_230,In_70);
and U803 (N_803,In_46,In_478);
nand U804 (N_804,In_971,In_123);
nor U805 (N_805,In_970,In_719);
nand U806 (N_806,In_714,In_473);
and U807 (N_807,In_869,In_335);
xor U808 (N_808,In_370,In_572);
or U809 (N_809,In_251,In_914);
nand U810 (N_810,In_257,In_501);
xnor U811 (N_811,In_425,In_490);
nor U812 (N_812,In_28,In_550);
nand U813 (N_813,In_232,In_785);
and U814 (N_814,In_862,In_725);
and U815 (N_815,In_869,In_410);
or U816 (N_816,In_697,In_969);
xnor U817 (N_817,In_617,In_639);
or U818 (N_818,In_38,In_846);
or U819 (N_819,In_111,In_728);
and U820 (N_820,In_590,In_900);
and U821 (N_821,In_471,In_880);
nand U822 (N_822,In_943,In_778);
and U823 (N_823,In_606,In_386);
nor U824 (N_824,In_365,In_735);
and U825 (N_825,In_54,In_783);
and U826 (N_826,In_442,In_372);
nand U827 (N_827,In_681,In_210);
and U828 (N_828,In_241,In_591);
nor U829 (N_829,In_816,In_428);
xor U830 (N_830,In_291,In_805);
and U831 (N_831,In_46,In_341);
and U832 (N_832,In_236,In_757);
or U833 (N_833,In_895,In_75);
and U834 (N_834,In_528,In_733);
or U835 (N_835,In_285,In_496);
nor U836 (N_836,In_855,In_206);
xnor U837 (N_837,In_962,In_127);
nor U838 (N_838,In_287,In_27);
or U839 (N_839,In_220,In_451);
nand U840 (N_840,In_50,In_235);
nand U841 (N_841,In_198,In_975);
nand U842 (N_842,In_724,In_975);
or U843 (N_843,In_903,In_20);
nand U844 (N_844,In_586,In_46);
nand U845 (N_845,In_643,In_135);
or U846 (N_846,In_739,In_968);
nor U847 (N_847,In_766,In_35);
nand U848 (N_848,In_894,In_113);
nand U849 (N_849,In_304,In_707);
or U850 (N_850,In_989,In_284);
nor U851 (N_851,In_952,In_134);
xnor U852 (N_852,In_873,In_692);
nor U853 (N_853,In_450,In_312);
or U854 (N_854,In_904,In_662);
xnor U855 (N_855,In_490,In_792);
and U856 (N_856,In_876,In_373);
and U857 (N_857,In_635,In_559);
or U858 (N_858,In_945,In_946);
nor U859 (N_859,In_126,In_244);
and U860 (N_860,In_879,In_105);
xor U861 (N_861,In_364,In_138);
nor U862 (N_862,In_900,In_568);
xnor U863 (N_863,In_582,In_699);
nor U864 (N_864,In_324,In_163);
nand U865 (N_865,In_965,In_748);
or U866 (N_866,In_408,In_119);
and U867 (N_867,In_671,In_956);
xor U868 (N_868,In_430,In_507);
nor U869 (N_869,In_308,In_693);
and U870 (N_870,In_220,In_512);
xor U871 (N_871,In_801,In_166);
nor U872 (N_872,In_719,In_433);
nor U873 (N_873,In_337,In_22);
nor U874 (N_874,In_755,In_636);
nand U875 (N_875,In_809,In_356);
nor U876 (N_876,In_616,In_859);
or U877 (N_877,In_847,In_349);
nand U878 (N_878,In_471,In_567);
nand U879 (N_879,In_112,In_589);
nor U880 (N_880,In_596,In_862);
xor U881 (N_881,In_900,In_380);
or U882 (N_882,In_262,In_949);
nor U883 (N_883,In_284,In_759);
xnor U884 (N_884,In_374,In_619);
nor U885 (N_885,In_758,In_936);
xnor U886 (N_886,In_858,In_839);
nand U887 (N_887,In_565,In_818);
or U888 (N_888,In_80,In_842);
nand U889 (N_889,In_531,In_327);
or U890 (N_890,In_683,In_370);
or U891 (N_891,In_928,In_428);
nand U892 (N_892,In_799,In_674);
and U893 (N_893,In_200,In_639);
nand U894 (N_894,In_101,In_928);
nor U895 (N_895,In_117,In_142);
nand U896 (N_896,In_114,In_307);
nand U897 (N_897,In_887,In_137);
or U898 (N_898,In_811,In_966);
or U899 (N_899,In_528,In_511);
nand U900 (N_900,In_858,In_431);
and U901 (N_901,In_491,In_970);
and U902 (N_902,In_813,In_368);
nand U903 (N_903,In_837,In_780);
nor U904 (N_904,In_995,In_142);
nor U905 (N_905,In_461,In_74);
and U906 (N_906,In_938,In_590);
nor U907 (N_907,In_891,In_849);
nor U908 (N_908,In_475,In_539);
and U909 (N_909,In_985,In_459);
nor U910 (N_910,In_928,In_722);
nand U911 (N_911,In_386,In_772);
nor U912 (N_912,In_988,In_745);
nor U913 (N_913,In_773,In_776);
nand U914 (N_914,In_282,In_573);
xor U915 (N_915,In_814,In_249);
or U916 (N_916,In_110,In_270);
nand U917 (N_917,In_939,In_654);
or U918 (N_918,In_437,In_600);
nand U919 (N_919,In_136,In_444);
nor U920 (N_920,In_244,In_758);
nand U921 (N_921,In_118,In_634);
nand U922 (N_922,In_514,In_77);
nor U923 (N_923,In_790,In_705);
and U924 (N_924,In_305,In_331);
nor U925 (N_925,In_902,In_764);
and U926 (N_926,In_596,In_247);
nand U927 (N_927,In_848,In_324);
nand U928 (N_928,In_378,In_571);
or U929 (N_929,In_314,In_396);
or U930 (N_930,In_343,In_184);
nor U931 (N_931,In_770,In_85);
nand U932 (N_932,In_698,In_154);
or U933 (N_933,In_261,In_397);
xnor U934 (N_934,In_380,In_912);
and U935 (N_935,In_185,In_995);
nor U936 (N_936,In_453,In_297);
nand U937 (N_937,In_280,In_536);
nand U938 (N_938,In_709,In_983);
nor U939 (N_939,In_438,In_959);
xnor U940 (N_940,In_973,In_449);
nand U941 (N_941,In_990,In_524);
or U942 (N_942,In_535,In_893);
and U943 (N_943,In_67,In_349);
and U944 (N_944,In_406,In_284);
and U945 (N_945,In_578,In_482);
nand U946 (N_946,In_143,In_847);
nor U947 (N_947,In_764,In_758);
xor U948 (N_948,In_581,In_816);
nand U949 (N_949,In_50,In_386);
or U950 (N_950,In_354,In_92);
or U951 (N_951,In_221,In_730);
nand U952 (N_952,In_413,In_110);
and U953 (N_953,In_631,In_196);
nor U954 (N_954,In_283,In_400);
and U955 (N_955,In_745,In_457);
xnor U956 (N_956,In_361,In_583);
or U957 (N_957,In_361,In_907);
and U958 (N_958,In_825,In_147);
nor U959 (N_959,In_575,In_262);
nand U960 (N_960,In_463,In_134);
nor U961 (N_961,In_177,In_946);
nor U962 (N_962,In_136,In_272);
and U963 (N_963,In_977,In_720);
and U964 (N_964,In_186,In_645);
nand U965 (N_965,In_510,In_870);
or U966 (N_966,In_319,In_534);
or U967 (N_967,In_724,In_329);
xnor U968 (N_968,In_986,In_334);
or U969 (N_969,In_261,In_316);
nand U970 (N_970,In_973,In_311);
or U971 (N_971,In_429,In_118);
and U972 (N_972,In_38,In_162);
nand U973 (N_973,In_169,In_253);
or U974 (N_974,In_925,In_462);
nand U975 (N_975,In_652,In_745);
nor U976 (N_976,In_728,In_884);
or U977 (N_977,In_582,In_901);
xnor U978 (N_978,In_250,In_148);
or U979 (N_979,In_158,In_966);
and U980 (N_980,In_343,In_585);
nor U981 (N_981,In_592,In_702);
nor U982 (N_982,In_215,In_572);
and U983 (N_983,In_585,In_471);
and U984 (N_984,In_121,In_377);
or U985 (N_985,In_641,In_846);
nor U986 (N_986,In_329,In_299);
and U987 (N_987,In_516,In_664);
and U988 (N_988,In_433,In_904);
or U989 (N_989,In_427,In_757);
nand U990 (N_990,In_184,In_416);
or U991 (N_991,In_162,In_714);
or U992 (N_992,In_190,In_374);
or U993 (N_993,In_611,In_877);
nand U994 (N_994,In_847,In_47);
and U995 (N_995,In_80,In_433);
and U996 (N_996,In_478,In_311);
and U997 (N_997,In_579,In_350);
or U998 (N_998,In_39,In_498);
nor U999 (N_999,In_98,In_561);
xor U1000 (N_1000,In_890,In_212);
nand U1001 (N_1001,In_613,In_572);
and U1002 (N_1002,In_602,In_316);
or U1003 (N_1003,In_144,In_443);
xnor U1004 (N_1004,In_235,In_510);
nor U1005 (N_1005,In_613,In_883);
nor U1006 (N_1006,In_11,In_803);
and U1007 (N_1007,In_86,In_981);
nand U1008 (N_1008,In_467,In_733);
and U1009 (N_1009,In_338,In_169);
and U1010 (N_1010,In_234,In_83);
and U1011 (N_1011,In_686,In_275);
or U1012 (N_1012,In_501,In_31);
and U1013 (N_1013,In_790,In_963);
nor U1014 (N_1014,In_707,In_486);
and U1015 (N_1015,In_635,In_236);
and U1016 (N_1016,In_714,In_589);
nor U1017 (N_1017,In_391,In_248);
and U1018 (N_1018,In_377,In_274);
nand U1019 (N_1019,In_710,In_402);
or U1020 (N_1020,In_794,In_266);
nand U1021 (N_1021,In_474,In_52);
and U1022 (N_1022,In_436,In_675);
nand U1023 (N_1023,In_495,In_525);
or U1024 (N_1024,In_871,In_309);
nor U1025 (N_1025,In_717,In_323);
or U1026 (N_1026,In_931,In_819);
nor U1027 (N_1027,In_437,In_534);
xor U1028 (N_1028,In_537,In_405);
nand U1029 (N_1029,In_345,In_456);
or U1030 (N_1030,In_234,In_367);
nand U1031 (N_1031,In_922,In_679);
or U1032 (N_1032,In_970,In_546);
nand U1033 (N_1033,In_68,In_448);
nand U1034 (N_1034,In_714,In_99);
nand U1035 (N_1035,In_569,In_715);
or U1036 (N_1036,In_202,In_526);
nor U1037 (N_1037,In_290,In_266);
nand U1038 (N_1038,In_155,In_324);
nor U1039 (N_1039,In_717,In_781);
or U1040 (N_1040,In_589,In_857);
nor U1041 (N_1041,In_184,In_104);
nand U1042 (N_1042,In_211,In_985);
nand U1043 (N_1043,In_56,In_514);
nor U1044 (N_1044,In_277,In_972);
xnor U1045 (N_1045,In_47,In_38);
nand U1046 (N_1046,In_250,In_760);
or U1047 (N_1047,In_852,In_783);
and U1048 (N_1048,In_545,In_859);
nor U1049 (N_1049,In_482,In_5);
nor U1050 (N_1050,In_304,In_919);
or U1051 (N_1051,In_242,In_120);
or U1052 (N_1052,In_248,In_457);
nor U1053 (N_1053,In_432,In_776);
nand U1054 (N_1054,In_906,In_34);
and U1055 (N_1055,In_244,In_220);
and U1056 (N_1056,In_626,In_899);
nor U1057 (N_1057,In_826,In_503);
nor U1058 (N_1058,In_318,In_423);
nand U1059 (N_1059,In_874,In_443);
and U1060 (N_1060,In_729,In_568);
nor U1061 (N_1061,In_401,In_722);
nand U1062 (N_1062,In_708,In_881);
or U1063 (N_1063,In_805,In_714);
or U1064 (N_1064,In_7,In_717);
nand U1065 (N_1065,In_697,In_243);
or U1066 (N_1066,In_917,In_972);
and U1067 (N_1067,In_790,In_897);
and U1068 (N_1068,In_874,In_177);
nor U1069 (N_1069,In_892,In_546);
nor U1070 (N_1070,In_789,In_943);
or U1071 (N_1071,In_950,In_925);
xnor U1072 (N_1072,In_534,In_757);
or U1073 (N_1073,In_264,In_163);
or U1074 (N_1074,In_938,In_860);
nor U1075 (N_1075,In_488,In_27);
nand U1076 (N_1076,In_846,In_136);
nand U1077 (N_1077,In_679,In_694);
nand U1078 (N_1078,In_814,In_698);
nand U1079 (N_1079,In_746,In_278);
nor U1080 (N_1080,In_375,In_434);
nor U1081 (N_1081,In_274,In_943);
nor U1082 (N_1082,In_29,In_633);
and U1083 (N_1083,In_906,In_915);
nand U1084 (N_1084,In_816,In_235);
nand U1085 (N_1085,In_989,In_861);
and U1086 (N_1086,In_106,In_631);
xnor U1087 (N_1087,In_375,In_923);
or U1088 (N_1088,In_12,In_829);
nor U1089 (N_1089,In_933,In_798);
xor U1090 (N_1090,In_140,In_570);
and U1091 (N_1091,In_179,In_736);
and U1092 (N_1092,In_203,In_299);
or U1093 (N_1093,In_772,In_402);
and U1094 (N_1094,In_344,In_438);
nor U1095 (N_1095,In_501,In_994);
nor U1096 (N_1096,In_143,In_181);
and U1097 (N_1097,In_960,In_429);
xnor U1098 (N_1098,In_310,In_266);
nand U1099 (N_1099,In_824,In_166);
nand U1100 (N_1100,In_204,In_11);
nor U1101 (N_1101,In_45,In_867);
xnor U1102 (N_1102,In_939,In_413);
xnor U1103 (N_1103,In_194,In_168);
nand U1104 (N_1104,In_790,In_462);
and U1105 (N_1105,In_817,In_231);
nand U1106 (N_1106,In_774,In_43);
and U1107 (N_1107,In_428,In_828);
nand U1108 (N_1108,In_495,In_479);
xor U1109 (N_1109,In_502,In_65);
or U1110 (N_1110,In_751,In_121);
and U1111 (N_1111,In_729,In_654);
and U1112 (N_1112,In_541,In_440);
nor U1113 (N_1113,In_111,In_447);
or U1114 (N_1114,In_588,In_424);
nor U1115 (N_1115,In_811,In_261);
or U1116 (N_1116,In_524,In_357);
nand U1117 (N_1117,In_926,In_487);
nor U1118 (N_1118,In_532,In_95);
and U1119 (N_1119,In_454,In_20);
or U1120 (N_1120,In_308,In_424);
or U1121 (N_1121,In_107,In_934);
or U1122 (N_1122,In_65,In_444);
nor U1123 (N_1123,In_224,In_26);
nand U1124 (N_1124,In_212,In_762);
xnor U1125 (N_1125,In_776,In_860);
and U1126 (N_1126,In_152,In_109);
or U1127 (N_1127,In_711,In_53);
or U1128 (N_1128,In_876,In_469);
nand U1129 (N_1129,In_906,In_495);
or U1130 (N_1130,In_392,In_458);
nand U1131 (N_1131,In_472,In_317);
nor U1132 (N_1132,In_255,In_771);
or U1133 (N_1133,In_507,In_756);
and U1134 (N_1134,In_413,In_707);
and U1135 (N_1135,In_146,In_235);
nor U1136 (N_1136,In_766,In_973);
or U1137 (N_1137,In_171,In_680);
nand U1138 (N_1138,In_513,In_294);
nand U1139 (N_1139,In_459,In_573);
or U1140 (N_1140,In_134,In_55);
nand U1141 (N_1141,In_455,In_155);
nand U1142 (N_1142,In_526,In_314);
xor U1143 (N_1143,In_664,In_638);
or U1144 (N_1144,In_485,In_913);
and U1145 (N_1145,In_654,In_870);
nand U1146 (N_1146,In_924,In_111);
and U1147 (N_1147,In_28,In_671);
xnor U1148 (N_1148,In_670,In_201);
nand U1149 (N_1149,In_499,In_191);
and U1150 (N_1150,In_820,In_717);
nand U1151 (N_1151,In_609,In_229);
xor U1152 (N_1152,In_556,In_736);
or U1153 (N_1153,In_801,In_248);
and U1154 (N_1154,In_581,In_780);
nand U1155 (N_1155,In_114,In_646);
or U1156 (N_1156,In_955,In_26);
or U1157 (N_1157,In_907,In_150);
nand U1158 (N_1158,In_374,In_801);
or U1159 (N_1159,In_771,In_198);
or U1160 (N_1160,In_576,In_813);
or U1161 (N_1161,In_476,In_639);
nor U1162 (N_1162,In_405,In_528);
nand U1163 (N_1163,In_24,In_246);
and U1164 (N_1164,In_402,In_586);
nor U1165 (N_1165,In_714,In_695);
nand U1166 (N_1166,In_971,In_651);
and U1167 (N_1167,In_195,In_973);
or U1168 (N_1168,In_154,In_772);
or U1169 (N_1169,In_588,In_151);
nor U1170 (N_1170,In_179,In_792);
nor U1171 (N_1171,In_934,In_386);
nor U1172 (N_1172,In_270,In_923);
nor U1173 (N_1173,In_754,In_375);
and U1174 (N_1174,In_926,In_895);
nor U1175 (N_1175,In_664,In_74);
and U1176 (N_1176,In_555,In_168);
xor U1177 (N_1177,In_890,In_374);
or U1178 (N_1178,In_316,In_785);
and U1179 (N_1179,In_927,In_188);
nand U1180 (N_1180,In_889,In_677);
nor U1181 (N_1181,In_958,In_356);
and U1182 (N_1182,In_655,In_3);
or U1183 (N_1183,In_497,In_673);
nand U1184 (N_1184,In_465,In_892);
xnor U1185 (N_1185,In_725,In_878);
xor U1186 (N_1186,In_801,In_448);
nor U1187 (N_1187,In_356,In_667);
xor U1188 (N_1188,In_488,In_484);
or U1189 (N_1189,In_27,In_831);
nand U1190 (N_1190,In_268,In_667);
nand U1191 (N_1191,In_441,In_395);
nor U1192 (N_1192,In_608,In_739);
nand U1193 (N_1193,In_663,In_449);
or U1194 (N_1194,In_765,In_724);
nand U1195 (N_1195,In_946,In_556);
xor U1196 (N_1196,In_592,In_924);
nor U1197 (N_1197,In_776,In_822);
nand U1198 (N_1198,In_723,In_613);
or U1199 (N_1199,In_278,In_274);
nand U1200 (N_1200,In_719,In_111);
nand U1201 (N_1201,In_481,In_987);
or U1202 (N_1202,In_178,In_404);
and U1203 (N_1203,In_388,In_10);
and U1204 (N_1204,In_460,In_864);
and U1205 (N_1205,In_72,In_967);
or U1206 (N_1206,In_359,In_724);
xnor U1207 (N_1207,In_218,In_784);
nor U1208 (N_1208,In_147,In_773);
and U1209 (N_1209,In_89,In_805);
nand U1210 (N_1210,In_507,In_269);
or U1211 (N_1211,In_377,In_707);
nand U1212 (N_1212,In_343,In_830);
nor U1213 (N_1213,In_742,In_933);
or U1214 (N_1214,In_870,In_523);
nand U1215 (N_1215,In_676,In_807);
or U1216 (N_1216,In_995,In_710);
xor U1217 (N_1217,In_912,In_904);
nand U1218 (N_1218,In_600,In_381);
or U1219 (N_1219,In_424,In_28);
and U1220 (N_1220,In_921,In_697);
nor U1221 (N_1221,In_795,In_280);
or U1222 (N_1222,In_297,In_218);
and U1223 (N_1223,In_870,In_506);
nand U1224 (N_1224,In_79,In_333);
and U1225 (N_1225,In_958,In_828);
nand U1226 (N_1226,In_625,In_173);
xor U1227 (N_1227,In_799,In_903);
xnor U1228 (N_1228,In_490,In_413);
or U1229 (N_1229,In_243,In_360);
and U1230 (N_1230,In_617,In_658);
or U1231 (N_1231,In_716,In_278);
nand U1232 (N_1232,In_833,In_677);
nor U1233 (N_1233,In_283,In_615);
nand U1234 (N_1234,In_194,In_796);
xnor U1235 (N_1235,In_906,In_639);
nand U1236 (N_1236,In_43,In_1);
or U1237 (N_1237,In_182,In_771);
xnor U1238 (N_1238,In_548,In_831);
or U1239 (N_1239,In_808,In_717);
or U1240 (N_1240,In_575,In_226);
and U1241 (N_1241,In_496,In_404);
nor U1242 (N_1242,In_169,In_438);
nor U1243 (N_1243,In_37,In_450);
nand U1244 (N_1244,In_463,In_278);
nor U1245 (N_1245,In_364,In_933);
and U1246 (N_1246,In_375,In_595);
or U1247 (N_1247,In_325,In_233);
or U1248 (N_1248,In_779,In_721);
nand U1249 (N_1249,In_600,In_720);
nor U1250 (N_1250,In_33,In_701);
nor U1251 (N_1251,In_162,In_734);
nand U1252 (N_1252,In_549,In_162);
xnor U1253 (N_1253,In_965,In_302);
nor U1254 (N_1254,In_342,In_686);
nand U1255 (N_1255,In_492,In_273);
nand U1256 (N_1256,In_316,In_12);
and U1257 (N_1257,In_201,In_787);
and U1258 (N_1258,In_51,In_300);
and U1259 (N_1259,In_898,In_549);
xnor U1260 (N_1260,In_903,In_451);
nand U1261 (N_1261,In_751,In_479);
nor U1262 (N_1262,In_913,In_2);
nand U1263 (N_1263,In_962,In_550);
nor U1264 (N_1264,In_151,In_465);
nor U1265 (N_1265,In_779,In_725);
nand U1266 (N_1266,In_435,In_564);
and U1267 (N_1267,In_210,In_553);
and U1268 (N_1268,In_882,In_568);
or U1269 (N_1269,In_972,In_172);
and U1270 (N_1270,In_685,In_934);
or U1271 (N_1271,In_986,In_528);
nand U1272 (N_1272,In_477,In_462);
nand U1273 (N_1273,In_502,In_58);
nor U1274 (N_1274,In_218,In_627);
nand U1275 (N_1275,In_895,In_580);
and U1276 (N_1276,In_992,In_118);
or U1277 (N_1277,In_240,In_173);
nand U1278 (N_1278,In_59,In_750);
xor U1279 (N_1279,In_209,In_646);
nand U1280 (N_1280,In_349,In_734);
and U1281 (N_1281,In_44,In_297);
nor U1282 (N_1282,In_329,In_518);
and U1283 (N_1283,In_380,In_714);
and U1284 (N_1284,In_663,In_852);
nor U1285 (N_1285,In_131,In_137);
and U1286 (N_1286,In_647,In_439);
nand U1287 (N_1287,In_14,In_514);
nor U1288 (N_1288,In_528,In_625);
xor U1289 (N_1289,In_226,In_970);
nand U1290 (N_1290,In_943,In_319);
and U1291 (N_1291,In_874,In_168);
nand U1292 (N_1292,In_524,In_878);
nand U1293 (N_1293,In_486,In_852);
and U1294 (N_1294,In_909,In_940);
and U1295 (N_1295,In_839,In_152);
and U1296 (N_1296,In_338,In_678);
nor U1297 (N_1297,In_24,In_677);
or U1298 (N_1298,In_737,In_281);
or U1299 (N_1299,In_669,In_924);
nand U1300 (N_1300,In_264,In_848);
and U1301 (N_1301,In_87,In_369);
nand U1302 (N_1302,In_273,In_420);
and U1303 (N_1303,In_703,In_723);
and U1304 (N_1304,In_121,In_235);
nor U1305 (N_1305,In_280,In_125);
or U1306 (N_1306,In_307,In_667);
or U1307 (N_1307,In_387,In_587);
or U1308 (N_1308,In_341,In_775);
nand U1309 (N_1309,In_985,In_147);
xnor U1310 (N_1310,In_743,In_993);
nor U1311 (N_1311,In_168,In_289);
xnor U1312 (N_1312,In_67,In_874);
nor U1313 (N_1313,In_820,In_923);
nand U1314 (N_1314,In_711,In_931);
or U1315 (N_1315,In_794,In_553);
xnor U1316 (N_1316,In_38,In_525);
and U1317 (N_1317,In_528,In_836);
and U1318 (N_1318,In_14,In_93);
nand U1319 (N_1319,In_478,In_262);
nand U1320 (N_1320,In_95,In_991);
and U1321 (N_1321,In_489,In_23);
or U1322 (N_1322,In_725,In_961);
or U1323 (N_1323,In_281,In_657);
xnor U1324 (N_1324,In_772,In_72);
and U1325 (N_1325,In_416,In_450);
or U1326 (N_1326,In_988,In_384);
or U1327 (N_1327,In_143,In_934);
nor U1328 (N_1328,In_343,In_176);
or U1329 (N_1329,In_124,In_204);
nand U1330 (N_1330,In_136,In_684);
xnor U1331 (N_1331,In_125,In_88);
nor U1332 (N_1332,In_211,In_171);
and U1333 (N_1333,In_317,In_554);
nor U1334 (N_1334,In_83,In_419);
or U1335 (N_1335,In_810,In_899);
nand U1336 (N_1336,In_493,In_217);
nand U1337 (N_1337,In_950,In_817);
or U1338 (N_1338,In_389,In_235);
nor U1339 (N_1339,In_854,In_541);
and U1340 (N_1340,In_312,In_532);
or U1341 (N_1341,In_295,In_646);
nor U1342 (N_1342,In_439,In_525);
nor U1343 (N_1343,In_542,In_986);
and U1344 (N_1344,In_757,In_129);
or U1345 (N_1345,In_247,In_794);
nor U1346 (N_1346,In_838,In_468);
and U1347 (N_1347,In_432,In_551);
or U1348 (N_1348,In_842,In_327);
nor U1349 (N_1349,In_812,In_420);
or U1350 (N_1350,In_786,In_943);
nor U1351 (N_1351,In_373,In_980);
and U1352 (N_1352,In_675,In_771);
and U1353 (N_1353,In_297,In_515);
and U1354 (N_1354,In_40,In_814);
or U1355 (N_1355,In_969,In_731);
or U1356 (N_1356,In_322,In_540);
or U1357 (N_1357,In_609,In_61);
or U1358 (N_1358,In_320,In_896);
xor U1359 (N_1359,In_818,In_115);
nor U1360 (N_1360,In_914,In_562);
and U1361 (N_1361,In_281,In_48);
and U1362 (N_1362,In_622,In_10);
nor U1363 (N_1363,In_778,In_367);
or U1364 (N_1364,In_812,In_117);
xnor U1365 (N_1365,In_252,In_917);
or U1366 (N_1366,In_661,In_860);
or U1367 (N_1367,In_297,In_552);
and U1368 (N_1368,In_550,In_538);
nand U1369 (N_1369,In_766,In_754);
nor U1370 (N_1370,In_379,In_402);
nand U1371 (N_1371,In_502,In_515);
nor U1372 (N_1372,In_843,In_442);
nor U1373 (N_1373,In_395,In_503);
and U1374 (N_1374,In_19,In_672);
or U1375 (N_1375,In_889,In_654);
and U1376 (N_1376,In_252,In_955);
xnor U1377 (N_1377,In_876,In_628);
and U1378 (N_1378,In_387,In_559);
nand U1379 (N_1379,In_666,In_150);
nand U1380 (N_1380,In_964,In_446);
nor U1381 (N_1381,In_786,In_474);
nand U1382 (N_1382,In_437,In_619);
and U1383 (N_1383,In_379,In_571);
and U1384 (N_1384,In_221,In_233);
and U1385 (N_1385,In_746,In_265);
nor U1386 (N_1386,In_751,In_456);
nand U1387 (N_1387,In_847,In_494);
nand U1388 (N_1388,In_790,In_854);
nand U1389 (N_1389,In_878,In_944);
nand U1390 (N_1390,In_703,In_358);
nor U1391 (N_1391,In_847,In_888);
nand U1392 (N_1392,In_604,In_602);
nor U1393 (N_1393,In_421,In_238);
or U1394 (N_1394,In_273,In_145);
or U1395 (N_1395,In_78,In_83);
and U1396 (N_1396,In_936,In_486);
nand U1397 (N_1397,In_11,In_860);
and U1398 (N_1398,In_864,In_8);
nand U1399 (N_1399,In_17,In_434);
or U1400 (N_1400,In_314,In_905);
and U1401 (N_1401,In_141,In_537);
and U1402 (N_1402,In_862,In_247);
nand U1403 (N_1403,In_394,In_431);
nand U1404 (N_1404,In_548,In_280);
xnor U1405 (N_1405,In_812,In_972);
or U1406 (N_1406,In_643,In_359);
nand U1407 (N_1407,In_993,In_215);
nand U1408 (N_1408,In_2,In_942);
nor U1409 (N_1409,In_264,In_469);
or U1410 (N_1410,In_20,In_978);
nand U1411 (N_1411,In_768,In_111);
nand U1412 (N_1412,In_37,In_69);
or U1413 (N_1413,In_294,In_742);
nand U1414 (N_1414,In_950,In_396);
nand U1415 (N_1415,In_950,In_836);
nor U1416 (N_1416,In_678,In_48);
xor U1417 (N_1417,In_376,In_175);
nor U1418 (N_1418,In_917,In_885);
nand U1419 (N_1419,In_680,In_421);
xnor U1420 (N_1420,In_417,In_499);
xor U1421 (N_1421,In_366,In_330);
nand U1422 (N_1422,In_232,In_932);
and U1423 (N_1423,In_506,In_968);
nor U1424 (N_1424,In_798,In_496);
or U1425 (N_1425,In_830,In_598);
xor U1426 (N_1426,In_161,In_292);
nand U1427 (N_1427,In_334,In_474);
nor U1428 (N_1428,In_937,In_589);
nand U1429 (N_1429,In_775,In_435);
or U1430 (N_1430,In_650,In_387);
or U1431 (N_1431,In_616,In_359);
or U1432 (N_1432,In_832,In_566);
or U1433 (N_1433,In_73,In_612);
nand U1434 (N_1434,In_225,In_867);
nor U1435 (N_1435,In_825,In_287);
or U1436 (N_1436,In_745,In_578);
and U1437 (N_1437,In_774,In_674);
nand U1438 (N_1438,In_558,In_687);
nor U1439 (N_1439,In_832,In_185);
nand U1440 (N_1440,In_41,In_450);
and U1441 (N_1441,In_406,In_586);
nand U1442 (N_1442,In_911,In_214);
and U1443 (N_1443,In_91,In_580);
nand U1444 (N_1444,In_960,In_497);
and U1445 (N_1445,In_850,In_174);
nand U1446 (N_1446,In_444,In_929);
xor U1447 (N_1447,In_402,In_372);
xor U1448 (N_1448,In_710,In_464);
xor U1449 (N_1449,In_510,In_356);
nor U1450 (N_1450,In_244,In_732);
or U1451 (N_1451,In_993,In_23);
and U1452 (N_1452,In_805,In_205);
and U1453 (N_1453,In_866,In_541);
and U1454 (N_1454,In_78,In_508);
xor U1455 (N_1455,In_577,In_464);
and U1456 (N_1456,In_950,In_208);
and U1457 (N_1457,In_644,In_757);
and U1458 (N_1458,In_235,In_588);
xnor U1459 (N_1459,In_188,In_391);
nand U1460 (N_1460,In_1,In_339);
nand U1461 (N_1461,In_654,In_519);
and U1462 (N_1462,In_122,In_626);
xor U1463 (N_1463,In_773,In_768);
xnor U1464 (N_1464,In_915,In_184);
or U1465 (N_1465,In_703,In_759);
nor U1466 (N_1466,In_519,In_665);
nand U1467 (N_1467,In_809,In_628);
nand U1468 (N_1468,In_551,In_733);
or U1469 (N_1469,In_258,In_594);
and U1470 (N_1470,In_808,In_78);
and U1471 (N_1471,In_935,In_467);
and U1472 (N_1472,In_309,In_304);
and U1473 (N_1473,In_42,In_106);
nand U1474 (N_1474,In_9,In_938);
and U1475 (N_1475,In_443,In_360);
nand U1476 (N_1476,In_153,In_444);
nor U1477 (N_1477,In_166,In_929);
and U1478 (N_1478,In_196,In_233);
nor U1479 (N_1479,In_421,In_310);
nor U1480 (N_1480,In_601,In_664);
nand U1481 (N_1481,In_554,In_413);
nor U1482 (N_1482,In_595,In_390);
and U1483 (N_1483,In_827,In_606);
and U1484 (N_1484,In_753,In_710);
nand U1485 (N_1485,In_58,In_302);
nor U1486 (N_1486,In_531,In_691);
nor U1487 (N_1487,In_789,In_937);
nor U1488 (N_1488,In_294,In_551);
nand U1489 (N_1489,In_11,In_897);
nor U1490 (N_1490,In_433,In_61);
nor U1491 (N_1491,In_369,In_429);
and U1492 (N_1492,In_123,In_215);
nor U1493 (N_1493,In_833,In_346);
and U1494 (N_1494,In_740,In_271);
and U1495 (N_1495,In_479,In_198);
xor U1496 (N_1496,In_916,In_257);
and U1497 (N_1497,In_924,In_211);
nand U1498 (N_1498,In_610,In_158);
nor U1499 (N_1499,In_211,In_428);
or U1500 (N_1500,In_964,In_304);
and U1501 (N_1501,In_322,In_328);
or U1502 (N_1502,In_295,In_266);
and U1503 (N_1503,In_973,In_700);
nand U1504 (N_1504,In_38,In_145);
and U1505 (N_1505,In_984,In_277);
nor U1506 (N_1506,In_503,In_814);
or U1507 (N_1507,In_896,In_168);
or U1508 (N_1508,In_277,In_854);
and U1509 (N_1509,In_862,In_546);
xor U1510 (N_1510,In_540,In_664);
and U1511 (N_1511,In_329,In_984);
nor U1512 (N_1512,In_274,In_646);
and U1513 (N_1513,In_325,In_110);
nand U1514 (N_1514,In_758,In_131);
nor U1515 (N_1515,In_35,In_505);
nor U1516 (N_1516,In_397,In_363);
nor U1517 (N_1517,In_297,In_235);
or U1518 (N_1518,In_877,In_313);
and U1519 (N_1519,In_415,In_967);
or U1520 (N_1520,In_847,In_993);
nand U1521 (N_1521,In_991,In_179);
nand U1522 (N_1522,In_662,In_532);
xnor U1523 (N_1523,In_650,In_599);
nand U1524 (N_1524,In_735,In_701);
and U1525 (N_1525,In_72,In_690);
nand U1526 (N_1526,In_225,In_460);
nand U1527 (N_1527,In_657,In_828);
nor U1528 (N_1528,In_257,In_198);
nor U1529 (N_1529,In_844,In_352);
or U1530 (N_1530,In_131,In_129);
nor U1531 (N_1531,In_940,In_638);
nand U1532 (N_1532,In_456,In_135);
xor U1533 (N_1533,In_2,In_126);
nand U1534 (N_1534,In_556,In_5);
or U1535 (N_1535,In_130,In_443);
or U1536 (N_1536,In_655,In_0);
or U1537 (N_1537,In_474,In_856);
or U1538 (N_1538,In_925,In_158);
nand U1539 (N_1539,In_76,In_103);
nor U1540 (N_1540,In_166,In_736);
nand U1541 (N_1541,In_846,In_429);
nor U1542 (N_1542,In_7,In_206);
nor U1543 (N_1543,In_193,In_460);
nor U1544 (N_1544,In_762,In_721);
nand U1545 (N_1545,In_272,In_96);
nand U1546 (N_1546,In_919,In_797);
or U1547 (N_1547,In_105,In_620);
or U1548 (N_1548,In_20,In_532);
nor U1549 (N_1549,In_446,In_549);
or U1550 (N_1550,In_964,In_56);
nand U1551 (N_1551,In_722,In_187);
or U1552 (N_1552,In_193,In_544);
nand U1553 (N_1553,In_37,In_981);
and U1554 (N_1554,In_832,In_349);
and U1555 (N_1555,In_491,In_621);
nand U1556 (N_1556,In_877,In_831);
nor U1557 (N_1557,In_2,In_750);
and U1558 (N_1558,In_230,In_67);
or U1559 (N_1559,In_535,In_918);
xnor U1560 (N_1560,In_199,In_521);
xnor U1561 (N_1561,In_292,In_484);
and U1562 (N_1562,In_694,In_375);
nand U1563 (N_1563,In_509,In_103);
nand U1564 (N_1564,In_390,In_944);
nor U1565 (N_1565,In_166,In_735);
nand U1566 (N_1566,In_772,In_178);
nand U1567 (N_1567,In_471,In_650);
nor U1568 (N_1568,In_923,In_757);
nor U1569 (N_1569,In_25,In_16);
or U1570 (N_1570,In_430,In_548);
nor U1571 (N_1571,In_181,In_715);
and U1572 (N_1572,In_592,In_467);
and U1573 (N_1573,In_657,In_92);
nand U1574 (N_1574,In_58,In_966);
nand U1575 (N_1575,In_2,In_930);
nor U1576 (N_1576,In_483,In_519);
nor U1577 (N_1577,In_414,In_30);
nor U1578 (N_1578,In_615,In_217);
xnor U1579 (N_1579,In_719,In_316);
nand U1580 (N_1580,In_250,In_419);
nand U1581 (N_1581,In_886,In_320);
nor U1582 (N_1582,In_498,In_761);
or U1583 (N_1583,In_999,In_130);
nor U1584 (N_1584,In_686,In_464);
and U1585 (N_1585,In_901,In_866);
or U1586 (N_1586,In_864,In_659);
and U1587 (N_1587,In_820,In_573);
xnor U1588 (N_1588,In_32,In_752);
and U1589 (N_1589,In_24,In_417);
or U1590 (N_1590,In_422,In_423);
or U1591 (N_1591,In_276,In_45);
nand U1592 (N_1592,In_336,In_127);
nand U1593 (N_1593,In_926,In_206);
nor U1594 (N_1594,In_436,In_948);
and U1595 (N_1595,In_795,In_19);
or U1596 (N_1596,In_57,In_55);
and U1597 (N_1597,In_920,In_290);
or U1598 (N_1598,In_718,In_12);
and U1599 (N_1599,In_437,In_572);
and U1600 (N_1600,In_556,In_727);
and U1601 (N_1601,In_910,In_526);
nand U1602 (N_1602,In_935,In_242);
and U1603 (N_1603,In_797,In_435);
xnor U1604 (N_1604,In_151,In_906);
and U1605 (N_1605,In_469,In_912);
nand U1606 (N_1606,In_687,In_794);
xnor U1607 (N_1607,In_792,In_129);
nand U1608 (N_1608,In_894,In_833);
and U1609 (N_1609,In_39,In_576);
nor U1610 (N_1610,In_243,In_0);
nand U1611 (N_1611,In_615,In_164);
nand U1612 (N_1612,In_272,In_974);
nor U1613 (N_1613,In_44,In_565);
nor U1614 (N_1614,In_268,In_308);
nor U1615 (N_1615,In_498,In_175);
xnor U1616 (N_1616,In_276,In_382);
nand U1617 (N_1617,In_765,In_729);
nand U1618 (N_1618,In_385,In_849);
xnor U1619 (N_1619,In_977,In_597);
or U1620 (N_1620,In_299,In_605);
or U1621 (N_1621,In_482,In_57);
and U1622 (N_1622,In_211,In_520);
and U1623 (N_1623,In_533,In_72);
nor U1624 (N_1624,In_999,In_169);
and U1625 (N_1625,In_389,In_820);
nor U1626 (N_1626,In_434,In_60);
nor U1627 (N_1627,In_208,In_391);
nand U1628 (N_1628,In_406,In_409);
nand U1629 (N_1629,In_688,In_406);
nand U1630 (N_1630,In_420,In_202);
nand U1631 (N_1631,In_675,In_441);
xor U1632 (N_1632,In_410,In_690);
nor U1633 (N_1633,In_66,In_987);
or U1634 (N_1634,In_73,In_345);
xor U1635 (N_1635,In_225,In_48);
and U1636 (N_1636,In_870,In_33);
nand U1637 (N_1637,In_903,In_448);
xor U1638 (N_1638,In_980,In_454);
nand U1639 (N_1639,In_241,In_550);
nor U1640 (N_1640,In_54,In_149);
nand U1641 (N_1641,In_25,In_436);
nor U1642 (N_1642,In_180,In_956);
nor U1643 (N_1643,In_611,In_607);
nand U1644 (N_1644,In_669,In_574);
nor U1645 (N_1645,In_991,In_987);
nand U1646 (N_1646,In_465,In_184);
nand U1647 (N_1647,In_233,In_172);
and U1648 (N_1648,In_772,In_22);
nand U1649 (N_1649,In_373,In_593);
or U1650 (N_1650,In_651,In_498);
and U1651 (N_1651,In_998,In_25);
nor U1652 (N_1652,In_773,In_5);
or U1653 (N_1653,In_428,In_57);
and U1654 (N_1654,In_566,In_108);
and U1655 (N_1655,In_687,In_514);
nor U1656 (N_1656,In_206,In_820);
and U1657 (N_1657,In_202,In_61);
nand U1658 (N_1658,In_379,In_759);
or U1659 (N_1659,In_324,In_150);
xor U1660 (N_1660,In_378,In_679);
or U1661 (N_1661,In_220,In_376);
xnor U1662 (N_1662,In_480,In_952);
nor U1663 (N_1663,In_374,In_93);
and U1664 (N_1664,In_965,In_997);
and U1665 (N_1665,In_978,In_849);
and U1666 (N_1666,In_650,In_333);
nand U1667 (N_1667,In_550,In_568);
nand U1668 (N_1668,In_50,In_88);
nor U1669 (N_1669,In_568,In_910);
nand U1670 (N_1670,In_559,In_625);
nor U1671 (N_1671,In_476,In_803);
and U1672 (N_1672,In_842,In_815);
or U1673 (N_1673,In_989,In_887);
and U1674 (N_1674,In_304,In_55);
and U1675 (N_1675,In_429,In_417);
nor U1676 (N_1676,In_125,In_501);
nor U1677 (N_1677,In_373,In_722);
and U1678 (N_1678,In_518,In_772);
nor U1679 (N_1679,In_158,In_35);
nand U1680 (N_1680,In_634,In_721);
and U1681 (N_1681,In_445,In_495);
xnor U1682 (N_1682,In_250,In_569);
and U1683 (N_1683,In_249,In_255);
or U1684 (N_1684,In_579,In_170);
nand U1685 (N_1685,In_806,In_715);
or U1686 (N_1686,In_676,In_295);
xor U1687 (N_1687,In_920,In_195);
nand U1688 (N_1688,In_485,In_155);
nand U1689 (N_1689,In_317,In_110);
and U1690 (N_1690,In_922,In_713);
or U1691 (N_1691,In_931,In_34);
nor U1692 (N_1692,In_14,In_360);
nand U1693 (N_1693,In_956,In_19);
and U1694 (N_1694,In_174,In_686);
or U1695 (N_1695,In_215,In_646);
nand U1696 (N_1696,In_150,In_250);
and U1697 (N_1697,In_733,In_278);
xor U1698 (N_1698,In_127,In_853);
and U1699 (N_1699,In_71,In_93);
or U1700 (N_1700,In_264,In_890);
or U1701 (N_1701,In_141,In_92);
and U1702 (N_1702,In_297,In_465);
and U1703 (N_1703,In_438,In_213);
and U1704 (N_1704,In_568,In_712);
xor U1705 (N_1705,In_2,In_322);
nand U1706 (N_1706,In_882,In_374);
nor U1707 (N_1707,In_424,In_501);
xnor U1708 (N_1708,In_159,In_826);
or U1709 (N_1709,In_500,In_29);
and U1710 (N_1710,In_568,In_607);
or U1711 (N_1711,In_549,In_592);
or U1712 (N_1712,In_308,In_162);
or U1713 (N_1713,In_875,In_750);
nor U1714 (N_1714,In_466,In_637);
nand U1715 (N_1715,In_536,In_482);
xor U1716 (N_1716,In_511,In_787);
or U1717 (N_1717,In_940,In_520);
nor U1718 (N_1718,In_2,In_853);
or U1719 (N_1719,In_982,In_478);
nand U1720 (N_1720,In_697,In_333);
nand U1721 (N_1721,In_776,In_344);
nor U1722 (N_1722,In_336,In_855);
nand U1723 (N_1723,In_383,In_395);
and U1724 (N_1724,In_285,In_566);
and U1725 (N_1725,In_835,In_781);
and U1726 (N_1726,In_632,In_361);
nor U1727 (N_1727,In_555,In_755);
nand U1728 (N_1728,In_0,In_23);
and U1729 (N_1729,In_23,In_243);
xor U1730 (N_1730,In_327,In_983);
and U1731 (N_1731,In_646,In_528);
and U1732 (N_1732,In_34,In_760);
nand U1733 (N_1733,In_30,In_215);
nor U1734 (N_1734,In_145,In_16);
nand U1735 (N_1735,In_313,In_647);
or U1736 (N_1736,In_74,In_453);
nor U1737 (N_1737,In_196,In_714);
or U1738 (N_1738,In_180,In_373);
xnor U1739 (N_1739,In_952,In_615);
nor U1740 (N_1740,In_496,In_395);
xor U1741 (N_1741,In_995,In_816);
nor U1742 (N_1742,In_331,In_740);
and U1743 (N_1743,In_512,In_954);
and U1744 (N_1744,In_968,In_382);
or U1745 (N_1745,In_354,In_305);
xor U1746 (N_1746,In_602,In_691);
or U1747 (N_1747,In_815,In_320);
xor U1748 (N_1748,In_24,In_834);
and U1749 (N_1749,In_431,In_727);
and U1750 (N_1750,In_784,In_167);
and U1751 (N_1751,In_327,In_607);
or U1752 (N_1752,In_149,In_324);
and U1753 (N_1753,In_12,In_800);
or U1754 (N_1754,In_622,In_346);
xor U1755 (N_1755,In_998,In_15);
nor U1756 (N_1756,In_60,In_518);
nand U1757 (N_1757,In_103,In_326);
nor U1758 (N_1758,In_400,In_422);
or U1759 (N_1759,In_395,In_256);
or U1760 (N_1760,In_447,In_85);
and U1761 (N_1761,In_313,In_862);
or U1762 (N_1762,In_589,In_881);
nor U1763 (N_1763,In_519,In_553);
or U1764 (N_1764,In_679,In_994);
or U1765 (N_1765,In_342,In_870);
nor U1766 (N_1766,In_797,In_454);
and U1767 (N_1767,In_368,In_933);
nand U1768 (N_1768,In_513,In_571);
or U1769 (N_1769,In_207,In_917);
nand U1770 (N_1770,In_778,In_430);
nand U1771 (N_1771,In_27,In_306);
nor U1772 (N_1772,In_822,In_660);
nor U1773 (N_1773,In_874,In_214);
or U1774 (N_1774,In_315,In_514);
nand U1775 (N_1775,In_997,In_156);
or U1776 (N_1776,In_355,In_555);
xor U1777 (N_1777,In_516,In_391);
nor U1778 (N_1778,In_386,In_615);
and U1779 (N_1779,In_253,In_795);
nor U1780 (N_1780,In_904,In_393);
nor U1781 (N_1781,In_962,In_73);
nand U1782 (N_1782,In_381,In_245);
nand U1783 (N_1783,In_970,In_58);
nand U1784 (N_1784,In_407,In_286);
nor U1785 (N_1785,In_321,In_370);
and U1786 (N_1786,In_154,In_795);
and U1787 (N_1787,In_768,In_734);
nor U1788 (N_1788,In_748,In_332);
or U1789 (N_1789,In_234,In_895);
and U1790 (N_1790,In_940,In_436);
and U1791 (N_1791,In_983,In_860);
or U1792 (N_1792,In_292,In_406);
and U1793 (N_1793,In_596,In_196);
and U1794 (N_1794,In_728,In_947);
nor U1795 (N_1795,In_564,In_38);
and U1796 (N_1796,In_910,In_355);
or U1797 (N_1797,In_497,In_260);
xor U1798 (N_1798,In_146,In_883);
nor U1799 (N_1799,In_659,In_317);
nand U1800 (N_1800,In_945,In_378);
nand U1801 (N_1801,In_592,In_972);
or U1802 (N_1802,In_546,In_778);
nand U1803 (N_1803,In_55,In_259);
nand U1804 (N_1804,In_570,In_70);
xnor U1805 (N_1805,In_561,In_223);
and U1806 (N_1806,In_980,In_549);
nor U1807 (N_1807,In_945,In_23);
and U1808 (N_1808,In_120,In_719);
xnor U1809 (N_1809,In_639,In_261);
or U1810 (N_1810,In_963,In_945);
or U1811 (N_1811,In_224,In_225);
or U1812 (N_1812,In_975,In_33);
and U1813 (N_1813,In_51,In_169);
or U1814 (N_1814,In_458,In_118);
nor U1815 (N_1815,In_653,In_276);
and U1816 (N_1816,In_275,In_265);
and U1817 (N_1817,In_637,In_49);
nand U1818 (N_1818,In_266,In_141);
xnor U1819 (N_1819,In_130,In_454);
or U1820 (N_1820,In_190,In_124);
and U1821 (N_1821,In_966,In_351);
nor U1822 (N_1822,In_700,In_459);
and U1823 (N_1823,In_691,In_714);
or U1824 (N_1824,In_493,In_229);
nand U1825 (N_1825,In_910,In_26);
and U1826 (N_1826,In_186,In_13);
and U1827 (N_1827,In_471,In_424);
and U1828 (N_1828,In_129,In_306);
nor U1829 (N_1829,In_643,In_929);
or U1830 (N_1830,In_512,In_117);
xor U1831 (N_1831,In_329,In_240);
and U1832 (N_1832,In_155,In_230);
nor U1833 (N_1833,In_493,In_920);
or U1834 (N_1834,In_611,In_600);
xnor U1835 (N_1835,In_763,In_144);
nand U1836 (N_1836,In_796,In_891);
and U1837 (N_1837,In_923,In_696);
xnor U1838 (N_1838,In_469,In_766);
nor U1839 (N_1839,In_795,In_538);
or U1840 (N_1840,In_660,In_14);
nor U1841 (N_1841,In_966,In_314);
and U1842 (N_1842,In_584,In_38);
or U1843 (N_1843,In_852,In_505);
nor U1844 (N_1844,In_327,In_810);
and U1845 (N_1845,In_92,In_533);
nand U1846 (N_1846,In_76,In_24);
nand U1847 (N_1847,In_564,In_263);
nand U1848 (N_1848,In_450,In_395);
nor U1849 (N_1849,In_762,In_618);
and U1850 (N_1850,In_527,In_265);
or U1851 (N_1851,In_908,In_14);
or U1852 (N_1852,In_681,In_45);
nor U1853 (N_1853,In_843,In_174);
nand U1854 (N_1854,In_595,In_978);
and U1855 (N_1855,In_715,In_869);
and U1856 (N_1856,In_164,In_479);
nand U1857 (N_1857,In_537,In_458);
and U1858 (N_1858,In_504,In_546);
nor U1859 (N_1859,In_185,In_426);
or U1860 (N_1860,In_101,In_444);
or U1861 (N_1861,In_911,In_385);
nor U1862 (N_1862,In_808,In_597);
and U1863 (N_1863,In_692,In_773);
xnor U1864 (N_1864,In_37,In_819);
or U1865 (N_1865,In_197,In_643);
nand U1866 (N_1866,In_422,In_101);
or U1867 (N_1867,In_451,In_266);
or U1868 (N_1868,In_633,In_598);
xnor U1869 (N_1869,In_883,In_159);
and U1870 (N_1870,In_188,In_758);
nor U1871 (N_1871,In_779,In_64);
or U1872 (N_1872,In_615,In_274);
nor U1873 (N_1873,In_173,In_75);
nor U1874 (N_1874,In_29,In_209);
nand U1875 (N_1875,In_308,In_305);
or U1876 (N_1876,In_683,In_260);
nand U1877 (N_1877,In_488,In_893);
nor U1878 (N_1878,In_728,In_576);
or U1879 (N_1879,In_876,In_962);
and U1880 (N_1880,In_641,In_271);
or U1881 (N_1881,In_502,In_95);
and U1882 (N_1882,In_613,In_703);
nor U1883 (N_1883,In_168,In_740);
or U1884 (N_1884,In_944,In_976);
nor U1885 (N_1885,In_287,In_918);
and U1886 (N_1886,In_39,In_336);
nor U1887 (N_1887,In_762,In_572);
and U1888 (N_1888,In_903,In_695);
and U1889 (N_1889,In_983,In_196);
and U1890 (N_1890,In_612,In_382);
or U1891 (N_1891,In_616,In_93);
or U1892 (N_1892,In_282,In_289);
nand U1893 (N_1893,In_950,In_921);
or U1894 (N_1894,In_851,In_755);
nand U1895 (N_1895,In_237,In_425);
or U1896 (N_1896,In_251,In_953);
and U1897 (N_1897,In_509,In_61);
nand U1898 (N_1898,In_577,In_446);
xor U1899 (N_1899,In_230,In_925);
xnor U1900 (N_1900,In_793,In_391);
nand U1901 (N_1901,In_935,In_12);
nor U1902 (N_1902,In_402,In_381);
nand U1903 (N_1903,In_165,In_504);
or U1904 (N_1904,In_636,In_829);
nor U1905 (N_1905,In_47,In_649);
nor U1906 (N_1906,In_547,In_344);
nor U1907 (N_1907,In_150,In_354);
and U1908 (N_1908,In_464,In_178);
or U1909 (N_1909,In_647,In_504);
xnor U1910 (N_1910,In_931,In_63);
nor U1911 (N_1911,In_753,In_892);
xnor U1912 (N_1912,In_196,In_283);
nor U1913 (N_1913,In_372,In_71);
and U1914 (N_1914,In_607,In_510);
nand U1915 (N_1915,In_243,In_520);
and U1916 (N_1916,In_688,In_783);
or U1917 (N_1917,In_454,In_895);
or U1918 (N_1918,In_94,In_609);
xnor U1919 (N_1919,In_712,In_66);
and U1920 (N_1920,In_672,In_907);
xnor U1921 (N_1921,In_281,In_446);
xor U1922 (N_1922,In_762,In_118);
and U1923 (N_1923,In_15,In_84);
or U1924 (N_1924,In_911,In_557);
or U1925 (N_1925,In_671,In_884);
nand U1926 (N_1926,In_970,In_639);
or U1927 (N_1927,In_540,In_545);
nor U1928 (N_1928,In_664,In_310);
nand U1929 (N_1929,In_567,In_312);
nor U1930 (N_1930,In_29,In_404);
xor U1931 (N_1931,In_277,In_346);
or U1932 (N_1932,In_757,In_707);
nand U1933 (N_1933,In_181,In_694);
nand U1934 (N_1934,In_326,In_676);
nor U1935 (N_1935,In_591,In_589);
nor U1936 (N_1936,In_67,In_422);
nor U1937 (N_1937,In_754,In_636);
or U1938 (N_1938,In_925,In_467);
and U1939 (N_1939,In_816,In_474);
nand U1940 (N_1940,In_776,In_500);
nor U1941 (N_1941,In_28,In_180);
nand U1942 (N_1942,In_40,In_210);
nor U1943 (N_1943,In_598,In_321);
nand U1944 (N_1944,In_691,In_583);
or U1945 (N_1945,In_724,In_507);
or U1946 (N_1946,In_493,In_906);
or U1947 (N_1947,In_711,In_624);
xnor U1948 (N_1948,In_586,In_982);
nand U1949 (N_1949,In_745,In_503);
nor U1950 (N_1950,In_109,In_531);
or U1951 (N_1951,In_10,In_252);
nor U1952 (N_1952,In_259,In_612);
nand U1953 (N_1953,In_948,In_38);
and U1954 (N_1954,In_171,In_157);
nor U1955 (N_1955,In_896,In_889);
and U1956 (N_1956,In_831,In_786);
nand U1957 (N_1957,In_326,In_995);
or U1958 (N_1958,In_764,In_561);
or U1959 (N_1959,In_438,In_316);
nand U1960 (N_1960,In_420,In_4);
nand U1961 (N_1961,In_549,In_46);
or U1962 (N_1962,In_941,In_221);
nand U1963 (N_1963,In_620,In_46);
or U1964 (N_1964,In_824,In_528);
xor U1965 (N_1965,In_404,In_348);
nor U1966 (N_1966,In_736,In_894);
and U1967 (N_1967,In_663,In_244);
nand U1968 (N_1968,In_696,In_435);
nor U1969 (N_1969,In_401,In_363);
nand U1970 (N_1970,In_553,In_485);
or U1971 (N_1971,In_142,In_68);
and U1972 (N_1972,In_928,In_96);
or U1973 (N_1973,In_208,In_517);
xnor U1974 (N_1974,In_656,In_4);
and U1975 (N_1975,In_827,In_836);
xor U1976 (N_1976,In_412,In_606);
nor U1977 (N_1977,In_388,In_665);
xor U1978 (N_1978,In_758,In_114);
nand U1979 (N_1979,In_833,In_799);
nand U1980 (N_1980,In_893,In_719);
and U1981 (N_1981,In_93,In_756);
nor U1982 (N_1982,In_995,In_754);
and U1983 (N_1983,In_22,In_839);
nand U1984 (N_1984,In_270,In_494);
and U1985 (N_1985,In_69,In_96);
or U1986 (N_1986,In_353,In_141);
and U1987 (N_1987,In_340,In_147);
or U1988 (N_1988,In_253,In_489);
or U1989 (N_1989,In_513,In_975);
nor U1990 (N_1990,In_0,In_344);
or U1991 (N_1991,In_662,In_707);
nand U1992 (N_1992,In_685,In_139);
and U1993 (N_1993,In_669,In_677);
and U1994 (N_1994,In_638,In_74);
or U1995 (N_1995,In_496,In_520);
nor U1996 (N_1996,In_947,In_424);
nor U1997 (N_1997,In_38,In_300);
and U1998 (N_1998,In_920,In_800);
xor U1999 (N_1999,In_406,In_604);
nand U2000 (N_2000,N_860,N_1851);
nand U2001 (N_2001,N_587,N_403);
or U2002 (N_2002,N_424,N_1737);
nor U2003 (N_2003,N_1452,N_489);
nor U2004 (N_2004,N_135,N_1540);
nand U2005 (N_2005,N_1509,N_1927);
xnor U2006 (N_2006,N_1777,N_1317);
nor U2007 (N_2007,N_166,N_399);
nand U2008 (N_2008,N_625,N_280);
or U2009 (N_2009,N_303,N_1002);
nor U2010 (N_2010,N_691,N_1235);
nand U2011 (N_2011,N_1579,N_51);
nand U2012 (N_2012,N_996,N_769);
nand U2013 (N_2013,N_277,N_900);
nand U2014 (N_2014,N_989,N_777);
and U2015 (N_2015,N_2,N_1888);
or U2016 (N_2016,N_984,N_1792);
nor U2017 (N_2017,N_1050,N_1342);
nand U2018 (N_2018,N_288,N_351);
or U2019 (N_2019,N_445,N_1121);
nor U2020 (N_2020,N_455,N_1323);
or U2021 (N_2021,N_1654,N_460);
xnor U2022 (N_2022,N_1392,N_862);
nor U2023 (N_2023,N_1192,N_606);
or U2024 (N_2024,N_1567,N_1784);
and U2025 (N_2025,N_114,N_1372);
nor U2026 (N_2026,N_884,N_1904);
nor U2027 (N_2027,N_1443,N_822);
xnor U2028 (N_2028,N_196,N_1412);
xnor U2029 (N_2029,N_440,N_975);
nand U2030 (N_2030,N_343,N_144);
nor U2031 (N_2031,N_1610,N_364);
and U2032 (N_2032,N_827,N_447);
and U2033 (N_2033,N_917,N_892);
nand U2034 (N_2034,N_1653,N_681);
and U2035 (N_2035,N_1755,N_700);
nand U2036 (N_2036,N_966,N_733);
xnor U2037 (N_2037,N_102,N_1574);
nand U2038 (N_2038,N_394,N_886);
and U2039 (N_2039,N_1467,N_395);
nand U2040 (N_2040,N_901,N_1133);
nand U2041 (N_2041,N_575,N_1001);
nor U2042 (N_2042,N_1542,N_744);
nand U2043 (N_2043,N_1606,N_1296);
xor U2044 (N_2044,N_1259,N_1332);
nand U2045 (N_2045,N_171,N_1781);
nor U2046 (N_2046,N_1665,N_1562);
nor U2047 (N_2047,N_520,N_1499);
nor U2048 (N_2048,N_168,N_1803);
and U2049 (N_2049,N_1080,N_95);
nor U2050 (N_2050,N_327,N_1544);
xnor U2051 (N_2051,N_956,N_300);
xor U2052 (N_2052,N_127,N_1970);
or U2053 (N_2053,N_1246,N_1437);
nand U2054 (N_2054,N_1686,N_1885);
and U2055 (N_2055,N_991,N_1575);
nor U2056 (N_2056,N_1295,N_845);
nor U2057 (N_2057,N_388,N_465);
or U2058 (N_2058,N_1596,N_1682);
nand U2059 (N_2059,N_41,N_1367);
nand U2060 (N_2060,N_1420,N_1361);
nand U2061 (N_2061,N_70,N_32);
or U2062 (N_2062,N_1961,N_1503);
xor U2063 (N_2063,N_1256,N_1478);
nor U2064 (N_2064,N_1331,N_368);
nand U2065 (N_2065,N_1647,N_940);
and U2066 (N_2066,N_45,N_220);
nor U2067 (N_2067,N_1841,N_1356);
nor U2068 (N_2068,N_232,N_1699);
nand U2069 (N_2069,N_215,N_672);
nor U2070 (N_2070,N_1,N_741);
and U2071 (N_2071,N_1787,N_354);
nand U2072 (N_2072,N_1152,N_407);
nand U2073 (N_2073,N_582,N_1563);
nor U2074 (N_2074,N_1740,N_67);
nand U2075 (N_2075,N_954,N_1585);
xor U2076 (N_2076,N_12,N_835);
nor U2077 (N_2077,N_1390,N_522);
nand U2078 (N_2078,N_1383,N_23);
or U2079 (N_2079,N_689,N_1117);
nand U2080 (N_2080,N_255,N_995);
nor U2081 (N_2081,N_1462,N_252);
or U2082 (N_2082,N_571,N_361);
and U2083 (N_2083,N_628,N_10);
nor U2084 (N_2084,N_1779,N_355);
nor U2085 (N_2085,N_1601,N_646);
or U2086 (N_2086,N_1400,N_273);
xor U2087 (N_2087,N_62,N_1962);
or U2088 (N_2088,N_1953,N_534);
xnor U2089 (N_2089,N_799,N_1111);
nor U2090 (N_2090,N_332,N_473);
nand U2091 (N_2091,N_627,N_307);
nand U2092 (N_2092,N_1382,N_1440);
nor U2093 (N_2093,N_226,N_269);
nand U2094 (N_2094,N_1725,N_877);
or U2095 (N_2095,N_1529,N_1285);
or U2096 (N_2096,N_1661,N_536);
nor U2097 (N_2097,N_205,N_561);
and U2098 (N_2098,N_391,N_1715);
xnor U2099 (N_2099,N_322,N_134);
and U2100 (N_2100,N_1243,N_65);
and U2101 (N_2101,N_1979,N_1046);
or U2102 (N_2102,N_920,N_640);
or U2103 (N_2103,N_420,N_314);
or U2104 (N_2104,N_339,N_1335);
nor U2105 (N_2105,N_239,N_551);
and U2106 (N_2106,N_129,N_121);
xor U2107 (N_2107,N_532,N_510);
nand U2108 (N_2108,N_804,N_519);
nand U2109 (N_2109,N_881,N_1968);
or U2110 (N_2110,N_1286,N_1198);
and U2111 (N_2111,N_1848,N_1639);
and U2112 (N_2112,N_1708,N_500);
xor U2113 (N_2113,N_1631,N_1265);
or U2114 (N_2114,N_1926,N_340);
or U2115 (N_2115,N_139,N_1778);
or U2116 (N_2116,N_1284,N_1195);
and U2117 (N_2117,N_1652,N_1569);
and U2118 (N_2118,N_308,N_1441);
or U2119 (N_2119,N_858,N_83);
nand U2120 (N_2120,N_1838,N_883);
or U2121 (N_2121,N_381,N_126);
xnor U2122 (N_2122,N_542,N_1869);
nor U2123 (N_2123,N_1860,N_44);
nand U2124 (N_2124,N_1167,N_371);
or U2125 (N_2125,N_7,N_410);
nand U2126 (N_2126,N_261,N_824);
and U2127 (N_2127,N_369,N_934);
and U2128 (N_2128,N_1809,N_1379);
xor U2129 (N_2129,N_572,N_1616);
nor U2130 (N_2130,N_665,N_1757);
nor U2131 (N_2131,N_1124,N_1621);
nor U2132 (N_2132,N_1608,N_1704);
and U2133 (N_2133,N_412,N_1615);
or U2134 (N_2134,N_1197,N_376);
nand U2135 (N_2135,N_604,N_1714);
or U2136 (N_2136,N_96,N_867);
nor U2137 (N_2137,N_1942,N_755);
nand U2138 (N_2138,N_1388,N_1836);
and U2139 (N_2139,N_1060,N_1173);
nand U2140 (N_2140,N_613,N_1721);
nor U2141 (N_2141,N_295,N_33);
and U2142 (N_2142,N_549,N_1224);
nand U2143 (N_2143,N_698,N_1157);
nand U2144 (N_2144,N_1949,N_1547);
nand U2145 (N_2145,N_298,N_885);
or U2146 (N_2146,N_999,N_91);
nor U2147 (N_2147,N_526,N_49);
xor U2148 (N_2148,N_1564,N_1552);
nor U2149 (N_2149,N_882,N_1933);
xor U2150 (N_2150,N_941,N_1957);
and U2151 (N_2151,N_1676,N_1096);
nand U2152 (N_2152,N_1716,N_262);
nor U2153 (N_2153,N_400,N_1360);
and U2154 (N_2154,N_1928,N_1186);
nand U2155 (N_2155,N_1166,N_710);
nand U2156 (N_2156,N_1067,N_406);
and U2157 (N_2157,N_229,N_37);
nand U2158 (N_2158,N_1362,N_964);
nand U2159 (N_2159,N_1255,N_776);
or U2160 (N_2160,N_939,N_1354);
and U2161 (N_2161,N_1233,N_1706);
or U2162 (N_2162,N_619,N_586);
nor U2163 (N_2163,N_1738,N_1930);
and U2164 (N_2164,N_231,N_1799);
or U2165 (N_2165,N_800,N_1808);
or U2166 (N_2166,N_1558,N_1835);
xnor U2167 (N_2167,N_1075,N_570);
or U2168 (N_2168,N_1132,N_50);
xnor U2169 (N_2169,N_1064,N_1000);
or U2170 (N_2170,N_1688,N_1758);
nand U2171 (N_2171,N_1883,N_396);
xor U2172 (N_2172,N_1505,N_1232);
and U2173 (N_2173,N_1022,N_1351);
xor U2174 (N_2174,N_1328,N_848);
nor U2175 (N_2175,N_812,N_1827);
and U2176 (N_2176,N_1076,N_417);
nand U2177 (N_2177,N_228,N_1833);
nand U2178 (N_2178,N_1346,N_1753);
xnor U2179 (N_2179,N_927,N_953);
or U2180 (N_2180,N_1998,N_1337);
nand U2181 (N_2181,N_1468,N_906);
and U2182 (N_2182,N_743,N_603);
or U2183 (N_2183,N_969,N_874);
and U2184 (N_2184,N_488,N_1845);
xor U2185 (N_2185,N_1685,N_1789);
or U2186 (N_2186,N_767,N_290);
and U2187 (N_2187,N_1782,N_285);
nand U2188 (N_2188,N_1710,N_1761);
xnor U2189 (N_2189,N_1153,N_260);
nand U2190 (N_2190,N_85,N_631);
and U2191 (N_2191,N_110,N_630);
nor U2192 (N_2192,N_955,N_1459);
and U2193 (N_2193,N_1625,N_1174);
and U2194 (N_2194,N_1967,N_1623);
or U2195 (N_2195,N_1150,N_543);
nor U2196 (N_2196,N_612,N_1774);
nand U2197 (N_2197,N_1538,N_1668);
nor U2198 (N_2198,N_516,N_1856);
and U2199 (N_2199,N_1539,N_1937);
or U2200 (N_2200,N_1965,N_1003);
xnor U2201 (N_2201,N_851,N_125);
and U2202 (N_2202,N_513,N_1450);
or U2203 (N_2203,N_373,N_187);
nand U2204 (N_2204,N_1023,N_374);
or U2205 (N_2205,N_912,N_1090);
xnor U2206 (N_2206,N_1029,N_584);
nand U2207 (N_2207,N_1995,N_1840);
nand U2208 (N_2208,N_1873,N_103);
nand U2209 (N_2209,N_263,N_819);
and U2210 (N_2210,N_347,N_1414);
nand U2211 (N_2211,N_1815,N_1047);
and U2212 (N_2212,N_676,N_820);
nor U2213 (N_2213,N_1274,N_565);
nand U2214 (N_2214,N_28,N_435);
or U2215 (N_2215,N_1911,N_1814);
nand U2216 (N_2216,N_734,N_358);
nor U2217 (N_2217,N_1674,N_1748);
xor U2218 (N_2218,N_133,N_1336);
nand U2219 (N_2219,N_1291,N_19);
xor U2220 (N_2220,N_1453,N_1999);
nor U2221 (N_2221,N_155,N_1822);
nor U2222 (N_2222,N_1614,N_605);
or U2223 (N_2223,N_1300,N_1093);
nand U2224 (N_2224,N_742,N_931);
or U2225 (N_2225,N_496,N_1726);
or U2226 (N_2226,N_1272,N_675);
or U2227 (N_2227,N_1791,N_1397);
xnor U2228 (N_2228,N_1380,N_1984);
or U2229 (N_2229,N_498,N_137);
nand U2230 (N_2230,N_1114,N_1294);
and U2231 (N_2231,N_740,N_384);
nor U2232 (N_2232,N_177,N_1470);
and U2233 (N_2233,N_1702,N_11);
nand U2234 (N_2234,N_1680,N_1363);
and U2235 (N_2235,N_952,N_1551);
nand U2236 (N_2236,N_366,N_538);
or U2237 (N_2237,N_926,N_1734);
nor U2238 (N_2238,N_596,N_1769);
or U2239 (N_2239,N_879,N_1182);
and U2240 (N_2240,N_1583,N_1496);
or U2241 (N_2241,N_1707,N_203);
or U2242 (N_2242,N_836,N_1430);
nor U2243 (N_2243,N_302,N_1333);
and U2244 (N_2244,N_1568,N_105);
and U2245 (N_2245,N_4,N_599);
and U2246 (N_2246,N_1491,N_1107);
and U2247 (N_2247,N_1048,N_1472);
and U2248 (N_2248,N_1550,N_705);
and U2249 (N_2249,N_722,N_1370);
xor U2250 (N_2250,N_1587,N_552);
nand U2251 (N_2251,N_1811,N_1717);
xnor U2252 (N_2252,N_1507,N_1994);
or U2253 (N_2253,N_897,N_271);
nor U2254 (N_2254,N_718,N_1749);
nand U2255 (N_2255,N_622,N_1905);
xor U2256 (N_2256,N_918,N_1410);
nor U2257 (N_2257,N_1655,N_1277);
nand U2258 (N_2258,N_701,N_1218);
and U2259 (N_2259,N_795,N_186);
nor U2260 (N_2260,N_462,N_773);
nor U2261 (N_2261,N_113,N_1373);
and U2262 (N_2262,N_1730,N_1896);
nand U2263 (N_2263,N_654,N_1626);
or U2264 (N_2264,N_1620,N_1693);
nor U2265 (N_2265,N_1508,N_1581);
or U2266 (N_2266,N_1502,N_1052);
or U2267 (N_2267,N_806,N_1040);
xor U2268 (N_2268,N_120,N_1057);
or U2269 (N_2269,N_1722,N_1215);
nor U2270 (N_2270,N_1698,N_1493);
or U2271 (N_2271,N_1490,N_1617);
nand U2272 (N_2272,N_1138,N_148);
nor U2273 (N_2273,N_1108,N_151);
and U2274 (N_2274,N_149,N_1591);
and U2275 (N_2275,N_1832,N_1872);
xor U2276 (N_2276,N_330,N_1589);
or U2277 (N_2277,N_1425,N_219);
and U2278 (N_2278,N_905,N_726);
nand U2279 (N_2279,N_1797,N_1104);
or U2280 (N_2280,N_567,N_1147);
nor U2281 (N_2281,N_725,N_241);
nor U2282 (N_2282,N_1555,N_224);
xnor U2283 (N_2283,N_1357,N_1062);
and U2284 (N_2284,N_1237,N_639);
or U2285 (N_2285,N_1011,N_559);
and U2286 (N_2286,N_1164,N_75);
and U2287 (N_2287,N_1162,N_1109);
nand U2288 (N_2288,N_175,N_79);
and U2289 (N_2289,N_1487,N_982);
and U2290 (N_2290,N_216,N_664);
or U2291 (N_2291,N_475,N_1158);
and U2292 (N_2292,N_974,N_1348);
nand U2293 (N_2293,N_658,N_1917);
and U2294 (N_2294,N_590,N_1433);
or U2295 (N_2295,N_833,N_597);
and U2296 (N_2296,N_257,N_641);
and U2297 (N_2297,N_317,N_674);
nor U2298 (N_2298,N_185,N_1458);
and U2299 (N_2299,N_1257,N_739);
and U2300 (N_2300,N_528,N_221);
nand U2301 (N_2301,N_181,N_1375);
or U2302 (N_2302,N_342,N_487);
and U2303 (N_2303,N_20,N_266);
nor U2304 (N_2304,N_404,N_985);
nand U2305 (N_2305,N_558,N_486);
nor U2306 (N_2306,N_1553,N_1130);
nor U2307 (N_2307,N_579,N_1514);
nor U2308 (N_2308,N_5,N_1322);
xor U2309 (N_2309,N_1353,N_1172);
or U2310 (N_2310,N_467,N_1584);
and U2311 (N_2311,N_1225,N_1184);
or U2312 (N_2312,N_1202,N_642);
and U2313 (N_2313,N_670,N_425);
and U2314 (N_2314,N_1878,N_682);
nand U2315 (N_2315,N_1679,N_1981);
nand U2316 (N_2316,N_1389,N_87);
and U2317 (N_2317,N_1033,N_306);
and U2318 (N_2318,N_1319,N_696);
xnor U2319 (N_2319,N_140,N_413);
nand U2320 (N_2320,N_873,N_1424);
nand U2321 (N_2321,N_1203,N_299);
and U2322 (N_2322,N_1051,N_461);
nor U2323 (N_2323,N_916,N_281);
nor U2324 (N_2324,N_169,N_711);
or U2325 (N_2325,N_297,N_1145);
or U2326 (N_2326,N_434,N_539);
or U2327 (N_2327,N_397,N_1220);
nor U2328 (N_2328,N_1398,N_1943);
nand U2329 (N_2329,N_53,N_673);
or U2330 (N_2330,N_826,N_1898);
or U2331 (N_2331,N_1377,N_786);
nor U2332 (N_2332,N_199,N_703);
or U2333 (N_2333,N_153,N_663);
and U2334 (N_2334,N_1670,N_644);
and U2335 (N_2335,N_1071,N_138);
or U2336 (N_2336,N_1985,N_762);
xnor U2337 (N_2337,N_1381,N_1513);
nor U2338 (N_2338,N_1316,N_1326);
xor U2339 (N_2339,N_1429,N_1149);
xor U2340 (N_2340,N_145,N_535);
nand U2341 (N_2341,N_1378,N_1207);
and U2342 (N_2342,N_1586,N_338);
nor U2343 (N_2343,N_1177,N_840);
nor U2344 (N_2344,N_24,N_1407);
and U2345 (N_2345,N_853,N_402);
nand U2346 (N_2346,N_1393,N_1650);
and U2347 (N_2347,N_207,N_182);
nand U2348 (N_2348,N_1746,N_1852);
nor U2349 (N_2349,N_328,N_1588);
nor U2350 (N_2350,N_379,N_1084);
nand U2351 (N_2351,N_1298,N_1276);
nor U2352 (N_2352,N_441,N_180);
nand U2353 (N_2353,N_1557,N_1906);
xor U2354 (N_2354,N_1719,N_1843);
xnor U2355 (N_2355,N_1580,N_1638);
nand U2356 (N_2356,N_1475,N_1387);
nor U2357 (N_2357,N_581,N_117);
and U2358 (N_2358,N_1973,N_1364);
and U2359 (N_2359,N_554,N_1017);
nor U2360 (N_2360,N_1773,N_1116);
nand U2361 (N_2361,N_1110,N_1573);
and U2362 (N_2362,N_1989,N_1030);
nor U2363 (N_2363,N_1221,N_815);
or U2364 (N_2364,N_1308,N_669);
nor U2365 (N_2365,N_1924,N_1305);
or U2366 (N_2366,N_1230,N_1528);
nor U2367 (N_2367,N_943,N_809);
nand U2368 (N_2368,N_1394,N_353);
or U2369 (N_2369,N_1947,N_191);
nor U2370 (N_2370,N_63,N_48);
or U2371 (N_2371,N_159,N_997);
or U2372 (N_2372,N_43,N_1935);
nor U2373 (N_2373,N_1582,N_1637);
nand U2374 (N_2374,N_794,N_1635);
and U2375 (N_2375,N_758,N_1537);
nand U2376 (N_2376,N_1471,N_1088);
or U2377 (N_2377,N_1341,N_1729);
and U2378 (N_2378,N_760,N_92);
and U2379 (N_2379,N_751,N_34);
nand U2380 (N_2380,N_408,N_202);
nand U2381 (N_2381,N_825,N_1253);
nor U2382 (N_2382,N_1828,N_1518);
nand U2383 (N_2383,N_278,N_385);
xnor U2384 (N_2384,N_1473,N_949);
nand U2385 (N_2385,N_1409,N_1325);
and U2386 (N_2386,N_1754,N_362);
nor U2387 (N_2387,N_1036,N_389);
or U2388 (N_2388,N_122,N_1194);
nor U2389 (N_2389,N_735,N_1061);
or U2390 (N_2390,N_1041,N_1783);
xor U2391 (N_2391,N_1549,N_1371);
or U2392 (N_2392,N_1876,N_651);
nor U2393 (N_2393,N_1115,N_783);
and U2394 (N_2394,N_1141,N_436);
nand U2395 (N_2395,N_1802,N_1849);
and U2396 (N_2396,N_1850,N_64);
or U2397 (N_2397,N_356,N_1599);
or U2398 (N_2398,N_501,N_1899);
nand U2399 (N_2399,N_282,N_188);
xnor U2400 (N_2400,N_1830,N_512);
nand U2401 (N_2401,N_337,N_275);
nand U2402 (N_2402,N_1098,N_763);
or U2403 (N_2403,N_732,N_1907);
xnor U2404 (N_2404,N_476,N_193);
and U2405 (N_2405,N_1408,N_878);
and U2406 (N_2406,N_1024,N_1415);
nor U2407 (N_2407,N_685,N_929);
and U2408 (N_2408,N_1442,N_68);
and U2409 (N_2409,N_248,N_284);
or U2410 (N_2410,N_707,N_198);
nand U2411 (N_2411,N_1870,N_678);
nor U2412 (N_2412,N_301,N_1944);
nand U2413 (N_2413,N_1511,N_1756);
or U2414 (N_2414,N_1660,N_1304);
nand U2415 (N_2415,N_118,N_1199);
nand U2416 (N_2416,N_178,N_258);
nor U2417 (N_2417,N_59,N_715);
xnor U2418 (N_2418,N_89,N_1500);
nor U2419 (N_2419,N_136,N_474);
nor U2420 (N_2420,N_946,N_1892);
nand U2421 (N_2421,N_1434,N_1628);
or U2422 (N_2422,N_429,N_1846);
and U2423 (N_2423,N_265,N_318);
nor U2424 (N_2424,N_1191,N_348);
and U2425 (N_2425,N_611,N_834);
and U2426 (N_2426,N_1212,N_268);
or U2427 (N_2427,N_405,N_1796);
nor U2428 (N_2428,N_57,N_1690);
xnor U2429 (N_2429,N_1504,N_923);
nand U2430 (N_2430,N_176,N_958);
nand U2431 (N_2431,N_1330,N_1603);
or U2432 (N_2432,N_932,N_1021);
nand U2433 (N_2433,N_1416,N_1054);
or U2434 (N_2434,N_771,N_158);
and U2435 (N_2435,N_810,N_1709);
nand U2436 (N_2436,N_545,N_93);
or U2437 (N_2437,N_1267,N_721);
or U2438 (N_2438,N_147,N_1066);
and U2439 (N_2439,N_30,N_1427);
or U2440 (N_2440,N_817,N_1403);
nand U2441 (N_2441,N_788,N_1019);
and U2442 (N_2442,N_1209,N_1079);
and U2443 (N_2443,N_914,N_709);
and U2444 (N_2444,N_244,N_451);
or U2445 (N_2445,N_54,N_1137);
or U2446 (N_2446,N_568,N_163);
xor U2447 (N_2447,N_1950,N_423);
nand U2448 (N_2448,N_1492,N_66);
and U2449 (N_2449,N_677,N_1893);
nand U2450 (N_2450,N_898,N_1085);
and U2451 (N_2451,N_1718,N_1517);
nand U2452 (N_2452,N_1735,N_1056);
and U2453 (N_2453,N_1094,N_609);
and U2454 (N_2454,N_1752,N_913);
nand U2455 (N_2455,N_1857,N_1102);
nand U2456 (N_2456,N_839,N_1775);
or U2457 (N_2457,N_872,N_1929);
or U2458 (N_2458,N_629,N_793);
nor U2459 (N_2459,N_666,N_1641);
or U2460 (N_2460,N_214,N_1432);
or U2461 (N_2461,N_1327,N_890);
nor U2462 (N_2462,N_1004,N_1572);
and U2463 (N_2463,N_904,N_1886);
and U2464 (N_2464,N_764,N_1270);
and U2465 (N_2465,N_1971,N_1163);
and U2466 (N_2466,N_1016,N_1687);
xor U2467 (N_2467,N_856,N_854);
nand U2468 (N_2468,N_576,N_218);
and U2469 (N_2469,N_493,N_547);
nor U2470 (N_2470,N_1692,N_320);
and U2471 (N_2471,N_598,N_1345);
or U2472 (N_2472,N_1651,N_1866);
nand U2473 (N_2473,N_1315,N_363);
or U2474 (N_2474,N_970,N_1519);
or U2475 (N_2475,N_1463,N_415);
or U2476 (N_2476,N_1607,N_72);
xor U2477 (N_2477,N_588,N_131);
or U2478 (N_2478,N_1139,N_1889);
or U2479 (N_2479,N_1854,N_1664);
nor U2480 (N_2480,N_687,N_124);
nor U2481 (N_2481,N_1684,N_1269);
or U2482 (N_2482,N_821,N_97);
nand U2483 (N_2483,N_1374,N_1307);
nor U2484 (N_2484,N_635,N_1210);
or U2485 (N_2485,N_1633,N_1352);
or U2486 (N_2486,N_1466,N_1701);
nand U2487 (N_2487,N_1855,N_1681);
nor U2488 (N_2488,N_387,N_1858);
nand U2489 (N_2489,N_1161,N_464);
or U2490 (N_2490,N_1421,N_756);
nor U2491 (N_2491,N_1444,N_164);
and U2492 (N_2492,N_645,N_620);
and U2493 (N_2493,N_1314,N_190);
nor U2494 (N_2494,N_1877,N_1489);
nor U2495 (N_2495,N_957,N_580);
or U2496 (N_2496,N_1622,N_1861);
and U2497 (N_2497,N_1891,N_1534);
or U2498 (N_2498,N_1086,N_312);
or U2499 (N_2499,N_1037,N_1901);
or U2500 (N_2500,N_660,N_1611);
and U2501 (N_2501,N_720,N_1329);
or U2502 (N_2502,N_1533,N_1077);
xor U2503 (N_2503,N_1015,N_1516);
and U2504 (N_2504,N_560,N_1816);
or U2505 (N_2505,N_1318,N_749);
xnor U2506 (N_2506,N_963,N_13);
nand U2507 (N_2507,N_1045,N_1188);
or U2508 (N_2508,N_935,N_1183);
nand U2509 (N_2509,N_1916,N_1101);
nor U2510 (N_2510,N_430,N_805);
nor U2511 (N_2511,N_1794,N_634);
nand U2512 (N_2512,N_1919,N_1988);
or U2513 (N_2513,N_761,N_1882);
or U2514 (N_2514,N_746,N_209);
or U2515 (N_2515,N_1922,N_1903);
nand U2516 (N_2516,N_1178,N_695);
and U2517 (N_2517,N_1831,N_514);
or U2518 (N_2518,N_1694,N_1275);
nor U2519 (N_2519,N_1909,N_69);
or U2520 (N_2520,N_52,N_279);
nand U2521 (N_2521,N_889,N_1629);
and U2522 (N_2522,N_1428,N_578);
or U2523 (N_2523,N_1880,N_1932);
xnor U2524 (N_2524,N_1966,N_1817);
xor U2525 (N_2525,N_792,N_71);
and U2526 (N_2526,N_6,N_1862);
nand U2527 (N_2527,N_1590,N_1165);
nor U2528 (N_2528,N_842,N_699);
nand U2529 (N_2529,N_1018,N_787);
and U2530 (N_2530,N_1663,N_837);
or U2531 (N_2531,N_1213,N_636);
or U2532 (N_2532,N_509,N_775);
nand U2533 (N_2533,N_523,N_504);
nor U2534 (N_2534,N_706,N_1271);
xnor U2535 (N_2535,N_36,N_615);
nand U2536 (N_2536,N_1785,N_123);
and U2537 (N_2537,N_1527,N_1081);
nor U2538 (N_2538,N_485,N_1894);
and U2539 (N_2539,N_195,N_716);
or U2540 (N_2540,N_1510,N_1595);
xor U2541 (N_2541,N_1642,N_3);
or U2542 (N_2542,N_1465,N_1263);
or U2543 (N_2543,N_1144,N_1495);
nand U2544 (N_2544,N_909,N_861);
and U2545 (N_2545,N_971,N_1645);
and U2546 (N_2546,N_111,N_938);
xor U2547 (N_2547,N_1560,N_668);
nor U2548 (N_2548,N_116,N_1282);
nand U2549 (N_2549,N_511,N_753);
or U2550 (N_2550,N_1273,N_84);
and U2551 (N_2551,N_1671,N_1405);
or U2552 (N_2552,N_564,N_1767);
nor U2553 (N_2553,N_911,N_1013);
nand U2554 (N_2554,N_823,N_1012);
and U2555 (N_2555,N_313,N_1454);
and U2556 (N_2556,N_1083,N_1976);
and U2557 (N_2557,N_1252,N_614);
and U2558 (N_2558,N_1804,N_569);
and U2559 (N_2559,N_1303,N_998);
nand U2560 (N_2560,N_200,N_637);
xor U2561 (N_2561,N_875,N_891);
or U2562 (N_2562,N_1234,N_211);
nand U2563 (N_2563,N_688,N_1727);
nand U2564 (N_2564,N_1853,N_1630);
nor U2565 (N_2565,N_1526,N_289);
nor U2566 (N_2566,N_1772,N_1521);
and U2567 (N_2567,N_1844,N_517);
or U2568 (N_2568,N_1820,N_375);
nor U2569 (N_2569,N_1447,N_871);
nor U2570 (N_2570,N_161,N_907);
and U2571 (N_2571,N_1515,N_350);
or U2572 (N_2572,N_194,N_1055);
and U2573 (N_2573,N_1476,N_254);
nand U2574 (N_2574,N_1936,N_479);
or U2575 (N_2575,N_903,N_1952);
nor U2576 (N_2576,N_1977,N_1187);
nand U2577 (N_2577,N_1993,N_316);
nand U2578 (N_2578,N_1597,N_212);
nor U2579 (N_2579,N_557,N_1460);
xor U2580 (N_2580,N_617,N_1657);
nand U2581 (N_2581,N_1897,N_272);
or U2582 (N_2582,N_548,N_784);
nor U2583 (N_2583,N_1605,N_1914);
nand U2584 (N_2584,N_736,N_1713);
xor U2585 (N_2585,N_236,N_1214);
or U2586 (N_2586,N_671,N_1535);
and U2587 (N_2587,N_1042,N_319);
nor U2588 (N_2588,N_1776,N_17);
nor U2589 (N_2589,N_1571,N_544);
nand U2590 (N_2590,N_392,N_1058);
nand U2591 (N_2591,N_253,N_492);
xor U2592 (N_2592,N_816,N_1455);
and U2593 (N_2593,N_1268,N_1078);
or U2594 (N_2594,N_179,N_1278);
nand U2595 (N_2595,N_1340,N_1097);
or U2596 (N_2596,N_1035,N_1324);
or U2597 (N_2597,N_1229,N_183);
or U2598 (N_2598,N_894,N_1739);
or U2599 (N_2599,N_811,N_1825);
and U2600 (N_2600,N_173,N_1819);
xor U2601 (N_2601,N_334,N_481);
or U2602 (N_2602,N_439,N_1531);
or U2603 (N_2603,N_1006,N_527);
nor U2604 (N_2604,N_270,N_657);
or U2605 (N_2605,N_1795,N_237);
and U2606 (N_2606,N_1826,N_141);
and U2607 (N_2607,N_508,N_745);
nand U2608 (N_2608,N_1546,N_55);
or U2609 (N_2609,N_684,N_448);
and U2610 (N_2610,N_372,N_1426);
or U2611 (N_2611,N_1823,N_915);
nor U2612 (N_2612,N_1250,N_1159);
xnor U2613 (N_2613,N_1673,N_1612);
nand U2614 (N_2614,N_101,N_723);
or U2615 (N_2615,N_1646,N_1643);
nor U2616 (N_2616,N_1020,N_1039);
and U2617 (N_2617,N_1180,N_325);
and U2618 (N_2618,N_469,N_1176);
or U2619 (N_2619,N_9,N_1910);
or U2620 (N_2620,N_852,N_108);
nor U2621 (N_2621,N_1921,N_843);
or U2622 (N_2622,N_1732,N_1992);
or U2623 (N_2623,N_647,N_1129);
and U2624 (N_2624,N_813,N_888);
nand U2625 (N_2625,N_808,N_650);
nand U2626 (N_2626,N_1223,N_478);
xnor U2627 (N_2627,N_1956,N_344);
nand U2628 (N_2628,N_1556,N_1120);
nor U2629 (N_2629,N_222,N_357);
nor U2630 (N_2630,N_1980,N_667);
nand U2631 (N_2631,N_1770,N_977);
and U2632 (N_2632,N_184,N_1868);
nor U2633 (N_2633,N_1010,N_1697);
xnor U2634 (N_2634,N_616,N_828);
nand U2635 (N_2635,N_22,N_201);
or U2636 (N_2636,N_814,N_694);
or U2637 (N_2637,N_531,N_1689);
nand U2638 (N_2638,N_770,N_1242);
or U2639 (N_2639,N_1244,N_1839);
nand U2640 (N_2640,N_1700,N_738);
and U2641 (N_2641,N_1695,N_1134);
and U2642 (N_2642,N_466,N_1175);
nand U2643 (N_2643,N_968,N_1640);
or U2644 (N_2644,N_359,N_1222);
and U2645 (N_2645,N_1963,N_274);
nor U2646 (N_2646,N_1406,N_855);
nor U2647 (N_2647,N_1297,N_765);
nor U2648 (N_2648,N_31,N_1376);
or U2649 (N_2649,N_1494,N_25);
nand U2650 (N_2650,N_367,N_789);
or U2651 (N_2651,N_990,N_1185);
nor U2652 (N_2652,N_757,N_595);
nand U2653 (N_2653,N_1321,N_233);
or U2654 (N_2654,N_458,N_1445);
nand U2655 (N_2655,N_311,N_782);
nor U2656 (N_2656,N_283,N_1292);
nand U2657 (N_2657,N_1760,N_1483);
and U2658 (N_2658,N_1997,N_80);
xnor U2659 (N_2659,N_1005,N_1481);
nand U2660 (N_2660,N_1578,N_494);
or U2661 (N_2661,N_382,N_618);
or U2662 (N_2662,N_1119,N_1865);
or U2663 (N_2663,N_1821,N_747);
nor U2664 (N_2664,N_1026,N_1813);
and U2665 (N_2665,N_1302,N_73);
or U2666 (N_2666,N_76,N_1594);
and U2667 (N_2667,N_591,N_1636);
and U2668 (N_2668,N_1609,N_1280);
nand U2669 (N_2669,N_1217,N_908);
nand U2670 (N_2670,N_421,N_143);
or U2671 (N_2671,N_1431,N_712);
nor U2672 (N_2672,N_142,N_1705);
nor U2673 (N_2673,N_1131,N_170);
nand U2674 (N_2674,N_592,N_1788);
and U2675 (N_2675,N_529,N_643);
or U2676 (N_2676,N_1320,N_1875);
or U2677 (N_2677,N_491,N_1920);
or U2678 (N_2678,N_1068,N_256);
or U2679 (N_2679,N_1128,N_331);
nand U2680 (N_2680,N_1879,N_1632);
nor U2681 (N_2681,N_1805,N_690);
nand U2682 (N_2682,N_1871,N_336);
and U2683 (N_2683,N_1190,N_602);
nor U2684 (N_2684,N_1874,N_109);
nand U2685 (N_2685,N_608,N_418);
or U2686 (N_2686,N_1247,N_468);
nand U2687 (N_2687,N_1764,N_1593);
nand U2688 (N_2688,N_1122,N_1436);
nor U2689 (N_2689,N_377,N_1951);
nand U2690 (N_2690,N_1073,N_1031);
nand U2691 (N_2691,N_1422,N_1368);
nor U2692 (N_2692,N_832,N_1565);
xnor U2693 (N_2693,N_1918,N_896);
nor U2694 (N_2694,N_208,N_1385);
or U2695 (N_2695,N_600,N_431);
nor U2696 (N_2696,N_1287,N_1859);
and U2697 (N_2697,N_1413,N_1863);
nand U2698 (N_2698,N_1954,N_150);
nand U2699 (N_2699,N_1448,N_1092);
and U2700 (N_2700,N_1105,N_981);
and U2701 (N_2701,N_1059,N_58);
xor U2702 (N_2702,N_422,N_1099);
nor U2703 (N_2703,N_589,N_1972);
and U2704 (N_2704,N_541,N_1522);
xor U2705 (N_2705,N_1238,N_1677);
nand U2706 (N_2706,N_802,N_730);
nor U2707 (N_2707,N_1485,N_1829);
nand U2708 (N_2708,N_1044,N_717);
xnor U2709 (N_2709,N_1662,N_94);
nand U2710 (N_2710,N_1142,N_238);
xor U2711 (N_2711,N_1154,N_1649);
nor U2712 (N_2712,N_223,N_986);
or U2713 (N_2713,N_1469,N_104);
nand U2714 (N_2714,N_880,N_15);
xnor U2715 (N_2715,N_1343,N_1310);
and U2716 (N_2716,N_457,N_35);
and U2717 (N_2717,N_1281,N_1895);
nand U2718 (N_2718,N_1106,N_1009);
nand U2719 (N_2719,N_1523,N_1386);
and U2720 (N_2720,N_919,N_454);
and U2721 (N_2721,N_728,N_774);
and U2722 (N_2722,N_293,N_1396);
or U2723 (N_2723,N_502,N_18);
xor U2724 (N_2724,N_895,N_1768);
and U2725 (N_2725,N_1125,N_1293);
nand U2726 (N_2726,N_638,N_398);
xnor U2727 (N_2727,N_1200,N_566);
or U2728 (N_2728,N_1712,N_1028);
and U2729 (N_2729,N_973,N_1211);
or U2730 (N_2730,N_495,N_1206);
or U2731 (N_2731,N_1309,N_1488);
nor U2732 (N_2732,N_294,N_585);
xnor U2733 (N_2733,N_1766,N_1241);
nor U2734 (N_2734,N_960,N_702);
nor U2735 (N_2735,N_246,N_778);
nor U2736 (N_2736,N_1344,N_443);
or U2737 (N_2737,N_383,N_74);
and U2738 (N_2738,N_937,N_1365);
or U2739 (N_2739,N_1912,N_1536);
and U2740 (N_2740,N_697,N_1554);
or U2741 (N_2741,N_525,N_1925);
nor U2742 (N_2742,N_1683,N_1745);
xnor U2743 (N_2743,N_98,N_1477);
or U2744 (N_2744,N_563,N_1498);
or U2745 (N_2745,N_950,N_521);
xnor U2746 (N_2746,N_727,N_530);
or U2747 (N_2747,N_1659,N_46);
or U2748 (N_2748,N_1658,N_1837);
xnor U2749 (N_2749,N_818,N_1226);
nor U2750 (N_2750,N_807,N_42);
xnor U2751 (N_2751,N_653,N_731);
nor U2752 (N_2752,N_21,N_1449);
and U2753 (N_2753,N_1627,N_1887);
and U2754 (N_2754,N_1990,N_887);
nand U2755 (N_2755,N_250,N_499);
nor U2756 (N_2756,N_1264,N_1369);
nand U2757 (N_2757,N_463,N_1451);
nand U2758 (N_2758,N_360,N_1669);
nor U2759 (N_2759,N_88,N_693);
or U2760 (N_2760,N_781,N_533);
nor U2761 (N_2761,N_719,N_1810);
nand U2762 (N_2762,N_857,N_1027);
and U2763 (N_2763,N_452,N_1359);
nand U2764 (N_2764,N_291,N_893);
or U2765 (N_2765,N_1982,N_1112);
nor U2766 (N_2766,N_1915,N_264);
or U2767 (N_2767,N_378,N_1931);
nor U2768 (N_2768,N_1366,N_1402);
nand U2769 (N_2769,N_456,N_661);
and U2770 (N_2770,N_1288,N_442);
nand U2771 (N_2771,N_780,N_555);
or U2772 (N_2772,N_107,N_1391);
and U2773 (N_2773,N_752,N_61);
nor U2774 (N_2774,N_1524,N_1228);
and U2775 (N_2775,N_1987,N_714);
nor U2776 (N_2776,N_483,N_962);
nand U2777 (N_2777,N_626,N_1100);
nand U2778 (N_2778,N_416,N_1559);
nor U2779 (N_2779,N_1945,N_988);
or U2780 (N_2780,N_1946,N_1148);
xor U2781 (N_2781,N_506,N_1543);
nand U2782 (N_2782,N_1762,N_1399);
and U2783 (N_2783,N_1975,N_865);
nand U2784 (N_2784,N_987,N_1736);
and U2785 (N_2785,N_662,N_1189);
nand U2786 (N_2786,N_1043,N_119);
nor U2787 (N_2787,N_1520,N_1251);
or U2788 (N_2788,N_1807,N_1666);
nand U2789 (N_2789,N_1063,N_1248);
nor U2790 (N_2790,N_945,N_1446);
nor U2791 (N_2791,N_965,N_944);
and U2792 (N_2792,N_1074,N_1461);
or U2793 (N_2793,N_82,N_922);
and U2794 (N_2794,N_1525,N_790);
and U2795 (N_2795,N_724,N_235);
nand U2796 (N_2796,N_829,N_132);
xnor U2797 (N_2797,N_772,N_1576);
and U2798 (N_2798,N_370,N_1236);
or U2799 (N_2799,N_924,N_868);
or U2800 (N_2800,N_1800,N_390);
or U2801 (N_2801,N_78,N_1260);
and U2802 (N_2802,N_1955,N_1978);
nand U2803 (N_2803,N_1618,N_1619);
or U2804 (N_2804,N_470,N_959);
nand U2805 (N_2805,N_785,N_713);
or U2806 (N_2806,N_480,N_798);
nand U2807 (N_2807,N_994,N_1939);
nor U2808 (N_2808,N_393,N_1008);
or U2809 (N_2809,N_249,N_863);
nor U2810 (N_2810,N_1890,N_686);
nand U2811 (N_2811,N_1742,N_1506);
nor U2812 (N_2812,N_1958,N_230);
xor U2813 (N_2813,N_1289,N_648);
or U2814 (N_2814,N_206,N_729);
and U2815 (N_2815,N_1497,N_902);
nand U2816 (N_2816,N_1457,N_1744);
or U2817 (N_2817,N_1349,N_482);
and U2818 (N_2818,N_1053,N_1723);
or U2819 (N_2819,N_1169,N_167);
or U2820 (N_2820,N_838,N_305);
nor U2821 (N_2821,N_1227,N_146);
and U2822 (N_2822,N_759,N_992);
nand U2823 (N_2823,N_1678,N_225);
nand U2824 (N_2824,N_979,N_1384);
nand U2825 (N_2825,N_56,N_1168);
nand U2826 (N_2826,N_1347,N_1007);
and U2827 (N_2827,N_1900,N_1991);
or U2828 (N_2828,N_1435,N_942);
nor U2829 (N_2829,N_621,N_1720);
nand U2830 (N_2830,N_1087,N_1983);
xor U2831 (N_2831,N_227,N_90);
nor U2832 (N_2832,N_948,N_870);
and U2833 (N_2833,N_160,N_128);
and U2834 (N_2834,N_8,N_1733);
nand U2835 (N_2835,N_333,N_38);
and U2836 (N_2836,N_1140,N_632);
xor U2837 (N_2837,N_1790,N_453);
nor U2838 (N_2838,N_1842,N_573);
or U2839 (N_2839,N_1548,N_1049);
or U2840 (N_2840,N_546,N_1486);
nand U2841 (N_2841,N_1118,N_321);
or U2842 (N_2842,N_309,N_287);
nand U2843 (N_2843,N_1334,N_1205);
nand U2844 (N_2844,N_490,N_40);
and U2845 (N_2845,N_518,N_515);
nand U2846 (N_2846,N_1171,N_1613);
nor U2847 (N_2847,N_1561,N_748);
nand U2848 (N_2848,N_1867,N_437);
nor U2849 (N_2849,N_1464,N_846);
or U2850 (N_2850,N_1941,N_39);
nor U2851 (N_2851,N_204,N_324);
or U2852 (N_2852,N_537,N_1239);
nand U2853 (N_2853,N_1566,N_323);
nor U2854 (N_2854,N_99,N_1069);
or U2855 (N_2855,N_26,N_704);
and U2856 (N_2856,N_234,N_503);
nor U2857 (N_2857,N_1401,N_1262);
nor U2858 (N_2858,N_976,N_245);
xor U2859 (N_2859,N_14,N_1751);
nand U2860 (N_2860,N_276,N_1313);
nand U2861 (N_2861,N_866,N_993);
or U2862 (N_2862,N_594,N_292);
or U2863 (N_2863,N_380,N_1179);
nand U2864 (N_2864,N_633,N_1201);
nor U2865 (N_2865,N_77,N_1884);
nand U2866 (N_2866,N_157,N_411);
nor U2867 (N_2867,N_623,N_779);
nor U2868 (N_2868,N_1032,N_1923);
xnor U2869 (N_2869,N_409,N_1741);
or U2870 (N_2870,N_1747,N_1986);
xor U2871 (N_2871,N_81,N_1072);
and U2872 (N_2872,N_1902,N_830);
or U2873 (N_2873,N_1765,N_251);
nand U2874 (N_2874,N_1691,N_910);
nor U2875 (N_2875,N_967,N_797);
and U2876 (N_2876,N_115,N_1103);
nor U2877 (N_2877,N_972,N_1411);
nand U2878 (N_2878,N_1404,N_1196);
nor U2879 (N_2879,N_1301,N_1731);
nand U2880 (N_2880,N_162,N_768);
or U2881 (N_2881,N_1350,N_1025);
and U2882 (N_2882,N_1193,N_1151);
nand U2883 (N_2883,N_692,N_1204);
and U2884 (N_2884,N_796,N_1113);
nor U2885 (N_2885,N_1245,N_1541);
or U2886 (N_2886,N_679,N_849);
xnor U2887 (N_2887,N_1763,N_1530);
nand U2888 (N_2888,N_1418,N_876);
nand U2889 (N_2889,N_864,N_1240);
nor U2890 (N_2890,N_1160,N_1419);
and U2891 (N_2891,N_1703,N_1570);
xnor U2892 (N_2892,N_1135,N_217);
nand U2893 (N_2893,N_1456,N_352);
nor U2894 (N_2894,N_1604,N_607);
nor U2895 (N_2895,N_1648,N_505);
nor U2896 (N_2896,N_152,N_477);
and U2897 (N_2897,N_583,N_346);
nor U2898 (N_2898,N_1780,N_401);
or U2899 (N_2899,N_1818,N_921);
nor U2900 (N_2900,N_296,N_1600);
xnor U2901 (N_2901,N_1219,N_553);
nor U2902 (N_2902,N_154,N_1996);
and U2903 (N_2903,N_267,N_438);
or U2904 (N_2904,N_593,N_1482);
and U2905 (N_2905,N_859,N_1266);
or U2906 (N_2906,N_1170,N_1156);
nor U2907 (N_2907,N_1501,N_1602);
nand U2908 (N_2908,N_310,N_414);
or U2909 (N_2909,N_1806,N_1290);
nand U2910 (N_2910,N_1306,N_189);
and U2911 (N_2911,N_1940,N_1771);
nand U2912 (N_2912,N_130,N_1395);
or U2913 (N_2913,N_192,N_1155);
nor U2914 (N_2914,N_850,N_930);
nor U2915 (N_2915,N_345,N_1338);
or U2916 (N_2916,N_1231,N_947);
nor U2917 (N_2917,N_286,N_649);
nor U2918 (N_2918,N_936,N_1095);
nor U2919 (N_2919,N_1249,N_1484);
nor U2920 (N_2920,N_315,N_1675);
nand U2921 (N_2921,N_326,N_961);
nand U2922 (N_2922,N_708,N_335);
and U2923 (N_2923,N_304,N_754);
and U2924 (N_2924,N_1801,N_624);
nor U2925 (N_2925,N_899,N_459);
or U2926 (N_2926,N_1592,N_341);
nand U2927 (N_2927,N_1798,N_47);
xor U2928 (N_2928,N_562,N_1038);
nor U2929 (N_2929,N_737,N_1793);
and U2930 (N_2930,N_1750,N_174);
nand U2931 (N_2931,N_329,N_165);
xnor U2932 (N_2932,N_801,N_213);
or U2933 (N_2933,N_1261,N_426);
nor U2934 (N_2934,N_1034,N_1964);
nor U2935 (N_2935,N_444,N_1123);
xor U2936 (N_2936,N_1938,N_1417);
and U2937 (N_2937,N_1014,N_1724);
and U2938 (N_2938,N_1091,N_766);
or U2939 (N_2939,N_610,N_1439);
or U2940 (N_2940,N_1146,N_240);
and U2941 (N_2941,N_1136,N_1743);
nand U2942 (N_2942,N_432,N_601);
and U2943 (N_2943,N_27,N_574);
nand U2944 (N_2944,N_869,N_1847);
xor U2945 (N_2945,N_1948,N_247);
or U2946 (N_2946,N_1143,N_1283);
or U2947 (N_2947,N_978,N_419);
nand U2948 (N_2948,N_197,N_156);
and U2949 (N_2949,N_1254,N_446);
and U2950 (N_2950,N_1624,N_349);
nand U2951 (N_2951,N_428,N_1181);
or U2952 (N_2952,N_841,N_16);
nand U2953 (N_2953,N_1834,N_1696);
or U2954 (N_2954,N_1127,N_550);
nor U2955 (N_2955,N_980,N_791);
nand U2956 (N_2956,N_577,N_1208);
or U2957 (N_2957,N_659,N_497);
xor U2958 (N_2958,N_1299,N_1339);
nand U2959 (N_2959,N_1082,N_484);
or U2960 (N_2960,N_1089,N_1812);
or U2961 (N_2961,N_1438,N_951);
nand U2962 (N_2962,N_1480,N_471);
and U2963 (N_2963,N_1598,N_1355);
nand U2964 (N_2964,N_1545,N_844);
or U2965 (N_2965,N_259,N_1423);
xnor U2966 (N_2966,N_524,N_210);
or U2967 (N_2967,N_683,N_655);
and U2968 (N_2968,N_1934,N_1759);
nor U2969 (N_2969,N_1960,N_1577);
or U2970 (N_2970,N_427,N_1312);
or U2971 (N_2971,N_60,N_1824);
and U2972 (N_2972,N_656,N_1913);
and U2973 (N_2973,N_933,N_1070);
nor U2974 (N_2974,N_1065,N_29);
nor U2975 (N_2975,N_556,N_1634);
nand U2976 (N_2976,N_1258,N_1969);
nand U2977 (N_2977,N_1311,N_925);
or U2978 (N_2978,N_242,N_1216);
or U2979 (N_2979,N_1474,N_507);
nor U2980 (N_2980,N_243,N_1864);
and U2981 (N_2981,N_86,N_1728);
or U2982 (N_2982,N_831,N_1959);
nor U2983 (N_2983,N_1512,N_540);
nor U2984 (N_2984,N_1786,N_365);
or U2985 (N_2985,N_1908,N_803);
or U2986 (N_2986,N_1672,N_983);
nor U2987 (N_2987,N_386,N_680);
nor U2988 (N_2988,N_750,N_1656);
and U2989 (N_2989,N_112,N_1644);
or U2990 (N_2990,N_1479,N_1711);
and U2991 (N_2991,N_433,N_1532);
and U2992 (N_2992,N_0,N_472);
or U2993 (N_2993,N_1667,N_1126);
xnor U2994 (N_2994,N_172,N_106);
nand U2995 (N_2995,N_652,N_1881);
nand U2996 (N_2996,N_1279,N_449);
or U2997 (N_2997,N_100,N_1974);
nor U2998 (N_2998,N_450,N_1358);
nor U2999 (N_2999,N_928,N_847);
nor U3000 (N_3000,N_1956,N_650);
nor U3001 (N_3001,N_754,N_1576);
and U3002 (N_3002,N_1873,N_160);
xnor U3003 (N_3003,N_503,N_1610);
nand U3004 (N_3004,N_1119,N_1980);
xnor U3005 (N_3005,N_1761,N_861);
nor U3006 (N_3006,N_1926,N_1364);
or U3007 (N_3007,N_1229,N_911);
or U3008 (N_3008,N_1123,N_912);
nor U3009 (N_3009,N_1377,N_428);
nand U3010 (N_3010,N_1996,N_1018);
xnor U3011 (N_3011,N_148,N_1152);
xnor U3012 (N_3012,N_1136,N_962);
nor U3013 (N_3013,N_1360,N_529);
or U3014 (N_3014,N_1783,N_971);
nand U3015 (N_3015,N_1027,N_154);
nor U3016 (N_3016,N_553,N_1735);
nor U3017 (N_3017,N_721,N_1505);
nor U3018 (N_3018,N_856,N_310);
nand U3019 (N_3019,N_436,N_1116);
nor U3020 (N_3020,N_1209,N_1116);
nand U3021 (N_3021,N_1544,N_865);
or U3022 (N_3022,N_1547,N_732);
and U3023 (N_3023,N_1411,N_611);
or U3024 (N_3024,N_432,N_72);
nand U3025 (N_3025,N_1647,N_1011);
xnor U3026 (N_3026,N_1861,N_679);
or U3027 (N_3027,N_685,N_869);
and U3028 (N_3028,N_302,N_314);
and U3029 (N_3029,N_839,N_1803);
nand U3030 (N_3030,N_1693,N_1767);
nand U3031 (N_3031,N_408,N_845);
nor U3032 (N_3032,N_1609,N_255);
or U3033 (N_3033,N_1665,N_1294);
nand U3034 (N_3034,N_429,N_1686);
or U3035 (N_3035,N_1809,N_428);
and U3036 (N_3036,N_1520,N_538);
or U3037 (N_3037,N_204,N_425);
nor U3038 (N_3038,N_1324,N_631);
nor U3039 (N_3039,N_1124,N_1766);
nand U3040 (N_3040,N_174,N_1914);
and U3041 (N_3041,N_565,N_184);
or U3042 (N_3042,N_312,N_1951);
nor U3043 (N_3043,N_1743,N_1503);
and U3044 (N_3044,N_1603,N_391);
xor U3045 (N_3045,N_542,N_1168);
xor U3046 (N_3046,N_1971,N_361);
and U3047 (N_3047,N_1618,N_1034);
xor U3048 (N_3048,N_765,N_346);
and U3049 (N_3049,N_1265,N_1811);
nand U3050 (N_3050,N_1187,N_1821);
nand U3051 (N_3051,N_873,N_503);
nand U3052 (N_3052,N_864,N_399);
and U3053 (N_3053,N_934,N_787);
nor U3054 (N_3054,N_1855,N_1165);
nand U3055 (N_3055,N_1440,N_581);
and U3056 (N_3056,N_939,N_1318);
nor U3057 (N_3057,N_129,N_1645);
or U3058 (N_3058,N_1777,N_1066);
or U3059 (N_3059,N_304,N_457);
or U3060 (N_3060,N_1336,N_1509);
and U3061 (N_3061,N_639,N_121);
xor U3062 (N_3062,N_504,N_1242);
nand U3063 (N_3063,N_495,N_407);
nand U3064 (N_3064,N_1092,N_1275);
and U3065 (N_3065,N_607,N_19);
nor U3066 (N_3066,N_1087,N_1192);
nor U3067 (N_3067,N_314,N_1097);
or U3068 (N_3068,N_1087,N_117);
and U3069 (N_3069,N_291,N_1107);
and U3070 (N_3070,N_1134,N_1273);
nand U3071 (N_3071,N_1870,N_743);
or U3072 (N_3072,N_754,N_1653);
nand U3073 (N_3073,N_885,N_1732);
nor U3074 (N_3074,N_538,N_286);
and U3075 (N_3075,N_246,N_1042);
or U3076 (N_3076,N_1625,N_581);
nor U3077 (N_3077,N_267,N_301);
or U3078 (N_3078,N_1229,N_1408);
nand U3079 (N_3079,N_906,N_1484);
nor U3080 (N_3080,N_1301,N_1746);
or U3081 (N_3081,N_911,N_615);
nor U3082 (N_3082,N_529,N_904);
xnor U3083 (N_3083,N_815,N_1111);
or U3084 (N_3084,N_23,N_1377);
or U3085 (N_3085,N_319,N_69);
and U3086 (N_3086,N_771,N_1895);
or U3087 (N_3087,N_520,N_1367);
and U3088 (N_3088,N_931,N_1239);
and U3089 (N_3089,N_442,N_1967);
xor U3090 (N_3090,N_1942,N_1021);
nor U3091 (N_3091,N_1029,N_362);
nor U3092 (N_3092,N_1674,N_1133);
nor U3093 (N_3093,N_1684,N_748);
nor U3094 (N_3094,N_1160,N_1286);
nor U3095 (N_3095,N_944,N_1570);
nand U3096 (N_3096,N_276,N_295);
nand U3097 (N_3097,N_760,N_1148);
or U3098 (N_3098,N_872,N_551);
and U3099 (N_3099,N_885,N_788);
or U3100 (N_3100,N_227,N_1940);
and U3101 (N_3101,N_1148,N_1096);
nand U3102 (N_3102,N_1448,N_349);
or U3103 (N_3103,N_85,N_369);
nand U3104 (N_3104,N_852,N_5);
and U3105 (N_3105,N_1920,N_509);
nand U3106 (N_3106,N_1981,N_1285);
nand U3107 (N_3107,N_912,N_1202);
nand U3108 (N_3108,N_746,N_492);
nand U3109 (N_3109,N_1039,N_739);
nand U3110 (N_3110,N_1561,N_583);
and U3111 (N_3111,N_1934,N_1343);
or U3112 (N_3112,N_102,N_247);
or U3113 (N_3113,N_638,N_752);
or U3114 (N_3114,N_552,N_1033);
nor U3115 (N_3115,N_282,N_110);
xor U3116 (N_3116,N_1394,N_1913);
and U3117 (N_3117,N_1269,N_1313);
and U3118 (N_3118,N_1979,N_1433);
or U3119 (N_3119,N_916,N_778);
or U3120 (N_3120,N_1503,N_1767);
xor U3121 (N_3121,N_77,N_769);
nand U3122 (N_3122,N_1675,N_739);
nor U3123 (N_3123,N_507,N_1090);
and U3124 (N_3124,N_1919,N_1227);
or U3125 (N_3125,N_1083,N_1682);
or U3126 (N_3126,N_763,N_943);
and U3127 (N_3127,N_403,N_1075);
nand U3128 (N_3128,N_1182,N_1941);
nand U3129 (N_3129,N_1449,N_1174);
or U3130 (N_3130,N_1702,N_1327);
nand U3131 (N_3131,N_1218,N_1450);
nand U3132 (N_3132,N_628,N_299);
nand U3133 (N_3133,N_1594,N_673);
or U3134 (N_3134,N_1945,N_246);
nor U3135 (N_3135,N_5,N_1662);
nor U3136 (N_3136,N_1415,N_988);
nand U3137 (N_3137,N_772,N_1044);
nor U3138 (N_3138,N_1883,N_381);
nor U3139 (N_3139,N_158,N_1853);
nand U3140 (N_3140,N_305,N_142);
xor U3141 (N_3141,N_250,N_52);
or U3142 (N_3142,N_1637,N_1706);
nor U3143 (N_3143,N_1615,N_488);
xor U3144 (N_3144,N_1105,N_626);
nand U3145 (N_3145,N_1295,N_851);
or U3146 (N_3146,N_968,N_1028);
nor U3147 (N_3147,N_220,N_1202);
nand U3148 (N_3148,N_543,N_897);
xnor U3149 (N_3149,N_1953,N_1008);
nand U3150 (N_3150,N_293,N_1403);
and U3151 (N_3151,N_149,N_1472);
or U3152 (N_3152,N_960,N_529);
and U3153 (N_3153,N_1645,N_1684);
or U3154 (N_3154,N_1513,N_1139);
or U3155 (N_3155,N_1240,N_67);
nand U3156 (N_3156,N_617,N_1046);
nor U3157 (N_3157,N_1233,N_27);
nand U3158 (N_3158,N_1948,N_1302);
nor U3159 (N_3159,N_1174,N_1705);
nand U3160 (N_3160,N_380,N_7);
nor U3161 (N_3161,N_1875,N_1656);
nor U3162 (N_3162,N_10,N_1200);
nand U3163 (N_3163,N_1357,N_1867);
or U3164 (N_3164,N_1224,N_1887);
or U3165 (N_3165,N_258,N_1408);
and U3166 (N_3166,N_172,N_1106);
or U3167 (N_3167,N_1027,N_1387);
nand U3168 (N_3168,N_193,N_108);
or U3169 (N_3169,N_897,N_1063);
nor U3170 (N_3170,N_1818,N_74);
nor U3171 (N_3171,N_528,N_1756);
and U3172 (N_3172,N_1570,N_156);
and U3173 (N_3173,N_1458,N_1066);
or U3174 (N_3174,N_939,N_1347);
nand U3175 (N_3175,N_470,N_1767);
and U3176 (N_3176,N_125,N_1097);
and U3177 (N_3177,N_492,N_1061);
xnor U3178 (N_3178,N_663,N_1683);
xor U3179 (N_3179,N_269,N_923);
or U3180 (N_3180,N_176,N_1271);
xor U3181 (N_3181,N_231,N_483);
and U3182 (N_3182,N_451,N_1270);
xor U3183 (N_3183,N_1638,N_393);
nor U3184 (N_3184,N_426,N_428);
xnor U3185 (N_3185,N_629,N_1339);
or U3186 (N_3186,N_1990,N_1082);
nor U3187 (N_3187,N_529,N_730);
nand U3188 (N_3188,N_1701,N_790);
xnor U3189 (N_3189,N_1724,N_1598);
nand U3190 (N_3190,N_1985,N_1997);
nand U3191 (N_3191,N_1803,N_1992);
and U3192 (N_3192,N_951,N_1656);
or U3193 (N_3193,N_1541,N_956);
or U3194 (N_3194,N_1512,N_1708);
nand U3195 (N_3195,N_1772,N_1196);
or U3196 (N_3196,N_1497,N_456);
or U3197 (N_3197,N_755,N_1497);
nand U3198 (N_3198,N_958,N_858);
nand U3199 (N_3199,N_595,N_862);
or U3200 (N_3200,N_698,N_796);
and U3201 (N_3201,N_837,N_75);
nor U3202 (N_3202,N_753,N_71);
nand U3203 (N_3203,N_930,N_1019);
and U3204 (N_3204,N_592,N_1970);
nand U3205 (N_3205,N_53,N_1197);
xor U3206 (N_3206,N_1938,N_1157);
nand U3207 (N_3207,N_1588,N_872);
or U3208 (N_3208,N_925,N_1650);
nand U3209 (N_3209,N_1542,N_1797);
nor U3210 (N_3210,N_1465,N_557);
and U3211 (N_3211,N_428,N_803);
and U3212 (N_3212,N_501,N_1168);
and U3213 (N_3213,N_1306,N_1206);
xor U3214 (N_3214,N_1525,N_165);
xor U3215 (N_3215,N_1080,N_1459);
xnor U3216 (N_3216,N_441,N_1426);
and U3217 (N_3217,N_1419,N_1817);
and U3218 (N_3218,N_950,N_1559);
and U3219 (N_3219,N_195,N_748);
nand U3220 (N_3220,N_932,N_298);
and U3221 (N_3221,N_291,N_607);
nand U3222 (N_3222,N_929,N_558);
xnor U3223 (N_3223,N_711,N_1045);
nor U3224 (N_3224,N_541,N_1796);
and U3225 (N_3225,N_340,N_4);
xnor U3226 (N_3226,N_960,N_1881);
xnor U3227 (N_3227,N_815,N_96);
nor U3228 (N_3228,N_32,N_1456);
nand U3229 (N_3229,N_1355,N_1138);
nor U3230 (N_3230,N_1261,N_1077);
nor U3231 (N_3231,N_541,N_100);
and U3232 (N_3232,N_1788,N_24);
or U3233 (N_3233,N_778,N_169);
nand U3234 (N_3234,N_549,N_364);
nand U3235 (N_3235,N_199,N_1956);
nor U3236 (N_3236,N_260,N_1669);
nor U3237 (N_3237,N_959,N_1502);
or U3238 (N_3238,N_49,N_1777);
or U3239 (N_3239,N_127,N_393);
nor U3240 (N_3240,N_554,N_1548);
xor U3241 (N_3241,N_1172,N_1850);
xor U3242 (N_3242,N_1446,N_1497);
or U3243 (N_3243,N_632,N_1911);
and U3244 (N_3244,N_1905,N_1954);
nand U3245 (N_3245,N_1694,N_1081);
xor U3246 (N_3246,N_1291,N_1699);
or U3247 (N_3247,N_138,N_1507);
xnor U3248 (N_3248,N_950,N_1275);
or U3249 (N_3249,N_202,N_669);
nand U3250 (N_3250,N_365,N_1695);
xnor U3251 (N_3251,N_41,N_327);
and U3252 (N_3252,N_471,N_1029);
nand U3253 (N_3253,N_1559,N_254);
and U3254 (N_3254,N_1272,N_159);
nor U3255 (N_3255,N_443,N_933);
nand U3256 (N_3256,N_185,N_1181);
or U3257 (N_3257,N_1633,N_198);
nor U3258 (N_3258,N_1858,N_1343);
nand U3259 (N_3259,N_1579,N_980);
nor U3260 (N_3260,N_438,N_806);
and U3261 (N_3261,N_446,N_892);
nor U3262 (N_3262,N_536,N_294);
xnor U3263 (N_3263,N_1275,N_1229);
or U3264 (N_3264,N_1949,N_1371);
nor U3265 (N_3265,N_1773,N_1428);
nand U3266 (N_3266,N_1034,N_477);
xnor U3267 (N_3267,N_1329,N_1811);
nand U3268 (N_3268,N_647,N_1895);
xnor U3269 (N_3269,N_1613,N_925);
nor U3270 (N_3270,N_1938,N_1527);
or U3271 (N_3271,N_519,N_591);
xnor U3272 (N_3272,N_705,N_1307);
nand U3273 (N_3273,N_1275,N_237);
nand U3274 (N_3274,N_489,N_277);
nand U3275 (N_3275,N_102,N_871);
nor U3276 (N_3276,N_75,N_1476);
and U3277 (N_3277,N_1649,N_1123);
or U3278 (N_3278,N_1599,N_1802);
nand U3279 (N_3279,N_1714,N_76);
nor U3280 (N_3280,N_1764,N_998);
xor U3281 (N_3281,N_1527,N_1749);
and U3282 (N_3282,N_1178,N_520);
xnor U3283 (N_3283,N_1304,N_1369);
nand U3284 (N_3284,N_1876,N_1066);
nor U3285 (N_3285,N_1287,N_1421);
nand U3286 (N_3286,N_157,N_879);
nand U3287 (N_3287,N_791,N_1188);
and U3288 (N_3288,N_945,N_1170);
nor U3289 (N_3289,N_170,N_1);
or U3290 (N_3290,N_1492,N_270);
nand U3291 (N_3291,N_1148,N_817);
or U3292 (N_3292,N_1692,N_573);
nor U3293 (N_3293,N_1123,N_1661);
xor U3294 (N_3294,N_494,N_1116);
nand U3295 (N_3295,N_136,N_1587);
and U3296 (N_3296,N_1417,N_1947);
nor U3297 (N_3297,N_1207,N_53);
and U3298 (N_3298,N_1722,N_1253);
and U3299 (N_3299,N_715,N_1113);
nand U3300 (N_3300,N_307,N_1479);
nor U3301 (N_3301,N_1920,N_1649);
and U3302 (N_3302,N_1936,N_937);
nor U3303 (N_3303,N_132,N_1699);
nand U3304 (N_3304,N_267,N_542);
nor U3305 (N_3305,N_191,N_54);
nor U3306 (N_3306,N_1989,N_619);
and U3307 (N_3307,N_490,N_1331);
xor U3308 (N_3308,N_343,N_515);
nor U3309 (N_3309,N_1320,N_1751);
and U3310 (N_3310,N_1913,N_1764);
nor U3311 (N_3311,N_1117,N_639);
or U3312 (N_3312,N_934,N_30);
xnor U3313 (N_3313,N_965,N_315);
or U3314 (N_3314,N_1178,N_1163);
and U3315 (N_3315,N_1499,N_401);
nand U3316 (N_3316,N_1376,N_815);
nor U3317 (N_3317,N_853,N_1500);
nor U3318 (N_3318,N_1159,N_992);
and U3319 (N_3319,N_604,N_768);
nand U3320 (N_3320,N_1425,N_911);
or U3321 (N_3321,N_710,N_848);
nand U3322 (N_3322,N_515,N_663);
xnor U3323 (N_3323,N_889,N_949);
nor U3324 (N_3324,N_1854,N_1413);
or U3325 (N_3325,N_215,N_1856);
xnor U3326 (N_3326,N_20,N_200);
or U3327 (N_3327,N_1699,N_445);
nand U3328 (N_3328,N_372,N_547);
and U3329 (N_3329,N_1439,N_1735);
and U3330 (N_3330,N_336,N_199);
nand U3331 (N_3331,N_1068,N_311);
and U3332 (N_3332,N_1219,N_1102);
nor U3333 (N_3333,N_687,N_1907);
and U3334 (N_3334,N_149,N_232);
nor U3335 (N_3335,N_1660,N_1047);
and U3336 (N_3336,N_725,N_1891);
and U3337 (N_3337,N_1060,N_1499);
nor U3338 (N_3338,N_1112,N_285);
and U3339 (N_3339,N_0,N_1006);
or U3340 (N_3340,N_1956,N_1981);
nor U3341 (N_3341,N_1574,N_1211);
and U3342 (N_3342,N_727,N_1533);
and U3343 (N_3343,N_1744,N_1809);
and U3344 (N_3344,N_531,N_1404);
or U3345 (N_3345,N_1528,N_40);
nor U3346 (N_3346,N_1974,N_126);
xnor U3347 (N_3347,N_1837,N_169);
or U3348 (N_3348,N_1657,N_779);
xor U3349 (N_3349,N_1676,N_1648);
or U3350 (N_3350,N_1866,N_292);
or U3351 (N_3351,N_291,N_196);
xor U3352 (N_3352,N_1202,N_1986);
and U3353 (N_3353,N_778,N_89);
nor U3354 (N_3354,N_1947,N_1570);
and U3355 (N_3355,N_1296,N_1213);
nand U3356 (N_3356,N_1172,N_90);
or U3357 (N_3357,N_976,N_840);
xnor U3358 (N_3358,N_1784,N_668);
and U3359 (N_3359,N_1424,N_456);
nand U3360 (N_3360,N_464,N_1544);
or U3361 (N_3361,N_659,N_1491);
or U3362 (N_3362,N_1719,N_1093);
or U3363 (N_3363,N_127,N_1699);
and U3364 (N_3364,N_142,N_307);
and U3365 (N_3365,N_646,N_1392);
nor U3366 (N_3366,N_405,N_646);
or U3367 (N_3367,N_1572,N_1702);
or U3368 (N_3368,N_413,N_1198);
or U3369 (N_3369,N_1109,N_1323);
nor U3370 (N_3370,N_1204,N_1870);
and U3371 (N_3371,N_316,N_716);
and U3372 (N_3372,N_1288,N_592);
nand U3373 (N_3373,N_608,N_151);
nand U3374 (N_3374,N_1059,N_1926);
and U3375 (N_3375,N_20,N_514);
or U3376 (N_3376,N_346,N_1155);
nor U3377 (N_3377,N_1189,N_756);
and U3378 (N_3378,N_1180,N_619);
nor U3379 (N_3379,N_440,N_837);
and U3380 (N_3380,N_1459,N_849);
or U3381 (N_3381,N_1441,N_1938);
and U3382 (N_3382,N_874,N_620);
nor U3383 (N_3383,N_889,N_1578);
nand U3384 (N_3384,N_447,N_298);
nor U3385 (N_3385,N_219,N_424);
or U3386 (N_3386,N_1572,N_848);
nand U3387 (N_3387,N_480,N_189);
nor U3388 (N_3388,N_776,N_1557);
and U3389 (N_3389,N_491,N_1308);
and U3390 (N_3390,N_1559,N_1535);
or U3391 (N_3391,N_1656,N_1413);
and U3392 (N_3392,N_1286,N_1623);
and U3393 (N_3393,N_365,N_28);
nor U3394 (N_3394,N_1478,N_367);
nand U3395 (N_3395,N_150,N_612);
and U3396 (N_3396,N_1850,N_1449);
nor U3397 (N_3397,N_978,N_662);
or U3398 (N_3398,N_401,N_1755);
and U3399 (N_3399,N_269,N_670);
nand U3400 (N_3400,N_1706,N_1374);
and U3401 (N_3401,N_97,N_837);
and U3402 (N_3402,N_314,N_789);
or U3403 (N_3403,N_507,N_441);
or U3404 (N_3404,N_317,N_557);
and U3405 (N_3405,N_1803,N_1048);
or U3406 (N_3406,N_1760,N_749);
xnor U3407 (N_3407,N_1287,N_1120);
nand U3408 (N_3408,N_564,N_1472);
and U3409 (N_3409,N_883,N_1602);
and U3410 (N_3410,N_1920,N_588);
nor U3411 (N_3411,N_1869,N_341);
or U3412 (N_3412,N_823,N_963);
xnor U3413 (N_3413,N_346,N_260);
nand U3414 (N_3414,N_1716,N_1976);
or U3415 (N_3415,N_1197,N_1938);
or U3416 (N_3416,N_48,N_197);
xor U3417 (N_3417,N_1298,N_1804);
or U3418 (N_3418,N_1341,N_1089);
and U3419 (N_3419,N_683,N_1876);
or U3420 (N_3420,N_1678,N_1829);
or U3421 (N_3421,N_1834,N_1564);
or U3422 (N_3422,N_1169,N_1943);
and U3423 (N_3423,N_1835,N_538);
nand U3424 (N_3424,N_726,N_603);
and U3425 (N_3425,N_288,N_1976);
or U3426 (N_3426,N_1624,N_1735);
and U3427 (N_3427,N_1287,N_1226);
and U3428 (N_3428,N_1165,N_1285);
and U3429 (N_3429,N_1633,N_1507);
nand U3430 (N_3430,N_1551,N_1916);
and U3431 (N_3431,N_1080,N_1616);
nor U3432 (N_3432,N_374,N_1232);
or U3433 (N_3433,N_890,N_225);
nand U3434 (N_3434,N_1254,N_270);
xor U3435 (N_3435,N_1982,N_1116);
nand U3436 (N_3436,N_298,N_1956);
xnor U3437 (N_3437,N_51,N_593);
nor U3438 (N_3438,N_1706,N_62);
nor U3439 (N_3439,N_698,N_598);
and U3440 (N_3440,N_363,N_1400);
or U3441 (N_3441,N_1842,N_1864);
and U3442 (N_3442,N_1323,N_1365);
nor U3443 (N_3443,N_32,N_751);
nor U3444 (N_3444,N_953,N_1732);
and U3445 (N_3445,N_1396,N_1769);
nand U3446 (N_3446,N_1946,N_1679);
xor U3447 (N_3447,N_68,N_1172);
nand U3448 (N_3448,N_524,N_822);
nand U3449 (N_3449,N_514,N_921);
or U3450 (N_3450,N_1136,N_550);
nor U3451 (N_3451,N_553,N_1321);
or U3452 (N_3452,N_1237,N_419);
xnor U3453 (N_3453,N_1983,N_181);
nor U3454 (N_3454,N_899,N_1139);
or U3455 (N_3455,N_1255,N_566);
or U3456 (N_3456,N_966,N_1004);
and U3457 (N_3457,N_1212,N_1766);
or U3458 (N_3458,N_1033,N_1227);
nand U3459 (N_3459,N_1981,N_1554);
nor U3460 (N_3460,N_326,N_1308);
or U3461 (N_3461,N_1247,N_1379);
or U3462 (N_3462,N_316,N_139);
xor U3463 (N_3463,N_847,N_1737);
or U3464 (N_3464,N_449,N_984);
or U3465 (N_3465,N_776,N_321);
nand U3466 (N_3466,N_1142,N_360);
and U3467 (N_3467,N_687,N_1663);
and U3468 (N_3468,N_188,N_365);
xnor U3469 (N_3469,N_1597,N_1003);
nor U3470 (N_3470,N_3,N_468);
nor U3471 (N_3471,N_1073,N_1660);
nand U3472 (N_3472,N_540,N_1660);
and U3473 (N_3473,N_1927,N_507);
nor U3474 (N_3474,N_67,N_479);
nand U3475 (N_3475,N_866,N_956);
or U3476 (N_3476,N_619,N_1074);
or U3477 (N_3477,N_1274,N_363);
and U3478 (N_3478,N_1737,N_1988);
nand U3479 (N_3479,N_460,N_1234);
xor U3480 (N_3480,N_1502,N_275);
and U3481 (N_3481,N_1140,N_1566);
nor U3482 (N_3482,N_46,N_1835);
nor U3483 (N_3483,N_593,N_1271);
and U3484 (N_3484,N_1945,N_1630);
and U3485 (N_3485,N_656,N_819);
and U3486 (N_3486,N_1818,N_537);
and U3487 (N_3487,N_1656,N_1692);
or U3488 (N_3488,N_652,N_1251);
nor U3489 (N_3489,N_510,N_1593);
nand U3490 (N_3490,N_1962,N_754);
nand U3491 (N_3491,N_807,N_920);
nor U3492 (N_3492,N_347,N_1548);
nand U3493 (N_3493,N_96,N_1027);
nand U3494 (N_3494,N_1029,N_563);
nand U3495 (N_3495,N_1668,N_821);
and U3496 (N_3496,N_1806,N_1312);
or U3497 (N_3497,N_739,N_481);
nor U3498 (N_3498,N_1251,N_177);
xor U3499 (N_3499,N_1517,N_786);
or U3500 (N_3500,N_266,N_1544);
nor U3501 (N_3501,N_1590,N_1759);
nor U3502 (N_3502,N_1753,N_446);
and U3503 (N_3503,N_1768,N_1071);
xnor U3504 (N_3504,N_382,N_1964);
or U3505 (N_3505,N_1273,N_1952);
xor U3506 (N_3506,N_1389,N_1370);
and U3507 (N_3507,N_175,N_1021);
and U3508 (N_3508,N_1433,N_880);
or U3509 (N_3509,N_358,N_1537);
nor U3510 (N_3510,N_443,N_1845);
or U3511 (N_3511,N_95,N_459);
nand U3512 (N_3512,N_181,N_1325);
or U3513 (N_3513,N_1995,N_404);
nand U3514 (N_3514,N_1156,N_205);
or U3515 (N_3515,N_1102,N_1326);
nand U3516 (N_3516,N_1719,N_812);
nand U3517 (N_3517,N_1311,N_302);
or U3518 (N_3518,N_1033,N_399);
nor U3519 (N_3519,N_234,N_212);
nand U3520 (N_3520,N_1884,N_1529);
and U3521 (N_3521,N_1700,N_281);
nand U3522 (N_3522,N_354,N_1174);
and U3523 (N_3523,N_53,N_1869);
and U3524 (N_3524,N_1794,N_503);
nor U3525 (N_3525,N_381,N_1718);
nand U3526 (N_3526,N_1735,N_110);
nor U3527 (N_3527,N_1550,N_1283);
nor U3528 (N_3528,N_885,N_1865);
or U3529 (N_3529,N_798,N_32);
or U3530 (N_3530,N_1157,N_1773);
nor U3531 (N_3531,N_919,N_42);
nand U3532 (N_3532,N_1904,N_55);
xor U3533 (N_3533,N_1669,N_739);
and U3534 (N_3534,N_1215,N_1298);
or U3535 (N_3535,N_1300,N_42);
nor U3536 (N_3536,N_1898,N_1584);
nor U3537 (N_3537,N_413,N_976);
and U3538 (N_3538,N_152,N_643);
or U3539 (N_3539,N_953,N_902);
and U3540 (N_3540,N_1289,N_1414);
nor U3541 (N_3541,N_1042,N_1283);
nor U3542 (N_3542,N_1699,N_1975);
xor U3543 (N_3543,N_384,N_1215);
nand U3544 (N_3544,N_936,N_447);
nor U3545 (N_3545,N_142,N_733);
or U3546 (N_3546,N_797,N_752);
and U3547 (N_3547,N_94,N_746);
and U3548 (N_3548,N_196,N_1674);
and U3549 (N_3549,N_1778,N_777);
nor U3550 (N_3550,N_812,N_1761);
nand U3551 (N_3551,N_18,N_1331);
nand U3552 (N_3552,N_787,N_1815);
nand U3553 (N_3553,N_561,N_606);
or U3554 (N_3554,N_1559,N_1988);
and U3555 (N_3555,N_1968,N_675);
nand U3556 (N_3556,N_785,N_191);
and U3557 (N_3557,N_627,N_322);
xnor U3558 (N_3558,N_1123,N_754);
nor U3559 (N_3559,N_972,N_458);
nor U3560 (N_3560,N_1432,N_1404);
or U3561 (N_3561,N_1209,N_191);
nor U3562 (N_3562,N_773,N_100);
or U3563 (N_3563,N_1740,N_1498);
nor U3564 (N_3564,N_647,N_1751);
and U3565 (N_3565,N_268,N_1202);
or U3566 (N_3566,N_1115,N_56);
or U3567 (N_3567,N_1524,N_933);
or U3568 (N_3568,N_261,N_1459);
xor U3569 (N_3569,N_212,N_1967);
and U3570 (N_3570,N_1524,N_1075);
nor U3571 (N_3571,N_1260,N_1229);
or U3572 (N_3572,N_32,N_349);
xnor U3573 (N_3573,N_978,N_1747);
and U3574 (N_3574,N_1086,N_1787);
and U3575 (N_3575,N_1617,N_1512);
nor U3576 (N_3576,N_1857,N_1710);
or U3577 (N_3577,N_1550,N_142);
xor U3578 (N_3578,N_1826,N_1318);
or U3579 (N_3579,N_173,N_953);
nand U3580 (N_3580,N_328,N_1561);
nand U3581 (N_3581,N_1508,N_515);
nor U3582 (N_3582,N_126,N_1464);
and U3583 (N_3583,N_1865,N_1279);
and U3584 (N_3584,N_1468,N_48);
nor U3585 (N_3585,N_1651,N_1035);
nand U3586 (N_3586,N_874,N_1262);
nor U3587 (N_3587,N_1430,N_1334);
nor U3588 (N_3588,N_1748,N_1450);
nor U3589 (N_3589,N_1038,N_953);
nor U3590 (N_3590,N_204,N_1237);
and U3591 (N_3591,N_524,N_1077);
nand U3592 (N_3592,N_466,N_1368);
or U3593 (N_3593,N_1779,N_262);
and U3594 (N_3594,N_1329,N_1814);
nor U3595 (N_3595,N_152,N_1269);
or U3596 (N_3596,N_1892,N_1430);
nand U3597 (N_3597,N_526,N_1822);
nand U3598 (N_3598,N_1121,N_945);
xor U3599 (N_3599,N_966,N_191);
nor U3600 (N_3600,N_141,N_795);
and U3601 (N_3601,N_299,N_1925);
and U3602 (N_3602,N_1641,N_38);
or U3603 (N_3603,N_1613,N_885);
or U3604 (N_3604,N_1156,N_1482);
nand U3605 (N_3605,N_1808,N_103);
nand U3606 (N_3606,N_1316,N_1573);
and U3607 (N_3607,N_1076,N_785);
and U3608 (N_3608,N_146,N_482);
or U3609 (N_3609,N_494,N_1094);
and U3610 (N_3610,N_1087,N_1282);
nand U3611 (N_3611,N_1781,N_933);
nand U3612 (N_3612,N_1209,N_1188);
nor U3613 (N_3613,N_1902,N_1463);
nand U3614 (N_3614,N_729,N_1910);
or U3615 (N_3615,N_744,N_1320);
nand U3616 (N_3616,N_1640,N_1663);
nor U3617 (N_3617,N_319,N_39);
and U3618 (N_3618,N_487,N_1166);
nand U3619 (N_3619,N_1917,N_134);
xor U3620 (N_3620,N_1402,N_388);
nand U3621 (N_3621,N_693,N_615);
or U3622 (N_3622,N_509,N_397);
xnor U3623 (N_3623,N_1875,N_1052);
nor U3624 (N_3624,N_570,N_603);
nor U3625 (N_3625,N_1382,N_1845);
and U3626 (N_3626,N_58,N_1180);
or U3627 (N_3627,N_403,N_1925);
nor U3628 (N_3628,N_1214,N_1808);
nor U3629 (N_3629,N_1364,N_1980);
nor U3630 (N_3630,N_1017,N_1464);
nor U3631 (N_3631,N_718,N_122);
nor U3632 (N_3632,N_556,N_202);
nand U3633 (N_3633,N_1730,N_1647);
and U3634 (N_3634,N_987,N_588);
and U3635 (N_3635,N_284,N_325);
xnor U3636 (N_3636,N_808,N_1568);
nor U3637 (N_3637,N_537,N_591);
nor U3638 (N_3638,N_96,N_753);
nor U3639 (N_3639,N_1591,N_1131);
nor U3640 (N_3640,N_1855,N_939);
nand U3641 (N_3641,N_1284,N_1640);
and U3642 (N_3642,N_1876,N_1690);
xnor U3643 (N_3643,N_307,N_1189);
or U3644 (N_3644,N_942,N_1850);
or U3645 (N_3645,N_447,N_899);
xor U3646 (N_3646,N_916,N_42);
or U3647 (N_3647,N_1157,N_472);
and U3648 (N_3648,N_1657,N_378);
nand U3649 (N_3649,N_1992,N_795);
nor U3650 (N_3650,N_1025,N_1227);
nor U3651 (N_3651,N_1212,N_1831);
nand U3652 (N_3652,N_1289,N_712);
nor U3653 (N_3653,N_1045,N_636);
nand U3654 (N_3654,N_1116,N_7);
or U3655 (N_3655,N_972,N_1232);
or U3656 (N_3656,N_1953,N_1974);
xor U3657 (N_3657,N_547,N_1919);
or U3658 (N_3658,N_1927,N_1484);
nor U3659 (N_3659,N_1218,N_1147);
nand U3660 (N_3660,N_1102,N_1665);
nor U3661 (N_3661,N_1152,N_1705);
or U3662 (N_3662,N_250,N_1823);
nor U3663 (N_3663,N_869,N_481);
and U3664 (N_3664,N_1385,N_251);
xor U3665 (N_3665,N_592,N_1755);
nand U3666 (N_3666,N_530,N_212);
nor U3667 (N_3667,N_1788,N_266);
nand U3668 (N_3668,N_1638,N_1647);
and U3669 (N_3669,N_719,N_1922);
or U3670 (N_3670,N_944,N_1851);
or U3671 (N_3671,N_560,N_1497);
nor U3672 (N_3672,N_1304,N_1866);
nor U3673 (N_3673,N_1343,N_608);
or U3674 (N_3674,N_1536,N_356);
or U3675 (N_3675,N_1278,N_1549);
and U3676 (N_3676,N_367,N_1598);
nor U3677 (N_3677,N_1290,N_122);
or U3678 (N_3678,N_1928,N_1324);
xnor U3679 (N_3679,N_173,N_749);
xor U3680 (N_3680,N_1355,N_1624);
xor U3681 (N_3681,N_495,N_880);
nand U3682 (N_3682,N_1296,N_475);
or U3683 (N_3683,N_723,N_1462);
or U3684 (N_3684,N_1334,N_455);
and U3685 (N_3685,N_755,N_1467);
nand U3686 (N_3686,N_708,N_1520);
or U3687 (N_3687,N_965,N_1826);
nand U3688 (N_3688,N_1938,N_1011);
or U3689 (N_3689,N_505,N_1834);
xor U3690 (N_3690,N_1487,N_1709);
xor U3691 (N_3691,N_725,N_924);
nand U3692 (N_3692,N_77,N_409);
or U3693 (N_3693,N_1968,N_66);
nand U3694 (N_3694,N_107,N_1824);
or U3695 (N_3695,N_1703,N_1496);
and U3696 (N_3696,N_1283,N_1437);
and U3697 (N_3697,N_555,N_1539);
xor U3698 (N_3698,N_969,N_1443);
nor U3699 (N_3699,N_1411,N_3);
nand U3700 (N_3700,N_379,N_1194);
nor U3701 (N_3701,N_1097,N_560);
or U3702 (N_3702,N_566,N_1086);
nand U3703 (N_3703,N_1168,N_1138);
nor U3704 (N_3704,N_305,N_1987);
nand U3705 (N_3705,N_490,N_1286);
and U3706 (N_3706,N_1862,N_778);
nand U3707 (N_3707,N_1015,N_508);
or U3708 (N_3708,N_1605,N_926);
nor U3709 (N_3709,N_540,N_1634);
or U3710 (N_3710,N_1651,N_922);
and U3711 (N_3711,N_736,N_1932);
and U3712 (N_3712,N_932,N_1556);
or U3713 (N_3713,N_1654,N_1234);
nand U3714 (N_3714,N_181,N_639);
or U3715 (N_3715,N_1874,N_636);
or U3716 (N_3716,N_321,N_1713);
or U3717 (N_3717,N_1449,N_479);
nand U3718 (N_3718,N_1163,N_166);
nor U3719 (N_3719,N_1138,N_1022);
and U3720 (N_3720,N_77,N_138);
nor U3721 (N_3721,N_824,N_686);
and U3722 (N_3722,N_106,N_1424);
and U3723 (N_3723,N_333,N_787);
or U3724 (N_3724,N_604,N_391);
nor U3725 (N_3725,N_25,N_45);
and U3726 (N_3726,N_335,N_902);
and U3727 (N_3727,N_1843,N_1603);
nor U3728 (N_3728,N_1625,N_1032);
or U3729 (N_3729,N_602,N_516);
nor U3730 (N_3730,N_1761,N_313);
nor U3731 (N_3731,N_1376,N_1665);
nor U3732 (N_3732,N_705,N_613);
nor U3733 (N_3733,N_306,N_1906);
or U3734 (N_3734,N_1007,N_1027);
nand U3735 (N_3735,N_447,N_552);
xnor U3736 (N_3736,N_188,N_1722);
or U3737 (N_3737,N_1637,N_43);
nand U3738 (N_3738,N_1275,N_1747);
and U3739 (N_3739,N_1914,N_951);
and U3740 (N_3740,N_1481,N_1477);
or U3741 (N_3741,N_581,N_352);
nand U3742 (N_3742,N_121,N_660);
or U3743 (N_3743,N_1529,N_1489);
or U3744 (N_3744,N_596,N_744);
or U3745 (N_3745,N_1698,N_549);
nand U3746 (N_3746,N_1227,N_1335);
or U3747 (N_3747,N_1334,N_1858);
nand U3748 (N_3748,N_659,N_1057);
and U3749 (N_3749,N_1593,N_738);
nor U3750 (N_3750,N_1159,N_1391);
or U3751 (N_3751,N_785,N_1638);
or U3752 (N_3752,N_1636,N_1938);
and U3753 (N_3753,N_1994,N_794);
and U3754 (N_3754,N_1621,N_1878);
and U3755 (N_3755,N_1137,N_1415);
or U3756 (N_3756,N_1876,N_769);
and U3757 (N_3757,N_152,N_972);
nand U3758 (N_3758,N_1532,N_65);
nor U3759 (N_3759,N_181,N_752);
xor U3760 (N_3760,N_844,N_1861);
nand U3761 (N_3761,N_1395,N_165);
nor U3762 (N_3762,N_1412,N_1551);
nor U3763 (N_3763,N_331,N_757);
nand U3764 (N_3764,N_224,N_1378);
and U3765 (N_3765,N_793,N_1782);
xnor U3766 (N_3766,N_1499,N_1111);
and U3767 (N_3767,N_475,N_1196);
nand U3768 (N_3768,N_553,N_115);
nand U3769 (N_3769,N_1633,N_1846);
xnor U3770 (N_3770,N_184,N_267);
or U3771 (N_3771,N_1203,N_1349);
and U3772 (N_3772,N_841,N_755);
and U3773 (N_3773,N_511,N_262);
or U3774 (N_3774,N_1946,N_1035);
nor U3775 (N_3775,N_1554,N_77);
or U3776 (N_3776,N_240,N_227);
or U3777 (N_3777,N_599,N_1585);
nand U3778 (N_3778,N_851,N_1762);
nor U3779 (N_3779,N_1375,N_1870);
and U3780 (N_3780,N_449,N_103);
xnor U3781 (N_3781,N_336,N_785);
or U3782 (N_3782,N_1315,N_878);
or U3783 (N_3783,N_270,N_892);
and U3784 (N_3784,N_1416,N_238);
or U3785 (N_3785,N_1550,N_796);
and U3786 (N_3786,N_1810,N_806);
and U3787 (N_3787,N_1330,N_1483);
xor U3788 (N_3788,N_1894,N_75);
or U3789 (N_3789,N_909,N_58);
or U3790 (N_3790,N_340,N_6);
or U3791 (N_3791,N_12,N_1551);
and U3792 (N_3792,N_870,N_320);
and U3793 (N_3793,N_400,N_1017);
or U3794 (N_3794,N_352,N_1540);
or U3795 (N_3795,N_1123,N_433);
and U3796 (N_3796,N_1915,N_369);
nand U3797 (N_3797,N_1691,N_430);
and U3798 (N_3798,N_1955,N_748);
xor U3799 (N_3799,N_1357,N_734);
and U3800 (N_3800,N_853,N_1955);
xor U3801 (N_3801,N_1695,N_510);
xnor U3802 (N_3802,N_212,N_1304);
nand U3803 (N_3803,N_944,N_1260);
or U3804 (N_3804,N_1215,N_1599);
and U3805 (N_3805,N_1915,N_605);
or U3806 (N_3806,N_1204,N_535);
nand U3807 (N_3807,N_1885,N_1284);
or U3808 (N_3808,N_1534,N_561);
and U3809 (N_3809,N_1401,N_1732);
nor U3810 (N_3810,N_1532,N_470);
nor U3811 (N_3811,N_543,N_1866);
or U3812 (N_3812,N_519,N_191);
nor U3813 (N_3813,N_1634,N_936);
xor U3814 (N_3814,N_865,N_1499);
nor U3815 (N_3815,N_1533,N_1947);
and U3816 (N_3816,N_1004,N_642);
or U3817 (N_3817,N_923,N_1953);
nor U3818 (N_3818,N_1668,N_80);
and U3819 (N_3819,N_1704,N_1766);
nor U3820 (N_3820,N_1968,N_1359);
and U3821 (N_3821,N_318,N_1138);
xor U3822 (N_3822,N_1701,N_54);
and U3823 (N_3823,N_910,N_1418);
nor U3824 (N_3824,N_1172,N_1821);
or U3825 (N_3825,N_458,N_366);
or U3826 (N_3826,N_566,N_100);
nor U3827 (N_3827,N_1912,N_1198);
or U3828 (N_3828,N_1100,N_746);
and U3829 (N_3829,N_303,N_425);
and U3830 (N_3830,N_590,N_1396);
or U3831 (N_3831,N_1757,N_975);
nor U3832 (N_3832,N_1391,N_1370);
nand U3833 (N_3833,N_428,N_59);
nor U3834 (N_3834,N_970,N_563);
xnor U3835 (N_3835,N_1164,N_562);
nand U3836 (N_3836,N_684,N_952);
or U3837 (N_3837,N_1015,N_1214);
nand U3838 (N_3838,N_323,N_1658);
nand U3839 (N_3839,N_980,N_1690);
nand U3840 (N_3840,N_1324,N_1478);
nand U3841 (N_3841,N_931,N_252);
or U3842 (N_3842,N_180,N_1314);
or U3843 (N_3843,N_1009,N_572);
and U3844 (N_3844,N_508,N_360);
nand U3845 (N_3845,N_773,N_359);
or U3846 (N_3846,N_675,N_670);
or U3847 (N_3847,N_1910,N_1227);
or U3848 (N_3848,N_101,N_14);
and U3849 (N_3849,N_548,N_167);
or U3850 (N_3850,N_397,N_357);
nor U3851 (N_3851,N_747,N_1222);
nand U3852 (N_3852,N_187,N_474);
nor U3853 (N_3853,N_627,N_1473);
nor U3854 (N_3854,N_1469,N_653);
nand U3855 (N_3855,N_1320,N_779);
xor U3856 (N_3856,N_639,N_1856);
nand U3857 (N_3857,N_1640,N_1271);
or U3858 (N_3858,N_553,N_917);
nor U3859 (N_3859,N_1776,N_1506);
and U3860 (N_3860,N_1780,N_817);
nor U3861 (N_3861,N_1606,N_341);
nor U3862 (N_3862,N_1513,N_1609);
xor U3863 (N_3863,N_62,N_1891);
nor U3864 (N_3864,N_1768,N_1167);
nor U3865 (N_3865,N_345,N_1599);
xor U3866 (N_3866,N_556,N_392);
or U3867 (N_3867,N_79,N_1288);
xor U3868 (N_3868,N_1681,N_457);
or U3869 (N_3869,N_1384,N_1040);
or U3870 (N_3870,N_954,N_925);
or U3871 (N_3871,N_61,N_96);
xnor U3872 (N_3872,N_386,N_53);
nor U3873 (N_3873,N_632,N_1269);
or U3874 (N_3874,N_364,N_1867);
nor U3875 (N_3875,N_1603,N_1461);
nand U3876 (N_3876,N_1342,N_404);
and U3877 (N_3877,N_609,N_1098);
and U3878 (N_3878,N_1847,N_665);
or U3879 (N_3879,N_1195,N_329);
and U3880 (N_3880,N_1935,N_1530);
nand U3881 (N_3881,N_1629,N_798);
nor U3882 (N_3882,N_1322,N_749);
and U3883 (N_3883,N_1621,N_775);
nor U3884 (N_3884,N_1819,N_211);
and U3885 (N_3885,N_743,N_1936);
nor U3886 (N_3886,N_1181,N_892);
or U3887 (N_3887,N_1862,N_1601);
nor U3888 (N_3888,N_368,N_839);
and U3889 (N_3889,N_1530,N_595);
or U3890 (N_3890,N_1119,N_547);
xnor U3891 (N_3891,N_497,N_908);
or U3892 (N_3892,N_467,N_633);
nand U3893 (N_3893,N_1790,N_1057);
or U3894 (N_3894,N_216,N_1207);
nor U3895 (N_3895,N_1282,N_1240);
nand U3896 (N_3896,N_421,N_1679);
nand U3897 (N_3897,N_176,N_1403);
or U3898 (N_3898,N_69,N_44);
or U3899 (N_3899,N_480,N_825);
nor U3900 (N_3900,N_349,N_1577);
nor U3901 (N_3901,N_573,N_45);
nor U3902 (N_3902,N_1626,N_1035);
or U3903 (N_3903,N_765,N_972);
nor U3904 (N_3904,N_1961,N_299);
and U3905 (N_3905,N_1856,N_1506);
and U3906 (N_3906,N_457,N_1425);
or U3907 (N_3907,N_600,N_724);
or U3908 (N_3908,N_749,N_472);
nor U3909 (N_3909,N_603,N_1746);
nand U3910 (N_3910,N_1242,N_1706);
nand U3911 (N_3911,N_1896,N_1900);
nand U3912 (N_3912,N_1094,N_199);
nor U3913 (N_3913,N_1357,N_660);
nand U3914 (N_3914,N_1345,N_1009);
nand U3915 (N_3915,N_1455,N_1750);
and U3916 (N_3916,N_648,N_616);
nand U3917 (N_3917,N_1634,N_1244);
or U3918 (N_3918,N_1801,N_1423);
nor U3919 (N_3919,N_1439,N_1322);
or U3920 (N_3920,N_1434,N_1651);
or U3921 (N_3921,N_131,N_1533);
nor U3922 (N_3922,N_37,N_570);
nor U3923 (N_3923,N_617,N_325);
nand U3924 (N_3924,N_165,N_599);
nor U3925 (N_3925,N_1646,N_9);
nor U3926 (N_3926,N_1727,N_1866);
and U3927 (N_3927,N_556,N_872);
nand U3928 (N_3928,N_264,N_1682);
and U3929 (N_3929,N_1739,N_873);
nand U3930 (N_3930,N_1741,N_1391);
nand U3931 (N_3931,N_964,N_464);
xor U3932 (N_3932,N_630,N_923);
or U3933 (N_3933,N_393,N_1623);
and U3934 (N_3934,N_1075,N_363);
nand U3935 (N_3935,N_760,N_1621);
nand U3936 (N_3936,N_1157,N_1513);
nand U3937 (N_3937,N_313,N_963);
nor U3938 (N_3938,N_1350,N_1483);
and U3939 (N_3939,N_1609,N_1691);
and U3940 (N_3940,N_819,N_619);
nor U3941 (N_3941,N_685,N_1052);
nor U3942 (N_3942,N_1878,N_260);
xnor U3943 (N_3943,N_850,N_59);
or U3944 (N_3944,N_724,N_1390);
and U3945 (N_3945,N_745,N_391);
or U3946 (N_3946,N_1498,N_14);
xor U3947 (N_3947,N_322,N_1634);
or U3948 (N_3948,N_747,N_324);
and U3949 (N_3949,N_1775,N_775);
nand U3950 (N_3950,N_1692,N_724);
nor U3951 (N_3951,N_1750,N_1640);
and U3952 (N_3952,N_506,N_508);
and U3953 (N_3953,N_110,N_539);
and U3954 (N_3954,N_1587,N_902);
and U3955 (N_3955,N_1235,N_1951);
or U3956 (N_3956,N_860,N_977);
or U3957 (N_3957,N_522,N_1700);
or U3958 (N_3958,N_340,N_76);
nor U3959 (N_3959,N_1629,N_1468);
or U3960 (N_3960,N_1312,N_1861);
xor U3961 (N_3961,N_650,N_338);
and U3962 (N_3962,N_36,N_1631);
nor U3963 (N_3963,N_114,N_1831);
or U3964 (N_3964,N_197,N_1389);
nor U3965 (N_3965,N_937,N_795);
or U3966 (N_3966,N_392,N_1502);
nand U3967 (N_3967,N_1226,N_364);
and U3968 (N_3968,N_531,N_109);
nor U3969 (N_3969,N_464,N_1538);
nand U3970 (N_3970,N_991,N_278);
and U3971 (N_3971,N_906,N_236);
nand U3972 (N_3972,N_742,N_1918);
nor U3973 (N_3973,N_864,N_235);
or U3974 (N_3974,N_1995,N_658);
nor U3975 (N_3975,N_1409,N_1719);
or U3976 (N_3976,N_291,N_732);
nor U3977 (N_3977,N_1275,N_1409);
nand U3978 (N_3978,N_1982,N_772);
or U3979 (N_3979,N_1955,N_1404);
nor U3980 (N_3980,N_633,N_1823);
and U3981 (N_3981,N_1699,N_701);
nor U3982 (N_3982,N_604,N_830);
nand U3983 (N_3983,N_431,N_1649);
xnor U3984 (N_3984,N_413,N_1721);
nor U3985 (N_3985,N_634,N_407);
and U3986 (N_3986,N_709,N_1061);
and U3987 (N_3987,N_91,N_992);
or U3988 (N_3988,N_84,N_1236);
xor U3989 (N_3989,N_748,N_566);
or U3990 (N_3990,N_249,N_1761);
and U3991 (N_3991,N_35,N_1808);
or U3992 (N_3992,N_736,N_414);
or U3993 (N_3993,N_1299,N_1362);
and U3994 (N_3994,N_833,N_682);
nor U3995 (N_3995,N_1229,N_162);
nor U3996 (N_3996,N_1352,N_492);
nand U3997 (N_3997,N_1476,N_1742);
and U3998 (N_3998,N_234,N_948);
nand U3999 (N_3999,N_1659,N_515);
nor U4000 (N_4000,N_3855,N_3733);
xor U4001 (N_4001,N_3259,N_3894);
xor U4002 (N_4002,N_3354,N_2455);
nor U4003 (N_4003,N_2874,N_2319);
and U4004 (N_4004,N_2994,N_2237);
nor U4005 (N_4005,N_2108,N_3079);
nand U4006 (N_4006,N_2304,N_3068);
and U4007 (N_4007,N_2200,N_2204);
nor U4008 (N_4008,N_2651,N_3388);
nor U4009 (N_4009,N_3747,N_3467);
or U4010 (N_4010,N_3436,N_2866);
or U4011 (N_4011,N_3590,N_3854);
nor U4012 (N_4012,N_3743,N_2184);
nand U4013 (N_4013,N_3604,N_2481);
or U4014 (N_4014,N_3153,N_3022);
nor U4015 (N_4015,N_3621,N_2381);
xnor U4016 (N_4016,N_2404,N_3111);
and U4017 (N_4017,N_2466,N_3638);
nand U4018 (N_4018,N_2389,N_2735);
or U4019 (N_4019,N_3714,N_2128);
and U4020 (N_4020,N_3701,N_3990);
or U4021 (N_4021,N_2152,N_2293);
nor U4022 (N_4022,N_2028,N_3293);
and U4023 (N_4023,N_3761,N_2654);
or U4024 (N_4024,N_3537,N_3924);
and U4025 (N_4025,N_2766,N_3702);
or U4026 (N_4026,N_3744,N_2121);
or U4027 (N_4027,N_3504,N_3502);
nand U4028 (N_4028,N_3035,N_2348);
nand U4029 (N_4029,N_3229,N_2221);
xor U4030 (N_4030,N_3023,N_3770);
and U4031 (N_4031,N_2551,N_2898);
nand U4032 (N_4032,N_3399,N_2934);
nand U4033 (N_4033,N_3807,N_3099);
nor U4034 (N_4034,N_2065,N_2828);
or U4035 (N_4035,N_2274,N_2497);
or U4036 (N_4036,N_2641,N_2194);
nand U4037 (N_4037,N_2008,N_2541);
or U4038 (N_4038,N_2837,N_3248);
and U4039 (N_4039,N_2003,N_2104);
or U4040 (N_4040,N_2281,N_2361);
xor U4041 (N_4041,N_3421,N_2212);
nor U4042 (N_4042,N_2145,N_3186);
nor U4043 (N_4043,N_3626,N_3199);
nor U4044 (N_4044,N_3599,N_3469);
and U4045 (N_4045,N_2075,N_3147);
nor U4046 (N_4046,N_3460,N_2933);
nand U4047 (N_4047,N_3908,N_3315);
or U4048 (N_4048,N_2462,N_2263);
nor U4049 (N_4049,N_3350,N_3085);
nand U4050 (N_4050,N_2567,N_3211);
nor U4051 (N_4051,N_3663,N_2329);
and U4052 (N_4052,N_3818,N_2115);
nor U4053 (N_4053,N_3528,N_2680);
and U4054 (N_4054,N_2671,N_3956);
or U4055 (N_4055,N_3535,N_2521);
nand U4056 (N_4056,N_3312,N_3672);
nand U4057 (N_4057,N_2364,N_3032);
and U4058 (N_4058,N_2538,N_3741);
and U4059 (N_4059,N_3786,N_3962);
nand U4060 (N_4060,N_3135,N_2816);
nor U4061 (N_4061,N_2313,N_3210);
or U4062 (N_4062,N_2801,N_3367);
xnor U4063 (N_4063,N_3907,N_3386);
and U4064 (N_4064,N_2725,N_2708);
and U4065 (N_4065,N_2129,N_2315);
or U4066 (N_4066,N_2949,N_2431);
and U4067 (N_4067,N_2130,N_3572);
or U4068 (N_4068,N_2970,N_3343);
or U4069 (N_4069,N_2147,N_3936);
and U4070 (N_4070,N_2211,N_3616);
nand U4071 (N_4071,N_3483,N_2048);
nor U4072 (N_4072,N_2303,N_3731);
nor U4073 (N_4073,N_3579,N_2367);
and U4074 (N_4074,N_3444,N_3014);
or U4075 (N_4075,N_3954,N_3719);
nand U4076 (N_4076,N_2001,N_3806);
or U4077 (N_4077,N_2771,N_2531);
nand U4078 (N_4078,N_2825,N_2318);
or U4079 (N_4079,N_3550,N_2167);
nand U4080 (N_4080,N_2421,N_2623);
nor U4081 (N_4081,N_2302,N_2442);
or U4082 (N_4082,N_3769,N_2457);
and U4083 (N_4083,N_2073,N_3285);
nor U4084 (N_4084,N_2287,N_2314);
or U4085 (N_4085,N_3425,N_3824);
nand U4086 (N_4086,N_3995,N_2446);
nand U4087 (N_4087,N_2209,N_2868);
nor U4088 (N_4088,N_3138,N_3008);
nand U4089 (N_4089,N_3815,N_3893);
or U4090 (N_4090,N_2344,N_2682);
nor U4091 (N_4091,N_2013,N_2330);
xnor U4092 (N_4092,N_3686,N_2443);
and U4093 (N_4093,N_2879,N_2526);
and U4094 (N_4094,N_3188,N_3557);
or U4095 (N_4095,N_2857,N_3143);
or U4096 (N_4096,N_2605,N_2203);
nand U4097 (N_4097,N_3179,N_2074);
nand U4098 (N_4098,N_3081,N_2935);
or U4099 (N_4099,N_2833,N_2743);
or U4100 (N_4100,N_2685,N_2723);
or U4101 (N_4101,N_2180,N_2175);
nand U4102 (N_4102,N_2402,N_3859);
or U4103 (N_4103,N_2757,N_3933);
nand U4104 (N_4104,N_3524,N_2620);
or U4105 (N_4105,N_3778,N_2822);
nand U4106 (N_4106,N_2405,N_3764);
and U4107 (N_4107,N_3843,N_2707);
nor U4108 (N_4108,N_3906,N_2829);
and U4109 (N_4109,N_2134,N_2997);
and U4110 (N_4110,N_3542,N_3307);
and U4111 (N_4111,N_3455,N_2440);
xnor U4112 (N_4112,N_3465,N_2226);
or U4113 (N_4113,N_3159,N_3586);
or U4114 (N_4114,N_3294,N_3250);
nor U4115 (N_4115,N_3348,N_3200);
xor U4116 (N_4116,N_3055,N_3074);
nor U4117 (N_4117,N_3495,N_2273);
and U4118 (N_4118,N_2909,N_3898);
nand U4119 (N_4119,N_2007,N_3453);
nand U4120 (N_4120,N_3264,N_2684);
xor U4121 (N_4121,N_2688,N_3998);
or U4122 (N_4122,N_2384,N_2876);
xnor U4123 (N_4123,N_2081,N_3351);
or U4124 (N_4124,N_3341,N_3570);
or U4125 (N_4125,N_2883,N_3031);
xnor U4126 (N_4126,N_2950,N_2550);
or U4127 (N_4127,N_2556,N_3493);
or U4128 (N_4128,N_3140,N_2573);
or U4129 (N_4129,N_2116,N_3652);
or U4130 (N_4130,N_3788,N_3768);
or U4131 (N_4131,N_3301,N_3739);
and U4132 (N_4132,N_3424,N_3072);
nand U4133 (N_4133,N_2610,N_3305);
or U4134 (N_4134,N_2679,N_2490);
nand U4135 (N_4135,N_2944,N_3693);
xnor U4136 (N_4136,N_2474,N_2590);
nor U4137 (N_4137,N_3271,N_3418);
nor U4138 (N_4138,N_2151,N_2247);
nand U4139 (N_4139,N_2845,N_2191);
nand U4140 (N_4140,N_2965,N_2699);
nor U4141 (N_4141,N_2911,N_2183);
xnor U4142 (N_4142,N_3345,N_2706);
and U4143 (N_4143,N_2705,N_3759);
nand U4144 (N_4144,N_2819,N_2505);
nor U4145 (N_4145,N_2905,N_2027);
or U4146 (N_4146,N_3710,N_3296);
or U4147 (N_4147,N_3848,N_3694);
and U4148 (N_4148,N_3204,N_2046);
or U4149 (N_4149,N_2842,N_3084);
nor U4150 (N_4150,N_3437,N_2818);
nand U4151 (N_4151,N_2020,N_3447);
xor U4152 (N_4152,N_2085,N_2185);
nor U4153 (N_4153,N_2892,N_2714);
or U4154 (N_4154,N_3158,N_3448);
nor U4155 (N_4155,N_3088,N_3239);
and U4156 (N_4156,N_3889,N_2710);
and U4157 (N_4157,N_2470,N_3593);
xor U4158 (N_4158,N_2327,N_3427);
nor U4159 (N_4159,N_3574,N_3949);
and U4160 (N_4160,N_3977,N_2496);
and U4161 (N_4161,N_3000,N_2830);
nand U4162 (N_4162,N_3887,N_2050);
or U4163 (N_4163,N_3878,N_2078);
nor U4164 (N_4164,N_2161,N_2214);
or U4165 (N_4165,N_3596,N_3266);
nor U4166 (N_4166,N_2037,N_3793);
xnor U4167 (N_4167,N_2370,N_3541);
nand U4168 (N_4168,N_2548,N_3505);
and U4169 (N_4169,N_3326,N_2500);
nor U4170 (N_4170,N_3454,N_3758);
or U4171 (N_4171,N_2345,N_3798);
xnor U4172 (N_4172,N_3221,N_2052);
nor U4173 (N_4173,N_2220,N_3641);
nor U4174 (N_4174,N_2125,N_2407);
nor U4175 (N_4175,N_2172,N_2042);
xor U4176 (N_4176,N_2087,N_2582);
and U4177 (N_4177,N_2778,N_2853);
xnor U4178 (N_4178,N_3582,N_2612);
nand U4179 (N_4179,N_2724,N_2810);
and U4180 (N_4180,N_2112,N_2750);
and U4181 (N_4181,N_2433,N_3944);
or U4182 (N_4182,N_2988,N_3830);
or U4183 (N_4183,N_2096,N_3241);
xnor U4184 (N_4184,N_2262,N_2346);
and U4185 (N_4185,N_2860,N_3531);
nor U4186 (N_4186,N_2117,N_3097);
and U4187 (N_4187,N_3857,N_2280);
nor U4188 (N_4188,N_3862,N_2337);
or U4189 (N_4189,N_2483,N_2607);
xnor U4190 (N_4190,N_2785,N_2992);
and U4191 (N_4191,N_3635,N_2264);
nand U4192 (N_4192,N_3985,N_3446);
and U4193 (N_4193,N_2712,N_3864);
and U4194 (N_4194,N_2228,N_2791);
or U4195 (N_4195,N_2176,N_3779);
or U4196 (N_4196,N_2762,N_3132);
nor U4197 (N_4197,N_3953,N_2924);
nor U4198 (N_4198,N_3858,N_2372);
nand U4199 (N_4199,N_3826,N_3829);
and U4200 (N_4200,N_3217,N_2197);
nor U4201 (N_4201,N_2529,N_2196);
and U4202 (N_4202,N_2578,N_2666);
or U4203 (N_4203,N_3161,N_3856);
and U4204 (N_4204,N_3036,N_3404);
nand U4205 (N_4205,N_3486,N_2864);
nor U4206 (N_4206,N_3080,N_3653);
nor U4207 (N_4207,N_2450,N_3920);
and U4208 (N_4208,N_2966,N_3613);
xnor U4209 (N_4209,N_2634,N_3005);
nor U4210 (N_4210,N_3627,N_3527);
or U4211 (N_4211,N_3601,N_2718);
nand U4212 (N_4212,N_2051,N_2608);
and U4213 (N_4213,N_3518,N_2164);
nand U4214 (N_4214,N_3822,N_3865);
nor U4215 (N_4215,N_3139,N_3397);
and U4216 (N_4216,N_2021,N_2993);
xor U4217 (N_4217,N_3766,N_3589);
xor U4218 (N_4218,N_2190,N_2388);
nand U4219 (N_4219,N_3196,N_2650);
or U4220 (N_4220,N_2296,N_3482);
or U4221 (N_4221,N_2459,N_2340);
nand U4222 (N_4222,N_3208,N_3152);
nand U4223 (N_4223,N_3162,N_2964);
or U4224 (N_4224,N_3654,N_3685);
nor U4225 (N_4225,N_2595,N_3246);
xor U4226 (N_4226,N_2011,N_2213);
and U4227 (N_4227,N_2035,N_3592);
and U4228 (N_4228,N_3511,N_3249);
or U4229 (N_4229,N_3958,N_2062);
nand U4230 (N_4230,N_3986,N_3915);
and U4231 (N_4231,N_3389,N_3109);
nand U4232 (N_4232,N_2544,N_3361);
or U4233 (N_4233,N_2435,N_2980);
xor U4234 (N_4234,N_3295,N_3522);
or U4235 (N_4235,N_2070,N_2336);
or U4236 (N_4236,N_2670,N_3255);
or U4237 (N_4237,N_3155,N_2923);
nand U4238 (N_4238,N_3882,N_3534);
or U4239 (N_4239,N_3148,N_3043);
nor U4240 (N_4240,N_2613,N_3580);
and U4241 (N_4241,N_3442,N_3061);
and U4242 (N_4242,N_2285,N_2292);
nand U4243 (N_4243,N_3930,N_2278);
xnor U4244 (N_4244,N_2297,N_2697);
and U4245 (N_4245,N_3879,N_2399);
and U4246 (N_4246,N_2787,N_3667);
nand U4247 (N_4247,N_3789,N_3019);
and U4248 (N_4248,N_2903,N_2234);
nand U4249 (N_4249,N_2254,N_2604);
and U4250 (N_4250,N_2764,N_2519);
and U4251 (N_4251,N_3607,N_2668);
nand U4252 (N_4252,N_2259,N_2417);
or U4253 (N_4253,N_3943,N_2797);
nand U4254 (N_4254,N_2458,N_3623);
nor U4255 (N_4255,N_2926,N_3165);
and U4256 (N_4256,N_3914,N_3921);
nand U4257 (N_4257,N_3608,N_2579);
and U4258 (N_4258,N_2646,N_2002);
xor U4259 (N_4259,N_2882,N_3844);
and U4260 (N_4260,N_2693,N_3318);
and U4261 (N_4261,N_2728,N_3538);
nand U4262 (N_4262,N_2132,N_2921);
nor U4263 (N_4263,N_2091,N_3996);
nand U4264 (N_4264,N_3674,N_2150);
or U4265 (N_4265,N_2835,N_2139);
nor U4266 (N_4266,N_3615,N_2657);
nor U4267 (N_4267,N_2324,N_2840);
or U4268 (N_4268,N_2746,N_2484);
nand U4269 (N_4269,N_2601,N_3838);
and U4270 (N_4270,N_3247,N_2979);
nor U4271 (N_4271,N_3431,N_2328);
and U4272 (N_4272,N_3683,N_2664);
nand U4273 (N_4273,N_2636,N_2502);
nor U4274 (N_4274,N_2506,N_2478);
nand U4275 (N_4275,N_2376,N_3317);
xor U4276 (N_4276,N_2454,N_2747);
and U4277 (N_4277,N_2959,N_2156);
or U4278 (N_4278,N_3587,N_3895);
and U4279 (N_4279,N_2198,N_2239);
nor U4280 (N_4280,N_3445,N_3716);
nor U4281 (N_4281,N_3902,N_2676);
nor U4282 (N_4282,N_2475,N_2437);
and U4283 (N_4283,N_3951,N_3380);
or U4284 (N_4284,N_2862,N_2080);
or U4285 (N_4285,N_3024,N_3414);
nor U4286 (N_4286,N_2887,N_2230);
nand U4287 (N_4287,N_2804,N_3910);
and U4288 (N_4288,N_3617,N_3082);
and U4289 (N_4289,N_2813,N_3365);
and U4290 (N_4290,N_2056,N_3491);
or U4291 (N_4291,N_2456,N_2990);
nand U4292 (N_4292,N_3321,N_3931);
xnor U4293 (N_4293,N_2106,N_2530);
nor U4294 (N_4294,N_2916,N_2918);
and U4295 (N_4295,N_3614,N_3034);
nand U4296 (N_4296,N_3959,N_3173);
or U4297 (N_4297,N_3720,N_2852);
nand U4298 (N_4298,N_2786,N_2510);
or U4299 (N_4299,N_2045,N_3157);
nand U4300 (N_4300,N_3556,N_3441);
nor U4301 (N_4301,N_2658,N_2795);
and U4302 (N_4302,N_3340,N_3984);
or U4303 (N_4303,N_2320,N_2186);
nand U4304 (N_4304,N_2991,N_3636);
nor U4305 (N_4305,N_2260,N_3863);
nand U4306 (N_4306,N_2626,N_2257);
nand U4307 (N_4307,N_3212,N_2754);
nand U4308 (N_4308,N_3098,N_3417);
and U4309 (N_4309,N_3410,N_3969);
nand U4310 (N_4310,N_3316,N_3176);
nand U4311 (N_4311,N_3497,N_3645);
and U4312 (N_4312,N_2339,N_2434);
xor U4313 (N_4313,N_3966,N_2071);
or U4314 (N_4314,N_2291,N_2107);
and U4315 (N_4315,N_2333,N_3237);
xor U4316 (N_4316,N_3029,N_3007);
or U4317 (N_4317,N_3228,N_3489);
and U4318 (N_4318,N_2914,N_2426);
and U4319 (N_4319,N_3642,N_2444);
or U4320 (N_4320,N_2597,N_2507);
or U4321 (N_4321,N_3001,N_2252);
or U4322 (N_4322,N_3840,N_3377);
nand U4323 (N_4323,N_3100,N_2794);
nor U4324 (N_4324,N_2188,N_2047);
nor U4325 (N_4325,N_2975,N_2669);
nor U4326 (N_4326,N_2967,N_2192);
nand U4327 (N_4327,N_2869,N_3265);
xnor U4328 (N_4328,N_2114,N_3332);
nor U4329 (N_4329,N_3868,N_2276);
or U4330 (N_4330,N_2583,N_3480);
nor U4331 (N_4331,N_2758,N_3922);
or U4332 (N_4332,N_2696,N_2479);
and U4333 (N_4333,N_2383,N_2890);
nor U4334 (N_4334,N_2266,N_3374);
nor U4335 (N_4335,N_3069,N_3578);
nand U4336 (N_4336,N_2585,N_3927);
nor U4337 (N_4337,N_2683,N_2839);
and U4338 (N_4338,N_3823,N_3884);
nor U4339 (N_4339,N_3835,N_3476);
nand U4340 (N_4340,N_2282,N_2588);
or U4341 (N_4341,N_2817,N_3320);
or U4342 (N_4342,N_2559,N_2148);
or U4343 (N_4343,N_3650,N_3089);
and U4344 (N_4344,N_2713,N_2557);
nor U4345 (N_4345,N_3117,N_3665);
and U4346 (N_4346,N_3494,N_3828);
nor U4347 (N_4347,N_3791,N_2201);
or U4348 (N_4348,N_2616,N_3867);
nand U4349 (N_4349,N_3408,N_3121);
or U4350 (N_4350,N_3633,N_3992);
or U4351 (N_4351,N_2784,N_3336);
and U4352 (N_4352,N_2289,N_3540);
and U4353 (N_4353,N_2773,N_3597);
nand U4354 (N_4354,N_2653,N_2373);
nor U4355 (N_4355,N_3192,N_2207);
and U4356 (N_4356,N_3968,N_2999);
xor U4357 (N_4357,N_3219,N_2981);
or U4358 (N_4358,N_3845,N_3214);
xor U4359 (N_4359,N_3370,N_3119);
nor U4360 (N_4360,N_3723,N_3359);
or U4361 (N_4361,N_3092,N_2902);
nand U4362 (N_4362,N_2017,N_3606);
and U4363 (N_4363,N_2393,N_2246);
nor U4364 (N_4364,N_3430,N_3429);
nand U4365 (N_4365,N_2897,N_3364);
nor U4366 (N_4366,N_2097,N_2820);
or U4367 (N_4367,N_3947,N_2467);
nor U4368 (N_4368,N_2033,N_3519);
and U4369 (N_4369,N_3649,N_2586);
nand U4370 (N_4370,N_3841,N_3175);
nand U4371 (N_4371,N_3393,N_3581);
nand U4372 (N_4372,N_2419,N_2102);
or U4373 (N_4373,N_2397,N_2546);
nor U4374 (N_4374,N_3141,N_2064);
and U4375 (N_4375,N_3630,N_3737);
nand U4376 (N_4376,N_3801,N_2625);
nand U4377 (N_4377,N_3971,N_3819);
xnor U4378 (N_4378,N_2218,N_3852);
nor U4379 (N_4379,N_2564,N_3349);
xor U4380 (N_4380,N_2301,N_3712);
or U4381 (N_4381,N_3763,N_3169);
nand U4382 (N_4382,N_3025,N_3328);
nand U4383 (N_4383,N_2572,N_3548);
nor U4384 (N_4384,N_2487,N_3094);
and U4385 (N_4385,N_2012,N_2555);
and U4386 (N_4386,N_3709,N_2776);
nor U4387 (N_4387,N_2424,N_3978);
nand U4388 (N_4388,N_3727,N_3565);
and U4389 (N_4389,N_2929,N_2652);
nand U4390 (N_4390,N_2495,N_3203);
and U4391 (N_4391,N_2503,N_2899);
or U4392 (N_4392,N_3989,N_2229);
xnor U4393 (N_4393,N_3136,N_2960);
or U4394 (N_4394,N_2089,N_3016);
nand U4395 (N_4395,N_2752,N_2602);
or U4396 (N_4396,N_2325,N_2870);
or U4397 (N_4397,N_2256,N_2760);
and U4398 (N_4398,N_3433,N_3485);
or U4399 (N_4399,N_2645,N_2974);
and U4400 (N_4400,N_3218,N_2912);
xnor U4401 (N_4401,N_3866,N_3960);
xor U4402 (N_4402,N_2423,N_2295);
nand U4403 (N_4403,N_3126,N_3258);
nor U4404 (N_4404,N_2629,N_2018);
nor U4405 (N_4405,N_2401,N_3748);
nor U4406 (N_4406,N_2733,N_3004);
nor U4407 (N_4407,N_2193,N_3813);
and U4408 (N_4408,N_2986,N_2379);
and U4409 (N_4409,N_3634,N_2343);
nand U4410 (N_4410,N_2086,N_2962);
or U4411 (N_4411,N_2195,N_3059);
nor U4412 (N_4412,N_3357,N_2181);
nand U4413 (N_4413,N_3583,N_3833);
nand U4414 (N_4414,N_2240,N_2943);
and U4415 (N_4415,N_2165,N_2957);
xor U4416 (N_4416,N_2800,N_3834);
and U4417 (N_4417,N_3803,N_2667);
nand U4418 (N_4418,N_2359,N_2334);
nor U4419 (N_4419,N_3553,N_2120);
xor U4420 (N_4420,N_2638,N_3591);
xnor U4421 (N_4421,N_2875,N_3780);
nor U4422 (N_4422,N_3595,N_2061);
nand U4423 (N_4423,N_3461,N_3901);
xor U4424 (N_4424,N_3892,N_2977);
or U4425 (N_4425,N_2730,N_3605);
nor U4426 (N_4426,N_3514,N_3568);
and U4427 (N_4427,N_2637,N_3288);
and U4428 (N_4428,N_3128,N_3525);
and U4429 (N_4429,N_2428,N_2335);
and U4430 (N_4430,N_2948,N_3205);
nor U4431 (N_4431,N_3206,N_3974);
or U4432 (N_4432,N_2231,N_3980);
and U4433 (N_4433,N_3718,N_3490);
nor U4434 (N_4434,N_2806,N_3101);
or U4435 (N_4435,N_3435,N_3302);
nand U4436 (N_4436,N_2332,N_3366);
nand U4437 (N_4437,N_3508,N_2138);
nand U4438 (N_4438,N_3782,N_2873);
and U4439 (N_4439,N_2631,N_2378);
xor U4440 (N_4440,N_3020,N_2076);
xnor U4441 (N_4441,N_2893,N_3888);
xor U4442 (N_4442,N_2749,N_2189);
nor U4443 (N_4443,N_2244,N_3010);
or U4444 (N_4444,N_2928,N_2931);
nand U4445 (N_4445,N_3213,N_3030);
nor U4446 (N_4446,N_3871,N_3276);
and U4447 (N_4447,N_3090,N_3821);
nand U4448 (N_4448,N_2382,N_2644);
and U4449 (N_4449,N_3096,N_3330);
nor U4450 (N_4450,N_2452,N_2844);
nor U4451 (N_4451,N_3679,N_3269);
nor U4452 (N_4452,N_3695,N_3073);
and U4453 (N_4453,N_2267,N_2031);
nand U4454 (N_4454,N_2169,N_2880);
and U4455 (N_4455,N_2512,N_2068);
xor U4456 (N_4456,N_3193,N_2177);
or U4457 (N_4457,N_2163,N_3347);
or U4458 (N_4458,N_2907,N_2751);
nand U4459 (N_4459,N_3479,N_2788);
nand U4460 (N_4460,N_3006,N_2700);
nand U4461 (N_4461,N_3167,N_3471);
nand U4462 (N_4462,N_3243,N_3095);
nor U4463 (N_4463,N_2662,N_2889);
or U4464 (N_4464,N_3911,N_2352);
nand U4465 (N_4465,N_3131,N_2577);
nor U4466 (N_4466,N_3837,N_2358);
and U4467 (N_4467,N_3286,N_3062);
or U4468 (N_4468,N_3227,N_3473);
nand U4469 (N_4469,N_3552,N_2400);
and U4470 (N_4470,N_3707,N_3263);
nand U4471 (N_4471,N_3053,N_2098);
nor U4472 (N_4472,N_3415,N_2111);
nand U4473 (N_4473,N_3372,N_3670);
nand U4474 (N_4474,N_2920,N_2524);
or U4475 (N_4475,N_2066,N_3929);
and U4476 (N_4476,N_2528,N_3245);
or U4477 (N_4477,N_2978,N_3260);
nor U4478 (N_4478,N_3297,N_3385);
or U4479 (N_4479,N_3232,N_3860);
xor U4480 (N_4480,N_2127,N_2354);
nand U4481 (N_4481,N_3506,N_3037);
nor U4482 (N_4482,N_2731,N_3164);
nor U4483 (N_4483,N_2554,N_2594);
or U4484 (N_4484,N_2611,N_3309);
nand U4485 (N_4485,N_3125,N_3198);
and U4486 (N_4486,N_3767,N_2691);
or U4487 (N_4487,N_2392,N_3403);
or U4488 (N_4488,N_3809,N_3182);
nor U4489 (N_4489,N_3017,N_2170);
and U4490 (N_4490,N_3820,N_2856);
nor U4491 (N_4491,N_3880,N_3439);
and U4492 (N_4492,N_2385,N_3935);
and U4493 (N_4493,N_3970,N_3598);
or U4494 (N_4494,N_2649,N_2398);
nor U4495 (N_4495,N_2729,N_2711);
xnor U4496 (N_4496,N_3280,N_3156);
and U4497 (N_4497,N_2469,N_3180);
nand U4498 (N_4498,N_2248,N_2004);
nand U4499 (N_4499,N_3734,N_3923);
nand U4500 (N_4500,N_3684,N_3640);
or U4501 (N_4501,N_3588,N_2242);
or U4502 (N_4502,N_2639,N_3805);
and U4503 (N_4503,N_2208,N_2223);
or U4504 (N_4504,N_3207,N_3492);
and U4505 (N_4505,N_2299,N_2672);
and U4506 (N_4506,N_2249,N_3725);
nor U4507 (N_4507,N_2438,N_2041);
and U4508 (N_4508,N_2896,N_3561);
or U4509 (N_4509,N_3774,N_2722);
and U4510 (N_4510,N_3515,N_3666);
and U4511 (N_4511,N_3178,N_3655);
and U4512 (N_4512,N_2095,N_3967);
and U4513 (N_4513,N_3470,N_3699);
or U4514 (N_4514,N_3040,N_3904);
and U4515 (N_4515,N_2686,N_2904);
nand U4516 (N_4516,N_3009,N_3499);
xnor U4517 (N_4517,N_3512,N_3762);
or U4518 (N_4518,N_2493,N_2351);
xor U4519 (N_4519,N_2298,N_2717);
or U4520 (N_4520,N_2692,N_3657);
nand U4521 (N_4521,N_2217,N_3532);
nor U4522 (N_4522,N_3831,N_2702);
or U4523 (N_4523,N_2775,N_3012);
xnor U4524 (N_4524,N_3790,N_3150);
nand U4525 (N_4525,N_3997,N_2961);
nor U4526 (N_4526,N_2362,N_3618);
or U4527 (N_4527,N_3609,N_2774);
nor U4528 (N_4528,N_2093,N_2251);
nor U4529 (N_4529,N_2803,N_3478);
or U4530 (N_4530,N_2741,N_2630);
nor U4531 (N_4531,N_2770,N_3406);
xnor U4532 (N_4532,N_2143,N_2411);
nand U4533 (N_4533,N_3919,N_2618);
nor U4534 (N_4534,N_2954,N_3477);
or U4535 (N_4535,N_2038,N_3335);
or U4536 (N_4536,N_2053,N_3475);
nand U4537 (N_4537,N_2353,N_2024);
nor U4538 (N_4538,N_3116,N_3058);
or U4539 (N_4539,N_3566,N_3190);
or U4540 (N_4540,N_3753,N_3544);
or U4541 (N_4541,N_3108,N_3802);
nor U4542 (N_4542,N_3344,N_2545);
nand U4543 (N_4543,N_3637,N_3594);
nor U4544 (N_4544,N_3104,N_2525);
nand U4545 (N_4545,N_3462,N_3571);
nor U4546 (N_4546,N_3209,N_3643);
xor U4547 (N_4547,N_3054,N_2738);
or U4548 (N_4548,N_2341,N_2827);
nand U4549 (N_4549,N_3401,N_2155);
or U4550 (N_4550,N_2678,N_3705);
or U4551 (N_4551,N_2025,N_3428);
or U4552 (N_4552,N_3622,N_2137);
nand U4553 (N_4553,N_3795,N_3463);
nor U4554 (N_4554,N_3869,N_3242);
nand U4555 (N_4555,N_2915,N_2006);
xor U4556 (N_4556,N_2782,N_2514);
or U4557 (N_4557,N_3808,N_2331);
or U4558 (N_4558,N_3963,N_3407);
or U4559 (N_4559,N_3692,N_3516);
nand U4560 (N_4560,N_2861,N_3191);
xnor U4561 (N_4561,N_3103,N_3015);
nand U4562 (N_4562,N_2609,N_2140);
xor U4563 (N_4563,N_2847,N_3554);
and U4564 (N_4564,N_3827,N_2836);
xor U4565 (N_4565,N_3771,N_3567);
nor U4566 (N_4566,N_2727,N_3662);
xor U4567 (N_4567,N_3353,N_2973);
nand U4568 (N_4568,N_2906,N_3262);
or U4569 (N_4569,N_3988,N_2072);
nand U4570 (N_4570,N_2060,N_2390);
or U4571 (N_4571,N_3839,N_3252);
nor U4572 (N_4572,N_2665,N_3458);
nand U4573 (N_4573,N_3575,N_3244);
and U4574 (N_4574,N_3027,N_2952);
nand U4575 (N_4575,N_2561,N_3375);
nand U4576 (N_4576,N_2917,N_3304);
or U4577 (N_4577,N_3419,N_2740);
nor U4578 (N_4578,N_3982,N_2034);
nor U4579 (N_4579,N_2371,N_3047);
xnor U4580 (N_4580,N_2360,N_2552);
or U4581 (N_4581,N_3691,N_3050);
and U4582 (N_4582,N_3913,N_3183);
nand U4583 (N_4583,N_2687,N_2511);
nor U4584 (N_4584,N_2241,N_2809);
or U4585 (N_4585,N_2537,N_2162);
nand U4586 (N_4586,N_2323,N_2342);
or U4587 (N_4587,N_3632,N_2461);
nor U4588 (N_4588,N_3577,N_3975);
xor U4589 (N_4589,N_3675,N_2569);
or U4590 (N_4590,N_2225,N_3273);
or U4591 (N_4591,N_3668,N_3500);
and U4592 (N_4592,N_2233,N_3781);
or U4593 (N_4593,N_3405,N_3450);
and U4594 (N_4594,N_3338,N_2798);
xnor U4595 (N_4595,N_2321,N_2306);
or U4596 (N_4596,N_2789,N_2279);
or U4597 (N_4597,N_2849,N_3170);
and U4598 (N_4598,N_3376,N_2640);
and U4599 (N_4599,N_3013,N_3171);
or U4600 (N_4600,N_2453,N_2886);
nor U4601 (N_4601,N_2811,N_2617);
nor U4602 (N_4602,N_3052,N_3003);
and U4603 (N_4603,N_3339,N_2480);
nor U4604 (N_4604,N_3311,N_3434);
nand U4605 (N_4605,N_2160,N_3742);
nor U4606 (N_4606,N_2542,N_3671);
nor U4607 (N_4607,N_3457,N_3925);
nand U4608 (N_4608,N_3750,N_3842);
nor U4609 (N_4609,N_3938,N_3091);
or U4610 (N_4610,N_2779,N_3137);
nand U4611 (N_4611,N_2491,N_3631);
or U4612 (N_4612,N_3130,N_2968);
nand U4613 (N_4613,N_2805,N_2584);
nand U4614 (N_4614,N_3698,N_3772);
nor U4615 (N_4615,N_3850,N_2998);
nand U4616 (N_4616,N_3939,N_2136);
xnor U4617 (N_4617,N_2855,N_2501);
nand U4618 (N_4618,N_3872,N_2149);
or U4619 (N_4619,N_2365,N_2473);
and U4620 (N_4620,N_2173,N_3950);
nand U4621 (N_4621,N_2739,N_2571);
nor U4622 (N_4622,N_2888,N_3539);
nor U4623 (N_4623,N_3903,N_3383);
and U4624 (N_4624,N_3373,N_3194);
nand U4625 (N_4625,N_2153,N_2633);
nand U4626 (N_4626,N_2049,N_2416);
nand U4627 (N_4627,N_2767,N_2808);
nor U4628 (N_4628,N_2562,N_2763);
or U4629 (N_4629,N_2566,N_2560);
or U4630 (N_4630,N_2759,N_3238);
nor U4631 (N_4631,N_3584,N_3323);
xnor U4632 (N_4632,N_2043,N_2614);
and U4633 (N_4633,N_3703,N_2937);
nand U4634 (N_4634,N_2308,N_2755);
and U4635 (N_4635,N_3049,N_2558);
nand U4636 (N_4636,N_3787,N_2901);
nor U4637 (N_4637,N_2698,N_2044);
or U4638 (N_4638,N_2236,N_3432);
xor U4639 (N_4639,N_2843,N_2420);
nand U4640 (N_4640,N_3275,N_2269);
or U4641 (N_4641,N_3289,N_2858);
or U4642 (N_4642,N_3585,N_3395);
xnor U4643 (N_4643,N_3382,N_3484);
nand U4644 (N_4644,N_3730,N_3660);
and U4645 (N_4645,N_3811,N_3378);
nor U4646 (N_4646,N_2347,N_2812);
and U4647 (N_4647,N_2326,N_3278);
and U4648 (N_4648,N_3077,N_3187);
and U4649 (N_4649,N_3379,N_3896);
xor U4650 (N_4650,N_2930,N_3422);
or U4651 (N_4651,N_2549,N_3449);
or U4652 (N_4652,N_2553,N_2987);
xor U4653 (N_4653,N_2425,N_2447);
and U4654 (N_4654,N_2356,N_3168);
nand U4655 (N_4655,N_3070,N_3426);
or U4656 (N_4656,N_3086,N_2309);
nand U4657 (N_4657,N_2159,N_3420);
nand U4658 (N_4658,N_3926,N_2720);
and U4659 (N_4659,N_2596,N_3521);
and U4660 (N_4660,N_3680,N_2799);
nand U4661 (N_4661,N_2290,N_3064);
nor U4662 (N_4662,N_3075,N_2941);
or U4663 (N_4663,N_2939,N_2971);
nor U4664 (N_4664,N_3051,N_3704);
nand U4665 (N_4665,N_2895,N_2777);
nand U4666 (N_4666,N_3481,N_2199);
nand U4667 (N_4667,N_2925,N_3371);
xnor U4668 (N_4668,N_3021,N_3682);
or U4669 (N_4669,N_3409,N_2515);
nand U4670 (N_4670,N_2821,N_2677);
nor U4671 (N_4671,N_3327,N_3142);
nand U4672 (N_4672,N_2059,N_3917);
nand U4673 (N_4673,N_3216,N_2872);
nor U4674 (N_4674,N_2848,N_3093);
xnor U4675 (N_4675,N_2756,N_3251);
xor U4676 (N_4676,N_3277,N_2831);
nor U4677 (N_4677,N_2891,N_3749);
nand U4678 (N_4678,N_2101,N_3932);
or U4679 (N_4679,N_3042,N_2488);
or U4680 (N_4680,N_3952,N_3543);
or U4681 (N_4681,N_3472,N_2029);
xnor U4682 (N_4682,N_2055,N_3078);
and U4683 (N_4683,N_2374,N_3310);
nand U4684 (N_4684,N_2058,N_2574);
xor U4685 (N_4685,N_2661,N_3724);
and U4686 (N_4686,N_2288,N_2570);
nand U4687 (N_4687,N_3533,N_3520);
nor U4688 (N_4688,N_2790,N_3715);
or U4689 (N_4689,N_3253,N_3154);
nor U4690 (N_4690,N_2219,N_3928);
nand U4691 (N_4691,N_2536,N_2030);
or U4692 (N_4692,N_3381,N_2947);
xor U4693 (N_4693,N_3905,N_3487);
and U4694 (N_4694,N_2632,N_2622);
nand U4695 (N_4695,N_3964,N_3981);
xor U4696 (N_4696,N_3303,N_2182);
and U4697 (N_4697,N_3751,N_3687);
nor U4698 (N_4698,N_2133,N_3112);
and U4699 (N_4699,N_3358,N_3324);
nand U4700 (N_4700,N_3284,N_2174);
or U4701 (N_4701,N_2413,N_3832);
and U4702 (N_4702,N_2235,N_2534);
nor U4703 (N_4703,N_2100,N_3777);
or U4704 (N_4704,N_2380,N_3038);
nand U4705 (N_4705,N_2039,N_3224);
or U4706 (N_4706,N_2863,N_2460);
or U4707 (N_4707,N_2753,N_2885);
nor U4708 (N_4708,N_3870,N_2412);
nor U4709 (N_4709,N_2591,N_2083);
and U4710 (N_4710,N_2019,N_2316);
or U4711 (N_4711,N_3267,N_2932);
nand U4712 (N_4712,N_3334,N_2465);
and U4713 (N_4713,N_2471,N_3392);
and U4714 (N_4714,N_2627,N_3438);
or U4715 (N_4715,N_3973,N_3713);
xor U4716 (N_4716,N_3817,N_2826);
nor U4717 (N_4717,N_2489,N_2377);
or U4718 (N_4718,N_2850,N_2258);
and U4719 (N_4719,N_2989,N_3503);
nor U4720 (N_4720,N_2772,N_2619);
or U4721 (N_4721,N_3222,N_3732);
and U4722 (N_4722,N_2386,N_3396);
or U4723 (N_4723,N_3387,N_2350);
or U4724 (N_4724,N_2090,N_3498);
or U4725 (N_4725,N_2294,N_2695);
nor U4726 (N_4726,N_2436,N_2283);
nand U4727 (N_4727,N_2126,N_3181);
nand U4728 (N_4728,N_2245,N_2761);
nor U4729 (N_4729,N_3127,N_3547);
or U4730 (N_4730,N_2187,N_3306);
and U4731 (N_4731,N_2409,N_2023);
or U4732 (N_4732,N_2508,N_2243);
nor U4733 (N_4733,N_3900,N_3110);
nor U4734 (N_4734,N_2224,N_2996);
and U4735 (N_4735,N_3402,N_2005);
nand U4736 (N_4736,N_3961,N_2284);
and U4737 (N_4737,N_3647,N_3257);
or U4738 (N_4738,N_2704,N_3390);
nor U4739 (N_4739,N_3279,N_3501);
nand U4740 (N_4740,N_3648,N_2307);
or U4741 (N_4741,N_2522,N_3885);
or U4742 (N_4742,N_2268,N_2009);
nor U4743 (N_4743,N_2834,N_2158);
and U4744 (N_4744,N_3600,N_2854);
and U4745 (N_4745,N_2222,N_2841);
or U4746 (N_4746,N_3861,N_3792);
or U4747 (N_4747,N_3063,N_3185);
nor U4748 (N_4748,N_3620,N_2026);
nor U4749 (N_4749,N_2509,N_2581);
or U4750 (N_4750,N_2092,N_2110);
nand U4751 (N_4751,N_3459,N_3646);
nand U4752 (N_4752,N_2387,N_3313);
nand U4753 (N_4753,N_2846,N_3440);
xnor U4754 (N_4754,N_3825,N_3048);
and U4755 (N_4755,N_3836,N_2468);
and U4756 (N_4756,N_2118,N_2871);
nor U4757 (N_4757,N_3282,N_3812);
or U4758 (N_4758,N_2832,N_2517);
nor U4759 (N_4759,N_2451,N_3268);
or U4760 (N_4760,N_3661,N_2580);
or U4761 (N_4761,N_2737,N_3177);
and U4762 (N_4762,N_3545,N_2851);
and U4763 (N_4763,N_2568,N_3717);
nor U4764 (N_4764,N_2768,N_2067);
and U4765 (N_4765,N_3184,N_3134);
nand U4766 (N_4766,N_3071,N_2205);
nand U4767 (N_4767,N_2464,N_3603);
nand U4768 (N_4768,N_3760,N_3994);
or U4769 (N_4769,N_2135,N_2540);
nand U4770 (N_4770,N_3890,N_2780);
or U4771 (N_4771,N_3509,N_2642);
or U4772 (N_4772,N_2927,N_3800);
nor U4773 (N_4773,N_3087,N_3172);
xnor U4774 (N_4774,N_2815,N_3847);
and U4775 (N_4775,N_3274,N_2485);
and U4776 (N_4776,N_3290,N_3225);
and U4777 (N_4777,N_2721,N_2748);
or U4778 (N_4778,N_2105,N_3083);
nand U4779 (N_4779,N_3233,N_3558);
xor U4780 (N_4780,N_3254,N_2410);
nand U4781 (N_4781,N_3851,N_2366);
and U4782 (N_4782,N_2995,N_2355);
or U4783 (N_4783,N_2069,N_2513);
nor U4784 (N_4784,N_2286,N_3876);
or U4785 (N_4785,N_3240,N_3105);
xor U4786 (N_4786,N_3816,N_3755);
nor U4787 (N_4787,N_2414,N_3883);
nor U4788 (N_4788,N_2403,N_3039);
nor U4789 (N_4789,N_3283,N_2271);
nand U4790 (N_4790,N_2951,N_2910);
xor U4791 (N_4791,N_3569,N_2124);
and U4792 (N_4792,N_3018,N_3765);
and U4793 (N_4793,N_3011,N_3756);
xor U4794 (N_4794,N_2432,N_3118);
and U4795 (N_4795,N_2216,N_3740);
and U4796 (N_4796,N_2593,N_3934);
and U4797 (N_4797,N_3270,N_2448);
nand U4798 (N_4798,N_2983,N_3783);
nor U4799 (N_4799,N_2363,N_2745);
nor U4800 (N_4800,N_3124,N_3735);
nor U4801 (N_4801,N_2716,N_3942);
nor U4802 (N_4802,N_2592,N_3496);
nand U4803 (N_4803,N_2215,N_2719);
and U4804 (N_4804,N_3160,N_3688);
and U4805 (N_4805,N_2206,N_2498);
nand U4806 (N_4806,N_3234,N_2824);
and U4807 (N_4807,N_3033,N_3067);
nor U4808 (N_4808,N_2422,N_3602);
and U4809 (N_4809,N_3689,N_2936);
and U4810 (N_4810,N_2322,N_3133);
or U4811 (N_4811,N_2010,N_2261);
and U4812 (N_4812,N_3452,N_2157);
and U4813 (N_4813,N_3976,N_3299);
nor U4814 (N_4814,N_3236,N_3106);
or U4815 (N_4815,N_3853,N_3423);
and U4816 (N_4816,N_3319,N_2624);
and U4817 (N_4817,N_2660,N_2171);
or U4818 (N_4818,N_3610,N_3729);
nand U4819 (N_4819,N_3026,N_3736);
nand U4820 (N_4820,N_2589,N_3002);
nand U4821 (N_4821,N_2565,N_2109);
or U4822 (N_4822,N_3291,N_2701);
or U4823 (N_4823,N_3559,N_3174);
or U4824 (N_4824,N_3530,N_3416);
nor U4825 (N_4825,N_3625,N_3965);
nand U4826 (N_4826,N_2765,N_3690);
or U4827 (N_4827,N_3115,N_2396);
nand U4828 (N_4828,N_3983,N_3363);
xor U4829 (N_4829,N_3322,N_2599);
and U4830 (N_4830,N_2603,N_2838);
or U4831 (N_4831,N_2504,N_3329);
or U4832 (N_4832,N_3849,N_2202);
nand U4833 (N_4833,N_3555,N_2094);
nor U4834 (N_4834,N_2945,N_3940);
or U4835 (N_4835,N_2270,N_3658);
or U4836 (N_4836,N_3368,N_2953);
nor U4837 (N_4837,N_2615,N_2429);
and U4838 (N_4838,N_2690,N_3757);
and U4839 (N_4839,N_3391,N_2166);
and U4840 (N_4840,N_3398,N_3411);
nor U4841 (N_4841,N_2877,N_3573);
nor U4842 (N_4842,N_2015,N_3738);
or U4843 (N_4843,N_3287,N_3536);
or U4844 (N_4844,N_2956,N_3700);
and U4845 (N_4845,N_3562,N_2305);
or U4846 (N_4846,N_2867,N_2349);
xor U4847 (N_4847,N_3202,N_2865);
nand U4848 (N_4848,N_2144,N_2476);
and U4849 (N_4849,N_3785,N_2919);
or U4850 (N_4850,N_2881,N_2958);
and U4851 (N_4851,N_3619,N_2972);
nand U4852 (N_4852,N_3369,N_3549);
nand U4853 (N_4853,N_2406,N_3560);
or U4854 (N_4854,N_3451,N_2338);
xnor U4855 (N_4855,N_3045,N_3551);
nor U4856 (N_4856,N_2709,N_3810);
nor U4857 (N_4857,N_2168,N_3065);
nand U4858 (N_4858,N_2913,N_3722);
and U4859 (N_4859,N_2922,N_2533);
xnor U4860 (N_4860,N_2940,N_3673);
nand U4861 (N_4861,N_3195,N_3948);
nor U4862 (N_4862,N_2946,N_2793);
and U4863 (N_4863,N_2694,N_3325);
or U4864 (N_4864,N_3728,N_2232);
nand U4865 (N_4865,N_2099,N_2985);
nand U4866 (N_4866,N_3362,N_3754);
or U4867 (N_4867,N_3355,N_2394);
nor U4868 (N_4868,N_3546,N_3991);
nand U4869 (N_4869,N_3796,N_2783);
and U4870 (N_4870,N_3281,N_3129);
xnor U4871 (N_4871,N_3874,N_3223);
and U4872 (N_4872,N_3197,N_3987);
nand U4873 (N_4873,N_3746,N_2310);
and U4874 (N_4874,N_3775,N_3916);
or U4875 (N_4875,N_3413,N_2859);
or U4876 (N_4876,N_3678,N_2648);
nand U4877 (N_4877,N_3563,N_3314);
or U4878 (N_4878,N_2781,N_3046);
nand U4879 (N_4879,N_2077,N_2178);
or U4880 (N_4880,N_2598,N_2703);
nand U4881 (N_4881,N_3526,N_3056);
or U4882 (N_4882,N_2663,N_3356);
or U4883 (N_4883,N_2357,N_3041);
or U4884 (N_4884,N_3576,N_2255);
or U4885 (N_4885,N_3897,N_2369);
nand U4886 (N_4886,N_3412,N_3201);
nor U4887 (N_4887,N_3629,N_3696);
nor U4888 (N_4888,N_2253,N_2732);
and U4889 (N_4889,N_2494,N_3726);
nand U4890 (N_4890,N_3028,N_3151);
nor U4891 (N_4891,N_3529,N_2814);
nand U4892 (N_4892,N_3333,N_2635);
and U4893 (N_4893,N_3466,N_3308);
and U4894 (N_4894,N_3189,N_3708);
and U4895 (N_4895,N_2472,N_2900);
xnor U4896 (N_4896,N_3122,N_2955);
and U4897 (N_4897,N_2391,N_3443);
nand U4898 (N_4898,N_2984,N_2445);
or U4899 (N_4899,N_2312,N_3149);
xnor U4900 (N_4900,N_3881,N_2982);
xnor U4901 (N_4901,N_3628,N_2942);
or U4902 (N_4902,N_2643,N_2499);
nor U4903 (N_4903,N_3298,N_2969);
xnor U4904 (N_4904,N_3517,N_3957);
or U4905 (N_4905,N_2057,N_3331);
xor U4906 (N_4906,N_2527,N_3799);
or U4907 (N_4907,N_2894,N_2113);
and U4908 (N_4908,N_2576,N_2415);
nor U4909 (N_4909,N_3464,N_2146);
or U4910 (N_4910,N_3697,N_3999);
xnor U4911 (N_4911,N_2088,N_2079);
nor U4912 (N_4912,N_2543,N_2647);
xor U4913 (N_4913,N_2621,N_2427);
and U4914 (N_4914,N_2275,N_3230);
and U4915 (N_4915,N_2792,N_3272);
nor U4916 (N_4916,N_2441,N_3231);
nand U4917 (N_4917,N_2884,N_3644);
nand U4918 (N_4918,N_3873,N_3474);
or U4919 (N_4919,N_3060,N_3346);
nor U4920 (N_4920,N_2532,N_3123);
nand U4921 (N_4921,N_2317,N_2547);
nor U4922 (N_4922,N_2368,N_2040);
and U4923 (N_4923,N_2179,N_2689);
or U4924 (N_4924,N_2520,N_3226);
or U4925 (N_4925,N_3342,N_3797);
nor U4926 (N_4926,N_2272,N_2655);
or U4927 (N_4927,N_3846,N_2154);
or U4928 (N_4928,N_3721,N_3513);
and U4929 (N_4929,N_2535,N_3877);
or U4930 (N_4930,N_2482,N_2014);
nand U4931 (N_4931,N_3773,N_2796);
and U4932 (N_4932,N_2575,N_3745);
nand U4933 (N_4933,N_3656,N_3510);
and U4934 (N_4934,N_2523,N_2054);
nor U4935 (N_4935,N_3163,N_2675);
nand U4936 (N_4936,N_2084,N_3235);
xor U4937 (N_4937,N_2938,N_2142);
nor U4938 (N_4938,N_2744,N_2736);
and U4939 (N_4939,N_3146,N_2131);
nor U4940 (N_4940,N_2300,N_3488);
or U4941 (N_4941,N_3972,N_3564);
and U4942 (N_4942,N_3360,N_3941);
nor U4943 (N_4943,N_3752,N_2518);
nor U4944 (N_4944,N_3113,N_3523);
or U4945 (N_4945,N_3706,N_2141);
nand U4946 (N_4946,N_3912,N_2082);
xor U4947 (N_4947,N_3044,N_2103);
and U4948 (N_4948,N_2022,N_3144);
and U4949 (N_4949,N_2734,N_3261);
and U4950 (N_4950,N_3120,N_3946);
nand U4951 (N_4951,N_3899,N_3384);
and U4952 (N_4952,N_3166,N_3784);
nor U4953 (N_4953,N_3611,N_3624);
and U4954 (N_4954,N_3794,N_2963);
nand U4955 (N_4955,N_2000,N_2210);
nand U4956 (N_4956,N_3114,N_2673);
nand U4957 (N_4957,N_2516,N_3300);
nand U4958 (N_4958,N_2122,N_2976);
nor U4959 (N_4959,N_3955,N_3215);
xnor U4960 (N_4960,N_3776,N_2606);
nor U4961 (N_4961,N_2726,N_3292);
nand U4962 (N_4962,N_2408,N_2563);
nand U4963 (N_4963,N_2477,N_3659);
and U4964 (N_4964,N_2823,N_3677);
nand U4965 (N_4965,N_3507,N_2656);
nor U4966 (N_4966,N_2659,N_2395);
nand U4967 (N_4967,N_2463,N_2628);
or U4968 (N_4968,N_2681,N_3107);
nor U4969 (N_4969,N_3102,N_3681);
nand U4970 (N_4970,N_3394,N_2277);
or U4971 (N_4971,N_2807,N_2742);
and U4972 (N_4972,N_2250,N_2587);
nand U4973 (N_4973,N_2238,N_2715);
nand U4974 (N_4974,N_2032,N_2486);
nor U4975 (N_4975,N_2539,N_3256);
nor U4976 (N_4976,N_2119,N_2600);
nor U4977 (N_4977,N_2375,N_3612);
and U4978 (N_4978,N_3891,N_3993);
and U4979 (N_4979,N_2878,N_3639);
and U4980 (N_4980,N_3066,N_2674);
or U4981 (N_4981,N_3804,N_3076);
nor U4982 (N_4982,N_3651,N_3669);
or U4983 (N_4983,N_2227,N_3711);
and U4984 (N_4984,N_3400,N_2802);
or U4985 (N_4985,N_2769,N_3909);
and U4986 (N_4986,N_2908,N_3057);
and U4987 (N_4987,N_3220,N_3886);
nor U4988 (N_4988,N_2449,N_3979);
or U4989 (N_4989,N_2265,N_2311);
or U4990 (N_4990,N_2430,N_3918);
nand U4991 (N_4991,N_3145,N_2063);
nor U4992 (N_4992,N_2439,N_2036);
and U4993 (N_4993,N_3937,N_2418);
and U4994 (N_4994,N_3875,N_3814);
xnor U4995 (N_4995,N_3945,N_3352);
nand U4996 (N_4996,N_2016,N_3468);
or U4997 (N_4997,N_2492,N_2123);
nand U4998 (N_4998,N_3337,N_3676);
nand U4999 (N_4999,N_3664,N_3456);
and U5000 (N_5000,N_2197,N_3273);
nand U5001 (N_5001,N_2419,N_3076);
nor U5002 (N_5002,N_3970,N_3533);
or U5003 (N_5003,N_2835,N_2493);
nor U5004 (N_5004,N_2719,N_2628);
and U5005 (N_5005,N_2511,N_3958);
nor U5006 (N_5006,N_3647,N_3938);
nand U5007 (N_5007,N_2939,N_3027);
xnor U5008 (N_5008,N_2642,N_2315);
nand U5009 (N_5009,N_3354,N_3192);
nand U5010 (N_5010,N_2608,N_2016);
nor U5011 (N_5011,N_3520,N_3108);
nor U5012 (N_5012,N_3488,N_3500);
or U5013 (N_5013,N_3717,N_2713);
nand U5014 (N_5014,N_3697,N_2421);
xor U5015 (N_5015,N_2045,N_3969);
and U5016 (N_5016,N_2854,N_2997);
xor U5017 (N_5017,N_3243,N_3432);
nand U5018 (N_5018,N_2784,N_3994);
or U5019 (N_5019,N_3778,N_3430);
nand U5020 (N_5020,N_3161,N_3386);
nor U5021 (N_5021,N_2593,N_2393);
nand U5022 (N_5022,N_3175,N_2065);
nor U5023 (N_5023,N_3311,N_2965);
and U5024 (N_5024,N_3432,N_3514);
nand U5025 (N_5025,N_2043,N_2609);
nand U5026 (N_5026,N_2666,N_2306);
or U5027 (N_5027,N_3157,N_3631);
nor U5028 (N_5028,N_2011,N_2023);
or U5029 (N_5029,N_3340,N_2148);
and U5030 (N_5030,N_2399,N_3544);
xor U5031 (N_5031,N_2565,N_3649);
xor U5032 (N_5032,N_2853,N_2293);
nand U5033 (N_5033,N_2805,N_3527);
xor U5034 (N_5034,N_3585,N_3678);
nand U5035 (N_5035,N_3401,N_3409);
nor U5036 (N_5036,N_3876,N_3640);
nor U5037 (N_5037,N_3188,N_3418);
xnor U5038 (N_5038,N_3533,N_3966);
nor U5039 (N_5039,N_2779,N_3590);
xnor U5040 (N_5040,N_2304,N_3239);
or U5041 (N_5041,N_2645,N_3867);
and U5042 (N_5042,N_2287,N_3660);
nand U5043 (N_5043,N_2966,N_2870);
and U5044 (N_5044,N_3309,N_3877);
nand U5045 (N_5045,N_2015,N_3022);
nor U5046 (N_5046,N_2569,N_2925);
and U5047 (N_5047,N_2490,N_3814);
and U5048 (N_5048,N_2157,N_3950);
xnor U5049 (N_5049,N_3426,N_3026);
or U5050 (N_5050,N_3973,N_3677);
nand U5051 (N_5051,N_2417,N_3179);
xnor U5052 (N_5052,N_3046,N_3716);
nand U5053 (N_5053,N_2972,N_2070);
nand U5054 (N_5054,N_3012,N_3382);
or U5055 (N_5055,N_2304,N_2175);
xor U5056 (N_5056,N_2855,N_2627);
and U5057 (N_5057,N_3061,N_2774);
or U5058 (N_5058,N_3938,N_2274);
nand U5059 (N_5059,N_2194,N_2567);
nor U5060 (N_5060,N_3220,N_2381);
nor U5061 (N_5061,N_3097,N_2609);
nor U5062 (N_5062,N_2461,N_3689);
and U5063 (N_5063,N_3404,N_3266);
or U5064 (N_5064,N_2185,N_2000);
xor U5065 (N_5065,N_2183,N_2990);
nor U5066 (N_5066,N_2556,N_2705);
or U5067 (N_5067,N_2708,N_2190);
xor U5068 (N_5068,N_2715,N_3910);
nand U5069 (N_5069,N_3332,N_2394);
xor U5070 (N_5070,N_3129,N_2944);
nor U5071 (N_5071,N_2916,N_3843);
xnor U5072 (N_5072,N_3700,N_2607);
nand U5073 (N_5073,N_2017,N_2167);
or U5074 (N_5074,N_3828,N_2909);
nand U5075 (N_5075,N_2002,N_3708);
and U5076 (N_5076,N_2817,N_2956);
or U5077 (N_5077,N_3321,N_2513);
nor U5078 (N_5078,N_3633,N_2539);
nor U5079 (N_5079,N_3626,N_3168);
nand U5080 (N_5080,N_2009,N_2501);
nor U5081 (N_5081,N_3903,N_2843);
or U5082 (N_5082,N_3426,N_2716);
nor U5083 (N_5083,N_3391,N_3957);
nand U5084 (N_5084,N_2753,N_3753);
nor U5085 (N_5085,N_3746,N_3449);
nor U5086 (N_5086,N_3906,N_2773);
xnor U5087 (N_5087,N_3107,N_2683);
or U5088 (N_5088,N_3191,N_2428);
or U5089 (N_5089,N_3481,N_2309);
nor U5090 (N_5090,N_3862,N_2477);
and U5091 (N_5091,N_2500,N_2528);
or U5092 (N_5092,N_2025,N_2786);
xor U5093 (N_5093,N_2433,N_3724);
or U5094 (N_5094,N_3817,N_2530);
and U5095 (N_5095,N_3494,N_2022);
or U5096 (N_5096,N_2623,N_3829);
xor U5097 (N_5097,N_2557,N_3368);
nor U5098 (N_5098,N_3963,N_3385);
and U5099 (N_5099,N_3307,N_3195);
and U5100 (N_5100,N_2370,N_2487);
nand U5101 (N_5101,N_3825,N_2566);
or U5102 (N_5102,N_3652,N_3624);
and U5103 (N_5103,N_3664,N_3957);
or U5104 (N_5104,N_2260,N_2808);
nand U5105 (N_5105,N_2573,N_3664);
nand U5106 (N_5106,N_2417,N_3635);
or U5107 (N_5107,N_2952,N_2950);
or U5108 (N_5108,N_3220,N_3978);
nand U5109 (N_5109,N_2024,N_2980);
xor U5110 (N_5110,N_3609,N_2873);
nand U5111 (N_5111,N_2964,N_3869);
and U5112 (N_5112,N_3898,N_3384);
xnor U5113 (N_5113,N_3326,N_2487);
nand U5114 (N_5114,N_3439,N_2532);
and U5115 (N_5115,N_3914,N_3102);
and U5116 (N_5116,N_2968,N_2497);
and U5117 (N_5117,N_2074,N_3384);
or U5118 (N_5118,N_3467,N_2864);
or U5119 (N_5119,N_3917,N_3695);
and U5120 (N_5120,N_3759,N_2344);
nor U5121 (N_5121,N_2791,N_3890);
or U5122 (N_5122,N_3852,N_3344);
nand U5123 (N_5123,N_3359,N_2344);
nand U5124 (N_5124,N_2200,N_3724);
and U5125 (N_5125,N_2402,N_2313);
nand U5126 (N_5126,N_2490,N_3805);
xnor U5127 (N_5127,N_3635,N_3884);
nand U5128 (N_5128,N_3347,N_2067);
and U5129 (N_5129,N_2165,N_2178);
nor U5130 (N_5130,N_3182,N_3606);
xor U5131 (N_5131,N_2199,N_2683);
nand U5132 (N_5132,N_3100,N_2644);
nor U5133 (N_5133,N_3999,N_2073);
nand U5134 (N_5134,N_2059,N_3976);
and U5135 (N_5135,N_2031,N_2795);
and U5136 (N_5136,N_2504,N_3772);
and U5137 (N_5137,N_3041,N_3791);
and U5138 (N_5138,N_3231,N_3168);
nand U5139 (N_5139,N_2779,N_3399);
or U5140 (N_5140,N_2777,N_2221);
nor U5141 (N_5141,N_2466,N_3439);
and U5142 (N_5142,N_2024,N_3197);
or U5143 (N_5143,N_3257,N_2739);
nor U5144 (N_5144,N_2585,N_2380);
nor U5145 (N_5145,N_3767,N_2989);
or U5146 (N_5146,N_2918,N_2867);
xnor U5147 (N_5147,N_2711,N_3949);
nor U5148 (N_5148,N_3123,N_3117);
nor U5149 (N_5149,N_2925,N_2826);
or U5150 (N_5150,N_3460,N_3699);
and U5151 (N_5151,N_2131,N_2182);
nor U5152 (N_5152,N_2957,N_3162);
nand U5153 (N_5153,N_3990,N_3658);
and U5154 (N_5154,N_3036,N_2005);
xor U5155 (N_5155,N_2935,N_2932);
xnor U5156 (N_5156,N_2011,N_2010);
and U5157 (N_5157,N_3853,N_2688);
nor U5158 (N_5158,N_3372,N_3317);
or U5159 (N_5159,N_3274,N_2479);
or U5160 (N_5160,N_3618,N_2958);
and U5161 (N_5161,N_2516,N_3997);
nand U5162 (N_5162,N_3830,N_2946);
and U5163 (N_5163,N_2484,N_3538);
nand U5164 (N_5164,N_2322,N_2582);
and U5165 (N_5165,N_2687,N_3567);
xnor U5166 (N_5166,N_3297,N_3248);
nand U5167 (N_5167,N_3785,N_2841);
nand U5168 (N_5168,N_3084,N_3604);
or U5169 (N_5169,N_2696,N_2988);
nand U5170 (N_5170,N_3516,N_2353);
and U5171 (N_5171,N_3860,N_2970);
or U5172 (N_5172,N_2769,N_3848);
nand U5173 (N_5173,N_3702,N_2864);
nand U5174 (N_5174,N_2946,N_2645);
nand U5175 (N_5175,N_3054,N_2902);
or U5176 (N_5176,N_3744,N_3901);
and U5177 (N_5177,N_3965,N_3646);
or U5178 (N_5178,N_2528,N_3956);
nor U5179 (N_5179,N_3462,N_2507);
and U5180 (N_5180,N_3219,N_3498);
xor U5181 (N_5181,N_2492,N_2077);
nand U5182 (N_5182,N_3358,N_3863);
nand U5183 (N_5183,N_2555,N_3694);
nand U5184 (N_5184,N_2709,N_3547);
nor U5185 (N_5185,N_2058,N_2021);
and U5186 (N_5186,N_2362,N_2496);
and U5187 (N_5187,N_2235,N_3629);
or U5188 (N_5188,N_2328,N_3342);
and U5189 (N_5189,N_3521,N_2593);
or U5190 (N_5190,N_2230,N_3149);
and U5191 (N_5191,N_2636,N_3322);
or U5192 (N_5192,N_2391,N_2749);
or U5193 (N_5193,N_2151,N_2693);
or U5194 (N_5194,N_3884,N_3899);
nor U5195 (N_5195,N_2133,N_2401);
nand U5196 (N_5196,N_2380,N_3650);
and U5197 (N_5197,N_2528,N_2716);
and U5198 (N_5198,N_3988,N_2844);
xor U5199 (N_5199,N_3863,N_2509);
or U5200 (N_5200,N_2239,N_2551);
and U5201 (N_5201,N_2083,N_2889);
and U5202 (N_5202,N_2824,N_2576);
and U5203 (N_5203,N_2559,N_3572);
nand U5204 (N_5204,N_2372,N_2497);
xnor U5205 (N_5205,N_3348,N_3663);
or U5206 (N_5206,N_3865,N_2813);
nor U5207 (N_5207,N_2102,N_2238);
and U5208 (N_5208,N_3650,N_2607);
nand U5209 (N_5209,N_3277,N_3505);
or U5210 (N_5210,N_2608,N_2170);
nand U5211 (N_5211,N_3907,N_3429);
nor U5212 (N_5212,N_3639,N_3356);
and U5213 (N_5213,N_2053,N_3798);
and U5214 (N_5214,N_2908,N_2976);
nor U5215 (N_5215,N_3321,N_2698);
nor U5216 (N_5216,N_2294,N_2867);
or U5217 (N_5217,N_2910,N_2341);
nand U5218 (N_5218,N_2569,N_3271);
nand U5219 (N_5219,N_2404,N_2594);
or U5220 (N_5220,N_2479,N_2572);
or U5221 (N_5221,N_2577,N_3069);
nand U5222 (N_5222,N_3080,N_3365);
and U5223 (N_5223,N_3662,N_2918);
xor U5224 (N_5224,N_2219,N_3524);
nor U5225 (N_5225,N_3527,N_3966);
and U5226 (N_5226,N_2394,N_2242);
or U5227 (N_5227,N_3452,N_3743);
or U5228 (N_5228,N_2648,N_3360);
or U5229 (N_5229,N_3905,N_2239);
nor U5230 (N_5230,N_3998,N_2280);
or U5231 (N_5231,N_2146,N_2103);
or U5232 (N_5232,N_3582,N_2135);
or U5233 (N_5233,N_3112,N_2205);
xor U5234 (N_5234,N_2350,N_2420);
nand U5235 (N_5235,N_3168,N_2819);
nand U5236 (N_5236,N_2010,N_2418);
nand U5237 (N_5237,N_3054,N_3540);
and U5238 (N_5238,N_3110,N_2789);
nand U5239 (N_5239,N_3744,N_3986);
or U5240 (N_5240,N_3952,N_2591);
or U5241 (N_5241,N_3776,N_2414);
xor U5242 (N_5242,N_3160,N_2178);
nor U5243 (N_5243,N_2065,N_3365);
nand U5244 (N_5244,N_3732,N_2368);
xor U5245 (N_5245,N_2931,N_2172);
nand U5246 (N_5246,N_2574,N_2815);
or U5247 (N_5247,N_2821,N_3998);
and U5248 (N_5248,N_2407,N_3619);
nand U5249 (N_5249,N_3642,N_3464);
nand U5250 (N_5250,N_2883,N_2021);
nor U5251 (N_5251,N_2811,N_2015);
nor U5252 (N_5252,N_2983,N_3908);
and U5253 (N_5253,N_3492,N_2719);
nor U5254 (N_5254,N_2193,N_2786);
nor U5255 (N_5255,N_3735,N_2091);
nand U5256 (N_5256,N_2215,N_3610);
xnor U5257 (N_5257,N_2671,N_3214);
xnor U5258 (N_5258,N_2944,N_2652);
nand U5259 (N_5259,N_2448,N_2909);
nor U5260 (N_5260,N_3586,N_2222);
and U5261 (N_5261,N_2919,N_3203);
xnor U5262 (N_5262,N_2387,N_2374);
nor U5263 (N_5263,N_3532,N_2294);
xor U5264 (N_5264,N_2563,N_3517);
or U5265 (N_5265,N_2715,N_2164);
nor U5266 (N_5266,N_3509,N_2866);
and U5267 (N_5267,N_3777,N_3436);
nand U5268 (N_5268,N_3662,N_2424);
or U5269 (N_5269,N_2511,N_3676);
and U5270 (N_5270,N_3642,N_3978);
or U5271 (N_5271,N_2205,N_3096);
and U5272 (N_5272,N_2869,N_2645);
xnor U5273 (N_5273,N_2698,N_3253);
nand U5274 (N_5274,N_3841,N_2991);
nand U5275 (N_5275,N_2227,N_3785);
and U5276 (N_5276,N_2936,N_2771);
and U5277 (N_5277,N_2713,N_2253);
or U5278 (N_5278,N_3876,N_2217);
nand U5279 (N_5279,N_2743,N_2270);
nand U5280 (N_5280,N_3972,N_3510);
or U5281 (N_5281,N_2359,N_2732);
or U5282 (N_5282,N_3588,N_2563);
and U5283 (N_5283,N_2965,N_2752);
and U5284 (N_5284,N_3666,N_2412);
or U5285 (N_5285,N_3373,N_3299);
xor U5286 (N_5286,N_3720,N_2891);
or U5287 (N_5287,N_2161,N_3067);
and U5288 (N_5288,N_3664,N_2788);
nor U5289 (N_5289,N_2699,N_3932);
or U5290 (N_5290,N_3224,N_2115);
or U5291 (N_5291,N_3226,N_2764);
or U5292 (N_5292,N_3421,N_3702);
nand U5293 (N_5293,N_2259,N_3209);
or U5294 (N_5294,N_3868,N_2463);
nor U5295 (N_5295,N_3599,N_3200);
nand U5296 (N_5296,N_3993,N_2663);
or U5297 (N_5297,N_3667,N_2821);
nand U5298 (N_5298,N_2835,N_2678);
nor U5299 (N_5299,N_2039,N_3279);
nor U5300 (N_5300,N_2713,N_3351);
nand U5301 (N_5301,N_3975,N_2822);
or U5302 (N_5302,N_2084,N_2461);
and U5303 (N_5303,N_3497,N_2856);
and U5304 (N_5304,N_2453,N_3642);
or U5305 (N_5305,N_3562,N_3315);
and U5306 (N_5306,N_2189,N_2938);
and U5307 (N_5307,N_2064,N_2278);
or U5308 (N_5308,N_2240,N_2848);
xor U5309 (N_5309,N_3323,N_3668);
xnor U5310 (N_5310,N_2795,N_3853);
or U5311 (N_5311,N_2132,N_3546);
nand U5312 (N_5312,N_2049,N_3751);
nand U5313 (N_5313,N_3339,N_2747);
xor U5314 (N_5314,N_3047,N_2424);
and U5315 (N_5315,N_3029,N_2426);
and U5316 (N_5316,N_2791,N_3757);
or U5317 (N_5317,N_3450,N_3585);
xor U5318 (N_5318,N_2812,N_2575);
nand U5319 (N_5319,N_2669,N_3009);
or U5320 (N_5320,N_2083,N_2184);
or U5321 (N_5321,N_3359,N_3221);
or U5322 (N_5322,N_2590,N_3352);
and U5323 (N_5323,N_3799,N_3292);
or U5324 (N_5324,N_2806,N_2340);
nand U5325 (N_5325,N_3305,N_3890);
xnor U5326 (N_5326,N_2512,N_3634);
nor U5327 (N_5327,N_2243,N_3857);
or U5328 (N_5328,N_3064,N_2484);
or U5329 (N_5329,N_3948,N_3564);
or U5330 (N_5330,N_2645,N_2073);
or U5331 (N_5331,N_3137,N_2954);
nand U5332 (N_5332,N_3790,N_2356);
and U5333 (N_5333,N_2705,N_2880);
or U5334 (N_5334,N_2490,N_2428);
xnor U5335 (N_5335,N_2232,N_2113);
or U5336 (N_5336,N_3164,N_2021);
nor U5337 (N_5337,N_2505,N_2124);
nand U5338 (N_5338,N_3369,N_3431);
or U5339 (N_5339,N_2281,N_2669);
nor U5340 (N_5340,N_3888,N_3237);
nor U5341 (N_5341,N_3758,N_2702);
nor U5342 (N_5342,N_3244,N_3092);
or U5343 (N_5343,N_2108,N_3616);
xnor U5344 (N_5344,N_3579,N_3496);
or U5345 (N_5345,N_2396,N_2514);
xnor U5346 (N_5346,N_2875,N_2789);
nor U5347 (N_5347,N_3227,N_3131);
xor U5348 (N_5348,N_3740,N_3889);
nand U5349 (N_5349,N_3899,N_2278);
nor U5350 (N_5350,N_2114,N_2317);
xnor U5351 (N_5351,N_2579,N_2990);
nor U5352 (N_5352,N_3751,N_2714);
nor U5353 (N_5353,N_3473,N_3609);
and U5354 (N_5354,N_3081,N_3003);
or U5355 (N_5355,N_2276,N_3126);
and U5356 (N_5356,N_2564,N_3879);
nand U5357 (N_5357,N_2880,N_3647);
and U5358 (N_5358,N_2660,N_2694);
nand U5359 (N_5359,N_2242,N_3234);
nor U5360 (N_5360,N_3586,N_3327);
and U5361 (N_5361,N_3868,N_3089);
nor U5362 (N_5362,N_3866,N_3844);
or U5363 (N_5363,N_3076,N_3266);
or U5364 (N_5364,N_2160,N_2306);
or U5365 (N_5365,N_2988,N_3445);
nand U5366 (N_5366,N_3976,N_3951);
nand U5367 (N_5367,N_2611,N_2364);
nor U5368 (N_5368,N_3512,N_2175);
and U5369 (N_5369,N_3549,N_3896);
and U5370 (N_5370,N_2491,N_3971);
or U5371 (N_5371,N_2983,N_3435);
nand U5372 (N_5372,N_3031,N_2101);
nor U5373 (N_5373,N_2429,N_2253);
and U5374 (N_5374,N_2294,N_2693);
or U5375 (N_5375,N_2388,N_2685);
and U5376 (N_5376,N_3788,N_2018);
or U5377 (N_5377,N_3838,N_3710);
nor U5378 (N_5378,N_2904,N_3963);
or U5379 (N_5379,N_2306,N_2892);
or U5380 (N_5380,N_2986,N_2236);
and U5381 (N_5381,N_2892,N_3024);
and U5382 (N_5382,N_3529,N_2218);
nor U5383 (N_5383,N_3178,N_3372);
nand U5384 (N_5384,N_2102,N_3373);
nand U5385 (N_5385,N_3394,N_2201);
nor U5386 (N_5386,N_2163,N_2124);
nand U5387 (N_5387,N_2313,N_2813);
and U5388 (N_5388,N_3983,N_3911);
or U5389 (N_5389,N_2036,N_3476);
and U5390 (N_5390,N_2831,N_3344);
nand U5391 (N_5391,N_2171,N_2360);
or U5392 (N_5392,N_3895,N_3200);
and U5393 (N_5393,N_3305,N_3419);
and U5394 (N_5394,N_3518,N_3770);
or U5395 (N_5395,N_2169,N_3892);
nor U5396 (N_5396,N_3070,N_3891);
or U5397 (N_5397,N_3749,N_3060);
nor U5398 (N_5398,N_3102,N_2263);
xor U5399 (N_5399,N_2966,N_2965);
nand U5400 (N_5400,N_3613,N_2549);
nand U5401 (N_5401,N_2619,N_2758);
and U5402 (N_5402,N_2387,N_2428);
and U5403 (N_5403,N_2656,N_2854);
or U5404 (N_5404,N_2846,N_2384);
nor U5405 (N_5405,N_2996,N_3994);
xnor U5406 (N_5406,N_3602,N_2884);
or U5407 (N_5407,N_2715,N_3307);
nor U5408 (N_5408,N_2076,N_3725);
or U5409 (N_5409,N_2422,N_3611);
or U5410 (N_5410,N_2964,N_2223);
nand U5411 (N_5411,N_2631,N_3503);
xnor U5412 (N_5412,N_3803,N_3740);
nand U5413 (N_5413,N_2590,N_2840);
nand U5414 (N_5414,N_2169,N_2275);
nand U5415 (N_5415,N_3236,N_3657);
nand U5416 (N_5416,N_2160,N_3682);
or U5417 (N_5417,N_3731,N_2294);
or U5418 (N_5418,N_3695,N_2020);
and U5419 (N_5419,N_3274,N_2763);
nor U5420 (N_5420,N_2584,N_3733);
nor U5421 (N_5421,N_3440,N_3713);
nor U5422 (N_5422,N_2757,N_2706);
nor U5423 (N_5423,N_3032,N_3239);
nor U5424 (N_5424,N_3318,N_3692);
nand U5425 (N_5425,N_2214,N_2261);
and U5426 (N_5426,N_3388,N_2914);
and U5427 (N_5427,N_3437,N_2225);
or U5428 (N_5428,N_3396,N_3815);
nand U5429 (N_5429,N_2366,N_2489);
nand U5430 (N_5430,N_2701,N_2886);
nor U5431 (N_5431,N_3508,N_2258);
or U5432 (N_5432,N_2550,N_2505);
and U5433 (N_5433,N_3442,N_3322);
nor U5434 (N_5434,N_3903,N_3065);
nor U5435 (N_5435,N_3132,N_2437);
nor U5436 (N_5436,N_2250,N_3524);
nor U5437 (N_5437,N_2146,N_3043);
and U5438 (N_5438,N_2616,N_3290);
xor U5439 (N_5439,N_2985,N_3389);
or U5440 (N_5440,N_3829,N_3308);
nand U5441 (N_5441,N_2390,N_3938);
nand U5442 (N_5442,N_2899,N_2280);
nor U5443 (N_5443,N_3435,N_2424);
and U5444 (N_5444,N_3352,N_3241);
nor U5445 (N_5445,N_2670,N_3600);
or U5446 (N_5446,N_3923,N_3429);
or U5447 (N_5447,N_2482,N_2336);
or U5448 (N_5448,N_3039,N_2010);
or U5449 (N_5449,N_3929,N_3234);
nor U5450 (N_5450,N_2410,N_3814);
or U5451 (N_5451,N_2027,N_2158);
nand U5452 (N_5452,N_2095,N_3470);
nand U5453 (N_5453,N_2757,N_3498);
or U5454 (N_5454,N_2518,N_3761);
or U5455 (N_5455,N_2503,N_3002);
nor U5456 (N_5456,N_3180,N_2463);
nor U5457 (N_5457,N_3525,N_3539);
or U5458 (N_5458,N_2684,N_2001);
xor U5459 (N_5459,N_3976,N_3143);
nand U5460 (N_5460,N_3373,N_2050);
and U5461 (N_5461,N_3816,N_2172);
nor U5462 (N_5462,N_3357,N_2423);
and U5463 (N_5463,N_2606,N_3492);
nand U5464 (N_5464,N_3556,N_3818);
nand U5465 (N_5465,N_3385,N_2484);
xor U5466 (N_5466,N_2733,N_2003);
or U5467 (N_5467,N_3050,N_2479);
nor U5468 (N_5468,N_2025,N_3287);
or U5469 (N_5469,N_3289,N_3738);
and U5470 (N_5470,N_2004,N_2556);
nand U5471 (N_5471,N_3979,N_3215);
or U5472 (N_5472,N_2606,N_2507);
nand U5473 (N_5473,N_2878,N_3220);
or U5474 (N_5474,N_2853,N_2257);
and U5475 (N_5475,N_2363,N_2913);
nand U5476 (N_5476,N_3081,N_2348);
and U5477 (N_5477,N_3623,N_3232);
or U5478 (N_5478,N_2207,N_2710);
and U5479 (N_5479,N_3558,N_3407);
xnor U5480 (N_5480,N_2157,N_2146);
and U5481 (N_5481,N_2313,N_3068);
nor U5482 (N_5482,N_3846,N_2590);
nand U5483 (N_5483,N_2558,N_3619);
nand U5484 (N_5484,N_3399,N_2528);
and U5485 (N_5485,N_2357,N_2290);
nor U5486 (N_5486,N_2278,N_2207);
or U5487 (N_5487,N_3010,N_3371);
nand U5488 (N_5488,N_3029,N_3462);
or U5489 (N_5489,N_2373,N_2811);
and U5490 (N_5490,N_2410,N_2387);
and U5491 (N_5491,N_2523,N_2209);
nand U5492 (N_5492,N_2824,N_2519);
nand U5493 (N_5493,N_3297,N_3625);
nand U5494 (N_5494,N_3531,N_3836);
nor U5495 (N_5495,N_3487,N_3416);
nand U5496 (N_5496,N_3058,N_2369);
nand U5497 (N_5497,N_2557,N_2947);
and U5498 (N_5498,N_2153,N_3209);
or U5499 (N_5499,N_3713,N_3967);
nand U5500 (N_5500,N_2079,N_2768);
or U5501 (N_5501,N_2045,N_2175);
and U5502 (N_5502,N_2448,N_2585);
nand U5503 (N_5503,N_2882,N_3088);
or U5504 (N_5504,N_3043,N_3615);
and U5505 (N_5505,N_2845,N_2045);
or U5506 (N_5506,N_2286,N_2745);
nor U5507 (N_5507,N_2502,N_2416);
nand U5508 (N_5508,N_2043,N_3537);
or U5509 (N_5509,N_2708,N_3536);
nand U5510 (N_5510,N_3738,N_2679);
and U5511 (N_5511,N_3195,N_2717);
or U5512 (N_5512,N_2481,N_3438);
nand U5513 (N_5513,N_3662,N_3620);
or U5514 (N_5514,N_2814,N_2638);
nor U5515 (N_5515,N_3177,N_3486);
nand U5516 (N_5516,N_2872,N_3878);
nand U5517 (N_5517,N_2759,N_2508);
and U5518 (N_5518,N_3615,N_2385);
and U5519 (N_5519,N_3283,N_2266);
and U5520 (N_5520,N_2255,N_3590);
or U5521 (N_5521,N_2071,N_2360);
and U5522 (N_5522,N_2935,N_2461);
or U5523 (N_5523,N_3532,N_3843);
and U5524 (N_5524,N_2976,N_2814);
nor U5525 (N_5525,N_2357,N_2261);
and U5526 (N_5526,N_3711,N_3684);
and U5527 (N_5527,N_3625,N_3180);
nor U5528 (N_5528,N_2654,N_2193);
nor U5529 (N_5529,N_3125,N_3765);
nor U5530 (N_5530,N_3795,N_2016);
nor U5531 (N_5531,N_3646,N_2213);
and U5532 (N_5532,N_2052,N_3040);
or U5533 (N_5533,N_3564,N_2233);
nor U5534 (N_5534,N_2549,N_2063);
nand U5535 (N_5535,N_2654,N_2232);
or U5536 (N_5536,N_2909,N_2446);
xor U5537 (N_5537,N_2287,N_2458);
or U5538 (N_5538,N_3057,N_3441);
nor U5539 (N_5539,N_3136,N_2263);
or U5540 (N_5540,N_3078,N_3162);
nand U5541 (N_5541,N_3540,N_2552);
and U5542 (N_5542,N_3581,N_3898);
nor U5543 (N_5543,N_3873,N_3602);
nor U5544 (N_5544,N_3251,N_2836);
nor U5545 (N_5545,N_3409,N_2238);
and U5546 (N_5546,N_2669,N_2690);
nor U5547 (N_5547,N_2518,N_3791);
nand U5548 (N_5548,N_2650,N_3142);
or U5549 (N_5549,N_2134,N_3368);
or U5550 (N_5550,N_3003,N_3258);
or U5551 (N_5551,N_2139,N_2049);
or U5552 (N_5552,N_2624,N_2218);
nand U5553 (N_5553,N_2625,N_3624);
xnor U5554 (N_5554,N_2667,N_2084);
nand U5555 (N_5555,N_3910,N_2023);
nand U5556 (N_5556,N_2944,N_3766);
nor U5557 (N_5557,N_2052,N_2128);
or U5558 (N_5558,N_2331,N_2216);
xor U5559 (N_5559,N_2233,N_2258);
and U5560 (N_5560,N_2598,N_3901);
nand U5561 (N_5561,N_2693,N_3339);
and U5562 (N_5562,N_2820,N_3554);
and U5563 (N_5563,N_3644,N_2026);
xnor U5564 (N_5564,N_2473,N_2509);
nor U5565 (N_5565,N_2643,N_2895);
and U5566 (N_5566,N_2226,N_3064);
and U5567 (N_5567,N_3760,N_3782);
nor U5568 (N_5568,N_2720,N_3538);
and U5569 (N_5569,N_3618,N_2871);
nor U5570 (N_5570,N_2395,N_2775);
nand U5571 (N_5571,N_3954,N_3555);
nor U5572 (N_5572,N_2197,N_2653);
and U5573 (N_5573,N_2971,N_2644);
or U5574 (N_5574,N_3824,N_2435);
nand U5575 (N_5575,N_2829,N_2018);
and U5576 (N_5576,N_3508,N_2038);
or U5577 (N_5577,N_3086,N_2386);
and U5578 (N_5578,N_2938,N_2921);
or U5579 (N_5579,N_3651,N_2196);
or U5580 (N_5580,N_2969,N_3968);
nor U5581 (N_5581,N_2498,N_3782);
nor U5582 (N_5582,N_3414,N_3395);
nand U5583 (N_5583,N_2610,N_3954);
or U5584 (N_5584,N_3040,N_3726);
nor U5585 (N_5585,N_3625,N_2369);
and U5586 (N_5586,N_2513,N_3128);
and U5587 (N_5587,N_2670,N_2338);
or U5588 (N_5588,N_3791,N_3459);
nor U5589 (N_5589,N_2523,N_2624);
and U5590 (N_5590,N_2366,N_3869);
and U5591 (N_5591,N_2609,N_3292);
or U5592 (N_5592,N_2990,N_2584);
nor U5593 (N_5593,N_3488,N_3243);
nor U5594 (N_5594,N_3321,N_3359);
nor U5595 (N_5595,N_2647,N_2968);
or U5596 (N_5596,N_2425,N_2074);
and U5597 (N_5597,N_2954,N_2239);
and U5598 (N_5598,N_2278,N_3438);
nor U5599 (N_5599,N_3146,N_2230);
nand U5600 (N_5600,N_3428,N_2845);
or U5601 (N_5601,N_2324,N_3960);
nor U5602 (N_5602,N_2789,N_2972);
nor U5603 (N_5603,N_3015,N_2358);
and U5604 (N_5604,N_3261,N_2214);
or U5605 (N_5605,N_2876,N_2539);
or U5606 (N_5606,N_2495,N_3589);
nand U5607 (N_5607,N_3729,N_2213);
nor U5608 (N_5608,N_2735,N_3262);
and U5609 (N_5609,N_2922,N_2246);
nor U5610 (N_5610,N_3029,N_3652);
nor U5611 (N_5611,N_3794,N_2430);
or U5612 (N_5612,N_3736,N_3555);
and U5613 (N_5613,N_2791,N_3009);
or U5614 (N_5614,N_3069,N_3835);
nor U5615 (N_5615,N_3440,N_3194);
or U5616 (N_5616,N_2206,N_3766);
or U5617 (N_5617,N_3815,N_2641);
and U5618 (N_5618,N_2336,N_2833);
or U5619 (N_5619,N_2352,N_3622);
or U5620 (N_5620,N_3934,N_3605);
xnor U5621 (N_5621,N_3695,N_2327);
nor U5622 (N_5622,N_2964,N_2185);
nand U5623 (N_5623,N_3077,N_2763);
or U5624 (N_5624,N_2042,N_2117);
nor U5625 (N_5625,N_2608,N_2780);
nor U5626 (N_5626,N_2275,N_2362);
and U5627 (N_5627,N_3113,N_2601);
nor U5628 (N_5628,N_3965,N_2845);
nand U5629 (N_5629,N_3125,N_3454);
or U5630 (N_5630,N_3875,N_2705);
nand U5631 (N_5631,N_3652,N_3547);
nor U5632 (N_5632,N_2800,N_2986);
nor U5633 (N_5633,N_2625,N_3831);
nand U5634 (N_5634,N_3038,N_2810);
and U5635 (N_5635,N_2827,N_3672);
nor U5636 (N_5636,N_3536,N_2984);
and U5637 (N_5637,N_2259,N_2455);
xor U5638 (N_5638,N_2546,N_2600);
and U5639 (N_5639,N_2431,N_2630);
and U5640 (N_5640,N_2860,N_2038);
or U5641 (N_5641,N_3022,N_2754);
and U5642 (N_5642,N_3079,N_2917);
and U5643 (N_5643,N_3624,N_2050);
nor U5644 (N_5644,N_3678,N_2938);
xnor U5645 (N_5645,N_3686,N_2641);
nand U5646 (N_5646,N_3454,N_2399);
nor U5647 (N_5647,N_3180,N_2821);
nor U5648 (N_5648,N_2430,N_2574);
and U5649 (N_5649,N_3948,N_3084);
nand U5650 (N_5650,N_2164,N_2267);
and U5651 (N_5651,N_2608,N_3051);
nor U5652 (N_5652,N_3530,N_3632);
nor U5653 (N_5653,N_3141,N_2839);
nand U5654 (N_5654,N_3730,N_2165);
nor U5655 (N_5655,N_2262,N_2104);
and U5656 (N_5656,N_2004,N_2349);
nand U5657 (N_5657,N_2652,N_3088);
nor U5658 (N_5658,N_2127,N_3487);
or U5659 (N_5659,N_3132,N_2841);
or U5660 (N_5660,N_3304,N_3049);
nor U5661 (N_5661,N_2029,N_3336);
and U5662 (N_5662,N_3998,N_3451);
nand U5663 (N_5663,N_2466,N_2556);
xor U5664 (N_5664,N_3337,N_3175);
or U5665 (N_5665,N_3936,N_2014);
nand U5666 (N_5666,N_3802,N_3944);
nor U5667 (N_5667,N_3122,N_3022);
xnor U5668 (N_5668,N_3457,N_2377);
nand U5669 (N_5669,N_2993,N_3885);
and U5670 (N_5670,N_2026,N_2158);
nand U5671 (N_5671,N_3741,N_3502);
nor U5672 (N_5672,N_2692,N_2223);
nand U5673 (N_5673,N_2996,N_2541);
and U5674 (N_5674,N_2694,N_2414);
nor U5675 (N_5675,N_3619,N_2329);
or U5676 (N_5676,N_2767,N_2910);
nand U5677 (N_5677,N_2839,N_3130);
nand U5678 (N_5678,N_2621,N_3398);
nor U5679 (N_5679,N_2049,N_2494);
or U5680 (N_5680,N_3926,N_3325);
nor U5681 (N_5681,N_3161,N_3882);
nor U5682 (N_5682,N_3066,N_3161);
nand U5683 (N_5683,N_2525,N_3166);
and U5684 (N_5684,N_3331,N_2634);
or U5685 (N_5685,N_3478,N_2989);
and U5686 (N_5686,N_2970,N_2757);
and U5687 (N_5687,N_2225,N_2648);
or U5688 (N_5688,N_3195,N_2716);
and U5689 (N_5689,N_3376,N_2716);
or U5690 (N_5690,N_2846,N_2508);
or U5691 (N_5691,N_3733,N_2856);
nand U5692 (N_5692,N_2423,N_3602);
nor U5693 (N_5693,N_3482,N_2493);
nor U5694 (N_5694,N_3511,N_3989);
or U5695 (N_5695,N_3285,N_2914);
or U5696 (N_5696,N_3776,N_3721);
nor U5697 (N_5697,N_3460,N_3091);
and U5698 (N_5698,N_3709,N_2030);
xor U5699 (N_5699,N_2208,N_3103);
nand U5700 (N_5700,N_2292,N_2406);
nor U5701 (N_5701,N_2242,N_3330);
nor U5702 (N_5702,N_3930,N_2460);
nor U5703 (N_5703,N_3036,N_2492);
nand U5704 (N_5704,N_2087,N_3297);
or U5705 (N_5705,N_3590,N_3573);
and U5706 (N_5706,N_2063,N_2333);
and U5707 (N_5707,N_3180,N_2020);
nor U5708 (N_5708,N_2165,N_2309);
nor U5709 (N_5709,N_3435,N_2388);
and U5710 (N_5710,N_2643,N_2070);
nand U5711 (N_5711,N_3588,N_3776);
and U5712 (N_5712,N_2433,N_2127);
nand U5713 (N_5713,N_3075,N_3430);
nand U5714 (N_5714,N_3704,N_3001);
and U5715 (N_5715,N_3326,N_3514);
and U5716 (N_5716,N_3560,N_2561);
xnor U5717 (N_5717,N_3907,N_3127);
nand U5718 (N_5718,N_2690,N_2116);
nand U5719 (N_5719,N_2306,N_3006);
nand U5720 (N_5720,N_2443,N_2313);
and U5721 (N_5721,N_3369,N_2385);
xor U5722 (N_5722,N_2595,N_3982);
xnor U5723 (N_5723,N_2502,N_3301);
xor U5724 (N_5724,N_3143,N_3674);
or U5725 (N_5725,N_3697,N_2330);
nor U5726 (N_5726,N_3388,N_2869);
nor U5727 (N_5727,N_2025,N_2941);
or U5728 (N_5728,N_2986,N_3542);
nand U5729 (N_5729,N_3647,N_3955);
and U5730 (N_5730,N_2511,N_2093);
nor U5731 (N_5731,N_3483,N_3327);
nor U5732 (N_5732,N_2473,N_2772);
and U5733 (N_5733,N_2791,N_2702);
xnor U5734 (N_5734,N_2882,N_3918);
nor U5735 (N_5735,N_3951,N_3067);
or U5736 (N_5736,N_2131,N_2286);
nand U5737 (N_5737,N_3638,N_3853);
nor U5738 (N_5738,N_3540,N_2672);
nand U5739 (N_5739,N_2810,N_3820);
or U5740 (N_5740,N_3719,N_2637);
nor U5741 (N_5741,N_3388,N_2382);
xnor U5742 (N_5742,N_3331,N_2082);
and U5743 (N_5743,N_3726,N_3987);
nor U5744 (N_5744,N_2491,N_3661);
nand U5745 (N_5745,N_2758,N_2186);
nor U5746 (N_5746,N_2254,N_2827);
nor U5747 (N_5747,N_2326,N_3185);
xnor U5748 (N_5748,N_3603,N_3122);
nor U5749 (N_5749,N_2498,N_3015);
nor U5750 (N_5750,N_3898,N_3648);
and U5751 (N_5751,N_3933,N_3224);
nor U5752 (N_5752,N_2651,N_2611);
or U5753 (N_5753,N_2366,N_2297);
or U5754 (N_5754,N_3860,N_2874);
or U5755 (N_5755,N_2919,N_2325);
nand U5756 (N_5756,N_2307,N_3214);
or U5757 (N_5757,N_2265,N_2809);
and U5758 (N_5758,N_3300,N_2273);
nand U5759 (N_5759,N_3281,N_3635);
nor U5760 (N_5760,N_2679,N_3234);
nor U5761 (N_5761,N_2767,N_3998);
xnor U5762 (N_5762,N_3135,N_2702);
nand U5763 (N_5763,N_2264,N_2628);
nor U5764 (N_5764,N_2953,N_2769);
or U5765 (N_5765,N_2082,N_3437);
nor U5766 (N_5766,N_3511,N_3466);
nand U5767 (N_5767,N_2474,N_3139);
nor U5768 (N_5768,N_2193,N_3250);
or U5769 (N_5769,N_2211,N_2201);
nor U5770 (N_5770,N_2096,N_3758);
nor U5771 (N_5771,N_2254,N_3240);
or U5772 (N_5772,N_2748,N_2889);
xor U5773 (N_5773,N_2039,N_2671);
or U5774 (N_5774,N_3660,N_2124);
xnor U5775 (N_5775,N_2721,N_2879);
nand U5776 (N_5776,N_2101,N_2140);
nand U5777 (N_5777,N_3456,N_2697);
nand U5778 (N_5778,N_2628,N_2400);
nand U5779 (N_5779,N_2711,N_3380);
nor U5780 (N_5780,N_2519,N_2654);
and U5781 (N_5781,N_3861,N_2386);
nand U5782 (N_5782,N_2928,N_2465);
nor U5783 (N_5783,N_3572,N_3993);
nor U5784 (N_5784,N_3658,N_2621);
nand U5785 (N_5785,N_2077,N_2479);
or U5786 (N_5786,N_2441,N_3461);
nand U5787 (N_5787,N_2948,N_3712);
or U5788 (N_5788,N_3674,N_3948);
and U5789 (N_5789,N_3046,N_3852);
or U5790 (N_5790,N_3371,N_2253);
nand U5791 (N_5791,N_3757,N_3292);
nand U5792 (N_5792,N_3578,N_3619);
and U5793 (N_5793,N_3355,N_3661);
xor U5794 (N_5794,N_2103,N_3912);
or U5795 (N_5795,N_2721,N_2618);
nor U5796 (N_5796,N_3854,N_3229);
and U5797 (N_5797,N_2996,N_2110);
nand U5798 (N_5798,N_3191,N_3488);
and U5799 (N_5799,N_2120,N_2152);
nand U5800 (N_5800,N_3273,N_3753);
and U5801 (N_5801,N_2175,N_3805);
nand U5802 (N_5802,N_2318,N_3689);
nor U5803 (N_5803,N_2878,N_2202);
nand U5804 (N_5804,N_2137,N_2701);
nand U5805 (N_5805,N_3240,N_2932);
nand U5806 (N_5806,N_2967,N_2840);
nand U5807 (N_5807,N_2480,N_3754);
nor U5808 (N_5808,N_3802,N_2808);
nand U5809 (N_5809,N_3969,N_2282);
or U5810 (N_5810,N_3100,N_2607);
and U5811 (N_5811,N_2782,N_2194);
or U5812 (N_5812,N_2229,N_3749);
or U5813 (N_5813,N_3973,N_3753);
nor U5814 (N_5814,N_3476,N_3302);
nor U5815 (N_5815,N_3150,N_2949);
nand U5816 (N_5816,N_2889,N_3766);
or U5817 (N_5817,N_3274,N_2481);
nand U5818 (N_5818,N_3382,N_2140);
nor U5819 (N_5819,N_3960,N_2645);
nand U5820 (N_5820,N_2811,N_3469);
or U5821 (N_5821,N_2517,N_3024);
and U5822 (N_5822,N_2575,N_2973);
nand U5823 (N_5823,N_3064,N_2771);
nor U5824 (N_5824,N_3766,N_3032);
and U5825 (N_5825,N_2742,N_2073);
and U5826 (N_5826,N_2689,N_2283);
or U5827 (N_5827,N_2877,N_2463);
and U5828 (N_5828,N_2607,N_3687);
and U5829 (N_5829,N_2674,N_2020);
nand U5830 (N_5830,N_2073,N_2724);
nor U5831 (N_5831,N_2945,N_2841);
nand U5832 (N_5832,N_2739,N_2400);
nor U5833 (N_5833,N_3914,N_2642);
or U5834 (N_5834,N_2201,N_2516);
or U5835 (N_5835,N_2691,N_2222);
nand U5836 (N_5836,N_3209,N_2394);
nand U5837 (N_5837,N_2416,N_3374);
nor U5838 (N_5838,N_2621,N_3259);
or U5839 (N_5839,N_2598,N_3904);
nor U5840 (N_5840,N_2120,N_3030);
nor U5841 (N_5841,N_2802,N_3649);
nor U5842 (N_5842,N_3209,N_2360);
nand U5843 (N_5843,N_2029,N_2500);
or U5844 (N_5844,N_2805,N_3113);
xnor U5845 (N_5845,N_2323,N_3257);
nor U5846 (N_5846,N_2378,N_2337);
nor U5847 (N_5847,N_3483,N_3500);
and U5848 (N_5848,N_3795,N_3431);
or U5849 (N_5849,N_3428,N_3967);
and U5850 (N_5850,N_3910,N_3247);
nor U5851 (N_5851,N_3153,N_2134);
and U5852 (N_5852,N_2260,N_3543);
or U5853 (N_5853,N_2239,N_2504);
nand U5854 (N_5854,N_3344,N_3264);
or U5855 (N_5855,N_3096,N_3862);
nor U5856 (N_5856,N_2010,N_2436);
nand U5857 (N_5857,N_3142,N_3204);
nand U5858 (N_5858,N_3549,N_2550);
xor U5859 (N_5859,N_3237,N_3454);
xor U5860 (N_5860,N_2282,N_2850);
and U5861 (N_5861,N_2007,N_2675);
xnor U5862 (N_5862,N_3786,N_3101);
and U5863 (N_5863,N_3037,N_2902);
and U5864 (N_5864,N_2291,N_3217);
and U5865 (N_5865,N_2457,N_3864);
and U5866 (N_5866,N_3407,N_3967);
xor U5867 (N_5867,N_3203,N_2998);
nor U5868 (N_5868,N_3988,N_2528);
or U5869 (N_5869,N_3639,N_3421);
nor U5870 (N_5870,N_3297,N_3819);
nor U5871 (N_5871,N_2874,N_3258);
or U5872 (N_5872,N_3850,N_2895);
nand U5873 (N_5873,N_3699,N_3828);
nand U5874 (N_5874,N_3411,N_3661);
or U5875 (N_5875,N_2694,N_3617);
or U5876 (N_5876,N_3917,N_3723);
or U5877 (N_5877,N_3517,N_2328);
xnor U5878 (N_5878,N_2738,N_3217);
nor U5879 (N_5879,N_2358,N_3228);
nor U5880 (N_5880,N_3713,N_3836);
or U5881 (N_5881,N_3415,N_3783);
nor U5882 (N_5882,N_3918,N_3023);
and U5883 (N_5883,N_3735,N_2276);
xor U5884 (N_5884,N_2402,N_2853);
and U5885 (N_5885,N_3583,N_2449);
or U5886 (N_5886,N_2162,N_3225);
nand U5887 (N_5887,N_2790,N_3582);
nor U5888 (N_5888,N_2736,N_3738);
or U5889 (N_5889,N_3027,N_2527);
or U5890 (N_5890,N_2713,N_2287);
nor U5891 (N_5891,N_3388,N_2187);
xor U5892 (N_5892,N_3698,N_2990);
nor U5893 (N_5893,N_2662,N_3747);
xor U5894 (N_5894,N_3973,N_2065);
xor U5895 (N_5895,N_3241,N_3236);
nand U5896 (N_5896,N_3203,N_2714);
nand U5897 (N_5897,N_3024,N_3403);
and U5898 (N_5898,N_2217,N_2737);
nand U5899 (N_5899,N_3221,N_2863);
nand U5900 (N_5900,N_3192,N_2248);
and U5901 (N_5901,N_2019,N_3546);
nor U5902 (N_5902,N_3275,N_3933);
nand U5903 (N_5903,N_3490,N_2651);
nor U5904 (N_5904,N_3500,N_2596);
nor U5905 (N_5905,N_3420,N_2973);
nor U5906 (N_5906,N_3618,N_3153);
nand U5907 (N_5907,N_2256,N_3363);
or U5908 (N_5908,N_3679,N_3976);
nand U5909 (N_5909,N_3487,N_3840);
nor U5910 (N_5910,N_3232,N_3889);
xor U5911 (N_5911,N_3864,N_2902);
nor U5912 (N_5912,N_2291,N_3913);
or U5913 (N_5913,N_2665,N_2137);
nand U5914 (N_5914,N_3815,N_3689);
nand U5915 (N_5915,N_2098,N_3183);
and U5916 (N_5916,N_3010,N_2488);
and U5917 (N_5917,N_2356,N_2564);
and U5918 (N_5918,N_3464,N_3852);
nor U5919 (N_5919,N_3216,N_2952);
or U5920 (N_5920,N_3309,N_3468);
nor U5921 (N_5921,N_3964,N_3527);
nor U5922 (N_5922,N_2659,N_3522);
nand U5923 (N_5923,N_2312,N_2065);
nand U5924 (N_5924,N_3896,N_2259);
nor U5925 (N_5925,N_2408,N_2329);
or U5926 (N_5926,N_2406,N_2714);
or U5927 (N_5927,N_3287,N_2023);
or U5928 (N_5928,N_3931,N_2143);
nand U5929 (N_5929,N_3935,N_2535);
or U5930 (N_5930,N_2725,N_2445);
nor U5931 (N_5931,N_2253,N_2107);
and U5932 (N_5932,N_3850,N_2535);
or U5933 (N_5933,N_3964,N_3586);
nor U5934 (N_5934,N_2325,N_3362);
and U5935 (N_5935,N_2380,N_2106);
or U5936 (N_5936,N_3202,N_2273);
or U5937 (N_5937,N_3859,N_3295);
nor U5938 (N_5938,N_2019,N_2020);
nor U5939 (N_5939,N_2384,N_2079);
or U5940 (N_5940,N_3256,N_3162);
xor U5941 (N_5941,N_3581,N_2094);
nor U5942 (N_5942,N_2804,N_3737);
nor U5943 (N_5943,N_2844,N_2732);
nand U5944 (N_5944,N_3050,N_2919);
nor U5945 (N_5945,N_3526,N_2683);
or U5946 (N_5946,N_3382,N_2478);
nand U5947 (N_5947,N_2468,N_2994);
nor U5948 (N_5948,N_3536,N_3062);
xnor U5949 (N_5949,N_2735,N_2141);
and U5950 (N_5950,N_3793,N_2703);
and U5951 (N_5951,N_2953,N_3606);
nor U5952 (N_5952,N_3337,N_3999);
and U5953 (N_5953,N_3657,N_3535);
and U5954 (N_5954,N_2184,N_2727);
or U5955 (N_5955,N_2333,N_3673);
nor U5956 (N_5956,N_3991,N_3402);
or U5957 (N_5957,N_3503,N_3041);
nor U5958 (N_5958,N_3698,N_3104);
and U5959 (N_5959,N_2548,N_3591);
and U5960 (N_5960,N_3922,N_2430);
and U5961 (N_5961,N_2991,N_3165);
nor U5962 (N_5962,N_3941,N_2277);
nor U5963 (N_5963,N_3928,N_3193);
and U5964 (N_5964,N_3532,N_3067);
and U5965 (N_5965,N_3336,N_3032);
nor U5966 (N_5966,N_2760,N_2075);
or U5967 (N_5967,N_2272,N_2529);
and U5968 (N_5968,N_3610,N_2475);
nor U5969 (N_5969,N_2716,N_3744);
nor U5970 (N_5970,N_2297,N_2980);
nor U5971 (N_5971,N_3959,N_2989);
and U5972 (N_5972,N_3992,N_3951);
and U5973 (N_5973,N_2994,N_3572);
xor U5974 (N_5974,N_2572,N_2093);
or U5975 (N_5975,N_3246,N_3239);
xor U5976 (N_5976,N_3777,N_3341);
and U5977 (N_5977,N_3536,N_3603);
or U5978 (N_5978,N_2731,N_3182);
nand U5979 (N_5979,N_2549,N_2143);
nand U5980 (N_5980,N_2962,N_2475);
nor U5981 (N_5981,N_2559,N_2086);
and U5982 (N_5982,N_2232,N_2052);
nand U5983 (N_5983,N_3160,N_2285);
or U5984 (N_5984,N_2865,N_2661);
nor U5985 (N_5985,N_2696,N_3610);
or U5986 (N_5986,N_2006,N_3716);
nand U5987 (N_5987,N_3179,N_3214);
nand U5988 (N_5988,N_3323,N_3725);
xor U5989 (N_5989,N_3476,N_3861);
and U5990 (N_5990,N_3390,N_3828);
xor U5991 (N_5991,N_2503,N_3865);
xor U5992 (N_5992,N_2453,N_2000);
and U5993 (N_5993,N_3743,N_3433);
nand U5994 (N_5994,N_2341,N_3725);
nor U5995 (N_5995,N_3165,N_3478);
or U5996 (N_5996,N_3641,N_2185);
nor U5997 (N_5997,N_2377,N_2972);
or U5998 (N_5998,N_3027,N_3025);
or U5999 (N_5999,N_2578,N_3485);
nor U6000 (N_6000,N_5248,N_5889);
nand U6001 (N_6001,N_5796,N_4776);
nor U6002 (N_6002,N_4275,N_5491);
nor U6003 (N_6003,N_4550,N_5792);
nand U6004 (N_6004,N_4520,N_4552);
nor U6005 (N_6005,N_4245,N_5830);
and U6006 (N_6006,N_5892,N_4518);
nor U6007 (N_6007,N_4419,N_5442);
nand U6008 (N_6008,N_5974,N_5269);
nand U6009 (N_6009,N_5591,N_5584);
xnor U6010 (N_6010,N_5682,N_5083);
or U6011 (N_6011,N_4535,N_5639);
nand U6012 (N_6012,N_4965,N_5913);
or U6013 (N_6013,N_4272,N_4584);
or U6014 (N_6014,N_5699,N_4841);
xor U6015 (N_6015,N_5355,N_5462);
nand U6016 (N_6016,N_4363,N_4753);
nor U6017 (N_6017,N_4096,N_5262);
or U6018 (N_6018,N_4129,N_4823);
and U6019 (N_6019,N_5800,N_5039);
or U6020 (N_6020,N_5516,N_5423);
nand U6021 (N_6021,N_4205,N_5100);
and U6022 (N_6022,N_5858,N_4058);
or U6023 (N_6023,N_4767,N_4549);
or U6024 (N_6024,N_5606,N_4143);
and U6025 (N_6025,N_5898,N_4571);
and U6026 (N_6026,N_5928,N_5727);
nor U6027 (N_6027,N_5365,N_5581);
nor U6028 (N_6028,N_4446,N_4087);
or U6029 (N_6029,N_4863,N_5971);
or U6030 (N_6030,N_4751,N_4404);
or U6031 (N_6031,N_4850,N_4531);
and U6032 (N_6032,N_5709,N_4939);
or U6033 (N_6033,N_5176,N_5774);
nand U6034 (N_6034,N_4542,N_4881);
nand U6035 (N_6035,N_4544,N_4144);
and U6036 (N_6036,N_4632,N_5067);
nand U6037 (N_6037,N_5945,N_5143);
nand U6038 (N_6038,N_4166,N_5424);
nand U6039 (N_6039,N_5759,N_4391);
nor U6040 (N_6040,N_5099,N_4495);
and U6041 (N_6041,N_5032,N_5194);
nor U6042 (N_6042,N_5702,N_5228);
nor U6043 (N_6043,N_5133,N_4278);
nor U6044 (N_6044,N_5661,N_4546);
nor U6045 (N_6045,N_5287,N_4053);
or U6046 (N_6046,N_5401,N_5022);
and U6047 (N_6047,N_5354,N_5327);
nand U6048 (N_6048,N_4007,N_5824);
xnor U6049 (N_6049,N_5587,N_5998);
or U6050 (N_6050,N_5562,N_4161);
nor U6051 (N_6051,N_4516,N_5125);
or U6052 (N_6052,N_4106,N_5675);
and U6053 (N_6053,N_4742,N_4985);
nor U6054 (N_6054,N_4423,N_5542);
and U6055 (N_6055,N_5166,N_5923);
and U6056 (N_6056,N_4757,N_5184);
nor U6057 (N_6057,N_5001,N_5488);
nor U6058 (N_6058,N_5225,N_5174);
or U6059 (N_6059,N_4226,N_5382);
xor U6060 (N_6060,N_4813,N_5209);
nand U6061 (N_6061,N_5130,N_5086);
xnor U6062 (N_6062,N_5038,N_4557);
and U6063 (N_6063,N_5873,N_4315);
or U6064 (N_6064,N_4020,N_4728);
or U6065 (N_6065,N_4924,N_5441);
nor U6066 (N_6066,N_5627,N_4147);
or U6067 (N_6067,N_5876,N_5852);
or U6068 (N_6068,N_5255,N_4054);
or U6069 (N_6069,N_5033,N_4969);
nand U6070 (N_6070,N_5743,N_5806);
and U6071 (N_6071,N_5678,N_4194);
and U6072 (N_6072,N_5929,N_5805);
or U6073 (N_6073,N_5741,N_4121);
nand U6074 (N_6074,N_4987,N_4956);
nand U6075 (N_6075,N_5358,N_5633);
or U6076 (N_6076,N_4216,N_4729);
and U6077 (N_6077,N_5050,N_4442);
nor U6078 (N_6078,N_4907,N_5431);
nand U6079 (N_6079,N_4262,N_4597);
and U6080 (N_6080,N_5908,N_4598);
nor U6081 (N_6081,N_4429,N_5791);
or U6082 (N_6082,N_5549,N_5981);
or U6083 (N_6083,N_4665,N_5839);
xor U6084 (N_6084,N_5959,N_5289);
and U6085 (N_6085,N_5245,N_5295);
or U6086 (N_6086,N_5626,N_5781);
or U6087 (N_6087,N_5135,N_5906);
nand U6088 (N_6088,N_5106,N_5413);
nor U6089 (N_6089,N_4893,N_5965);
and U6090 (N_6090,N_4803,N_4354);
nor U6091 (N_6091,N_5617,N_5217);
and U6092 (N_6092,N_4524,N_5416);
nand U6093 (N_6093,N_5063,N_4876);
nand U6094 (N_6094,N_5089,N_4156);
or U6095 (N_6095,N_4328,N_5250);
or U6096 (N_6096,N_5241,N_5771);
xnor U6097 (N_6097,N_4212,N_4703);
or U6098 (N_6098,N_5676,N_4569);
and U6099 (N_6099,N_4393,N_4774);
nand U6100 (N_6100,N_5569,N_4739);
xor U6101 (N_6101,N_5218,N_4478);
and U6102 (N_6102,N_4555,N_4621);
nand U6103 (N_6103,N_5803,N_4130);
nand U6104 (N_6104,N_5234,N_5211);
or U6105 (N_6105,N_5614,N_5812);
nand U6106 (N_6106,N_5943,N_5762);
and U6107 (N_6107,N_4692,N_5470);
xnor U6108 (N_6108,N_5304,N_5527);
nand U6109 (N_6109,N_4910,N_4761);
and U6110 (N_6110,N_4829,N_4459);
or U6111 (N_6111,N_4000,N_4292);
xor U6112 (N_6112,N_4438,N_5153);
or U6113 (N_6113,N_4983,N_5685);
or U6114 (N_6114,N_4668,N_4947);
nand U6115 (N_6115,N_5119,N_4655);
or U6116 (N_6116,N_5026,N_4826);
or U6117 (N_6117,N_4341,N_5132);
nand U6118 (N_6118,N_5029,N_5095);
nor U6119 (N_6119,N_4385,N_4526);
nand U6120 (N_6120,N_5126,N_5819);
or U6121 (N_6121,N_5129,N_4406);
nand U6122 (N_6122,N_5979,N_5170);
or U6123 (N_6123,N_5880,N_4674);
or U6124 (N_6124,N_5392,N_5473);
nor U6125 (N_6125,N_4968,N_5318);
nand U6126 (N_6126,N_5668,N_4502);
nor U6127 (N_6127,N_4172,N_4136);
nand U6128 (N_6128,N_4624,N_4101);
and U6129 (N_6129,N_5875,N_5298);
and U6130 (N_6130,N_5993,N_4013);
or U6131 (N_6131,N_5193,N_4330);
or U6132 (N_6132,N_4326,N_5565);
nor U6133 (N_6133,N_5109,N_4709);
xor U6134 (N_6134,N_5673,N_4426);
and U6135 (N_6135,N_4783,N_5181);
and U6136 (N_6136,N_5897,N_4248);
nor U6137 (N_6137,N_4891,N_5788);
nand U6138 (N_6138,N_5911,N_4455);
nor U6139 (N_6139,N_5256,N_4022);
nor U6140 (N_6140,N_4199,N_4937);
nand U6141 (N_6141,N_5249,N_4859);
nor U6142 (N_6142,N_4238,N_4119);
nor U6143 (N_6143,N_5749,N_5813);
nand U6144 (N_6144,N_4862,N_5436);
or U6145 (N_6145,N_4168,N_4439);
nand U6146 (N_6146,N_5932,N_5016);
xor U6147 (N_6147,N_4333,N_4152);
nand U6148 (N_6148,N_5021,N_5294);
or U6149 (N_6149,N_4998,N_5058);
nor U6150 (N_6150,N_5122,N_4454);
nor U6151 (N_6151,N_5780,N_4314);
and U6152 (N_6152,N_5448,N_4795);
and U6153 (N_6153,N_4941,N_5237);
and U6154 (N_6154,N_5097,N_4900);
and U6155 (N_6155,N_4425,N_5390);
and U6156 (N_6156,N_4160,N_5112);
nand U6157 (N_6157,N_4277,N_4734);
or U6158 (N_6158,N_5013,N_4599);
or U6159 (N_6159,N_5550,N_4094);
and U6160 (N_6160,N_4573,N_4180);
xor U6161 (N_6161,N_4801,N_4304);
and U6162 (N_6162,N_4722,N_4055);
nor U6163 (N_6163,N_4320,N_5272);
or U6164 (N_6164,N_5487,N_5758);
nor U6165 (N_6165,N_4828,N_5251);
nand U6166 (N_6166,N_5017,N_5930);
nor U6167 (N_6167,N_5007,N_4731);
nand U6168 (N_6168,N_5235,N_4994);
or U6169 (N_6169,N_4435,N_5994);
and U6170 (N_6170,N_4636,N_5964);
nand U6171 (N_6171,N_4580,N_4352);
or U6172 (N_6172,N_5395,N_4892);
or U6173 (N_6173,N_5629,N_4733);
nor U6174 (N_6174,N_5656,N_4511);
and U6175 (N_6175,N_4456,N_4611);
or U6176 (N_6176,N_5275,N_4851);
or U6177 (N_6177,N_4360,N_4149);
nand U6178 (N_6178,N_4268,N_4402);
xor U6179 (N_6179,N_5389,N_4252);
nor U6180 (N_6180,N_5385,N_5090);
nor U6181 (N_6181,N_4556,N_5212);
or U6182 (N_6182,N_4752,N_4362);
xor U6183 (N_6183,N_4128,N_5798);
xnor U6184 (N_6184,N_4564,N_4612);
or U6185 (N_6185,N_4817,N_5185);
nand U6186 (N_6186,N_5186,N_5331);
and U6187 (N_6187,N_4650,N_4291);
and U6188 (N_6188,N_5522,N_5918);
xnor U6189 (N_6189,N_5443,N_5620);
nor U6190 (N_6190,N_4297,N_5207);
or U6191 (N_6191,N_4343,N_5432);
or U6192 (N_6192,N_5836,N_5474);
or U6193 (N_6193,N_4035,N_5040);
and U6194 (N_6194,N_5430,N_5794);
nand U6195 (N_6195,N_5146,N_4713);
and U6196 (N_6196,N_5963,N_5479);
and U6197 (N_6197,N_5180,N_5232);
nand U6198 (N_6198,N_4600,N_4079);
nor U6199 (N_6199,N_4107,N_5793);
or U6200 (N_6200,N_5951,N_4327);
xnor U6201 (N_6201,N_4133,N_5757);
and U6202 (N_6202,N_4635,N_5383);
and U6203 (N_6203,N_5982,N_4777);
nand U6204 (N_6204,N_5961,N_4953);
nand U6205 (N_6205,N_5051,N_5374);
or U6206 (N_6206,N_4176,N_5841);
and U6207 (N_6207,N_4280,N_4463);
or U6208 (N_6208,N_5764,N_5924);
or U6209 (N_6209,N_4477,N_5192);
xor U6210 (N_6210,N_4517,N_4942);
or U6211 (N_6211,N_4097,N_5730);
nand U6212 (N_6212,N_5069,N_5739);
nor U6213 (N_6213,N_4701,N_5801);
and U6214 (N_6214,N_5429,N_5098);
xor U6215 (N_6215,N_4529,N_4561);
nand U6216 (N_6216,N_5005,N_4848);
xnor U6217 (N_6217,N_5704,N_4800);
nor U6218 (N_6218,N_4902,N_5667);
nand U6219 (N_6219,N_5992,N_4451);
nor U6220 (N_6220,N_5168,N_5446);
or U6221 (N_6221,N_5641,N_4479);
or U6222 (N_6222,N_4081,N_4652);
or U6223 (N_6223,N_5990,N_5322);
and U6224 (N_6224,N_5818,N_5457);
nor U6225 (N_6225,N_5782,N_5349);
and U6226 (N_6226,N_5975,N_5418);
and U6227 (N_6227,N_4418,N_5552);
or U6228 (N_6228,N_5871,N_4835);
and U6229 (N_6229,N_4559,N_5242);
xnor U6230 (N_6230,N_5236,N_5362);
xnor U6231 (N_6231,N_5490,N_4875);
nor U6232 (N_6232,N_5905,N_4061);
or U6233 (N_6233,N_5970,N_5597);
and U6234 (N_6234,N_5283,N_5159);
and U6235 (N_6235,N_4576,N_4037);
nand U6236 (N_6236,N_4618,N_4504);
or U6237 (N_6237,N_5397,N_5078);
and U6238 (N_6238,N_4141,N_5957);
nor U6239 (N_6239,N_4880,N_5976);
xnor U6240 (N_6240,N_5154,N_5030);
and U6241 (N_6241,N_5199,N_5938);
nor U6242 (N_6242,N_5411,N_4240);
nand U6243 (N_6243,N_5915,N_5885);
and U6244 (N_6244,N_4434,N_5266);
nand U6245 (N_6245,N_4990,N_4579);
and U6246 (N_6246,N_4492,N_4702);
and U6247 (N_6247,N_5213,N_5364);
nor U6248 (N_6248,N_5074,N_5393);
nor U6249 (N_6249,N_5557,N_4369);
nand U6250 (N_6250,N_5605,N_4042);
nand U6251 (N_6251,N_4657,N_4613);
nand U6252 (N_6252,N_5453,N_4308);
nor U6253 (N_6253,N_4026,N_4588);
nor U6254 (N_6254,N_4833,N_5169);
or U6255 (N_6255,N_5291,N_5972);
and U6256 (N_6256,N_5150,N_5366);
nand U6257 (N_6257,N_5138,N_4629);
nand U6258 (N_6258,N_4715,N_4028);
or U6259 (N_6259,N_5151,N_4532);
nor U6260 (N_6260,N_4646,N_5046);
or U6261 (N_6261,N_5577,N_5348);
nand U6262 (N_6262,N_5271,N_5282);
nor U6263 (N_6263,N_5088,N_4789);
nor U6264 (N_6264,N_4215,N_5816);
xor U6265 (N_6265,N_4617,N_4250);
or U6266 (N_6266,N_5533,N_5837);
and U6267 (N_6267,N_5220,N_5137);
and U6268 (N_6268,N_5690,N_4979);
or U6269 (N_6269,N_4162,N_5080);
or U6270 (N_6270,N_5723,N_4689);
nor U6271 (N_6271,N_4491,N_5092);
nor U6272 (N_6272,N_4699,N_5761);
or U6273 (N_6273,N_5657,N_5303);
nor U6274 (N_6274,N_4620,N_4666);
and U6275 (N_6275,N_5601,N_5882);
and U6276 (N_6276,N_5848,N_4116);
and U6277 (N_6277,N_5301,N_4260);
nor U6278 (N_6278,N_4086,N_5216);
or U6279 (N_6279,N_4938,N_4148);
or U6280 (N_6280,N_4911,N_5261);
or U6281 (N_6281,N_4978,N_5486);
xor U6282 (N_6282,N_4973,N_4267);
nand U6283 (N_6283,N_4787,N_5440);
xnor U6284 (N_6284,N_5607,N_4895);
and U6285 (N_6285,N_4006,N_4640);
xor U6286 (N_6286,N_4029,N_5464);
nor U6287 (N_6287,N_4688,N_5623);
or U6288 (N_6288,N_5011,N_4548);
and U6289 (N_6289,N_5728,N_5091);
nor U6290 (N_6290,N_4645,N_5373);
nand U6291 (N_6291,N_5611,N_4401);
and U6292 (N_6292,N_4972,N_5305);
nand U6293 (N_6293,N_5113,N_4189);
or U6294 (N_6294,N_4461,N_4452);
xor U6295 (N_6295,N_5960,N_5452);
or U6296 (N_6296,N_5378,N_5953);
and U6297 (N_6297,N_5043,N_5855);
and U6298 (N_6298,N_4306,N_4344);
and U6299 (N_6299,N_5901,N_4812);
and U6300 (N_6300,N_4592,N_4122);
nor U6301 (N_6301,N_4410,N_4541);
nor U6302 (N_6302,N_4912,N_4105);
xnor U6303 (N_6303,N_4553,N_4188);
or U6304 (N_6304,N_4788,N_4970);
and U6305 (N_6305,N_4609,N_5618);
nand U6306 (N_6306,N_4732,N_5094);
or U6307 (N_6307,N_5712,N_5564);
or U6308 (N_6308,N_4021,N_5344);
nor U6309 (N_6309,N_4533,N_4497);
nand U6310 (N_6310,N_4080,N_5028);
nand U6311 (N_6311,N_5031,N_4347);
xor U6312 (N_6312,N_5934,N_5459);
nand U6313 (N_6313,N_5888,N_4236);
or U6314 (N_6314,N_4551,N_5454);
nand U6315 (N_6315,N_5517,N_4882);
nor U6316 (N_6316,N_4323,N_4868);
or U6317 (N_6317,N_5570,N_4485);
xnor U6318 (N_6318,N_5206,N_5695);
xor U6319 (N_6319,N_4432,N_5731);
and U6320 (N_6320,N_4897,N_4887);
or U6321 (N_6321,N_5650,N_5346);
nand U6322 (N_6322,N_5360,N_4415);
nor U6323 (N_6323,N_4174,N_4510);
or U6324 (N_6324,N_5336,N_5502);
or U6325 (N_6325,N_5654,N_5802);
or U6326 (N_6326,N_5164,N_4033);
nor U6327 (N_6327,N_5447,N_4390);
or U6328 (N_6328,N_4676,N_5000);
or U6329 (N_6329,N_5115,N_5408);
nor U6330 (N_6330,N_4179,N_5489);
nor U6331 (N_6331,N_5958,N_5073);
or U6332 (N_6332,N_5504,N_4679);
or U6333 (N_6333,N_4717,N_4693);
nor U6334 (N_6334,N_4445,N_5573);
or U6335 (N_6335,N_5535,N_5689);
or U6336 (N_6336,N_4224,N_5735);
nor U6337 (N_6337,N_5404,N_4376);
xor U6338 (N_6338,N_5425,N_5740);
nor U6339 (N_6339,N_4669,N_5785);
nor U6340 (N_6340,N_4568,N_5345);
nor U6341 (N_6341,N_4755,N_5854);
or U6342 (N_6342,N_4927,N_5002);
and U6343 (N_6343,N_5696,N_4462);
and U6344 (N_6344,N_4460,N_4349);
and U6345 (N_6345,N_5684,N_4339);
nor U6346 (N_6346,N_5257,N_5477);
nor U6347 (N_6347,N_4575,N_5868);
nor U6348 (N_6348,N_5296,N_5514);
nand U6349 (N_6349,N_4486,N_4771);
and U6350 (N_6350,N_5369,N_5285);
or U6351 (N_6351,N_5510,N_5104);
and U6352 (N_6352,N_5077,N_4871);
and U6353 (N_6353,N_4616,N_4831);
nand U6354 (N_6354,N_4483,N_4293);
nand U6355 (N_6355,N_4473,N_4299);
and U6356 (N_6356,N_4470,N_5920);
and U6357 (N_6357,N_4951,N_4190);
nor U6358 (N_6358,N_4749,N_4986);
nand U6359 (N_6359,N_4324,N_5664);
nor U6360 (N_6360,N_5907,N_4537);
or U6361 (N_6361,N_4971,N_4678);
nand U6362 (N_6362,N_4405,N_4667);
and U6363 (N_6363,N_5281,N_5658);
xnor U6364 (N_6364,N_4608,N_4301);
xnor U6365 (N_6365,N_4220,N_5526);
nor U6366 (N_6366,N_5053,N_4849);
or U6367 (N_6367,N_5226,N_4222);
nand U6368 (N_6368,N_4276,N_4332);
nand U6369 (N_6369,N_4720,N_5341);
nor U6370 (N_6370,N_4158,N_4412);
nand U6371 (N_6371,N_4244,N_4254);
nor U6372 (N_6372,N_4498,N_4527);
and U6373 (N_6373,N_4984,N_5507);
and U6374 (N_6374,N_4433,N_4719);
nor U6375 (N_6375,N_5027,N_5989);
nor U6376 (N_6376,N_5280,N_5763);
and U6377 (N_6377,N_4231,N_5127);
or U6378 (N_6378,N_5671,N_5978);
or U6379 (N_6379,N_5461,N_4832);
or U6380 (N_6380,N_5288,N_4059);
nor U6381 (N_6381,N_4772,N_4992);
nand U6382 (N_6382,N_4488,N_5324);
nor U6383 (N_6383,N_4858,N_5518);
nand U6384 (N_6384,N_5386,N_4449);
and U6385 (N_6385,N_5316,N_4905);
or U6386 (N_6386,N_4980,N_4329);
and U6387 (N_6387,N_4536,N_4458);
nor U6388 (N_6388,N_5578,N_4241);
or U6389 (N_6389,N_4214,N_5773);
and U6390 (N_6390,N_5846,N_5456);
and U6391 (N_6391,N_4554,N_4310);
nand U6392 (N_6392,N_5683,N_5279);
xor U6393 (N_6393,N_4103,N_4099);
nor U6394 (N_6394,N_5445,N_5265);
nor U6395 (N_6395,N_5198,N_5914);
or U6396 (N_6396,N_5415,N_5356);
and U6397 (N_6397,N_5553,N_5037);
and U6398 (N_6398,N_4440,N_5505);
xnor U6399 (N_6399,N_4077,N_5851);
nor U6400 (N_6400,N_4457,N_5222);
nand U6401 (N_6401,N_5352,N_4847);
and U6402 (N_6402,N_4325,N_5273);
xor U6403 (N_6403,N_5219,N_5546);
nand U6404 (N_6404,N_5939,N_5317);
or U6405 (N_6405,N_4145,N_4539);
nand U6406 (N_6406,N_5659,N_4844);
nor U6407 (N_6407,N_5861,N_4196);
nor U6408 (N_6408,N_4705,N_4184);
nand U6409 (N_6409,N_5760,N_5024);
and U6410 (N_6410,N_5519,N_5530);
and U6411 (N_6411,N_5034,N_5622);
nand U6412 (N_6412,N_4857,N_5863);
nand U6413 (N_6413,N_4091,N_4137);
xnor U6414 (N_6414,N_5320,N_4836);
or U6415 (N_6415,N_4672,N_4223);
and U6416 (N_6416,N_4869,N_4371);
nor U6417 (N_6417,N_4109,N_4048);
nand U6418 (N_6418,N_5850,N_5534);
or U6419 (N_6419,N_5538,N_4919);
nand U6420 (N_6420,N_5828,N_4270);
and U6421 (N_6421,N_5059,N_5835);
or U6422 (N_6422,N_4114,N_5734);
nor U6423 (N_6423,N_5493,N_4071);
nor U6424 (N_6424,N_4258,N_4167);
or U6425 (N_6425,N_5902,N_4387);
nand U6426 (N_6426,N_5047,N_4353);
and U6427 (N_6427,N_5465,N_4273);
xnor U6428 (N_6428,N_4860,N_5506);
or U6429 (N_6429,N_4159,N_5595);
or U6430 (N_6430,N_4030,N_5379);
and U6431 (N_6431,N_4027,N_4493);
or U6432 (N_6432,N_4139,N_5867);
and U6433 (N_6433,N_4044,N_5665);
xor U6434 (N_6434,N_5776,N_4453);
and U6435 (N_6435,N_5121,N_4377);
and U6436 (N_6436,N_5302,N_4750);
or U6437 (N_6437,N_4818,N_4695);
and U6438 (N_6438,N_4845,N_4601);
nand U6439 (N_6439,N_4480,N_4637);
and U6440 (N_6440,N_5375,N_4842);
and U6441 (N_6441,N_4639,N_5596);
nand U6442 (N_6442,N_5496,N_4078);
nor U6443 (N_6443,N_5779,N_5935);
nand U6444 (N_6444,N_4589,N_4906);
nor U6445 (N_6445,N_5093,N_5149);
nor U6446 (N_6446,N_5883,N_5869);
or U6447 (N_6447,N_4878,N_4274);
or U6448 (N_6448,N_4102,N_5847);
nor U6449 (N_6449,N_5574,N_4092);
and U6450 (N_6450,N_4981,N_5598);
nor U6451 (N_6451,N_4475,N_4368);
nor U6452 (N_6452,N_4051,N_5434);
and U6453 (N_6453,N_5608,N_5815);
xor U6454 (N_6454,N_5720,N_5380);
nor U6455 (N_6455,N_4700,N_4976);
nor U6456 (N_6456,N_5361,N_4118);
nor U6457 (N_6457,N_5402,N_4500);
nand U6458 (N_6458,N_4685,N_4411);
and U6459 (N_6459,N_4560,N_5191);
xnor U6460 (N_6460,N_4681,N_5381);
nor U6461 (N_6461,N_4530,N_4481);
or U6462 (N_6462,N_5893,N_5692);
nor U6463 (N_6463,N_5229,N_4995);
or U6464 (N_6464,N_4271,N_5060);
and U6465 (N_6465,N_5756,N_4745);
or U6466 (N_6466,N_4773,N_4759);
nand U6467 (N_6467,N_4988,N_4762);
nand U6468 (N_6468,N_5177,N_4361);
nor U6469 (N_6469,N_5466,N_5777);
and U6470 (N_6470,N_4177,N_4586);
nor U6471 (N_6471,N_5772,N_4286);
nand U6472 (N_6472,N_4181,N_4697);
nand U6473 (N_6473,N_5637,N_5955);
and U6474 (N_6474,N_4744,N_4945);
xnor U6475 (N_6475,N_5997,N_5697);
and U6476 (N_6476,N_5586,N_5956);
nand U6477 (N_6477,N_5922,N_4596);
or U6478 (N_6478,N_5260,N_5148);
nand U6479 (N_6479,N_4644,N_4738);
and U6480 (N_6480,N_5107,N_4735);
nand U6481 (N_6481,N_4183,N_5925);
and U6482 (N_6482,N_4038,N_4658);
or U6483 (N_6483,N_5309,N_5082);
nand U6484 (N_6484,N_4201,N_4113);
nand U6485 (N_6485,N_5700,N_4023);
nand U6486 (N_6486,N_4337,N_4202);
and U6487 (N_6487,N_4820,N_5335);
or U6488 (N_6488,N_4436,N_4928);
nor U6489 (N_6489,N_4378,N_5579);
xor U6490 (N_6490,N_5768,N_4740);
or U6491 (N_6491,N_5543,N_5455);
nand U6492 (N_6492,N_4512,N_4151);
xor U6493 (N_6493,N_5014,N_4358);
nor U6494 (N_6494,N_5252,N_4946);
nor U6495 (N_6495,N_4631,N_4009);
and U6496 (N_6496,N_5221,N_5588);
and U6497 (N_6497,N_4318,N_4019);
and U6498 (N_6498,N_4002,N_5246);
and U6499 (N_6499,N_5931,N_5726);
nand U6500 (N_6500,N_5103,N_4394);
nor U6501 (N_6501,N_4798,N_4232);
and U6502 (N_6502,N_4756,N_5710);
xor U6503 (N_6503,N_4545,N_5559);
nand U6504 (N_6504,N_4816,N_4966);
nor U6505 (N_6505,N_5162,N_4175);
nor U6506 (N_6506,N_5267,N_5172);
xor U6507 (N_6507,N_4359,N_4853);
nand U6508 (N_6508,N_5227,N_5576);
and U6509 (N_6509,N_5766,N_4138);
nor U6510 (N_6510,N_4997,N_5722);
nand U6511 (N_6511,N_4960,N_4623);
nand U6512 (N_6512,N_4521,N_5311);
and U6513 (N_6513,N_4065,N_5532);
nand U6514 (N_6514,N_4581,N_4540);
or U6515 (N_6515,N_5437,N_5062);
and U6516 (N_6516,N_5200,N_5008);
or U6517 (N_6517,N_5536,N_5117);
and U6518 (N_6518,N_4170,N_5342);
and U6519 (N_6519,N_5746,N_4437);
nand U6520 (N_6520,N_5156,N_4785);
and U6521 (N_6521,N_4721,N_5811);
xor U6522 (N_6522,N_4283,N_5544);
or U6523 (N_6523,N_4111,N_4153);
or U6524 (N_6524,N_4302,N_4572);
xor U6525 (N_6525,N_5865,N_4164);
nor U6526 (N_6526,N_5903,N_4944);
xor U6527 (N_6527,N_4888,N_5625);
and U6528 (N_6528,N_4335,N_5253);
nand U6529 (N_6529,N_4351,N_4642);
and U6530 (N_6530,N_4468,N_4040);
nor U6531 (N_6531,N_5711,N_4661);
and U6532 (N_6532,N_4977,N_5128);
nor U6533 (N_6533,N_4193,N_5463);
and U6534 (N_6534,N_4603,N_5645);
and U6535 (N_6535,N_4256,N_5843);
and U6536 (N_6536,N_5314,N_5838);
nand U6537 (N_6537,N_4088,N_4627);
xor U6538 (N_6538,N_4577,N_5895);
nor U6539 (N_6539,N_5340,N_4522);
and U6540 (N_6540,N_5421,N_5438);
and U6541 (N_6541,N_4913,N_4422);
or U6542 (N_6542,N_5387,N_4748);
and U6543 (N_6543,N_5941,N_4294);
or U6544 (N_6544,N_5909,N_5844);
and U6545 (N_6545,N_5478,N_5142);
xnor U6546 (N_6546,N_4684,N_4959);
or U6547 (N_6547,N_5555,N_5359);
or U6548 (N_6548,N_4169,N_5713);
nand U6549 (N_6549,N_5394,N_4594);
and U6550 (N_6550,N_4769,N_4659);
nand U6551 (N_6551,N_5315,N_5243);
or U6552 (N_6552,N_5558,N_4707);
nor U6553 (N_6553,N_5054,N_4694);
or U6554 (N_6554,N_5520,N_5482);
or U6555 (N_6555,N_4999,N_4754);
nand U6556 (N_6556,N_5744,N_4443);
xor U6557 (N_6557,N_5593,N_4482);
nor U6558 (N_6558,N_4210,N_4253);
and U6559 (N_6559,N_4610,N_4355);
xnor U6560 (N_6560,N_5977,N_4766);
or U6561 (N_6561,N_5714,N_4125);
nor U6562 (N_6562,N_5560,N_5274);
or U6563 (N_6563,N_5350,N_5208);
nand U6564 (N_6564,N_4723,N_5259);
or U6565 (N_6565,N_4962,N_5286);
nor U6566 (N_6566,N_5524,N_4896);
or U6567 (N_6567,N_5767,N_5602);
nor U6568 (N_6568,N_4626,N_4200);
nor U6569 (N_6569,N_5247,N_4806);
and U6570 (N_6570,N_4673,N_5691);
nand U6571 (N_6571,N_4487,N_4501);
or U6572 (N_6572,N_5368,N_5006);
nor U6573 (N_6573,N_4025,N_5049);
nor U6574 (N_6574,N_5334,N_4993);
or U6575 (N_6575,N_5891,N_5114);
nand U6576 (N_6576,N_5343,N_4916);
and U6577 (N_6577,N_4047,N_5084);
and U6578 (N_6578,N_4414,N_5540);
nor U6579 (N_6579,N_4441,N_4949);
and U6580 (N_6580,N_4003,N_4380);
and U6581 (N_6581,N_4146,N_5609);
nor U6582 (N_6582,N_4954,N_4649);
nor U6583 (N_6583,N_4259,N_5666);
or U6584 (N_6584,N_4225,N_5655);
and U6585 (N_6585,N_4614,N_4124);
nand U6586 (N_6586,N_5663,N_4211);
nor U6587 (N_6587,N_4063,N_4641);
or U6588 (N_6588,N_5102,N_5188);
or U6589 (N_6589,N_5653,N_5745);
nand U6590 (N_6590,N_4663,N_5621);
xor U6591 (N_6591,N_5210,N_5825);
or U6592 (N_6592,N_5707,N_4898);
xor U6593 (N_6593,N_5231,N_5525);
nand U6594 (N_6594,N_5980,N_5567);
and U6595 (N_6595,N_5996,N_5313);
nor U6596 (N_6596,N_4534,N_5571);
and U6597 (N_6597,N_4711,N_5398);
nor U6598 (N_6598,N_4288,N_4187);
nand U6599 (N_6599,N_5646,N_4367);
nand U6600 (N_6600,N_4045,N_5983);
and U6601 (N_6601,N_4760,N_5900);
and U6602 (N_6602,N_4108,N_4309);
nor U6603 (N_6603,N_4062,N_4587);
and U6604 (N_6604,N_5284,N_5705);
nor U6605 (N_6605,N_5827,N_5268);
nor U6606 (N_6606,N_5632,N_5224);
or U6607 (N_6607,N_5879,N_4290);
nand U6608 (N_6608,N_5312,N_5881);
or U6609 (N_6609,N_4034,N_4014);
nor U6610 (N_6610,N_5715,N_4243);
or U6611 (N_6611,N_4024,N_4780);
or U6612 (N_6612,N_4852,N_4628);
or U6613 (N_6613,N_5775,N_4373);
or U6614 (N_6614,N_4682,N_4383);
or U6615 (N_6615,N_4300,N_4316);
nand U6616 (N_6616,N_4269,N_5233);
or U6617 (N_6617,N_4651,N_4567);
nand U6618 (N_6618,N_5498,N_5672);
and U6619 (N_6619,N_4523,N_4922);
nor U6620 (N_6620,N_5857,N_5449);
nor U6621 (N_6621,N_4925,N_5950);
nor U6622 (N_6622,N_5009,N_4991);
nand U6623 (N_6623,N_5333,N_5561);
and U6624 (N_6624,N_4313,N_5933);
or U6625 (N_6625,N_4221,N_4933);
or U6626 (N_6626,N_4010,N_4467);
or U6627 (N_6627,N_4036,N_4073);
and U6628 (N_6628,N_4213,N_4538);
or U6629 (N_6629,N_5787,N_5919);
xor U6630 (N_6630,N_4049,N_5419);
nand U6631 (N_6631,N_5652,N_4282);
nand U6632 (N_6632,N_4403,N_5681);
or U6633 (N_6633,N_4696,N_5277);
nor U6634 (N_6634,N_5969,N_5214);
xnor U6635 (N_6635,N_4515,N_4476);
or U6636 (N_6636,N_4604,N_4076);
or U6637 (N_6637,N_5173,N_5012);
or U6638 (N_6638,N_5842,N_4957);
and U6639 (N_6639,N_5035,N_4727);
or U6640 (N_6640,N_5718,N_4011);
or U6641 (N_6641,N_4619,N_4931);
nand U6642 (N_6642,N_5111,N_4743);
nor U6643 (N_6643,N_5991,N_4856);
xor U6644 (N_6644,N_4710,N_4615);
nand U6645 (N_6645,N_4284,N_5458);
and U6646 (N_6646,N_5729,N_5332);
nor U6647 (N_6647,N_5161,N_5420);
or U6648 (N_6648,N_4864,N_4165);
nand U6649 (N_6649,N_4570,N_5004);
and U6650 (N_6650,N_4295,N_4778);
and U6651 (N_6651,N_5946,N_5822);
nand U6652 (N_6652,N_5019,N_5644);
xor U6653 (N_6653,N_5660,N_4814);
nand U6654 (N_6654,N_4506,N_5503);
nor U6655 (N_6655,N_4104,N_5531);
nand U6656 (N_6656,N_5765,N_4822);
and U6657 (N_6657,N_5239,N_4012);
nor U6658 (N_6658,N_5254,N_4499);
nand U6659 (N_6659,N_4322,N_4375);
nand U6660 (N_6660,N_4431,N_4872);
nand U6661 (N_6661,N_5377,N_5784);
xnor U6662 (N_6662,N_5160,N_5703);
nand U6663 (N_6663,N_5515,N_5747);
nand U6664 (N_6664,N_5849,N_4574);
and U6665 (N_6665,N_4825,N_5426);
and U6666 (N_6666,N_5936,N_5649);
nor U6667 (N_6667,N_5856,N_4131);
or U6668 (N_6668,N_4648,N_5679);
and U6669 (N_6669,N_5541,N_4914);
nor U6670 (N_6670,N_4675,N_4364);
nor U6671 (N_6671,N_5351,N_4208);
xnor U6672 (N_6672,N_5912,N_5399);
nand U6673 (N_6673,N_4069,N_5179);
nor U6674 (N_6674,N_4056,N_4416);
or U6675 (N_6675,N_5197,N_5619);
nand U6676 (N_6676,N_5372,N_5613);
or U6677 (N_6677,N_4725,N_4289);
or U6678 (N_6678,N_5300,N_4765);
or U6679 (N_6679,N_5292,N_5783);
or U6680 (N_6680,N_4001,N_5509);
or U6681 (N_6681,N_4296,N_4417);
or U6682 (N_6682,N_5409,N_4197);
nor U6683 (N_6683,N_5870,N_5003);
or U6684 (N_6684,N_5737,N_5769);
nor U6685 (N_6685,N_5890,N_4095);
nand U6686 (N_6686,N_5986,N_4582);
nor U6687 (N_6687,N_5833,N_5116);
and U6688 (N_6688,N_5821,N_4809);
nor U6689 (N_6689,N_4861,N_5643);
or U6690 (N_6690,N_5708,N_5278);
nor U6691 (N_6691,N_4963,N_4961);
and U6692 (N_6692,N_4039,N_5495);
and U6693 (N_6693,N_4839,N_4528);
or U6694 (N_6694,N_5163,N_4312);
nor U6695 (N_6695,N_4543,N_5968);
xnor U6696 (N_6696,N_5831,N_5648);
nand U6697 (N_6697,N_4348,N_5147);
nand U6698 (N_6698,N_4607,N_4654);
nor U6699 (N_6699,N_5556,N_4421);
and U6700 (N_6700,N_5887,N_5428);
or U6701 (N_6701,N_5190,N_5338);
nor U6702 (N_6702,N_5189,N_4591);
and U6703 (N_6703,N_4894,N_5450);
nand U6704 (N_6704,N_4217,N_5944);
or U6705 (N_6705,N_5508,N_5123);
and U6706 (N_6706,N_4932,N_5910);
nor U6707 (N_6707,N_4389,N_5642);
nor U6708 (N_6708,N_5752,N_5144);
and U6709 (N_6709,N_4660,N_4249);
and U6710 (N_6710,N_4903,N_4228);
and U6711 (N_6711,N_4775,N_4790);
or U6712 (N_6712,N_4072,N_4142);
xnor U6713 (N_6713,N_4219,N_5721);
and U6714 (N_6714,N_5451,N_4192);
and U6715 (N_6715,N_5799,N_5947);
or U6716 (N_6716,N_5706,N_5949);
or U6717 (N_6717,N_5065,N_4671);
xor U6718 (N_6718,N_4186,N_4683);
and U6719 (N_6719,N_5545,N_4251);
nand U6720 (N_6720,N_5636,N_4182);
or U6721 (N_6721,N_4396,N_5329);
nor U6722 (N_6722,N_5751,N_5085);
or U6723 (N_6723,N_4824,N_5750);
xor U6724 (N_6724,N_4808,N_4712);
nand U6725 (N_6725,N_4008,N_4730);
nand U6726 (N_6726,N_5045,N_4366);
nand U6727 (N_6727,N_4889,N_5677);
and U6728 (N_6728,N_4100,N_5537);
nand U6729 (N_6729,N_4815,N_4741);
and U6730 (N_6730,N_5845,N_4514);
nor U6731 (N_6731,N_4321,N_4909);
nor U6732 (N_6732,N_4068,N_4837);
nand U6733 (N_6733,N_5042,N_4593);
xor U6734 (N_6734,N_4634,N_5572);
or U6735 (N_6735,N_5539,N_4602);
xor U6736 (N_6736,N_4031,N_5804);
nor U6737 (N_6737,N_5435,N_4625);
and U6738 (N_6738,N_5973,N_4915);
nand U6739 (N_6739,N_5962,N_5319);
or U6740 (N_6740,N_5874,N_4005);
or U6741 (N_6741,N_4067,N_5583);
and U6742 (N_6742,N_5554,N_5238);
nand U6743 (N_6743,N_5215,N_4855);
nand U6744 (N_6744,N_5674,N_4154);
and U6745 (N_6745,N_4714,N_4469);
and U6746 (N_6746,N_4890,N_4768);
xor U6747 (N_6747,N_4305,N_5670);
nor U6748 (N_6748,N_5410,N_4943);
or U6749 (N_6749,N_5719,N_4395);
nand U6750 (N_6750,N_5308,N_4662);
nand U6751 (N_6751,N_4303,N_4066);
and U6752 (N_6752,N_4585,N_5020);
xor U6753 (N_6753,N_4901,N_5158);
nor U6754 (N_6754,N_4004,N_4398);
xor U6755 (N_6755,N_5422,N_5071);
nor U6756 (N_6756,N_4886,N_4605);
xor U6757 (N_6757,N_4866,N_5070);
nor U6758 (N_6758,N_5339,N_5202);
or U6759 (N_6759,N_5615,N_4018);
or U6760 (N_6760,N_4792,N_4680);
or U6761 (N_6761,N_4317,N_4865);
and U6762 (N_6762,N_4185,N_4811);
nor U6763 (N_6763,N_4921,N_4017);
nor U6764 (N_6764,N_4140,N_4266);
xor U6765 (N_6765,N_5631,N_5987);
nor U6766 (N_6766,N_4677,N_4899);
nor U6767 (N_6767,N_5575,N_5927);
nor U6768 (N_6768,N_4247,N_5439);
and U6769 (N_6769,N_4690,N_4737);
or U6770 (N_6770,N_5196,N_5662);
xnor U6771 (N_6771,N_5600,N_4281);
or U6772 (N_6772,N_5264,N_4950);
and U6773 (N_6773,N_4448,N_5832);
or U6774 (N_6774,N_4370,N_5433);
nand U6775 (N_6775,N_4797,N_5594);
or U6776 (N_6776,N_5732,N_5717);
or U6777 (N_6777,N_4505,N_5444);
or U6778 (N_6778,N_5786,N_4948);
and U6779 (N_6779,N_4873,N_4198);
xor U6780 (N_6780,N_5693,N_4408);
nor U6781 (N_6781,N_5321,N_4770);
nand U6782 (N_6782,N_5101,N_5651);
or U6783 (N_6783,N_5954,N_5948);
and U6784 (N_6784,N_5391,N_4331);
xor U6785 (N_6785,N_5187,N_4206);
nand U6786 (N_6786,N_5647,N_5630);
xor U6787 (N_6787,N_4547,N_5823);
nor U6788 (N_6788,N_4257,N_4490);
nand U6789 (N_6789,N_4934,N_5388);
nand U6790 (N_6790,N_4209,N_4940);
or U6791 (N_6791,N_4235,N_4885);
nor U6792 (N_6792,N_4583,N_5635);
nor U6793 (N_6793,N_5323,N_4239);
and U6794 (N_6794,N_5079,N_4746);
nand U6795 (N_6795,N_4397,N_4195);
xnor U6796 (N_6796,N_4653,N_4508);
nand U6797 (N_6797,N_4098,N_5480);
nand U6798 (N_6798,N_5817,N_5738);
xor U6799 (N_6799,N_5396,N_4127);
and U6800 (N_6800,N_5736,N_4233);
and U6801 (N_6801,N_4084,N_5886);
and U6802 (N_6802,N_4074,N_5795);
or U6803 (N_6803,N_4126,N_5068);
xor U6804 (N_6804,N_4474,N_5789);
or U6805 (N_6805,N_4043,N_5603);
or U6806 (N_6806,N_4466,N_5853);
and U6807 (N_6807,N_4178,N_4708);
nor U6808 (N_6808,N_4342,N_4287);
nor U6809 (N_6809,N_5694,N_4120);
nor U6810 (N_6810,N_5328,N_4428);
or U6811 (N_6811,N_5500,N_5367);
xor U6812 (N_6812,N_4726,N_5604);
nor U6813 (N_6813,N_5809,N_5995);
xor U6814 (N_6814,N_4484,N_4085);
and U6815 (N_6815,N_5155,N_5357);
and U6816 (N_6816,N_5263,N_5528);
or U6817 (N_6817,N_5064,N_5165);
nor U6818 (N_6818,N_4918,N_5896);
nand U6819 (N_6819,N_5347,N_5460);
nor U6820 (N_6820,N_4399,N_5952);
nand U6821 (N_6821,N_4409,N_5904);
nand U6822 (N_6822,N_5494,N_4255);
nand U6823 (N_6823,N_4563,N_5018);
nor U6824 (N_6824,N_5417,N_5589);
nand U6825 (N_6825,N_5669,N_5167);
nand U6826 (N_6826,N_4704,N_5403);
nor U6827 (N_6827,N_4687,N_5427);
nor U6828 (N_6828,N_5688,N_4372);
or U6829 (N_6829,N_4843,N_4338);
and U6830 (N_6830,N_5297,N_5081);
xor U6831 (N_6831,N_5066,N_5223);
xnor U6832 (N_6832,N_4562,N_5599);
or U6833 (N_6833,N_4388,N_4791);
and U6834 (N_6834,N_4670,N_4227);
and U6835 (N_6835,N_4464,N_5511);
and U6836 (N_6836,N_4279,N_5864);
xor U6837 (N_6837,N_5894,N_4050);
nand U6838 (N_6838,N_5076,N_5862);
nor U6839 (N_6839,N_4975,N_5108);
and U6840 (N_6840,N_4763,N_4203);
and U6841 (N_6841,N_5290,N_5778);
nand U6842 (N_6842,N_5044,N_4716);
and U6843 (N_6843,N_5306,N_4496);
nand U6844 (N_6844,N_4041,N_5940);
and U6845 (N_6845,N_5497,N_5686);
and U6846 (N_6846,N_5866,N_4032);
nand U6847 (N_6847,N_4996,N_4656);
nor U6848 (N_6848,N_4334,N_4307);
or U6849 (N_6849,N_4724,N_5725);
or U6850 (N_6850,N_4263,N_5325);
nor U6851 (N_6851,N_4191,N_5701);
nor U6852 (N_6852,N_4503,N_4786);
and U6853 (N_6853,N_5384,N_4346);
or U6854 (N_6854,N_4664,N_4319);
xor U6855 (N_6855,N_4157,N_5742);
or U6856 (N_6856,N_5547,N_5551);
nor U6857 (N_6857,N_5025,N_4877);
and U6858 (N_6858,N_4691,N_4229);
or U6859 (N_6859,N_4345,N_5204);
nor U6860 (N_6860,N_5770,N_5310);
and U6861 (N_6861,N_4879,N_4513);
nor U6862 (N_6862,N_4793,N_4465);
and U6863 (N_6863,N_4509,N_5899);
xor U6864 (N_6864,N_4923,N_5628);
or U6865 (N_6865,N_4171,N_4955);
and U6866 (N_6866,N_5467,N_5716);
nand U6867 (N_6867,N_4821,N_4016);
nor U6868 (N_6868,N_5376,N_4311);
or U6869 (N_6869,N_5754,N_4336);
and U6870 (N_6870,N_4357,N_4494);
or U6871 (N_6871,N_4840,N_4883);
nand U6872 (N_6872,N_4952,N_4237);
and U6873 (N_6873,N_4870,N_4747);
xnor U6874 (N_6874,N_5353,N_5937);
or U6875 (N_6875,N_5917,N_4430);
nand U6876 (N_6876,N_5872,N_4150);
and U6877 (N_6877,N_4647,N_5640);
and U6878 (N_6878,N_5139,N_5337);
or U6879 (N_6879,N_4392,N_5136);
nor U6880 (N_6880,N_4173,N_4796);
nand U6881 (N_6881,N_5134,N_5612);
nand U6882 (N_6882,N_4781,N_4935);
nand U6883 (N_6883,N_4057,N_4758);
nand U6884 (N_6884,N_4830,N_5178);
xor U6885 (N_6885,N_4155,N_5878);
xnor U6886 (N_6886,N_5140,N_4779);
or U6887 (N_6887,N_4374,N_4736);
nand U6888 (N_6888,N_4565,N_5240);
and U6889 (N_6889,N_5807,N_5157);
nand U6890 (N_6890,N_5826,N_4424);
or U6891 (N_6891,N_5814,N_4117);
nor U6892 (N_6892,N_5131,N_5481);
and U6893 (N_6893,N_4132,N_4929);
nand U6894 (N_6894,N_5840,N_5967);
nor U6895 (N_6895,N_4519,N_4218);
nand U6896 (N_6896,N_4884,N_4135);
nor U6897 (N_6897,N_5056,N_5610);
or U6898 (N_6898,N_4089,N_5860);
or U6899 (N_6899,N_4958,N_4234);
or U6900 (N_6900,N_5036,N_4874);
xor U6901 (N_6901,N_5624,N_4386);
nand U6902 (N_6902,N_5407,N_5884);
and U6903 (N_6903,N_4936,N_5513);
nand U6904 (N_6904,N_5307,N_4590);
or U6905 (N_6905,N_5244,N_4163);
and U6906 (N_6906,N_5563,N_4810);
nor U6907 (N_6907,N_5171,N_5055);
nand U6908 (N_6908,N_4638,N_5152);
nor U6909 (N_6909,N_5820,N_5468);
nand U6910 (N_6910,N_4230,N_4015);
and U6911 (N_6911,N_5985,N_4447);
or U6912 (N_6912,N_4110,N_5370);
nand U6913 (N_6913,N_5475,N_5472);
nand U6914 (N_6914,N_4784,N_5755);
and U6915 (N_6915,N_5182,N_4381);
nand U6916 (N_6916,N_5145,N_4926);
nand U6917 (N_6917,N_4264,N_5057);
nand U6918 (N_6918,N_5687,N_4807);
and U6919 (N_6919,N_4794,N_4340);
nand U6920 (N_6920,N_4246,N_4413);
nor U6921 (N_6921,N_5293,N_5270);
and U6922 (N_6922,N_5201,N_5921);
and U6923 (N_6923,N_4052,N_4471);
and U6924 (N_6924,N_4706,N_4686);
nand U6925 (N_6925,N_5175,N_4964);
or U6926 (N_6926,N_5568,N_4382);
nor U6927 (N_6927,N_5048,N_5141);
nand U6928 (N_6928,N_4242,N_4630);
xnor U6929 (N_6929,N_4090,N_5501);
nand U6930 (N_6930,N_5371,N_5521);
or U6931 (N_6931,N_4595,N_5299);
nand U6932 (N_6932,N_4407,N_5808);
or U6933 (N_6933,N_4379,N_5999);
and U6934 (N_6934,N_5499,N_4207);
xor U6935 (N_6935,N_4908,N_5523);
nor U6936 (N_6936,N_4578,N_4060);
nand U6937 (N_6937,N_5916,N_4400);
or U6938 (N_6938,N_5733,N_4046);
or U6939 (N_6939,N_5834,N_4920);
and U6940 (N_6940,N_5829,N_5492);
nor U6941 (N_6941,N_4123,N_4365);
nand U6942 (N_6942,N_4064,N_5406);
nor U6943 (N_6943,N_4350,N_5988);
xor U6944 (N_6944,N_5548,N_4917);
nor U6945 (N_6945,N_5585,N_5118);
nor U6946 (N_6946,N_4782,N_5859);
nand U6947 (N_6947,N_5790,N_5590);
xor U6948 (N_6948,N_5023,N_4093);
xor U6949 (N_6949,N_4606,N_4298);
nand U6950 (N_6950,N_5195,N_5276);
nand U6951 (N_6951,N_5926,N_4261);
or U6952 (N_6952,N_5984,N_5797);
nand U6953 (N_6953,N_4265,N_4799);
nand U6954 (N_6954,N_5580,N_5124);
and U6955 (N_6955,N_5414,N_4082);
or U6956 (N_6956,N_4112,N_5616);
xor U6957 (N_6957,N_4834,N_4507);
nor U6958 (N_6958,N_4974,N_4838);
or U6959 (N_6959,N_5330,N_4764);
nor U6960 (N_6960,N_5634,N_4427);
nor U6961 (N_6961,N_4930,N_4989);
and U6962 (N_6962,N_5326,N_5484);
or U6963 (N_6963,N_4802,N_5566);
and U6964 (N_6964,N_4083,N_5110);
nand U6965 (N_6965,N_4819,N_5592);
nor U6966 (N_6966,N_5183,N_5680);
nor U6967 (N_6967,N_4356,N_5363);
nand U6968 (N_6968,N_5698,N_4444);
or U6969 (N_6969,N_5485,N_4472);
or U6970 (N_6970,N_5405,N_5010);
nand U6971 (N_6971,N_4070,N_5205);
or U6972 (N_6972,N_5412,N_5512);
and U6973 (N_6973,N_4804,N_5087);
and U6974 (N_6974,N_4867,N_4134);
xor U6975 (N_6975,N_5105,N_5753);
and U6976 (N_6976,N_4420,N_4204);
nor U6977 (N_6977,N_5075,N_5469);
or U6978 (N_6978,N_5041,N_4827);
nand U6979 (N_6979,N_5072,N_5400);
or U6980 (N_6980,N_5638,N_5582);
or U6981 (N_6981,N_5748,N_4525);
nor U6982 (N_6982,N_5877,N_4285);
or U6983 (N_6983,N_4854,N_4718);
xor U6984 (N_6984,N_4450,N_5529);
nand U6985 (N_6985,N_5476,N_4622);
xnor U6986 (N_6986,N_5724,N_5015);
and U6987 (N_6987,N_4982,N_5096);
or U6988 (N_6988,N_5942,N_5471);
and U6989 (N_6989,N_4558,N_5052);
nor U6990 (N_6990,N_4115,N_5230);
and U6991 (N_6991,N_5483,N_5258);
and U6992 (N_6992,N_4566,N_4967);
nor U6993 (N_6993,N_4384,N_5203);
or U6994 (N_6994,N_5120,N_5810);
and U6995 (N_6995,N_4904,N_4805);
nand U6996 (N_6996,N_4075,N_4698);
nand U6997 (N_6997,N_4643,N_4633);
and U6998 (N_6998,N_4846,N_4489);
or U6999 (N_6999,N_5966,N_5061);
or U7000 (N_7000,N_5627,N_4577);
or U7001 (N_7001,N_4553,N_4907);
or U7002 (N_7002,N_4791,N_5828);
nand U7003 (N_7003,N_4814,N_5617);
nor U7004 (N_7004,N_4099,N_4683);
nor U7005 (N_7005,N_4769,N_5334);
nor U7006 (N_7006,N_5691,N_5538);
and U7007 (N_7007,N_5834,N_5195);
and U7008 (N_7008,N_4425,N_4569);
nor U7009 (N_7009,N_4682,N_4608);
xnor U7010 (N_7010,N_5472,N_4588);
or U7011 (N_7011,N_4235,N_5100);
and U7012 (N_7012,N_4232,N_5118);
or U7013 (N_7013,N_5376,N_5395);
and U7014 (N_7014,N_5325,N_4534);
nor U7015 (N_7015,N_4623,N_5135);
nor U7016 (N_7016,N_4700,N_5205);
nor U7017 (N_7017,N_4387,N_5655);
nand U7018 (N_7018,N_4213,N_4373);
nor U7019 (N_7019,N_5188,N_5586);
and U7020 (N_7020,N_4195,N_4581);
xnor U7021 (N_7021,N_4727,N_5972);
nand U7022 (N_7022,N_5614,N_5462);
and U7023 (N_7023,N_5311,N_5665);
nor U7024 (N_7024,N_4979,N_5761);
and U7025 (N_7025,N_4812,N_4971);
and U7026 (N_7026,N_5842,N_5397);
or U7027 (N_7027,N_4024,N_5151);
or U7028 (N_7028,N_5067,N_5867);
or U7029 (N_7029,N_5913,N_4947);
and U7030 (N_7030,N_5147,N_5118);
and U7031 (N_7031,N_5460,N_5031);
nand U7032 (N_7032,N_4547,N_4247);
or U7033 (N_7033,N_4015,N_5299);
and U7034 (N_7034,N_5470,N_4909);
xor U7035 (N_7035,N_4744,N_5043);
nor U7036 (N_7036,N_4205,N_4736);
nor U7037 (N_7037,N_4133,N_4582);
nor U7038 (N_7038,N_4596,N_4873);
nand U7039 (N_7039,N_4709,N_4754);
or U7040 (N_7040,N_5709,N_5200);
nand U7041 (N_7041,N_5526,N_5054);
nand U7042 (N_7042,N_5702,N_5438);
nand U7043 (N_7043,N_4438,N_4226);
nor U7044 (N_7044,N_4161,N_4619);
and U7045 (N_7045,N_4385,N_5990);
and U7046 (N_7046,N_5970,N_4750);
and U7047 (N_7047,N_5203,N_5680);
or U7048 (N_7048,N_5455,N_5850);
and U7049 (N_7049,N_5855,N_5963);
nor U7050 (N_7050,N_5366,N_5675);
and U7051 (N_7051,N_5686,N_5366);
nor U7052 (N_7052,N_5901,N_5536);
nand U7053 (N_7053,N_5235,N_4571);
nand U7054 (N_7054,N_4931,N_4570);
or U7055 (N_7055,N_5077,N_5310);
nand U7056 (N_7056,N_4587,N_5170);
and U7057 (N_7057,N_5184,N_4044);
nor U7058 (N_7058,N_5846,N_5390);
nand U7059 (N_7059,N_4187,N_4499);
nor U7060 (N_7060,N_5910,N_4643);
nand U7061 (N_7061,N_5240,N_4871);
and U7062 (N_7062,N_4843,N_4570);
or U7063 (N_7063,N_4259,N_5513);
and U7064 (N_7064,N_5183,N_5461);
and U7065 (N_7065,N_4425,N_4455);
nor U7066 (N_7066,N_4015,N_4714);
or U7067 (N_7067,N_4436,N_5412);
or U7068 (N_7068,N_4309,N_4426);
and U7069 (N_7069,N_4772,N_4425);
and U7070 (N_7070,N_4642,N_5573);
and U7071 (N_7071,N_5103,N_5172);
nor U7072 (N_7072,N_4583,N_5707);
nor U7073 (N_7073,N_4029,N_4762);
nor U7074 (N_7074,N_5650,N_4705);
nor U7075 (N_7075,N_4150,N_5958);
nor U7076 (N_7076,N_4297,N_5580);
nor U7077 (N_7077,N_4808,N_5380);
nor U7078 (N_7078,N_4772,N_5610);
or U7079 (N_7079,N_4153,N_5874);
and U7080 (N_7080,N_5684,N_4302);
or U7081 (N_7081,N_4730,N_5694);
xnor U7082 (N_7082,N_5571,N_4667);
nand U7083 (N_7083,N_4870,N_5944);
or U7084 (N_7084,N_5268,N_5033);
nor U7085 (N_7085,N_4198,N_5933);
nor U7086 (N_7086,N_5068,N_5859);
nand U7087 (N_7087,N_4190,N_4678);
nand U7088 (N_7088,N_5235,N_4142);
and U7089 (N_7089,N_4881,N_5232);
or U7090 (N_7090,N_5852,N_5092);
nor U7091 (N_7091,N_4078,N_4539);
nor U7092 (N_7092,N_4408,N_5280);
and U7093 (N_7093,N_5803,N_5481);
nor U7094 (N_7094,N_4305,N_5332);
xor U7095 (N_7095,N_5364,N_5667);
nor U7096 (N_7096,N_4441,N_5997);
nand U7097 (N_7097,N_5346,N_5778);
xor U7098 (N_7098,N_5565,N_5357);
xnor U7099 (N_7099,N_5872,N_4994);
nand U7100 (N_7100,N_5343,N_5064);
and U7101 (N_7101,N_5281,N_4290);
nand U7102 (N_7102,N_4929,N_5581);
and U7103 (N_7103,N_4005,N_5337);
and U7104 (N_7104,N_5176,N_5217);
nor U7105 (N_7105,N_5775,N_4792);
xor U7106 (N_7106,N_5174,N_5949);
or U7107 (N_7107,N_4542,N_5489);
nor U7108 (N_7108,N_4270,N_5025);
and U7109 (N_7109,N_5418,N_5534);
or U7110 (N_7110,N_4983,N_5422);
or U7111 (N_7111,N_5238,N_5073);
nand U7112 (N_7112,N_5084,N_5543);
xnor U7113 (N_7113,N_4832,N_5607);
nand U7114 (N_7114,N_5330,N_5630);
or U7115 (N_7115,N_4572,N_4833);
nand U7116 (N_7116,N_4457,N_5195);
nor U7117 (N_7117,N_5543,N_5940);
nand U7118 (N_7118,N_5484,N_4422);
nand U7119 (N_7119,N_4241,N_5735);
or U7120 (N_7120,N_5880,N_5569);
nand U7121 (N_7121,N_4397,N_4624);
and U7122 (N_7122,N_4126,N_5864);
nor U7123 (N_7123,N_4387,N_5086);
or U7124 (N_7124,N_4522,N_5715);
and U7125 (N_7125,N_4721,N_5129);
nor U7126 (N_7126,N_5760,N_5628);
nor U7127 (N_7127,N_5440,N_4263);
and U7128 (N_7128,N_4088,N_4124);
or U7129 (N_7129,N_4487,N_4218);
nand U7130 (N_7130,N_5797,N_5243);
xor U7131 (N_7131,N_4700,N_5498);
or U7132 (N_7132,N_4779,N_5609);
nor U7133 (N_7133,N_5197,N_5996);
or U7134 (N_7134,N_5480,N_4706);
nor U7135 (N_7135,N_4433,N_5815);
xor U7136 (N_7136,N_5292,N_4728);
nor U7137 (N_7137,N_5136,N_4618);
nand U7138 (N_7138,N_5741,N_4680);
xor U7139 (N_7139,N_5320,N_5076);
or U7140 (N_7140,N_4986,N_4993);
and U7141 (N_7141,N_5435,N_5364);
nor U7142 (N_7142,N_5362,N_4680);
nand U7143 (N_7143,N_5924,N_4333);
or U7144 (N_7144,N_4849,N_5720);
xor U7145 (N_7145,N_5281,N_5183);
nand U7146 (N_7146,N_4506,N_5034);
nor U7147 (N_7147,N_4731,N_4083);
or U7148 (N_7148,N_5932,N_5140);
nand U7149 (N_7149,N_4468,N_5889);
and U7150 (N_7150,N_5651,N_5902);
nor U7151 (N_7151,N_5052,N_4712);
nand U7152 (N_7152,N_5409,N_5431);
and U7153 (N_7153,N_4666,N_5520);
or U7154 (N_7154,N_5467,N_4988);
nand U7155 (N_7155,N_4166,N_5213);
nand U7156 (N_7156,N_5916,N_5542);
xnor U7157 (N_7157,N_4960,N_4553);
and U7158 (N_7158,N_5629,N_4228);
nor U7159 (N_7159,N_4375,N_4649);
nor U7160 (N_7160,N_4325,N_5705);
nor U7161 (N_7161,N_5333,N_4942);
nand U7162 (N_7162,N_4479,N_5014);
xor U7163 (N_7163,N_4324,N_4789);
and U7164 (N_7164,N_4722,N_5716);
nand U7165 (N_7165,N_4966,N_4900);
or U7166 (N_7166,N_4254,N_5446);
nand U7167 (N_7167,N_4635,N_5417);
and U7168 (N_7168,N_5175,N_4291);
or U7169 (N_7169,N_4053,N_5711);
nand U7170 (N_7170,N_5596,N_4959);
xnor U7171 (N_7171,N_4744,N_5933);
nand U7172 (N_7172,N_5137,N_5685);
nand U7173 (N_7173,N_4188,N_4880);
nand U7174 (N_7174,N_5585,N_4499);
and U7175 (N_7175,N_4921,N_4117);
or U7176 (N_7176,N_4523,N_4976);
or U7177 (N_7177,N_4575,N_4712);
and U7178 (N_7178,N_5646,N_4924);
nor U7179 (N_7179,N_4915,N_5582);
xor U7180 (N_7180,N_5338,N_5289);
and U7181 (N_7181,N_4401,N_4465);
and U7182 (N_7182,N_4284,N_4400);
and U7183 (N_7183,N_5033,N_4594);
nand U7184 (N_7184,N_5995,N_5442);
nand U7185 (N_7185,N_4788,N_5238);
nor U7186 (N_7186,N_4896,N_4265);
xnor U7187 (N_7187,N_5095,N_4011);
nor U7188 (N_7188,N_4284,N_5109);
nor U7189 (N_7189,N_4782,N_5785);
nor U7190 (N_7190,N_4568,N_4862);
xnor U7191 (N_7191,N_5542,N_4290);
and U7192 (N_7192,N_4735,N_4697);
and U7193 (N_7193,N_5145,N_5285);
xor U7194 (N_7194,N_4354,N_5653);
or U7195 (N_7195,N_5948,N_5992);
and U7196 (N_7196,N_5793,N_5582);
xnor U7197 (N_7197,N_4351,N_4010);
and U7198 (N_7198,N_4493,N_5977);
nand U7199 (N_7199,N_5985,N_4921);
nor U7200 (N_7200,N_5051,N_5521);
and U7201 (N_7201,N_4186,N_4034);
nor U7202 (N_7202,N_4089,N_4328);
nand U7203 (N_7203,N_4922,N_4517);
nand U7204 (N_7204,N_4981,N_5533);
nand U7205 (N_7205,N_4104,N_4066);
nand U7206 (N_7206,N_5816,N_4169);
nor U7207 (N_7207,N_5731,N_4656);
and U7208 (N_7208,N_4610,N_4771);
nand U7209 (N_7209,N_4148,N_5260);
xnor U7210 (N_7210,N_5564,N_4747);
nand U7211 (N_7211,N_5991,N_4588);
and U7212 (N_7212,N_4923,N_5299);
and U7213 (N_7213,N_5338,N_5762);
and U7214 (N_7214,N_4750,N_5356);
nor U7215 (N_7215,N_5092,N_4685);
or U7216 (N_7216,N_5459,N_4956);
and U7217 (N_7217,N_4508,N_4749);
and U7218 (N_7218,N_5909,N_4723);
or U7219 (N_7219,N_4234,N_5448);
and U7220 (N_7220,N_5270,N_4312);
and U7221 (N_7221,N_5681,N_4109);
nor U7222 (N_7222,N_4730,N_4752);
or U7223 (N_7223,N_5681,N_5141);
and U7224 (N_7224,N_4910,N_4412);
or U7225 (N_7225,N_4028,N_4159);
nand U7226 (N_7226,N_5527,N_5235);
xnor U7227 (N_7227,N_4269,N_5274);
nand U7228 (N_7228,N_4605,N_4227);
nand U7229 (N_7229,N_4624,N_4650);
and U7230 (N_7230,N_5694,N_4067);
or U7231 (N_7231,N_5743,N_4175);
or U7232 (N_7232,N_5086,N_5548);
nor U7233 (N_7233,N_4383,N_5366);
nor U7234 (N_7234,N_4136,N_4050);
nor U7235 (N_7235,N_5889,N_4451);
or U7236 (N_7236,N_4836,N_4612);
or U7237 (N_7237,N_5997,N_5123);
nand U7238 (N_7238,N_5595,N_5012);
nand U7239 (N_7239,N_5556,N_5723);
nor U7240 (N_7240,N_4538,N_4167);
and U7241 (N_7241,N_4522,N_5895);
or U7242 (N_7242,N_4414,N_5225);
nand U7243 (N_7243,N_4136,N_4392);
and U7244 (N_7244,N_4792,N_4697);
or U7245 (N_7245,N_4174,N_4773);
nand U7246 (N_7246,N_4617,N_5534);
nand U7247 (N_7247,N_4688,N_5622);
nor U7248 (N_7248,N_5489,N_4899);
xnor U7249 (N_7249,N_4918,N_4707);
nand U7250 (N_7250,N_4687,N_4272);
xnor U7251 (N_7251,N_5829,N_4211);
and U7252 (N_7252,N_4972,N_4943);
and U7253 (N_7253,N_4373,N_5784);
nand U7254 (N_7254,N_4773,N_5085);
nand U7255 (N_7255,N_5609,N_5926);
xor U7256 (N_7256,N_4183,N_4650);
or U7257 (N_7257,N_4784,N_5714);
nor U7258 (N_7258,N_4634,N_4305);
or U7259 (N_7259,N_4308,N_4824);
and U7260 (N_7260,N_5208,N_4506);
nand U7261 (N_7261,N_4339,N_4458);
and U7262 (N_7262,N_4269,N_4799);
nand U7263 (N_7263,N_5628,N_5067);
nand U7264 (N_7264,N_4444,N_4477);
nand U7265 (N_7265,N_5238,N_5620);
nor U7266 (N_7266,N_4899,N_5677);
or U7267 (N_7267,N_4793,N_4381);
nor U7268 (N_7268,N_5463,N_5982);
nand U7269 (N_7269,N_4484,N_4194);
or U7270 (N_7270,N_5631,N_4015);
nand U7271 (N_7271,N_5698,N_4469);
nor U7272 (N_7272,N_5275,N_5313);
xor U7273 (N_7273,N_5717,N_4573);
nand U7274 (N_7274,N_4274,N_5217);
xnor U7275 (N_7275,N_4556,N_5948);
and U7276 (N_7276,N_4035,N_4892);
or U7277 (N_7277,N_4276,N_5755);
or U7278 (N_7278,N_5375,N_4894);
xor U7279 (N_7279,N_5602,N_5258);
and U7280 (N_7280,N_5027,N_5622);
and U7281 (N_7281,N_4963,N_4392);
nand U7282 (N_7282,N_4576,N_5527);
and U7283 (N_7283,N_5097,N_4822);
nand U7284 (N_7284,N_4512,N_5369);
and U7285 (N_7285,N_4258,N_5077);
nand U7286 (N_7286,N_5279,N_4045);
nand U7287 (N_7287,N_4177,N_5195);
xnor U7288 (N_7288,N_4085,N_5176);
or U7289 (N_7289,N_4974,N_5810);
nor U7290 (N_7290,N_5197,N_5355);
xor U7291 (N_7291,N_4249,N_5502);
or U7292 (N_7292,N_5584,N_5941);
or U7293 (N_7293,N_4939,N_5721);
nand U7294 (N_7294,N_5836,N_4130);
or U7295 (N_7295,N_4475,N_4204);
and U7296 (N_7296,N_5714,N_4334);
or U7297 (N_7297,N_4855,N_4999);
nand U7298 (N_7298,N_4062,N_5358);
or U7299 (N_7299,N_4830,N_5245);
or U7300 (N_7300,N_5884,N_4727);
nand U7301 (N_7301,N_4520,N_5438);
nor U7302 (N_7302,N_5962,N_4711);
or U7303 (N_7303,N_4935,N_5844);
nand U7304 (N_7304,N_5502,N_5920);
nor U7305 (N_7305,N_4340,N_5883);
or U7306 (N_7306,N_5358,N_5609);
nand U7307 (N_7307,N_5938,N_4510);
and U7308 (N_7308,N_5397,N_5871);
and U7309 (N_7309,N_4997,N_4531);
and U7310 (N_7310,N_5308,N_4067);
nand U7311 (N_7311,N_5733,N_4241);
and U7312 (N_7312,N_4688,N_4306);
nor U7313 (N_7313,N_4858,N_5774);
and U7314 (N_7314,N_5429,N_5498);
nand U7315 (N_7315,N_5525,N_5208);
or U7316 (N_7316,N_4697,N_4124);
xnor U7317 (N_7317,N_4986,N_5573);
or U7318 (N_7318,N_5377,N_5925);
and U7319 (N_7319,N_5100,N_4203);
nand U7320 (N_7320,N_4354,N_4766);
xnor U7321 (N_7321,N_5817,N_5502);
and U7322 (N_7322,N_4080,N_5572);
and U7323 (N_7323,N_5593,N_5800);
xor U7324 (N_7324,N_5484,N_4130);
xor U7325 (N_7325,N_5986,N_4614);
nand U7326 (N_7326,N_4112,N_5092);
nor U7327 (N_7327,N_4243,N_4072);
and U7328 (N_7328,N_5479,N_5272);
or U7329 (N_7329,N_5026,N_4258);
nor U7330 (N_7330,N_5994,N_5953);
nor U7331 (N_7331,N_5213,N_4510);
and U7332 (N_7332,N_5428,N_4094);
or U7333 (N_7333,N_5776,N_4634);
or U7334 (N_7334,N_5743,N_4543);
nand U7335 (N_7335,N_4969,N_4181);
nor U7336 (N_7336,N_5155,N_5606);
or U7337 (N_7337,N_5781,N_4288);
and U7338 (N_7338,N_5503,N_5577);
or U7339 (N_7339,N_4394,N_4059);
nor U7340 (N_7340,N_4196,N_4024);
or U7341 (N_7341,N_5858,N_4554);
nor U7342 (N_7342,N_4984,N_5075);
or U7343 (N_7343,N_5064,N_4689);
or U7344 (N_7344,N_5498,N_4536);
nand U7345 (N_7345,N_5995,N_4686);
nand U7346 (N_7346,N_5970,N_5656);
or U7347 (N_7347,N_4710,N_4498);
xnor U7348 (N_7348,N_4860,N_5746);
xnor U7349 (N_7349,N_5430,N_4917);
or U7350 (N_7350,N_5468,N_4928);
nand U7351 (N_7351,N_5923,N_4858);
nand U7352 (N_7352,N_5447,N_5806);
nand U7353 (N_7353,N_4250,N_4256);
nor U7354 (N_7354,N_4211,N_5297);
nor U7355 (N_7355,N_4447,N_5009);
or U7356 (N_7356,N_4870,N_4454);
nand U7357 (N_7357,N_5731,N_5257);
or U7358 (N_7358,N_4095,N_5818);
or U7359 (N_7359,N_5429,N_4514);
xnor U7360 (N_7360,N_5130,N_4886);
or U7361 (N_7361,N_5853,N_5969);
and U7362 (N_7362,N_4185,N_4679);
xor U7363 (N_7363,N_4706,N_4968);
nand U7364 (N_7364,N_5011,N_5127);
nor U7365 (N_7365,N_5081,N_4396);
nor U7366 (N_7366,N_4988,N_4817);
nor U7367 (N_7367,N_5492,N_4234);
or U7368 (N_7368,N_4974,N_5690);
xnor U7369 (N_7369,N_4515,N_4610);
or U7370 (N_7370,N_4871,N_4866);
xor U7371 (N_7371,N_5847,N_4865);
and U7372 (N_7372,N_5555,N_4591);
nand U7373 (N_7373,N_5210,N_4517);
nand U7374 (N_7374,N_4319,N_5363);
nor U7375 (N_7375,N_5407,N_5449);
nand U7376 (N_7376,N_5976,N_5725);
nand U7377 (N_7377,N_4125,N_5205);
xor U7378 (N_7378,N_4447,N_4106);
and U7379 (N_7379,N_4025,N_5827);
or U7380 (N_7380,N_4324,N_4582);
or U7381 (N_7381,N_4697,N_4643);
nand U7382 (N_7382,N_4716,N_4601);
nand U7383 (N_7383,N_4904,N_4070);
or U7384 (N_7384,N_5508,N_5893);
nor U7385 (N_7385,N_4389,N_4642);
nor U7386 (N_7386,N_4217,N_5193);
xnor U7387 (N_7387,N_4280,N_4187);
and U7388 (N_7388,N_5679,N_4860);
nor U7389 (N_7389,N_5607,N_5111);
nand U7390 (N_7390,N_4716,N_5169);
and U7391 (N_7391,N_4382,N_5971);
nand U7392 (N_7392,N_4763,N_4175);
and U7393 (N_7393,N_5222,N_5849);
nand U7394 (N_7394,N_4234,N_4924);
and U7395 (N_7395,N_4985,N_5548);
and U7396 (N_7396,N_5922,N_5653);
nor U7397 (N_7397,N_4392,N_5079);
nand U7398 (N_7398,N_4599,N_4339);
nand U7399 (N_7399,N_5650,N_4824);
or U7400 (N_7400,N_5299,N_5190);
nor U7401 (N_7401,N_5406,N_4910);
nor U7402 (N_7402,N_4838,N_4325);
and U7403 (N_7403,N_5282,N_4084);
nand U7404 (N_7404,N_5980,N_5427);
xnor U7405 (N_7405,N_5948,N_4501);
nand U7406 (N_7406,N_4291,N_4855);
and U7407 (N_7407,N_5874,N_5429);
or U7408 (N_7408,N_5158,N_4848);
and U7409 (N_7409,N_4714,N_5965);
nor U7410 (N_7410,N_5392,N_4479);
xnor U7411 (N_7411,N_5143,N_5976);
and U7412 (N_7412,N_4887,N_5861);
and U7413 (N_7413,N_4714,N_5953);
nor U7414 (N_7414,N_5415,N_4769);
nor U7415 (N_7415,N_4930,N_4599);
xor U7416 (N_7416,N_4451,N_5629);
or U7417 (N_7417,N_4004,N_5936);
nor U7418 (N_7418,N_4721,N_5858);
and U7419 (N_7419,N_5587,N_4974);
and U7420 (N_7420,N_4337,N_5352);
or U7421 (N_7421,N_4685,N_4449);
or U7422 (N_7422,N_5874,N_4845);
or U7423 (N_7423,N_5544,N_4456);
or U7424 (N_7424,N_4988,N_5979);
or U7425 (N_7425,N_5840,N_5737);
nand U7426 (N_7426,N_5935,N_4224);
nor U7427 (N_7427,N_4131,N_5371);
and U7428 (N_7428,N_4401,N_5188);
nor U7429 (N_7429,N_4929,N_5678);
nand U7430 (N_7430,N_4217,N_4174);
and U7431 (N_7431,N_4894,N_5515);
or U7432 (N_7432,N_4070,N_5243);
or U7433 (N_7433,N_5836,N_4846);
or U7434 (N_7434,N_4194,N_5071);
nand U7435 (N_7435,N_4704,N_4457);
or U7436 (N_7436,N_5580,N_4964);
nor U7437 (N_7437,N_4047,N_5949);
nor U7438 (N_7438,N_4059,N_5121);
and U7439 (N_7439,N_5816,N_5964);
or U7440 (N_7440,N_5947,N_5790);
nand U7441 (N_7441,N_4001,N_4015);
nor U7442 (N_7442,N_5175,N_5456);
or U7443 (N_7443,N_4237,N_5891);
or U7444 (N_7444,N_5289,N_5433);
or U7445 (N_7445,N_5358,N_5549);
xnor U7446 (N_7446,N_4601,N_4025);
and U7447 (N_7447,N_4817,N_5154);
and U7448 (N_7448,N_4063,N_4501);
or U7449 (N_7449,N_5986,N_5720);
or U7450 (N_7450,N_4561,N_4240);
nor U7451 (N_7451,N_5796,N_5785);
nand U7452 (N_7452,N_4629,N_5644);
nand U7453 (N_7453,N_5862,N_4418);
and U7454 (N_7454,N_4245,N_5952);
nor U7455 (N_7455,N_5370,N_5309);
and U7456 (N_7456,N_5064,N_5821);
and U7457 (N_7457,N_5694,N_5684);
nand U7458 (N_7458,N_5527,N_4405);
or U7459 (N_7459,N_4970,N_5475);
or U7460 (N_7460,N_5315,N_5553);
xnor U7461 (N_7461,N_4639,N_4594);
and U7462 (N_7462,N_4532,N_5005);
nand U7463 (N_7463,N_5175,N_4666);
nand U7464 (N_7464,N_5331,N_4967);
and U7465 (N_7465,N_5477,N_5088);
and U7466 (N_7466,N_5494,N_4670);
and U7467 (N_7467,N_5530,N_4754);
nand U7468 (N_7468,N_4925,N_5676);
xor U7469 (N_7469,N_4589,N_5774);
nand U7470 (N_7470,N_5535,N_5777);
and U7471 (N_7471,N_4569,N_5132);
nor U7472 (N_7472,N_5835,N_4005);
nand U7473 (N_7473,N_4090,N_4761);
nor U7474 (N_7474,N_4235,N_4918);
and U7475 (N_7475,N_4714,N_4556);
or U7476 (N_7476,N_4799,N_5879);
nand U7477 (N_7477,N_4980,N_5889);
or U7478 (N_7478,N_5832,N_4831);
and U7479 (N_7479,N_5115,N_5512);
nand U7480 (N_7480,N_5100,N_5894);
nor U7481 (N_7481,N_5166,N_5532);
xnor U7482 (N_7482,N_4844,N_5640);
nor U7483 (N_7483,N_4222,N_5580);
nand U7484 (N_7484,N_4691,N_4386);
and U7485 (N_7485,N_5897,N_5530);
nor U7486 (N_7486,N_5644,N_5713);
and U7487 (N_7487,N_5720,N_4591);
nor U7488 (N_7488,N_5945,N_4620);
and U7489 (N_7489,N_5920,N_5301);
and U7490 (N_7490,N_4849,N_4122);
nand U7491 (N_7491,N_4149,N_4983);
nand U7492 (N_7492,N_5481,N_4927);
and U7493 (N_7493,N_4178,N_5373);
nand U7494 (N_7494,N_4708,N_4307);
and U7495 (N_7495,N_5387,N_5678);
nand U7496 (N_7496,N_5476,N_4940);
nor U7497 (N_7497,N_5924,N_4644);
nor U7498 (N_7498,N_5751,N_4410);
nor U7499 (N_7499,N_5764,N_4369);
and U7500 (N_7500,N_4311,N_4675);
or U7501 (N_7501,N_4772,N_4172);
and U7502 (N_7502,N_4904,N_5093);
nand U7503 (N_7503,N_4418,N_5935);
xor U7504 (N_7504,N_4026,N_4232);
nor U7505 (N_7505,N_4151,N_4400);
nor U7506 (N_7506,N_5461,N_5529);
or U7507 (N_7507,N_5865,N_4132);
or U7508 (N_7508,N_4194,N_4278);
nand U7509 (N_7509,N_5639,N_4069);
nand U7510 (N_7510,N_5465,N_4205);
nand U7511 (N_7511,N_5861,N_4161);
nand U7512 (N_7512,N_5248,N_4305);
nor U7513 (N_7513,N_5277,N_4715);
or U7514 (N_7514,N_5757,N_4965);
or U7515 (N_7515,N_5764,N_5072);
or U7516 (N_7516,N_4102,N_5709);
and U7517 (N_7517,N_4862,N_4573);
nand U7518 (N_7518,N_4028,N_4980);
xor U7519 (N_7519,N_4573,N_4731);
nor U7520 (N_7520,N_5047,N_4662);
and U7521 (N_7521,N_4310,N_4270);
nor U7522 (N_7522,N_4562,N_5288);
or U7523 (N_7523,N_5092,N_4839);
nand U7524 (N_7524,N_5380,N_4567);
nor U7525 (N_7525,N_5516,N_4846);
and U7526 (N_7526,N_4124,N_4696);
and U7527 (N_7527,N_5193,N_5298);
nor U7528 (N_7528,N_5870,N_5810);
and U7529 (N_7529,N_5861,N_5552);
and U7530 (N_7530,N_4637,N_5768);
and U7531 (N_7531,N_4084,N_4236);
xor U7532 (N_7532,N_4526,N_4894);
nand U7533 (N_7533,N_4142,N_5532);
and U7534 (N_7534,N_5663,N_4568);
and U7535 (N_7535,N_5250,N_4022);
nor U7536 (N_7536,N_4736,N_5268);
xor U7537 (N_7537,N_5753,N_5261);
xor U7538 (N_7538,N_5855,N_4521);
nand U7539 (N_7539,N_4674,N_4238);
nor U7540 (N_7540,N_4087,N_4445);
nand U7541 (N_7541,N_4704,N_4728);
nand U7542 (N_7542,N_4756,N_5449);
and U7543 (N_7543,N_5538,N_4064);
nand U7544 (N_7544,N_5929,N_5310);
nand U7545 (N_7545,N_4036,N_4566);
nor U7546 (N_7546,N_5773,N_4043);
and U7547 (N_7547,N_4802,N_4939);
nor U7548 (N_7548,N_4400,N_5767);
nor U7549 (N_7549,N_4529,N_5298);
nor U7550 (N_7550,N_4144,N_4067);
or U7551 (N_7551,N_4889,N_4405);
nand U7552 (N_7552,N_5035,N_4675);
xnor U7553 (N_7553,N_5796,N_5213);
xnor U7554 (N_7554,N_4956,N_4735);
and U7555 (N_7555,N_5977,N_4004);
or U7556 (N_7556,N_4657,N_5921);
nor U7557 (N_7557,N_4017,N_5812);
and U7558 (N_7558,N_4828,N_4771);
xor U7559 (N_7559,N_4483,N_4926);
xor U7560 (N_7560,N_4058,N_5420);
nand U7561 (N_7561,N_4075,N_4279);
xnor U7562 (N_7562,N_5636,N_4726);
nor U7563 (N_7563,N_5132,N_5002);
and U7564 (N_7564,N_4080,N_4975);
nand U7565 (N_7565,N_4501,N_5233);
xor U7566 (N_7566,N_5388,N_4038);
xnor U7567 (N_7567,N_4947,N_4352);
and U7568 (N_7568,N_5787,N_4179);
xnor U7569 (N_7569,N_5004,N_4592);
nand U7570 (N_7570,N_4888,N_4113);
nand U7571 (N_7571,N_5127,N_5543);
and U7572 (N_7572,N_4120,N_5163);
nor U7573 (N_7573,N_4303,N_4425);
or U7574 (N_7574,N_5372,N_4580);
or U7575 (N_7575,N_4498,N_5085);
and U7576 (N_7576,N_4145,N_5715);
nand U7577 (N_7577,N_4509,N_5669);
and U7578 (N_7578,N_4146,N_5389);
nand U7579 (N_7579,N_4475,N_5903);
xor U7580 (N_7580,N_5656,N_4958);
nor U7581 (N_7581,N_4718,N_4913);
nand U7582 (N_7582,N_4339,N_5738);
nand U7583 (N_7583,N_5726,N_5680);
nor U7584 (N_7584,N_5123,N_5729);
and U7585 (N_7585,N_4376,N_4425);
or U7586 (N_7586,N_5396,N_4378);
xnor U7587 (N_7587,N_5046,N_4144);
nor U7588 (N_7588,N_4533,N_4544);
and U7589 (N_7589,N_5155,N_5482);
and U7590 (N_7590,N_4697,N_4261);
nand U7591 (N_7591,N_5630,N_5669);
nor U7592 (N_7592,N_5290,N_5601);
nand U7593 (N_7593,N_5673,N_4485);
nor U7594 (N_7594,N_5757,N_5201);
or U7595 (N_7595,N_5828,N_5286);
nor U7596 (N_7596,N_4933,N_4875);
nor U7597 (N_7597,N_5800,N_5168);
or U7598 (N_7598,N_5504,N_5910);
nor U7599 (N_7599,N_4309,N_4420);
xnor U7600 (N_7600,N_5803,N_4832);
and U7601 (N_7601,N_5412,N_5242);
or U7602 (N_7602,N_5028,N_4248);
nand U7603 (N_7603,N_5562,N_5212);
or U7604 (N_7604,N_5330,N_4758);
and U7605 (N_7605,N_4885,N_5057);
nand U7606 (N_7606,N_4087,N_4798);
nand U7607 (N_7607,N_4770,N_4516);
or U7608 (N_7608,N_5615,N_5902);
or U7609 (N_7609,N_4527,N_5618);
or U7610 (N_7610,N_5542,N_5125);
or U7611 (N_7611,N_4828,N_4113);
or U7612 (N_7612,N_5083,N_4328);
nor U7613 (N_7613,N_4525,N_4235);
and U7614 (N_7614,N_4967,N_5892);
nand U7615 (N_7615,N_5191,N_4170);
and U7616 (N_7616,N_4639,N_5193);
nand U7617 (N_7617,N_5147,N_5817);
or U7618 (N_7618,N_5635,N_5985);
and U7619 (N_7619,N_4157,N_4939);
nand U7620 (N_7620,N_4975,N_4759);
nor U7621 (N_7621,N_5433,N_5857);
xnor U7622 (N_7622,N_5908,N_4839);
or U7623 (N_7623,N_5804,N_4392);
and U7624 (N_7624,N_5208,N_5989);
or U7625 (N_7625,N_5651,N_4281);
and U7626 (N_7626,N_5461,N_5997);
and U7627 (N_7627,N_5607,N_5639);
nand U7628 (N_7628,N_5348,N_4596);
and U7629 (N_7629,N_5926,N_5818);
nand U7630 (N_7630,N_5739,N_4962);
and U7631 (N_7631,N_5025,N_5557);
and U7632 (N_7632,N_5954,N_5955);
nor U7633 (N_7633,N_4366,N_4220);
nand U7634 (N_7634,N_5456,N_4363);
and U7635 (N_7635,N_5518,N_5896);
nand U7636 (N_7636,N_4199,N_5100);
nand U7637 (N_7637,N_5836,N_5665);
or U7638 (N_7638,N_5249,N_5258);
and U7639 (N_7639,N_4491,N_4543);
nor U7640 (N_7640,N_4968,N_5651);
nand U7641 (N_7641,N_5929,N_4888);
xor U7642 (N_7642,N_5569,N_5838);
nand U7643 (N_7643,N_4373,N_4443);
nand U7644 (N_7644,N_5571,N_4095);
or U7645 (N_7645,N_5815,N_5291);
nor U7646 (N_7646,N_4850,N_5454);
and U7647 (N_7647,N_4346,N_5161);
or U7648 (N_7648,N_5011,N_4920);
and U7649 (N_7649,N_4860,N_5522);
nand U7650 (N_7650,N_4817,N_5975);
or U7651 (N_7651,N_4883,N_4858);
nand U7652 (N_7652,N_5113,N_5292);
or U7653 (N_7653,N_5518,N_4730);
nor U7654 (N_7654,N_5799,N_4971);
nor U7655 (N_7655,N_4909,N_5721);
and U7656 (N_7656,N_4262,N_5855);
or U7657 (N_7657,N_4364,N_5252);
xor U7658 (N_7658,N_4493,N_4344);
and U7659 (N_7659,N_5363,N_5152);
nor U7660 (N_7660,N_4693,N_4414);
xor U7661 (N_7661,N_4106,N_4842);
or U7662 (N_7662,N_4835,N_4091);
nand U7663 (N_7663,N_4564,N_5200);
or U7664 (N_7664,N_4778,N_4245);
nor U7665 (N_7665,N_4766,N_4063);
or U7666 (N_7666,N_4692,N_5399);
nand U7667 (N_7667,N_5442,N_5906);
nor U7668 (N_7668,N_4848,N_5553);
or U7669 (N_7669,N_5179,N_5437);
nand U7670 (N_7670,N_5040,N_4985);
or U7671 (N_7671,N_5600,N_5524);
or U7672 (N_7672,N_4735,N_4903);
nand U7673 (N_7673,N_4367,N_5521);
xnor U7674 (N_7674,N_5118,N_5571);
nand U7675 (N_7675,N_4717,N_4986);
nor U7676 (N_7676,N_5429,N_5129);
or U7677 (N_7677,N_4346,N_5271);
nor U7678 (N_7678,N_5210,N_5681);
xor U7679 (N_7679,N_5063,N_5629);
nand U7680 (N_7680,N_4724,N_5370);
nand U7681 (N_7681,N_5076,N_4377);
nand U7682 (N_7682,N_5664,N_5459);
or U7683 (N_7683,N_4357,N_5056);
or U7684 (N_7684,N_4154,N_5615);
or U7685 (N_7685,N_4379,N_5198);
and U7686 (N_7686,N_4136,N_4821);
and U7687 (N_7687,N_4828,N_5106);
nor U7688 (N_7688,N_5948,N_4590);
xnor U7689 (N_7689,N_4938,N_4591);
or U7690 (N_7690,N_4930,N_5647);
or U7691 (N_7691,N_4233,N_5656);
or U7692 (N_7692,N_5551,N_5563);
nand U7693 (N_7693,N_5796,N_4237);
nand U7694 (N_7694,N_5292,N_4991);
xnor U7695 (N_7695,N_4472,N_4695);
or U7696 (N_7696,N_5895,N_5965);
or U7697 (N_7697,N_5722,N_4307);
and U7698 (N_7698,N_5528,N_4559);
nor U7699 (N_7699,N_5341,N_5184);
or U7700 (N_7700,N_4967,N_5690);
or U7701 (N_7701,N_4238,N_5283);
nand U7702 (N_7702,N_5803,N_5003);
and U7703 (N_7703,N_4052,N_4515);
or U7704 (N_7704,N_5384,N_5417);
nor U7705 (N_7705,N_5613,N_4543);
nor U7706 (N_7706,N_4147,N_5670);
xnor U7707 (N_7707,N_4905,N_5503);
nand U7708 (N_7708,N_4160,N_5604);
nand U7709 (N_7709,N_5950,N_5363);
nor U7710 (N_7710,N_5708,N_4445);
xnor U7711 (N_7711,N_5012,N_4052);
nand U7712 (N_7712,N_4873,N_4920);
or U7713 (N_7713,N_4624,N_4147);
or U7714 (N_7714,N_5033,N_5041);
nand U7715 (N_7715,N_4220,N_5422);
and U7716 (N_7716,N_4145,N_5932);
xor U7717 (N_7717,N_4712,N_4448);
nand U7718 (N_7718,N_4275,N_5339);
nand U7719 (N_7719,N_4747,N_5622);
nor U7720 (N_7720,N_4027,N_5335);
and U7721 (N_7721,N_4277,N_4707);
or U7722 (N_7722,N_4757,N_5981);
and U7723 (N_7723,N_5919,N_4382);
or U7724 (N_7724,N_5792,N_4144);
nand U7725 (N_7725,N_4229,N_5074);
and U7726 (N_7726,N_4030,N_5258);
nor U7727 (N_7727,N_5810,N_5514);
xnor U7728 (N_7728,N_5479,N_5206);
xnor U7729 (N_7729,N_5081,N_5409);
nor U7730 (N_7730,N_5624,N_5122);
nand U7731 (N_7731,N_5275,N_5383);
and U7732 (N_7732,N_5694,N_4814);
xnor U7733 (N_7733,N_4753,N_5552);
nand U7734 (N_7734,N_4548,N_4248);
and U7735 (N_7735,N_5978,N_5094);
nor U7736 (N_7736,N_4460,N_4141);
xor U7737 (N_7737,N_4633,N_5919);
nand U7738 (N_7738,N_4805,N_4849);
or U7739 (N_7739,N_5040,N_5995);
nor U7740 (N_7740,N_5360,N_4142);
nand U7741 (N_7741,N_4706,N_4434);
nor U7742 (N_7742,N_5479,N_5291);
xor U7743 (N_7743,N_5782,N_5070);
nor U7744 (N_7744,N_4897,N_4264);
nand U7745 (N_7745,N_5339,N_5640);
nand U7746 (N_7746,N_4737,N_4317);
nor U7747 (N_7747,N_4178,N_5177);
and U7748 (N_7748,N_4634,N_5744);
nand U7749 (N_7749,N_4908,N_4647);
nand U7750 (N_7750,N_4454,N_4421);
nand U7751 (N_7751,N_5351,N_4234);
nand U7752 (N_7752,N_4091,N_5020);
and U7753 (N_7753,N_5130,N_5104);
nand U7754 (N_7754,N_4162,N_4433);
nand U7755 (N_7755,N_5374,N_4371);
xor U7756 (N_7756,N_5405,N_4219);
nor U7757 (N_7757,N_5039,N_5161);
or U7758 (N_7758,N_4652,N_5605);
and U7759 (N_7759,N_5417,N_4429);
nor U7760 (N_7760,N_4264,N_5475);
or U7761 (N_7761,N_5784,N_4066);
or U7762 (N_7762,N_4739,N_4711);
or U7763 (N_7763,N_5384,N_5677);
nor U7764 (N_7764,N_4645,N_5097);
and U7765 (N_7765,N_4258,N_4801);
or U7766 (N_7766,N_4891,N_5804);
nand U7767 (N_7767,N_4692,N_4534);
nor U7768 (N_7768,N_4634,N_4140);
or U7769 (N_7769,N_5033,N_4933);
nand U7770 (N_7770,N_4792,N_5306);
nand U7771 (N_7771,N_4997,N_5457);
nor U7772 (N_7772,N_5021,N_4969);
xnor U7773 (N_7773,N_5352,N_5086);
nor U7774 (N_7774,N_4166,N_4542);
or U7775 (N_7775,N_4446,N_4176);
nand U7776 (N_7776,N_5962,N_5655);
xnor U7777 (N_7777,N_5968,N_5444);
nand U7778 (N_7778,N_5985,N_5266);
and U7779 (N_7779,N_5388,N_5022);
nand U7780 (N_7780,N_4795,N_5466);
nand U7781 (N_7781,N_4459,N_5134);
or U7782 (N_7782,N_4778,N_5363);
or U7783 (N_7783,N_5680,N_5581);
xnor U7784 (N_7784,N_4727,N_5570);
nor U7785 (N_7785,N_5394,N_5078);
nor U7786 (N_7786,N_5996,N_5606);
nand U7787 (N_7787,N_4379,N_5586);
and U7788 (N_7788,N_5621,N_4613);
nor U7789 (N_7789,N_5440,N_4640);
nor U7790 (N_7790,N_4595,N_5052);
nand U7791 (N_7791,N_4183,N_4269);
nand U7792 (N_7792,N_4213,N_4708);
nand U7793 (N_7793,N_5529,N_4147);
and U7794 (N_7794,N_4454,N_4532);
and U7795 (N_7795,N_5750,N_5914);
xnor U7796 (N_7796,N_5206,N_4181);
nor U7797 (N_7797,N_5674,N_4063);
and U7798 (N_7798,N_5979,N_5665);
xor U7799 (N_7799,N_4892,N_5319);
xnor U7800 (N_7800,N_5996,N_4254);
and U7801 (N_7801,N_5924,N_5628);
or U7802 (N_7802,N_5536,N_5489);
and U7803 (N_7803,N_5399,N_5438);
or U7804 (N_7804,N_5522,N_5775);
nand U7805 (N_7805,N_4038,N_5874);
or U7806 (N_7806,N_4885,N_5962);
and U7807 (N_7807,N_5476,N_4250);
and U7808 (N_7808,N_5677,N_5025);
nor U7809 (N_7809,N_5641,N_5984);
and U7810 (N_7810,N_4627,N_5679);
and U7811 (N_7811,N_5273,N_4930);
nor U7812 (N_7812,N_4865,N_5082);
and U7813 (N_7813,N_5049,N_4134);
xnor U7814 (N_7814,N_4503,N_4181);
or U7815 (N_7815,N_4459,N_4416);
nor U7816 (N_7816,N_5903,N_5275);
or U7817 (N_7817,N_4267,N_4817);
nand U7818 (N_7818,N_5008,N_5066);
and U7819 (N_7819,N_4615,N_4982);
nor U7820 (N_7820,N_5913,N_5928);
and U7821 (N_7821,N_5357,N_4636);
nor U7822 (N_7822,N_4237,N_5211);
nand U7823 (N_7823,N_4270,N_4340);
and U7824 (N_7824,N_4261,N_5627);
and U7825 (N_7825,N_4350,N_4831);
nand U7826 (N_7826,N_4029,N_4552);
nand U7827 (N_7827,N_4635,N_4782);
nor U7828 (N_7828,N_5959,N_4656);
xor U7829 (N_7829,N_4615,N_5274);
xor U7830 (N_7830,N_4128,N_4533);
nor U7831 (N_7831,N_4150,N_5667);
or U7832 (N_7832,N_5469,N_5672);
nor U7833 (N_7833,N_5471,N_4800);
or U7834 (N_7834,N_4590,N_5472);
xnor U7835 (N_7835,N_4164,N_4801);
nand U7836 (N_7836,N_5477,N_5028);
nor U7837 (N_7837,N_4465,N_4165);
xor U7838 (N_7838,N_5154,N_5957);
nand U7839 (N_7839,N_4584,N_4423);
or U7840 (N_7840,N_4650,N_4592);
and U7841 (N_7841,N_5852,N_5468);
and U7842 (N_7842,N_4346,N_4850);
nand U7843 (N_7843,N_5275,N_4212);
nor U7844 (N_7844,N_5023,N_5664);
nand U7845 (N_7845,N_4599,N_4522);
xor U7846 (N_7846,N_4689,N_5261);
or U7847 (N_7847,N_4981,N_5103);
nor U7848 (N_7848,N_4168,N_4525);
nor U7849 (N_7849,N_4294,N_5979);
or U7850 (N_7850,N_5525,N_5092);
nand U7851 (N_7851,N_5426,N_5393);
nand U7852 (N_7852,N_5488,N_5281);
nor U7853 (N_7853,N_5619,N_5694);
nand U7854 (N_7854,N_5628,N_4285);
xnor U7855 (N_7855,N_5525,N_5161);
nand U7856 (N_7856,N_4361,N_5539);
nor U7857 (N_7857,N_5144,N_4909);
and U7858 (N_7858,N_4717,N_5559);
nor U7859 (N_7859,N_4791,N_4279);
nor U7860 (N_7860,N_5768,N_4080);
nand U7861 (N_7861,N_5226,N_4333);
or U7862 (N_7862,N_5456,N_4677);
nand U7863 (N_7863,N_5623,N_5259);
nor U7864 (N_7864,N_5605,N_4544);
nand U7865 (N_7865,N_4693,N_4809);
or U7866 (N_7866,N_5111,N_4848);
or U7867 (N_7867,N_4766,N_4591);
nor U7868 (N_7868,N_5013,N_5880);
and U7869 (N_7869,N_4670,N_4638);
nor U7870 (N_7870,N_5462,N_5687);
nor U7871 (N_7871,N_4192,N_5508);
nand U7872 (N_7872,N_4661,N_4428);
nand U7873 (N_7873,N_4091,N_4441);
xor U7874 (N_7874,N_5782,N_4625);
nor U7875 (N_7875,N_4135,N_4154);
and U7876 (N_7876,N_5612,N_4476);
or U7877 (N_7877,N_5969,N_4326);
nor U7878 (N_7878,N_5161,N_5648);
nor U7879 (N_7879,N_4965,N_4434);
nand U7880 (N_7880,N_4085,N_5334);
and U7881 (N_7881,N_5256,N_4922);
and U7882 (N_7882,N_5892,N_5410);
and U7883 (N_7883,N_5608,N_5855);
and U7884 (N_7884,N_4470,N_5947);
xor U7885 (N_7885,N_5981,N_5405);
nand U7886 (N_7886,N_4978,N_5135);
or U7887 (N_7887,N_4507,N_5364);
xnor U7888 (N_7888,N_4639,N_5351);
and U7889 (N_7889,N_5712,N_4355);
and U7890 (N_7890,N_5061,N_4952);
or U7891 (N_7891,N_4789,N_5692);
or U7892 (N_7892,N_5803,N_4131);
or U7893 (N_7893,N_5949,N_5491);
or U7894 (N_7894,N_5111,N_4421);
or U7895 (N_7895,N_4557,N_4627);
nand U7896 (N_7896,N_4467,N_5660);
nand U7897 (N_7897,N_5371,N_4211);
nand U7898 (N_7898,N_5507,N_5484);
nor U7899 (N_7899,N_5939,N_5698);
or U7900 (N_7900,N_4531,N_5094);
nor U7901 (N_7901,N_5436,N_4118);
nor U7902 (N_7902,N_5509,N_4119);
or U7903 (N_7903,N_4805,N_5622);
or U7904 (N_7904,N_5423,N_5614);
nor U7905 (N_7905,N_4640,N_5883);
and U7906 (N_7906,N_4047,N_4291);
and U7907 (N_7907,N_4772,N_5237);
nand U7908 (N_7908,N_5310,N_5043);
or U7909 (N_7909,N_5130,N_5153);
xnor U7910 (N_7910,N_5784,N_4843);
nand U7911 (N_7911,N_5817,N_4344);
and U7912 (N_7912,N_5107,N_5348);
or U7913 (N_7913,N_4251,N_5326);
and U7914 (N_7914,N_4351,N_4157);
and U7915 (N_7915,N_4191,N_4837);
xor U7916 (N_7916,N_5746,N_4673);
or U7917 (N_7917,N_4311,N_5443);
nor U7918 (N_7918,N_4839,N_5203);
nand U7919 (N_7919,N_4090,N_5384);
xnor U7920 (N_7920,N_5659,N_5307);
nand U7921 (N_7921,N_5820,N_5467);
nand U7922 (N_7922,N_4334,N_5121);
nor U7923 (N_7923,N_4264,N_4876);
nand U7924 (N_7924,N_4458,N_5463);
and U7925 (N_7925,N_5993,N_4116);
nor U7926 (N_7926,N_5716,N_4323);
and U7927 (N_7927,N_4362,N_4151);
or U7928 (N_7928,N_4637,N_5975);
xor U7929 (N_7929,N_4619,N_5899);
and U7930 (N_7930,N_5278,N_4313);
nand U7931 (N_7931,N_4361,N_5139);
or U7932 (N_7932,N_4865,N_4147);
nor U7933 (N_7933,N_4094,N_4725);
nor U7934 (N_7934,N_4100,N_4982);
nand U7935 (N_7935,N_4748,N_5383);
or U7936 (N_7936,N_4850,N_4062);
and U7937 (N_7937,N_4381,N_4635);
nand U7938 (N_7938,N_5205,N_4548);
and U7939 (N_7939,N_5227,N_4241);
and U7940 (N_7940,N_4480,N_5118);
nor U7941 (N_7941,N_4058,N_5593);
nor U7942 (N_7942,N_4543,N_5436);
nor U7943 (N_7943,N_4088,N_4982);
nor U7944 (N_7944,N_4442,N_5343);
nor U7945 (N_7945,N_4490,N_4944);
or U7946 (N_7946,N_5570,N_4493);
nor U7947 (N_7947,N_5887,N_4719);
or U7948 (N_7948,N_5463,N_5847);
and U7949 (N_7949,N_4314,N_5920);
nand U7950 (N_7950,N_5117,N_5644);
or U7951 (N_7951,N_4238,N_4027);
nor U7952 (N_7952,N_5716,N_4410);
nor U7953 (N_7953,N_4112,N_5157);
nor U7954 (N_7954,N_4301,N_5932);
nor U7955 (N_7955,N_4943,N_5568);
and U7956 (N_7956,N_5220,N_4241);
nand U7957 (N_7957,N_4255,N_5642);
and U7958 (N_7958,N_4132,N_5309);
or U7959 (N_7959,N_5418,N_4968);
nand U7960 (N_7960,N_4071,N_5982);
or U7961 (N_7961,N_4501,N_4396);
or U7962 (N_7962,N_5695,N_4417);
nor U7963 (N_7963,N_4730,N_5592);
or U7964 (N_7964,N_4828,N_4429);
nor U7965 (N_7965,N_4726,N_4869);
or U7966 (N_7966,N_4138,N_5704);
and U7967 (N_7967,N_4622,N_5596);
nand U7968 (N_7968,N_5790,N_5503);
and U7969 (N_7969,N_5643,N_4798);
nand U7970 (N_7970,N_5274,N_5361);
xor U7971 (N_7971,N_4971,N_4141);
and U7972 (N_7972,N_4836,N_5224);
nand U7973 (N_7973,N_5729,N_4553);
nor U7974 (N_7974,N_5096,N_5978);
and U7975 (N_7975,N_5998,N_4843);
xnor U7976 (N_7976,N_4159,N_4424);
and U7977 (N_7977,N_5785,N_5410);
nand U7978 (N_7978,N_4884,N_4266);
and U7979 (N_7979,N_4519,N_4769);
or U7980 (N_7980,N_5414,N_4489);
and U7981 (N_7981,N_4830,N_4907);
nor U7982 (N_7982,N_4376,N_5738);
xnor U7983 (N_7983,N_5258,N_5606);
nor U7984 (N_7984,N_5787,N_5225);
nor U7985 (N_7985,N_4383,N_4486);
or U7986 (N_7986,N_5580,N_4476);
or U7987 (N_7987,N_5170,N_5810);
nand U7988 (N_7988,N_5559,N_5925);
or U7989 (N_7989,N_5114,N_4262);
and U7990 (N_7990,N_4796,N_5081);
xor U7991 (N_7991,N_4810,N_5441);
or U7992 (N_7992,N_4458,N_4633);
or U7993 (N_7993,N_4941,N_4574);
nand U7994 (N_7994,N_5616,N_5338);
nand U7995 (N_7995,N_5196,N_5215);
xor U7996 (N_7996,N_4905,N_5964);
or U7997 (N_7997,N_4058,N_4422);
xnor U7998 (N_7998,N_5832,N_4884);
or U7999 (N_7999,N_4867,N_4128);
nand U8000 (N_8000,N_7084,N_6751);
nor U8001 (N_8001,N_6284,N_6255);
and U8002 (N_8002,N_7061,N_6880);
nand U8003 (N_8003,N_6786,N_7695);
nand U8004 (N_8004,N_7292,N_7488);
nor U8005 (N_8005,N_6574,N_7907);
and U8006 (N_8006,N_6458,N_7252);
or U8007 (N_8007,N_7428,N_6316);
and U8008 (N_8008,N_7881,N_7307);
or U8009 (N_8009,N_7944,N_7107);
nor U8010 (N_8010,N_6748,N_7694);
and U8011 (N_8011,N_7476,N_6913);
nor U8012 (N_8012,N_7301,N_6842);
nand U8013 (N_8013,N_7576,N_7072);
and U8014 (N_8014,N_7284,N_7261);
xor U8015 (N_8015,N_6171,N_6404);
nor U8016 (N_8016,N_7866,N_6761);
nand U8017 (N_8017,N_6460,N_7958);
nor U8018 (N_8018,N_7533,N_7677);
and U8019 (N_8019,N_7348,N_6765);
or U8020 (N_8020,N_7779,N_7721);
or U8021 (N_8021,N_6432,N_6985);
and U8022 (N_8022,N_6421,N_6799);
nand U8023 (N_8023,N_7995,N_6602);
nand U8024 (N_8024,N_6057,N_7080);
nand U8025 (N_8025,N_7420,N_6577);
or U8026 (N_8026,N_6587,N_7273);
nand U8027 (N_8027,N_7376,N_7947);
nand U8028 (N_8028,N_6904,N_7829);
or U8029 (N_8029,N_7041,N_7039);
and U8030 (N_8030,N_6716,N_6134);
nand U8031 (N_8031,N_6355,N_6506);
nor U8032 (N_8032,N_6152,N_6860);
and U8033 (N_8033,N_6031,N_6168);
xor U8034 (N_8034,N_6147,N_6244);
or U8035 (N_8035,N_6154,N_6770);
nor U8036 (N_8036,N_7042,N_7014);
nor U8037 (N_8037,N_6241,N_7153);
or U8038 (N_8038,N_6091,N_6254);
nand U8039 (N_8039,N_6320,N_6337);
nor U8040 (N_8040,N_6328,N_7063);
nand U8041 (N_8041,N_7641,N_6935);
nand U8042 (N_8042,N_6314,N_6148);
or U8043 (N_8043,N_7055,N_6085);
xnor U8044 (N_8044,N_7959,N_6215);
nor U8045 (N_8045,N_6982,N_7706);
and U8046 (N_8046,N_7492,N_7398);
and U8047 (N_8047,N_6968,N_6830);
or U8048 (N_8048,N_6219,N_6781);
nand U8049 (N_8049,N_7158,N_7358);
xor U8050 (N_8050,N_6586,N_6089);
nand U8051 (N_8051,N_7387,N_6112);
and U8052 (N_8052,N_6302,N_7154);
nor U8053 (N_8053,N_6056,N_7555);
nor U8054 (N_8054,N_7506,N_7047);
or U8055 (N_8055,N_7734,N_6654);
nor U8056 (N_8056,N_6275,N_7577);
nor U8057 (N_8057,N_6109,N_6507);
nor U8058 (N_8058,N_6005,N_7874);
nand U8059 (N_8059,N_6167,N_7513);
and U8060 (N_8060,N_6103,N_6519);
nor U8061 (N_8061,N_6657,N_7226);
or U8062 (N_8062,N_6349,N_7889);
or U8063 (N_8063,N_6995,N_6819);
nor U8064 (N_8064,N_7051,N_7361);
or U8065 (N_8065,N_6445,N_6090);
or U8066 (N_8066,N_7350,N_6868);
or U8067 (N_8067,N_7705,N_6703);
xor U8068 (N_8068,N_7174,N_6266);
or U8069 (N_8069,N_6196,N_6132);
nand U8070 (N_8070,N_6644,N_7755);
nor U8071 (N_8071,N_7128,N_7979);
nand U8072 (N_8072,N_6719,N_6382);
and U8073 (N_8073,N_6755,N_6209);
or U8074 (N_8074,N_7928,N_6508);
or U8075 (N_8075,N_6925,N_6475);
or U8076 (N_8076,N_7386,N_7535);
and U8077 (N_8077,N_6601,N_6802);
xnor U8078 (N_8078,N_6212,N_6263);
or U8079 (N_8079,N_6310,N_6652);
nor U8080 (N_8080,N_7544,N_7227);
and U8081 (N_8081,N_6386,N_7332);
nor U8082 (N_8082,N_7700,N_6502);
or U8083 (N_8083,N_7201,N_7207);
and U8084 (N_8084,N_6710,N_7383);
nor U8085 (N_8085,N_6855,N_7581);
nand U8086 (N_8086,N_6501,N_6231);
and U8087 (N_8087,N_6495,N_7624);
and U8088 (N_8088,N_7658,N_7263);
or U8089 (N_8089,N_7161,N_6608);
nor U8090 (N_8090,N_7120,N_6669);
nor U8091 (N_8091,N_6983,N_7426);
nor U8092 (N_8092,N_6564,N_6364);
nor U8093 (N_8093,N_6286,N_7208);
nand U8094 (N_8094,N_7241,N_6481);
xor U8095 (N_8095,N_7300,N_7032);
and U8096 (N_8096,N_7353,N_7841);
or U8097 (N_8097,N_7699,N_6838);
or U8098 (N_8098,N_6815,N_7186);
and U8099 (N_8099,N_7433,N_7481);
nand U8100 (N_8100,N_6332,N_6711);
or U8101 (N_8101,N_7271,N_6232);
and U8102 (N_8102,N_7642,N_7045);
nand U8103 (N_8103,N_6032,N_6008);
or U8104 (N_8104,N_6415,N_6299);
or U8105 (N_8105,N_6561,N_6324);
nor U8106 (N_8106,N_7996,N_7341);
or U8107 (N_8107,N_6172,N_7654);
nand U8108 (N_8108,N_6503,N_6156);
and U8109 (N_8109,N_6833,N_7501);
or U8110 (N_8110,N_6978,N_6185);
or U8111 (N_8111,N_6377,N_7843);
nor U8112 (N_8112,N_7598,N_7122);
or U8113 (N_8113,N_6319,N_6997);
or U8114 (N_8114,N_6537,N_7343);
or U8115 (N_8115,N_7693,N_6173);
and U8116 (N_8116,N_7758,N_7988);
nor U8117 (N_8117,N_6407,N_7251);
or U8118 (N_8118,N_7138,N_7140);
or U8119 (N_8119,N_6965,N_6006);
nor U8120 (N_8120,N_6891,N_6462);
or U8121 (N_8121,N_6028,N_6294);
or U8122 (N_8122,N_7955,N_7649);
nand U8123 (N_8123,N_6672,N_7737);
or U8124 (N_8124,N_7732,N_7751);
and U8125 (N_8125,N_7983,N_7670);
nand U8126 (N_8126,N_7421,N_7191);
nand U8127 (N_8127,N_6214,N_7038);
and U8128 (N_8128,N_6067,N_6927);
or U8129 (N_8129,N_6202,N_7452);
nand U8130 (N_8130,N_6308,N_6443);
nor U8131 (N_8131,N_7915,N_7809);
or U8132 (N_8132,N_7526,N_6246);
nand U8133 (N_8133,N_6902,N_6426);
or U8134 (N_8134,N_6225,N_6051);
nor U8135 (N_8135,N_6081,N_6914);
xnor U8136 (N_8136,N_7180,N_7612);
nand U8137 (N_8137,N_7902,N_7171);
nor U8138 (N_8138,N_7470,N_7108);
nor U8139 (N_8139,N_7026,N_7280);
nor U8140 (N_8140,N_7689,N_7089);
nor U8141 (N_8141,N_7636,N_7132);
and U8142 (N_8142,N_6516,N_7002);
nand U8143 (N_8143,N_6844,N_7805);
nor U8144 (N_8144,N_7491,N_7438);
and U8145 (N_8145,N_6182,N_6797);
nand U8146 (N_8146,N_6963,N_7363);
nand U8147 (N_8147,N_6581,N_7609);
or U8148 (N_8148,N_6964,N_6446);
nand U8149 (N_8149,N_7010,N_7976);
nand U8150 (N_8150,N_7236,N_6835);
nand U8151 (N_8151,N_7957,N_7857);
nor U8152 (N_8152,N_6151,N_6281);
and U8153 (N_8153,N_6774,N_6694);
nor U8154 (N_8154,N_6200,N_6492);
and U8155 (N_8155,N_7580,N_7659);
xnor U8156 (N_8156,N_6705,N_7033);
or U8157 (N_8157,N_7534,N_6724);
nor U8158 (N_8158,N_7401,N_6124);
nor U8159 (N_8159,N_7255,N_7901);
nand U8160 (N_8160,N_7391,N_6754);
or U8161 (N_8161,N_7244,N_6823);
and U8162 (N_8162,N_7018,N_6878);
nand U8163 (N_8163,N_7661,N_7664);
xnor U8164 (N_8164,N_7075,N_7222);
nand U8165 (N_8165,N_6230,N_7112);
or U8166 (N_8166,N_6875,N_7011);
xor U8167 (N_8167,N_7604,N_7647);
xnor U8168 (N_8168,N_6312,N_6920);
or U8169 (N_8169,N_6114,N_6846);
nor U8170 (N_8170,N_7621,N_7449);
nor U8171 (N_8171,N_6380,N_7337);
or U8172 (N_8172,N_6301,N_7774);
or U8173 (N_8173,N_7825,N_6059);
or U8174 (N_8174,N_7757,N_7672);
xor U8175 (N_8175,N_7950,N_7557);
nand U8176 (N_8176,N_6113,N_6526);
or U8177 (N_8177,N_6367,N_6276);
or U8178 (N_8178,N_7323,N_7136);
nand U8179 (N_8179,N_6375,N_7188);
nor U8180 (N_8180,N_7134,N_7594);
nand U8181 (N_8181,N_7970,N_7893);
nand U8182 (N_8182,N_6697,N_7772);
nand U8183 (N_8183,N_6779,N_7121);
xor U8184 (N_8184,N_7308,N_7105);
nor U8185 (N_8185,N_6767,N_6606);
nand U8186 (N_8186,N_6698,N_6749);
or U8187 (N_8187,N_6735,N_6289);
nor U8188 (N_8188,N_7130,N_6674);
nor U8189 (N_8189,N_7742,N_6422);
or U8190 (N_8190,N_7220,N_6464);
nor U8191 (N_8191,N_6951,N_7842);
and U8192 (N_8192,N_6045,N_6122);
or U8193 (N_8193,N_6750,N_7137);
or U8194 (N_8194,N_6226,N_6341);
nor U8195 (N_8195,N_6473,N_7611);
nor U8196 (N_8196,N_7827,N_6100);
nand U8197 (N_8197,N_7927,N_7560);
nand U8198 (N_8198,N_7539,N_6262);
or U8199 (N_8199,N_6543,N_7152);
nor U8200 (N_8200,N_6769,N_7034);
or U8201 (N_8201,N_7217,N_7623);
nand U8202 (N_8202,N_7200,N_6723);
or U8203 (N_8203,N_7456,N_7898);
and U8204 (N_8204,N_6398,N_6149);
or U8205 (N_8205,N_7109,N_6327);
xor U8206 (N_8206,N_6903,N_7613);
nor U8207 (N_8207,N_6768,N_6102);
nor U8208 (N_8208,N_6290,N_6696);
xor U8209 (N_8209,N_7726,N_6208);
and U8210 (N_8210,N_6335,N_7865);
xor U8211 (N_8211,N_6737,N_7524);
nand U8212 (N_8212,N_7464,N_7910);
nand U8213 (N_8213,N_6718,N_7318);
and U8214 (N_8214,N_6949,N_7389);
and U8215 (N_8215,N_7060,N_6420);
nor U8216 (N_8216,N_7322,N_7744);
or U8217 (N_8217,N_6092,N_7087);
or U8218 (N_8218,N_6794,N_7093);
and U8219 (N_8219,N_7028,N_6198);
nor U8220 (N_8220,N_6472,N_6670);
nand U8221 (N_8221,N_6720,N_6228);
and U8222 (N_8222,N_7913,N_7753);
or U8223 (N_8223,N_7442,N_7097);
and U8224 (N_8224,N_7943,N_6677);
nand U8225 (N_8225,N_6030,N_7116);
and U8226 (N_8226,N_7936,N_6717);
or U8227 (N_8227,N_7044,N_6683);
xor U8228 (N_8228,N_6379,N_6583);
and U8229 (N_8229,N_6591,N_7472);
or U8230 (N_8230,N_7615,N_6594);
nor U8231 (N_8231,N_7293,N_6036);
nand U8232 (N_8232,N_7561,N_7720);
xnor U8233 (N_8233,N_7756,N_7259);
or U8234 (N_8234,N_6614,N_7740);
nand U8235 (N_8235,N_7287,N_6000);
and U8236 (N_8236,N_7931,N_7704);
nand U8237 (N_8237,N_7748,N_6605);
nor U8238 (N_8238,N_7864,N_6107);
nor U8239 (N_8239,N_7940,N_7845);
and U8240 (N_8240,N_7202,N_6653);
or U8241 (N_8241,N_6947,N_6663);
nor U8242 (N_8242,N_7733,N_6133);
and U8243 (N_8243,N_6932,N_7823);
xor U8244 (N_8244,N_7321,N_6104);
or U8245 (N_8245,N_7074,N_7590);
or U8246 (N_8246,N_6267,N_6394);
nand U8247 (N_8247,N_6017,N_6952);
nand U8248 (N_8248,N_7338,N_6865);
nor U8249 (N_8249,N_7967,N_6634);
nor U8250 (N_8250,N_6162,N_6343);
or U8251 (N_8251,N_6848,N_6626);
nor U8252 (N_8252,N_7606,N_6117);
nor U8253 (N_8253,N_7745,N_6551);
or U8254 (N_8254,N_6814,N_6144);
and U8255 (N_8255,N_6476,N_7754);
or U8256 (N_8256,N_7462,N_7738);
nor U8257 (N_8257,N_6480,N_6692);
nor U8258 (N_8258,N_6268,N_7495);
xnor U8259 (N_8259,N_7368,N_6139);
and U8260 (N_8260,N_7596,N_7268);
nand U8261 (N_8261,N_7730,N_6513);
and U8262 (N_8262,N_6595,N_7903);
or U8263 (N_8263,N_7616,N_7556);
nor U8264 (N_8264,N_7545,N_7270);
or U8265 (N_8265,N_7406,N_7148);
xnor U8266 (N_8266,N_6201,N_7454);
nand U8267 (N_8267,N_6108,N_7531);
or U8268 (N_8268,N_7231,N_6962);
nand U8269 (N_8269,N_6259,N_7373);
nand U8270 (N_8270,N_7269,N_6269);
nand U8271 (N_8271,N_6953,N_7546);
nand U8272 (N_8272,N_6592,N_6961);
nand U8273 (N_8273,N_7599,N_7530);
and U8274 (N_8274,N_7768,N_7876);
nor U8275 (N_8275,N_6186,N_7848);
nor U8276 (N_8276,N_6659,N_6093);
nor U8277 (N_8277,N_7708,N_6027);
nand U8278 (N_8278,N_6489,N_7991);
nor U8279 (N_8279,N_6646,N_6673);
nor U8280 (N_8280,N_7894,N_6552);
xnor U8281 (N_8281,N_7766,N_6509);
and U8282 (N_8282,N_6690,N_6866);
and U8283 (N_8283,N_6498,N_7146);
xor U8284 (N_8284,N_6300,N_7838);
nor U8285 (N_8285,N_6493,N_6417);
or U8286 (N_8286,N_6374,N_6699);
xnor U8287 (N_8287,N_6371,N_6544);
nor U8288 (N_8288,N_7379,N_6528);
or U8289 (N_8289,N_7216,N_6740);
and U8290 (N_8290,N_6998,N_7582);
xor U8291 (N_8291,N_6060,N_6011);
nand U8292 (N_8292,N_6832,N_7938);
and U8293 (N_8293,N_7209,N_6378);
xnor U8294 (N_8294,N_7573,N_6971);
xnor U8295 (N_8295,N_7887,N_6900);
nand U8296 (N_8296,N_6485,N_7071);
nand U8297 (N_8297,N_6119,N_7219);
nor U8298 (N_8298,N_7818,N_7836);
and U8299 (N_8299,N_7572,N_6403);
nand U8300 (N_8300,N_6427,N_6365);
nor U8301 (N_8301,N_7265,N_7163);
nor U8302 (N_8302,N_7584,N_7416);
nand U8303 (N_8303,N_7298,N_7629);
xnor U8304 (N_8304,N_7666,N_7895);
or U8305 (N_8305,N_7870,N_7349);
or U8306 (N_8306,N_6658,N_7179);
nor U8307 (N_8307,N_6063,N_6897);
or U8308 (N_8308,N_6418,N_7320);
xnor U8309 (N_8309,N_7850,N_6477);
and U8310 (N_8310,N_6725,N_6410);
nand U8311 (N_8311,N_6869,N_7998);
and U8312 (N_8312,N_6707,N_7884);
nor U8313 (N_8313,N_7315,N_7485);
xor U8314 (N_8314,N_7834,N_7739);
or U8315 (N_8315,N_6466,N_7500);
nand U8316 (N_8316,N_6972,N_6023);
and U8317 (N_8317,N_6068,N_7528);
xor U8318 (N_8318,N_7242,N_6545);
nor U8319 (N_8319,N_7684,N_6682);
nand U8320 (N_8320,N_7115,N_7691);
nor U8321 (N_8321,N_7354,N_6923);
nor U8322 (N_8322,N_6976,N_7961);
nor U8323 (N_8323,N_7412,N_6448);
nor U8324 (N_8324,N_7079,N_6457);
or U8325 (N_8325,N_7478,N_7329);
nor U8326 (N_8326,N_6954,N_7213);
nand U8327 (N_8327,N_7388,N_7548);
xnor U8328 (N_8328,N_6298,N_6497);
nor U8329 (N_8329,N_7133,N_6907);
nor U8330 (N_8330,N_6331,N_7990);
xnor U8331 (N_8331,N_6070,N_6950);
nand U8332 (N_8332,N_7453,N_6397);
and U8333 (N_8333,N_7062,N_7094);
nor U8334 (N_8334,N_6096,N_6412);
and U8335 (N_8335,N_7973,N_7731);
or U8336 (N_8336,N_6265,N_6282);
or U8337 (N_8337,N_6204,N_7396);
nand U8338 (N_8338,N_6478,N_7106);
nor U8339 (N_8339,N_7125,N_7111);
nor U8340 (N_8340,N_6729,N_7741);
nor U8341 (N_8341,N_7776,N_7477);
nor U8342 (N_8342,N_6055,N_7685);
and U8343 (N_8343,N_6560,N_7637);
nor U8344 (N_8344,N_7735,N_6854);
and U8345 (N_8345,N_7160,N_7247);
nand U8346 (N_8346,N_7331,N_6073);
or U8347 (N_8347,N_7775,N_7319);
nand U8348 (N_8348,N_6222,N_7429);
or U8349 (N_8349,N_6809,N_7668);
nand U8350 (N_8350,N_6536,N_7618);
nor U8351 (N_8351,N_6471,N_7662);
nand U8352 (N_8352,N_7372,N_7777);
nand U8353 (N_8353,N_6990,N_6181);
or U8354 (N_8354,N_6447,N_7496);
nand U8355 (N_8355,N_6392,N_7926);
xnor U8356 (N_8356,N_7088,N_6039);
nor U8357 (N_8357,N_6992,N_7814);
nor U8358 (N_8358,N_6839,N_7399);
or U8359 (N_8359,N_6571,N_7288);
nand U8360 (N_8360,N_6727,N_6981);
and U8361 (N_8361,N_6701,N_7067);
and U8362 (N_8362,N_7951,N_7035);
and U8363 (N_8363,N_6129,N_7709);
and U8364 (N_8364,N_6853,N_7614);
nor U8365 (N_8365,N_7245,N_7053);
or U8366 (N_8366,N_6213,N_7183);
nand U8367 (N_8367,N_7306,N_6484);
or U8368 (N_8368,N_7415,N_7409);
nand U8369 (N_8369,N_7494,N_7274);
or U8370 (N_8370,N_6714,N_7862);
or U8371 (N_8371,N_7169,N_6730);
and U8372 (N_8372,N_7295,N_6272);
nand U8373 (N_8373,N_7291,N_6456);
and U8374 (N_8374,N_7040,N_7559);
nand U8375 (N_8375,N_7460,N_7225);
nor U8376 (N_8376,N_7224,N_7583);
nand U8377 (N_8377,N_6496,N_7682);
nand U8378 (N_8378,N_7000,N_6243);
xor U8379 (N_8379,N_6632,N_6239);
nand U8380 (N_8380,N_6675,N_6373);
and U8381 (N_8381,N_7212,N_6655);
nor U8382 (N_8382,N_7487,N_7999);
and U8383 (N_8383,N_7486,N_6434);
and U8384 (N_8384,N_7339,N_6603);
and U8385 (N_8385,N_6199,N_6895);
or U8386 (N_8386,N_6851,N_7633);
or U8387 (N_8387,N_7811,N_7165);
and U8388 (N_8388,N_7064,N_6015);
nand U8389 (N_8389,N_6311,N_6522);
nand U8390 (N_8390,N_7313,N_6306);
nor U8391 (N_8391,N_7457,N_6431);
nor U8392 (N_8392,N_7591,N_7875);
and U8393 (N_8393,N_6049,N_6074);
or U8394 (N_8394,N_6285,N_6195);
nand U8395 (N_8395,N_7819,N_6323);
nand U8396 (N_8396,N_7982,N_7211);
or U8397 (N_8397,N_7853,N_7031);
and U8398 (N_8398,N_6487,N_7450);
nand U8399 (N_8399,N_7786,N_7005);
and U8400 (N_8400,N_6598,N_7840);
nor U8401 (N_8401,N_7930,N_6671);
nand U8402 (N_8402,N_7346,N_6926);
or U8403 (N_8403,N_7317,N_6034);
or U8404 (N_8404,N_7916,N_6633);
and U8405 (N_8405,N_6229,N_7170);
or U8406 (N_8406,N_6001,N_7248);
and U8407 (N_8407,N_7256,N_7505);
nand U8408 (N_8408,N_6890,N_7669);
nand U8409 (N_8409,N_7816,N_7059);
and U8410 (N_8410,N_7986,N_6731);
xor U8411 (N_8411,N_6021,N_7327);
or U8412 (N_8412,N_7027,N_7276);
and U8413 (N_8413,N_6676,N_6256);
nand U8414 (N_8414,N_7340,N_7538);
or U8415 (N_8415,N_6288,N_6106);
and U8416 (N_8416,N_6510,N_6530);
nand U8417 (N_8417,N_6419,N_7172);
or U8418 (N_8418,N_6296,N_7871);
nand U8419 (N_8419,N_6557,N_6816);
nand U8420 (N_8420,N_6918,N_6430);
nand U8421 (N_8421,N_7254,N_6077);
and U8422 (N_8422,N_7397,N_6338);
nand U8423 (N_8423,N_6123,N_7001);
nor U8424 (N_8424,N_6624,N_7490);
or U8425 (N_8425,N_6504,N_6879);
and U8426 (N_8426,N_7960,N_6798);
and U8427 (N_8427,N_7168,N_7223);
nor U8428 (N_8428,N_6389,N_6153);
nand U8429 (N_8429,N_7029,N_7634);
nand U8430 (N_8430,N_6183,N_7956);
nand U8431 (N_8431,N_7597,N_7952);
or U8432 (N_8432,N_6469,N_6121);
nor U8433 (N_8433,N_6511,N_6192);
or U8434 (N_8434,N_7182,N_7810);
nor U8435 (N_8435,N_6082,N_6402);
nand U8436 (N_8436,N_6930,N_6479);
nand U8437 (N_8437,N_7083,N_6079);
or U8438 (N_8438,N_6884,N_7418);
and U8439 (N_8439,N_6381,N_6597);
nor U8440 (N_8440,N_6746,N_6463);
nand U8441 (N_8441,N_7414,N_6680);
and U8442 (N_8442,N_7003,N_7844);
xor U8443 (N_8443,N_7728,N_6040);
nand U8444 (N_8444,N_6163,N_7997);
and U8445 (N_8445,N_6007,N_7362);
nor U8446 (N_8446,N_7863,N_7184);
nand U8447 (N_8447,N_7724,N_7607);
nand U8448 (N_8448,N_6116,N_6344);
and U8449 (N_8449,N_7965,N_6763);
or U8450 (N_8450,N_6414,N_6157);
or U8451 (N_8451,N_6333,N_7833);
and U8452 (N_8452,N_6554,N_7085);
or U8453 (N_8453,N_6709,N_6347);
or U8454 (N_8454,N_6946,N_6859);
nand U8455 (N_8455,N_6205,N_6126);
or U8456 (N_8456,N_6631,N_6396);
nor U8457 (N_8457,N_7156,N_6589);
and U8458 (N_8458,N_7714,N_6881);
or U8459 (N_8459,N_6086,N_6960);
nand U8460 (N_8460,N_7365,N_6191);
nand U8461 (N_8461,N_7806,N_7065);
nand U8462 (N_8462,N_6339,N_7830);
and U8463 (N_8463,N_7963,N_7086);
nor U8464 (N_8464,N_7360,N_6621);
xor U8465 (N_8465,N_7050,N_7906);
and U8466 (N_8466,N_7335,N_6309);
nor U8467 (N_8467,N_6388,N_6732);
nand U8468 (N_8468,N_7303,N_7007);
nand U8469 (N_8469,N_6733,N_6812);
nand U8470 (N_8470,N_7824,N_7802);
and U8471 (N_8471,N_6973,N_7729);
nor U8472 (N_8472,N_6649,N_7417);
and U8473 (N_8473,N_6250,N_7448);
or U8474 (N_8474,N_7297,N_7512);
and U8475 (N_8475,N_7603,N_6840);
and U8476 (N_8476,N_6906,N_7764);
xnor U8477 (N_8477,N_6297,N_6428);
nand U8478 (N_8478,N_7826,N_7888);
nor U8479 (N_8479,N_7879,N_7181);
and U8480 (N_8480,N_7037,N_7283);
xnor U8481 (N_8481,N_6570,N_7474);
nand U8482 (N_8482,N_6098,N_7459);
or U8483 (N_8483,N_7124,N_7872);
nand U8484 (N_8484,N_6505,N_7068);
nor U8485 (N_8485,N_6776,N_6569);
nand U8486 (N_8486,N_7446,N_7855);
or U8487 (N_8487,N_7859,N_6087);
or U8488 (N_8488,N_6974,N_7984);
or U8489 (N_8489,N_6363,N_7278);
nor U8490 (N_8490,N_7886,N_7762);
or U8491 (N_8491,N_7314,N_6637);
nor U8492 (N_8492,N_7195,N_6957);
nor U8493 (N_8493,N_7574,N_6722);
nor U8494 (N_8494,N_7994,N_7655);
or U8495 (N_8495,N_6650,N_6617);
and U8496 (N_8496,N_7192,N_7765);
and U8497 (N_8497,N_6042,N_7054);
and U8498 (N_8498,N_6177,N_7852);
nand U8499 (N_8499,N_6628,N_6449);
or U8500 (N_8500,N_6712,N_6206);
xor U8501 (N_8501,N_7366,N_7868);
nand U8502 (N_8502,N_6662,N_6071);
and U8503 (N_8503,N_7954,N_7550);
and U8504 (N_8504,N_7511,N_7800);
or U8505 (N_8505,N_6488,N_7403);
and U8506 (N_8506,N_6211,N_6980);
nor U8507 (N_8507,N_6541,N_7791);
nand U8508 (N_8508,N_7780,N_6894);
or U8509 (N_8509,N_6736,N_7344);
nand U8510 (N_8510,N_6384,N_6576);
and U8511 (N_8511,N_6189,N_6416);
nor U8512 (N_8512,N_6494,N_6529);
nand U8513 (N_8513,N_6977,N_6304);
nand U8514 (N_8514,N_6870,N_6280);
nor U8515 (N_8515,N_7917,N_6486);
nand U8516 (N_8516,N_7392,N_6877);
or U8517 (N_8517,N_7324,N_6958);
nand U8518 (N_8518,N_6041,N_7939);
nor U8519 (N_8519,N_7921,N_6235);
nand U8520 (N_8520,N_7056,N_6066);
xnor U8521 (N_8521,N_6058,N_6578);
and U8522 (N_8522,N_7126,N_7413);
nor U8523 (N_8523,N_6169,N_7568);
xor U8524 (N_8524,N_6274,N_7012);
or U8525 (N_8525,N_7395,N_6945);
nand U8526 (N_8526,N_7914,N_7521);
nor U8527 (N_8527,N_7718,N_7869);
nand U8528 (N_8528,N_6567,N_7626);
or U8529 (N_8529,N_7817,N_6801);
or U8530 (N_8530,N_6004,N_7030);
nor U8531 (N_8531,N_6630,N_6987);
nor U8532 (N_8532,N_6700,N_6715);
nor U8533 (N_8533,N_6467,N_6666);
nand U8534 (N_8534,N_7667,N_7411);
nor U8535 (N_8535,N_7197,N_7380);
nor U8536 (N_8536,N_6785,N_6979);
or U8537 (N_8537,N_7102,N_6721);
and U8538 (N_8538,N_6824,N_6013);
xnor U8539 (N_8539,N_6563,N_7281);
or U8540 (N_8540,N_7799,N_6783);
and U8541 (N_8541,N_7972,N_6889);
nor U8542 (N_8542,N_6546,N_6790);
or U8543 (N_8543,N_6534,N_6165);
and U8544 (N_8544,N_7905,N_6207);
or U8545 (N_8545,N_6756,N_6138);
and U8546 (N_8546,N_7282,N_6849);
and U8547 (N_8547,N_7267,N_7123);
nor U8548 (N_8548,N_7193,N_7650);
and U8549 (N_8549,N_6967,N_7347);
and U8550 (N_8550,N_7767,N_6622);
or U8551 (N_8551,N_6858,N_7937);
nor U8552 (N_8552,N_7540,N_7977);
nor U8553 (N_8553,N_7974,N_6002);
nor U8554 (N_8554,N_7419,N_7257);
and U8555 (N_8555,N_7790,N_6899);
and U8556 (N_8556,N_6353,N_7385);
nor U8557 (N_8557,N_7543,N_7141);
and U8558 (N_8558,N_7230,N_7356);
and U8559 (N_8559,N_6739,N_7746);
xor U8560 (N_8560,N_6588,N_6704);
and U8561 (N_8561,N_7069,N_7899);
or U8562 (N_8562,N_7378,N_6413);
or U8563 (N_8563,N_7432,N_6242);
nor U8564 (N_8564,N_7253,N_7801);
or U8565 (N_8565,N_7569,N_7567);
or U8566 (N_8566,N_6641,N_7769);
or U8567 (N_8567,N_7966,N_7911);
xor U8568 (N_8568,N_7214,N_6257);
and U8569 (N_8569,N_6385,N_7510);
nand U8570 (N_8570,N_7233,N_7727);
nand U8571 (N_8571,N_7407,N_6292);
or U8572 (N_8572,N_7514,N_6164);
xnor U8573 (N_8573,N_6796,N_7820);
xnor U8574 (N_8574,N_7600,N_6179);
or U8575 (N_8575,N_6273,N_6346);
nand U8576 (N_8576,N_6053,N_7479);
and U8577 (N_8577,N_6455,N_6532);
nand U8578 (N_8578,N_6253,N_7877);
or U8579 (N_8579,N_7964,N_6155);
and U8580 (N_8580,N_6661,N_7110);
xnor U8581 (N_8581,N_7553,N_6806);
nor U8582 (N_8582,N_6782,N_6887);
nor U8583 (N_8583,N_7676,N_6223);
nand U8584 (N_8584,N_7675,N_7578);
or U8585 (N_8585,N_6623,N_7628);
and U8586 (N_8586,N_7631,N_6094);
or U8587 (N_8587,N_7499,N_7919);
nor U8588 (N_8588,N_7326,N_7294);
nand U8589 (N_8589,N_6237,N_6161);
and U8590 (N_8590,N_7444,N_6792);
nor U8591 (N_8591,N_6533,N_6135);
nand U8592 (N_8592,N_6743,N_7155);
nand U8593 (N_8593,N_7458,N_6220);
nor U8594 (N_8594,N_6937,N_7713);
nor U8595 (N_8595,N_7683,N_6318);
and U8596 (N_8596,N_7143,N_7686);
or U8597 (N_8597,N_6643,N_6635);
nand U8598 (N_8598,N_6753,N_6482);
and U8599 (N_8599,N_7285,N_6009);
or U8600 (N_8600,N_7542,N_6616);
xor U8601 (N_8601,N_7882,N_6856);
and U8602 (N_8602,N_7046,N_6829);
and U8603 (N_8603,N_7250,N_7440);
nand U8604 (N_8604,N_6127,N_7503);
nand U8605 (N_8605,N_7529,N_7400);
or U8606 (N_8606,N_7784,N_7517);
nand U8607 (N_8607,N_7532,N_7175);
nand U8608 (N_8608,N_6787,N_7861);
nand U8609 (N_8609,N_6465,N_6831);
nor U8610 (N_8610,N_6627,N_6905);
nand U8611 (N_8611,N_7277,N_7364);
nand U8612 (N_8612,N_6047,N_7229);
nand U8613 (N_8613,N_6726,N_7405);
xnor U8614 (N_8614,N_6647,N_6584);
or U8615 (N_8615,N_6742,N_7052);
nor U8616 (N_8616,N_7646,N_6638);
nor U8617 (N_8617,N_7837,N_6453);
nand U8618 (N_8618,N_7760,N_7203);
xor U8619 (N_8619,N_7422,N_6249);
xnor U8620 (N_8620,N_7497,N_7638);
and U8621 (N_8621,N_7374,N_6372);
and U8622 (N_8622,N_6876,N_6811);
and U8623 (N_8623,N_6037,N_6325);
nor U8624 (N_8624,N_7867,N_7509);
or U8625 (N_8625,N_6305,N_6411);
xnor U8626 (N_8626,N_7920,N_7665);
or U8627 (N_8627,N_7463,N_6395);
xnor U8628 (N_8628,N_6350,N_6454);
and U8629 (N_8629,N_6245,N_6864);
nor U8630 (N_8630,N_6956,N_6523);
and U8631 (N_8631,N_6857,N_6996);
xnor U8632 (N_8632,N_6793,N_7151);
nor U8633 (N_8633,N_7880,N_7190);
nand U8634 (N_8634,N_7342,N_6216);
nor U8635 (N_8635,N_6270,N_7796);
nor U8636 (N_8636,N_6713,N_6908);
and U8637 (N_8637,N_7436,N_6025);
nor U8638 (N_8638,N_6120,N_6293);
nand U8639 (N_8639,N_7092,N_6029);
and U8640 (N_8640,N_6170,N_6766);
nand U8641 (N_8641,N_6582,N_6224);
or U8642 (N_8642,N_7073,N_7289);
xor U8643 (N_8643,N_7098,N_6777);
nand U8644 (N_8644,N_7377,N_7846);
nor U8645 (N_8645,N_7246,N_7725);
or U8646 (N_8646,N_7632,N_6143);
or U8647 (N_8647,N_7541,N_6159);
or U8648 (N_8648,N_7260,N_7258);
nor U8649 (N_8649,N_7466,N_6942);
nand U8650 (N_8650,N_6818,N_7443);
nand U8651 (N_8651,N_6264,N_7167);
nand U8652 (N_8652,N_6251,N_7286);
xor U8653 (N_8653,N_7674,N_7924);
or U8654 (N_8654,N_7264,N_7483);
nand U8655 (N_8655,N_7653,N_7832);
nor U8656 (N_8656,N_6440,N_6391);
xor U8657 (N_8657,N_7187,N_6834);
nor U8658 (N_8658,N_6757,N_6019);
and U8659 (N_8659,N_6515,N_6745);
and U8660 (N_8660,N_7770,N_6210);
and U8661 (N_8661,N_6444,N_6130);
and U8662 (N_8662,N_6874,N_7992);
nand U8663 (N_8663,N_6836,N_6620);
nand U8664 (N_8664,N_7563,N_7302);
nand U8665 (N_8665,N_6681,N_7839);
and U8666 (N_8666,N_6929,N_7129);
and U8667 (N_8667,N_7352,N_6401);
nand U8668 (N_8668,N_7431,N_7797);
nand U8669 (N_8669,N_6468,N_6033);
and U8670 (N_8670,N_6408,N_6227);
and U8671 (N_8671,N_6277,N_6795);
nor U8672 (N_8672,N_7475,N_6354);
nor U8673 (N_8673,N_6863,N_6283);
nand U8674 (N_8674,N_7334,N_6741);
and U8675 (N_8675,N_6760,N_7602);
nand U8676 (N_8676,N_7657,N_6994);
or U8677 (N_8677,N_7237,N_7159);
and U8678 (N_8678,N_6307,N_6636);
or U8679 (N_8679,N_7325,N_7210);
and U8680 (N_8680,N_6804,N_7369);
nand U8681 (N_8681,N_6565,N_7673);
nor U8682 (N_8682,N_7570,N_6691);
nor U8683 (N_8683,N_6105,N_7077);
and U8684 (N_8684,N_6520,N_7763);
and U8685 (N_8685,N_6573,N_6236);
nand U8686 (N_8686,N_7985,N_7687);
and U8687 (N_8687,N_6807,N_6648);
or U8688 (N_8688,N_7166,N_6321);
and U8689 (N_8689,N_7849,N_7610);
or U8690 (N_8690,N_7644,N_7547);
or U8691 (N_8691,N_6771,N_7113);
nand U8692 (N_8692,N_6791,N_6861);
xnor U8693 (N_8693,N_7015,N_6639);
nor U8694 (N_8694,N_6539,N_7150);
and U8695 (N_8695,N_7807,N_7423);
nor U8696 (N_8696,N_6922,N_6991);
or U8697 (N_8697,N_6252,N_7723);
or U8698 (N_8698,N_7923,N_7328);
nand U8699 (N_8699,N_6376,N_7371);
and U8700 (N_8700,N_7147,N_7017);
and U8701 (N_8701,N_7434,N_6668);
xor U8702 (N_8702,N_7468,N_7139);
or U8703 (N_8703,N_7480,N_7789);
nand U8704 (N_8704,N_6590,N_6762);
or U8705 (N_8705,N_7803,N_6828);
nor U8706 (N_8706,N_7484,N_7081);
nor U8707 (N_8707,N_7177,N_6140);
or U8708 (N_8708,N_7473,N_7145);
nor U8709 (N_8709,N_7945,N_6424);
nand U8710 (N_8710,N_7091,N_6514);
or U8711 (N_8711,N_7099,N_7892);
nor U8712 (N_8712,N_6238,N_7275);
or U8713 (N_8713,N_7272,N_7831);
xor U8714 (N_8714,N_6178,N_7698);
or U8715 (N_8715,N_6014,N_7185);
nand U8716 (N_8716,N_6429,N_7671);
xor U8717 (N_8717,N_6368,N_7394);
nand U8718 (N_8718,N_7447,N_6706);
xnor U8719 (N_8719,N_6362,N_6313);
and U8720 (N_8720,N_7828,N_7873);
or U8721 (N_8721,N_7912,N_7461);
nor U8722 (N_8722,N_7660,N_6400);
nor U8723 (N_8723,N_6048,N_6759);
and U8724 (N_8724,N_7009,N_7643);
or U8725 (N_8725,N_6131,N_6640);
or U8726 (N_8726,N_7424,N_6218);
xor U8727 (N_8727,N_6559,N_7847);
nor U8728 (N_8728,N_6483,N_6340);
or U8729 (N_8729,N_7240,N_6271);
nor U8730 (N_8730,N_6435,N_7502);
nor U8731 (N_8731,N_6970,N_7941);
or U8732 (N_8732,N_7717,N_7878);
and U8733 (N_8733,N_6158,N_6330);
nor U8734 (N_8734,N_6518,N_7451);
nor U8735 (N_8735,N_7142,N_7228);
nor U8736 (N_8736,N_7345,N_7971);
nand U8737 (N_8737,N_7605,N_7309);
xnor U8738 (N_8738,N_7575,N_6531);
nand U8739 (N_8739,N_6012,N_7640);
nand U8740 (N_8740,N_7617,N_7096);
xor U8741 (N_8741,N_7696,N_7587);
nor U8742 (N_8742,N_6336,N_7144);
nor U8743 (N_8743,N_6010,N_6651);
xnor U8744 (N_8744,N_7507,N_7057);
and U8745 (N_8745,N_6500,N_7523);
nor U8746 (N_8746,N_7891,N_6088);
and U8747 (N_8747,N_7962,N_6820);
nand U8748 (N_8748,N_6176,N_6708);
nor U8749 (N_8749,N_6035,N_6084);
or U8750 (N_8750,N_6826,N_7043);
and U8751 (N_8751,N_7773,N_6451);
nand U8752 (N_8752,N_6989,N_7290);
and U8753 (N_8753,N_7697,N_6425);
nand U8754 (N_8754,N_6685,N_6642);
or U8755 (N_8755,N_7858,N_7249);
and U8756 (N_8756,N_6910,N_7552);
nand U8757 (N_8757,N_6575,N_6695);
xnor U8758 (N_8758,N_6044,N_7885);
or U8759 (N_8759,N_6061,N_6279);
nand U8760 (N_8760,N_7622,N_6303);
xnor U8761 (N_8761,N_6822,N_6043);
or U8762 (N_8762,N_6247,N_7678);
and U8763 (N_8763,N_6568,N_7589);
or U8764 (N_8764,N_7465,N_7218);
and U8765 (N_8765,N_7922,N_7117);
or U8766 (N_8766,N_6160,N_7608);
nor U8767 (N_8767,N_7189,N_6941);
and U8768 (N_8768,N_7100,N_7648);
or U8769 (N_8769,N_6083,N_6442);
nand U8770 (N_8770,N_7311,N_6898);
nor U8771 (N_8771,N_6261,N_6988);
and U8772 (N_8772,N_7627,N_6450);
nand U8773 (N_8773,N_6909,N_7375);
nor U8774 (N_8774,N_7048,N_6805);
and U8775 (N_8775,N_7482,N_7204);
and U8776 (N_8776,N_7639,N_6615);
nand U8777 (N_8777,N_6825,N_7722);
or U8778 (N_8778,N_7620,N_6194);
nor U8779 (N_8779,N_6097,N_6610);
or U8780 (N_8780,N_7215,N_6540);
nand U8781 (N_8781,N_7390,N_7795);
or U8782 (N_8782,N_6490,N_6524);
xnor U8783 (N_8783,N_7794,N_7131);
or U8784 (N_8784,N_7101,N_7680);
nand U8785 (N_8785,N_6020,N_7164);
nor U8786 (N_8786,N_6003,N_7355);
and U8787 (N_8787,N_6775,N_7856);
and U8788 (N_8788,N_6837,N_6054);
nor U8789 (N_8789,N_7656,N_7761);
nand U8790 (N_8790,N_7262,N_7571);
and U8791 (N_8791,N_7205,N_6933);
and U8792 (N_8792,N_7948,N_7565);
nand U8793 (N_8793,N_6934,N_6187);
xor U8794 (N_8794,N_7707,N_6438);
or U8795 (N_8795,N_7402,N_7785);
nand U8796 (N_8796,N_6873,N_6550);
and U8797 (N_8797,N_6069,N_7783);
or U8798 (N_8798,N_7357,N_7929);
xor U8799 (N_8799,N_6702,N_7330);
or U8800 (N_8800,N_7425,N_7467);
or U8801 (N_8801,N_7066,N_6137);
and U8802 (N_8802,N_6248,N_6291);
nand U8803 (N_8803,N_7968,N_6050);
or U8804 (N_8804,N_7715,N_6625);
nand U8805 (N_8805,N_6491,N_7221);
or U8806 (N_8806,N_7750,N_6882);
and U8807 (N_8807,N_7798,N_7537);
or U8808 (N_8808,N_6038,N_6499);
or U8809 (N_8809,N_7243,N_6984);
and U8810 (N_8810,N_6888,N_7981);
or U8811 (N_8811,N_6689,N_6234);
xor U8812 (N_8812,N_6474,N_6203);
nand U8813 (N_8813,N_6780,N_6145);
and U8814 (N_8814,N_7897,N_6315);
nor U8815 (N_8815,N_7013,N_6146);
and U8816 (N_8816,N_7078,N_6441);
nand U8817 (N_8817,N_7975,N_7987);
nand U8818 (N_8818,N_6764,N_7021);
nand U8819 (N_8819,N_7006,N_7381);
and U8820 (N_8820,N_6517,N_7821);
nor U8821 (N_8821,N_7359,N_7703);
nand U8822 (N_8822,N_6948,N_6852);
and U8823 (N_8823,N_6738,N_7519);
nand U8824 (N_8824,N_7980,N_7804);
or U8825 (N_8825,N_7493,N_7367);
xnor U8826 (N_8826,N_7688,N_6558);
or U8827 (N_8827,N_6599,N_6461);
or U8828 (N_8828,N_7808,N_6399);
nor U8829 (N_8829,N_6969,N_7525);
nor U8830 (N_8830,N_6433,N_6184);
or U8831 (N_8831,N_6062,N_6549);
nor U8832 (N_8832,N_6393,N_7989);
nor U8833 (N_8833,N_6600,N_6911);
nor U8834 (N_8834,N_6101,N_6886);
and U8835 (N_8835,N_6287,N_6629);
nand U8836 (N_8836,N_6052,N_6521);
and U8837 (N_8837,N_6405,N_7909);
or U8838 (N_8838,N_6525,N_7393);
nor U8839 (N_8839,N_7566,N_6150);
and U8840 (N_8840,N_7551,N_6572);
and U8841 (N_8841,N_7601,N_7635);
or U8842 (N_8842,N_6190,N_6885);
nand U8843 (N_8843,N_7196,N_6562);
nor U8844 (N_8844,N_7679,N_7908);
and U8845 (N_8845,N_6175,N_7114);
or U8846 (N_8846,N_6197,N_6018);
nand U8847 (N_8847,N_6387,N_6022);
nor U8848 (N_8848,N_6871,N_7558);
and U8849 (N_8849,N_7925,N_6026);
or U8850 (N_8850,N_7441,N_7504);
or U8851 (N_8851,N_7812,N_7299);
or U8852 (N_8852,N_6611,N_6136);
or U8853 (N_8853,N_6361,N_7781);
nor U8854 (N_8854,N_6656,N_6512);
and U8855 (N_8855,N_6095,N_6752);
or U8856 (N_8856,N_6841,N_6358);
and U8857 (N_8857,N_7935,N_7793);
nand U8858 (N_8858,N_7508,N_7822);
or U8859 (N_8859,N_7969,N_6660);
nor U8860 (N_8860,N_7408,N_6278);
or U8861 (N_8861,N_6188,N_7934);
and U8862 (N_8862,N_7384,N_7854);
and U8863 (N_8863,N_7199,N_6679);
nor U8864 (N_8864,N_7835,N_6437);
nand U8865 (N_8865,N_6111,N_6326);
and U8866 (N_8866,N_7518,N_6917);
and U8867 (N_8867,N_6688,N_7351);
nand U8868 (N_8868,N_7238,N_6217);
and U8869 (N_8869,N_7119,N_7946);
and U8870 (N_8870,N_7586,N_7692);
and U8871 (N_8871,N_7070,N_6317);
nor U8872 (N_8872,N_7536,N_7206);
or U8873 (N_8873,N_6553,N_6548);
and U8874 (N_8874,N_6110,N_7410);
and U8875 (N_8875,N_6999,N_6436);
or U8876 (N_8876,N_6687,N_7455);
and U8877 (N_8877,N_7333,N_7194);
and U8878 (N_8878,N_6943,N_6423);
nor U8879 (N_8879,N_7792,N_7176);
or U8880 (N_8880,N_7949,N_7736);
nor U8881 (N_8881,N_6115,N_6645);
or U8882 (N_8882,N_6128,N_6915);
or U8883 (N_8883,N_6619,N_6604);
xnor U8884 (N_8884,N_6221,N_7058);
nand U8885 (N_8885,N_7522,N_7787);
nand U8886 (N_8886,N_6938,N_7004);
nand U8887 (N_8887,N_6406,N_7942);
xor U8888 (N_8888,N_7716,N_6329);
nand U8889 (N_8889,N_6747,N_7149);
nor U8890 (N_8890,N_6813,N_6744);
nor U8891 (N_8891,N_6607,N_6609);
or U8892 (N_8892,N_6193,N_6409);
nor U8893 (N_8893,N_7025,N_6896);
nand U8894 (N_8894,N_6470,N_7782);
or U8895 (N_8895,N_6665,N_7022);
nand U8896 (N_8896,N_7469,N_6585);
nor U8897 (N_8897,N_6940,N_6535);
and U8898 (N_8898,N_7016,N_6556);
or U8899 (N_8899,N_7815,N_7173);
or U8900 (N_8900,N_6901,N_7860);
nand U8901 (N_8901,N_7036,N_6348);
nor U8902 (N_8902,N_7118,N_6370);
xor U8903 (N_8903,N_6803,N_7279);
or U8904 (N_8904,N_7933,N_7681);
and U8905 (N_8905,N_6596,N_6064);
nand U8906 (N_8906,N_6921,N_7890);
nor U8907 (N_8907,N_6142,N_6352);
nor U8908 (N_8908,N_7593,N_6808);
or U8909 (N_8909,N_7430,N_7234);
nor U8910 (N_8910,N_6357,N_7564);
nand U8911 (N_8911,N_7024,N_7771);
and U8912 (N_8912,N_6240,N_7310);
and U8913 (N_8913,N_7515,N_6919);
or U8914 (N_8914,N_6847,N_7435);
and U8915 (N_8915,N_6555,N_6916);
nand U8916 (N_8916,N_7630,N_7953);
nand U8917 (N_8917,N_6593,N_6788);
nor U8918 (N_8918,N_7896,N_6345);
or U8919 (N_8919,N_7316,N_6728);
or U8920 (N_8920,N_6174,N_6075);
or U8921 (N_8921,N_6986,N_7759);
or U8922 (N_8922,N_6360,N_7645);
nor U8923 (N_8923,N_6924,N_6351);
and U8924 (N_8924,N_6867,N_6773);
and U8925 (N_8925,N_7993,N_7932);
and U8926 (N_8926,N_6612,N_7082);
xor U8927 (N_8927,N_6580,N_7498);
or U8928 (N_8928,N_7437,N_6295);
nand U8929 (N_8929,N_7336,N_6664);
and U8930 (N_8930,N_6686,N_6452);
nand U8931 (N_8931,N_7918,N_6359);
and U8932 (N_8932,N_7020,N_6993);
nand U8933 (N_8933,N_7239,N_6538);
xnor U8934 (N_8934,N_6966,N_6383);
or U8935 (N_8935,N_6778,N_7579);
nor U8936 (N_8936,N_7439,N_6233);
nand U8937 (N_8937,N_7127,N_7049);
and U8938 (N_8938,N_6459,N_6693);
nor U8939 (N_8939,N_6862,N_6356);
nor U8940 (N_8940,N_6893,N_7305);
xnor U8941 (N_8941,N_7978,N_6141);
nand U8942 (N_8942,N_6258,N_7711);
nand U8943 (N_8943,N_7549,N_6613);
and U8944 (N_8944,N_6678,N_7813);
nand U8945 (N_8945,N_7019,N_7690);
nand U8946 (N_8946,N_6579,N_7900);
nand U8947 (N_8947,N_6439,N_6850);
or U8948 (N_8948,N_6928,N_7619);
nor U8949 (N_8949,N_6892,N_6065);
and U8950 (N_8950,N_6800,N_7104);
nor U8951 (N_8951,N_6166,N_7235);
nor U8952 (N_8952,N_7625,N_7562);
and U8953 (N_8953,N_6975,N_7585);
or U8954 (N_8954,N_7719,N_7904);
or U8955 (N_8955,N_6024,N_6527);
nor U8956 (N_8956,N_6872,N_6936);
and U8957 (N_8957,N_7651,N_6076);
nor U8958 (N_8958,N_6072,N_6016);
nor U8959 (N_8959,N_7471,N_7489);
nand U8960 (N_8960,N_7095,N_7090);
nand U8961 (N_8961,N_7370,N_6180);
and U8962 (N_8962,N_7788,N_7232);
nor U8963 (N_8963,N_6944,N_7752);
and U8964 (N_8964,N_7312,N_7445);
xor U8965 (N_8965,N_6322,N_6566);
or U8966 (N_8966,N_6810,N_6080);
nand U8967 (N_8967,N_6758,N_7702);
nand U8968 (N_8968,N_7023,N_6618);
nor U8969 (N_8969,N_6939,N_7520);
nand U8970 (N_8970,N_7135,N_7554);
xor U8971 (N_8971,N_7588,N_6684);
nand U8972 (N_8972,N_7304,N_7178);
and U8973 (N_8973,N_6542,N_7076);
nand U8974 (N_8974,N_7103,N_7008);
or U8975 (N_8975,N_7701,N_6931);
and U8976 (N_8976,N_7712,N_6845);
xor U8977 (N_8977,N_7851,N_6342);
and U8978 (N_8978,N_7595,N_6334);
xor U8979 (N_8979,N_6955,N_7162);
or U8980 (N_8980,N_6547,N_6959);
nand U8981 (N_8981,N_6260,N_6827);
or U8982 (N_8982,N_7710,N_7527);
and U8983 (N_8983,N_6369,N_7198);
and U8984 (N_8984,N_7296,N_6772);
and U8985 (N_8985,N_6817,N_7592);
nand U8986 (N_8986,N_7778,N_7427);
or U8987 (N_8987,N_6843,N_6821);
nand U8988 (N_8988,N_7743,N_6125);
nor U8989 (N_8989,N_6784,N_6366);
nand U8990 (N_8990,N_7747,N_6789);
and U8991 (N_8991,N_6912,N_7652);
or U8992 (N_8992,N_6078,N_6667);
nor U8993 (N_8993,N_7516,N_7663);
nor U8994 (N_8994,N_7266,N_7749);
nor U8995 (N_8995,N_7157,N_6099);
nand U8996 (N_8996,N_6734,N_6883);
nor U8997 (N_8997,N_7883,N_7382);
and U8998 (N_8998,N_6390,N_7404);
nand U8999 (N_8999,N_6118,N_6046);
or U9000 (N_9000,N_6456,N_6620);
or U9001 (N_9001,N_6553,N_7766);
or U9002 (N_9002,N_7758,N_6755);
and U9003 (N_9003,N_7890,N_7872);
and U9004 (N_9004,N_6272,N_7566);
and U9005 (N_9005,N_6292,N_6928);
nand U9006 (N_9006,N_6256,N_6890);
xor U9007 (N_9007,N_7727,N_6333);
and U9008 (N_9008,N_6634,N_6891);
nand U9009 (N_9009,N_6729,N_7265);
xor U9010 (N_9010,N_7738,N_7605);
nor U9011 (N_9011,N_7931,N_7428);
or U9012 (N_9012,N_6233,N_6068);
or U9013 (N_9013,N_6779,N_6542);
nand U9014 (N_9014,N_6322,N_7125);
or U9015 (N_9015,N_6795,N_6049);
and U9016 (N_9016,N_7118,N_6484);
nor U9017 (N_9017,N_6705,N_6981);
and U9018 (N_9018,N_7175,N_6860);
xnor U9019 (N_9019,N_7567,N_6215);
nand U9020 (N_9020,N_6845,N_7300);
or U9021 (N_9021,N_7852,N_7099);
and U9022 (N_9022,N_7395,N_6530);
and U9023 (N_9023,N_6766,N_6588);
nand U9024 (N_9024,N_6581,N_7637);
nand U9025 (N_9025,N_6142,N_6888);
and U9026 (N_9026,N_6590,N_6799);
and U9027 (N_9027,N_6370,N_7680);
or U9028 (N_9028,N_7381,N_7823);
and U9029 (N_9029,N_6560,N_6021);
and U9030 (N_9030,N_7458,N_6587);
or U9031 (N_9031,N_6780,N_7295);
and U9032 (N_9032,N_6417,N_6247);
nand U9033 (N_9033,N_7372,N_7138);
or U9034 (N_9034,N_7723,N_7516);
nor U9035 (N_9035,N_7885,N_6884);
and U9036 (N_9036,N_6786,N_7256);
and U9037 (N_9037,N_7696,N_7277);
nor U9038 (N_9038,N_7818,N_6747);
xor U9039 (N_9039,N_7553,N_7369);
and U9040 (N_9040,N_7049,N_7530);
and U9041 (N_9041,N_6723,N_7140);
nand U9042 (N_9042,N_6153,N_7680);
and U9043 (N_9043,N_7573,N_6106);
nor U9044 (N_9044,N_7494,N_6317);
or U9045 (N_9045,N_7015,N_7342);
and U9046 (N_9046,N_6410,N_7242);
and U9047 (N_9047,N_6451,N_7661);
or U9048 (N_9048,N_6439,N_6646);
nand U9049 (N_9049,N_6356,N_7073);
nand U9050 (N_9050,N_6645,N_6303);
nand U9051 (N_9051,N_6033,N_6221);
and U9052 (N_9052,N_7099,N_7084);
and U9053 (N_9053,N_7347,N_6128);
or U9054 (N_9054,N_6104,N_7353);
nand U9055 (N_9055,N_7843,N_7191);
nor U9056 (N_9056,N_6610,N_6797);
or U9057 (N_9057,N_6498,N_6036);
xor U9058 (N_9058,N_7865,N_6987);
nand U9059 (N_9059,N_7941,N_7226);
nand U9060 (N_9060,N_6493,N_6216);
and U9061 (N_9061,N_7878,N_7341);
xor U9062 (N_9062,N_6797,N_7867);
or U9063 (N_9063,N_6752,N_6136);
or U9064 (N_9064,N_7995,N_6576);
nand U9065 (N_9065,N_7700,N_6852);
or U9066 (N_9066,N_7577,N_6153);
nor U9067 (N_9067,N_6345,N_7291);
nor U9068 (N_9068,N_7766,N_7026);
nor U9069 (N_9069,N_6075,N_6853);
or U9070 (N_9070,N_6275,N_6352);
or U9071 (N_9071,N_6768,N_7320);
nand U9072 (N_9072,N_7490,N_7248);
nand U9073 (N_9073,N_7358,N_7629);
nor U9074 (N_9074,N_6529,N_7258);
nor U9075 (N_9075,N_7126,N_7403);
xnor U9076 (N_9076,N_7315,N_7711);
xnor U9077 (N_9077,N_7283,N_6953);
nand U9078 (N_9078,N_7217,N_7057);
nand U9079 (N_9079,N_6048,N_6631);
or U9080 (N_9080,N_7432,N_6478);
and U9081 (N_9081,N_6336,N_6037);
xor U9082 (N_9082,N_7571,N_7037);
and U9083 (N_9083,N_6970,N_7419);
or U9084 (N_9084,N_7913,N_6334);
and U9085 (N_9085,N_7594,N_6768);
nor U9086 (N_9086,N_6971,N_6997);
and U9087 (N_9087,N_6244,N_7751);
nand U9088 (N_9088,N_7773,N_6885);
xor U9089 (N_9089,N_7736,N_7155);
or U9090 (N_9090,N_6140,N_7490);
nor U9091 (N_9091,N_6116,N_6680);
or U9092 (N_9092,N_7279,N_7818);
nand U9093 (N_9093,N_7035,N_6430);
xor U9094 (N_9094,N_7012,N_6286);
or U9095 (N_9095,N_6520,N_7648);
nor U9096 (N_9096,N_6969,N_7318);
nor U9097 (N_9097,N_7271,N_6048);
nor U9098 (N_9098,N_6533,N_7913);
nand U9099 (N_9099,N_7459,N_7761);
and U9100 (N_9100,N_6314,N_6904);
nor U9101 (N_9101,N_7965,N_6581);
nor U9102 (N_9102,N_7691,N_6988);
nor U9103 (N_9103,N_7201,N_7725);
nand U9104 (N_9104,N_6833,N_7345);
or U9105 (N_9105,N_6334,N_6166);
and U9106 (N_9106,N_7477,N_6952);
and U9107 (N_9107,N_6043,N_6794);
and U9108 (N_9108,N_6705,N_6038);
nand U9109 (N_9109,N_6795,N_6093);
nor U9110 (N_9110,N_6769,N_7283);
nand U9111 (N_9111,N_7168,N_7258);
xnor U9112 (N_9112,N_6400,N_6623);
or U9113 (N_9113,N_6216,N_7607);
and U9114 (N_9114,N_7544,N_7485);
nor U9115 (N_9115,N_7328,N_6404);
xor U9116 (N_9116,N_6843,N_7939);
and U9117 (N_9117,N_6396,N_6603);
nor U9118 (N_9118,N_7883,N_7332);
nand U9119 (N_9119,N_7090,N_6539);
nor U9120 (N_9120,N_7143,N_6378);
or U9121 (N_9121,N_6572,N_7344);
nand U9122 (N_9122,N_7892,N_6464);
and U9123 (N_9123,N_7944,N_7688);
xnor U9124 (N_9124,N_6762,N_7080);
or U9125 (N_9125,N_6034,N_7653);
nand U9126 (N_9126,N_7587,N_7074);
nor U9127 (N_9127,N_7606,N_6704);
nand U9128 (N_9128,N_7817,N_7798);
or U9129 (N_9129,N_7625,N_6890);
xnor U9130 (N_9130,N_6344,N_7969);
and U9131 (N_9131,N_7557,N_7802);
and U9132 (N_9132,N_6444,N_6963);
nor U9133 (N_9133,N_7493,N_6705);
nand U9134 (N_9134,N_7426,N_7550);
or U9135 (N_9135,N_7824,N_6330);
and U9136 (N_9136,N_6957,N_6380);
or U9137 (N_9137,N_6989,N_6904);
nor U9138 (N_9138,N_6489,N_7675);
or U9139 (N_9139,N_6464,N_7138);
nand U9140 (N_9140,N_6192,N_6942);
nor U9141 (N_9141,N_7013,N_7140);
xnor U9142 (N_9142,N_7701,N_7741);
and U9143 (N_9143,N_7137,N_7381);
nor U9144 (N_9144,N_7884,N_6443);
nand U9145 (N_9145,N_7645,N_6527);
nor U9146 (N_9146,N_7766,N_6309);
and U9147 (N_9147,N_6140,N_6749);
or U9148 (N_9148,N_6085,N_6140);
nor U9149 (N_9149,N_6101,N_7870);
and U9150 (N_9150,N_7363,N_6635);
nand U9151 (N_9151,N_7203,N_7116);
and U9152 (N_9152,N_7958,N_7032);
and U9153 (N_9153,N_7807,N_7651);
and U9154 (N_9154,N_6936,N_7848);
nor U9155 (N_9155,N_6801,N_6355);
nand U9156 (N_9156,N_6286,N_6848);
nor U9157 (N_9157,N_6555,N_7615);
nor U9158 (N_9158,N_7827,N_7207);
nand U9159 (N_9159,N_6662,N_6455);
or U9160 (N_9160,N_6592,N_6373);
or U9161 (N_9161,N_7643,N_6709);
nand U9162 (N_9162,N_6202,N_6155);
and U9163 (N_9163,N_7347,N_7966);
nand U9164 (N_9164,N_7179,N_7409);
or U9165 (N_9165,N_6280,N_6059);
nand U9166 (N_9166,N_6340,N_6649);
xnor U9167 (N_9167,N_6836,N_7069);
nor U9168 (N_9168,N_7194,N_7744);
or U9169 (N_9169,N_6548,N_6781);
nor U9170 (N_9170,N_7139,N_7639);
nor U9171 (N_9171,N_6089,N_7171);
nand U9172 (N_9172,N_6682,N_6099);
xor U9173 (N_9173,N_6804,N_6225);
xor U9174 (N_9174,N_6661,N_6676);
nor U9175 (N_9175,N_6994,N_6223);
nand U9176 (N_9176,N_7644,N_7269);
or U9177 (N_9177,N_7212,N_7069);
or U9178 (N_9178,N_6539,N_6152);
and U9179 (N_9179,N_6707,N_7599);
nand U9180 (N_9180,N_7395,N_6721);
and U9181 (N_9181,N_7722,N_7401);
and U9182 (N_9182,N_6490,N_7593);
nand U9183 (N_9183,N_7756,N_6940);
or U9184 (N_9184,N_6034,N_6851);
nand U9185 (N_9185,N_7212,N_7594);
xnor U9186 (N_9186,N_7053,N_7305);
nand U9187 (N_9187,N_7389,N_7025);
nor U9188 (N_9188,N_6792,N_6471);
or U9189 (N_9189,N_6669,N_6616);
nand U9190 (N_9190,N_6214,N_7797);
nor U9191 (N_9191,N_7230,N_6714);
xnor U9192 (N_9192,N_7973,N_7460);
and U9193 (N_9193,N_7072,N_6000);
xor U9194 (N_9194,N_7232,N_7492);
or U9195 (N_9195,N_6601,N_7344);
nand U9196 (N_9196,N_7360,N_6703);
xnor U9197 (N_9197,N_6579,N_7798);
and U9198 (N_9198,N_7126,N_7534);
or U9199 (N_9199,N_7029,N_6302);
nor U9200 (N_9200,N_7424,N_7946);
or U9201 (N_9201,N_6292,N_7072);
nand U9202 (N_9202,N_7864,N_6329);
nor U9203 (N_9203,N_6259,N_6347);
or U9204 (N_9204,N_7833,N_7744);
nor U9205 (N_9205,N_7637,N_7130);
nand U9206 (N_9206,N_6918,N_6082);
nand U9207 (N_9207,N_6337,N_6715);
and U9208 (N_9208,N_7456,N_6368);
and U9209 (N_9209,N_6982,N_7201);
and U9210 (N_9210,N_6224,N_6965);
and U9211 (N_9211,N_6777,N_7022);
nand U9212 (N_9212,N_7787,N_6950);
nand U9213 (N_9213,N_7604,N_6835);
nor U9214 (N_9214,N_6689,N_7681);
or U9215 (N_9215,N_7784,N_6866);
nor U9216 (N_9216,N_6048,N_7652);
and U9217 (N_9217,N_7193,N_6766);
and U9218 (N_9218,N_7279,N_7951);
xor U9219 (N_9219,N_7529,N_7967);
or U9220 (N_9220,N_7477,N_7410);
and U9221 (N_9221,N_7138,N_7839);
and U9222 (N_9222,N_7509,N_6332);
or U9223 (N_9223,N_6279,N_6803);
xor U9224 (N_9224,N_6985,N_6637);
or U9225 (N_9225,N_7338,N_6738);
xnor U9226 (N_9226,N_6095,N_6151);
nand U9227 (N_9227,N_7303,N_6592);
or U9228 (N_9228,N_7201,N_6639);
nor U9229 (N_9229,N_7422,N_6460);
nor U9230 (N_9230,N_6129,N_6758);
nand U9231 (N_9231,N_6198,N_7151);
or U9232 (N_9232,N_6622,N_7712);
nor U9233 (N_9233,N_6605,N_6191);
nand U9234 (N_9234,N_6747,N_6830);
nor U9235 (N_9235,N_6799,N_6562);
nand U9236 (N_9236,N_6837,N_7598);
nor U9237 (N_9237,N_7040,N_7239);
xnor U9238 (N_9238,N_7614,N_7317);
nand U9239 (N_9239,N_6045,N_6490);
or U9240 (N_9240,N_6251,N_7856);
nor U9241 (N_9241,N_6123,N_6056);
and U9242 (N_9242,N_7022,N_7141);
nand U9243 (N_9243,N_7399,N_6467);
nor U9244 (N_9244,N_6728,N_7494);
or U9245 (N_9245,N_7395,N_7697);
and U9246 (N_9246,N_7573,N_7694);
nor U9247 (N_9247,N_7483,N_6279);
or U9248 (N_9248,N_7422,N_7857);
or U9249 (N_9249,N_6034,N_6318);
and U9250 (N_9250,N_7915,N_6092);
xnor U9251 (N_9251,N_6741,N_7350);
nor U9252 (N_9252,N_7097,N_7982);
nor U9253 (N_9253,N_6689,N_6282);
or U9254 (N_9254,N_7762,N_7463);
nand U9255 (N_9255,N_6112,N_7134);
xor U9256 (N_9256,N_7734,N_6436);
and U9257 (N_9257,N_7766,N_6854);
nand U9258 (N_9258,N_6883,N_6814);
xnor U9259 (N_9259,N_7314,N_6928);
nor U9260 (N_9260,N_6700,N_7263);
xnor U9261 (N_9261,N_6819,N_7141);
and U9262 (N_9262,N_7575,N_6879);
and U9263 (N_9263,N_7555,N_7918);
nand U9264 (N_9264,N_6208,N_6211);
nor U9265 (N_9265,N_7128,N_7515);
nor U9266 (N_9266,N_6273,N_7640);
xnor U9267 (N_9267,N_7433,N_6253);
xor U9268 (N_9268,N_7488,N_7257);
xor U9269 (N_9269,N_7714,N_7744);
nand U9270 (N_9270,N_7054,N_7210);
or U9271 (N_9271,N_7005,N_7863);
nand U9272 (N_9272,N_7965,N_7314);
nand U9273 (N_9273,N_6488,N_6548);
nor U9274 (N_9274,N_6289,N_6500);
and U9275 (N_9275,N_7607,N_6463);
xor U9276 (N_9276,N_7741,N_7412);
or U9277 (N_9277,N_7783,N_7735);
or U9278 (N_9278,N_6316,N_7992);
or U9279 (N_9279,N_7238,N_6764);
xnor U9280 (N_9280,N_7489,N_6917);
nor U9281 (N_9281,N_7724,N_6640);
nor U9282 (N_9282,N_6248,N_6988);
nor U9283 (N_9283,N_7898,N_6332);
xor U9284 (N_9284,N_6655,N_6193);
and U9285 (N_9285,N_7808,N_6688);
and U9286 (N_9286,N_7863,N_6399);
and U9287 (N_9287,N_6748,N_7766);
xor U9288 (N_9288,N_7452,N_7186);
or U9289 (N_9289,N_6968,N_7171);
or U9290 (N_9290,N_7494,N_7858);
nor U9291 (N_9291,N_7762,N_6532);
or U9292 (N_9292,N_6597,N_6188);
or U9293 (N_9293,N_6797,N_7229);
or U9294 (N_9294,N_7049,N_7567);
or U9295 (N_9295,N_7273,N_7474);
nand U9296 (N_9296,N_6885,N_6878);
nor U9297 (N_9297,N_6572,N_6154);
and U9298 (N_9298,N_6615,N_6137);
nand U9299 (N_9299,N_7286,N_6562);
and U9300 (N_9300,N_7337,N_6862);
nand U9301 (N_9301,N_6662,N_7897);
nor U9302 (N_9302,N_6272,N_7084);
nor U9303 (N_9303,N_7389,N_6907);
nor U9304 (N_9304,N_7088,N_7618);
nor U9305 (N_9305,N_6491,N_6824);
and U9306 (N_9306,N_6037,N_7408);
nand U9307 (N_9307,N_7695,N_6767);
xor U9308 (N_9308,N_6066,N_7005);
or U9309 (N_9309,N_7923,N_7570);
nor U9310 (N_9310,N_6922,N_6499);
or U9311 (N_9311,N_6124,N_7297);
nand U9312 (N_9312,N_7872,N_6062);
or U9313 (N_9313,N_6029,N_7732);
nor U9314 (N_9314,N_7240,N_7834);
nor U9315 (N_9315,N_7170,N_7442);
nor U9316 (N_9316,N_6061,N_6149);
xor U9317 (N_9317,N_7678,N_6665);
or U9318 (N_9318,N_7843,N_6506);
and U9319 (N_9319,N_7190,N_7267);
xnor U9320 (N_9320,N_6934,N_7164);
or U9321 (N_9321,N_6056,N_7450);
nor U9322 (N_9322,N_6243,N_6849);
or U9323 (N_9323,N_6446,N_7981);
and U9324 (N_9324,N_6594,N_6302);
nand U9325 (N_9325,N_7806,N_6135);
or U9326 (N_9326,N_7184,N_7615);
and U9327 (N_9327,N_6012,N_6043);
nor U9328 (N_9328,N_6712,N_6979);
nand U9329 (N_9329,N_6159,N_7499);
nand U9330 (N_9330,N_7282,N_7103);
nor U9331 (N_9331,N_6596,N_6821);
and U9332 (N_9332,N_6574,N_6257);
nor U9333 (N_9333,N_7967,N_6106);
and U9334 (N_9334,N_6957,N_6148);
and U9335 (N_9335,N_7122,N_6318);
nor U9336 (N_9336,N_7678,N_6608);
or U9337 (N_9337,N_6131,N_7568);
and U9338 (N_9338,N_6960,N_6022);
or U9339 (N_9339,N_7454,N_6717);
xnor U9340 (N_9340,N_6758,N_7690);
and U9341 (N_9341,N_7533,N_6078);
nor U9342 (N_9342,N_7660,N_6022);
or U9343 (N_9343,N_7704,N_7006);
nand U9344 (N_9344,N_7906,N_6130);
nor U9345 (N_9345,N_7924,N_6369);
and U9346 (N_9346,N_7582,N_7089);
and U9347 (N_9347,N_6759,N_7051);
or U9348 (N_9348,N_7316,N_7199);
nor U9349 (N_9349,N_7259,N_6186);
or U9350 (N_9350,N_6629,N_6002);
and U9351 (N_9351,N_6229,N_6103);
or U9352 (N_9352,N_7554,N_7975);
and U9353 (N_9353,N_6897,N_6771);
and U9354 (N_9354,N_7132,N_7715);
nand U9355 (N_9355,N_7816,N_7518);
nor U9356 (N_9356,N_7838,N_7925);
nor U9357 (N_9357,N_6857,N_7320);
nand U9358 (N_9358,N_6477,N_6302);
xor U9359 (N_9359,N_6520,N_7874);
nor U9360 (N_9360,N_7112,N_7375);
nor U9361 (N_9361,N_7283,N_7553);
nand U9362 (N_9362,N_7077,N_6403);
xnor U9363 (N_9363,N_6273,N_6988);
xnor U9364 (N_9364,N_7150,N_6755);
and U9365 (N_9365,N_7834,N_6965);
nand U9366 (N_9366,N_6393,N_7335);
or U9367 (N_9367,N_7389,N_6232);
nand U9368 (N_9368,N_6708,N_7374);
or U9369 (N_9369,N_7615,N_6609);
and U9370 (N_9370,N_6312,N_7127);
and U9371 (N_9371,N_6234,N_7112);
or U9372 (N_9372,N_6615,N_6410);
or U9373 (N_9373,N_6773,N_6145);
and U9374 (N_9374,N_7240,N_7916);
or U9375 (N_9375,N_7083,N_7618);
or U9376 (N_9376,N_6671,N_6624);
xnor U9377 (N_9377,N_7341,N_6876);
and U9378 (N_9378,N_7109,N_6624);
or U9379 (N_9379,N_6133,N_6461);
nor U9380 (N_9380,N_7388,N_6767);
nand U9381 (N_9381,N_6233,N_7133);
xnor U9382 (N_9382,N_6162,N_7354);
nor U9383 (N_9383,N_7807,N_6670);
and U9384 (N_9384,N_7876,N_6461);
xor U9385 (N_9385,N_7191,N_7713);
nor U9386 (N_9386,N_7220,N_6270);
xnor U9387 (N_9387,N_7002,N_6398);
nand U9388 (N_9388,N_7364,N_6474);
or U9389 (N_9389,N_6930,N_7265);
or U9390 (N_9390,N_7451,N_7634);
and U9391 (N_9391,N_6556,N_6139);
xor U9392 (N_9392,N_7782,N_6820);
nor U9393 (N_9393,N_7848,N_6690);
or U9394 (N_9394,N_7620,N_7608);
or U9395 (N_9395,N_7147,N_6452);
xnor U9396 (N_9396,N_6823,N_7020);
or U9397 (N_9397,N_6928,N_6311);
nand U9398 (N_9398,N_6620,N_6194);
or U9399 (N_9399,N_6939,N_6483);
or U9400 (N_9400,N_6567,N_6393);
nor U9401 (N_9401,N_6284,N_6155);
xnor U9402 (N_9402,N_6211,N_7201);
nor U9403 (N_9403,N_6166,N_6877);
and U9404 (N_9404,N_6009,N_7464);
nand U9405 (N_9405,N_6919,N_7574);
nand U9406 (N_9406,N_6959,N_6740);
nor U9407 (N_9407,N_7470,N_6839);
xor U9408 (N_9408,N_6496,N_7243);
and U9409 (N_9409,N_7623,N_7340);
nand U9410 (N_9410,N_6552,N_7822);
nor U9411 (N_9411,N_6213,N_6302);
nand U9412 (N_9412,N_6851,N_7082);
xor U9413 (N_9413,N_6809,N_7006);
or U9414 (N_9414,N_7532,N_7525);
xnor U9415 (N_9415,N_7040,N_7466);
nand U9416 (N_9416,N_6532,N_6696);
or U9417 (N_9417,N_7670,N_7149);
and U9418 (N_9418,N_7024,N_6179);
nand U9419 (N_9419,N_7929,N_7199);
nor U9420 (N_9420,N_6077,N_6724);
or U9421 (N_9421,N_6260,N_7920);
xnor U9422 (N_9422,N_6101,N_7550);
or U9423 (N_9423,N_6587,N_6738);
and U9424 (N_9424,N_7461,N_7319);
or U9425 (N_9425,N_7185,N_6683);
or U9426 (N_9426,N_7612,N_6992);
or U9427 (N_9427,N_6993,N_6463);
nand U9428 (N_9428,N_6973,N_6035);
nor U9429 (N_9429,N_7401,N_6912);
xor U9430 (N_9430,N_6515,N_6757);
nand U9431 (N_9431,N_6524,N_6967);
or U9432 (N_9432,N_7207,N_7548);
nor U9433 (N_9433,N_6002,N_7290);
or U9434 (N_9434,N_7781,N_7774);
nand U9435 (N_9435,N_6969,N_6592);
nor U9436 (N_9436,N_7066,N_7394);
nor U9437 (N_9437,N_6651,N_7867);
or U9438 (N_9438,N_7480,N_7539);
and U9439 (N_9439,N_7609,N_7680);
nor U9440 (N_9440,N_6606,N_6320);
xnor U9441 (N_9441,N_7864,N_7776);
or U9442 (N_9442,N_6838,N_7138);
nand U9443 (N_9443,N_7294,N_7613);
xnor U9444 (N_9444,N_6137,N_6483);
nor U9445 (N_9445,N_6266,N_7025);
or U9446 (N_9446,N_7134,N_7021);
and U9447 (N_9447,N_7779,N_6189);
or U9448 (N_9448,N_6231,N_6732);
nor U9449 (N_9449,N_7676,N_7522);
or U9450 (N_9450,N_7842,N_7908);
nand U9451 (N_9451,N_6875,N_7068);
nand U9452 (N_9452,N_7714,N_6697);
xor U9453 (N_9453,N_7026,N_6400);
nand U9454 (N_9454,N_7805,N_6269);
or U9455 (N_9455,N_7479,N_6588);
and U9456 (N_9456,N_6282,N_7448);
nand U9457 (N_9457,N_7782,N_6233);
or U9458 (N_9458,N_7292,N_6246);
or U9459 (N_9459,N_7623,N_7726);
and U9460 (N_9460,N_6464,N_6193);
nor U9461 (N_9461,N_6616,N_7088);
and U9462 (N_9462,N_6321,N_7382);
or U9463 (N_9463,N_6225,N_7822);
and U9464 (N_9464,N_6826,N_6119);
nand U9465 (N_9465,N_7746,N_7089);
nor U9466 (N_9466,N_7017,N_6183);
and U9467 (N_9467,N_6466,N_6329);
and U9468 (N_9468,N_7497,N_7905);
nand U9469 (N_9469,N_6214,N_6676);
nor U9470 (N_9470,N_6880,N_6358);
nand U9471 (N_9471,N_6895,N_6885);
and U9472 (N_9472,N_6929,N_6074);
xnor U9473 (N_9473,N_7803,N_7381);
or U9474 (N_9474,N_6667,N_6844);
nor U9475 (N_9475,N_7465,N_7089);
nor U9476 (N_9476,N_7753,N_7774);
nand U9477 (N_9477,N_6175,N_7618);
nand U9478 (N_9478,N_6799,N_7493);
xor U9479 (N_9479,N_6707,N_6322);
nor U9480 (N_9480,N_6800,N_6243);
or U9481 (N_9481,N_7335,N_7158);
xnor U9482 (N_9482,N_6001,N_7245);
and U9483 (N_9483,N_6836,N_7170);
nor U9484 (N_9484,N_7746,N_6718);
nand U9485 (N_9485,N_6655,N_6519);
or U9486 (N_9486,N_7529,N_6889);
or U9487 (N_9487,N_6739,N_7043);
or U9488 (N_9488,N_7164,N_7743);
nand U9489 (N_9489,N_6928,N_7843);
or U9490 (N_9490,N_7173,N_6756);
and U9491 (N_9491,N_7296,N_6835);
and U9492 (N_9492,N_7482,N_7256);
nor U9493 (N_9493,N_6900,N_7141);
or U9494 (N_9494,N_7819,N_6993);
nor U9495 (N_9495,N_7631,N_6729);
nand U9496 (N_9496,N_6860,N_6210);
or U9497 (N_9497,N_6827,N_6837);
and U9498 (N_9498,N_6143,N_6389);
nand U9499 (N_9499,N_7387,N_7144);
nor U9500 (N_9500,N_7794,N_6041);
xnor U9501 (N_9501,N_7571,N_7620);
or U9502 (N_9502,N_6818,N_6831);
nor U9503 (N_9503,N_6446,N_6406);
nand U9504 (N_9504,N_7081,N_7200);
and U9505 (N_9505,N_6710,N_7771);
or U9506 (N_9506,N_6008,N_7593);
nor U9507 (N_9507,N_7650,N_6278);
nor U9508 (N_9508,N_7160,N_6126);
or U9509 (N_9509,N_7779,N_7688);
or U9510 (N_9510,N_6406,N_7065);
nor U9511 (N_9511,N_6847,N_7748);
xnor U9512 (N_9512,N_7721,N_6876);
and U9513 (N_9513,N_6905,N_6271);
and U9514 (N_9514,N_6049,N_7739);
nor U9515 (N_9515,N_6666,N_6383);
or U9516 (N_9516,N_6463,N_7894);
nand U9517 (N_9517,N_7375,N_6892);
nor U9518 (N_9518,N_6866,N_7651);
and U9519 (N_9519,N_6688,N_7688);
or U9520 (N_9520,N_6247,N_6922);
or U9521 (N_9521,N_7263,N_6279);
or U9522 (N_9522,N_6778,N_6382);
nand U9523 (N_9523,N_6544,N_6116);
xor U9524 (N_9524,N_7454,N_7207);
nor U9525 (N_9525,N_7940,N_6987);
and U9526 (N_9526,N_6722,N_7080);
or U9527 (N_9527,N_6038,N_7004);
xor U9528 (N_9528,N_6993,N_6975);
and U9529 (N_9529,N_6341,N_6375);
nand U9530 (N_9530,N_6021,N_6352);
and U9531 (N_9531,N_7950,N_6353);
nand U9532 (N_9532,N_6768,N_7398);
and U9533 (N_9533,N_7637,N_6153);
nand U9534 (N_9534,N_7748,N_6002);
nor U9535 (N_9535,N_6148,N_6845);
nor U9536 (N_9536,N_6767,N_6216);
nor U9537 (N_9537,N_6754,N_6433);
nor U9538 (N_9538,N_6807,N_7829);
and U9539 (N_9539,N_7852,N_6566);
nand U9540 (N_9540,N_6371,N_7481);
or U9541 (N_9541,N_7960,N_6031);
and U9542 (N_9542,N_6434,N_6436);
or U9543 (N_9543,N_6722,N_6511);
and U9544 (N_9544,N_6978,N_7707);
or U9545 (N_9545,N_6376,N_6555);
and U9546 (N_9546,N_6179,N_7666);
nand U9547 (N_9547,N_7828,N_7154);
and U9548 (N_9548,N_7193,N_7544);
xor U9549 (N_9549,N_7433,N_6525);
nand U9550 (N_9550,N_7418,N_6137);
nor U9551 (N_9551,N_7454,N_6637);
and U9552 (N_9552,N_6131,N_7707);
nand U9553 (N_9553,N_7652,N_7039);
nor U9554 (N_9554,N_6892,N_6471);
and U9555 (N_9555,N_7490,N_6450);
nand U9556 (N_9556,N_7237,N_6507);
or U9557 (N_9557,N_7703,N_6174);
or U9558 (N_9558,N_6840,N_7305);
nor U9559 (N_9559,N_7901,N_6516);
nor U9560 (N_9560,N_6877,N_6517);
nand U9561 (N_9561,N_6998,N_7298);
xor U9562 (N_9562,N_6750,N_6299);
or U9563 (N_9563,N_6183,N_6339);
xnor U9564 (N_9564,N_7172,N_6086);
xnor U9565 (N_9565,N_7461,N_7915);
or U9566 (N_9566,N_6174,N_7132);
and U9567 (N_9567,N_7926,N_6263);
and U9568 (N_9568,N_7486,N_6226);
or U9569 (N_9569,N_7243,N_6229);
and U9570 (N_9570,N_6252,N_7820);
nand U9571 (N_9571,N_6214,N_7511);
nand U9572 (N_9572,N_7137,N_7354);
xor U9573 (N_9573,N_7116,N_6614);
xor U9574 (N_9574,N_6847,N_6298);
or U9575 (N_9575,N_6778,N_7747);
nor U9576 (N_9576,N_6378,N_6972);
and U9577 (N_9577,N_7904,N_6809);
nand U9578 (N_9578,N_6645,N_6182);
nor U9579 (N_9579,N_6555,N_7271);
nor U9580 (N_9580,N_7153,N_7636);
and U9581 (N_9581,N_7485,N_7887);
and U9582 (N_9582,N_6901,N_7920);
and U9583 (N_9583,N_7117,N_6492);
xor U9584 (N_9584,N_6270,N_6478);
xor U9585 (N_9585,N_7841,N_7562);
or U9586 (N_9586,N_6224,N_6899);
and U9587 (N_9587,N_7280,N_7694);
nand U9588 (N_9588,N_6192,N_7669);
and U9589 (N_9589,N_6256,N_7831);
nor U9590 (N_9590,N_6187,N_6021);
nand U9591 (N_9591,N_7247,N_7417);
xnor U9592 (N_9592,N_7342,N_6549);
nand U9593 (N_9593,N_6018,N_6354);
and U9594 (N_9594,N_6042,N_6475);
and U9595 (N_9595,N_7353,N_7154);
nand U9596 (N_9596,N_7109,N_6349);
or U9597 (N_9597,N_6975,N_7981);
nor U9598 (N_9598,N_7645,N_6037);
and U9599 (N_9599,N_7971,N_6180);
nand U9600 (N_9600,N_7576,N_6765);
nor U9601 (N_9601,N_6923,N_7755);
nor U9602 (N_9602,N_6667,N_7594);
xnor U9603 (N_9603,N_6762,N_7603);
or U9604 (N_9604,N_7668,N_7320);
xnor U9605 (N_9605,N_6408,N_6793);
and U9606 (N_9606,N_7445,N_7411);
and U9607 (N_9607,N_6552,N_7389);
nor U9608 (N_9608,N_7365,N_7703);
nor U9609 (N_9609,N_7365,N_6810);
and U9610 (N_9610,N_7467,N_7138);
nand U9611 (N_9611,N_6708,N_7399);
and U9612 (N_9612,N_7390,N_7448);
xor U9613 (N_9613,N_7471,N_6648);
nor U9614 (N_9614,N_7583,N_7143);
nor U9615 (N_9615,N_6456,N_7916);
nor U9616 (N_9616,N_6408,N_6310);
and U9617 (N_9617,N_6435,N_6548);
nor U9618 (N_9618,N_7061,N_6286);
nor U9619 (N_9619,N_6423,N_6575);
nor U9620 (N_9620,N_7400,N_7771);
and U9621 (N_9621,N_6407,N_7337);
nor U9622 (N_9622,N_6802,N_6707);
or U9623 (N_9623,N_7154,N_6127);
nor U9624 (N_9624,N_7869,N_7654);
nand U9625 (N_9625,N_7226,N_7537);
nand U9626 (N_9626,N_6211,N_6704);
xnor U9627 (N_9627,N_7341,N_7770);
and U9628 (N_9628,N_6579,N_6710);
or U9629 (N_9629,N_6321,N_7367);
or U9630 (N_9630,N_6167,N_6899);
nand U9631 (N_9631,N_6492,N_6785);
or U9632 (N_9632,N_7435,N_6399);
or U9633 (N_9633,N_7831,N_7325);
or U9634 (N_9634,N_6973,N_7124);
nand U9635 (N_9635,N_6208,N_7611);
or U9636 (N_9636,N_7680,N_7097);
and U9637 (N_9637,N_7047,N_6286);
and U9638 (N_9638,N_7656,N_6805);
nand U9639 (N_9639,N_7010,N_7563);
and U9640 (N_9640,N_7431,N_6963);
and U9641 (N_9641,N_6003,N_6010);
and U9642 (N_9642,N_7786,N_6940);
or U9643 (N_9643,N_6769,N_7981);
or U9644 (N_9644,N_6062,N_6235);
nor U9645 (N_9645,N_7472,N_7849);
xnor U9646 (N_9646,N_7864,N_6250);
nor U9647 (N_9647,N_6306,N_6029);
and U9648 (N_9648,N_7501,N_7566);
nand U9649 (N_9649,N_6293,N_7730);
and U9650 (N_9650,N_6133,N_7618);
and U9651 (N_9651,N_6195,N_6755);
or U9652 (N_9652,N_7209,N_7959);
and U9653 (N_9653,N_7565,N_6668);
or U9654 (N_9654,N_6807,N_6758);
or U9655 (N_9655,N_7083,N_6146);
and U9656 (N_9656,N_7760,N_7608);
xnor U9657 (N_9657,N_6507,N_6255);
nor U9658 (N_9658,N_7851,N_7493);
or U9659 (N_9659,N_6812,N_7557);
nand U9660 (N_9660,N_7371,N_6358);
or U9661 (N_9661,N_6974,N_7542);
and U9662 (N_9662,N_6910,N_6496);
nand U9663 (N_9663,N_7431,N_6006);
or U9664 (N_9664,N_6446,N_7903);
or U9665 (N_9665,N_6992,N_7178);
nor U9666 (N_9666,N_7787,N_6697);
or U9667 (N_9667,N_6436,N_6585);
nor U9668 (N_9668,N_7584,N_7455);
or U9669 (N_9669,N_7153,N_6377);
or U9670 (N_9670,N_7380,N_7389);
or U9671 (N_9671,N_6941,N_6925);
nor U9672 (N_9672,N_7497,N_7451);
or U9673 (N_9673,N_7866,N_6409);
nor U9674 (N_9674,N_6941,N_6531);
nand U9675 (N_9675,N_7698,N_6227);
nand U9676 (N_9676,N_6551,N_6529);
nor U9677 (N_9677,N_7587,N_6801);
nand U9678 (N_9678,N_6738,N_7673);
and U9679 (N_9679,N_6307,N_7142);
or U9680 (N_9680,N_7461,N_7292);
nor U9681 (N_9681,N_7262,N_6168);
xor U9682 (N_9682,N_6013,N_6968);
nor U9683 (N_9683,N_7122,N_7017);
nand U9684 (N_9684,N_6936,N_6648);
nor U9685 (N_9685,N_6978,N_6992);
nand U9686 (N_9686,N_7252,N_6883);
nand U9687 (N_9687,N_6411,N_6767);
and U9688 (N_9688,N_6624,N_6695);
xor U9689 (N_9689,N_6390,N_7170);
nand U9690 (N_9690,N_6667,N_7117);
or U9691 (N_9691,N_7826,N_6606);
or U9692 (N_9692,N_7896,N_7245);
nand U9693 (N_9693,N_6252,N_6848);
nand U9694 (N_9694,N_7394,N_7982);
or U9695 (N_9695,N_6374,N_6294);
nand U9696 (N_9696,N_7751,N_6708);
nand U9697 (N_9697,N_6259,N_7057);
xnor U9698 (N_9698,N_6609,N_6261);
nor U9699 (N_9699,N_7168,N_7113);
or U9700 (N_9700,N_6044,N_7189);
and U9701 (N_9701,N_6340,N_6164);
nor U9702 (N_9702,N_6217,N_6711);
xor U9703 (N_9703,N_6854,N_6976);
nand U9704 (N_9704,N_6663,N_6123);
xnor U9705 (N_9705,N_6564,N_7871);
or U9706 (N_9706,N_6929,N_6153);
or U9707 (N_9707,N_6601,N_7548);
and U9708 (N_9708,N_7765,N_6560);
nor U9709 (N_9709,N_6862,N_7246);
and U9710 (N_9710,N_7365,N_6368);
and U9711 (N_9711,N_7974,N_7719);
and U9712 (N_9712,N_7078,N_6123);
nor U9713 (N_9713,N_7353,N_7670);
nand U9714 (N_9714,N_6152,N_7565);
nor U9715 (N_9715,N_7101,N_7820);
xnor U9716 (N_9716,N_6992,N_6648);
nand U9717 (N_9717,N_7608,N_7698);
or U9718 (N_9718,N_6091,N_6049);
or U9719 (N_9719,N_7816,N_6212);
or U9720 (N_9720,N_6132,N_7953);
and U9721 (N_9721,N_7952,N_7427);
nand U9722 (N_9722,N_6235,N_7977);
xnor U9723 (N_9723,N_7339,N_6607);
nand U9724 (N_9724,N_7988,N_6841);
or U9725 (N_9725,N_6574,N_7184);
or U9726 (N_9726,N_7415,N_6089);
and U9727 (N_9727,N_7212,N_7094);
or U9728 (N_9728,N_7147,N_7238);
and U9729 (N_9729,N_7044,N_7284);
or U9730 (N_9730,N_7127,N_6737);
nor U9731 (N_9731,N_6191,N_7071);
or U9732 (N_9732,N_6423,N_6692);
nor U9733 (N_9733,N_6314,N_6739);
or U9734 (N_9734,N_6628,N_7634);
and U9735 (N_9735,N_6465,N_6477);
nand U9736 (N_9736,N_6915,N_7502);
and U9737 (N_9737,N_7746,N_6839);
nand U9738 (N_9738,N_7609,N_6035);
or U9739 (N_9739,N_6153,N_7956);
and U9740 (N_9740,N_6277,N_6261);
or U9741 (N_9741,N_6040,N_7962);
and U9742 (N_9742,N_6074,N_6693);
nand U9743 (N_9743,N_6606,N_6242);
and U9744 (N_9744,N_7448,N_7073);
and U9745 (N_9745,N_7615,N_6546);
and U9746 (N_9746,N_7294,N_6574);
and U9747 (N_9747,N_7894,N_6438);
and U9748 (N_9748,N_7024,N_6507);
xnor U9749 (N_9749,N_6072,N_6619);
xnor U9750 (N_9750,N_7350,N_7226);
nor U9751 (N_9751,N_7931,N_7294);
or U9752 (N_9752,N_6583,N_6553);
nor U9753 (N_9753,N_6121,N_7180);
nand U9754 (N_9754,N_7894,N_7820);
nor U9755 (N_9755,N_6848,N_7259);
nor U9756 (N_9756,N_6851,N_6450);
nor U9757 (N_9757,N_6444,N_7832);
nand U9758 (N_9758,N_6643,N_7690);
nor U9759 (N_9759,N_6198,N_7941);
nor U9760 (N_9760,N_7637,N_6327);
and U9761 (N_9761,N_6616,N_6958);
or U9762 (N_9762,N_7622,N_6092);
nand U9763 (N_9763,N_7460,N_7447);
or U9764 (N_9764,N_6086,N_6874);
and U9765 (N_9765,N_6204,N_6133);
nand U9766 (N_9766,N_6423,N_6147);
nand U9767 (N_9767,N_7300,N_7677);
or U9768 (N_9768,N_6687,N_7796);
or U9769 (N_9769,N_6371,N_7027);
xnor U9770 (N_9770,N_7599,N_7915);
or U9771 (N_9771,N_6033,N_7357);
or U9772 (N_9772,N_6414,N_6998);
and U9773 (N_9773,N_7450,N_7122);
xnor U9774 (N_9774,N_6825,N_7222);
nor U9775 (N_9775,N_6450,N_6033);
or U9776 (N_9776,N_7506,N_6576);
nor U9777 (N_9777,N_7757,N_6180);
and U9778 (N_9778,N_6178,N_7531);
nand U9779 (N_9779,N_7637,N_7767);
nand U9780 (N_9780,N_6128,N_7798);
nand U9781 (N_9781,N_7517,N_7450);
nand U9782 (N_9782,N_7900,N_7611);
nand U9783 (N_9783,N_7038,N_7288);
nor U9784 (N_9784,N_6549,N_6219);
nor U9785 (N_9785,N_6680,N_6878);
nand U9786 (N_9786,N_7159,N_7279);
nand U9787 (N_9787,N_7998,N_6308);
nand U9788 (N_9788,N_7671,N_6734);
nand U9789 (N_9789,N_7027,N_6287);
or U9790 (N_9790,N_6424,N_7690);
and U9791 (N_9791,N_6147,N_7236);
nand U9792 (N_9792,N_7033,N_6986);
nor U9793 (N_9793,N_6040,N_6545);
and U9794 (N_9794,N_7868,N_7421);
nand U9795 (N_9795,N_7039,N_7756);
and U9796 (N_9796,N_7795,N_7900);
nand U9797 (N_9797,N_6363,N_7726);
or U9798 (N_9798,N_7880,N_7426);
nor U9799 (N_9799,N_7900,N_6381);
or U9800 (N_9800,N_7955,N_6661);
or U9801 (N_9801,N_7690,N_6342);
and U9802 (N_9802,N_6045,N_6233);
nand U9803 (N_9803,N_7753,N_6802);
and U9804 (N_9804,N_7766,N_6118);
xnor U9805 (N_9805,N_6694,N_6883);
or U9806 (N_9806,N_6347,N_6003);
or U9807 (N_9807,N_7271,N_6642);
nand U9808 (N_9808,N_7408,N_6524);
xor U9809 (N_9809,N_6821,N_7513);
or U9810 (N_9810,N_7900,N_7729);
nor U9811 (N_9811,N_7365,N_7664);
and U9812 (N_9812,N_7789,N_7936);
nand U9813 (N_9813,N_7596,N_6607);
nor U9814 (N_9814,N_6262,N_7858);
xnor U9815 (N_9815,N_7905,N_7044);
nor U9816 (N_9816,N_7885,N_6068);
or U9817 (N_9817,N_7589,N_6880);
nand U9818 (N_9818,N_7031,N_6734);
xnor U9819 (N_9819,N_6578,N_7609);
nand U9820 (N_9820,N_6061,N_6701);
or U9821 (N_9821,N_6456,N_7963);
nand U9822 (N_9822,N_7010,N_7941);
or U9823 (N_9823,N_7080,N_7885);
nand U9824 (N_9824,N_7451,N_6488);
nand U9825 (N_9825,N_7208,N_6928);
xor U9826 (N_9826,N_6561,N_6547);
or U9827 (N_9827,N_7661,N_7383);
or U9828 (N_9828,N_6028,N_6358);
and U9829 (N_9829,N_7859,N_6060);
xor U9830 (N_9830,N_6257,N_7616);
and U9831 (N_9831,N_6351,N_7083);
nand U9832 (N_9832,N_6823,N_6738);
nor U9833 (N_9833,N_7255,N_6898);
nor U9834 (N_9834,N_6078,N_6874);
and U9835 (N_9835,N_6731,N_6151);
and U9836 (N_9836,N_6464,N_7413);
and U9837 (N_9837,N_7262,N_7597);
nand U9838 (N_9838,N_6013,N_7697);
or U9839 (N_9839,N_6623,N_6381);
nand U9840 (N_9840,N_6923,N_6259);
and U9841 (N_9841,N_6312,N_6117);
nor U9842 (N_9842,N_6980,N_6907);
nand U9843 (N_9843,N_6709,N_7182);
nor U9844 (N_9844,N_7545,N_7340);
nand U9845 (N_9845,N_7882,N_6170);
and U9846 (N_9846,N_6636,N_7681);
nor U9847 (N_9847,N_7823,N_6112);
or U9848 (N_9848,N_7732,N_7217);
xnor U9849 (N_9849,N_6847,N_7764);
or U9850 (N_9850,N_6825,N_7115);
xor U9851 (N_9851,N_6931,N_6569);
nand U9852 (N_9852,N_7605,N_6333);
or U9853 (N_9853,N_7251,N_6994);
nand U9854 (N_9854,N_6902,N_7190);
nor U9855 (N_9855,N_7760,N_6895);
or U9856 (N_9856,N_6438,N_6550);
or U9857 (N_9857,N_6119,N_7236);
nor U9858 (N_9858,N_7921,N_6495);
and U9859 (N_9859,N_6480,N_7506);
xor U9860 (N_9860,N_6734,N_6268);
or U9861 (N_9861,N_7806,N_6081);
nand U9862 (N_9862,N_7965,N_6713);
nor U9863 (N_9863,N_6179,N_7681);
or U9864 (N_9864,N_6668,N_6139);
xnor U9865 (N_9865,N_6588,N_7638);
or U9866 (N_9866,N_7879,N_6503);
nand U9867 (N_9867,N_6983,N_7822);
nand U9868 (N_9868,N_7238,N_7365);
nand U9869 (N_9869,N_6766,N_6799);
xnor U9870 (N_9870,N_6524,N_6371);
and U9871 (N_9871,N_6531,N_6097);
and U9872 (N_9872,N_7737,N_6596);
or U9873 (N_9873,N_7240,N_7670);
xor U9874 (N_9874,N_6304,N_6145);
nor U9875 (N_9875,N_7587,N_7677);
nor U9876 (N_9876,N_7523,N_7485);
nand U9877 (N_9877,N_6182,N_7441);
or U9878 (N_9878,N_7861,N_7745);
xnor U9879 (N_9879,N_6824,N_6757);
or U9880 (N_9880,N_7667,N_6233);
xnor U9881 (N_9881,N_7248,N_6016);
and U9882 (N_9882,N_7745,N_7836);
nor U9883 (N_9883,N_7038,N_6761);
or U9884 (N_9884,N_6839,N_7507);
nor U9885 (N_9885,N_7198,N_7931);
xor U9886 (N_9886,N_7491,N_6858);
and U9887 (N_9887,N_6598,N_7796);
and U9888 (N_9888,N_6195,N_7999);
nand U9889 (N_9889,N_6388,N_7392);
xnor U9890 (N_9890,N_6573,N_6882);
and U9891 (N_9891,N_7330,N_6481);
and U9892 (N_9892,N_7883,N_7321);
and U9893 (N_9893,N_6607,N_7468);
nand U9894 (N_9894,N_6719,N_6893);
or U9895 (N_9895,N_7451,N_6821);
nand U9896 (N_9896,N_6374,N_6908);
nor U9897 (N_9897,N_7550,N_7131);
or U9898 (N_9898,N_6084,N_6205);
or U9899 (N_9899,N_7606,N_6187);
xor U9900 (N_9900,N_7266,N_7599);
or U9901 (N_9901,N_6110,N_7130);
or U9902 (N_9902,N_7693,N_6741);
and U9903 (N_9903,N_6181,N_7522);
and U9904 (N_9904,N_7416,N_7127);
nand U9905 (N_9905,N_6286,N_7015);
nand U9906 (N_9906,N_6911,N_7399);
or U9907 (N_9907,N_6032,N_6801);
nor U9908 (N_9908,N_6347,N_7787);
nor U9909 (N_9909,N_7236,N_6697);
or U9910 (N_9910,N_7929,N_6588);
nand U9911 (N_9911,N_7086,N_7788);
and U9912 (N_9912,N_6798,N_6008);
nand U9913 (N_9913,N_7129,N_6854);
nor U9914 (N_9914,N_7280,N_7244);
or U9915 (N_9915,N_7234,N_6754);
nand U9916 (N_9916,N_7577,N_6660);
and U9917 (N_9917,N_7184,N_7017);
nand U9918 (N_9918,N_7133,N_6046);
nand U9919 (N_9919,N_6676,N_6680);
nand U9920 (N_9920,N_6702,N_6934);
xor U9921 (N_9921,N_7170,N_7763);
or U9922 (N_9922,N_7388,N_6496);
xnor U9923 (N_9923,N_6631,N_6255);
or U9924 (N_9924,N_6455,N_6133);
nor U9925 (N_9925,N_7792,N_7260);
nor U9926 (N_9926,N_6671,N_7174);
xor U9927 (N_9927,N_7162,N_6107);
or U9928 (N_9928,N_7768,N_6237);
nor U9929 (N_9929,N_7798,N_7505);
nand U9930 (N_9930,N_6849,N_6283);
nand U9931 (N_9931,N_6070,N_6701);
nand U9932 (N_9932,N_6013,N_7392);
or U9933 (N_9933,N_7145,N_7719);
nor U9934 (N_9934,N_6681,N_6258);
nand U9935 (N_9935,N_6302,N_7754);
nand U9936 (N_9936,N_7967,N_7002);
and U9937 (N_9937,N_6989,N_7401);
nand U9938 (N_9938,N_6873,N_6359);
nand U9939 (N_9939,N_7840,N_7770);
nand U9940 (N_9940,N_6087,N_7804);
or U9941 (N_9941,N_6337,N_7185);
and U9942 (N_9942,N_6421,N_7459);
and U9943 (N_9943,N_7650,N_7130);
xnor U9944 (N_9944,N_6691,N_7707);
nand U9945 (N_9945,N_6589,N_6723);
nand U9946 (N_9946,N_6990,N_7085);
and U9947 (N_9947,N_6051,N_7534);
and U9948 (N_9948,N_7739,N_6288);
nand U9949 (N_9949,N_7312,N_7288);
xor U9950 (N_9950,N_7122,N_7955);
xnor U9951 (N_9951,N_7273,N_7773);
nand U9952 (N_9952,N_6044,N_6659);
or U9953 (N_9953,N_7058,N_7876);
or U9954 (N_9954,N_6439,N_7431);
and U9955 (N_9955,N_7658,N_7265);
nor U9956 (N_9956,N_6935,N_6529);
and U9957 (N_9957,N_6950,N_7863);
xor U9958 (N_9958,N_6573,N_7831);
or U9959 (N_9959,N_7880,N_7571);
or U9960 (N_9960,N_7946,N_6407);
or U9961 (N_9961,N_7615,N_6632);
nand U9962 (N_9962,N_6018,N_6677);
or U9963 (N_9963,N_7329,N_6273);
nor U9964 (N_9964,N_6841,N_7651);
or U9965 (N_9965,N_7470,N_7776);
and U9966 (N_9966,N_7460,N_6481);
or U9967 (N_9967,N_6182,N_6987);
or U9968 (N_9968,N_6562,N_7047);
nor U9969 (N_9969,N_6782,N_7178);
nor U9970 (N_9970,N_7568,N_6145);
or U9971 (N_9971,N_6020,N_6860);
and U9972 (N_9972,N_7981,N_7060);
xnor U9973 (N_9973,N_6781,N_6986);
or U9974 (N_9974,N_7051,N_6166);
xnor U9975 (N_9975,N_7304,N_7537);
nor U9976 (N_9976,N_6769,N_6681);
or U9977 (N_9977,N_6469,N_7648);
xor U9978 (N_9978,N_7322,N_6725);
nand U9979 (N_9979,N_6849,N_7701);
nor U9980 (N_9980,N_6908,N_7485);
and U9981 (N_9981,N_7739,N_7107);
or U9982 (N_9982,N_7565,N_7810);
or U9983 (N_9983,N_6320,N_7979);
xnor U9984 (N_9984,N_7350,N_7200);
nand U9985 (N_9985,N_6916,N_6073);
xor U9986 (N_9986,N_7685,N_7018);
nor U9987 (N_9987,N_7621,N_7683);
nor U9988 (N_9988,N_6424,N_7952);
nor U9989 (N_9989,N_7280,N_6491);
or U9990 (N_9990,N_6761,N_6572);
xnor U9991 (N_9991,N_6379,N_7535);
nand U9992 (N_9992,N_7446,N_7960);
nand U9993 (N_9993,N_7717,N_6271);
nand U9994 (N_9994,N_6290,N_7567);
nand U9995 (N_9995,N_6065,N_6116);
nor U9996 (N_9996,N_6163,N_7497);
xnor U9997 (N_9997,N_6390,N_6363);
nand U9998 (N_9998,N_7685,N_7520);
xor U9999 (N_9999,N_7679,N_7191);
nand UO_0 (O_0,N_9429,N_8550);
nand UO_1 (O_1,N_8376,N_9671);
and UO_2 (O_2,N_9492,N_8829);
nor UO_3 (O_3,N_9768,N_8728);
and UO_4 (O_4,N_9423,N_9898);
or UO_5 (O_5,N_8016,N_8722);
nand UO_6 (O_6,N_8235,N_9915);
nand UO_7 (O_7,N_9640,N_8735);
or UO_8 (O_8,N_9719,N_9757);
nand UO_9 (O_9,N_8055,N_8684);
and UO_10 (O_10,N_9311,N_8551);
nand UO_11 (O_11,N_8600,N_9954);
nand UO_12 (O_12,N_9211,N_8514);
nand UO_13 (O_13,N_9329,N_8881);
and UO_14 (O_14,N_9636,N_8632);
nand UO_15 (O_15,N_9210,N_9814);
nor UO_16 (O_16,N_8814,N_8380);
xnor UO_17 (O_17,N_8003,N_9914);
and UO_18 (O_18,N_9341,N_9100);
nand UO_19 (O_19,N_8367,N_9616);
nand UO_20 (O_20,N_9782,N_8953);
and UO_21 (O_21,N_9012,N_9978);
or UO_22 (O_22,N_8199,N_8081);
nand UO_23 (O_23,N_8863,N_8145);
and UO_24 (O_24,N_8272,N_9183);
nand UO_25 (O_25,N_8714,N_8713);
nor UO_26 (O_26,N_8628,N_9314);
xnor UO_27 (O_27,N_8783,N_9910);
and UO_28 (O_28,N_9494,N_8737);
and UO_29 (O_29,N_8321,N_9824);
nor UO_30 (O_30,N_9245,N_9375);
or UO_31 (O_31,N_9922,N_9597);
nand UO_32 (O_32,N_9785,N_9904);
or UO_33 (O_33,N_8390,N_8398);
nand UO_34 (O_34,N_8712,N_9647);
nand UO_35 (O_35,N_8416,N_9909);
nand UO_36 (O_36,N_9927,N_9026);
or UO_37 (O_37,N_9382,N_9158);
xnor UO_38 (O_38,N_8257,N_8212);
nor UO_39 (O_39,N_8732,N_8138);
or UO_40 (O_40,N_9749,N_9422);
or UO_41 (O_41,N_9400,N_8511);
nor UO_42 (O_42,N_9637,N_9251);
and UO_43 (O_43,N_8271,N_8778);
and UO_44 (O_44,N_9555,N_9133);
or UO_45 (O_45,N_8149,N_9857);
and UO_46 (O_46,N_9434,N_8054);
nor UO_47 (O_47,N_8805,N_8729);
or UO_48 (O_48,N_8370,N_9651);
nand UO_49 (O_49,N_8912,N_8608);
xnor UO_50 (O_50,N_9846,N_9541);
or UO_51 (O_51,N_9103,N_8485);
or UO_52 (O_52,N_8520,N_8825);
and UO_53 (O_53,N_9425,N_9090);
nand UO_54 (O_54,N_9352,N_9034);
xnor UO_55 (O_55,N_9209,N_8685);
nand UO_56 (O_56,N_9713,N_8964);
nand UO_57 (O_57,N_8837,N_9143);
nor UO_58 (O_58,N_9615,N_9728);
or UO_59 (O_59,N_9379,N_8818);
nor UO_60 (O_60,N_9495,N_9943);
xnor UO_61 (O_61,N_8965,N_8372);
nand UO_62 (O_62,N_9661,N_9729);
xnor UO_63 (O_63,N_9124,N_9725);
and UO_64 (O_64,N_8404,N_8816);
and UO_65 (O_65,N_8426,N_9003);
nand UO_66 (O_66,N_8447,N_9854);
nor UO_67 (O_67,N_8413,N_9754);
nand UO_68 (O_68,N_8762,N_9006);
and UO_69 (O_69,N_8353,N_8446);
nand UO_70 (O_70,N_8696,N_8553);
or UO_71 (O_71,N_8549,N_8085);
and UO_72 (O_72,N_9081,N_9624);
and UO_73 (O_73,N_8217,N_9086);
nand UO_74 (O_74,N_8092,N_9182);
nor UO_75 (O_75,N_8640,N_8099);
nand UO_76 (O_76,N_9313,N_8113);
and UO_77 (O_77,N_8284,N_9044);
or UO_78 (O_78,N_8435,N_8342);
nand UO_79 (O_79,N_8229,N_9902);
nand UO_80 (O_80,N_8689,N_9256);
and UO_81 (O_81,N_9803,N_8038);
nand UO_82 (O_82,N_9703,N_8682);
or UO_83 (O_83,N_8823,N_8977);
or UO_84 (O_84,N_8868,N_9377);
nor UO_85 (O_85,N_9859,N_9482);
nand UO_86 (O_86,N_8898,N_8343);
nor UO_87 (O_87,N_9087,N_8754);
xnor UO_88 (O_88,N_9232,N_8817);
or UO_89 (O_89,N_8688,N_9459);
or UO_90 (O_90,N_9206,N_8335);
or UO_91 (O_91,N_9126,N_9589);
nand UO_92 (O_92,N_8704,N_9069);
nand UO_93 (O_93,N_8958,N_9746);
xnor UO_94 (O_94,N_9146,N_8176);
nor UO_95 (O_95,N_8623,N_9947);
and UO_96 (O_96,N_9498,N_8862);
nor UO_97 (O_97,N_8593,N_8503);
nand UO_98 (O_98,N_9769,N_8559);
nor UO_99 (O_99,N_9410,N_9856);
and UO_100 (O_100,N_8281,N_8811);
nand UO_101 (O_101,N_9617,N_9469);
or UO_102 (O_102,N_9140,N_8356);
and UO_103 (O_103,N_9448,N_8359);
or UO_104 (O_104,N_8207,N_9024);
nor UO_105 (O_105,N_8261,N_9796);
nand UO_106 (O_106,N_8674,N_9432);
and UO_107 (O_107,N_9505,N_9391);
xor UO_108 (O_108,N_9295,N_8601);
nor UO_109 (O_109,N_8761,N_9384);
nor UO_110 (O_110,N_8245,N_8961);
or UO_111 (O_111,N_9600,N_8455);
xor UO_112 (O_112,N_8901,N_8213);
nor UO_113 (O_113,N_9831,N_8334);
nor UO_114 (O_114,N_8889,N_9860);
or UO_115 (O_115,N_8570,N_9554);
xnor UO_116 (O_116,N_9243,N_8987);
nor UO_117 (O_117,N_9507,N_8209);
xnor UO_118 (O_118,N_8646,N_9581);
nor UO_119 (O_119,N_9586,N_9468);
xnor UO_120 (O_120,N_8107,N_9950);
nor UO_121 (O_121,N_8386,N_9663);
or UO_122 (O_122,N_9350,N_9395);
and UO_123 (O_123,N_8399,N_9948);
and UO_124 (O_124,N_8848,N_9317);
or UO_125 (O_125,N_8239,N_8440);
or UO_126 (O_126,N_9548,N_8385);
and UO_127 (O_127,N_9489,N_8530);
or UO_128 (O_128,N_9791,N_8153);
and UO_129 (O_129,N_9602,N_8341);
nor UO_130 (O_130,N_9771,N_8833);
or UO_131 (O_131,N_8289,N_9956);
and UO_132 (O_132,N_8915,N_8585);
or UO_133 (O_133,N_9825,N_9903);
nand UO_134 (O_134,N_9986,N_8957);
and UO_135 (O_135,N_9532,N_9763);
or UO_136 (O_136,N_9009,N_8716);
and UO_137 (O_137,N_8617,N_9918);
and UO_138 (O_138,N_8127,N_9237);
nand UO_139 (O_139,N_9940,N_8998);
and UO_140 (O_140,N_8676,N_8132);
nand UO_141 (O_141,N_9335,N_9573);
nor UO_142 (O_142,N_9453,N_9166);
nor UO_143 (O_143,N_8523,N_8673);
and UO_144 (O_144,N_9184,N_8088);
nor UO_145 (O_145,N_9307,N_9518);
nor UO_146 (O_146,N_9715,N_9439);
and UO_147 (O_147,N_9040,N_9582);
nand UO_148 (O_148,N_8610,N_9996);
and UO_149 (O_149,N_8846,N_8906);
nor UO_150 (O_150,N_9125,N_8799);
and UO_151 (O_151,N_8109,N_9113);
and UO_152 (O_152,N_8793,N_9116);
nand UO_153 (O_153,N_9850,N_9955);
nor UO_154 (O_154,N_9818,N_8950);
and UO_155 (O_155,N_9449,N_9576);
nand UO_156 (O_156,N_9369,N_8001);
and UO_157 (O_157,N_8519,N_9110);
nand UO_158 (O_158,N_8219,N_8744);
nor UO_159 (O_159,N_8711,N_9755);
nor UO_160 (O_160,N_9465,N_8798);
and UO_161 (O_161,N_9111,N_8467);
nand UO_162 (O_162,N_8120,N_8108);
or UO_163 (O_163,N_8642,N_8845);
and UO_164 (O_164,N_8963,N_8122);
nor UO_165 (O_165,N_8432,N_8715);
and UO_166 (O_166,N_8720,N_8922);
nand UO_167 (O_167,N_8489,N_9225);
or UO_168 (O_168,N_8202,N_9679);
or UO_169 (O_169,N_8659,N_9741);
nor UO_170 (O_170,N_9889,N_8899);
nor UO_171 (O_171,N_8086,N_9753);
and UO_172 (O_172,N_9957,N_8575);
nor UO_173 (O_173,N_9928,N_8832);
nand UO_174 (O_174,N_9406,N_8537);
and UO_175 (O_175,N_9745,N_9320);
nor UO_176 (O_176,N_9872,N_8885);
nor UO_177 (O_177,N_8100,N_8460);
and UO_178 (O_178,N_9387,N_8923);
or UO_179 (O_179,N_9230,N_8782);
or UO_180 (O_180,N_8547,N_9809);
or UO_181 (O_181,N_8792,N_9858);
nor UO_182 (O_182,N_8278,N_8206);
nand UO_183 (O_183,N_8952,N_8328);
nor UO_184 (O_184,N_9207,N_8017);
nor UO_185 (O_185,N_8116,N_9515);
nor UO_186 (O_186,N_8363,N_8044);
nor UO_187 (O_187,N_9490,N_9901);
xnor UO_188 (O_188,N_9523,N_8077);
nor UO_189 (O_189,N_9319,N_9897);
or UO_190 (O_190,N_8855,N_9007);
nor UO_191 (O_191,N_8415,N_9421);
nor UO_192 (O_192,N_8581,N_8701);
nand UO_193 (O_193,N_8766,N_9951);
and UO_194 (O_194,N_9936,N_8903);
nor UO_195 (O_195,N_9273,N_8591);
or UO_196 (O_196,N_8477,N_8238);
nor UO_197 (O_197,N_9804,N_9798);
nand UO_198 (O_198,N_9260,N_9051);
nor UO_199 (O_199,N_8373,N_8430);
and UO_200 (O_200,N_8663,N_9266);
nand UO_201 (O_201,N_8752,N_9974);
and UO_202 (O_202,N_8412,N_8204);
nand UO_203 (O_203,N_8164,N_8645);
nand UO_204 (O_204,N_8548,N_9175);
nand UO_205 (O_205,N_8369,N_8037);
and UO_206 (O_206,N_8558,N_8210);
xor UO_207 (O_207,N_8327,N_8853);
nand UO_208 (O_208,N_9851,N_9519);
and UO_209 (O_209,N_9185,N_9000);
and UO_210 (O_210,N_9281,N_9149);
nor UO_211 (O_211,N_9073,N_8170);
and UO_212 (O_212,N_8956,N_8536);
nor UO_213 (O_213,N_8280,N_9438);
and UO_214 (O_214,N_8118,N_8546);
nor UO_215 (O_215,N_8942,N_9134);
or UO_216 (O_216,N_8203,N_8764);
nand UO_217 (O_217,N_9873,N_8566);
and UO_218 (O_218,N_9466,N_9562);
and UO_219 (O_219,N_9911,N_9217);
or UO_220 (O_220,N_8142,N_8187);
nor UO_221 (O_221,N_8756,N_8189);
or UO_222 (O_222,N_8264,N_9843);
nor UO_223 (O_223,N_8790,N_9348);
nor UO_224 (O_224,N_9393,N_9062);
nand UO_225 (O_225,N_8258,N_8618);
or UO_226 (O_226,N_9349,N_9070);
or UO_227 (O_227,N_8025,N_9257);
xor UO_228 (O_228,N_8510,N_9655);
nor UO_229 (O_229,N_9611,N_9205);
xor UO_230 (O_230,N_9526,N_9998);
or UO_231 (O_231,N_8910,N_9992);
nand UO_232 (O_232,N_8686,N_9222);
nand UO_233 (O_233,N_9574,N_8653);
nor UO_234 (O_234,N_9267,N_8499);
or UO_235 (O_235,N_9037,N_9659);
xnor UO_236 (O_236,N_9138,N_8158);
or UO_237 (O_237,N_8246,N_9157);
and UO_238 (O_238,N_8345,N_8268);
or UO_239 (O_239,N_8864,N_8567);
or UO_240 (O_240,N_8733,N_8131);
nand UO_241 (O_241,N_9830,N_9264);
or UO_242 (O_242,N_9591,N_9446);
and UO_243 (O_243,N_8568,N_8362);
nor UO_244 (O_244,N_9463,N_8178);
nor UO_245 (O_245,N_9837,N_8887);
and UO_246 (O_246,N_9645,N_9683);
nand UO_247 (O_247,N_8808,N_9008);
nand UO_248 (O_248,N_9742,N_8418);
and UO_249 (O_249,N_8115,N_8332);
and UO_250 (O_250,N_8597,N_9443);
nand UO_251 (O_251,N_9388,N_8014);
nand UO_252 (O_252,N_9359,N_9935);
nor UO_253 (O_253,N_9360,N_8456);
nor UO_254 (O_254,N_8384,N_9983);
and UO_255 (O_255,N_9845,N_9164);
nor UO_256 (O_256,N_8616,N_9822);
or UO_257 (O_257,N_8441,N_8773);
nor UO_258 (O_258,N_9789,N_8710);
xor UO_259 (O_259,N_8660,N_9622);
nand UO_260 (O_260,N_9826,N_9170);
and UO_261 (O_261,N_8594,N_8927);
nor UO_262 (O_262,N_8505,N_8040);
nor UO_263 (O_263,N_8005,N_9265);
or UO_264 (O_264,N_9867,N_9345);
nor UO_265 (O_265,N_9542,N_9670);
nand UO_266 (O_266,N_9714,N_9297);
xnor UO_267 (O_267,N_8255,N_9118);
xor UO_268 (O_268,N_9487,N_9631);
nor UO_269 (O_269,N_8249,N_9474);
nand UO_270 (O_270,N_9543,N_9799);
or UO_271 (O_271,N_8725,N_8454);
and UO_272 (O_272,N_9832,N_9476);
or UO_273 (O_273,N_8218,N_9180);
nor UO_274 (O_274,N_8981,N_8847);
nand UO_275 (O_275,N_8333,N_8709);
nor UO_276 (O_276,N_8532,N_9968);
nor UO_277 (O_277,N_9629,N_8070);
or UO_278 (O_278,N_8986,N_8797);
and UO_279 (O_279,N_9296,N_9560);
nor UO_280 (O_280,N_8091,N_8495);
or UO_281 (O_281,N_9112,N_8233);
or UO_282 (O_282,N_8168,N_8061);
nor UO_283 (O_283,N_8290,N_9022);
xnor UO_284 (O_284,N_8379,N_9275);
nand UO_285 (O_285,N_8259,N_9326);
and UO_286 (O_286,N_9578,N_9106);
and UO_287 (O_287,N_9479,N_8033);
nor UO_288 (O_288,N_8350,N_8724);
nand UO_289 (O_289,N_8105,N_8397);
nand UO_290 (O_290,N_8672,N_8090);
nor UO_291 (O_291,N_8216,N_8631);
nand UO_292 (O_292,N_8396,N_9480);
nor UO_293 (O_293,N_9838,N_9279);
nand UO_294 (O_294,N_9450,N_9056);
nand UO_295 (O_295,N_9751,N_8726);
nor UO_296 (O_296,N_9471,N_8262);
xnor UO_297 (O_297,N_8188,N_8442);
and UO_298 (O_298,N_8087,N_8308);
nand UO_299 (O_299,N_8926,N_9707);
or UO_300 (O_300,N_9065,N_9414);
or UO_301 (O_301,N_9031,N_9972);
xnor UO_302 (O_302,N_9372,N_8789);
or UO_303 (O_303,N_9292,N_9351);
or UO_304 (O_304,N_9626,N_8096);
nand UO_305 (O_305,N_8179,N_8163);
nand UO_306 (O_306,N_8529,N_8298);
nor UO_307 (O_307,N_9870,N_9949);
nor UO_308 (O_308,N_8946,N_9530);
nor UO_309 (O_309,N_9906,N_9148);
or UO_310 (O_310,N_8195,N_8637);
nor UO_311 (O_311,N_8746,N_8892);
nor UO_312 (O_312,N_8437,N_9458);
nand UO_313 (O_313,N_9340,N_9131);
nor UO_314 (O_314,N_9756,N_9710);
nand UO_315 (O_315,N_9231,N_8776);
xnor UO_316 (O_316,N_8155,N_9963);
xor UO_317 (O_317,N_8995,N_9685);
xor UO_318 (O_318,N_9130,N_8895);
nor UO_319 (O_319,N_8433,N_8484);
nand UO_320 (O_320,N_9718,N_9033);
and UO_321 (O_321,N_8858,N_8731);
nor UO_322 (O_322,N_8161,N_8473);
nor UO_323 (O_323,N_9780,N_8666);
and UO_324 (O_324,N_8313,N_9942);
nor UO_325 (O_325,N_8072,N_8482);
nor UO_326 (O_326,N_9969,N_9398);
nor UO_327 (O_327,N_8602,N_8143);
nor UO_328 (O_328,N_9535,N_9248);
xor UO_329 (O_329,N_9058,N_8757);
and UO_330 (O_330,N_8747,N_8664);
or UO_331 (O_331,N_9484,N_9899);
and UO_332 (O_332,N_9876,N_9516);
nor UO_333 (O_333,N_9499,N_9332);
nor UO_334 (O_334,N_9945,N_8854);
nor UO_335 (O_335,N_8525,N_9862);
or UO_336 (O_336,N_9061,N_8315);
nand UO_337 (O_337,N_8027,N_9364);
nand UO_338 (O_338,N_8322,N_8665);
nand UO_339 (O_339,N_9967,N_8411);
nand UO_340 (O_340,N_8137,N_9977);
nor UO_341 (O_341,N_9921,N_8326);
or UO_342 (O_342,N_9738,N_8064);
nor UO_343 (O_343,N_9151,N_9533);
and UO_344 (O_344,N_9177,N_8114);
or UO_345 (O_345,N_8364,N_9762);
nand UO_346 (O_346,N_9045,N_9202);
nand UO_347 (O_347,N_9805,N_9765);
nand UO_348 (O_348,N_8535,N_8821);
nand UO_349 (O_349,N_9570,N_8967);
nor UO_350 (O_350,N_9353,N_9861);
or UO_351 (O_351,N_8828,N_9268);
or UO_352 (O_352,N_9575,N_9152);
nor UO_353 (O_353,N_9868,N_8047);
or UO_354 (O_354,N_9141,N_9588);
or UO_355 (O_355,N_9917,N_8374);
nor UO_356 (O_356,N_8966,N_8448);
and UO_357 (O_357,N_9551,N_9559);
or UO_358 (O_358,N_9189,N_9706);
and UO_359 (O_359,N_8011,N_9156);
or UO_360 (O_360,N_8497,N_9440);
xnor UO_361 (O_361,N_8924,N_8121);
nand UO_362 (O_362,N_9092,N_8338);
and UO_363 (O_363,N_9531,N_9455);
or UO_364 (O_364,N_9962,N_9964);
and UO_365 (O_365,N_8633,N_9052);
nor UO_366 (O_366,N_9696,N_8555);
nand UO_367 (O_367,N_8826,N_8771);
nor UO_368 (O_368,N_9386,N_8299);
and UO_369 (O_369,N_9853,N_8948);
nand UO_370 (O_370,N_8148,N_8656);
nand UO_371 (O_371,N_8867,N_8480);
and UO_372 (O_372,N_8586,N_9654);
or UO_373 (O_373,N_8339,N_8159);
xor UO_374 (O_374,N_9633,N_8311);
and UO_375 (O_375,N_9593,N_8928);
nor UO_376 (O_376,N_8777,N_8968);
or UO_377 (O_377,N_8220,N_9430);
or UO_378 (O_378,N_8650,N_9283);
and UO_379 (O_379,N_8208,N_9041);
xor UO_380 (O_380,N_8989,N_8531);
and UO_381 (O_381,N_8836,N_9833);
nor UO_382 (O_382,N_9653,N_9773);
and UO_383 (O_383,N_9192,N_9381);
or UO_384 (O_384,N_9431,N_9117);
nor UO_385 (O_385,N_8010,N_8034);
and UO_386 (O_386,N_8355,N_9527);
or UO_387 (O_387,N_8340,N_8068);
nor UO_388 (O_388,N_9563,N_8106);
nor UO_389 (O_389,N_8389,N_8655);
xnor UO_390 (O_390,N_8395,N_8151);
or UO_391 (O_391,N_8425,N_9885);
nand UO_392 (O_392,N_8812,N_8392);
and UO_393 (O_393,N_9958,N_8850);
and UO_394 (O_394,N_9509,N_8443);
and UO_395 (O_395,N_9054,N_9036);
and UO_396 (O_396,N_8649,N_9788);
and UO_397 (O_397,N_8282,N_8742);
nand UO_398 (O_398,N_9304,N_9988);
or UO_399 (O_399,N_9635,N_8580);
or UO_400 (O_400,N_8439,N_8994);
xnor UO_401 (O_401,N_8226,N_9094);
nor UO_402 (O_402,N_9668,N_9770);
and UO_403 (O_403,N_8045,N_9428);
nor UO_404 (O_404,N_8346,N_9380);
nor UO_405 (O_405,N_8059,N_9540);
or UO_406 (O_406,N_9068,N_9959);
xnor UO_407 (O_407,N_8751,N_8933);
nand UO_408 (O_408,N_8139,N_8078);
or UO_409 (O_409,N_9179,N_8075);
or UO_410 (O_410,N_8932,N_9737);
or UO_411 (O_411,N_8427,N_8694);
nand UO_412 (O_412,N_9887,N_9306);
and UO_413 (O_413,N_9881,N_9966);
nand UO_414 (O_414,N_8699,N_8893);
or UO_415 (O_415,N_9212,N_8561);
or UO_416 (O_416,N_8702,N_8288);
and UO_417 (O_417,N_8234,N_8622);
nand UO_418 (O_418,N_8611,N_8976);
or UO_419 (O_419,N_8669,N_8486);
nand UO_420 (O_420,N_8063,N_8174);
or UO_421 (O_421,N_9999,N_9486);
nand UO_422 (O_422,N_8972,N_8509);
and UO_423 (O_423,N_8675,N_8302);
or UO_424 (O_424,N_9253,N_9362);
and UO_425 (O_425,N_8574,N_8658);
nand UO_426 (O_426,N_8423,N_8554);
nand UO_427 (O_427,N_8569,N_8490);
nand UO_428 (O_428,N_9700,N_8755);
or UO_429 (O_429,N_9652,N_9167);
or UO_430 (O_430,N_8450,N_8030);
or UO_431 (O_431,N_8273,N_9059);
and UO_432 (O_432,N_8939,N_8760);
or UO_433 (O_433,N_8117,N_9472);
nor UO_434 (O_434,N_8110,N_9135);
or UO_435 (O_435,N_9539,N_9627);
or UO_436 (O_436,N_8344,N_8721);
nor UO_437 (O_437,N_8629,N_9067);
and UO_438 (O_438,N_8609,N_8224);
nand UO_439 (O_439,N_9643,N_8648);
nand UO_440 (O_440,N_9288,N_8706);
nand UO_441 (O_441,N_9869,N_8074);
xnor UO_442 (O_442,N_8232,N_9368);
and UO_443 (O_443,N_9286,N_9121);
or UO_444 (O_444,N_8644,N_9339);
nand UO_445 (O_445,N_8573,N_8079);
or UO_446 (O_446,N_8013,N_9373);
nor UO_447 (O_447,N_9794,N_8331);
and UO_448 (O_448,N_8407,N_8408);
or UO_449 (O_449,N_9077,N_8300);
nor UO_450 (O_450,N_9470,N_8461);
nand UO_451 (O_451,N_8800,N_9196);
nor UO_452 (O_452,N_8102,N_8677);
and UO_453 (O_453,N_9721,N_8381);
and UO_454 (O_454,N_9650,N_9800);
nor UO_455 (O_455,N_9673,N_9587);
or UO_456 (O_456,N_9993,N_8310);
and UO_457 (O_457,N_9247,N_9767);
or UO_458 (O_458,N_9970,N_8604);
nand UO_459 (O_459,N_9987,N_9418);
and UO_460 (O_460,N_8022,N_8896);
nor UO_461 (O_461,N_9473,N_9150);
and UO_462 (O_462,N_9628,N_8275);
or UO_463 (O_463,N_9776,N_8157);
nor UO_464 (O_464,N_9401,N_9119);
nor UO_465 (O_465,N_8784,N_9667);
nor UO_466 (O_466,N_8371,N_8316);
nand UO_467 (O_467,N_8857,N_9161);
xor UO_468 (O_468,N_8270,N_8588);
nand UO_469 (O_469,N_8919,N_9249);
nor UO_470 (O_470,N_9517,N_8431);
nor UO_471 (O_471,N_9690,N_8860);
or UO_472 (O_472,N_8791,N_8545);
or UO_473 (O_473,N_9405,N_9107);
nor UO_474 (O_474,N_8834,N_9774);
nand UO_475 (O_475,N_8572,N_9960);
nand UO_476 (O_476,N_9178,N_8329);
nand UO_477 (O_477,N_9584,N_8947);
or UO_478 (O_478,N_9656,N_9242);
or UO_479 (O_479,N_9464,N_8167);
and UO_480 (O_480,N_9736,N_9282);
nor UO_481 (O_481,N_8035,N_9089);
nand UO_482 (O_482,N_8513,N_9608);
nor UO_483 (O_483,N_8518,N_8596);
nand UO_484 (O_484,N_8842,N_8652);
and UO_485 (O_485,N_9408,N_9743);
nand UO_486 (O_486,N_8165,N_8459);
and UO_487 (O_487,N_8508,N_8719);
and UO_488 (O_488,N_9879,N_9865);
nand UO_489 (O_489,N_9493,N_8815);
and UO_490 (O_490,N_8662,N_9079);
or UO_491 (O_491,N_8683,N_9649);
and UO_492 (O_492,N_9975,N_8657);
nor UO_493 (O_493,N_8293,N_9366);
nand UO_494 (O_494,N_9254,N_8292);
nand UO_495 (O_495,N_8587,N_8521);
nand UO_496 (O_496,N_8227,N_9389);
or UO_497 (O_497,N_9807,N_9760);
nor UO_498 (O_498,N_9613,N_9336);
nand UO_499 (O_499,N_8758,N_9604);
or UO_500 (O_500,N_8094,N_8865);
or UO_501 (O_501,N_9337,N_8565);
and UO_502 (O_502,N_8879,N_9614);
nor UO_503 (O_503,N_8717,N_9739);
and UO_504 (O_504,N_8058,N_8781);
nor UO_505 (O_505,N_8471,N_9692);
nor UO_506 (O_506,N_8890,N_8191);
and UO_507 (O_507,N_9424,N_9334);
nor UO_508 (O_508,N_9096,N_8681);
or UO_509 (O_509,N_8563,N_9404);
xnor UO_510 (O_510,N_8813,N_9488);
or UO_511 (O_511,N_9016,N_8740);
or UO_512 (O_512,N_9203,N_8774);
nand UO_513 (O_513,N_8500,N_9731);
nand UO_514 (O_514,N_8806,N_8730);
or UO_515 (O_515,N_9447,N_9971);
xor UO_516 (O_516,N_9732,N_9137);
or UO_517 (O_517,N_8126,N_9990);
nor UO_518 (O_518,N_9644,N_9290);
or UO_519 (O_519,N_9734,N_9585);
nor UO_520 (O_520,N_8827,N_9042);
nand UO_521 (O_521,N_9634,N_8612);
nor UO_522 (O_522,N_8241,N_8351);
and UO_523 (O_523,N_9050,N_8544);
nor UO_524 (O_524,N_8228,N_9727);
or UO_525 (O_525,N_8162,N_9566);
and UO_526 (O_526,N_8388,N_9842);
or UO_527 (O_527,N_8366,N_9095);
or UO_528 (O_528,N_8852,N_9529);
nor UO_529 (O_529,N_9356,N_8905);
or UO_530 (O_530,N_9343,N_9565);
nor UO_531 (O_531,N_8621,N_8123);
nor UO_532 (O_532,N_9011,N_9017);
nor UO_533 (O_533,N_8267,N_8820);
xnor UO_534 (O_534,N_8651,N_9664);
nor UO_535 (O_535,N_9015,N_9699);
xor UO_536 (O_536,N_8065,N_9609);
nand UO_537 (O_537,N_8775,N_8285);
or UO_538 (O_538,N_9145,N_9630);
and UO_539 (O_539,N_9893,N_9129);
nor UO_540 (O_540,N_9923,N_9048);
xor UO_541 (O_541,N_8944,N_8048);
xor UO_542 (O_542,N_9181,N_9127);
and UO_543 (O_543,N_8481,N_8135);
and UO_544 (O_544,N_9160,N_8348);
and UO_545 (O_545,N_8184,N_8046);
or UO_546 (O_546,N_8318,N_8197);
and UO_547 (O_547,N_9330,N_8802);
nand UO_548 (O_548,N_9702,N_9813);
or UO_549 (O_549,N_8974,N_9099);
nand UO_550 (O_550,N_8301,N_8200);
nor UO_551 (O_551,N_9847,N_8767);
xor UO_552 (O_552,N_9852,N_9220);
and UO_553 (O_553,N_9528,N_9772);
nor UO_554 (O_554,N_8136,N_9503);
or UO_555 (O_555,N_9801,N_9605);
and UO_556 (O_556,N_9658,N_8071);
or UO_557 (O_557,N_8835,N_9695);
nor UO_558 (O_558,N_9001,N_9550);
and UO_559 (O_559,N_8470,N_9811);
xnor UO_560 (O_560,N_8449,N_8266);
and UO_561 (O_561,N_9510,N_8453);
and UO_562 (O_562,N_9213,N_8607);
and UO_563 (O_563,N_9437,N_9402);
or UO_564 (O_564,N_9717,N_8043);
or UO_565 (O_565,N_8172,N_8603);
or UO_566 (O_566,N_8739,N_9173);
and UO_567 (O_567,N_9929,N_8538);
xnor UO_568 (O_568,N_9142,N_9994);
and UO_569 (O_569,N_8929,N_9835);
nor UO_570 (O_570,N_8982,N_9674);
nand UO_571 (O_571,N_9412,N_9687);
nand UO_572 (O_572,N_8349,N_8129);
and UO_573 (O_573,N_9420,N_9299);
nor UO_574 (O_574,N_8036,N_9396);
and UO_575 (O_575,N_8562,N_8076);
and UO_576 (O_576,N_8305,N_9483);
xnor UO_577 (O_577,N_8937,N_8417);
nand UO_578 (O_578,N_8578,N_8391);
and UO_579 (O_579,N_8307,N_8504);
or UO_580 (O_580,N_8250,N_9285);
nand UO_581 (O_581,N_8768,N_8401);
nor UO_582 (O_582,N_8883,N_8985);
nand UO_583 (O_583,N_9002,N_9808);
nand UO_584 (O_584,N_8062,N_8183);
or UO_585 (O_585,N_8051,N_8907);
or UO_586 (O_586,N_9888,N_8256);
nand UO_587 (O_587,N_8613,N_9102);
nand UO_588 (O_588,N_8671,N_8274);
nand UO_589 (O_589,N_8787,N_9195);
nor UO_590 (O_590,N_8357,N_8993);
nor UO_591 (O_591,N_9938,N_9165);
or UO_592 (O_592,N_8943,N_8287);
or UO_593 (O_593,N_9797,N_9980);
nand UO_594 (O_594,N_9445,N_9525);
nor UO_595 (O_595,N_8186,N_9442);
nor UO_596 (O_596,N_9705,N_8175);
nor UO_597 (O_597,N_8377,N_9315);
or UO_598 (O_598,N_9301,N_8457);
or UO_599 (O_599,N_8844,N_8991);
or UO_600 (O_600,N_9639,N_9657);
nor UO_601 (O_601,N_8406,N_8492);
or UO_602 (O_602,N_9097,N_9924);
and UO_603 (O_603,N_8026,N_8534);
or UO_604 (O_604,N_9750,N_9669);
and UO_605 (O_605,N_9312,N_9930);
and UO_606 (O_606,N_9701,N_9892);
or UO_607 (O_607,N_8996,N_9976);
or UO_608 (O_608,N_9973,N_8522);
xnor UO_609 (O_609,N_9919,N_8277);
or UO_610 (O_610,N_8630,N_9748);
or UO_611 (O_611,N_9567,N_9619);
nor UO_612 (O_612,N_9905,N_9777);
nor UO_613 (O_613,N_8524,N_8387);
nand UO_614 (O_614,N_9194,N_9091);
and UO_615 (O_615,N_8474,N_9623);
nand UO_616 (O_616,N_9200,N_8019);
and UO_617 (O_617,N_9778,N_9747);
nand UO_618 (O_618,N_8909,N_8097);
and UO_619 (O_619,N_8668,N_8002);
and UO_620 (O_620,N_9171,N_8738);
and UO_621 (O_621,N_9435,N_9163);
xnor UO_622 (O_622,N_8103,N_9357);
and UO_623 (O_623,N_8082,N_8917);
and UO_624 (O_624,N_9105,N_8007);
or UO_625 (O_625,N_8498,N_9638);
and UO_626 (O_626,N_9277,N_8445);
nor UO_627 (O_627,N_9478,N_8780);
nor UO_628 (O_628,N_9467,N_8698);
or UO_629 (O_629,N_9263,N_9761);
and UO_630 (O_630,N_8619,N_8723);
nand UO_631 (O_631,N_8727,N_9840);
and UO_632 (O_632,N_8934,N_9907);
nand UO_633 (O_633,N_8247,N_8325);
and UO_634 (O_634,N_8634,N_9891);
nor UO_635 (O_635,N_8691,N_9908);
nand UO_636 (O_636,N_8788,N_9328);
and UO_637 (O_637,N_9561,N_8743);
and UO_638 (O_638,N_9595,N_8589);
nor UO_639 (O_639,N_8251,N_9219);
and UO_640 (O_640,N_8626,N_8080);
nand UO_641 (O_641,N_9278,N_8067);
or UO_642 (O_642,N_9564,N_8337);
or UO_643 (O_643,N_8215,N_8980);
or UO_644 (O_644,N_9779,N_9709);
nor UO_645 (O_645,N_9764,N_9271);
xnor UO_646 (O_646,N_8223,N_9694);
nor UO_647 (O_647,N_8252,N_8819);
xor UO_648 (O_648,N_9444,N_9894);
nand UO_649 (O_649,N_9612,N_9259);
and UO_650 (O_650,N_9795,N_8557);
and UO_651 (O_651,N_8703,N_9758);
and UO_652 (O_652,N_9361,N_8697);
nand UO_653 (O_653,N_9224,N_9427);
or UO_654 (O_654,N_9855,N_8999);
nor UO_655 (O_655,N_9269,N_8667);
nand UO_656 (O_656,N_9433,N_9025);
or UO_657 (O_657,N_9303,N_9169);
nor UO_658 (O_658,N_9035,N_8309);
or UO_659 (O_659,N_8056,N_8152);
nor UO_660 (O_660,N_9198,N_8900);
and UO_661 (O_661,N_8501,N_9226);
or UO_662 (O_662,N_9932,N_8941);
nand UO_663 (O_663,N_8479,N_8133);
nand UO_664 (O_664,N_9816,N_8419);
nor UO_665 (O_665,N_9864,N_8375);
nand UO_666 (O_666,N_9153,N_8705);
nand UO_667 (O_667,N_9937,N_9144);
or UO_668 (O_668,N_8749,N_9641);
nand UO_669 (O_669,N_9060,N_8198);
nand UO_670 (O_670,N_9896,N_9123);
xor UO_671 (O_671,N_9817,N_9538);
nand UO_672 (O_672,N_9759,N_8765);
or UO_673 (O_673,N_9895,N_8839);
or UO_674 (O_674,N_8759,N_8541);
nand UO_675 (O_675,N_9255,N_8801);
nor UO_676 (O_676,N_8785,N_9392);
or UO_677 (O_677,N_9646,N_8491);
nor UO_678 (O_678,N_8809,N_8069);
or UO_679 (O_679,N_8354,N_8225);
or UO_680 (O_680,N_9740,N_9325);
xnor UO_681 (O_681,N_8269,N_8983);
or UO_682 (O_682,N_8244,N_8810);
and UO_683 (O_683,N_9046,N_9810);
nor UO_684 (O_684,N_9675,N_9187);
nor UO_685 (O_685,N_9632,N_9316);
nor UO_686 (O_686,N_9302,N_9227);
and UO_687 (O_687,N_9537,N_9512);
nor UO_688 (O_688,N_9039,N_9394);
or UO_689 (O_689,N_8921,N_8945);
or UO_690 (O_690,N_8741,N_9027);
nand UO_691 (O_691,N_9884,N_9413);
nand UO_692 (O_692,N_8690,N_9240);
or UO_693 (O_693,N_8358,N_9716);
nor UO_694 (O_694,N_9071,N_9601);
nor UO_695 (O_695,N_9934,N_8084);
and UO_696 (O_696,N_8347,N_8506);
nor UO_697 (O_697,N_9558,N_8049);
nor UO_698 (O_698,N_9358,N_9115);
nor UO_699 (O_699,N_8496,N_8978);
nor UO_700 (O_700,N_8475,N_9075);
nor UO_701 (O_701,N_8517,N_9298);
and UO_702 (O_702,N_9534,N_9252);
xnor UO_703 (O_703,N_9677,N_9557);
nor UO_704 (O_704,N_9204,N_8422);
nand UO_705 (O_705,N_9965,N_9122);
xor UO_706 (O_706,N_8276,N_8483);
and UO_707 (O_707,N_8466,N_8462);
or UO_708 (O_708,N_8196,N_8969);
and UO_709 (O_709,N_9363,N_9766);
nor UO_710 (O_710,N_8973,N_8954);
and UO_711 (O_711,N_9383,N_8997);
or UO_712 (O_712,N_8319,N_9261);
nor UO_713 (O_713,N_9441,N_8112);
nand UO_714 (O_714,N_9621,N_9436);
or UO_715 (O_715,N_9193,N_8627);
or UO_716 (O_716,N_9590,N_8294);
and UO_717 (O_717,N_8263,N_9462);
or UO_718 (O_718,N_8193,N_9839);
nor UO_719 (O_719,N_9981,N_8936);
nor UO_720 (O_720,N_9191,N_9088);
or UO_721 (O_721,N_8296,N_8872);
or UO_722 (O_722,N_8970,N_8057);
nor UO_723 (O_723,N_8089,N_9053);
and UO_724 (O_724,N_9323,N_8098);
xor UO_725 (O_725,N_9724,N_9961);
nor UO_726 (O_726,N_8150,N_9333);
nor UO_727 (O_727,N_9886,N_8911);
and UO_728 (O_728,N_9524,N_8312);
or UO_729 (O_729,N_9686,N_9544);
nand UO_730 (O_730,N_8796,N_9244);
and UO_731 (O_731,N_9933,N_8050);
nand UO_732 (O_732,N_8598,N_9580);
nor UO_733 (O_733,N_9072,N_8303);
nand UO_734 (O_734,N_9596,N_8494);
nor UO_735 (O_735,N_9010,N_9790);
nor UO_736 (O_736,N_8458,N_9502);
and UO_737 (O_737,N_9409,N_9294);
or UO_738 (O_738,N_9270,N_8542);
and UO_739 (O_739,N_9300,N_8891);
nor UO_740 (O_740,N_9834,N_9064);
nand UO_741 (O_741,N_8795,N_9367);
nor UO_742 (O_742,N_9258,N_8680);
nand UO_743 (O_743,N_8861,N_9521);
or UO_744 (O_744,N_8032,N_9390);
nand UO_745 (O_745,N_8876,N_8147);
and UO_746 (O_746,N_9374,N_8830);
or UO_747 (O_747,N_8360,N_8878);
and UO_748 (O_748,N_9598,N_9085);
and UO_749 (O_749,N_8125,N_8493);
nand UO_750 (O_750,N_8527,N_8214);
nor UO_751 (O_751,N_9208,N_9004);
nor UO_752 (O_752,N_9370,N_8211);
nand UO_753 (O_753,N_8695,N_8979);
or UO_754 (O_754,N_8822,N_9890);
nor UO_755 (O_755,N_9076,N_9322);
nand UO_756 (O_756,N_8786,N_8181);
nor UO_757 (O_757,N_8866,N_8564);
or UO_758 (O_758,N_8066,N_9188);
nand UO_759 (O_759,N_9504,N_9666);
and UO_760 (O_760,N_8590,N_9931);
nor UO_761 (O_761,N_9572,N_9403);
xor UO_762 (O_762,N_9744,N_8421);
nand UO_763 (O_763,N_8383,N_8297);
and UO_764 (O_764,N_9104,N_8643);
nand UO_765 (O_765,N_9376,N_8291);
and UO_766 (O_766,N_9783,N_8478);
nor UO_767 (O_767,N_8476,N_9355);
or UO_768 (O_768,N_8888,N_8434);
or UO_769 (O_769,N_9606,N_8378);
nor UO_770 (O_770,N_8678,N_8571);
nor UO_771 (O_771,N_9925,N_9172);
nand UO_772 (O_772,N_8595,N_9218);
xnor UO_773 (O_773,N_8410,N_8849);
nand UO_774 (O_774,N_8940,N_9711);
and UO_775 (O_775,N_8831,N_9197);
or UO_776 (O_776,N_9057,N_8951);
and UO_777 (O_777,N_9820,N_9216);
or UO_778 (O_778,N_8577,N_8185);
or UO_779 (O_779,N_8488,N_8988);
or UO_780 (O_780,N_9599,N_9520);
and UO_781 (O_781,N_9344,N_8753);
nor UO_782 (O_782,N_9583,N_9168);
nor UO_783 (O_783,N_8770,N_8707);
or UO_784 (O_784,N_8750,N_9098);
or UO_785 (O_785,N_8886,N_9477);
and UO_786 (O_786,N_9781,N_8824);
and UO_787 (O_787,N_9176,N_9829);
nand UO_788 (O_788,N_9234,N_8242);
xor UO_789 (O_789,N_8237,N_8420);
or UO_790 (O_790,N_8654,N_9511);
nor UO_791 (O_791,N_8254,N_8052);
or UO_792 (O_792,N_8444,N_9214);
nor UO_793 (O_793,N_9802,N_9055);
nand UO_794 (O_794,N_9223,N_8230);
nand UO_795 (O_795,N_8884,N_8201);
nand UO_796 (O_796,N_9607,N_8984);
nor UO_797 (O_797,N_9722,N_8243);
nor UO_798 (O_798,N_8873,N_8779);
nor UO_799 (O_799,N_8539,N_8472);
or UO_800 (O_800,N_9648,N_8039);
nor UO_801 (O_801,N_8083,N_8582);
nor UO_802 (O_802,N_8794,N_9289);
nor UO_803 (O_803,N_8130,N_8146);
or UO_804 (O_804,N_8962,N_8745);
or UO_805 (O_805,N_9114,N_8870);
nor UO_806 (O_806,N_9309,N_9452);
nor UO_807 (O_807,N_9536,N_9926);
and UO_808 (O_808,N_9331,N_9941);
nand UO_809 (O_809,N_9665,N_9723);
or UO_810 (O_810,N_9508,N_8400);
and UO_811 (O_811,N_9871,N_9018);
nor UO_812 (O_812,N_9276,N_9883);
nand UO_813 (O_813,N_8543,N_8295);
xor UO_814 (O_814,N_8205,N_8516);
or UO_815 (O_815,N_8841,N_8869);
or UO_816 (O_816,N_8236,N_9792);
nand UO_817 (O_817,N_9416,N_9233);
and UO_818 (O_818,N_9132,N_8960);
nand UO_819 (O_819,N_9155,N_8772);
or UO_820 (O_820,N_8012,N_8992);
and UO_821 (O_821,N_9235,N_9354);
nor UO_822 (O_822,N_8576,N_9793);
nor UO_823 (O_823,N_9752,N_9877);
or UO_824 (O_824,N_8882,N_9082);
or UO_825 (O_825,N_9426,N_8382);
nand UO_826 (O_826,N_9457,N_8194);
nor UO_827 (O_827,N_8606,N_8515);
or UO_828 (O_828,N_8166,N_8605);
xor UO_829 (O_829,N_9944,N_9828);
nor UO_830 (O_830,N_9407,N_9109);
xnor UO_831 (O_831,N_8000,N_8324);
and UO_832 (O_832,N_8429,N_8336);
or UO_833 (O_833,N_8286,N_8041);
nand UO_834 (O_834,N_8931,N_8190);
nand UO_835 (O_835,N_9577,N_8248);
and UO_836 (O_836,N_8368,N_9399);
nand UO_837 (O_837,N_8317,N_9120);
or UO_838 (O_838,N_9878,N_9844);
and UO_839 (O_839,N_8718,N_8914);
nor UO_840 (O_840,N_9848,N_8222);
nor UO_841 (O_841,N_9662,N_8856);
or UO_842 (O_842,N_8894,N_8949);
nand UO_843 (O_843,N_8024,N_8807);
nand UO_844 (O_844,N_8330,N_9678);
nor UO_845 (O_845,N_8851,N_9063);
or UO_846 (O_846,N_8708,N_8009);
nand UO_847 (O_847,N_9556,N_8679);
and UO_848 (O_848,N_9849,N_9346);
or UO_849 (O_849,N_8560,N_9347);
nand UO_850 (O_850,N_8902,N_9461);
nor UO_851 (O_851,N_9074,N_8647);
nor UO_852 (O_852,N_9841,N_9819);
and UO_853 (O_853,N_9496,N_8990);
or UO_854 (O_854,N_8240,N_8405);
nand UO_855 (O_855,N_8859,N_8692);
and UO_856 (O_856,N_8583,N_9952);
nand UO_857 (O_857,N_8004,N_9456);
nor UO_858 (O_858,N_9522,N_8639);
or UO_859 (O_859,N_9787,N_8635);
and UO_860 (O_860,N_9823,N_8700);
and UO_861 (O_861,N_9704,N_8661);
xnor UO_862 (O_862,N_8614,N_9660);
nand UO_863 (O_863,N_8073,N_8804);
or UO_864 (O_864,N_9274,N_9417);
or UO_865 (O_865,N_8502,N_9239);
nor UO_866 (O_866,N_8468,N_9047);
and UO_867 (O_867,N_9821,N_9946);
nor UO_868 (O_868,N_9338,N_9900);
or UO_869 (O_869,N_8528,N_8279);
nor UO_870 (O_870,N_8880,N_8053);
xnor UO_871 (O_871,N_8436,N_8060);
nor UO_872 (O_872,N_9023,N_9997);
and UO_873 (O_873,N_8925,N_8424);
or UO_874 (O_874,N_8414,N_9162);
and UO_875 (O_875,N_8023,N_9318);
or UO_876 (O_876,N_9215,N_9365);
nor UO_877 (O_877,N_9592,N_8265);
nand UO_878 (O_878,N_8177,N_8959);
or UO_879 (O_879,N_9827,N_9836);
or UO_880 (O_880,N_9989,N_8955);
nand UO_881 (O_881,N_9712,N_9579);
and UO_882 (O_882,N_9571,N_8556);
and UO_883 (O_883,N_9547,N_8104);
nand UO_884 (O_884,N_9618,N_8253);
nor UO_885 (O_885,N_9460,N_8320);
nor UO_886 (O_886,N_9280,N_9775);
nor UO_887 (O_887,N_9680,N_9038);
or UO_888 (O_888,N_8095,N_8624);
or UO_889 (O_889,N_9939,N_8128);
or UO_890 (O_890,N_9698,N_9866);
xor UO_891 (O_891,N_8393,N_9620);
or UO_892 (O_892,N_9689,N_8160);
nor UO_893 (O_893,N_8451,N_9190);
nand UO_894 (O_894,N_9342,N_9863);
or UO_895 (O_895,N_8840,N_8464);
nand UO_896 (O_896,N_9108,N_8918);
nand UO_897 (O_897,N_9093,N_9491);
nand UO_898 (O_898,N_9284,N_8428);
or UO_899 (O_899,N_9066,N_9481);
nand UO_900 (O_900,N_9238,N_9730);
or UO_901 (O_901,N_9625,N_9693);
nor UO_902 (O_902,N_9552,N_8463);
nand UO_903 (O_903,N_8144,N_8134);
and UO_904 (O_904,N_9726,N_8540);
xor UO_905 (O_905,N_9083,N_9310);
or UO_906 (O_906,N_9327,N_8365);
and UO_907 (O_907,N_9101,N_9397);
or UO_908 (O_908,N_9991,N_9419);
or UO_909 (O_909,N_8018,N_9411);
xnor UO_910 (O_910,N_8438,N_8031);
nand UO_911 (O_911,N_9672,N_8394);
and UO_912 (O_912,N_8938,N_8409);
nor UO_913 (O_913,N_9953,N_8638);
or UO_914 (O_914,N_8042,N_8687);
or UO_915 (O_915,N_8871,N_9174);
or UO_916 (O_916,N_9982,N_9913);
nor UO_917 (O_917,N_8156,N_8182);
or UO_918 (O_918,N_8736,N_9681);
nand UO_919 (O_919,N_8920,N_9228);
nor UO_920 (O_920,N_8140,N_9241);
or UO_921 (O_921,N_9642,N_8625);
nor UO_922 (O_922,N_9594,N_9021);
nor UO_923 (O_923,N_8403,N_8533);
nor UO_924 (O_924,N_9735,N_9308);
or UO_925 (O_925,N_8192,N_8975);
or UO_926 (O_926,N_9497,N_8734);
nand UO_927 (O_927,N_9676,N_8124);
nand UO_928 (O_928,N_9272,N_8971);
or UO_929 (O_929,N_8916,N_9691);
nor UO_930 (O_930,N_9139,N_9159);
nand UO_931 (O_931,N_9043,N_9553);
nor UO_932 (O_932,N_8935,N_9733);
and UO_933 (O_933,N_8620,N_8008);
and UO_934 (O_934,N_9875,N_9032);
and UO_935 (O_935,N_9028,N_8843);
and UO_936 (O_936,N_9603,N_8763);
nand UO_937 (O_937,N_8615,N_9199);
and UO_938 (O_938,N_9305,N_9545);
nor UO_939 (O_939,N_9049,N_9697);
or UO_940 (O_940,N_9084,N_8323);
nand UO_941 (O_941,N_9250,N_9128);
nand UO_942 (O_942,N_8465,N_9610);
nand UO_943 (O_943,N_9201,N_8875);
or UO_944 (O_944,N_8306,N_9029);
and UO_945 (O_945,N_9324,N_8169);
nor UO_946 (O_946,N_8897,N_9378);
and UO_947 (O_947,N_8260,N_9506);
and UO_948 (O_948,N_8636,N_8507);
nor UO_949 (O_949,N_9720,N_8111);
and UO_950 (O_950,N_8029,N_9568);
nor UO_951 (O_951,N_8579,N_8093);
nand UO_952 (O_952,N_8171,N_8101);
or UO_953 (O_953,N_8020,N_8221);
nor UO_954 (O_954,N_9916,N_9500);
nand UO_955 (O_955,N_9451,N_9501);
nor UO_956 (O_956,N_9546,N_9815);
nand UO_957 (O_957,N_9291,N_8526);
and UO_958 (O_958,N_9880,N_8838);
and UO_959 (O_959,N_9786,N_9154);
xnor UO_960 (O_960,N_9030,N_9080);
and UO_961 (O_961,N_8361,N_8469);
nor UO_962 (O_962,N_8452,N_9985);
nor UO_963 (O_963,N_9013,N_9784);
and UO_964 (O_964,N_8693,N_9995);
or UO_965 (O_965,N_8592,N_9684);
or UO_966 (O_966,N_9005,N_9874);
or UO_967 (O_967,N_9920,N_9371);
nor UO_968 (O_968,N_9221,N_9514);
xnor UO_969 (O_969,N_8930,N_8584);
nand UO_970 (O_970,N_8599,N_8283);
nor UO_971 (O_971,N_9569,N_9147);
and UO_972 (O_972,N_9688,N_8180);
xnor UO_973 (O_973,N_9262,N_9454);
or UO_974 (O_974,N_9287,N_9912);
and UO_975 (O_975,N_8015,N_8314);
or UO_976 (O_976,N_8402,N_9708);
nor UO_977 (O_977,N_9475,N_8908);
or UO_978 (O_978,N_8803,N_9415);
and UO_979 (O_979,N_8769,N_9186);
nand UO_980 (O_980,N_8874,N_9229);
nand UO_981 (O_981,N_9020,N_9136);
nand UO_982 (O_982,N_8352,N_9321);
and UO_983 (O_983,N_8231,N_9293);
nand UO_984 (O_984,N_8487,N_9246);
xor UO_985 (O_985,N_8913,N_8006);
xnor UO_986 (O_986,N_9812,N_8670);
and UO_987 (O_987,N_9682,N_9236);
or UO_988 (O_988,N_9979,N_9549);
and UO_989 (O_989,N_8904,N_9014);
nand UO_990 (O_990,N_8119,N_8141);
and UO_991 (O_991,N_9984,N_8304);
nand UO_992 (O_992,N_8154,N_9882);
nor UO_993 (O_993,N_8028,N_9513);
or UO_994 (O_994,N_8021,N_9485);
nand UO_995 (O_995,N_8748,N_9806);
nand UO_996 (O_996,N_8512,N_9019);
and UO_997 (O_997,N_8173,N_8641);
nand UO_998 (O_998,N_9078,N_9385);
nand UO_999 (O_999,N_8877,N_8552);
or UO_1000 (O_1000,N_9196,N_8445);
and UO_1001 (O_1001,N_8245,N_9887);
or UO_1002 (O_1002,N_8063,N_9287);
nand UO_1003 (O_1003,N_8600,N_9701);
nor UO_1004 (O_1004,N_8192,N_8750);
and UO_1005 (O_1005,N_8102,N_9409);
nand UO_1006 (O_1006,N_9424,N_9892);
or UO_1007 (O_1007,N_9022,N_8343);
xor UO_1008 (O_1008,N_8718,N_8414);
xnor UO_1009 (O_1009,N_9868,N_9554);
and UO_1010 (O_1010,N_9551,N_9736);
and UO_1011 (O_1011,N_8532,N_8247);
nor UO_1012 (O_1012,N_9469,N_9265);
nor UO_1013 (O_1013,N_9482,N_9978);
or UO_1014 (O_1014,N_9903,N_9680);
and UO_1015 (O_1015,N_9509,N_9907);
or UO_1016 (O_1016,N_9395,N_8002);
xnor UO_1017 (O_1017,N_8032,N_8904);
nand UO_1018 (O_1018,N_8311,N_8953);
nor UO_1019 (O_1019,N_8484,N_8337);
nor UO_1020 (O_1020,N_8201,N_8230);
nand UO_1021 (O_1021,N_9940,N_9799);
or UO_1022 (O_1022,N_8487,N_9765);
nand UO_1023 (O_1023,N_8966,N_8200);
nor UO_1024 (O_1024,N_8140,N_9196);
or UO_1025 (O_1025,N_8830,N_9552);
nor UO_1026 (O_1026,N_9892,N_9311);
and UO_1027 (O_1027,N_9989,N_9340);
and UO_1028 (O_1028,N_9993,N_8667);
nand UO_1029 (O_1029,N_9223,N_9476);
or UO_1030 (O_1030,N_9466,N_8443);
nor UO_1031 (O_1031,N_8355,N_9447);
and UO_1032 (O_1032,N_9813,N_8577);
xor UO_1033 (O_1033,N_9923,N_9075);
nor UO_1034 (O_1034,N_9506,N_9833);
nor UO_1035 (O_1035,N_8203,N_9488);
and UO_1036 (O_1036,N_9105,N_8002);
nand UO_1037 (O_1037,N_8535,N_9332);
nand UO_1038 (O_1038,N_8389,N_9063);
or UO_1039 (O_1039,N_9804,N_8425);
nor UO_1040 (O_1040,N_9784,N_9123);
or UO_1041 (O_1041,N_8461,N_9614);
and UO_1042 (O_1042,N_8118,N_8001);
or UO_1043 (O_1043,N_9302,N_8555);
and UO_1044 (O_1044,N_8505,N_9218);
or UO_1045 (O_1045,N_9926,N_9540);
nor UO_1046 (O_1046,N_9026,N_9718);
nor UO_1047 (O_1047,N_8340,N_9993);
nand UO_1048 (O_1048,N_8243,N_9032);
nand UO_1049 (O_1049,N_8010,N_9686);
or UO_1050 (O_1050,N_8253,N_9815);
nor UO_1051 (O_1051,N_9191,N_8121);
or UO_1052 (O_1052,N_9322,N_8297);
nand UO_1053 (O_1053,N_8583,N_9514);
nand UO_1054 (O_1054,N_8580,N_9782);
and UO_1055 (O_1055,N_9648,N_9393);
xor UO_1056 (O_1056,N_9333,N_9911);
and UO_1057 (O_1057,N_8130,N_9361);
nand UO_1058 (O_1058,N_9927,N_9068);
nand UO_1059 (O_1059,N_8661,N_8619);
nor UO_1060 (O_1060,N_8240,N_8358);
nor UO_1061 (O_1061,N_9908,N_8431);
or UO_1062 (O_1062,N_9202,N_9014);
nand UO_1063 (O_1063,N_8194,N_8610);
nand UO_1064 (O_1064,N_8062,N_8509);
or UO_1065 (O_1065,N_9439,N_9037);
nor UO_1066 (O_1066,N_9350,N_9475);
and UO_1067 (O_1067,N_9318,N_9395);
nor UO_1068 (O_1068,N_9637,N_9382);
nand UO_1069 (O_1069,N_9652,N_8376);
or UO_1070 (O_1070,N_8281,N_9895);
nor UO_1071 (O_1071,N_8315,N_9413);
nand UO_1072 (O_1072,N_9013,N_8920);
nor UO_1073 (O_1073,N_9585,N_8981);
xor UO_1074 (O_1074,N_9493,N_8000);
and UO_1075 (O_1075,N_9781,N_9716);
or UO_1076 (O_1076,N_8149,N_8840);
nand UO_1077 (O_1077,N_8755,N_8463);
and UO_1078 (O_1078,N_8769,N_9214);
or UO_1079 (O_1079,N_9362,N_8378);
and UO_1080 (O_1080,N_8228,N_9389);
and UO_1081 (O_1081,N_9192,N_8751);
and UO_1082 (O_1082,N_8367,N_8758);
nand UO_1083 (O_1083,N_9898,N_8942);
and UO_1084 (O_1084,N_9873,N_8156);
or UO_1085 (O_1085,N_9283,N_8298);
and UO_1086 (O_1086,N_9177,N_9684);
and UO_1087 (O_1087,N_9964,N_8746);
nor UO_1088 (O_1088,N_9105,N_9229);
nor UO_1089 (O_1089,N_9762,N_9230);
and UO_1090 (O_1090,N_8553,N_9877);
or UO_1091 (O_1091,N_8769,N_8860);
or UO_1092 (O_1092,N_8420,N_8742);
nor UO_1093 (O_1093,N_8103,N_8705);
xor UO_1094 (O_1094,N_8687,N_8181);
xnor UO_1095 (O_1095,N_8955,N_9954);
nor UO_1096 (O_1096,N_8713,N_8338);
xnor UO_1097 (O_1097,N_8967,N_9155);
nor UO_1098 (O_1098,N_9755,N_9632);
or UO_1099 (O_1099,N_9674,N_9611);
nor UO_1100 (O_1100,N_8851,N_8652);
and UO_1101 (O_1101,N_9956,N_8690);
nand UO_1102 (O_1102,N_8938,N_8702);
xnor UO_1103 (O_1103,N_8848,N_8768);
nand UO_1104 (O_1104,N_9037,N_9880);
and UO_1105 (O_1105,N_8603,N_9765);
or UO_1106 (O_1106,N_8740,N_8683);
and UO_1107 (O_1107,N_9130,N_9594);
or UO_1108 (O_1108,N_8389,N_8218);
nor UO_1109 (O_1109,N_8770,N_9987);
nand UO_1110 (O_1110,N_8312,N_9497);
or UO_1111 (O_1111,N_9995,N_8499);
or UO_1112 (O_1112,N_9227,N_9893);
or UO_1113 (O_1113,N_8447,N_9879);
nor UO_1114 (O_1114,N_9445,N_9364);
nor UO_1115 (O_1115,N_8910,N_8241);
or UO_1116 (O_1116,N_9665,N_8772);
nor UO_1117 (O_1117,N_9353,N_8719);
nand UO_1118 (O_1118,N_9434,N_8238);
xnor UO_1119 (O_1119,N_8599,N_8475);
nand UO_1120 (O_1120,N_8593,N_9434);
or UO_1121 (O_1121,N_9901,N_9071);
nand UO_1122 (O_1122,N_8472,N_9734);
and UO_1123 (O_1123,N_8166,N_8762);
nand UO_1124 (O_1124,N_8278,N_9815);
nor UO_1125 (O_1125,N_9243,N_9759);
nor UO_1126 (O_1126,N_9769,N_9833);
xnor UO_1127 (O_1127,N_9889,N_8236);
or UO_1128 (O_1128,N_9890,N_9023);
nor UO_1129 (O_1129,N_9565,N_9670);
and UO_1130 (O_1130,N_8344,N_8487);
and UO_1131 (O_1131,N_8624,N_9807);
nand UO_1132 (O_1132,N_9121,N_8926);
xnor UO_1133 (O_1133,N_9923,N_9621);
nor UO_1134 (O_1134,N_8492,N_8887);
and UO_1135 (O_1135,N_8550,N_9576);
and UO_1136 (O_1136,N_8491,N_9594);
or UO_1137 (O_1137,N_8976,N_9791);
nor UO_1138 (O_1138,N_8862,N_8839);
and UO_1139 (O_1139,N_9466,N_9060);
or UO_1140 (O_1140,N_8953,N_9366);
xnor UO_1141 (O_1141,N_8141,N_9000);
nor UO_1142 (O_1142,N_8213,N_8378);
and UO_1143 (O_1143,N_8894,N_8957);
and UO_1144 (O_1144,N_8449,N_9299);
nand UO_1145 (O_1145,N_9578,N_9504);
xor UO_1146 (O_1146,N_8834,N_9302);
and UO_1147 (O_1147,N_8737,N_8193);
nand UO_1148 (O_1148,N_9802,N_8762);
or UO_1149 (O_1149,N_9312,N_8953);
nor UO_1150 (O_1150,N_9250,N_8991);
and UO_1151 (O_1151,N_9196,N_8334);
nor UO_1152 (O_1152,N_8715,N_9586);
or UO_1153 (O_1153,N_8381,N_8785);
nand UO_1154 (O_1154,N_8473,N_8716);
and UO_1155 (O_1155,N_9062,N_8545);
and UO_1156 (O_1156,N_8114,N_9170);
or UO_1157 (O_1157,N_9223,N_9167);
or UO_1158 (O_1158,N_9588,N_8051);
nor UO_1159 (O_1159,N_8273,N_9001);
nor UO_1160 (O_1160,N_9305,N_8584);
nand UO_1161 (O_1161,N_8823,N_9973);
nand UO_1162 (O_1162,N_9200,N_8082);
xnor UO_1163 (O_1163,N_9357,N_9892);
nor UO_1164 (O_1164,N_9090,N_8085);
xnor UO_1165 (O_1165,N_8717,N_8612);
nand UO_1166 (O_1166,N_8307,N_9415);
or UO_1167 (O_1167,N_9545,N_8964);
and UO_1168 (O_1168,N_9122,N_8076);
or UO_1169 (O_1169,N_8107,N_8039);
nand UO_1170 (O_1170,N_8124,N_9201);
xnor UO_1171 (O_1171,N_9152,N_9219);
and UO_1172 (O_1172,N_8108,N_8811);
nand UO_1173 (O_1173,N_9176,N_9492);
nand UO_1174 (O_1174,N_9668,N_9717);
nor UO_1175 (O_1175,N_8961,N_8437);
nor UO_1176 (O_1176,N_8456,N_9921);
nor UO_1177 (O_1177,N_8735,N_9508);
xor UO_1178 (O_1178,N_8995,N_8585);
nor UO_1179 (O_1179,N_9520,N_8793);
nor UO_1180 (O_1180,N_8291,N_9180);
nor UO_1181 (O_1181,N_8059,N_9272);
and UO_1182 (O_1182,N_8269,N_9521);
nor UO_1183 (O_1183,N_9748,N_9149);
nor UO_1184 (O_1184,N_9695,N_8730);
nand UO_1185 (O_1185,N_8399,N_9127);
and UO_1186 (O_1186,N_8317,N_8026);
xor UO_1187 (O_1187,N_8670,N_9940);
or UO_1188 (O_1188,N_8108,N_9897);
or UO_1189 (O_1189,N_8576,N_8407);
nor UO_1190 (O_1190,N_9679,N_9727);
xnor UO_1191 (O_1191,N_8732,N_9851);
nand UO_1192 (O_1192,N_9583,N_8757);
xnor UO_1193 (O_1193,N_8638,N_8717);
nor UO_1194 (O_1194,N_9240,N_9856);
or UO_1195 (O_1195,N_8824,N_8079);
nand UO_1196 (O_1196,N_9251,N_8600);
nand UO_1197 (O_1197,N_9053,N_8147);
nor UO_1198 (O_1198,N_9872,N_9224);
nand UO_1199 (O_1199,N_8520,N_8178);
nand UO_1200 (O_1200,N_8549,N_8093);
and UO_1201 (O_1201,N_8443,N_9220);
nor UO_1202 (O_1202,N_9900,N_8086);
and UO_1203 (O_1203,N_8015,N_8657);
nand UO_1204 (O_1204,N_8443,N_8403);
nor UO_1205 (O_1205,N_8380,N_9855);
nand UO_1206 (O_1206,N_9841,N_8266);
nor UO_1207 (O_1207,N_8855,N_8256);
or UO_1208 (O_1208,N_9110,N_8251);
and UO_1209 (O_1209,N_8117,N_8924);
nor UO_1210 (O_1210,N_8712,N_8718);
nor UO_1211 (O_1211,N_9953,N_8891);
nor UO_1212 (O_1212,N_9029,N_9762);
nor UO_1213 (O_1213,N_9401,N_9410);
nor UO_1214 (O_1214,N_9338,N_9573);
or UO_1215 (O_1215,N_8168,N_9505);
nand UO_1216 (O_1216,N_8774,N_9337);
nor UO_1217 (O_1217,N_9092,N_9561);
or UO_1218 (O_1218,N_8375,N_8404);
or UO_1219 (O_1219,N_9585,N_8554);
nor UO_1220 (O_1220,N_9203,N_8584);
nand UO_1221 (O_1221,N_8380,N_8668);
and UO_1222 (O_1222,N_8720,N_9265);
nor UO_1223 (O_1223,N_8814,N_9889);
nor UO_1224 (O_1224,N_8855,N_9966);
or UO_1225 (O_1225,N_8153,N_9233);
or UO_1226 (O_1226,N_9043,N_8031);
xor UO_1227 (O_1227,N_9478,N_9355);
and UO_1228 (O_1228,N_8913,N_8924);
xnor UO_1229 (O_1229,N_8408,N_8073);
or UO_1230 (O_1230,N_8791,N_9596);
and UO_1231 (O_1231,N_8649,N_9296);
or UO_1232 (O_1232,N_9556,N_9425);
or UO_1233 (O_1233,N_9414,N_9699);
xor UO_1234 (O_1234,N_8347,N_9746);
nand UO_1235 (O_1235,N_9300,N_8128);
nor UO_1236 (O_1236,N_8095,N_8961);
nor UO_1237 (O_1237,N_9082,N_9836);
nor UO_1238 (O_1238,N_8210,N_9952);
nor UO_1239 (O_1239,N_8765,N_9465);
nor UO_1240 (O_1240,N_8308,N_8204);
nand UO_1241 (O_1241,N_8520,N_8592);
or UO_1242 (O_1242,N_9710,N_9527);
nor UO_1243 (O_1243,N_8120,N_9437);
nor UO_1244 (O_1244,N_8721,N_9027);
nor UO_1245 (O_1245,N_9528,N_9742);
and UO_1246 (O_1246,N_8935,N_8357);
or UO_1247 (O_1247,N_8216,N_8928);
and UO_1248 (O_1248,N_9140,N_8209);
nor UO_1249 (O_1249,N_8629,N_9240);
or UO_1250 (O_1250,N_8594,N_8564);
and UO_1251 (O_1251,N_8029,N_8112);
or UO_1252 (O_1252,N_8385,N_9202);
or UO_1253 (O_1253,N_8565,N_9045);
or UO_1254 (O_1254,N_8141,N_8718);
and UO_1255 (O_1255,N_9721,N_9535);
or UO_1256 (O_1256,N_9580,N_9824);
and UO_1257 (O_1257,N_8467,N_8172);
and UO_1258 (O_1258,N_9937,N_8006);
or UO_1259 (O_1259,N_9192,N_8396);
nor UO_1260 (O_1260,N_8788,N_9957);
or UO_1261 (O_1261,N_9405,N_8904);
and UO_1262 (O_1262,N_9734,N_8894);
and UO_1263 (O_1263,N_9921,N_8670);
nand UO_1264 (O_1264,N_8892,N_8589);
nor UO_1265 (O_1265,N_8992,N_8068);
or UO_1266 (O_1266,N_8307,N_9329);
nor UO_1267 (O_1267,N_8396,N_8857);
nor UO_1268 (O_1268,N_8694,N_8918);
nor UO_1269 (O_1269,N_9521,N_9047);
or UO_1270 (O_1270,N_9372,N_9874);
xor UO_1271 (O_1271,N_9989,N_9924);
nand UO_1272 (O_1272,N_9202,N_9561);
nor UO_1273 (O_1273,N_8894,N_9551);
nor UO_1274 (O_1274,N_8664,N_8452);
xnor UO_1275 (O_1275,N_9945,N_9381);
nand UO_1276 (O_1276,N_8634,N_9560);
nand UO_1277 (O_1277,N_9312,N_9569);
and UO_1278 (O_1278,N_8294,N_9548);
or UO_1279 (O_1279,N_8011,N_9885);
nand UO_1280 (O_1280,N_9737,N_9571);
xor UO_1281 (O_1281,N_9010,N_8779);
or UO_1282 (O_1282,N_8403,N_8259);
xnor UO_1283 (O_1283,N_9070,N_8623);
or UO_1284 (O_1284,N_8180,N_9657);
nor UO_1285 (O_1285,N_8791,N_8981);
and UO_1286 (O_1286,N_9874,N_8424);
or UO_1287 (O_1287,N_8851,N_9657);
xnor UO_1288 (O_1288,N_8366,N_9368);
nor UO_1289 (O_1289,N_8805,N_8006);
nand UO_1290 (O_1290,N_8396,N_8210);
nor UO_1291 (O_1291,N_8602,N_9947);
and UO_1292 (O_1292,N_8578,N_9191);
nand UO_1293 (O_1293,N_8220,N_8787);
nor UO_1294 (O_1294,N_8172,N_9055);
or UO_1295 (O_1295,N_8492,N_8786);
and UO_1296 (O_1296,N_9818,N_8592);
nand UO_1297 (O_1297,N_9296,N_9750);
or UO_1298 (O_1298,N_9186,N_8935);
or UO_1299 (O_1299,N_9467,N_8949);
or UO_1300 (O_1300,N_9473,N_8025);
nand UO_1301 (O_1301,N_9238,N_9810);
or UO_1302 (O_1302,N_9707,N_9098);
nor UO_1303 (O_1303,N_8535,N_9221);
nor UO_1304 (O_1304,N_8535,N_9020);
nor UO_1305 (O_1305,N_8261,N_8696);
nand UO_1306 (O_1306,N_8901,N_9883);
and UO_1307 (O_1307,N_9519,N_8731);
nor UO_1308 (O_1308,N_9181,N_9403);
nor UO_1309 (O_1309,N_9082,N_9173);
nand UO_1310 (O_1310,N_9466,N_8461);
nor UO_1311 (O_1311,N_8597,N_9740);
nand UO_1312 (O_1312,N_9141,N_9620);
and UO_1313 (O_1313,N_9223,N_8010);
nor UO_1314 (O_1314,N_9971,N_9820);
and UO_1315 (O_1315,N_8245,N_8643);
and UO_1316 (O_1316,N_8181,N_9097);
and UO_1317 (O_1317,N_9346,N_9618);
nand UO_1318 (O_1318,N_8487,N_8829);
nor UO_1319 (O_1319,N_9021,N_8298);
and UO_1320 (O_1320,N_8841,N_8597);
or UO_1321 (O_1321,N_8035,N_8666);
and UO_1322 (O_1322,N_8508,N_9114);
and UO_1323 (O_1323,N_9008,N_9213);
nor UO_1324 (O_1324,N_9151,N_9494);
and UO_1325 (O_1325,N_8391,N_9768);
or UO_1326 (O_1326,N_8495,N_9634);
and UO_1327 (O_1327,N_8371,N_8729);
or UO_1328 (O_1328,N_9978,N_8607);
and UO_1329 (O_1329,N_9603,N_8540);
nand UO_1330 (O_1330,N_8612,N_9618);
and UO_1331 (O_1331,N_8794,N_9560);
and UO_1332 (O_1332,N_9642,N_8808);
or UO_1333 (O_1333,N_9916,N_9719);
and UO_1334 (O_1334,N_9010,N_8499);
xnor UO_1335 (O_1335,N_8070,N_8633);
nand UO_1336 (O_1336,N_8348,N_9988);
nand UO_1337 (O_1337,N_9451,N_8461);
or UO_1338 (O_1338,N_9484,N_8737);
xor UO_1339 (O_1339,N_8643,N_8131);
nand UO_1340 (O_1340,N_8599,N_8986);
xnor UO_1341 (O_1341,N_8299,N_8613);
and UO_1342 (O_1342,N_8144,N_8080);
and UO_1343 (O_1343,N_8444,N_9720);
nor UO_1344 (O_1344,N_9991,N_9407);
nand UO_1345 (O_1345,N_9815,N_9159);
nor UO_1346 (O_1346,N_8972,N_9787);
nand UO_1347 (O_1347,N_9309,N_9596);
and UO_1348 (O_1348,N_9088,N_9525);
nand UO_1349 (O_1349,N_9866,N_8057);
or UO_1350 (O_1350,N_8860,N_9818);
nand UO_1351 (O_1351,N_8144,N_9065);
xor UO_1352 (O_1352,N_9531,N_8601);
and UO_1353 (O_1353,N_9585,N_8423);
nor UO_1354 (O_1354,N_8737,N_9310);
and UO_1355 (O_1355,N_9707,N_8078);
and UO_1356 (O_1356,N_9409,N_8783);
or UO_1357 (O_1357,N_9593,N_8089);
or UO_1358 (O_1358,N_8007,N_9818);
and UO_1359 (O_1359,N_9945,N_8330);
and UO_1360 (O_1360,N_8153,N_9346);
nor UO_1361 (O_1361,N_9503,N_9709);
and UO_1362 (O_1362,N_8284,N_8656);
or UO_1363 (O_1363,N_8928,N_8823);
nor UO_1364 (O_1364,N_9845,N_8628);
and UO_1365 (O_1365,N_9925,N_9194);
and UO_1366 (O_1366,N_9971,N_9337);
nand UO_1367 (O_1367,N_8901,N_8884);
or UO_1368 (O_1368,N_8630,N_9566);
and UO_1369 (O_1369,N_9567,N_9983);
and UO_1370 (O_1370,N_9282,N_8887);
and UO_1371 (O_1371,N_9712,N_9324);
xor UO_1372 (O_1372,N_8889,N_8696);
and UO_1373 (O_1373,N_8673,N_8688);
nand UO_1374 (O_1374,N_8815,N_8200);
or UO_1375 (O_1375,N_8530,N_8490);
xnor UO_1376 (O_1376,N_9689,N_9385);
nor UO_1377 (O_1377,N_9263,N_9262);
nor UO_1378 (O_1378,N_9966,N_9543);
nand UO_1379 (O_1379,N_9375,N_8800);
nor UO_1380 (O_1380,N_8745,N_8842);
nand UO_1381 (O_1381,N_8954,N_9196);
nor UO_1382 (O_1382,N_8094,N_9190);
nor UO_1383 (O_1383,N_9157,N_8310);
or UO_1384 (O_1384,N_9548,N_9200);
and UO_1385 (O_1385,N_9429,N_8010);
or UO_1386 (O_1386,N_9253,N_9456);
or UO_1387 (O_1387,N_8864,N_9286);
or UO_1388 (O_1388,N_8754,N_9026);
nor UO_1389 (O_1389,N_9779,N_9876);
and UO_1390 (O_1390,N_8491,N_8464);
nand UO_1391 (O_1391,N_8031,N_9999);
nand UO_1392 (O_1392,N_8585,N_9138);
or UO_1393 (O_1393,N_9231,N_9538);
nand UO_1394 (O_1394,N_9822,N_9880);
xnor UO_1395 (O_1395,N_8501,N_9731);
nand UO_1396 (O_1396,N_8844,N_8539);
and UO_1397 (O_1397,N_9700,N_8000);
and UO_1398 (O_1398,N_9047,N_8359);
xnor UO_1399 (O_1399,N_8042,N_8796);
nand UO_1400 (O_1400,N_9245,N_9796);
xor UO_1401 (O_1401,N_8510,N_8458);
nor UO_1402 (O_1402,N_9737,N_8282);
nor UO_1403 (O_1403,N_8466,N_8120);
and UO_1404 (O_1404,N_8024,N_8537);
or UO_1405 (O_1405,N_8511,N_9586);
xor UO_1406 (O_1406,N_8619,N_9940);
or UO_1407 (O_1407,N_8268,N_9235);
or UO_1408 (O_1408,N_8490,N_9808);
or UO_1409 (O_1409,N_8146,N_8013);
nand UO_1410 (O_1410,N_8160,N_9578);
nor UO_1411 (O_1411,N_9601,N_9008);
nor UO_1412 (O_1412,N_8274,N_8461);
or UO_1413 (O_1413,N_9304,N_8503);
nor UO_1414 (O_1414,N_9585,N_8446);
xor UO_1415 (O_1415,N_9379,N_9039);
and UO_1416 (O_1416,N_9015,N_9114);
or UO_1417 (O_1417,N_9879,N_8000);
and UO_1418 (O_1418,N_9028,N_8423);
nor UO_1419 (O_1419,N_8845,N_8307);
nand UO_1420 (O_1420,N_9632,N_9635);
and UO_1421 (O_1421,N_8398,N_9856);
or UO_1422 (O_1422,N_8507,N_8113);
nand UO_1423 (O_1423,N_8127,N_8640);
or UO_1424 (O_1424,N_9584,N_9837);
or UO_1425 (O_1425,N_8516,N_9943);
nand UO_1426 (O_1426,N_9544,N_9187);
or UO_1427 (O_1427,N_9485,N_9190);
and UO_1428 (O_1428,N_8089,N_8959);
nor UO_1429 (O_1429,N_9112,N_9995);
and UO_1430 (O_1430,N_9330,N_9902);
or UO_1431 (O_1431,N_9884,N_9125);
nor UO_1432 (O_1432,N_9053,N_8978);
or UO_1433 (O_1433,N_8807,N_9713);
or UO_1434 (O_1434,N_9900,N_9343);
nand UO_1435 (O_1435,N_9695,N_9082);
or UO_1436 (O_1436,N_8687,N_9825);
or UO_1437 (O_1437,N_8889,N_9886);
and UO_1438 (O_1438,N_9031,N_9306);
nand UO_1439 (O_1439,N_8614,N_8356);
or UO_1440 (O_1440,N_8546,N_9233);
or UO_1441 (O_1441,N_8725,N_9491);
or UO_1442 (O_1442,N_9766,N_8324);
or UO_1443 (O_1443,N_9310,N_8975);
xor UO_1444 (O_1444,N_8858,N_9886);
and UO_1445 (O_1445,N_8663,N_8764);
nor UO_1446 (O_1446,N_9361,N_9451);
or UO_1447 (O_1447,N_9164,N_9140);
nand UO_1448 (O_1448,N_9752,N_8555);
or UO_1449 (O_1449,N_9794,N_8065);
or UO_1450 (O_1450,N_9515,N_8913);
or UO_1451 (O_1451,N_8330,N_9883);
nor UO_1452 (O_1452,N_8209,N_9237);
nand UO_1453 (O_1453,N_8357,N_9063);
or UO_1454 (O_1454,N_9458,N_8398);
and UO_1455 (O_1455,N_9673,N_9084);
or UO_1456 (O_1456,N_8030,N_8353);
nor UO_1457 (O_1457,N_9154,N_9218);
or UO_1458 (O_1458,N_9863,N_9541);
xor UO_1459 (O_1459,N_9861,N_9103);
or UO_1460 (O_1460,N_8554,N_8182);
nand UO_1461 (O_1461,N_8690,N_9101);
or UO_1462 (O_1462,N_8696,N_8320);
and UO_1463 (O_1463,N_8955,N_9588);
nor UO_1464 (O_1464,N_8090,N_8198);
and UO_1465 (O_1465,N_8726,N_9461);
nand UO_1466 (O_1466,N_8754,N_8612);
or UO_1467 (O_1467,N_8424,N_8855);
nand UO_1468 (O_1468,N_9371,N_9647);
or UO_1469 (O_1469,N_9976,N_8135);
nor UO_1470 (O_1470,N_8427,N_9220);
nand UO_1471 (O_1471,N_8203,N_9426);
nand UO_1472 (O_1472,N_9840,N_8632);
and UO_1473 (O_1473,N_9132,N_9979);
and UO_1474 (O_1474,N_9368,N_8903);
nand UO_1475 (O_1475,N_8753,N_9040);
nor UO_1476 (O_1476,N_8900,N_9342);
nand UO_1477 (O_1477,N_8379,N_9220);
nor UO_1478 (O_1478,N_9531,N_8835);
nor UO_1479 (O_1479,N_8397,N_8234);
nor UO_1480 (O_1480,N_8764,N_8305);
and UO_1481 (O_1481,N_8518,N_8047);
nand UO_1482 (O_1482,N_9530,N_9267);
nand UO_1483 (O_1483,N_8569,N_9910);
or UO_1484 (O_1484,N_8354,N_8786);
nor UO_1485 (O_1485,N_8830,N_8033);
nor UO_1486 (O_1486,N_9890,N_9595);
nor UO_1487 (O_1487,N_9778,N_8634);
or UO_1488 (O_1488,N_8405,N_9798);
or UO_1489 (O_1489,N_8470,N_9670);
nand UO_1490 (O_1490,N_9687,N_9509);
and UO_1491 (O_1491,N_8171,N_8665);
nand UO_1492 (O_1492,N_8366,N_9456);
nor UO_1493 (O_1493,N_8757,N_8258);
and UO_1494 (O_1494,N_9272,N_9397);
nand UO_1495 (O_1495,N_8390,N_9221);
nand UO_1496 (O_1496,N_8321,N_8853);
or UO_1497 (O_1497,N_8165,N_8874);
or UO_1498 (O_1498,N_8274,N_9627);
or UO_1499 (O_1499,N_8580,N_8285);
endmodule