module basic_750_5000_1000_2_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2501,N_2502,N_2503,N_2504,N_2506,N_2507,N_2508,N_2510,N_2511,N_2513,N_2514,N_2515,N_2516,N_2518,N_2519,N_2521,N_2522,N_2523,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2538,N_2539,N_2540,N_2541,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2551,N_2552,N_2553,N_2554,N_2555,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2567,N_2568,N_2569,N_2570,N_2572,N_2574,N_2575,N_2576,N_2577,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2595,N_2597,N_2598,N_2599,N_2601,N_2602,N_2604,N_2605,N_2606,N_2607,N_2609,N_2610,N_2612,N_2613,N_2614,N_2616,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2627,N_2628,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2643,N_2644,N_2645,N_2647,N_2648,N_2649,N_2652,N_2653,N_2654,N_2655,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2665,N_2666,N_2667,N_2669,N_2670,N_2671,N_2672,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2698,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2733,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2743,N_2745,N_2746,N_2748,N_2750,N_2751,N_2753,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2790,N_2791,N_2792,N_2793,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2802,N_2803,N_2804,N_2806,N_2808,N_2809,N_2810,N_2812,N_2813,N_2815,N_2816,N_2818,N_2821,N_2822,N_2823,N_2824,N_2825,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2865,N_2866,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2899,N_2900,N_2901,N_2902,N_2903,N_2905,N_2906,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2932,N_2934,N_2935,N_2936,N_2937,N_2938,N_2940,N_2941,N_2942,N_2943,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2963,N_2964,N_2965,N_2968,N_2969,N_2970,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2981,N_2982,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3023,N_3024,N_3026,N_3027,N_3028,N_3029,N_3030,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3049,N_3050,N_3053,N_3054,N_3055,N_3056,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3102,N_3103,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3115,N_3116,N_3119,N_3120,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3130,N_3131,N_3132,N_3133,N_3134,N_3136,N_3138,N_3139,N_3140,N_3141,N_3142,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3162,N_3164,N_3165,N_3166,N_3168,N_3170,N_3171,N_3172,N_3173,N_3174,N_3176,N_3177,N_3179,N_3180,N_3181,N_3183,N_3185,N_3186,N_3187,N_3188,N_3189,N_3191,N_3192,N_3193,N_3194,N_3195,N_3197,N_3198,N_3199,N_3201,N_3202,N_3204,N_3205,N_3207,N_3210,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3268,N_3270,N_3271,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3281,N_3282,N_3283,N_3284,N_3286,N_3287,N_3288,N_3289,N_3290,N_3292,N_3293,N_3294,N_3295,N_3297,N_3298,N_3300,N_3301,N_3303,N_3304,N_3305,N_3306,N_3307,N_3310,N_3311,N_3313,N_3314,N_3315,N_3316,N_3317,N_3319,N_3322,N_3323,N_3324,N_3328,N_3329,N_3330,N_3331,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3343,N_3344,N_3345,N_3346,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3365,N_3366,N_3367,N_3368,N_3369,N_3372,N_3373,N_3375,N_3376,N_3377,N_3379,N_3380,N_3382,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3403,N_3405,N_3406,N_3408,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3422,N_3424,N_3425,N_3426,N_3427,N_3428,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3441,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3468,N_3469,N_3470,N_3471,N_3473,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3487,N_3490,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3503,N_3504,N_3505,N_3506,N_3507,N_3509,N_3511,N_3513,N_3514,N_3515,N_3516,N_3518,N_3519,N_3520,N_3522,N_3523,N_3524,N_3525,N_3526,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3547,N_3548,N_3550,N_3551,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3576,N_3577,N_3579,N_3580,N_3581,N_3583,N_3584,N_3586,N_3587,N_3588,N_3589,N_3590,N_3592,N_3593,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3603,N_3604,N_3605,N_3606,N_3608,N_3610,N_3611,N_3612,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3632,N_3633,N_3634,N_3635,N_3636,N_3638,N_3639,N_3641,N_3643,N_3645,N_3646,N_3647,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3663,N_3664,N_3666,N_3667,N_3668,N_3669,N_3671,N_3672,N_3674,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3714,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3735,N_3736,N_3737,N_3739,N_3741,N_3742,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3752,N_3753,N_3754,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3764,N_3766,N_3767,N_3768,N_3769,N_3770,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3781,N_3782,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3793,N_3794,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3813,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3830,N_3831,N_3833,N_3834,N_3835,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3848,N_3849,N_3850,N_3852,N_3853,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3867,N_3868,N_3869,N_3870,N_3871,N_3873,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3894,N_3895,N_3897,N_3898,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3910,N_3911,N_3912,N_3913,N_3914,N_3916,N_3918,N_3919,N_3921,N_3923,N_3924,N_3925,N_3926,N_3928,N_3929,N_3931,N_3932,N_3933,N_3934,N_3936,N_3937,N_3938,N_3939,N_3940,N_3942,N_3944,N_3945,N_3946,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3957,N_3958,N_3959,N_3960,N_3962,N_3963,N_3964,N_3965,N_3966,N_3968,N_3969,N_3970,N_3976,N_3977,N_3978,N_3979,N_3982,N_3983,N_3984,N_3986,N_3987,N_3990,N_3991,N_3992,N_3993,N_3994,N_3996,N_3997,N_4000,N_4001,N_4002,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4011,N_4012,N_4013,N_4014,N_4017,N_4019,N_4020,N_4023,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4048,N_4049,N_4050,N_4051,N_4052,N_4055,N_4056,N_4057,N_4059,N_4061,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4079,N_4081,N_4083,N_4084,N_4085,N_4086,N_4087,N_4089,N_4091,N_4094,N_4095,N_4096,N_4097,N_4099,N_4100,N_4101,N_4103,N_4104,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4125,N_4126,N_4127,N_4128,N_4130,N_4132,N_4133,N_4134,N_4135,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4155,N_4156,N_4157,N_4158,N_4159,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4173,N_4174,N_4175,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4184,N_4186,N_4187,N_4189,N_4190,N_4191,N_4192,N_4193,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4220,N_4221,N_4222,N_4223,N_4225,N_4226,N_4228,N_4230,N_4231,N_4233,N_4234,N_4236,N_4237,N_4238,N_4241,N_4242,N_4246,N_4249,N_4251,N_4254,N_4255,N_4256,N_4257,N_4259,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4277,N_4278,N_4280,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4297,N_4299,N_4300,N_4301,N_4302,N_4303,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4314,N_4315,N_4316,N_4317,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4328,N_4329,N_4330,N_4332,N_4333,N_4334,N_4335,N_4337,N_4339,N_4340,N_4341,N_4343,N_4346,N_4347,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4363,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4394,N_4395,N_4396,N_4398,N_4399,N_4400,N_4402,N_4406,N_4408,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4417,N_4418,N_4420,N_4421,N_4422,N_4423,N_4424,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4436,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4453,N_4454,N_4455,N_4456,N_4457,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4496,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4506,N_4508,N_4509,N_4510,N_4511,N_4512,N_4514,N_4515,N_4519,N_4521,N_4522,N_4523,N_4524,N_4526,N_4527,N_4528,N_4530,N_4531,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4541,N_4542,N_4543,N_4544,N_4545,N_4548,N_4549,N_4551,N_4552,N_4553,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4602,N_4603,N_4604,N_4606,N_4607,N_4609,N_4610,N_4612,N_4614,N_4616,N_4617,N_4619,N_4620,N_4622,N_4623,N_4624,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4634,N_4636,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4659,N_4660,N_4661,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4693,N_4694,N_4696,N_4697,N_4699,N_4701,N_4702,N_4706,N_4707,N_4708,N_4710,N_4712,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4744,N_4745,N_4747,N_4749,N_4750,N_4751,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4773,N_4774,N_4775,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4790,N_4793,N_4794,N_4795,N_4796,N_4797,N_4800,N_4801,N_4803,N_4804,N_4805,N_4806,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4840,N_4841,N_4842,N_4844,N_4845,N_4846,N_4847,N_4848,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4860,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4875,N_4877,N_4879,N_4880,N_4882,N_4883,N_4884,N_4888,N_4889,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4927,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4938,N_4940,N_4941,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4997,N_4998;
nand U0 (N_0,In_692,In_544);
or U1 (N_1,In_353,In_284);
and U2 (N_2,In_177,In_426);
nand U3 (N_3,In_256,In_263);
nor U4 (N_4,In_142,In_86);
nand U5 (N_5,In_210,In_701);
nand U6 (N_6,In_209,In_718);
nor U7 (N_7,In_387,In_83);
or U8 (N_8,In_439,In_524);
nor U9 (N_9,In_190,In_447);
and U10 (N_10,In_286,In_516);
nand U11 (N_11,In_249,In_272);
or U12 (N_12,In_366,In_265);
nand U13 (N_13,In_116,In_258);
nor U14 (N_14,In_234,In_480);
nand U15 (N_15,In_499,In_505);
nand U16 (N_16,In_342,In_324);
nand U17 (N_17,In_181,In_160);
xor U18 (N_18,In_720,In_734);
nand U19 (N_19,In_625,In_332);
or U20 (N_20,In_185,In_397);
or U21 (N_21,In_440,In_235);
nor U22 (N_22,In_42,In_64);
and U23 (N_23,In_11,In_128);
or U24 (N_24,In_77,In_647);
nor U25 (N_25,In_50,In_436);
nor U26 (N_26,In_261,In_512);
nor U27 (N_27,In_129,In_489);
or U28 (N_28,In_56,In_451);
or U29 (N_29,In_427,In_333);
nand U30 (N_30,In_737,In_199);
nor U31 (N_31,In_291,In_595);
or U32 (N_32,In_541,In_111);
nand U33 (N_33,In_742,In_497);
nand U34 (N_34,In_279,In_58);
nor U35 (N_35,In_183,In_375);
and U36 (N_36,In_721,In_309);
or U37 (N_37,In_98,In_206);
or U38 (N_38,In_578,In_144);
nor U39 (N_39,In_556,In_457);
nor U40 (N_40,In_171,In_748);
nor U41 (N_41,In_507,In_93);
or U42 (N_42,In_695,In_669);
nor U43 (N_43,In_271,In_422);
nor U44 (N_44,In_255,In_450);
nand U45 (N_45,In_562,In_310);
and U46 (N_46,In_697,In_51);
nand U47 (N_47,In_322,In_545);
nor U48 (N_48,In_109,In_338);
xor U49 (N_49,In_400,In_317);
and U50 (N_50,In_722,In_155);
nor U51 (N_51,In_605,In_501);
nor U52 (N_52,In_285,In_574);
nand U53 (N_53,In_632,In_491);
nor U54 (N_54,In_303,In_84);
and U55 (N_55,In_604,In_319);
or U56 (N_56,In_301,In_461);
nor U57 (N_57,In_484,In_627);
and U58 (N_58,In_67,In_577);
nor U59 (N_59,In_148,In_719);
nor U60 (N_60,In_386,In_33);
or U61 (N_61,In_736,In_389);
nor U62 (N_62,In_471,In_334);
nand U63 (N_63,In_442,In_66);
and U64 (N_64,In_108,In_671);
and U65 (N_65,In_602,In_292);
or U66 (N_66,In_2,In_470);
nand U67 (N_67,In_394,In_415);
nand U68 (N_68,In_641,In_483);
and U69 (N_69,In_127,In_566);
xnor U70 (N_70,In_438,In_664);
nand U71 (N_71,In_479,In_268);
nor U72 (N_72,In_216,In_132);
and U73 (N_73,In_162,In_4);
nand U74 (N_74,In_462,In_367);
nor U75 (N_75,In_237,In_28);
or U76 (N_76,In_619,In_223);
nand U77 (N_77,In_659,In_633);
nor U78 (N_78,In_746,In_145);
nand U79 (N_79,In_196,In_328);
and U80 (N_80,In_147,In_246);
or U81 (N_81,In_20,In_260);
nor U82 (N_82,In_276,In_563);
nand U83 (N_83,In_321,In_494);
nor U84 (N_84,In_110,In_75);
or U85 (N_85,In_526,In_548);
nor U86 (N_86,In_730,In_599);
or U87 (N_87,In_305,In_165);
nand U88 (N_88,In_363,In_735);
and U89 (N_89,In_38,In_421);
nand U90 (N_90,In_112,In_26);
nor U91 (N_91,In_60,In_296);
nor U92 (N_92,In_537,In_682);
and U93 (N_93,In_732,In_115);
or U94 (N_94,In_253,In_161);
or U95 (N_95,In_226,In_652);
or U96 (N_96,In_531,In_738);
or U97 (N_97,In_404,In_335);
nor U98 (N_98,In_76,In_217);
and U99 (N_99,In_549,In_481);
nor U100 (N_100,In_673,In_374);
nor U101 (N_101,In_337,In_509);
nand U102 (N_102,In_178,In_449);
or U103 (N_103,In_488,In_413);
nor U104 (N_104,In_74,In_472);
nor U105 (N_105,In_740,In_518);
nand U106 (N_106,In_355,In_612);
and U107 (N_107,In_248,In_198);
nor U108 (N_108,In_368,In_267);
nor U109 (N_109,In_243,In_675);
and U110 (N_110,In_616,In_113);
nand U111 (N_111,In_684,In_159);
or U112 (N_112,In_495,In_350);
xor U113 (N_113,In_238,In_716);
or U114 (N_114,In_24,In_608);
nor U115 (N_115,In_666,In_559);
and U116 (N_116,In_430,In_141);
nand U117 (N_117,In_362,In_583);
nor U118 (N_118,In_358,In_107);
or U119 (N_119,In_14,In_496);
and U120 (N_120,In_406,In_204);
nand U121 (N_121,In_273,In_62);
nand U122 (N_122,In_661,In_48);
xor U123 (N_123,In_278,In_408);
or U124 (N_124,In_651,In_525);
nor U125 (N_125,In_90,In_607);
or U126 (N_126,In_345,In_711);
nand U127 (N_127,In_19,In_176);
nand U128 (N_128,In_52,In_281);
nor U129 (N_129,In_7,In_553);
nor U130 (N_130,In_139,In_274);
and U131 (N_131,In_739,In_468);
nor U132 (N_132,In_392,In_679);
nor U133 (N_133,In_289,In_411);
and U134 (N_134,In_244,In_254);
nand U135 (N_135,In_596,In_663);
nand U136 (N_136,In_320,In_713);
or U137 (N_137,In_687,In_435);
and U138 (N_138,In_224,In_54);
nand U139 (N_139,In_463,In_382);
nand U140 (N_140,In_402,In_403);
or U141 (N_141,In_569,In_710);
nand U142 (N_142,In_469,In_529);
nand U143 (N_143,In_519,In_15);
nor U144 (N_144,In_433,In_175);
nand U145 (N_145,In_207,In_43);
and U146 (N_146,In_61,In_347);
and U147 (N_147,In_242,In_180);
and U148 (N_148,In_114,In_360);
nor U149 (N_149,In_637,In_580);
nor U150 (N_150,In_87,In_493);
xnor U151 (N_151,In_466,In_448);
nor U152 (N_152,In_137,In_588);
or U153 (N_153,In_589,In_726);
nand U154 (N_154,In_700,In_476);
nand U155 (N_155,In_94,In_47);
and U156 (N_156,In_485,In_197);
or U157 (N_157,In_568,In_146);
nor U158 (N_158,In_508,In_65);
and U159 (N_159,In_552,In_629);
and U160 (N_160,In_646,In_655);
or U161 (N_161,In_89,In_540);
nor U162 (N_162,In_245,In_369);
nor U163 (N_163,In_203,In_228);
and U164 (N_164,In_189,In_662);
and U165 (N_165,In_564,In_225);
or U166 (N_166,In_151,In_68);
or U167 (N_167,In_215,In_167);
nor U168 (N_168,In_704,In_150);
nand U169 (N_169,In_723,In_365);
or U170 (N_170,In_391,In_288);
or U171 (N_171,In_455,In_354);
or U172 (N_172,In_174,In_229);
or U173 (N_173,In_192,In_85);
or U174 (N_174,In_572,In_538);
nor U175 (N_175,In_70,In_379);
and U176 (N_176,In_714,In_573);
nand U177 (N_177,In_80,In_584);
and U178 (N_178,In_547,In_743);
xnor U179 (N_179,In_688,In_314);
nand U180 (N_180,In_282,In_25);
nand U181 (N_181,In_221,In_532);
or U182 (N_182,In_346,In_280);
and U183 (N_183,In_533,In_393);
nor U184 (N_184,In_46,In_418);
nand U185 (N_185,In_414,In_100);
or U186 (N_186,In_377,In_709);
nand U187 (N_187,In_517,In_97);
or U188 (N_188,In_638,In_21);
xor U189 (N_189,In_315,In_49);
nand U190 (N_190,In_744,In_262);
or U191 (N_191,In_428,In_269);
or U192 (N_192,In_95,In_172);
or U193 (N_193,In_120,In_364);
and U194 (N_194,In_741,In_648);
nor U195 (N_195,In_313,In_191);
nand U196 (N_196,In_498,In_745);
and U197 (N_197,In_571,In_103);
and U198 (N_198,In_560,In_611);
and U199 (N_199,In_45,In_643);
nor U200 (N_200,In_41,In_401);
nor U201 (N_201,In_478,In_445);
nor U202 (N_202,In_521,In_446);
nand U203 (N_203,In_264,In_644);
and U204 (N_204,In_130,In_444);
and U205 (N_205,In_339,In_318);
nand U206 (N_206,In_640,In_570);
and U207 (N_207,In_283,In_515);
and U208 (N_208,In_654,In_373);
nor U209 (N_209,In_536,In_678);
nor U210 (N_210,In_676,In_708);
nor U211 (N_211,In_606,In_691);
nand U212 (N_212,In_69,In_157);
nand U213 (N_213,In_205,In_376);
or U214 (N_214,In_169,In_307);
and U215 (N_215,In_561,In_555);
nand U216 (N_216,In_92,In_399);
and U217 (N_217,In_681,In_121);
or U218 (N_218,In_8,In_13);
and U219 (N_219,In_639,In_17);
nand U220 (N_220,In_275,In_585);
nand U221 (N_221,In_81,In_405);
nor U222 (N_222,In_236,In_630);
or U223 (N_223,In_166,In_635);
or U224 (N_224,In_591,In_696);
or U225 (N_225,In_452,In_618);
nand U226 (N_226,In_118,In_59);
xor U227 (N_227,In_441,In_617);
nand U228 (N_228,In_657,In_717);
xnor U229 (N_229,In_523,In_214);
and U230 (N_230,In_300,In_194);
and U231 (N_231,In_326,In_417);
and U232 (N_232,In_308,In_133);
and U233 (N_233,In_163,In_384);
or U234 (N_234,In_614,In_725);
or U235 (N_235,In_232,In_590);
or U236 (N_236,In_551,In_443);
nor U237 (N_237,In_705,In_672);
and U238 (N_238,In_27,In_135);
or U239 (N_239,In_188,In_527);
and U240 (N_240,In_201,In_327);
nand U241 (N_241,In_82,In_312);
or U242 (N_242,In_34,In_513);
nor U243 (N_243,In_610,In_252);
nor U244 (N_244,In_336,In_23);
xor U245 (N_245,In_727,In_567);
nand U246 (N_246,In_32,In_410);
nand U247 (N_247,In_550,In_510);
or U248 (N_248,In_212,In_636);
nor U249 (N_249,In_173,In_409);
or U250 (N_250,In_259,In_156);
or U251 (N_251,In_143,In_88);
and U252 (N_252,In_434,In_728);
and U253 (N_253,In_656,In_359);
or U254 (N_254,In_306,In_693);
nand U255 (N_255,In_594,In_477);
nor U256 (N_256,In_371,In_558);
nand U257 (N_257,In_357,In_153);
nand U258 (N_258,In_431,In_348);
nand U259 (N_259,In_294,In_395);
nand U260 (N_260,In_603,In_105);
or U261 (N_261,In_35,In_323);
or U262 (N_262,In_168,In_658);
and U263 (N_263,In_707,In_241);
and U264 (N_264,In_474,In_240);
nor U265 (N_265,In_609,In_706);
nor U266 (N_266,In_535,In_304);
nor U267 (N_267,In_44,In_287);
or U268 (N_268,In_557,In_715);
or U269 (N_269,In_668,In_257);
or U270 (N_270,In_615,In_486);
nand U271 (N_271,In_425,In_601);
and U272 (N_272,In_195,In_372);
or U273 (N_273,In_125,In_220);
nand U274 (N_274,In_208,In_520);
or U275 (N_275,In_0,In_134);
nor U276 (N_276,In_660,In_482);
nor U277 (N_277,In_329,In_747);
or U278 (N_278,In_534,In_302);
or U279 (N_279,In_247,In_233);
xnor U280 (N_280,In_119,In_10);
and U281 (N_281,In_502,In_492);
or U282 (N_282,In_543,In_597);
nand U283 (N_283,In_613,In_352);
and U284 (N_284,In_152,In_295);
nand U285 (N_285,In_218,In_124);
or U286 (N_286,In_40,In_749);
and U287 (N_287,In_412,In_230);
nor U288 (N_288,In_12,In_419);
and U289 (N_289,In_634,In_398);
or U290 (N_290,In_138,In_653);
or U291 (N_291,In_645,In_164);
or U292 (N_292,In_624,In_702);
or U293 (N_293,In_3,In_1);
nand U294 (N_294,In_349,In_79);
and U295 (N_295,In_102,In_378);
nor U296 (N_296,In_9,In_187);
and U297 (N_297,In_694,In_642);
nor U298 (N_298,In_733,In_293);
nand U299 (N_299,In_53,In_424);
nor U300 (N_300,In_490,In_351);
nor U301 (N_301,In_622,In_16);
nor U302 (N_302,In_674,In_123);
or U303 (N_303,In_628,In_385);
and U304 (N_304,In_454,In_649);
and U305 (N_305,In_453,In_670);
and U306 (N_306,In_182,In_202);
or U307 (N_307,In_677,In_731);
nor U308 (N_308,In_689,In_222);
nand U309 (N_309,In_72,In_343);
nor U310 (N_310,In_6,In_131);
nand U311 (N_311,In_325,In_460);
and U312 (N_312,In_542,In_703);
and U313 (N_313,In_511,In_73);
nor U314 (N_314,In_620,In_341);
or U315 (N_315,In_390,In_37);
nand U316 (N_316,In_231,In_227);
and U317 (N_317,In_311,In_593);
or U318 (N_318,In_55,In_250);
and U319 (N_319,In_546,In_184);
nor U320 (N_320,In_437,In_154);
nor U321 (N_321,In_429,In_600);
nand U322 (N_322,In_5,In_140);
nor U323 (N_323,In_631,In_299);
nor U324 (N_324,In_39,In_370);
nand U325 (N_325,In_104,In_239);
or U326 (N_326,In_298,In_487);
nor U327 (N_327,In_514,In_330);
and U328 (N_328,In_686,In_396);
or U329 (N_329,In_456,In_465);
or U330 (N_330,In_581,In_500);
or U331 (N_331,In_626,In_504);
or U332 (N_332,In_586,In_667);
nor U333 (N_333,In_106,In_122);
or U334 (N_334,In_136,In_213);
xnor U335 (N_335,In_71,In_598);
nand U336 (N_336,In_416,In_149);
nand U337 (N_337,In_356,In_316);
and U338 (N_338,In_78,In_592);
or U339 (N_339,In_18,In_29);
and U340 (N_340,In_698,In_63);
or U341 (N_341,In_587,In_565);
nand U342 (N_342,In_530,In_712);
nor U343 (N_343,In_36,In_623);
nor U344 (N_344,In_270,In_650);
and U345 (N_345,In_528,In_458);
nor U346 (N_346,In_117,In_729);
nand U347 (N_347,In_724,In_576);
nand U348 (N_348,In_383,In_22);
or U349 (N_349,In_554,In_432);
or U350 (N_350,In_388,In_340);
or U351 (N_351,In_193,In_331);
nand U352 (N_352,In_158,In_251);
nand U353 (N_353,In_683,In_91);
and U354 (N_354,In_96,In_179);
nand U355 (N_355,In_361,In_30);
nor U356 (N_356,In_503,In_665);
nand U357 (N_357,In_475,In_467);
nor U358 (N_358,In_579,In_200);
nand U359 (N_359,In_699,In_266);
nor U360 (N_360,In_186,In_506);
or U361 (N_361,In_621,In_277);
or U362 (N_362,In_99,In_459);
or U363 (N_363,In_473,In_582);
nor U364 (N_364,In_539,In_575);
nor U365 (N_365,In_381,In_57);
nor U366 (N_366,In_126,In_380);
and U367 (N_367,In_464,In_101);
and U368 (N_368,In_211,In_31);
and U369 (N_369,In_344,In_423);
nor U370 (N_370,In_685,In_297);
or U371 (N_371,In_290,In_170);
nand U372 (N_372,In_407,In_420);
nand U373 (N_373,In_522,In_690);
or U374 (N_374,In_680,In_219);
or U375 (N_375,In_435,In_160);
nand U376 (N_376,In_317,In_47);
and U377 (N_377,In_51,In_648);
or U378 (N_378,In_323,In_368);
nor U379 (N_379,In_615,In_60);
nor U380 (N_380,In_244,In_720);
nor U381 (N_381,In_462,In_591);
and U382 (N_382,In_276,In_181);
and U383 (N_383,In_286,In_108);
or U384 (N_384,In_254,In_286);
and U385 (N_385,In_93,In_417);
nand U386 (N_386,In_416,In_684);
nand U387 (N_387,In_236,In_365);
and U388 (N_388,In_655,In_501);
nor U389 (N_389,In_72,In_646);
nor U390 (N_390,In_94,In_602);
or U391 (N_391,In_543,In_477);
nor U392 (N_392,In_137,In_591);
and U393 (N_393,In_395,In_71);
nand U394 (N_394,In_529,In_250);
nand U395 (N_395,In_126,In_385);
and U396 (N_396,In_676,In_522);
and U397 (N_397,In_713,In_201);
or U398 (N_398,In_626,In_11);
nand U399 (N_399,In_729,In_626);
nor U400 (N_400,In_495,In_86);
and U401 (N_401,In_396,In_570);
nor U402 (N_402,In_411,In_149);
or U403 (N_403,In_245,In_227);
nor U404 (N_404,In_589,In_445);
nand U405 (N_405,In_112,In_440);
and U406 (N_406,In_27,In_401);
or U407 (N_407,In_475,In_555);
nand U408 (N_408,In_480,In_648);
nor U409 (N_409,In_134,In_57);
nor U410 (N_410,In_745,In_270);
nor U411 (N_411,In_363,In_323);
or U412 (N_412,In_555,In_143);
xnor U413 (N_413,In_393,In_744);
nor U414 (N_414,In_521,In_714);
or U415 (N_415,In_613,In_367);
nand U416 (N_416,In_478,In_291);
and U417 (N_417,In_522,In_536);
or U418 (N_418,In_376,In_186);
nand U419 (N_419,In_10,In_197);
xnor U420 (N_420,In_60,In_77);
nand U421 (N_421,In_169,In_69);
or U422 (N_422,In_644,In_299);
or U423 (N_423,In_302,In_351);
nor U424 (N_424,In_625,In_456);
or U425 (N_425,In_255,In_456);
nand U426 (N_426,In_151,In_491);
and U427 (N_427,In_421,In_158);
and U428 (N_428,In_294,In_30);
nor U429 (N_429,In_27,In_132);
nor U430 (N_430,In_315,In_363);
and U431 (N_431,In_579,In_691);
nand U432 (N_432,In_92,In_44);
or U433 (N_433,In_83,In_240);
xnor U434 (N_434,In_329,In_284);
nand U435 (N_435,In_47,In_379);
nand U436 (N_436,In_599,In_447);
and U437 (N_437,In_740,In_462);
or U438 (N_438,In_592,In_51);
nor U439 (N_439,In_114,In_422);
and U440 (N_440,In_643,In_635);
nor U441 (N_441,In_405,In_478);
and U442 (N_442,In_403,In_296);
and U443 (N_443,In_38,In_374);
nor U444 (N_444,In_444,In_110);
xnor U445 (N_445,In_337,In_588);
nand U446 (N_446,In_118,In_689);
nor U447 (N_447,In_407,In_529);
nand U448 (N_448,In_225,In_638);
and U449 (N_449,In_728,In_368);
and U450 (N_450,In_443,In_488);
or U451 (N_451,In_280,In_534);
nand U452 (N_452,In_375,In_178);
nand U453 (N_453,In_136,In_57);
nand U454 (N_454,In_468,In_540);
or U455 (N_455,In_299,In_689);
nand U456 (N_456,In_686,In_71);
nor U457 (N_457,In_737,In_505);
and U458 (N_458,In_22,In_253);
nand U459 (N_459,In_61,In_479);
nand U460 (N_460,In_251,In_18);
or U461 (N_461,In_270,In_385);
nand U462 (N_462,In_309,In_731);
or U463 (N_463,In_665,In_96);
or U464 (N_464,In_488,In_569);
and U465 (N_465,In_688,In_283);
or U466 (N_466,In_211,In_541);
nor U467 (N_467,In_164,In_49);
nand U468 (N_468,In_486,In_647);
or U469 (N_469,In_658,In_255);
nand U470 (N_470,In_652,In_605);
and U471 (N_471,In_140,In_395);
and U472 (N_472,In_556,In_521);
or U473 (N_473,In_410,In_45);
or U474 (N_474,In_370,In_75);
and U475 (N_475,In_535,In_406);
and U476 (N_476,In_575,In_740);
nor U477 (N_477,In_283,In_133);
nand U478 (N_478,In_80,In_726);
and U479 (N_479,In_203,In_322);
nand U480 (N_480,In_68,In_194);
nand U481 (N_481,In_216,In_91);
or U482 (N_482,In_15,In_74);
or U483 (N_483,In_97,In_167);
nand U484 (N_484,In_116,In_256);
nand U485 (N_485,In_550,In_0);
nand U486 (N_486,In_362,In_109);
nor U487 (N_487,In_56,In_430);
and U488 (N_488,In_165,In_150);
or U489 (N_489,In_576,In_358);
nor U490 (N_490,In_717,In_26);
and U491 (N_491,In_111,In_142);
or U492 (N_492,In_115,In_250);
or U493 (N_493,In_22,In_501);
xor U494 (N_494,In_50,In_666);
and U495 (N_495,In_488,In_470);
nor U496 (N_496,In_722,In_656);
nor U497 (N_497,In_343,In_392);
and U498 (N_498,In_679,In_397);
nor U499 (N_499,In_171,In_447);
or U500 (N_500,In_432,In_279);
nand U501 (N_501,In_471,In_429);
nor U502 (N_502,In_57,In_507);
or U503 (N_503,In_416,In_712);
or U504 (N_504,In_400,In_20);
nor U505 (N_505,In_29,In_47);
or U506 (N_506,In_634,In_723);
nor U507 (N_507,In_314,In_376);
or U508 (N_508,In_620,In_220);
nand U509 (N_509,In_200,In_577);
or U510 (N_510,In_60,In_309);
and U511 (N_511,In_385,In_211);
nor U512 (N_512,In_122,In_74);
nand U513 (N_513,In_287,In_492);
nand U514 (N_514,In_235,In_522);
or U515 (N_515,In_508,In_374);
nand U516 (N_516,In_347,In_486);
and U517 (N_517,In_404,In_257);
nor U518 (N_518,In_354,In_245);
or U519 (N_519,In_269,In_533);
nor U520 (N_520,In_96,In_571);
nor U521 (N_521,In_697,In_594);
and U522 (N_522,In_359,In_78);
nor U523 (N_523,In_330,In_232);
and U524 (N_524,In_432,In_29);
nor U525 (N_525,In_603,In_657);
nor U526 (N_526,In_586,In_585);
nand U527 (N_527,In_590,In_288);
and U528 (N_528,In_82,In_52);
and U529 (N_529,In_78,In_437);
nor U530 (N_530,In_666,In_282);
nor U531 (N_531,In_360,In_444);
nand U532 (N_532,In_454,In_602);
nor U533 (N_533,In_619,In_69);
and U534 (N_534,In_438,In_167);
nand U535 (N_535,In_37,In_270);
nor U536 (N_536,In_666,In_639);
and U537 (N_537,In_75,In_188);
or U538 (N_538,In_80,In_656);
nor U539 (N_539,In_168,In_508);
or U540 (N_540,In_392,In_266);
and U541 (N_541,In_17,In_98);
or U542 (N_542,In_595,In_192);
nor U543 (N_543,In_396,In_80);
or U544 (N_544,In_691,In_159);
nand U545 (N_545,In_300,In_181);
nand U546 (N_546,In_588,In_641);
or U547 (N_547,In_477,In_357);
or U548 (N_548,In_426,In_113);
or U549 (N_549,In_635,In_232);
xor U550 (N_550,In_708,In_272);
nor U551 (N_551,In_176,In_105);
or U552 (N_552,In_443,In_469);
or U553 (N_553,In_476,In_397);
nor U554 (N_554,In_411,In_567);
and U555 (N_555,In_119,In_402);
nand U556 (N_556,In_429,In_498);
xor U557 (N_557,In_65,In_256);
nor U558 (N_558,In_714,In_424);
or U559 (N_559,In_233,In_304);
nand U560 (N_560,In_423,In_119);
nor U561 (N_561,In_414,In_79);
or U562 (N_562,In_89,In_158);
or U563 (N_563,In_35,In_61);
or U564 (N_564,In_569,In_610);
and U565 (N_565,In_566,In_316);
or U566 (N_566,In_346,In_224);
or U567 (N_567,In_367,In_93);
and U568 (N_568,In_687,In_694);
and U569 (N_569,In_383,In_10);
xor U570 (N_570,In_413,In_173);
and U571 (N_571,In_503,In_276);
nor U572 (N_572,In_178,In_576);
nor U573 (N_573,In_590,In_303);
nor U574 (N_574,In_382,In_683);
or U575 (N_575,In_112,In_713);
or U576 (N_576,In_571,In_606);
and U577 (N_577,In_93,In_164);
or U578 (N_578,In_355,In_121);
nor U579 (N_579,In_493,In_37);
or U580 (N_580,In_437,In_6);
nor U581 (N_581,In_556,In_564);
nor U582 (N_582,In_378,In_588);
and U583 (N_583,In_402,In_5);
nand U584 (N_584,In_92,In_512);
nor U585 (N_585,In_250,In_650);
nand U586 (N_586,In_636,In_267);
xnor U587 (N_587,In_328,In_573);
or U588 (N_588,In_12,In_51);
and U589 (N_589,In_230,In_719);
or U590 (N_590,In_608,In_733);
and U591 (N_591,In_51,In_580);
or U592 (N_592,In_543,In_147);
and U593 (N_593,In_225,In_304);
nand U594 (N_594,In_172,In_659);
and U595 (N_595,In_531,In_533);
xnor U596 (N_596,In_607,In_105);
xnor U597 (N_597,In_517,In_92);
xor U598 (N_598,In_35,In_156);
and U599 (N_599,In_312,In_637);
and U600 (N_600,In_118,In_376);
or U601 (N_601,In_357,In_114);
or U602 (N_602,In_411,In_469);
and U603 (N_603,In_678,In_690);
or U604 (N_604,In_150,In_229);
or U605 (N_605,In_148,In_197);
nor U606 (N_606,In_614,In_156);
nand U607 (N_607,In_512,In_19);
and U608 (N_608,In_263,In_61);
and U609 (N_609,In_239,In_453);
nor U610 (N_610,In_474,In_82);
and U611 (N_611,In_648,In_411);
nand U612 (N_612,In_534,In_703);
and U613 (N_613,In_521,In_34);
nor U614 (N_614,In_230,In_144);
nor U615 (N_615,In_102,In_300);
nor U616 (N_616,In_138,In_348);
nor U617 (N_617,In_657,In_461);
nand U618 (N_618,In_681,In_713);
nor U619 (N_619,In_98,In_483);
and U620 (N_620,In_469,In_684);
or U621 (N_621,In_585,In_61);
or U622 (N_622,In_494,In_159);
and U623 (N_623,In_246,In_202);
xor U624 (N_624,In_117,In_301);
or U625 (N_625,In_490,In_662);
and U626 (N_626,In_417,In_457);
nor U627 (N_627,In_261,In_291);
and U628 (N_628,In_197,In_465);
nand U629 (N_629,In_450,In_682);
and U630 (N_630,In_564,In_171);
nand U631 (N_631,In_364,In_746);
nand U632 (N_632,In_321,In_27);
nand U633 (N_633,In_25,In_193);
nor U634 (N_634,In_431,In_319);
or U635 (N_635,In_452,In_272);
nor U636 (N_636,In_744,In_55);
nor U637 (N_637,In_60,In_635);
nand U638 (N_638,In_464,In_85);
nand U639 (N_639,In_365,In_212);
or U640 (N_640,In_499,In_240);
nor U641 (N_641,In_192,In_25);
or U642 (N_642,In_686,In_122);
and U643 (N_643,In_668,In_48);
nand U644 (N_644,In_541,In_118);
xor U645 (N_645,In_436,In_264);
or U646 (N_646,In_291,In_564);
and U647 (N_647,In_81,In_374);
or U648 (N_648,In_599,In_168);
nand U649 (N_649,In_41,In_457);
nor U650 (N_650,In_683,In_343);
and U651 (N_651,In_416,In_136);
nor U652 (N_652,In_214,In_163);
and U653 (N_653,In_64,In_28);
or U654 (N_654,In_427,In_98);
nor U655 (N_655,In_261,In_405);
or U656 (N_656,In_75,In_277);
nor U657 (N_657,In_410,In_46);
nand U658 (N_658,In_702,In_187);
and U659 (N_659,In_253,In_224);
nand U660 (N_660,In_479,In_197);
nor U661 (N_661,In_346,In_112);
nor U662 (N_662,In_422,In_78);
xnor U663 (N_663,In_262,In_235);
and U664 (N_664,In_685,In_534);
nand U665 (N_665,In_347,In_207);
nor U666 (N_666,In_496,In_285);
nor U667 (N_667,In_71,In_283);
and U668 (N_668,In_270,In_279);
or U669 (N_669,In_423,In_151);
or U670 (N_670,In_538,In_730);
nand U671 (N_671,In_380,In_478);
and U672 (N_672,In_504,In_512);
nand U673 (N_673,In_0,In_685);
nand U674 (N_674,In_553,In_639);
and U675 (N_675,In_78,In_122);
nor U676 (N_676,In_704,In_587);
and U677 (N_677,In_131,In_183);
nand U678 (N_678,In_493,In_110);
nand U679 (N_679,In_366,In_476);
and U680 (N_680,In_145,In_397);
or U681 (N_681,In_360,In_78);
xor U682 (N_682,In_178,In_175);
and U683 (N_683,In_550,In_716);
or U684 (N_684,In_60,In_625);
nand U685 (N_685,In_378,In_119);
and U686 (N_686,In_641,In_708);
or U687 (N_687,In_265,In_38);
nand U688 (N_688,In_695,In_255);
and U689 (N_689,In_577,In_6);
and U690 (N_690,In_325,In_500);
nor U691 (N_691,In_492,In_270);
nand U692 (N_692,In_570,In_638);
nand U693 (N_693,In_733,In_507);
nor U694 (N_694,In_317,In_198);
nand U695 (N_695,In_443,In_410);
and U696 (N_696,In_557,In_560);
and U697 (N_697,In_672,In_402);
and U698 (N_698,In_194,In_39);
nand U699 (N_699,In_715,In_47);
and U700 (N_700,In_721,In_470);
nand U701 (N_701,In_627,In_271);
and U702 (N_702,In_368,In_409);
xor U703 (N_703,In_159,In_585);
and U704 (N_704,In_143,In_102);
and U705 (N_705,In_39,In_38);
or U706 (N_706,In_444,In_612);
and U707 (N_707,In_425,In_263);
nand U708 (N_708,In_742,In_152);
nor U709 (N_709,In_724,In_334);
or U710 (N_710,In_233,In_651);
or U711 (N_711,In_496,In_306);
nand U712 (N_712,In_504,In_47);
nor U713 (N_713,In_692,In_384);
nor U714 (N_714,In_407,In_589);
and U715 (N_715,In_659,In_101);
or U716 (N_716,In_418,In_520);
nand U717 (N_717,In_589,In_105);
nand U718 (N_718,In_547,In_103);
nor U719 (N_719,In_235,In_690);
nand U720 (N_720,In_607,In_178);
nand U721 (N_721,In_322,In_149);
nor U722 (N_722,In_260,In_712);
and U723 (N_723,In_492,In_434);
nand U724 (N_724,In_481,In_708);
nor U725 (N_725,In_20,In_35);
nor U726 (N_726,In_218,In_362);
or U727 (N_727,In_742,In_22);
or U728 (N_728,In_192,In_66);
and U729 (N_729,In_468,In_397);
nor U730 (N_730,In_240,In_82);
nor U731 (N_731,In_558,In_160);
or U732 (N_732,In_310,In_702);
and U733 (N_733,In_347,In_390);
or U734 (N_734,In_249,In_315);
or U735 (N_735,In_16,In_243);
nand U736 (N_736,In_490,In_721);
nand U737 (N_737,In_175,In_630);
and U738 (N_738,In_321,In_723);
nor U739 (N_739,In_198,In_732);
xor U740 (N_740,In_60,In_287);
and U741 (N_741,In_668,In_512);
or U742 (N_742,In_140,In_397);
nand U743 (N_743,In_391,In_270);
or U744 (N_744,In_13,In_513);
nor U745 (N_745,In_679,In_161);
nand U746 (N_746,In_167,In_415);
or U747 (N_747,In_53,In_694);
and U748 (N_748,In_57,In_731);
nand U749 (N_749,In_527,In_325);
or U750 (N_750,In_46,In_459);
nand U751 (N_751,In_372,In_698);
and U752 (N_752,In_136,In_168);
nor U753 (N_753,In_628,In_620);
nor U754 (N_754,In_725,In_399);
or U755 (N_755,In_611,In_3);
or U756 (N_756,In_624,In_19);
nor U757 (N_757,In_166,In_704);
and U758 (N_758,In_646,In_180);
nor U759 (N_759,In_484,In_624);
and U760 (N_760,In_620,In_496);
and U761 (N_761,In_481,In_12);
or U762 (N_762,In_449,In_437);
or U763 (N_763,In_374,In_747);
xor U764 (N_764,In_487,In_15);
or U765 (N_765,In_572,In_637);
and U766 (N_766,In_84,In_202);
nand U767 (N_767,In_356,In_261);
and U768 (N_768,In_244,In_149);
nand U769 (N_769,In_747,In_63);
nand U770 (N_770,In_131,In_646);
nor U771 (N_771,In_63,In_280);
or U772 (N_772,In_102,In_290);
or U773 (N_773,In_206,In_332);
nand U774 (N_774,In_477,In_271);
nand U775 (N_775,In_171,In_120);
nand U776 (N_776,In_389,In_399);
xnor U777 (N_777,In_581,In_354);
or U778 (N_778,In_157,In_67);
nor U779 (N_779,In_606,In_551);
or U780 (N_780,In_311,In_409);
or U781 (N_781,In_90,In_326);
xor U782 (N_782,In_573,In_484);
xnor U783 (N_783,In_364,In_439);
or U784 (N_784,In_130,In_61);
nor U785 (N_785,In_652,In_740);
and U786 (N_786,In_511,In_317);
nor U787 (N_787,In_500,In_146);
nand U788 (N_788,In_284,In_233);
or U789 (N_789,In_370,In_480);
or U790 (N_790,In_438,In_396);
nand U791 (N_791,In_652,In_540);
nor U792 (N_792,In_727,In_521);
or U793 (N_793,In_322,In_732);
or U794 (N_794,In_686,In_508);
or U795 (N_795,In_545,In_191);
or U796 (N_796,In_228,In_626);
nor U797 (N_797,In_702,In_116);
nor U798 (N_798,In_659,In_66);
nor U799 (N_799,In_378,In_411);
nor U800 (N_800,In_324,In_554);
nand U801 (N_801,In_373,In_186);
or U802 (N_802,In_448,In_671);
or U803 (N_803,In_315,In_238);
and U804 (N_804,In_91,In_313);
nor U805 (N_805,In_600,In_286);
or U806 (N_806,In_631,In_475);
nor U807 (N_807,In_578,In_279);
nand U808 (N_808,In_404,In_387);
and U809 (N_809,In_208,In_326);
nor U810 (N_810,In_388,In_683);
nor U811 (N_811,In_377,In_289);
and U812 (N_812,In_141,In_4);
nor U813 (N_813,In_144,In_350);
nand U814 (N_814,In_419,In_430);
or U815 (N_815,In_72,In_152);
or U816 (N_816,In_652,In_160);
nand U817 (N_817,In_183,In_228);
and U818 (N_818,In_39,In_506);
nand U819 (N_819,In_474,In_383);
and U820 (N_820,In_467,In_187);
and U821 (N_821,In_89,In_454);
nor U822 (N_822,In_421,In_687);
and U823 (N_823,In_375,In_454);
nand U824 (N_824,In_337,In_733);
and U825 (N_825,In_600,In_525);
nor U826 (N_826,In_287,In_290);
or U827 (N_827,In_386,In_507);
nor U828 (N_828,In_447,In_309);
or U829 (N_829,In_627,In_119);
nand U830 (N_830,In_158,In_587);
nor U831 (N_831,In_642,In_264);
nor U832 (N_832,In_517,In_581);
nand U833 (N_833,In_523,In_301);
or U834 (N_834,In_239,In_102);
and U835 (N_835,In_561,In_458);
or U836 (N_836,In_289,In_452);
and U837 (N_837,In_684,In_511);
or U838 (N_838,In_513,In_620);
nand U839 (N_839,In_127,In_424);
and U840 (N_840,In_170,In_749);
nor U841 (N_841,In_180,In_144);
and U842 (N_842,In_11,In_646);
or U843 (N_843,In_706,In_676);
and U844 (N_844,In_446,In_381);
nor U845 (N_845,In_679,In_53);
nor U846 (N_846,In_143,In_600);
and U847 (N_847,In_17,In_316);
nand U848 (N_848,In_240,In_374);
and U849 (N_849,In_36,In_630);
nor U850 (N_850,In_406,In_484);
and U851 (N_851,In_342,In_638);
or U852 (N_852,In_728,In_290);
or U853 (N_853,In_413,In_408);
or U854 (N_854,In_643,In_280);
nand U855 (N_855,In_390,In_610);
nor U856 (N_856,In_178,In_494);
xor U857 (N_857,In_595,In_657);
nor U858 (N_858,In_209,In_620);
and U859 (N_859,In_45,In_512);
and U860 (N_860,In_380,In_544);
and U861 (N_861,In_6,In_51);
or U862 (N_862,In_245,In_510);
or U863 (N_863,In_714,In_208);
nand U864 (N_864,In_253,In_608);
and U865 (N_865,In_357,In_514);
nand U866 (N_866,In_73,In_241);
nor U867 (N_867,In_34,In_676);
or U868 (N_868,In_475,In_558);
nand U869 (N_869,In_248,In_191);
nand U870 (N_870,In_656,In_156);
nor U871 (N_871,In_18,In_351);
nand U872 (N_872,In_58,In_552);
or U873 (N_873,In_94,In_689);
nand U874 (N_874,In_382,In_80);
nor U875 (N_875,In_658,In_217);
or U876 (N_876,In_32,In_732);
and U877 (N_877,In_421,In_684);
or U878 (N_878,In_460,In_549);
nand U879 (N_879,In_389,In_617);
and U880 (N_880,In_356,In_669);
nor U881 (N_881,In_242,In_737);
or U882 (N_882,In_392,In_623);
nor U883 (N_883,In_474,In_550);
nand U884 (N_884,In_117,In_702);
or U885 (N_885,In_720,In_706);
nor U886 (N_886,In_346,In_48);
and U887 (N_887,In_421,In_225);
or U888 (N_888,In_240,In_284);
and U889 (N_889,In_640,In_359);
nor U890 (N_890,In_16,In_60);
nor U891 (N_891,In_273,In_485);
nand U892 (N_892,In_740,In_738);
nor U893 (N_893,In_708,In_516);
or U894 (N_894,In_664,In_604);
nor U895 (N_895,In_279,In_590);
xnor U896 (N_896,In_192,In_328);
or U897 (N_897,In_611,In_495);
nor U898 (N_898,In_191,In_612);
nand U899 (N_899,In_676,In_426);
or U900 (N_900,In_308,In_123);
or U901 (N_901,In_522,In_585);
and U902 (N_902,In_123,In_473);
or U903 (N_903,In_642,In_393);
xnor U904 (N_904,In_364,In_545);
or U905 (N_905,In_650,In_389);
nor U906 (N_906,In_38,In_698);
or U907 (N_907,In_92,In_563);
nor U908 (N_908,In_81,In_513);
nand U909 (N_909,In_222,In_47);
and U910 (N_910,In_131,In_136);
or U911 (N_911,In_199,In_597);
nand U912 (N_912,In_577,In_366);
or U913 (N_913,In_401,In_19);
nand U914 (N_914,In_242,In_477);
nand U915 (N_915,In_143,In_164);
nand U916 (N_916,In_291,In_686);
nand U917 (N_917,In_409,In_265);
and U918 (N_918,In_465,In_105);
and U919 (N_919,In_372,In_688);
or U920 (N_920,In_633,In_591);
and U921 (N_921,In_738,In_286);
nand U922 (N_922,In_463,In_676);
and U923 (N_923,In_74,In_424);
xor U924 (N_924,In_550,In_294);
nor U925 (N_925,In_194,In_608);
nand U926 (N_926,In_520,In_122);
nor U927 (N_927,In_397,In_478);
or U928 (N_928,In_500,In_219);
or U929 (N_929,In_602,In_695);
nor U930 (N_930,In_694,In_15);
or U931 (N_931,In_352,In_329);
and U932 (N_932,In_65,In_569);
nand U933 (N_933,In_593,In_299);
or U934 (N_934,In_569,In_108);
or U935 (N_935,In_642,In_319);
and U936 (N_936,In_91,In_177);
and U937 (N_937,In_175,In_499);
or U938 (N_938,In_226,In_676);
and U939 (N_939,In_743,In_191);
or U940 (N_940,In_34,In_145);
nand U941 (N_941,In_535,In_385);
nand U942 (N_942,In_274,In_104);
and U943 (N_943,In_456,In_381);
nor U944 (N_944,In_284,In_579);
and U945 (N_945,In_418,In_320);
or U946 (N_946,In_193,In_645);
or U947 (N_947,In_453,In_739);
or U948 (N_948,In_708,In_661);
or U949 (N_949,In_131,In_336);
or U950 (N_950,In_445,In_476);
nor U951 (N_951,In_199,In_581);
nand U952 (N_952,In_328,In_95);
and U953 (N_953,In_132,In_243);
nor U954 (N_954,In_294,In_364);
and U955 (N_955,In_41,In_215);
nor U956 (N_956,In_55,In_571);
nand U957 (N_957,In_729,In_702);
nor U958 (N_958,In_9,In_32);
nand U959 (N_959,In_458,In_104);
and U960 (N_960,In_95,In_408);
nand U961 (N_961,In_50,In_59);
and U962 (N_962,In_170,In_175);
nand U963 (N_963,In_495,In_18);
nand U964 (N_964,In_600,In_387);
nand U965 (N_965,In_718,In_527);
nand U966 (N_966,In_195,In_402);
and U967 (N_967,In_627,In_148);
or U968 (N_968,In_664,In_335);
nand U969 (N_969,In_15,In_335);
or U970 (N_970,In_109,In_470);
nand U971 (N_971,In_390,In_669);
nand U972 (N_972,In_123,In_244);
nand U973 (N_973,In_468,In_347);
nand U974 (N_974,In_484,In_555);
or U975 (N_975,In_102,In_181);
nand U976 (N_976,In_421,In_734);
nor U977 (N_977,In_220,In_485);
and U978 (N_978,In_237,In_130);
or U979 (N_979,In_555,In_91);
nor U980 (N_980,In_210,In_572);
nand U981 (N_981,In_356,In_83);
or U982 (N_982,In_343,In_470);
and U983 (N_983,In_464,In_717);
nor U984 (N_984,In_649,In_717);
nand U985 (N_985,In_178,In_93);
nand U986 (N_986,In_560,In_480);
nand U987 (N_987,In_255,In_167);
and U988 (N_988,In_81,In_371);
nor U989 (N_989,In_186,In_436);
nor U990 (N_990,In_158,In_658);
and U991 (N_991,In_745,In_244);
nor U992 (N_992,In_506,In_301);
nand U993 (N_993,In_663,In_728);
nor U994 (N_994,In_126,In_128);
nand U995 (N_995,In_15,In_331);
nand U996 (N_996,In_676,In_716);
nand U997 (N_997,In_194,In_590);
or U998 (N_998,In_533,In_120);
or U999 (N_999,In_362,In_736);
and U1000 (N_1000,In_369,In_670);
and U1001 (N_1001,In_267,In_749);
nor U1002 (N_1002,In_180,In_585);
nor U1003 (N_1003,In_241,In_88);
nand U1004 (N_1004,In_285,In_55);
nor U1005 (N_1005,In_117,In_573);
nand U1006 (N_1006,In_318,In_226);
or U1007 (N_1007,In_154,In_707);
nor U1008 (N_1008,In_458,In_461);
nor U1009 (N_1009,In_144,In_488);
nand U1010 (N_1010,In_596,In_574);
or U1011 (N_1011,In_386,In_503);
or U1012 (N_1012,In_697,In_273);
or U1013 (N_1013,In_492,In_553);
nand U1014 (N_1014,In_621,In_41);
and U1015 (N_1015,In_666,In_425);
or U1016 (N_1016,In_417,In_209);
nor U1017 (N_1017,In_730,In_73);
and U1018 (N_1018,In_213,In_111);
nand U1019 (N_1019,In_508,In_319);
nor U1020 (N_1020,In_646,In_302);
nor U1021 (N_1021,In_543,In_334);
and U1022 (N_1022,In_40,In_406);
nor U1023 (N_1023,In_736,In_12);
nor U1024 (N_1024,In_58,In_79);
or U1025 (N_1025,In_575,In_38);
and U1026 (N_1026,In_122,In_548);
nand U1027 (N_1027,In_186,In_631);
and U1028 (N_1028,In_78,In_130);
nor U1029 (N_1029,In_192,In_265);
or U1030 (N_1030,In_398,In_40);
nand U1031 (N_1031,In_431,In_422);
nand U1032 (N_1032,In_102,In_115);
and U1033 (N_1033,In_149,In_424);
or U1034 (N_1034,In_604,In_169);
xnor U1035 (N_1035,In_126,In_573);
and U1036 (N_1036,In_198,In_41);
nor U1037 (N_1037,In_367,In_151);
and U1038 (N_1038,In_236,In_459);
nor U1039 (N_1039,In_75,In_84);
nor U1040 (N_1040,In_449,In_23);
nor U1041 (N_1041,In_588,In_283);
nand U1042 (N_1042,In_291,In_725);
and U1043 (N_1043,In_505,In_608);
and U1044 (N_1044,In_606,In_662);
and U1045 (N_1045,In_519,In_491);
nand U1046 (N_1046,In_726,In_330);
nand U1047 (N_1047,In_344,In_542);
and U1048 (N_1048,In_255,In_199);
nand U1049 (N_1049,In_52,In_669);
nor U1050 (N_1050,In_77,In_739);
or U1051 (N_1051,In_249,In_374);
and U1052 (N_1052,In_70,In_663);
nor U1053 (N_1053,In_511,In_243);
nand U1054 (N_1054,In_59,In_523);
nor U1055 (N_1055,In_475,In_679);
or U1056 (N_1056,In_706,In_343);
and U1057 (N_1057,In_81,In_594);
or U1058 (N_1058,In_134,In_639);
nand U1059 (N_1059,In_450,In_73);
nand U1060 (N_1060,In_722,In_587);
or U1061 (N_1061,In_63,In_184);
and U1062 (N_1062,In_532,In_467);
or U1063 (N_1063,In_671,In_700);
xor U1064 (N_1064,In_656,In_410);
nand U1065 (N_1065,In_470,In_305);
nand U1066 (N_1066,In_7,In_441);
nor U1067 (N_1067,In_380,In_509);
or U1068 (N_1068,In_109,In_466);
nor U1069 (N_1069,In_169,In_640);
nand U1070 (N_1070,In_71,In_104);
nor U1071 (N_1071,In_387,In_731);
xnor U1072 (N_1072,In_481,In_455);
or U1073 (N_1073,In_107,In_591);
nand U1074 (N_1074,In_240,In_441);
and U1075 (N_1075,In_564,In_212);
xor U1076 (N_1076,In_342,In_174);
nor U1077 (N_1077,In_549,In_717);
nand U1078 (N_1078,In_555,In_551);
nor U1079 (N_1079,In_692,In_512);
nand U1080 (N_1080,In_381,In_220);
or U1081 (N_1081,In_81,In_634);
and U1082 (N_1082,In_73,In_603);
or U1083 (N_1083,In_554,In_644);
or U1084 (N_1084,In_581,In_582);
nor U1085 (N_1085,In_599,In_289);
and U1086 (N_1086,In_265,In_304);
and U1087 (N_1087,In_554,In_187);
or U1088 (N_1088,In_407,In_592);
or U1089 (N_1089,In_324,In_521);
and U1090 (N_1090,In_358,In_411);
or U1091 (N_1091,In_716,In_732);
nand U1092 (N_1092,In_547,In_92);
and U1093 (N_1093,In_144,In_132);
or U1094 (N_1094,In_399,In_384);
and U1095 (N_1095,In_166,In_535);
nor U1096 (N_1096,In_558,In_41);
nor U1097 (N_1097,In_301,In_185);
nor U1098 (N_1098,In_327,In_276);
nor U1099 (N_1099,In_734,In_215);
nor U1100 (N_1100,In_259,In_384);
or U1101 (N_1101,In_717,In_333);
nor U1102 (N_1102,In_359,In_602);
nor U1103 (N_1103,In_306,In_553);
and U1104 (N_1104,In_501,In_499);
and U1105 (N_1105,In_661,In_327);
or U1106 (N_1106,In_528,In_335);
nand U1107 (N_1107,In_146,In_361);
nand U1108 (N_1108,In_399,In_138);
nand U1109 (N_1109,In_198,In_342);
and U1110 (N_1110,In_283,In_214);
or U1111 (N_1111,In_114,In_520);
nor U1112 (N_1112,In_418,In_217);
and U1113 (N_1113,In_499,In_704);
nand U1114 (N_1114,In_237,In_683);
or U1115 (N_1115,In_122,In_491);
or U1116 (N_1116,In_422,In_457);
xor U1117 (N_1117,In_41,In_159);
nand U1118 (N_1118,In_687,In_372);
and U1119 (N_1119,In_213,In_627);
or U1120 (N_1120,In_546,In_453);
or U1121 (N_1121,In_195,In_711);
and U1122 (N_1122,In_471,In_217);
or U1123 (N_1123,In_681,In_731);
nand U1124 (N_1124,In_409,In_587);
or U1125 (N_1125,In_261,In_307);
nand U1126 (N_1126,In_436,In_510);
nor U1127 (N_1127,In_430,In_454);
nor U1128 (N_1128,In_284,In_92);
or U1129 (N_1129,In_655,In_44);
or U1130 (N_1130,In_80,In_420);
and U1131 (N_1131,In_134,In_132);
or U1132 (N_1132,In_685,In_99);
nor U1133 (N_1133,In_504,In_164);
nand U1134 (N_1134,In_436,In_138);
nand U1135 (N_1135,In_480,In_556);
nor U1136 (N_1136,In_257,In_740);
or U1137 (N_1137,In_202,In_24);
or U1138 (N_1138,In_317,In_55);
and U1139 (N_1139,In_173,In_716);
or U1140 (N_1140,In_389,In_692);
or U1141 (N_1141,In_281,In_420);
nor U1142 (N_1142,In_561,In_413);
and U1143 (N_1143,In_688,In_26);
nand U1144 (N_1144,In_217,In_563);
and U1145 (N_1145,In_336,In_506);
nor U1146 (N_1146,In_145,In_136);
nor U1147 (N_1147,In_276,In_580);
xnor U1148 (N_1148,In_276,In_119);
nor U1149 (N_1149,In_74,In_429);
nand U1150 (N_1150,In_123,In_563);
or U1151 (N_1151,In_626,In_592);
or U1152 (N_1152,In_595,In_690);
or U1153 (N_1153,In_237,In_159);
nor U1154 (N_1154,In_86,In_697);
and U1155 (N_1155,In_598,In_657);
nand U1156 (N_1156,In_11,In_725);
nor U1157 (N_1157,In_105,In_267);
nor U1158 (N_1158,In_116,In_480);
and U1159 (N_1159,In_234,In_344);
nand U1160 (N_1160,In_182,In_452);
nand U1161 (N_1161,In_706,In_372);
and U1162 (N_1162,In_11,In_247);
xnor U1163 (N_1163,In_339,In_133);
nand U1164 (N_1164,In_591,In_658);
and U1165 (N_1165,In_10,In_115);
or U1166 (N_1166,In_29,In_69);
nand U1167 (N_1167,In_145,In_637);
and U1168 (N_1168,In_628,In_108);
nand U1169 (N_1169,In_632,In_151);
and U1170 (N_1170,In_412,In_120);
xnor U1171 (N_1171,In_400,In_623);
nor U1172 (N_1172,In_664,In_430);
nand U1173 (N_1173,In_135,In_178);
and U1174 (N_1174,In_600,In_239);
or U1175 (N_1175,In_669,In_242);
nor U1176 (N_1176,In_427,In_181);
and U1177 (N_1177,In_650,In_687);
and U1178 (N_1178,In_10,In_124);
and U1179 (N_1179,In_0,In_672);
or U1180 (N_1180,In_517,In_3);
or U1181 (N_1181,In_550,In_97);
and U1182 (N_1182,In_508,In_455);
and U1183 (N_1183,In_547,In_442);
and U1184 (N_1184,In_201,In_55);
nand U1185 (N_1185,In_19,In_627);
or U1186 (N_1186,In_418,In_601);
nand U1187 (N_1187,In_478,In_43);
or U1188 (N_1188,In_78,In_74);
nor U1189 (N_1189,In_263,In_580);
and U1190 (N_1190,In_138,In_524);
xor U1191 (N_1191,In_383,In_481);
nand U1192 (N_1192,In_74,In_69);
or U1193 (N_1193,In_457,In_468);
or U1194 (N_1194,In_209,In_658);
nor U1195 (N_1195,In_490,In_125);
nand U1196 (N_1196,In_486,In_491);
or U1197 (N_1197,In_479,In_307);
or U1198 (N_1198,In_666,In_582);
nand U1199 (N_1199,In_341,In_673);
and U1200 (N_1200,In_229,In_589);
nand U1201 (N_1201,In_270,In_328);
nand U1202 (N_1202,In_173,In_379);
nor U1203 (N_1203,In_736,In_714);
or U1204 (N_1204,In_241,In_206);
or U1205 (N_1205,In_700,In_162);
and U1206 (N_1206,In_685,In_431);
or U1207 (N_1207,In_745,In_742);
nor U1208 (N_1208,In_287,In_579);
nand U1209 (N_1209,In_116,In_527);
nor U1210 (N_1210,In_318,In_359);
xor U1211 (N_1211,In_304,In_543);
or U1212 (N_1212,In_401,In_116);
and U1213 (N_1213,In_1,In_138);
nand U1214 (N_1214,In_408,In_598);
or U1215 (N_1215,In_383,In_577);
nand U1216 (N_1216,In_143,In_342);
nor U1217 (N_1217,In_199,In_273);
nand U1218 (N_1218,In_277,In_211);
nor U1219 (N_1219,In_311,In_661);
and U1220 (N_1220,In_281,In_333);
or U1221 (N_1221,In_95,In_416);
and U1222 (N_1222,In_381,In_287);
or U1223 (N_1223,In_259,In_134);
or U1224 (N_1224,In_594,In_250);
and U1225 (N_1225,In_62,In_374);
nand U1226 (N_1226,In_16,In_203);
nand U1227 (N_1227,In_130,In_414);
or U1228 (N_1228,In_100,In_427);
nand U1229 (N_1229,In_26,In_310);
and U1230 (N_1230,In_303,In_400);
or U1231 (N_1231,In_448,In_14);
and U1232 (N_1232,In_448,In_386);
nand U1233 (N_1233,In_547,In_647);
nor U1234 (N_1234,In_738,In_569);
nor U1235 (N_1235,In_334,In_277);
or U1236 (N_1236,In_100,In_713);
or U1237 (N_1237,In_343,In_594);
and U1238 (N_1238,In_221,In_40);
nand U1239 (N_1239,In_571,In_411);
or U1240 (N_1240,In_456,In_686);
nand U1241 (N_1241,In_443,In_480);
nor U1242 (N_1242,In_551,In_712);
or U1243 (N_1243,In_260,In_358);
xor U1244 (N_1244,In_556,In_686);
or U1245 (N_1245,In_216,In_295);
nand U1246 (N_1246,In_485,In_275);
or U1247 (N_1247,In_670,In_696);
and U1248 (N_1248,In_1,In_711);
nand U1249 (N_1249,In_592,In_234);
or U1250 (N_1250,In_438,In_558);
nor U1251 (N_1251,In_342,In_58);
and U1252 (N_1252,In_365,In_195);
nor U1253 (N_1253,In_50,In_745);
nand U1254 (N_1254,In_745,In_603);
and U1255 (N_1255,In_620,In_379);
nand U1256 (N_1256,In_517,In_556);
or U1257 (N_1257,In_706,In_165);
nand U1258 (N_1258,In_146,In_72);
nor U1259 (N_1259,In_146,In_2);
nand U1260 (N_1260,In_301,In_631);
or U1261 (N_1261,In_117,In_296);
and U1262 (N_1262,In_13,In_247);
nor U1263 (N_1263,In_188,In_173);
nor U1264 (N_1264,In_43,In_667);
nand U1265 (N_1265,In_498,In_114);
nand U1266 (N_1266,In_96,In_489);
nand U1267 (N_1267,In_280,In_501);
nand U1268 (N_1268,In_1,In_582);
nor U1269 (N_1269,In_215,In_368);
nand U1270 (N_1270,In_631,In_341);
or U1271 (N_1271,In_165,In_157);
xnor U1272 (N_1272,In_214,In_387);
nor U1273 (N_1273,In_27,In_533);
nand U1274 (N_1274,In_281,In_101);
nand U1275 (N_1275,In_412,In_113);
and U1276 (N_1276,In_701,In_611);
nor U1277 (N_1277,In_748,In_449);
and U1278 (N_1278,In_676,In_232);
and U1279 (N_1279,In_688,In_566);
and U1280 (N_1280,In_383,In_566);
and U1281 (N_1281,In_140,In_363);
or U1282 (N_1282,In_342,In_426);
or U1283 (N_1283,In_291,In_619);
xor U1284 (N_1284,In_177,In_151);
or U1285 (N_1285,In_191,In_501);
and U1286 (N_1286,In_705,In_29);
nor U1287 (N_1287,In_192,In_300);
and U1288 (N_1288,In_160,In_405);
nor U1289 (N_1289,In_445,In_680);
nand U1290 (N_1290,In_418,In_581);
nor U1291 (N_1291,In_271,In_154);
nand U1292 (N_1292,In_117,In_201);
nor U1293 (N_1293,In_475,In_165);
and U1294 (N_1294,In_451,In_337);
nand U1295 (N_1295,In_327,In_257);
nand U1296 (N_1296,In_49,In_98);
or U1297 (N_1297,In_527,In_724);
or U1298 (N_1298,In_126,In_357);
nand U1299 (N_1299,In_426,In_598);
nand U1300 (N_1300,In_154,In_370);
nand U1301 (N_1301,In_279,In_671);
xnor U1302 (N_1302,In_20,In_306);
nand U1303 (N_1303,In_346,In_192);
nor U1304 (N_1304,In_0,In_482);
xor U1305 (N_1305,In_524,In_414);
or U1306 (N_1306,In_30,In_323);
nand U1307 (N_1307,In_151,In_249);
and U1308 (N_1308,In_117,In_53);
or U1309 (N_1309,In_307,In_154);
xor U1310 (N_1310,In_89,In_196);
or U1311 (N_1311,In_500,In_433);
nand U1312 (N_1312,In_332,In_212);
and U1313 (N_1313,In_85,In_77);
and U1314 (N_1314,In_459,In_683);
nand U1315 (N_1315,In_17,In_96);
nand U1316 (N_1316,In_678,In_350);
nand U1317 (N_1317,In_15,In_12);
nand U1318 (N_1318,In_133,In_149);
nand U1319 (N_1319,In_151,In_88);
nor U1320 (N_1320,In_633,In_6);
or U1321 (N_1321,In_366,In_244);
and U1322 (N_1322,In_536,In_392);
or U1323 (N_1323,In_618,In_373);
or U1324 (N_1324,In_476,In_345);
nand U1325 (N_1325,In_230,In_316);
xor U1326 (N_1326,In_664,In_294);
nand U1327 (N_1327,In_26,In_466);
and U1328 (N_1328,In_317,In_376);
nor U1329 (N_1329,In_424,In_430);
or U1330 (N_1330,In_729,In_5);
and U1331 (N_1331,In_96,In_635);
nor U1332 (N_1332,In_280,In_450);
or U1333 (N_1333,In_696,In_337);
and U1334 (N_1334,In_138,In_491);
nand U1335 (N_1335,In_131,In_218);
nand U1336 (N_1336,In_703,In_182);
nor U1337 (N_1337,In_589,In_489);
or U1338 (N_1338,In_659,In_222);
or U1339 (N_1339,In_553,In_672);
and U1340 (N_1340,In_378,In_226);
and U1341 (N_1341,In_600,In_653);
xnor U1342 (N_1342,In_467,In_102);
nor U1343 (N_1343,In_478,In_140);
nand U1344 (N_1344,In_246,In_733);
nor U1345 (N_1345,In_616,In_169);
nand U1346 (N_1346,In_664,In_238);
nand U1347 (N_1347,In_495,In_459);
nor U1348 (N_1348,In_328,In_691);
xnor U1349 (N_1349,In_41,In_306);
nor U1350 (N_1350,In_641,In_689);
and U1351 (N_1351,In_263,In_275);
or U1352 (N_1352,In_282,In_149);
nand U1353 (N_1353,In_94,In_548);
or U1354 (N_1354,In_370,In_331);
nor U1355 (N_1355,In_653,In_114);
or U1356 (N_1356,In_262,In_53);
nand U1357 (N_1357,In_711,In_371);
or U1358 (N_1358,In_174,In_407);
nor U1359 (N_1359,In_578,In_336);
nor U1360 (N_1360,In_681,In_406);
and U1361 (N_1361,In_488,In_347);
and U1362 (N_1362,In_86,In_71);
nand U1363 (N_1363,In_667,In_672);
nand U1364 (N_1364,In_454,In_521);
or U1365 (N_1365,In_517,In_440);
nor U1366 (N_1366,In_189,In_618);
and U1367 (N_1367,In_391,In_626);
nor U1368 (N_1368,In_591,In_30);
xnor U1369 (N_1369,In_183,In_28);
nand U1370 (N_1370,In_125,In_594);
nor U1371 (N_1371,In_424,In_145);
and U1372 (N_1372,In_272,In_423);
nor U1373 (N_1373,In_499,In_593);
nor U1374 (N_1374,In_0,In_264);
xnor U1375 (N_1375,In_64,In_353);
nand U1376 (N_1376,In_495,In_596);
nor U1377 (N_1377,In_128,In_314);
nand U1378 (N_1378,In_206,In_142);
and U1379 (N_1379,In_456,In_629);
or U1380 (N_1380,In_727,In_333);
nand U1381 (N_1381,In_398,In_399);
nand U1382 (N_1382,In_122,In_197);
or U1383 (N_1383,In_697,In_737);
nor U1384 (N_1384,In_518,In_390);
and U1385 (N_1385,In_68,In_224);
and U1386 (N_1386,In_303,In_115);
and U1387 (N_1387,In_292,In_625);
nor U1388 (N_1388,In_87,In_80);
and U1389 (N_1389,In_269,In_289);
or U1390 (N_1390,In_604,In_705);
or U1391 (N_1391,In_394,In_637);
and U1392 (N_1392,In_232,In_432);
and U1393 (N_1393,In_701,In_128);
nor U1394 (N_1394,In_251,In_544);
nor U1395 (N_1395,In_118,In_359);
nand U1396 (N_1396,In_315,In_253);
nor U1397 (N_1397,In_40,In_492);
nand U1398 (N_1398,In_222,In_68);
or U1399 (N_1399,In_604,In_470);
nor U1400 (N_1400,In_641,In_235);
and U1401 (N_1401,In_511,In_650);
and U1402 (N_1402,In_473,In_22);
nand U1403 (N_1403,In_43,In_233);
or U1404 (N_1404,In_177,In_468);
and U1405 (N_1405,In_637,In_79);
and U1406 (N_1406,In_728,In_301);
and U1407 (N_1407,In_354,In_516);
and U1408 (N_1408,In_149,In_188);
nand U1409 (N_1409,In_68,In_713);
or U1410 (N_1410,In_98,In_411);
nor U1411 (N_1411,In_447,In_616);
and U1412 (N_1412,In_92,In_270);
nand U1413 (N_1413,In_137,In_720);
nor U1414 (N_1414,In_2,In_463);
and U1415 (N_1415,In_147,In_402);
or U1416 (N_1416,In_130,In_181);
nand U1417 (N_1417,In_464,In_277);
and U1418 (N_1418,In_326,In_731);
or U1419 (N_1419,In_403,In_593);
and U1420 (N_1420,In_237,In_105);
or U1421 (N_1421,In_580,In_469);
nor U1422 (N_1422,In_358,In_210);
or U1423 (N_1423,In_439,In_631);
and U1424 (N_1424,In_538,In_286);
and U1425 (N_1425,In_655,In_385);
nand U1426 (N_1426,In_443,In_610);
nor U1427 (N_1427,In_13,In_420);
or U1428 (N_1428,In_1,In_647);
or U1429 (N_1429,In_276,In_404);
nor U1430 (N_1430,In_117,In_246);
or U1431 (N_1431,In_290,In_421);
and U1432 (N_1432,In_274,In_744);
nand U1433 (N_1433,In_57,In_349);
or U1434 (N_1434,In_601,In_676);
or U1435 (N_1435,In_288,In_396);
or U1436 (N_1436,In_299,In_496);
and U1437 (N_1437,In_636,In_591);
nand U1438 (N_1438,In_223,In_517);
and U1439 (N_1439,In_244,In_545);
nand U1440 (N_1440,In_478,In_0);
nor U1441 (N_1441,In_554,In_361);
nand U1442 (N_1442,In_267,In_63);
nor U1443 (N_1443,In_413,In_235);
and U1444 (N_1444,In_287,In_129);
or U1445 (N_1445,In_408,In_467);
nor U1446 (N_1446,In_295,In_648);
or U1447 (N_1447,In_320,In_686);
nand U1448 (N_1448,In_410,In_608);
or U1449 (N_1449,In_499,In_259);
nor U1450 (N_1450,In_654,In_596);
nor U1451 (N_1451,In_728,In_59);
nand U1452 (N_1452,In_152,In_303);
or U1453 (N_1453,In_75,In_427);
nand U1454 (N_1454,In_697,In_332);
and U1455 (N_1455,In_419,In_272);
nor U1456 (N_1456,In_220,In_175);
nand U1457 (N_1457,In_550,In_4);
or U1458 (N_1458,In_27,In_396);
nor U1459 (N_1459,In_715,In_736);
and U1460 (N_1460,In_68,In_156);
nor U1461 (N_1461,In_127,In_159);
or U1462 (N_1462,In_570,In_66);
or U1463 (N_1463,In_400,In_513);
or U1464 (N_1464,In_506,In_675);
and U1465 (N_1465,In_709,In_289);
nand U1466 (N_1466,In_180,In_113);
or U1467 (N_1467,In_275,In_39);
nor U1468 (N_1468,In_151,In_711);
and U1469 (N_1469,In_213,In_658);
nor U1470 (N_1470,In_340,In_557);
or U1471 (N_1471,In_720,In_308);
xnor U1472 (N_1472,In_195,In_296);
nor U1473 (N_1473,In_317,In_278);
and U1474 (N_1474,In_591,In_490);
nor U1475 (N_1475,In_327,In_676);
and U1476 (N_1476,In_527,In_485);
and U1477 (N_1477,In_170,In_63);
or U1478 (N_1478,In_369,In_73);
or U1479 (N_1479,In_50,In_669);
nand U1480 (N_1480,In_464,In_313);
and U1481 (N_1481,In_134,In_679);
nor U1482 (N_1482,In_183,In_120);
and U1483 (N_1483,In_394,In_538);
or U1484 (N_1484,In_427,In_472);
xor U1485 (N_1485,In_717,In_199);
nand U1486 (N_1486,In_130,In_569);
and U1487 (N_1487,In_127,In_398);
nand U1488 (N_1488,In_330,In_634);
nand U1489 (N_1489,In_191,In_374);
nand U1490 (N_1490,In_115,In_241);
and U1491 (N_1491,In_475,In_210);
or U1492 (N_1492,In_704,In_605);
or U1493 (N_1493,In_369,In_365);
nand U1494 (N_1494,In_623,In_725);
nor U1495 (N_1495,In_315,In_374);
and U1496 (N_1496,In_514,In_28);
nand U1497 (N_1497,In_18,In_300);
and U1498 (N_1498,In_56,In_396);
or U1499 (N_1499,In_717,In_120);
nand U1500 (N_1500,In_695,In_138);
nor U1501 (N_1501,In_693,In_242);
nand U1502 (N_1502,In_624,In_171);
nand U1503 (N_1503,In_452,In_569);
or U1504 (N_1504,In_187,In_595);
nand U1505 (N_1505,In_135,In_109);
nand U1506 (N_1506,In_677,In_586);
nand U1507 (N_1507,In_510,In_540);
nor U1508 (N_1508,In_245,In_254);
nand U1509 (N_1509,In_11,In_501);
nand U1510 (N_1510,In_460,In_51);
or U1511 (N_1511,In_123,In_294);
nand U1512 (N_1512,In_495,In_288);
nand U1513 (N_1513,In_134,In_743);
and U1514 (N_1514,In_741,In_606);
and U1515 (N_1515,In_64,In_449);
nor U1516 (N_1516,In_423,In_581);
nand U1517 (N_1517,In_212,In_417);
and U1518 (N_1518,In_725,In_482);
or U1519 (N_1519,In_44,In_694);
nor U1520 (N_1520,In_349,In_437);
or U1521 (N_1521,In_670,In_710);
nor U1522 (N_1522,In_174,In_600);
nor U1523 (N_1523,In_136,In_33);
and U1524 (N_1524,In_373,In_743);
or U1525 (N_1525,In_327,In_739);
nand U1526 (N_1526,In_333,In_174);
and U1527 (N_1527,In_409,In_710);
nor U1528 (N_1528,In_234,In_616);
and U1529 (N_1529,In_731,In_360);
nor U1530 (N_1530,In_737,In_325);
and U1531 (N_1531,In_340,In_479);
and U1532 (N_1532,In_474,In_324);
nor U1533 (N_1533,In_374,In_85);
nor U1534 (N_1534,In_667,In_740);
nand U1535 (N_1535,In_364,In_390);
and U1536 (N_1536,In_713,In_195);
nor U1537 (N_1537,In_743,In_262);
and U1538 (N_1538,In_703,In_725);
nand U1539 (N_1539,In_288,In_309);
xor U1540 (N_1540,In_62,In_474);
nand U1541 (N_1541,In_442,In_244);
or U1542 (N_1542,In_101,In_488);
and U1543 (N_1543,In_692,In_34);
or U1544 (N_1544,In_437,In_484);
nor U1545 (N_1545,In_442,In_500);
xnor U1546 (N_1546,In_184,In_480);
nor U1547 (N_1547,In_369,In_528);
nor U1548 (N_1548,In_544,In_257);
nor U1549 (N_1549,In_534,In_316);
nand U1550 (N_1550,In_534,In_397);
and U1551 (N_1551,In_93,In_307);
nand U1552 (N_1552,In_291,In_104);
and U1553 (N_1553,In_740,In_524);
or U1554 (N_1554,In_514,In_654);
nor U1555 (N_1555,In_402,In_475);
nor U1556 (N_1556,In_735,In_287);
xnor U1557 (N_1557,In_481,In_654);
nor U1558 (N_1558,In_700,In_81);
and U1559 (N_1559,In_183,In_550);
nor U1560 (N_1560,In_126,In_234);
or U1561 (N_1561,In_373,In_437);
and U1562 (N_1562,In_277,In_186);
nand U1563 (N_1563,In_248,In_49);
or U1564 (N_1564,In_129,In_121);
or U1565 (N_1565,In_675,In_145);
nor U1566 (N_1566,In_77,In_597);
or U1567 (N_1567,In_303,In_435);
and U1568 (N_1568,In_36,In_708);
nor U1569 (N_1569,In_626,In_314);
and U1570 (N_1570,In_643,In_460);
or U1571 (N_1571,In_45,In_590);
nor U1572 (N_1572,In_448,In_738);
nor U1573 (N_1573,In_735,In_239);
and U1574 (N_1574,In_210,In_11);
nor U1575 (N_1575,In_681,In_741);
and U1576 (N_1576,In_180,In_248);
nor U1577 (N_1577,In_667,In_666);
and U1578 (N_1578,In_41,In_671);
and U1579 (N_1579,In_428,In_313);
or U1580 (N_1580,In_462,In_635);
or U1581 (N_1581,In_468,In_426);
nor U1582 (N_1582,In_534,In_730);
nor U1583 (N_1583,In_127,In_519);
and U1584 (N_1584,In_522,In_540);
and U1585 (N_1585,In_351,In_49);
nor U1586 (N_1586,In_354,In_97);
xnor U1587 (N_1587,In_62,In_51);
or U1588 (N_1588,In_389,In_314);
or U1589 (N_1589,In_539,In_69);
and U1590 (N_1590,In_638,In_191);
and U1591 (N_1591,In_442,In_376);
nor U1592 (N_1592,In_631,In_536);
and U1593 (N_1593,In_263,In_674);
nand U1594 (N_1594,In_135,In_487);
nand U1595 (N_1595,In_514,In_648);
and U1596 (N_1596,In_110,In_381);
or U1597 (N_1597,In_457,In_168);
or U1598 (N_1598,In_716,In_598);
nand U1599 (N_1599,In_437,In_36);
nor U1600 (N_1600,In_520,In_234);
or U1601 (N_1601,In_218,In_262);
or U1602 (N_1602,In_538,In_5);
nand U1603 (N_1603,In_443,In_138);
or U1604 (N_1604,In_98,In_389);
nor U1605 (N_1605,In_620,In_633);
or U1606 (N_1606,In_480,In_523);
nor U1607 (N_1607,In_727,In_746);
nor U1608 (N_1608,In_512,In_246);
nor U1609 (N_1609,In_550,In_356);
nor U1610 (N_1610,In_69,In_77);
or U1611 (N_1611,In_49,In_193);
or U1612 (N_1612,In_704,In_396);
and U1613 (N_1613,In_219,In_264);
or U1614 (N_1614,In_110,In_125);
nand U1615 (N_1615,In_169,In_249);
nor U1616 (N_1616,In_337,In_121);
or U1617 (N_1617,In_475,In_316);
nand U1618 (N_1618,In_451,In_323);
and U1619 (N_1619,In_668,In_247);
nor U1620 (N_1620,In_67,In_613);
nor U1621 (N_1621,In_372,In_480);
nor U1622 (N_1622,In_219,In_728);
nor U1623 (N_1623,In_650,In_90);
nor U1624 (N_1624,In_292,In_603);
or U1625 (N_1625,In_71,In_628);
or U1626 (N_1626,In_87,In_68);
nand U1627 (N_1627,In_495,In_137);
or U1628 (N_1628,In_644,In_255);
and U1629 (N_1629,In_193,In_323);
nor U1630 (N_1630,In_202,In_36);
or U1631 (N_1631,In_358,In_378);
nand U1632 (N_1632,In_59,In_622);
and U1633 (N_1633,In_271,In_504);
nand U1634 (N_1634,In_195,In_709);
or U1635 (N_1635,In_560,In_126);
nor U1636 (N_1636,In_348,In_213);
nor U1637 (N_1637,In_727,In_305);
and U1638 (N_1638,In_507,In_635);
nand U1639 (N_1639,In_524,In_20);
nand U1640 (N_1640,In_737,In_96);
nand U1641 (N_1641,In_419,In_198);
or U1642 (N_1642,In_294,In_377);
or U1643 (N_1643,In_259,In_734);
nand U1644 (N_1644,In_190,In_710);
or U1645 (N_1645,In_301,In_576);
nand U1646 (N_1646,In_280,In_126);
nor U1647 (N_1647,In_388,In_76);
and U1648 (N_1648,In_635,In_156);
and U1649 (N_1649,In_581,In_497);
nand U1650 (N_1650,In_604,In_467);
nand U1651 (N_1651,In_26,In_669);
nor U1652 (N_1652,In_262,In_499);
xnor U1653 (N_1653,In_400,In_259);
and U1654 (N_1654,In_376,In_734);
nand U1655 (N_1655,In_191,In_418);
and U1656 (N_1656,In_737,In_291);
nand U1657 (N_1657,In_622,In_224);
nor U1658 (N_1658,In_191,In_553);
nand U1659 (N_1659,In_628,In_577);
and U1660 (N_1660,In_588,In_333);
nand U1661 (N_1661,In_232,In_580);
or U1662 (N_1662,In_147,In_477);
nand U1663 (N_1663,In_314,In_658);
nand U1664 (N_1664,In_572,In_330);
nor U1665 (N_1665,In_25,In_434);
nand U1666 (N_1666,In_14,In_73);
or U1667 (N_1667,In_687,In_522);
or U1668 (N_1668,In_25,In_704);
nand U1669 (N_1669,In_429,In_198);
or U1670 (N_1670,In_299,In_356);
nand U1671 (N_1671,In_730,In_323);
and U1672 (N_1672,In_711,In_464);
nor U1673 (N_1673,In_690,In_434);
nand U1674 (N_1674,In_84,In_218);
or U1675 (N_1675,In_707,In_173);
nor U1676 (N_1676,In_247,In_340);
or U1677 (N_1677,In_500,In_10);
nand U1678 (N_1678,In_374,In_50);
nor U1679 (N_1679,In_285,In_623);
nor U1680 (N_1680,In_397,In_609);
nor U1681 (N_1681,In_325,In_121);
and U1682 (N_1682,In_746,In_94);
nand U1683 (N_1683,In_480,In_282);
and U1684 (N_1684,In_235,In_338);
and U1685 (N_1685,In_672,In_467);
nand U1686 (N_1686,In_357,In_748);
or U1687 (N_1687,In_142,In_365);
and U1688 (N_1688,In_517,In_351);
or U1689 (N_1689,In_626,In_703);
nor U1690 (N_1690,In_280,In_284);
or U1691 (N_1691,In_647,In_524);
and U1692 (N_1692,In_586,In_459);
and U1693 (N_1693,In_725,In_409);
nor U1694 (N_1694,In_400,In_362);
and U1695 (N_1695,In_332,In_655);
nand U1696 (N_1696,In_277,In_489);
and U1697 (N_1697,In_377,In_555);
nand U1698 (N_1698,In_404,In_629);
and U1699 (N_1699,In_577,In_328);
and U1700 (N_1700,In_549,In_356);
nand U1701 (N_1701,In_597,In_249);
and U1702 (N_1702,In_470,In_583);
and U1703 (N_1703,In_200,In_42);
nand U1704 (N_1704,In_542,In_255);
nor U1705 (N_1705,In_477,In_262);
nand U1706 (N_1706,In_585,In_559);
nor U1707 (N_1707,In_70,In_383);
nand U1708 (N_1708,In_87,In_165);
and U1709 (N_1709,In_419,In_520);
or U1710 (N_1710,In_195,In_468);
or U1711 (N_1711,In_265,In_346);
nor U1712 (N_1712,In_232,In_460);
and U1713 (N_1713,In_189,In_440);
nor U1714 (N_1714,In_451,In_740);
nor U1715 (N_1715,In_312,In_118);
nand U1716 (N_1716,In_328,In_320);
or U1717 (N_1717,In_746,In_76);
or U1718 (N_1718,In_684,In_536);
nand U1719 (N_1719,In_513,In_387);
and U1720 (N_1720,In_361,In_338);
or U1721 (N_1721,In_658,In_621);
nand U1722 (N_1722,In_232,In_594);
nor U1723 (N_1723,In_2,In_85);
nor U1724 (N_1724,In_371,In_482);
nand U1725 (N_1725,In_503,In_480);
and U1726 (N_1726,In_398,In_580);
and U1727 (N_1727,In_379,In_236);
or U1728 (N_1728,In_713,In_226);
and U1729 (N_1729,In_26,In_393);
nand U1730 (N_1730,In_207,In_247);
nor U1731 (N_1731,In_186,In_579);
or U1732 (N_1732,In_238,In_198);
nand U1733 (N_1733,In_244,In_360);
nand U1734 (N_1734,In_96,In_144);
or U1735 (N_1735,In_647,In_141);
or U1736 (N_1736,In_148,In_642);
nand U1737 (N_1737,In_263,In_613);
nor U1738 (N_1738,In_259,In_368);
and U1739 (N_1739,In_72,In_32);
or U1740 (N_1740,In_10,In_480);
nor U1741 (N_1741,In_635,In_602);
nor U1742 (N_1742,In_650,In_507);
nand U1743 (N_1743,In_378,In_101);
nor U1744 (N_1744,In_207,In_41);
and U1745 (N_1745,In_232,In_310);
and U1746 (N_1746,In_655,In_677);
and U1747 (N_1747,In_201,In_305);
and U1748 (N_1748,In_209,In_107);
xor U1749 (N_1749,In_676,In_495);
nor U1750 (N_1750,In_713,In_476);
and U1751 (N_1751,In_575,In_3);
or U1752 (N_1752,In_463,In_426);
or U1753 (N_1753,In_161,In_671);
nor U1754 (N_1754,In_189,In_475);
or U1755 (N_1755,In_328,In_172);
nor U1756 (N_1756,In_340,In_187);
nor U1757 (N_1757,In_425,In_118);
nand U1758 (N_1758,In_95,In_318);
or U1759 (N_1759,In_406,In_172);
nor U1760 (N_1760,In_251,In_499);
or U1761 (N_1761,In_58,In_224);
nand U1762 (N_1762,In_507,In_458);
and U1763 (N_1763,In_608,In_546);
nand U1764 (N_1764,In_268,In_568);
or U1765 (N_1765,In_548,In_392);
and U1766 (N_1766,In_55,In_277);
nor U1767 (N_1767,In_546,In_529);
or U1768 (N_1768,In_407,In_442);
nor U1769 (N_1769,In_62,In_616);
nand U1770 (N_1770,In_740,In_174);
and U1771 (N_1771,In_66,In_302);
and U1772 (N_1772,In_571,In_252);
nand U1773 (N_1773,In_280,In_399);
nor U1774 (N_1774,In_657,In_560);
nor U1775 (N_1775,In_124,In_453);
or U1776 (N_1776,In_222,In_324);
and U1777 (N_1777,In_267,In_378);
nor U1778 (N_1778,In_604,In_721);
nor U1779 (N_1779,In_3,In_233);
and U1780 (N_1780,In_449,In_448);
nand U1781 (N_1781,In_649,In_350);
and U1782 (N_1782,In_729,In_428);
nand U1783 (N_1783,In_493,In_510);
or U1784 (N_1784,In_662,In_539);
and U1785 (N_1785,In_68,In_361);
nand U1786 (N_1786,In_634,In_388);
nand U1787 (N_1787,In_52,In_596);
or U1788 (N_1788,In_572,In_334);
nand U1789 (N_1789,In_686,In_494);
nor U1790 (N_1790,In_627,In_612);
nor U1791 (N_1791,In_541,In_520);
and U1792 (N_1792,In_198,In_623);
and U1793 (N_1793,In_23,In_703);
and U1794 (N_1794,In_439,In_605);
nor U1795 (N_1795,In_547,In_513);
nor U1796 (N_1796,In_405,In_46);
and U1797 (N_1797,In_455,In_87);
nand U1798 (N_1798,In_710,In_592);
nand U1799 (N_1799,In_123,In_158);
nand U1800 (N_1800,In_722,In_611);
nand U1801 (N_1801,In_202,In_194);
and U1802 (N_1802,In_550,In_360);
or U1803 (N_1803,In_519,In_346);
and U1804 (N_1804,In_675,In_210);
and U1805 (N_1805,In_426,In_211);
or U1806 (N_1806,In_354,In_688);
nor U1807 (N_1807,In_432,In_566);
nand U1808 (N_1808,In_635,In_14);
or U1809 (N_1809,In_693,In_748);
or U1810 (N_1810,In_232,In_673);
nor U1811 (N_1811,In_437,In_177);
xor U1812 (N_1812,In_68,In_512);
nand U1813 (N_1813,In_633,In_531);
nor U1814 (N_1814,In_355,In_418);
and U1815 (N_1815,In_613,In_511);
or U1816 (N_1816,In_417,In_407);
and U1817 (N_1817,In_261,In_193);
xor U1818 (N_1818,In_122,In_288);
or U1819 (N_1819,In_325,In_12);
and U1820 (N_1820,In_632,In_272);
nand U1821 (N_1821,In_217,In_675);
nor U1822 (N_1822,In_426,In_209);
or U1823 (N_1823,In_98,In_346);
nor U1824 (N_1824,In_346,In_585);
nor U1825 (N_1825,In_527,In_233);
and U1826 (N_1826,In_295,In_417);
nand U1827 (N_1827,In_216,In_663);
nand U1828 (N_1828,In_628,In_461);
nand U1829 (N_1829,In_583,In_628);
nor U1830 (N_1830,In_8,In_28);
and U1831 (N_1831,In_437,In_548);
nand U1832 (N_1832,In_106,In_614);
or U1833 (N_1833,In_339,In_593);
xor U1834 (N_1834,In_122,In_600);
nand U1835 (N_1835,In_550,In_48);
nor U1836 (N_1836,In_666,In_307);
and U1837 (N_1837,In_735,In_133);
nand U1838 (N_1838,In_276,In_94);
and U1839 (N_1839,In_133,In_531);
or U1840 (N_1840,In_356,In_682);
nand U1841 (N_1841,In_328,In_39);
or U1842 (N_1842,In_14,In_296);
nor U1843 (N_1843,In_418,In_683);
nor U1844 (N_1844,In_128,In_185);
nand U1845 (N_1845,In_348,In_50);
nand U1846 (N_1846,In_85,In_748);
nand U1847 (N_1847,In_300,In_571);
or U1848 (N_1848,In_615,In_272);
nor U1849 (N_1849,In_676,In_743);
or U1850 (N_1850,In_168,In_19);
or U1851 (N_1851,In_135,In_624);
nand U1852 (N_1852,In_302,In_313);
nand U1853 (N_1853,In_32,In_534);
or U1854 (N_1854,In_547,In_368);
nor U1855 (N_1855,In_45,In_739);
or U1856 (N_1856,In_724,In_409);
and U1857 (N_1857,In_568,In_59);
nor U1858 (N_1858,In_223,In_450);
or U1859 (N_1859,In_508,In_655);
or U1860 (N_1860,In_513,In_665);
or U1861 (N_1861,In_605,In_209);
and U1862 (N_1862,In_719,In_322);
or U1863 (N_1863,In_714,In_400);
nand U1864 (N_1864,In_251,In_197);
or U1865 (N_1865,In_746,In_711);
nor U1866 (N_1866,In_656,In_341);
nor U1867 (N_1867,In_305,In_569);
or U1868 (N_1868,In_525,In_506);
or U1869 (N_1869,In_427,In_734);
nor U1870 (N_1870,In_398,In_437);
or U1871 (N_1871,In_517,In_425);
or U1872 (N_1872,In_587,In_674);
and U1873 (N_1873,In_682,In_107);
and U1874 (N_1874,In_271,In_18);
xor U1875 (N_1875,In_385,In_645);
and U1876 (N_1876,In_470,In_354);
or U1877 (N_1877,In_638,In_372);
nand U1878 (N_1878,In_183,In_155);
nor U1879 (N_1879,In_193,In_570);
nand U1880 (N_1880,In_351,In_561);
and U1881 (N_1881,In_176,In_662);
and U1882 (N_1882,In_160,In_376);
or U1883 (N_1883,In_272,In_403);
nor U1884 (N_1884,In_498,In_683);
and U1885 (N_1885,In_577,In_80);
and U1886 (N_1886,In_18,In_733);
nand U1887 (N_1887,In_537,In_685);
or U1888 (N_1888,In_460,In_589);
or U1889 (N_1889,In_343,In_595);
nand U1890 (N_1890,In_737,In_631);
xor U1891 (N_1891,In_551,In_480);
nor U1892 (N_1892,In_302,In_425);
and U1893 (N_1893,In_590,In_729);
or U1894 (N_1894,In_150,In_36);
nor U1895 (N_1895,In_458,In_558);
nand U1896 (N_1896,In_538,In_151);
nor U1897 (N_1897,In_623,In_501);
or U1898 (N_1898,In_660,In_88);
or U1899 (N_1899,In_6,In_39);
nand U1900 (N_1900,In_448,In_355);
nor U1901 (N_1901,In_53,In_324);
and U1902 (N_1902,In_319,In_713);
or U1903 (N_1903,In_380,In_387);
nor U1904 (N_1904,In_680,In_234);
or U1905 (N_1905,In_592,In_702);
or U1906 (N_1906,In_119,In_744);
and U1907 (N_1907,In_43,In_458);
nor U1908 (N_1908,In_522,In_281);
nor U1909 (N_1909,In_290,In_384);
nand U1910 (N_1910,In_288,In_121);
nand U1911 (N_1911,In_320,In_205);
nand U1912 (N_1912,In_117,In_123);
or U1913 (N_1913,In_569,In_495);
or U1914 (N_1914,In_44,In_331);
and U1915 (N_1915,In_643,In_347);
nor U1916 (N_1916,In_659,In_375);
and U1917 (N_1917,In_491,In_296);
nand U1918 (N_1918,In_632,In_177);
nor U1919 (N_1919,In_373,In_36);
nor U1920 (N_1920,In_614,In_424);
nor U1921 (N_1921,In_646,In_281);
nor U1922 (N_1922,In_134,In_524);
nor U1923 (N_1923,In_110,In_43);
nor U1924 (N_1924,In_437,In_721);
or U1925 (N_1925,In_229,In_48);
nor U1926 (N_1926,In_4,In_606);
nor U1927 (N_1927,In_477,In_614);
xnor U1928 (N_1928,In_23,In_237);
or U1929 (N_1929,In_502,In_264);
nand U1930 (N_1930,In_314,In_635);
nand U1931 (N_1931,In_382,In_450);
or U1932 (N_1932,In_327,In_177);
and U1933 (N_1933,In_446,In_615);
and U1934 (N_1934,In_298,In_49);
or U1935 (N_1935,In_624,In_210);
nor U1936 (N_1936,In_319,In_533);
nor U1937 (N_1937,In_349,In_456);
and U1938 (N_1938,In_167,In_61);
nor U1939 (N_1939,In_56,In_724);
xnor U1940 (N_1940,In_704,In_33);
nor U1941 (N_1941,In_436,In_62);
or U1942 (N_1942,In_388,In_82);
and U1943 (N_1943,In_67,In_482);
or U1944 (N_1944,In_493,In_690);
nor U1945 (N_1945,In_347,In_678);
and U1946 (N_1946,In_43,In_747);
nand U1947 (N_1947,In_154,In_535);
and U1948 (N_1948,In_378,In_106);
nand U1949 (N_1949,In_686,In_339);
and U1950 (N_1950,In_638,In_289);
or U1951 (N_1951,In_285,In_728);
nand U1952 (N_1952,In_387,In_77);
and U1953 (N_1953,In_450,In_127);
nor U1954 (N_1954,In_643,In_240);
or U1955 (N_1955,In_77,In_228);
and U1956 (N_1956,In_310,In_115);
and U1957 (N_1957,In_273,In_203);
xor U1958 (N_1958,In_700,In_228);
nand U1959 (N_1959,In_21,In_140);
nor U1960 (N_1960,In_417,In_325);
or U1961 (N_1961,In_551,In_507);
nand U1962 (N_1962,In_226,In_555);
and U1963 (N_1963,In_316,In_270);
nand U1964 (N_1964,In_622,In_498);
nor U1965 (N_1965,In_625,In_242);
and U1966 (N_1966,In_396,In_370);
and U1967 (N_1967,In_55,In_2);
and U1968 (N_1968,In_264,In_23);
nand U1969 (N_1969,In_409,In_251);
nand U1970 (N_1970,In_640,In_122);
or U1971 (N_1971,In_605,In_83);
or U1972 (N_1972,In_489,In_418);
nand U1973 (N_1973,In_488,In_663);
or U1974 (N_1974,In_385,In_436);
nor U1975 (N_1975,In_670,In_425);
or U1976 (N_1976,In_386,In_151);
and U1977 (N_1977,In_183,In_267);
nand U1978 (N_1978,In_169,In_228);
nor U1979 (N_1979,In_256,In_79);
nand U1980 (N_1980,In_34,In_343);
and U1981 (N_1981,In_366,In_587);
and U1982 (N_1982,In_147,In_96);
or U1983 (N_1983,In_13,In_437);
or U1984 (N_1984,In_638,In_336);
or U1985 (N_1985,In_266,In_434);
nor U1986 (N_1986,In_468,In_171);
nand U1987 (N_1987,In_711,In_322);
nor U1988 (N_1988,In_67,In_114);
and U1989 (N_1989,In_248,In_463);
nand U1990 (N_1990,In_374,In_160);
or U1991 (N_1991,In_579,In_484);
and U1992 (N_1992,In_252,In_483);
nor U1993 (N_1993,In_281,In_521);
and U1994 (N_1994,In_81,In_696);
or U1995 (N_1995,In_173,In_419);
nand U1996 (N_1996,In_183,In_532);
and U1997 (N_1997,In_375,In_204);
nor U1998 (N_1998,In_452,In_543);
nor U1999 (N_1999,In_723,In_115);
nor U2000 (N_2000,In_42,In_296);
and U2001 (N_2001,In_557,In_389);
nor U2002 (N_2002,In_372,In_657);
nor U2003 (N_2003,In_2,In_666);
nand U2004 (N_2004,In_14,In_675);
or U2005 (N_2005,In_382,In_84);
nand U2006 (N_2006,In_537,In_524);
nor U2007 (N_2007,In_726,In_486);
or U2008 (N_2008,In_363,In_548);
or U2009 (N_2009,In_582,In_49);
nand U2010 (N_2010,In_202,In_47);
or U2011 (N_2011,In_558,In_360);
nor U2012 (N_2012,In_485,In_280);
nand U2013 (N_2013,In_21,In_31);
or U2014 (N_2014,In_224,In_641);
nand U2015 (N_2015,In_296,In_710);
nand U2016 (N_2016,In_716,In_554);
nor U2017 (N_2017,In_569,In_422);
or U2018 (N_2018,In_223,In_154);
and U2019 (N_2019,In_149,In_80);
nand U2020 (N_2020,In_706,In_436);
nor U2021 (N_2021,In_691,In_98);
or U2022 (N_2022,In_339,In_269);
or U2023 (N_2023,In_525,In_465);
nor U2024 (N_2024,In_625,In_390);
or U2025 (N_2025,In_320,In_354);
nand U2026 (N_2026,In_230,In_413);
nor U2027 (N_2027,In_136,In_643);
nand U2028 (N_2028,In_688,In_495);
and U2029 (N_2029,In_491,In_72);
or U2030 (N_2030,In_342,In_233);
and U2031 (N_2031,In_648,In_313);
and U2032 (N_2032,In_741,In_565);
and U2033 (N_2033,In_431,In_358);
nor U2034 (N_2034,In_495,In_278);
nor U2035 (N_2035,In_237,In_129);
and U2036 (N_2036,In_579,In_328);
nand U2037 (N_2037,In_88,In_705);
and U2038 (N_2038,In_288,In_125);
or U2039 (N_2039,In_300,In_163);
and U2040 (N_2040,In_545,In_311);
nor U2041 (N_2041,In_134,In_136);
and U2042 (N_2042,In_80,In_696);
and U2043 (N_2043,In_357,In_643);
or U2044 (N_2044,In_74,In_7);
xnor U2045 (N_2045,In_510,In_342);
and U2046 (N_2046,In_326,In_61);
and U2047 (N_2047,In_330,In_612);
nand U2048 (N_2048,In_469,In_527);
nand U2049 (N_2049,In_45,In_61);
nor U2050 (N_2050,In_524,In_6);
nor U2051 (N_2051,In_19,In_12);
xnor U2052 (N_2052,In_124,In_614);
and U2053 (N_2053,In_626,In_699);
nand U2054 (N_2054,In_491,In_726);
nand U2055 (N_2055,In_401,In_92);
and U2056 (N_2056,In_597,In_667);
nor U2057 (N_2057,In_669,In_571);
or U2058 (N_2058,In_66,In_236);
or U2059 (N_2059,In_426,In_197);
nor U2060 (N_2060,In_749,In_104);
nand U2061 (N_2061,In_634,In_110);
and U2062 (N_2062,In_224,In_737);
or U2063 (N_2063,In_265,In_330);
or U2064 (N_2064,In_692,In_212);
xnor U2065 (N_2065,In_242,In_448);
and U2066 (N_2066,In_581,In_741);
or U2067 (N_2067,In_569,In_535);
nor U2068 (N_2068,In_161,In_412);
and U2069 (N_2069,In_541,In_49);
or U2070 (N_2070,In_611,In_614);
or U2071 (N_2071,In_139,In_437);
nand U2072 (N_2072,In_595,In_691);
and U2073 (N_2073,In_368,In_242);
nand U2074 (N_2074,In_197,In_357);
xor U2075 (N_2075,In_598,In_728);
nor U2076 (N_2076,In_577,In_539);
nand U2077 (N_2077,In_713,In_24);
or U2078 (N_2078,In_116,In_10);
and U2079 (N_2079,In_307,In_596);
and U2080 (N_2080,In_586,In_58);
nand U2081 (N_2081,In_424,In_194);
nand U2082 (N_2082,In_622,In_139);
nor U2083 (N_2083,In_209,In_253);
or U2084 (N_2084,In_567,In_668);
nor U2085 (N_2085,In_284,In_460);
nor U2086 (N_2086,In_696,In_487);
and U2087 (N_2087,In_220,In_22);
nand U2088 (N_2088,In_431,In_162);
or U2089 (N_2089,In_452,In_713);
nor U2090 (N_2090,In_664,In_261);
nand U2091 (N_2091,In_214,In_557);
and U2092 (N_2092,In_677,In_380);
and U2093 (N_2093,In_490,In_522);
or U2094 (N_2094,In_167,In_710);
or U2095 (N_2095,In_255,In_152);
and U2096 (N_2096,In_46,In_386);
or U2097 (N_2097,In_315,In_146);
nand U2098 (N_2098,In_247,In_725);
nor U2099 (N_2099,In_27,In_729);
and U2100 (N_2100,In_68,In_745);
and U2101 (N_2101,In_340,In_625);
or U2102 (N_2102,In_686,In_455);
nor U2103 (N_2103,In_604,In_39);
or U2104 (N_2104,In_596,In_430);
or U2105 (N_2105,In_314,In_103);
or U2106 (N_2106,In_75,In_245);
or U2107 (N_2107,In_193,In_717);
nand U2108 (N_2108,In_90,In_264);
or U2109 (N_2109,In_580,In_497);
or U2110 (N_2110,In_287,In_546);
nor U2111 (N_2111,In_226,In_719);
or U2112 (N_2112,In_443,In_650);
and U2113 (N_2113,In_99,In_249);
nand U2114 (N_2114,In_609,In_252);
or U2115 (N_2115,In_125,In_642);
nor U2116 (N_2116,In_231,In_328);
nor U2117 (N_2117,In_529,In_730);
and U2118 (N_2118,In_594,In_515);
and U2119 (N_2119,In_586,In_113);
or U2120 (N_2120,In_126,In_257);
and U2121 (N_2121,In_303,In_337);
nand U2122 (N_2122,In_145,In_739);
nand U2123 (N_2123,In_710,In_66);
or U2124 (N_2124,In_189,In_471);
and U2125 (N_2125,In_250,In_539);
xor U2126 (N_2126,In_527,In_699);
and U2127 (N_2127,In_88,In_147);
nand U2128 (N_2128,In_211,In_30);
and U2129 (N_2129,In_224,In_216);
nor U2130 (N_2130,In_266,In_570);
xnor U2131 (N_2131,In_619,In_632);
nand U2132 (N_2132,In_395,In_104);
nand U2133 (N_2133,In_412,In_411);
nand U2134 (N_2134,In_47,In_201);
and U2135 (N_2135,In_112,In_196);
nand U2136 (N_2136,In_568,In_483);
and U2137 (N_2137,In_605,In_436);
or U2138 (N_2138,In_141,In_329);
or U2139 (N_2139,In_508,In_519);
nor U2140 (N_2140,In_379,In_133);
or U2141 (N_2141,In_27,In_653);
and U2142 (N_2142,In_370,In_669);
and U2143 (N_2143,In_455,In_412);
and U2144 (N_2144,In_689,In_201);
and U2145 (N_2145,In_667,In_164);
nor U2146 (N_2146,In_119,In_234);
nand U2147 (N_2147,In_205,In_0);
nor U2148 (N_2148,In_616,In_121);
and U2149 (N_2149,In_253,In_46);
nand U2150 (N_2150,In_49,In_225);
nand U2151 (N_2151,In_657,In_215);
or U2152 (N_2152,In_711,In_545);
nand U2153 (N_2153,In_485,In_218);
and U2154 (N_2154,In_184,In_305);
nor U2155 (N_2155,In_438,In_624);
nand U2156 (N_2156,In_78,In_317);
nand U2157 (N_2157,In_207,In_98);
or U2158 (N_2158,In_389,In_307);
nand U2159 (N_2159,In_733,In_354);
or U2160 (N_2160,In_602,In_323);
and U2161 (N_2161,In_51,In_282);
nor U2162 (N_2162,In_96,In_624);
nand U2163 (N_2163,In_332,In_419);
nor U2164 (N_2164,In_207,In_551);
or U2165 (N_2165,In_613,In_453);
or U2166 (N_2166,In_61,In_39);
nor U2167 (N_2167,In_589,In_264);
and U2168 (N_2168,In_689,In_135);
or U2169 (N_2169,In_730,In_696);
nor U2170 (N_2170,In_202,In_678);
nor U2171 (N_2171,In_169,In_332);
and U2172 (N_2172,In_689,In_360);
or U2173 (N_2173,In_14,In_438);
nand U2174 (N_2174,In_392,In_33);
and U2175 (N_2175,In_248,In_9);
and U2176 (N_2176,In_132,In_627);
nand U2177 (N_2177,In_425,In_221);
and U2178 (N_2178,In_143,In_328);
nand U2179 (N_2179,In_182,In_88);
or U2180 (N_2180,In_505,In_450);
and U2181 (N_2181,In_116,In_622);
nor U2182 (N_2182,In_251,In_562);
or U2183 (N_2183,In_558,In_353);
and U2184 (N_2184,In_634,In_114);
or U2185 (N_2185,In_268,In_120);
and U2186 (N_2186,In_317,In_4);
and U2187 (N_2187,In_183,In_471);
nand U2188 (N_2188,In_249,In_704);
or U2189 (N_2189,In_346,In_343);
or U2190 (N_2190,In_732,In_514);
nor U2191 (N_2191,In_737,In_43);
nand U2192 (N_2192,In_725,In_94);
or U2193 (N_2193,In_78,In_51);
nor U2194 (N_2194,In_321,In_663);
and U2195 (N_2195,In_535,In_24);
nor U2196 (N_2196,In_319,In_597);
nand U2197 (N_2197,In_644,In_58);
or U2198 (N_2198,In_245,In_343);
nor U2199 (N_2199,In_471,In_267);
and U2200 (N_2200,In_691,In_341);
nand U2201 (N_2201,In_515,In_353);
or U2202 (N_2202,In_497,In_331);
and U2203 (N_2203,In_602,In_324);
or U2204 (N_2204,In_545,In_157);
xnor U2205 (N_2205,In_65,In_372);
nand U2206 (N_2206,In_681,In_214);
or U2207 (N_2207,In_492,In_611);
xnor U2208 (N_2208,In_160,In_593);
nand U2209 (N_2209,In_395,In_632);
and U2210 (N_2210,In_612,In_155);
and U2211 (N_2211,In_558,In_568);
and U2212 (N_2212,In_352,In_240);
and U2213 (N_2213,In_31,In_485);
nor U2214 (N_2214,In_238,In_258);
or U2215 (N_2215,In_93,In_484);
xnor U2216 (N_2216,In_180,In_0);
or U2217 (N_2217,In_80,In_635);
and U2218 (N_2218,In_632,In_63);
nand U2219 (N_2219,In_422,In_417);
nor U2220 (N_2220,In_265,In_397);
or U2221 (N_2221,In_271,In_731);
nand U2222 (N_2222,In_41,In_144);
nand U2223 (N_2223,In_37,In_640);
nand U2224 (N_2224,In_8,In_291);
nor U2225 (N_2225,In_369,In_442);
nor U2226 (N_2226,In_683,In_10);
or U2227 (N_2227,In_170,In_512);
or U2228 (N_2228,In_8,In_482);
nor U2229 (N_2229,In_665,In_85);
nor U2230 (N_2230,In_510,In_377);
nand U2231 (N_2231,In_305,In_437);
or U2232 (N_2232,In_536,In_43);
and U2233 (N_2233,In_400,In_291);
nand U2234 (N_2234,In_135,In_590);
nor U2235 (N_2235,In_420,In_65);
nor U2236 (N_2236,In_497,In_659);
nor U2237 (N_2237,In_424,In_250);
and U2238 (N_2238,In_229,In_441);
nand U2239 (N_2239,In_87,In_334);
and U2240 (N_2240,In_388,In_352);
xnor U2241 (N_2241,In_114,In_23);
nand U2242 (N_2242,In_443,In_507);
nor U2243 (N_2243,In_390,In_152);
and U2244 (N_2244,In_355,In_663);
or U2245 (N_2245,In_434,In_497);
nand U2246 (N_2246,In_627,In_348);
nor U2247 (N_2247,In_611,In_38);
nand U2248 (N_2248,In_285,In_29);
nand U2249 (N_2249,In_584,In_211);
or U2250 (N_2250,In_383,In_97);
xor U2251 (N_2251,In_679,In_135);
and U2252 (N_2252,In_130,In_257);
xnor U2253 (N_2253,In_433,In_179);
or U2254 (N_2254,In_202,In_467);
and U2255 (N_2255,In_212,In_677);
nand U2256 (N_2256,In_82,In_617);
or U2257 (N_2257,In_498,In_256);
or U2258 (N_2258,In_511,In_88);
and U2259 (N_2259,In_80,In_555);
and U2260 (N_2260,In_506,In_730);
or U2261 (N_2261,In_461,In_267);
and U2262 (N_2262,In_257,In_147);
nor U2263 (N_2263,In_80,In_436);
or U2264 (N_2264,In_666,In_649);
or U2265 (N_2265,In_95,In_298);
or U2266 (N_2266,In_84,In_702);
nor U2267 (N_2267,In_400,In_682);
nor U2268 (N_2268,In_279,In_249);
nand U2269 (N_2269,In_231,In_731);
or U2270 (N_2270,In_220,In_607);
or U2271 (N_2271,In_438,In_82);
or U2272 (N_2272,In_134,In_443);
or U2273 (N_2273,In_213,In_56);
and U2274 (N_2274,In_539,In_296);
nand U2275 (N_2275,In_618,In_153);
or U2276 (N_2276,In_163,In_38);
nor U2277 (N_2277,In_413,In_387);
nand U2278 (N_2278,In_487,In_453);
nand U2279 (N_2279,In_33,In_595);
nand U2280 (N_2280,In_69,In_416);
and U2281 (N_2281,In_526,In_279);
and U2282 (N_2282,In_545,In_424);
nor U2283 (N_2283,In_656,In_737);
and U2284 (N_2284,In_561,In_184);
and U2285 (N_2285,In_397,In_528);
or U2286 (N_2286,In_279,In_163);
xor U2287 (N_2287,In_706,In_304);
nand U2288 (N_2288,In_636,In_575);
nor U2289 (N_2289,In_336,In_431);
or U2290 (N_2290,In_373,In_252);
nor U2291 (N_2291,In_627,In_452);
or U2292 (N_2292,In_181,In_568);
or U2293 (N_2293,In_12,In_18);
nor U2294 (N_2294,In_483,In_315);
and U2295 (N_2295,In_169,In_389);
or U2296 (N_2296,In_613,In_297);
nand U2297 (N_2297,In_149,In_477);
nor U2298 (N_2298,In_16,In_719);
or U2299 (N_2299,In_283,In_478);
nor U2300 (N_2300,In_84,In_244);
nand U2301 (N_2301,In_134,In_209);
or U2302 (N_2302,In_638,In_589);
nor U2303 (N_2303,In_172,In_289);
nand U2304 (N_2304,In_687,In_689);
or U2305 (N_2305,In_173,In_444);
and U2306 (N_2306,In_712,In_333);
nor U2307 (N_2307,In_325,In_2);
and U2308 (N_2308,In_495,In_237);
or U2309 (N_2309,In_471,In_192);
or U2310 (N_2310,In_399,In_715);
nor U2311 (N_2311,In_626,In_458);
or U2312 (N_2312,In_414,In_289);
nand U2313 (N_2313,In_198,In_177);
nor U2314 (N_2314,In_653,In_315);
and U2315 (N_2315,In_190,In_504);
and U2316 (N_2316,In_533,In_242);
and U2317 (N_2317,In_80,In_502);
nor U2318 (N_2318,In_569,In_36);
nand U2319 (N_2319,In_57,In_690);
nand U2320 (N_2320,In_699,In_42);
nor U2321 (N_2321,In_511,In_492);
xor U2322 (N_2322,In_416,In_2);
or U2323 (N_2323,In_253,In_651);
nor U2324 (N_2324,In_51,In_354);
xor U2325 (N_2325,In_317,In_132);
or U2326 (N_2326,In_240,In_726);
nand U2327 (N_2327,In_217,In_578);
nor U2328 (N_2328,In_141,In_64);
or U2329 (N_2329,In_77,In_737);
and U2330 (N_2330,In_626,In_661);
or U2331 (N_2331,In_531,In_198);
or U2332 (N_2332,In_295,In_416);
nand U2333 (N_2333,In_452,In_114);
and U2334 (N_2334,In_265,In_112);
or U2335 (N_2335,In_156,In_320);
nor U2336 (N_2336,In_49,In_136);
and U2337 (N_2337,In_693,In_594);
nand U2338 (N_2338,In_372,In_169);
or U2339 (N_2339,In_567,In_135);
nor U2340 (N_2340,In_596,In_34);
nor U2341 (N_2341,In_470,In_9);
or U2342 (N_2342,In_144,In_642);
or U2343 (N_2343,In_665,In_571);
nor U2344 (N_2344,In_246,In_418);
and U2345 (N_2345,In_606,In_325);
and U2346 (N_2346,In_290,In_374);
and U2347 (N_2347,In_5,In_90);
xnor U2348 (N_2348,In_572,In_136);
nor U2349 (N_2349,In_138,In_74);
nor U2350 (N_2350,In_667,In_425);
and U2351 (N_2351,In_719,In_319);
or U2352 (N_2352,In_631,In_705);
nor U2353 (N_2353,In_194,In_286);
and U2354 (N_2354,In_684,In_191);
nand U2355 (N_2355,In_440,In_9);
nand U2356 (N_2356,In_383,In_466);
nand U2357 (N_2357,In_149,In_707);
nand U2358 (N_2358,In_71,In_261);
nor U2359 (N_2359,In_124,In_92);
xnor U2360 (N_2360,In_99,In_78);
and U2361 (N_2361,In_544,In_78);
and U2362 (N_2362,In_594,In_447);
nor U2363 (N_2363,In_497,In_535);
xor U2364 (N_2364,In_268,In_270);
and U2365 (N_2365,In_540,In_128);
nand U2366 (N_2366,In_68,In_78);
or U2367 (N_2367,In_511,In_642);
nand U2368 (N_2368,In_128,In_581);
or U2369 (N_2369,In_347,In_0);
and U2370 (N_2370,In_441,In_625);
nor U2371 (N_2371,In_154,In_610);
nand U2372 (N_2372,In_183,In_224);
nor U2373 (N_2373,In_120,In_441);
nand U2374 (N_2374,In_358,In_39);
or U2375 (N_2375,In_741,In_253);
nor U2376 (N_2376,In_699,In_690);
or U2377 (N_2377,In_314,In_330);
nand U2378 (N_2378,In_237,In_224);
nand U2379 (N_2379,In_416,In_729);
xnor U2380 (N_2380,In_496,In_101);
or U2381 (N_2381,In_71,In_430);
nand U2382 (N_2382,In_367,In_78);
and U2383 (N_2383,In_93,In_704);
nand U2384 (N_2384,In_289,In_454);
and U2385 (N_2385,In_126,In_272);
or U2386 (N_2386,In_523,In_251);
or U2387 (N_2387,In_408,In_164);
or U2388 (N_2388,In_176,In_35);
and U2389 (N_2389,In_647,In_64);
and U2390 (N_2390,In_243,In_108);
and U2391 (N_2391,In_405,In_526);
and U2392 (N_2392,In_220,In_280);
or U2393 (N_2393,In_161,In_171);
and U2394 (N_2394,In_383,In_204);
or U2395 (N_2395,In_211,In_427);
and U2396 (N_2396,In_723,In_401);
or U2397 (N_2397,In_243,In_358);
nand U2398 (N_2398,In_707,In_230);
or U2399 (N_2399,In_67,In_120);
nand U2400 (N_2400,In_627,In_74);
nand U2401 (N_2401,In_358,In_707);
and U2402 (N_2402,In_118,In_319);
and U2403 (N_2403,In_704,In_701);
and U2404 (N_2404,In_324,In_304);
and U2405 (N_2405,In_374,In_682);
or U2406 (N_2406,In_114,In_24);
nand U2407 (N_2407,In_196,In_722);
nand U2408 (N_2408,In_574,In_121);
or U2409 (N_2409,In_247,In_734);
or U2410 (N_2410,In_336,In_214);
nor U2411 (N_2411,In_474,In_539);
and U2412 (N_2412,In_360,In_246);
and U2413 (N_2413,In_332,In_456);
nor U2414 (N_2414,In_688,In_654);
nor U2415 (N_2415,In_746,In_602);
nand U2416 (N_2416,In_733,In_483);
and U2417 (N_2417,In_471,In_573);
nand U2418 (N_2418,In_386,In_45);
and U2419 (N_2419,In_165,In_260);
or U2420 (N_2420,In_69,In_403);
nand U2421 (N_2421,In_73,In_99);
or U2422 (N_2422,In_273,In_298);
nor U2423 (N_2423,In_297,In_717);
or U2424 (N_2424,In_215,In_309);
nand U2425 (N_2425,In_99,In_406);
nor U2426 (N_2426,In_302,In_218);
or U2427 (N_2427,In_596,In_443);
nand U2428 (N_2428,In_407,In_218);
and U2429 (N_2429,In_1,In_531);
nor U2430 (N_2430,In_267,In_354);
and U2431 (N_2431,In_577,In_96);
nor U2432 (N_2432,In_368,In_386);
nand U2433 (N_2433,In_705,In_568);
or U2434 (N_2434,In_706,In_98);
nor U2435 (N_2435,In_684,In_168);
nand U2436 (N_2436,In_406,In_464);
or U2437 (N_2437,In_76,In_370);
and U2438 (N_2438,In_282,In_606);
nor U2439 (N_2439,In_316,In_96);
nand U2440 (N_2440,In_260,In_4);
and U2441 (N_2441,In_35,In_172);
or U2442 (N_2442,In_607,In_667);
or U2443 (N_2443,In_653,In_257);
or U2444 (N_2444,In_507,In_665);
nand U2445 (N_2445,In_713,In_661);
and U2446 (N_2446,In_224,In_69);
nand U2447 (N_2447,In_74,In_164);
nor U2448 (N_2448,In_357,In_510);
or U2449 (N_2449,In_600,In_104);
nor U2450 (N_2450,In_43,In_92);
and U2451 (N_2451,In_589,In_584);
nand U2452 (N_2452,In_733,In_703);
and U2453 (N_2453,In_460,In_640);
or U2454 (N_2454,In_595,In_97);
nor U2455 (N_2455,In_408,In_109);
nand U2456 (N_2456,In_141,In_439);
or U2457 (N_2457,In_249,In_598);
and U2458 (N_2458,In_360,In_191);
nor U2459 (N_2459,In_291,In_110);
or U2460 (N_2460,In_301,In_551);
and U2461 (N_2461,In_372,In_739);
or U2462 (N_2462,In_360,In_89);
and U2463 (N_2463,In_21,In_542);
nor U2464 (N_2464,In_623,In_484);
nand U2465 (N_2465,In_641,In_113);
nor U2466 (N_2466,In_557,In_10);
nor U2467 (N_2467,In_61,In_639);
nand U2468 (N_2468,In_155,In_67);
nor U2469 (N_2469,In_233,In_120);
nand U2470 (N_2470,In_305,In_600);
nor U2471 (N_2471,In_433,In_326);
and U2472 (N_2472,In_470,In_571);
nor U2473 (N_2473,In_77,In_255);
and U2474 (N_2474,In_252,In_467);
nor U2475 (N_2475,In_17,In_389);
nor U2476 (N_2476,In_165,In_687);
and U2477 (N_2477,In_428,In_146);
nand U2478 (N_2478,In_184,In_644);
nor U2479 (N_2479,In_518,In_166);
and U2480 (N_2480,In_568,In_690);
nor U2481 (N_2481,In_695,In_469);
nand U2482 (N_2482,In_54,In_181);
nand U2483 (N_2483,In_327,In_31);
nand U2484 (N_2484,In_331,In_182);
or U2485 (N_2485,In_474,In_94);
or U2486 (N_2486,In_551,In_74);
nand U2487 (N_2487,In_548,In_297);
or U2488 (N_2488,In_15,In_309);
nand U2489 (N_2489,In_623,In_105);
nor U2490 (N_2490,In_486,In_332);
or U2491 (N_2491,In_153,In_115);
or U2492 (N_2492,In_708,In_119);
nand U2493 (N_2493,In_294,In_593);
or U2494 (N_2494,In_659,In_264);
or U2495 (N_2495,In_69,In_432);
and U2496 (N_2496,In_53,In_354);
or U2497 (N_2497,In_237,In_627);
and U2498 (N_2498,In_338,In_674);
and U2499 (N_2499,In_510,In_654);
nor U2500 (N_2500,N_2035,N_1733);
and U2501 (N_2501,N_742,N_779);
nand U2502 (N_2502,N_1017,N_1022);
xor U2503 (N_2503,N_2091,N_1661);
nand U2504 (N_2504,N_1204,N_1942);
nand U2505 (N_2505,N_1485,N_1548);
or U2506 (N_2506,N_2203,N_2077);
nand U2507 (N_2507,N_2134,N_1918);
and U2508 (N_2508,N_1000,N_1177);
or U2509 (N_2509,N_808,N_2308);
nor U2510 (N_2510,N_1365,N_998);
or U2511 (N_2511,N_612,N_1531);
nor U2512 (N_2512,N_1262,N_1974);
nor U2513 (N_2513,N_2194,N_1642);
or U2514 (N_2514,N_1805,N_465);
nand U2515 (N_2515,N_1307,N_928);
nor U2516 (N_2516,N_226,N_1156);
nand U2517 (N_2517,N_2000,N_127);
and U2518 (N_2518,N_90,N_851);
and U2519 (N_2519,N_1081,N_1471);
nor U2520 (N_2520,N_2206,N_64);
nand U2521 (N_2521,N_369,N_1046);
and U2522 (N_2522,N_2027,N_2098);
and U2523 (N_2523,N_2058,N_1199);
nor U2524 (N_2524,N_953,N_1764);
or U2525 (N_2525,N_221,N_1317);
or U2526 (N_2526,N_914,N_2127);
nand U2527 (N_2527,N_403,N_1804);
nand U2528 (N_2528,N_721,N_730);
nand U2529 (N_2529,N_380,N_1864);
or U2530 (N_2530,N_1814,N_1419);
nor U2531 (N_2531,N_2030,N_2217);
or U2532 (N_2532,N_151,N_1565);
and U2533 (N_2533,N_1694,N_1519);
nor U2534 (N_2534,N_659,N_315);
and U2535 (N_2535,N_1171,N_1710);
and U2536 (N_2536,N_2479,N_1477);
and U2537 (N_2537,N_655,N_1491);
and U2538 (N_2538,N_1053,N_1076);
nor U2539 (N_2539,N_2079,N_1372);
nor U2540 (N_2540,N_1023,N_2310);
or U2541 (N_2541,N_1408,N_871);
nand U2542 (N_2542,N_1225,N_1851);
nand U2543 (N_2543,N_2063,N_2270);
nor U2544 (N_2544,N_699,N_1559);
nor U2545 (N_2545,N_1265,N_115);
or U2546 (N_2546,N_430,N_2008);
or U2547 (N_2547,N_932,N_680);
and U2548 (N_2548,N_373,N_844);
nor U2549 (N_2549,N_60,N_1861);
nor U2550 (N_2550,N_378,N_2484);
xor U2551 (N_2551,N_139,N_1097);
nand U2552 (N_2552,N_2138,N_452);
nand U2553 (N_2553,N_76,N_392);
nand U2554 (N_2554,N_1673,N_459);
or U2555 (N_2555,N_2325,N_2234);
and U2556 (N_2556,N_1292,N_1042);
and U2557 (N_2557,N_2344,N_2119);
or U2558 (N_2558,N_1068,N_1459);
and U2559 (N_2559,N_1366,N_1179);
nor U2560 (N_2560,N_184,N_455);
and U2561 (N_2561,N_581,N_695);
and U2562 (N_2562,N_1065,N_2353);
or U2563 (N_2563,N_2470,N_792);
nand U2564 (N_2564,N_687,N_623);
and U2565 (N_2565,N_2297,N_747);
nor U2566 (N_2566,N_1868,N_120);
and U2567 (N_2567,N_1035,N_1810);
nor U2568 (N_2568,N_864,N_2427);
and U2569 (N_2569,N_1625,N_571);
nand U2570 (N_2570,N_1211,N_2362);
or U2571 (N_2571,N_1461,N_729);
nand U2572 (N_2572,N_239,N_400);
or U2573 (N_2573,N_1950,N_2496);
xnor U2574 (N_2574,N_2354,N_1396);
nor U2575 (N_2575,N_2,N_762);
nand U2576 (N_2576,N_838,N_1669);
and U2577 (N_2577,N_189,N_2277);
and U2578 (N_2578,N_652,N_2154);
or U2579 (N_2579,N_1062,N_18);
nand U2580 (N_2580,N_19,N_794);
nand U2581 (N_2581,N_1364,N_1321);
nand U2582 (N_2582,N_944,N_70);
nand U2583 (N_2583,N_304,N_519);
nand U2584 (N_2584,N_546,N_2378);
nand U2585 (N_2585,N_2117,N_5);
nor U2586 (N_2586,N_2320,N_147);
and U2587 (N_2587,N_1487,N_67);
or U2588 (N_2588,N_183,N_422);
nor U2589 (N_2589,N_1128,N_795);
nand U2590 (N_2590,N_2491,N_807);
or U2591 (N_2591,N_1351,N_2057);
and U2592 (N_2592,N_446,N_566);
nand U2593 (N_2593,N_520,N_2005);
nand U2594 (N_2594,N_1412,N_1938);
and U2595 (N_2595,N_2169,N_717);
and U2596 (N_2596,N_1391,N_1212);
or U2597 (N_2597,N_1497,N_2156);
nand U2598 (N_2598,N_752,N_621);
nand U2599 (N_2599,N_1650,N_1976);
nand U2600 (N_2600,N_2246,N_2275);
or U2601 (N_2601,N_1045,N_309);
and U2602 (N_2602,N_1582,N_278);
nor U2603 (N_2603,N_957,N_1560);
nor U2604 (N_2604,N_1369,N_2348);
nand U2605 (N_2605,N_899,N_763);
nand U2606 (N_2606,N_178,N_2139);
nand U2607 (N_2607,N_122,N_2120);
or U2608 (N_2608,N_1618,N_2274);
or U2609 (N_2609,N_166,N_1812);
or U2610 (N_2610,N_274,N_2421);
or U2611 (N_2611,N_534,N_31);
nor U2612 (N_2612,N_1198,N_2490);
nand U2613 (N_2613,N_934,N_1755);
and U2614 (N_2614,N_1882,N_1374);
and U2615 (N_2615,N_2214,N_2272);
nor U2616 (N_2616,N_1756,N_1239);
nand U2617 (N_2617,N_1324,N_1168);
or U2618 (N_2618,N_2341,N_2021);
or U2619 (N_2619,N_1146,N_170);
nand U2620 (N_2620,N_1305,N_1186);
and U2621 (N_2621,N_2465,N_2413);
and U2622 (N_2622,N_1534,N_2279);
and U2623 (N_2623,N_2287,N_219);
and U2624 (N_2624,N_458,N_992);
and U2625 (N_2625,N_1278,N_1542);
or U2626 (N_2626,N_1946,N_2480);
nor U2627 (N_2627,N_856,N_2438);
or U2628 (N_2628,N_467,N_1201);
nor U2629 (N_2629,N_2195,N_37);
nand U2630 (N_2630,N_440,N_1009);
nor U2631 (N_2631,N_884,N_2369);
or U2632 (N_2632,N_319,N_2104);
nand U2633 (N_2633,N_2386,N_1348);
or U2634 (N_2634,N_694,N_310);
and U2635 (N_2635,N_135,N_999);
nor U2636 (N_2636,N_2249,N_1993);
or U2637 (N_2637,N_1909,N_2061);
nand U2638 (N_2638,N_16,N_1453);
nand U2639 (N_2639,N_2345,N_575);
nand U2640 (N_2640,N_1706,N_404);
and U2641 (N_2641,N_1313,N_266);
nor U2642 (N_2642,N_574,N_216);
nor U2643 (N_2643,N_771,N_1202);
nand U2644 (N_2644,N_1149,N_732);
nor U2645 (N_2645,N_2442,N_751);
and U2646 (N_2646,N_890,N_1256);
nand U2647 (N_2647,N_665,N_2226);
and U2648 (N_2648,N_937,N_2422);
nand U2649 (N_2649,N_114,N_2242);
or U2650 (N_2650,N_2135,N_1871);
and U2651 (N_2651,N_2307,N_287);
nand U2652 (N_2652,N_2295,N_1914);
nand U2653 (N_2653,N_1210,N_1008);
nand U2654 (N_2654,N_1304,N_333);
nand U2655 (N_2655,N_1511,N_949);
nand U2656 (N_2656,N_1589,N_273);
or U2657 (N_2657,N_619,N_200);
nor U2658 (N_2658,N_74,N_736);
xor U2659 (N_2659,N_1218,N_1912);
and U2660 (N_2660,N_470,N_1306);
nand U2661 (N_2661,N_1230,N_1486);
or U2662 (N_2662,N_965,N_669);
or U2663 (N_2663,N_568,N_1352);
or U2664 (N_2664,N_1482,N_1344);
or U2665 (N_2665,N_785,N_714);
nand U2666 (N_2666,N_1513,N_223);
and U2667 (N_2667,N_1298,N_414);
and U2668 (N_2668,N_1085,N_1508);
nand U2669 (N_2669,N_2164,N_169);
or U2670 (N_2670,N_161,N_285);
nor U2671 (N_2671,N_2253,N_2048);
or U2672 (N_2672,N_1113,N_107);
or U2673 (N_2673,N_2073,N_1613);
or U2674 (N_2674,N_155,N_1088);
nand U2675 (N_2675,N_1853,N_2471);
or U2676 (N_2676,N_1049,N_2261);
and U2677 (N_2677,N_1931,N_1879);
and U2678 (N_2678,N_1108,N_224);
nor U2679 (N_2679,N_1677,N_53);
or U2680 (N_2680,N_1185,N_2283);
nor U2681 (N_2681,N_1796,N_1852);
nor U2682 (N_2682,N_335,N_2290);
nand U2683 (N_2683,N_1518,N_782);
nor U2684 (N_2684,N_1243,N_1702);
and U2685 (N_2685,N_2267,N_739);
nand U2686 (N_2686,N_1099,N_875);
nand U2687 (N_2687,N_14,N_225);
and U2688 (N_2688,N_1908,N_723);
or U2689 (N_2689,N_1176,N_1446);
nand U2690 (N_2690,N_1464,N_1577);
nor U2691 (N_2691,N_1060,N_1214);
and U2692 (N_2692,N_2399,N_2131);
or U2693 (N_2693,N_1536,N_1789);
or U2694 (N_2694,N_398,N_1147);
and U2695 (N_2695,N_28,N_69);
nand U2696 (N_2696,N_578,N_1215);
and U2697 (N_2697,N_1300,N_1194);
or U2698 (N_2698,N_206,N_1255);
and U2699 (N_2699,N_447,N_502);
nor U2700 (N_2700,N_2163,N_1945);
nor U2701 (N_2701,N_2266,N_840);
and U2702 (N_2702,N_1737,N_1140);
nand U2703 (N_2703,N_2312,N_1657);
nor U2704 (N_2704,N_437,N_491);
or U2705 (N_2705,N_1430,N_1303);
nor U2706 (N_2706,N_1203,N_2268);
nand U2707 (N_2707,N_2288,N_952);
and U2708 (N_2708,N_1449,N_1285);
nor U2709 (N_2709,N_2296,N_2282);
nor U2710 (N_2710,N_765,N_203);
or U2711 (N_2711,N_306,N_343);
nand U2712 (N_2712,N_2271,N_1037);
nor U2713 (N_2713,N_1987,N_126);
or U2714 (N_2714,N_783,N_49);
nand U2715 (N_2715,N_980,N_1696);
nor U2716 (N_2716,N_997,N_1570);
and U2717 (N_2717,N_1715,N_2196);
nand U2718 (N_2718,N_462,N_2410);
and U2719 (N_2719,N_1318,N_2055);
nor U2720 (N_2720,N_681,N_1824);
nor U2721 (N_2721,N_754,N_1493);
and U2722 (N_2722,N_1898,N_716);
and U2723 (N_2723,N_2276,N_2435);
nand U2724 (N_2724,N_187,N_961);
nand U2725 (N_2725,N_1213,N_1728);
nand U2726 (N_2726,N_466,N_208);
and U2727 (N_2727,N_331,N_393);
and U2728 (N_2728,N_603,N_1547);
or U2729 (N_2729,N_173,N_889);
nand U2730 (N_2730,N_1221,N_51);
and U2731 (N_2731,N_2425,N_507);
or U2732 (N_2732,N_1995,N_1415);
or U2733 (N_2733,N_2467,N_2199);
or U2734 (N_2734,N_560,N_407);
nor U2735 (N_2735,N_84,N_1837);
nor U2736 (N_2736,N_2423,N_1356);
nand U2737 (N_2737,N_58,N_4);
nand U2738 (N_2738,N_711,N_2444);
or U2739 (N_2739,N_2106,N_313);
and U2740 (N_2740,N_325,N_715);
and U2741 (N_2741,N_371,N_872);
or U2742 (N_2742,N_210,N_1746);
or U2743 (N_2743,N_709,N_2319);
and U2744 (N_2744,N_1601,N_1575);
and U2745 (N_2745,N_833,N_1674);
nand U2746 (N_2746,N_246,N_731);
or U2747 (N_2747,N_235,N_2034);
nand U2748 (N_2748,N_826,N_1709);
nand U2749 (N_2749,N_2437,N_1752);
nand U2750 (N_2750,N_190,N_2094);
or U2751 (N_2751,N_1116,N_2291);
nand U2752 (N_2752,N_2250,N_260);
nand U2753 (N_2753,N_1970,N_1659);
or U2754 (N_2754,N_234,N_1118);
nor U2755 (N_2755,N_2218,N_2004);
nand U2756 (N_2756,N_958,N_1041);
or U2757 (N_2757,N_175,N_913);
nand U2758 (N_2758,N_2232,N_734);
or U2759 (N_2759,N_968,N_1001);
or U2760 (N_2760,N_148,N_1635);
xnor U2761 (N_2761,N_516,N_1828);
or U2762 (N_2762,N_2356,N_453);
nor U2763 (N_2763,N_1167,N_1533);
and U2764 (N_2764,N_1546,N_1341);
nor U2765 (N_2765,N_790,N_2492);
nand U2766 (N_2766,N_1863,N_286);
nor U2767 (N_2767,N_117,N_391);
nor U2768 (N_2768,N_1539,N_2498);
nand U2769 (N_2769,N_485,N_249);
nor U2770 (N_2770,N_355,N_2204);
and U2771 (N_2771,N_172,N_891);
nand U2772 (N_2772,N_1893,N_803);
nor U2773 (N_2773,N_2280,N_1421);
nor U2774 (N_2774,N_1978,N_701);
or U2775 (N_2775,N_1857,N_1878);
nand U2776 (N_2776,N_129,N_128);
or U2777 (N_2777,N_909,N_1721);
and U2778 (N_2778,N_912,N_1526);
or U2779 (N_2779,N_1345,N_1339);
or U2780 (N_2780,N_666,N_1250);
nor U2781 (N_2781,N_387,N_1242);
xor U2782 (N_2782,N_558,N_859);
or U2783 (N_2783,N_2269,N_352);
and U2784 (N_2784,N_1792,N_2306);
or U2785 (N_2785,N_56,N_1395);
and U2786 (N_2786,N_1791,N_641);
nand U2787 (N_2787,N_908,N_1059);
nand U2788 (N_2788,N_198,N_1111);
nand U2789 (N_2789,N_1585,N_229);
xor U2790 (N_2790,N_2334,N_451);
and U2791 (N_2791,N_1916,N_57);
nor U2792 (N_2792,N_479,N_945);
or U2793 (N_2793,N_760,N_1667);
or U2794 (N_2794,N_1957,N_631);
or U2795 (N_2795,N_743,N_1478);
xor U2796 (N_2796,N_1438,N_1398);
nand U2797 (N_2797,N_1574,N_2256);
nand U2798 (N_2798,N_1774,N_113);
or U2799 (N_2799,N_825,N_674);
nand U2800 (N_2800,N_1802,N_1907);
nor U2801 (N_2801,N_543,N_2301);
nand U2802 (N_2802,N_2247,N_599);
or U2803 (N_2803,N_1143,N_71);
nand U2804 (N_2804,N_1921,N_1722);
and U2805 (N_2805,N_1846,N_679);
and U2806 (N_2806,N_1170,N_1377);
nor U2807 (N_2807,N_1785,N_116);
nand U2808 (N_2808,N_1034,N_1953);
nor U2809 (N_2809,N_529,N_1161);
or U2810 (N_2810,N_2244,N_2191);
nand U2811 (N_2811,N_2285,N_513);
or U2812 (N_2812,N_684,N_326);
or U2813 (N_2813,N_98,N_106);
and U2814 (N_2814,N_1284,N_1514);
or U2815 (N_2815,N_737,N_887);
nand U2816 (N_2816,N_1102,N_1675);
and U2817 (N_2817,N_1549,N_1460);
xnor U2818 (N_2818,N_2110,N_522);
or U2819 (N_2819,N_237,N_528);
or U2820 (N_2820,N_580,N_539);
nor U2821 (N_2821,N_1819,N_2023);
nand U2822 (N_2822,N_920,N_1189);
nor U2823 (N_2823,N_531,N_441);
nand U2824 (N_2824,N_1747,N_435);
or U2825 (N_2825,N_2182,N_1279);
nor U2826 (N_2826,N_1855,N_654);
and U2827 (N_2827,N_846,N_1763);
nand U2828 (N_2828,N_1287,N_2177);
nor U2829 (N_2829,N_2248,N_881);
or U2830 (N_2830,N_2109,N_259);
or U2831 (N_2831,N_308,N_2017);
nand U2832 (N_2832,N_1586,N_1556);
and U2833 (N_2833,N_1439,N_445);
or U2834 (N_2834,N_395,N_2001);
nor U2835 (N_2835,N_2443,N_426);
nand U2836 (N_2836,N_2167,N_1952);
nand U2837 (N_2837,N_570,N_1761);
nand U2838 (N_2838,N_2309,N_1012);
or U2839 (N_2839,N_427,N_2188);
nor U2840 (N_2840,N_500,N_2014);
and U2841 (N_2841,N_1823,N_2144);
and U2842 (N_2842,N_1644,N_1492);
and U2843 (N_2843,N_1749,N_1688);
nor U2844 (N_2844,N_2497,N_1768);
or U2845 (N_2845,N_2045,N_1915);
nor U2846 (N_2846,N_2153,N_630);
and U2847 (N_2847,N_1136,N_1454);
nor U2848 (N_2848,N_2458,N_1757);
nand U2849 (N_2849,N_1293,N_2180);
nand U2850 (N_2850,N_2054,N_1616);
and U2851 (N_2851,N_201,N_1386);
and U2852 (N_2852,N_617,N_1106);
or U2853 (N_2853,N_29,N_1748);
and U2854 (N_2854,N_828,N_2033);
nand U2855 (N_2855,N_1399,N_1891);
or U2856 (N_2856,N_359,N_1164);
nand U2857 (N_2857,N_586,N_2405);
nand U2858 (N_2858,N_2389,N_941);
nor U2859 (N_2859,N_270,N_608);
or U2860 (N_2860,N_2221,N_1150);
and U2861 (N_2861,N_1063,N_984);
or U2862 (N_2862,N_2192,N_349);
nor U2863 (N_2863,N_1251,N_152);
and U2864 (N_2864,N_2365,N_1444);
or U2865 (N_2865,N_2315,N_1154);
nand U2866 (N_2866,N_1571,N_653);
nor U2867 (N_2867,N_88,N_2383);
xnor U2868 (N_2868,N_2464,N_1397);
nor U2869 (N_2869,N_950,N_2474);
nor U2870 (N_2870,N_2255,N_1922);
and U2871 (N_2871,N_448,N_1114);
and U2872 (N_2872,N_428,N_2254);
and U2873 (N_2873,N_1658,N_1940);
nand U2874 (N_2874,N_9,N_425);
and U2875 (N_2875,N_677,N_801);
and U2876 (N_2876,N_2097,N_1173);
nor U2877 (N_2877,N_1456,N_1959);
and U2878 (N_2878,N_1742,N_837);
nand U2879 (N_2879,N_1363,N_640);
or U2880 (N_2880,N_17,N_1992);
or U2881 (N_2881,N_690,N_2032);
or U2882 (N_2882,N_2259,N_741);
or U2883 (N_2883,N_15,N_423);
and U2884 (N_2884,N_1594,N_2174);
and U2885 (N_2885,N_2468,N_2323);
nand U2886 (N_2886,N_1765,N_275);
nor U2887 (N_2887,N_2379,N_1902);
and U2888 (N_2888,N_2324,N_1236);
or U2889 (N_2889,N_1445,N_2116);
and U2890 (N_2890,N_1268,N_2143);
and U2891 (N_2891,N_493,N_2393);
and U2892 (N_2892,N_1754,N_664);
or U2893 (N_2893,N_774,N_1316);
nor U2894 (N_2894,N_1467,N_2078);
nor U2895 (N_2895,N_244,N_2476);
nor U2896 (N_2896,N_2111,N_1196);
nand U2897 (N_2897,N_1540,N_2210);
and U2898 (N_2898,N_1528,N_670);
and U2899 (N_2899,N_1943,N_988);
nand U2900 (N_2900,N_1676,N_2229);
xor U2901 (N_2901,N_499,N_2463);
or U2902 (N_2902,N_873,N_409);
nand U2903 (N_2903,N_1649,N_1271);
nor U2904 (N_2904,N_697,N_27);
or U2905 (N_2905,N_854,N_550);
or U2906 (N_2906,N_2322,N_990);
nand U2907 (N_2907,N_993,N_924);
nand U2908 (N_2908,N_689,N_726);
or U2909 (N_2909,N_150,N_1044);
xor U2910 (N_2910,N_1554,N_2370);
nor U2911 (N_2911,N_1101,N_2408);
or U2912 (N_2912,N_1580,N_457);
or U2913 (N_2913,N_177,N_501);
or U2914 (N_2914,N_962,N_727);
nand U2915 (N_2915,N_514,N_291);
nand U2916 (N_2916,N_394,N_1414);
and U2917 (N_2917,N_1431,N_1277);
and U2918 (N_2918,N_607,N_1608);
nor U2919 (N_2919,N_787,N_1329);
nor U2920 (N_2920,N_1323,N_816);
nand U2921 (N_2921,N_1342,N_518);
or U2922 (N_2922,N_613,N_2342);
nor U2923 (N_2923,N_158,N_673);
or U2924 (N_2924,N_853,N_2209);
nand U2925 (N_2925,N_1087,N_938);
and U2926 (N_2926,N_1355,N_1772);
and U2927 (N_2927,N_1744,N_929);
and U2928 (N_2928,N_1520,N_554);
and U2929 (N_2929,N_1964,N_1730);
or U2930 (N_2930,N_830,N_1672);
and U2931 (N_2931,N_1564,N_1848);
or U2932 (N_2932,N_1979,N_2241);
and U2933 (N_2933,N_1260,N_1032);
or U2934 (N_2934,N_1014,N_2022);
and U2935 (N_2935,N_1603,N_939);
nor U2936 (N_2936,N_1235,N_1296);
nand U2937 (N_2937,N_1172,N_2071);
or U2938 (N_2938,N_10,N_363);
nand U2939 (N_2939,N_2380,N_1423);
nor U2940 (N_2940,N_1019,N_777);
nand U2941 (N_2941,N_2317,N_632);
nand U2942 (N_2942,N_1226,N_2440);
or U2943 (N_2943,N_2028,N_1027);
nor U2944 (N_2944,N_1731,N_2049);
nand U2945 (N_2945,N_1311,N_2136);
and U2946 (N_2946,N_1617,N_649);
and U2947 (N_2947,N_1003,N_2065);
nor U2948 (N_2948,N_211,N_975);
or U2949 (N_2949,N_524,N_1400);
nor U2950 (N_2950,N_671,N_1832);
nor U2951 (N_2951,N_906,N_2327);
nand U2952 (N_2952,N_1484,N_1054);
nand U2953 (N_2953,N_271,N_587);
or U2954 (N_2954,N_643,N_2239);
or U2955 (N_2955,N_512,N_138);
and U2956 (N_2956,N_776,N_1894);
xor U2957 (N_2957,N_645,N_1205);
and U2958 (N_2958,N_2260,N_1822);
nor U2959 (N_2959,N_1025,N_1157);
nor U2960 (N_2960,N_1346,N_1130);
nand U2961 (N_2961,N_2299,N_1495);
or U2962 (N_2962,N_2070,N_2103);
nand U2963 (N_2963,N_324,N_1117);
nand U2964 (N_2964,N_2371,N_1083);
nor U2965 (N_2965,N_1077,N_861);
nor U2966 (N_2966,N_280,N_2355);
nand U2967 (N_2967,N_439,N_367);
nor U2968 (N_2968,N_26,N_1407);
or U2969 (N_2969,N_2224,N_1634);
nor U2970 (N_2970,N_537,N_842);
and U2971 (N_2971,N_231,N_517);
or U2972 (N_2972,N_1184,N_1375);
and U2973 (N_2973,N_136,N_12);
nand U2974 (N_2974,N_1900,N_540);
and U2975 (N_2975,N_417,N_2251);
nor U2976 (N_2976,N_1443,N_1666);
nor U2977 (N_2977,N_1434,N_2385);
or U2978 (N_2978,N_511,N_882);
xnor U2979 (N_2979,N_637,N_2024);
nand U2980 (N_2980,N_1137,N_1138);
nand U2981 (N_2981,N_1240,N_691);
or U2982 (N_2982,N_969,N_636);
nor U2983 (N_2983,N_443,N_2346);
nand U2984 (N_2984,N_207,N_1052);
nor U2985 (N_2985,N_946,N_2457);
nor U2986 (N_2986,N_1858,N_1602);
nand U2987 (N_2987,N_2446,N_1558);
nand U2988 (N_2988,N_1680,N_305);
nor U2989 (N_2989,N_2085,N_1562);
nor U2990 (N_2990,N_2363,N_1120);
nor U2991 (N_2991,N_1839,N_2434);
and U2992 (N_2992,N_1927,N_769);
nor U2993 (N_2993,N_0,N_2121);
and U2994 (N_2994,N_1773,N_415);
nor U2995 (N_2995,N_433,N_1521);
nand U2996 (N_2996,N_2012,N_66);
and U2997 (N_2997,N_806,N_1159);
xnor U2998 (N_2998,N_1084,N_1537);
nor U2999 (N_2999,N_2060,N_1835);
or U3000 (N_3000,N_954,N_788);
nor U3001 (N_3001,N_1849,N_960);
nand U3002 (N_3002,N_2436,N_2125);
and U3003 (N_3003,N_284,N_916);
nand U3004 (N_3004,N_888,N_1280);
nand U3005 (N_3005,N_490,N_1093);
or U3006 (N_3006,N_294,N_1217);
nand U3007 (N_3007,N_103,N_1751);
and U3008 (N_3008,N_756,N_109);
nor U3009 (N_3009,N_967,N_989);
nor U3010 (N_3010,N_1998,N_1187);
or U3011 (N_3011,N_1289,N_1647);
or U3012 (N_3012,N_2108,N_898);
and U3013 (N_3013,N_46,N_921);
or U3014 (N_3014,N_2102,N_277);
or U3015 (N_3015,N_1402,N_281);
nor U3016 (N_3016,N_434,N_1178);
nor U3017 (N_3017,N_2200,N_2157);
and U3018 (N_3018,N_1104,N_827);
or U3019 (N_3019,N_633,N_1843);
or U3020 (N_3020,N_2066,N_356);
or U3021 (N_3021,N_2489,N_44);
nor U3022 (N_3022,N_1836,N_710);
nor U3023 (N_3023,N_365,N_2473);
and U3024 (N_3024,N_1247,N_2416);
and U3025 (N_3025,N_923,N_693);
nand U3026 (N_3026,N_2373,N_1145);
or U3027 (N_3027,N_866,N_1462);
and U3028 (N_3028,N_2316,N_2168);
or U3029 (N_3029,N_1328,N_1132);
nor U3030 (N_3030,N_209,N_296);
nand U3031 (N_3031,N_1646,N_896);
nand U3032 (N_3032,N_1831,N_2185);
xor U3033 (N_3033,N_94,N_1566);
or U3034 (N_3034,N_2140,N_1030);
nor U3035 (N_3035,N_903,N_1246);
and U3036 (N_3036,N_1457,N_597);
or U3037 (N_3037,N_885,N_1762);
nor U3038 (N_3038,N_13,N_1779);
or U3039 (N_3039,N_344,N_1631);
nand U3040 (N_3040,N_2340,N_1686);
or U3041 (N_3041,N_629,N_241);
nor U3042 (N_3042,N_1692,N_1623);
xnor U3043 (N_3043,N_1568,N_1840);
nor U3044 (N_3044,N_1472,N_1904);
and U3045 (N_3045,N_591,N_2088);
or U3046 (N_3046,N_484,N_657);
and U3047 (N_3047,N_1379,N_1219);
nor U3048 (N_3048,N_994,N_180);
or U3049 (N_3049,N_222,N_215);
or U3050 (N_3050,N_1640,N_548);
nor U3051 (N_3051,N_402,N_2313);
and U3052 (N_3052,N_559,N_978);
or U3053 (N_3053,N_1689,N_567);
nor U3054 (N_3054,N_65,N_11);
nand U3055 (N_3055,N_660,N_541);
and U3056 (N_3056,N_25,N_974);
or U3057 (N_3057,N_1801,N_2150);
nor U3058 (N_3058,N_411,N_2100);
nor U3059 (N_3059,N_2284,N_2069);
or U3060 (N_3060,N_667,N_1958);
nor U3061 (N_3061,N_1227,N_1335);
nand U3062 (N_3062,N_1082,N_2430);
or U3063 (N_3063,N_2096,N_809);
and U3064 (N_3064,N_1643,N_883);
and U3065 (N_3065,N_2335,N_2074);
nand U3066 (N_3066,N_1139,N_1523);
or U3067 (N_3067,N_1162,N_1195);
nand U3068 (N_3068,N_1869,N_54);
nand U3069 (N_3069,N_1725,N_1126);
or U3070 (N_3070,N_746,N_647);
or U3071 (N_3071,N_1133,N_89);
or U3072 (N_3072,N_656,N_1770);
and U3073 (N_3073,N_1451,N_41);
nor U3074 (N_3074,N_1270,N_572);
or U3075 (N_3075,N_1687,N_1413);
nor U3076 (N_3076,N_1693,N_1877);
and U3077 (N_3077,N_1955,N_959);
and U3078 (N_3078,N_703,N_1645);
or U3079 (N_3079,N_1516,N_2238);
nand U3080 (N_3080,N_341,N_893);
and U3081 (N_3081,N_243,N_1781);
or U3082 (N_3082,N_579,N_2148);
or U3083 (N_3083,N_1653,N_1237);
or U3084 (N_3084,N_1919,N_922);
or U3085 (N_3085,N_753,N_1923);
or U3086 (N_3086,N_1652,N_1109);
nand U3087 (N_3087,N_220,N_386);
nor U3088 (N_3088,N_1127,N_644);
nor U3089 (N_3089,N_1967,N_1895);
nor U3090 (N_3090,N_1018,N_2113);
and U3091 (N_3091,N_1639,N_1986);
nand U3092 (N_3092,N_1411,N_1174);
and U3093 (N_3093,N_1338,N_2231);
nor U3094 (N_3094,N_2447,N_2172);
nand U3095 (N_3095,N_1929,N_1718);
nor U3096 (N_3096,N_1690,N_1392);
or U3097 (N_3097,N_1538,N_1257);
xnor U3098 (N_3098,N_263,N_1954);
nor U3099 (N_3099,N_1678,N_347);
or U3100 (N_3100,N_351,N_1142);
nand U3101 (N_3101,N_2126,N_1119);
or U3102 (N_3102,N_2456,N_1947);
nor U3103 (N_3103,N_1975,N_2429);
nor U3104 (N_3104,N_81,N_545);
and U3105 (N_3105,N_1830,N_719);
nand U3106 (N_3106,N_1036,N_2377);
nor U3107 (N_3107,N_880,N_1224);
and U3108 (N_3108,N_1253,N_2162);
or U3109 (N_3109,N_910,N_1778);
nor U3110 (N_3110,N_460,N_1665);
nor U3111 (N_3111,N_904,N_1825);
nor U3112 (N_3112,N_1557,N_101);
nor U3113 (N_3113,N_1681,N_86);
nand U3114 (N_3114,N_1319,N_804);
nor U3115 (N_3115,N_892,N_2129);
and U3116 (N_3116,N_544,N_1357);
or U3117 (N_3117,N_1656,N_2486);
nor U3118 (N_3118,N_1982,N_1498);
or U3119 (N_3119,N_1435,N_1481);
nor U3120 (N_3120,N_1021,N_1604);
and U3121 (N_3121,N_824,N_2459);
and U3122 (N_3122,N_1735,N_1005);
nor U3123 (N_3123,N_966,N_1787);
nand U3124 (N_3124,N_2382,N_1913);
and U3125 (N_3125,N_1527,N_2026);
nand U3126 (N_3126,N_1409,N_2499);
and U3127 (N_3127,N_2469,N_1719);
nor U3128 (N_3128,N_1269,N_7);
or U3129 (N_3129,N_800,N_886);
nor U3130 (N_3130,N_565,N_764);
nand U3131 (N_3131,N_1968,N_1884);
nor U3132 (N_3132,N_174,N_2205);
nand U3133 (N_3133,N_1888,N_111);
or U3134 (N_3134,N_2064,N_2417);
or U3135 (N_3135,N_661,N_272);
or U3136 (N_3136,N_1977,N_2009);
nor U3137 (N_3137,N_628,N_1865);
and U3138 (N_3138,N_1784,N_2332);
and U3139 (N_3139,N_2123,N_1026);
and U3140 (N_3140,N_1070,N_1885);
or U3141 (N_3141,N_770,N_685);
and U3142 (N_3142,N_228,N_1160);
and U3143 (N_3143,N_812,N_102);
and U3144 (N_3144,N_668,N_142);
nor U3145 (N_3145,N_1960,N_1295);
or U3146 (N_3146,N_2197,N_1881);
nand U3147 (N_3147,N_706,N_2132);
or U3148 (N_3148,N_230,N_1932);
or U3149 (N_3149,N_2453,N_382);
or U3150 (N_3150,N_21,N_1833);
and U3151 (N_3151,N_2003,N_1309);
and U3152 (N_3152,N_2056,N_2047);
or U3153 (N_3153,N_925,N_1743);
or U3154 (N_3154,N_2240,N_733);
nor U3155 (N_3155,N_100,N_1264);
nor U3156 (N_3156,N_1314,N_1510);
or U3157 (N_3157,N_2015,N_2493);
and U3158 (N_3158,N_2043,N_829);
nand U3159 (N_3159,N_317,N_482);
or U3160 (N_3160,N_1552,N_2178);
or U3161 (N_3161,N_469,N_1803);
and U3162 (N_3162,N_553,N_1624);
nor U3163 (N_3163,N_2477,N_564);
nand U3164 (N_3164,N_1595,N_879);
nand U3165 (N_3165,N_1800,N_329);
nor U3166 (N_3166,N_683,N_345);
nor U3167 (N_3167,N_1630,N_1734);
nor U3168 (N_3168,N_1874,N_639);
and U3169 (N_3169,N_2173,N_1254);
or U3170 (N_3170,N_1432,N_204);
nor U3171 (N_3171,N_1697,N_1965);
nand U3172 (N_3172,N_2412,N_2114);
xor U3173 (N_3173,N_2245,N_238);
nand U3174 (N_3174,N_334,N_2392);
and U3175 (N_3175,N_1131,N_533);
and U3176 (N_3176,N_1880,N_682);
or U3177 (N_3177,N_1427,N_1067);
and U3178 (N_3178,N_497,N_802);
and U3179 (N_3179,N_1206,N_354);
nand U3180 (N_3180,N_817,N_1302);
and U3181 (N_3181,N_124,N_255);
nand U3182 (N_3182,N_1726,N_104);
or U3183 (N_3183,N_551,N_2038);
nand U3184 (N_3184,N_948,N_312);
or U3185 (N_3185,N_1222,N_268);
and U3186 (N_3186,N_1561,N_2390);
nor U3187 (N_3187,N_964,N_449);
and U3188 (N_3188,N_2146,N_562);
and U3189 (N_3189,N_55,N_410);
nand U3190 (N_3190,N_1197,N_860);
nor U3191 (N_3191,N_2462,N_379);
nor U3192 (N_3192,N_542,N_1820);
nor U3193 (N_3193,N_2011,N_374);
and U3194 (N_3194,N_444,N_253);
nand U3195 (N_3195,N_463,N_390);
nor U3196 (N_3196,N_602,N_905);
or U3197 (N_3197,N_563,N_1286);
nand U3198 (N_3198,N_2040,N_620);
nor U3199 (N_3199,N_527,N_2328);
nand U3200 (N_3200,N_573,N_595);
or U3201 (N_3201,N_1576,N_1739);
nor U3202 (N_3202,N_2031,N_2292);
or U3203 (N_3203,N_1758,N_987);
and U3204 (N_3204,N_1827,N_577);
nor U3205 (N_3205,N_2432,N_2395);
or U3206 (N_3206,N_381,N_1337);
nand U3207 (N_3207,N_1961,N_1079);
nor U3208 (N_3208,N_845,N_1591);
nor U3209 (N_3209,N_168,N_2130);
and U3210 (N_3210,N_1169,N_2142);
and U3211 (N_3211,N_614,N_865);
or U3212 (N_3212,N_2020,N_610);
nor U3213 (N_3213,N_1682,N_194);
and U3214 (N_3214,N_429,N_1078);
nor U3215 (N_3215,N_530,N_1347);
or U3216 (N_3216,N_2166,N_1361);
nor U3217 (N_3217,N_757,N_1183);
nand U3218 (N_3218,N_1385,N_160);
nand U3219 (N_3219,N_1416,N_450);
nor U3220 (N_3220,N_1043,N_1935);
nor U3221 (N_3221,N_773,N_2212);
nand U3222 (N_3222,N_1550,N_1860);
nand U3223 (N_3223,N_982,N_320);
and U3224 (N_3224,N_97,N_298);
or U3225 (N_3225,N_2149,N_863);
and U3226 (N_3226,N_646,N_2225);
or U3227 (N_3227,N_2258,N_1308);
nor U3228 (N_3228,N_165,N_972);
and U3229 (N_3229,N_508,N_191);
nor U3230 (N_3230,N_1966,N_2409);
nor U3231 (N_3231,N_80,N_834);
or U3232 (N_3232,N_1906,N_1532);
nand U3233 (N_3233,N_2137,N_1442);
nor U3234 (N_3234,N_181,N_408);
and U3235 (N_3235,N_705,N_532);
or U3236 (N_3236,N_1588,N_1073);
and U3237 (N_3237,N_798,N_2046);
xnor U3238 (N_3238,N_338,N_432);
or U3239 (N_3239,N_34,N_2118);
nand U3240 (N_3240,N_2228,N_47);
or U3241 (N_3241,N_366,N_658);
nand U3242 (N_3242,N_2075,N_1098);
nand U3243 (N_3243,N_1807,N_68);
nand U3244 (N_3244,N_1469,N_596);
or U3245 (N_3245,N_1433,N_1340);
and U3246 (N_3246,N_1597,N_588);
and U3247 (N_3247,N_869,N_1699);
nand U3248 (N_3248,N_1994,N_503);
or U3249 (N_3249,N_2461,N_819);
and U3250 (N_3250,N_2018,N_1892);
nor U3251 (N_3251,N_538,N_1641);
and U3252 (N_3252,N_1473,N_1515);
nor U3253 (N_3253,N_799,N_438);
nor U3254 (N_3254,N_1732,N_2414);
and U3255 (N_3255,N_461,N_1368);
nor U3256 (N_3256,N_2401,N_2304);
nand U3257 (N_3257,N_2067,N_384);
nand U3258 (N_3258,N_130,N_1889);
nand U3259 (N_3259,N_2080,N_2068);
and U3260 (N_3260,N_1191,N_525);
nor U3261 (N_3261,N_2029,N_1683);
and U3262 (N_3262,N_791,N_1474);
nor U3263 (N_3263,N_1750,N_1782);
or U3264 (N_3264,N_282,N_1301);
nor U3265 (N_3265,N_1121,N_73);
nand U3266 (N_3266,N_1272,N_836);
xnor U3267 (N_3267,N_1029,N_1809);
or U3268 (N_3268,N_1816,N_1050);
and U3269 (N_3269,N_626,N_2398);
nand U3270 (N_3270,N_991,N_722);
nor U3271 (N_3271,N_2059,N_2286);
nand U3272 (N_3272,N_943,N_1753);
xnor U3273 (N_3273,N_1315,N_676);
nor U3274 (N_3274,N_6,N_2350);
or U3275 (N_3275,N_2273,N_328);
or U3276 (N_3276,N_1700,N_841);
or U3277 (N_3277,N_1327,N_456);
nand U3278 (N_3278,N_915,N_778);
or U3279 (N_3279,N_1793,N_63);
and U3280 (N_3280,N_894,N_604);
and U3281 (N_3281,N_748,N_2211);
or U3282 (N_3282,N_651,N_2081);
xnor U3283 (N_3283,N_1040,N_2329);
and U3284 (N_3284,N_1638,N_618);
nor U3285 (N_3285,N_1403,N_72);
nand U3286 (N_3286,N_2007,N_1910);
and U3287 (N_3287,N_2361,N_1371);
nand U3288 (N_3288,N_1332,N_735);
nand U3289 (N_3289,N_625,N_2343);
or U3290 (N_3290,N_1283,N_1760);
nor U3291 (N_3291,N_2230,N_2128);
nand U3292 (N_3292,N_153,N_1583);
nand U3293 (N_3293,N_1780,N_171);
or U3294 (N_3294,N_442,N_156);
or U3295 (N_3295,N_2396,N_1507);
nor U3296 (N_3296,N_119,N_1563);
or U3297 (N_3297,N_1297,N_2155);
xor U3298 (N_3298,N_1627,N_1592);
nor U3299 (N_3299,N_2101,N_1129);
xor U3300 (N_3300,N_627,N_1829);
and U3301 (N_3301,N_1382,N_1530);
nand U3302 (N_3302,N_2302,N_793);
nand U3303 (N_3303,N_2053,N_535);
nand U3304 (N_3304,N_1263,N_377);
or U3305 (N_3305,N_358,N_1636);
nor U3306 (N_3306,N_2494,N_1723);
and U3307 (N_3307,N_1811,N_99);
xor U3308 (N_3308,N_303,N_1766);
or U3309 (N_3309,N_321,N_496);
or U3310 (N_3310,N_1972,N_416);
nand U3311 (N_3311,N_1244,N_1578);
or U3312 (N_3312,N_79,N_2141);
nor U3313 (N_3313,N_876,N_718);
and U3314 (N_3314,N_1428,N_1024);
nand U3315 (N_3315,N_1038,N_1890);
or U3316 (N_3316,N_1500,N_1980);
or U3317 (N_3317,N_2419,N_2159);
nand U3318 (N_3318,N_1695,N_2051);
nand U3319 (N_3319,N_1939,N_1872);
or U3320 (N_3320,N_1394,N_1876);
nor U3321 (N_3321,N_1016,N_2449);
or U3322 (N_3322,N_2006,N_1163);
xor U3323 (N_3323,N_1175,N_96);
nor U3324 (N_3324,N_1933,N_1590);
and U3325 (N_3325,N_2388,N_1973);
or U3326 (N_3326,N_1740,N_1545);
and U3327 (N_3327,N_36,N_1859);
or U3328 (N_3328,N_1358,N_1465);
and U3329 (N_3329,N_813,N_1596);
and U3330 (N_3330,N_164,N_372);
nor U3331 (N_3331,N_781,N_1847);
or U3332 (N_3332,N_2044,N_1007);
nand U3333 (N_3333,N_2107,N_1867);
or U3334 (N_3334,N_1112,N_388);
or U3335 (N_3335,N_1887,N_1671);
and U3336 (N_3336,N_217,N_2072);
and U3337 (N_3337,N_2481,N_1422);
and U3338 (N_3338,N_137,N_1384);
and U3339 (N_3339,N_2036,N_772);
nor U3340 (N_3340,N_1670,N_279);
nand U3341 (N_3341,N_1663,N_849);
nor U3342 (N_3342,N_1662,N_202);
nor U3343 (N_3343,N_40,N_1238);
and U3344 (N_3344,N_1405,N_598);
and U3345 (N_3345,N_1182,N_248);
nor U3346 (N_3346,N_1095,N_32);
nand U3347 (N_3347,N_1155,N_1153);
nor U3348 (N_3348,N_134,N_1506);
nor U3349 (N_3349,N_1870,N_820);
nor U3350 (N_3350,N_698,N_339);
or U3351 (N_3351,N_1241,N_789);
nand U3352 (N_3352,N_133,N_2175);
and U3353 (N_3353,N_1135,N_1541);
or U3354 (N_3354,N_2237,N_1759);
nand U3355 (N_3355,N_2472,N_1004);
xnor U3356 (N_3356,N_1231,N_163);
nor U3357 (N_3357,N_1981,N_2441);
nand U3358 (N_3358,N_1479,N_301);
or U3359 (N_3359,N_1614,N_1370);
nor U3360 (N_3360,N_125,N_2165);
or U3361 (N_3361,N_963,N_1741);
nand U3362 (N_3362,N_1600,N_233);
or U3363 (N_3363,N_2431,N_2219);
nor U3364 (N_3364,N_942,N_2339);
xnor U3365 (N_3365,N_118,N_141);
and U3366 (N_3366,N_877,N_1767);
nor U3367 (N_3367,N_1813,N_1209);
nand U3368 (N_3368,N_1899,N_105);
and U3369 (N_3369,N_1158,N_1841);
and U3370 (N_3370,N_1607,N_144);
nor U3371 (N_3371,N_1075,N_1320);
and U3372 (N_3372,N_2411,N_2152);
nor U3373 (N_3373,N_2158,N_1941);
and U3374 (N_3374,N_1448,N_1333);
or U3375 (N_3375,N_1124,N_39);
or U3376 (N_3376,N_725,N_1134);
and U3377 (N_3377,N_1996,N_1911);
and U3378 (N_3378,N_199,N_1367);
or U3379 (N_3379,N_1387,N_82);
and U3380 (N_3380,N_1,N_1061);
nand U3381 (N_3381,N_2087,N_1745);
nand U3382 (N_3382,N_1794,N_1798);
or U3383 (N_3383,N_364,N_675);
or U3384 (N_3384,N_1660,N_22);
xnor U3385 (N_3385,N_454,N_2351);
nor U3386 (N_3386,N_323,N_1208);
or U3387 (N_3387,N_261,N_985);
xor U3388 (N_3388,N_1509,N_672);
nor U3389 (N_3389,N_650,N_1714);
nand U3390 (N_3390,N_638,N_401);
nand U3391 (N_3391,N_786,N_1069);
or U3392 (N_3392,N_123,N_1089);
nor U3393 (N_3393,N_796,N_855);
and U3394 (N_3394,N_288,N_1092);
or U3395 (N_3395,N_1336,N_2337);
or U3396 (N_3396,N_1572,N_1425);
or U3397 (N_3397,N_1010,N_2407);
and U3398 (N_3398,N_918,N_1633);
or U3399 (N_3399,N_1410,N_399);
or U3400 (N_3400,N_146,N_1584);
nand U3401 (N_3401,N_2321,N_768);
nand U3402 (N_3402,N_1684,N_2368);
xor U3403 (N_3403,N_289,N_1223);
nor U3404 (N_3404,N_1901,N_8);
or U3405 (N_3405,N_2220,N_132);
xor U3406 (N_3406,N_1248,N_474);
xor U3407 (N_3407,N_1654,N_1944);
or U3408 (N_3408,N_196,N_2099);
nand U3409 (N_3409,N_755,N_322);
nand U3410 (N_3410,N_1875,N_1736);
nand U3411 (N_3411,N_917,N_1249);
nand U3412 (N_3412,N_977,N_254);
or U3413 (N_3413,N_188,N_1937);
or U3414 (N_3414,N_1086,N_2406);
and U3415 (N_3415,N_1928,N_1380);
and U3416 (N_3416,N_1229,N_1488);
or U3417 (N_3417,N_1969,N_2170);
nand U3418 (N_3418,N_1844,N_2424);
xor U3419 (N_3419,N_1529,N_2124);
or U3420 (N_3420,N_340,N_468);
and U3421 (N_3421,N_902,N_1883);
nand U3422 (N_3422,N_1512,N_1808);
nor U3423 (N_3423,N_1252,N_707);
or U3424 (N_3424,N_1951,N_252);
or U3425 (N_3425,N_162,N_557);
nor U3426 (N_3426,N_1389,N_475);
nand U3427 (N_3427,N_635,N_1406);
or U3428 (N_3428,N_337,N_2298);
or U3429 (N_3429,N_526,N_406);
nor U3430 (N_3430,N_1276,N_911);
nand U3431 (N_3431,N_1468,N_42);
nor U3432 (N_3432,N_307,N_1245);
nand U3433 (N_3433,N_1123,N_1393);
xor U3434 (N_3434,N_1873,N_1096);
and U3435 (N_3435,N_23,N_1326);
nand U3436 (N_3436,N_823,N_1115);
and U3437 (N_3437,N_1417,N_370);
or U3438 (N_3438,N_1897,N_2095);
nand U3439 (N_3439,N_1144,N_1266);
and U3440 (N_3440,N_1325,N_2208);
or U3441 (N_3441,N_121,N_1080);
and U3442 (N_3442,N_227,N_2293);
and U3443 (N_3443,N_2336,N_2404);
and U3444 (N_3444,N_2198,N_1299);
nor U3445 (N_3445,N_784,N_1729);
nand U3446 (N_3446,N_2300,N_1771);
or U3447 (N_3447,N_245,N_2460);
nand U3448 (N_3448,N_900,N_2019);
nand U3449 (N_3449,N_510,N_357);
and U3450 (N_3450,N_1622,N_2330);
nor U3451 (N_3451,N_292,N_405);
nor U3452 (N_3452,N_1612,N_1281);
and U3453 (N_3453,N_1216,N_936);
or U3454 (N_3454,N_1418,N_302);
nand U3455 (N_3455,N_1103,N_740);
nand U3456 (N_3456,N_2455,N_336);
or U3457 (N_3457,N_583,N_780);
and U3458 (N_3458,N_92,N_981);
nand U3459 (N_3459,N_728,N_1048);
or U3460 (N_3460,N_2133,N_1817);
nor U3461 (N_3461,N_43,N_745);
nor U3462 (N_3462,N_1983,N_131);
nor U3463 (N_3463,N_2190,N_1997);
nand U3464 (N_3464,N_1390,N_1551);
nor U3465 (N_3465,N_868,N_688);
nand U3466 (N_3466,N_1166,N_1525);
or U3467 (N_3467,N_1151,N_2227);
and U3468 (N_3468,N_2454,N_605);
xor U3469 (N_3469,N_761,N_1383);
or U3470 (N_3470,N_973,N_1990);
nor U3471 (N_3471,N_1517,N_648);
or U3472 (N_3472,N_811,N_2400);
nand U3473 (N_3473,N_2050,N_83);
nand U3474 (N_3474,N_478,N_75);
nand U3475 (N_3475,N_814,N_1152);
nand U3476 (N_3476,N_720,N_1629);
or U3477 (N_3477,N_492,N_205);
nand U3478 (N_3478,N_1795,N_2483);
xnor U3479 (N_3479,N_311,N_2262);
nor U3480 (N_3480,N_185,N_1619);
and U3481 (N_3481,N_2090,N_2387);
nor U3482 (N_3482,N_267,N_2189);
nor U3483 (N_3483,N_480,N_1424);
and U3484 (N_3484,N_1834,N_3);
and U3485 (N_3485,N_1360,N_1055);
nand U3486 (N_3486,N_663,N_1776);
nand U3487 (N_3487,N_330,N_368);
nand U3488 (N_3488,N_2176,N_2193);
xnor U3489 (N_3489,N_2145,N_195);
or U3490 (N_3490,N_1051,N_197);
and U3491 (N_3491,N_1610,N_1499);
nand U3492 (N_3492,N_2235,N_283);
nor U3493 (N_3493,N_112,N_2147);
or U3494 (N_3494,N_2016,N_1006);
or U3495 (N_3495,N_383,N_1930);
and U3496 (N_3496,N_2452,N_2418);
or U3497 (N_3497,N_1651,N_61);
nor U3498 (N_3498,N_1567,N_1200);
and U3499 (N_3499,N_2161,N_2105);
and U3500 (N_3500,N_2381,N_2376);
nor U3501 (N_3501,N_2375,N_176);
or U3502 (N_3502,N_878,N_2384);
and U3503 (N_3503,N_1388,N_996);
or U3504 (N_3504,N_375,N_2184);
nand U3505 (N_3505,N_592,N_1555);
or U3506 (N_3506,N_489,N_264);
nand U3507 (N_3507,N_569,N_1193);
nand U3508 (N_3508,N_505,N_1015);
or U3509 (N_3509,N_2367,N_498);
or U3510 (N_3510,N_1886,N_1100);
nor U3511 (N_3511,N_476,N_1963);
and U3512 (N_3512,N_1593,N_486);
nand U3513 (N_3513,N_1605,N_1553);
nor U3514 (N_3514,N_256,N_750);
or U3515 (N_3515,N_1181,N_1543);
or U3516 (N_3516,N_2372,N_1141);
or U3517 (N_3517,N_2347,N_1628);
nor U3518 (N_3518,N_77,N_933);
or U3519 (N_3519,N_2358,N_473);
nor U3520 (N_3520,N_2338,N_1701);
nand U3521 (N_3521,N_1790,N_593);
nand U3522 (N_3522,N_1799,N_1232);
nor U3523 (N_3523,N_2252,N_240);
and U3524 (N_3524,N_1125,N_2326);
and U3525 (N_3525,N_874,N_831);
nor U3526 (N_3526,N_1259,N_488);
nand U3527 (N_3527,N_1903,N_1991);
nand U3528 (N_3528,N_2093,N_145);
or U3529 (N_3529,N_346,N_696);
nor U3530 (N_3530,N_1441,N_515);
nand U3531 (N_3531,N_1727,N_549);
or U3532 (N_3532,N_1826,N_2482);
and U3533 (N_3533,N_1496,N_212);
xor U3534 (N_3534,N_1420,N_556);
nor U3535 (N_3535,N_2397,N_2311);
and U3536 (N_3536,N_1039,N_2223);
or U3537 (N_3537,N_108,N_1579);
xnor U3538 (N_3538,N_2305,N_858);
and U3539 (N_3539,N_353,N_2428);
nand U3540 (N_3540,N_1349,N_2037);
and U3541 (N_3541,N_193,N_1359);
nand U3542 (N_3542,N_2331,N_850);
nand U3543 (N_3543,N_1632,N_1426);
or U3544 (N_3544,N_947,N_1905);
and U3545 (N_3545,N_547,N_1948);
nor U3546 (N_3546,N_1107,N_1956);
nand U3547 (N_3547,N_2403,N_2089);
nand U3548 (N_3548,N_361,N_300);
nor U3549 (N_3549,N_1988,N_2112);
or U3550 (N_3550,N_2216,N_2318);
and U3551 (N_3551,N_1777,N_1717);
nand U3552 (N_3552,N_1926,N_1288);
nand U3553 (N_3553,N_2233,N_2084);
and U3554 (N_3554,N_477,N_1373);
and U3555 (N_3555,N_1738,N_2086);
or U3556 (N_3556,N_257,N_1587);
nand U3557 (N_3557,N_269,N_2041);
nand U3558 (N_3558,N_1999,N_1188);
and U3559 (N_3559,N_362,N_1331);
nor U3560 (N_3560,N_1330,N_1936);
or U3561 (N_3561,N_1707,N_232);
nand U3562 (N_3562,N_2222,N_1064);
and U3563 (N_3563,N_1343,N_951);
nand U3564 (N_3564,N_1463,N_1668);
nor U3565 (N_3565,N_1708,N_1148);
nand U3566 (N_3566,N_1524,N_686);
and U3567 (N_3567,N_927,N_634);
nor U3568 (N_3568,N_919,N_1866);
or U3569 (N_3569,N_38,N_431);
nand U3570 (N_3570,N_471,N_1720);
and U3571 (N_3571,N_2010,N_389);
and U3572 (N_3572,N_1985,N_1440);
nand U3573 (N_3573,N_1769,N_2115);
nand U3574 (N_3574,N_766,N_419);
xor U3575 (N_3575,N_1071,N_1028);
or U3576 (N_3576,N_1002,N_738);
nand U3577 (N_3577,N_713,N_662);
xor U3578 (N_3578,N_297,N_385);
nand U3579 (N_3579,N_1962,N_1648);
nand U3580 (N_3580,N_2366,N_2487);
or U3581 (N_3581,N_396,N_1502);
nor U3582 (N_3582,N_1854,N_436);
or U3583 (N_3583,N_167,N_1606);
nand U3584 (N_3584,N_509,N_236);
nand U3585 (N_3585,N_2002,N_1476);
nand U3586 (N_3586,N_708,N_2202);
nand U3587 (N_3587,N_1786,N_1845);
or U3588 (N_3588,N_582,N_897);
nor U3589 (N_3589,N_376,N_1234);
and U3590 (N_3590,N_360,N_2083);
or U3591 (N_3591,N_143,N_555);
nor U3592 (N_3592,N_1470,N_1261);
and U3593 (N_3593,N_724,N_2264);
nor U3594 (N_3594,N_744,N_624);
nor U3595 (N_3595,N_1294,N_749);
and U3596 (N_3596,N_2303,N_995);
or U3597 (N_3597,N_412,N_1489);
or U3598 (N_3598,N_1850,N_843);
nand U3599 (N_3599,N_420,N_1621);
nand U3600 (N_3600,N_702,N_1452);
and U3601 (N_3601,N_332,N_2263);
nor U3602 (N_3602,N_1362,N_1934);
nor U3603 (N_3603,N_1310,N_2186);
and U3604 (N_3604,N_1450,N_1569);
or U3605 (N_3605,N_1376,N_1455);
and U3606 (N_3606,N_2391,N_970);
nor U3607 (N_3607,N_584,N_1458);
nor U3608 (N_3608,N_870,N_1783);
nand U3609 (N_3609,N_157,N_1581);
nor U3610 (N_3610,N_1437,N_1685);
nand U3611 (N_3611,N_472,N_1703);
and U3612 (N_3612,N_956,N_2183);
or U3613 (N_3613,N_318,N_2201);
nor U3614 (N_3614,N_2360,N_1711);
or U3615 (N_3615,N_1378,N_1258);
and U3616 (N_3616,N_418,N_1074);
and U3617 (N_3617,N_600,N_867);
or U3618 (N_3618,N_45,N_1072);
and U3619 (N_3619,N_523,N_1282);
and U3620 (N_3620,N_536,N_775);
xnor U3621 (N_3621,N_2179,N_1856);
nand U3622 (N_3622,N_622,N_2475);
nor U3623 (N_3623,N_85,N_33);
or U3624 (N_3624,N_327,N_1312);
nor U3625 (N_3625,N_2207,N_1058);
xnor U3626 (N_3626,N_1090,N_1704);
nand U3627 (N_3627,N_611,N_1504);
nand U3628 (N_3628,N_62,N_1599);
nand U3629 (N_3629,N_931,N_2445);
nor U3630 (N_3630,N_759,N_615);
or U3631 (N_3631,N_1190,N_2265);
nand U3632 (N_3632,N_1122,N_606);
or U3633 (N_3633,N_1522,N_2451);
and U3634 (N_3634,N_1655,N_1291);
xor U3635 (N_3635,N_1483,N_2213);
nor U3636 (N_3636,N_293,N_822);
nand U3637 (N_3637,N_2426,N_2402);
and U3638 (N_3638,N_20,N_862);
nand U3639 (N_3639,N_1447,N_110);
nor U3640 (N_3640,N_159,N_1788);
nor U3641 (N_3641,N_1698,N_1322);
nand U3642 (N_3642,N_805,N_1267);
nand U3643 (N_3643,N_589,N_930);
xnor U3644 (N_3644,N_1047,N_926);
nand U3645 (N_3645,N_87,N_1066);
and U3646 (N_3646,N_1724,N_1091);
nand U3647 (N_3647,N_242,N_1679);
or U3648 (N_3648,N_1056,N_1598);
or U3649 (N_3649,N_1404,N_1350);
nor U3650 (N_3650,N_692,N_213);
and U3651 (N_3651,N_2052,N_397);
or U3652 (N_3652,N_810,N_935);
or U3653 (N_3653,N_2478,N_2495);
or U3654 (N_3654,N_1381,N_2349);
nor U3655 (N_3655,N_797,N_182);
nor U3656 (N_3656,N_1013,N_2042);
and U3657 (N_3657,N_95,N_1949);
and U3658 (N_3658,N_1057,N_1334);
and U3659 (N_3659,N_1626,N_1818);
and U3660 (N_3660,N_91,N_1611);
and U3661 (N_3661,N_1691,N_839);
and U3662 (N_3662,N_642,N_895);
nor U3663 (N_3663,N_2122,N_1637);
nor U3664 (N_3664,N_483,N_848);
and U3665 (N_3665,N_186,N_1031);
nor U3666 (N_3666,N_1984,N_2281);
nor U3667 (N_3667,N_265,N_258);
nor U3668 (N_3668,N_506,N_2394);
and U3669 (N_3669,N_2076,N_1505);
nor U3670 (N_3670,N_262,N_2013);
and U3671 (N_3671,N_2160,N_1664);
nor U3672 (N_3672,N_299,N_986);
nand U3673 (N_3673,N_295,N_2466);
nand U3674 (N_3674,N_971,N_2359);
and U3675 (N_3675,N_1228,N_576);
nor U3676 (N_3676,N_2433,N_857);
and U3677 (N_3677,N_2448,N_2488);
or U3678 (N_3678,N_504,N_2278);
nor U3679 (N_3679,N_1925,N_758);
nor U3680 (N_3680,N_2215,N_601);
nor U3681 (N_3681,N_2082,N_1233);
nand U3682 (N_3682,N_1705,N_594);
nor U3683 (N_3683,N_179,N_1020);
or U3684 (N_3684,N_2294,N_1180);
or U3685 (N_3685,N_1503,N_494);
or U3686 (N_3686,N_1713,N_247);
xnor U3687 (N_3687,N_342,N_2236);
or U3688 (N_3688,N_276,N_712);
nor U3689 (N_3689,N_1429,N_2357);
and U3690 (N_3690,N_678,N_1466);
or U3691 (N_3691,N_487,N_1494);
and U3692 (N_3692,N_1480,N_940);
nand U3693 (N_3693,N_1609,N_1436);
and U3694 (N_3694,N_2181,N_1712);
nand U3695 (N_3695,N_1838,N_2257);
or U3696 (N_3696,N_552,N_616);
and U3697 (N_3697,N_350,N_154);
nor U3698 (N_3698,N_2092,N_835);
nor U3699 (N_3699,N_1896,N_1924);
nor U3700 (N_3700,N_1716,N_140);
nor U3701 (N_3701,N_1917,N_821);
nand U3702 (N_3702,N_2352,N_1033);
nor U3703 (N_3703,N_1920,N_2374);
and U3704 (N_3704,N_2364,N_214);
and U3705 (N_3705,N_314,N_1971);
nor U3706 (N_3706,N_290,N_1275);
nand U3707 (N_3707,N_1815,N_1862);
and U3708 (N_3708,N_1165,N_52);
nor U3709 (N_3709,N_250,N_852);
and U3710 (N_3710,N_832,N_1220);
nor U3711 (N_3711,N_1501,N_1797);
nand U3712 (N_3712,N_2025,N_1105);
or U3713 (N_3713,N_1989,N_590);
or U3714 (N_3714,N_251,N_976);
and U3715 (N_3715,N_1094,N_316);
or U3716 (N_3716,N_421,N_35);
and U3717 (N_3717,N_1544,N_481);
nor U3718 (N_3718,N_1620,N_585);
and U3719 (N_3719,N_1354,N_1490);
and U3720 (N_3720,N_2039,N_2450);
nor U3721 (N_3721,N_1842,N_1353);
or U3722 (N_3722,N_78,N_955);
and U3723 (N_3723,N_979,N_1806);
nand U3724 (N_3724,N_1192,N_2439);
and U3725 (N_3725,N_983,N_2062);
xnor U3726 (N_3726,N_1110,N_24);
and U3727 (N_3727,N_93,N_1475);
nand U3728 (N_3728,N_1207,N_2333);
nor U3729 (N_3729,N_609,N_192);
nand U3730 (N_3730,N_413,N_767);
nand U3731 (N_3731,N_2171,N_561);
or U3732 (N_3732,N_2314,N_2187);
nand U3733 (N_3733,N_847,N_2151);
and U3734 (N_3734,N_48,N_464);
nor U3735 (N_3735,N_1535,N_495);
and U3736 (N_3736,N_59,N_521);
nand U3737 (N_3737,N_1615,N_818);
and U3738 (N_3738,N_2420,N_815);
or U3739 (N_3739,N_2289,N_704);
nor U3740 (N_3740,N_901,N_1011);
and U3741 (N_3741,N_1290,N_218);
nor U3742 (N_3742,N_30,N_1775);
or U3743 (N_3743,N_2415,N_2485);
or U3744 (N_3744,N_1573,N_1401);
xor U3745 (N_3745,N_1273,N_149);
nor U3746 (N_3746,N_424,N_1821);
nor U3747 (N_3747,N_2243,N_348);
or U3748 (N_3748,N_700,N_50);
nand U3749 (N_3749,N_1274,N_907);
or U3750 (N_3750,N_2044,N_1077);
and U3751 (N_3751,N_802,N_1183);
and U3752 (N_3752,N_509,N_197);
nand U3753 (N_3753,N_1854,N_1773);
or U3754 (N_3754,N_1965,N_2283);
or U3755 (N_3755,N_215,N_296);
nand U3756 (N_3756,N_1025,N_1686);
or U3757 (N_3757,N_279,N_57);
or U3758 (N_3758,N_1831,N_1479);
nand U3759 (N_3759,N_1016,N_2245);
or U3760 (N_3760,N_339,N_2326);
nor U3761 (N_3761,N_1693,N_1175);
and U3762 (N_3762,N_118,N_369);
or U3763 (N_3763,N_136,N_535);
nand U3764 (N_3764,N_1656,N_1562);
or U3765 (N_3765,N_2492,N_1238);
and U3766 (N_3766,N_1775,N_1896);
or U3767 (N_3767,N_1244,N_1698);
or U3768 (N_3768,N_1098,N_1621);
nand U3769 (N_3769,N_1416,N_2309);
and U3770 (N_3770,N_971,N_2253);
nor U3771 (N_3771,N_1875,N_2252);
nor U3772 (N_3772,N_1495,N_1374);
and U3773 (N_3773,N_1602,N_2099);
nor U3774 (N_3774,N_1050,N_1714);
nor U3775 (N_3775,N_501,N_1526);
nand U3776 (N_3776,N_166,N_773);
nor U3777 (N_3777,N_1042,N_1195);
and U3778 (N_3778,N_1309,N_858);
and U3779 (N_3779,N_2363,N_26);
nand U3780 (N_3780,N_822,N_377);
or U3781 (N_3781,N_787,N_654);
nor U3782 (N_3782,N_749,N_436);
nor U3783 (N_3783,N_18,N_76);
nor U3784 (N_3784,N_1277,N_1898);
or U3785 (N_3785,N_34,N_481);
nor U3786 (N_3786,N_892,N_2403);
and U3787 (N_3787,N_2226,N_1411);
nand U3788 (N_3788,N_2491,N_810);
or U3789 (N_3789,N_2190,N_1532);
or U3790 (N_3790,N_549,N_2028);
nor U3791 (N_3791,N_806,N_1546);
nor U3792 (N_3792,N_1434,N_1397);
nor U3793 (N_3793,N_158,N_1177);
and U3794 (N_3794,N_1361,N_1008);
nor U3795 (N_3795,N_875,N_2095);
nand U3796 (N_3796,N_1612,N_1541);
or U3797 (N_3797,N_1451,N_864);
or U3798 (N_3798,N_1356,N_477);
or U3799 (N_3799,N_1758,N_836);
nand U3800 (N_3800,N_1579,N_289);
and U3801 (N_3801,N_808,N_2136);
nor U3802 (N_3802,N_321,N_2470);
nand U3803 (N_3803,N_1075,N_2225);
xnor U3804 (N_3804,N_159,N_2034);
and U3805 (N_3805,N_1012,N_1160);
nand U3806 (N_3806,N_1069,N_2372);
and U3807 (N_3807,N_1851,N_244);
nor U3808 (N_3808,N_1946,N_535);
nor U3809 (N_3809,N_1255,N_1269);
and U3810 (N_3810,N_1633,N_491);
or U3811 (N_3811,N_2163,N_291);
nor U3812 (N_3812,N_1654,N_1507);
or U3813 (N_3813,N_1969,N_2053);
or U3814 (N_3814,N_1633,N_2007);
nand U3815 (N_3815,N_1911,N_1146);
nor U3816 (N_3816,N_873,N_1110);
or U3817 (N_3817,N_1878,N_66);
nand U3818 (N_3818,N_959,N_2094);
nor U3819 (N_3819,N_1398,N_1012);
or U3820 (N_3820,N_604,N_1461);
and U3821 (N_3821,N_735,N_1170);
and U3822 (N_3822,N_2133,N_1347);
and U3823 (N_3823,N_811,N_174);
nand U3824 (N_3824,N_2042,N_1669);
or U3825 (N_3825,N_1165,N_2435);
nand U3826 (N_3826,N_2102,N_115);
nor U3827 (N_3827,N_2109,N_2049);
nand U3828 (N_3828,N_957,N_674);
nor U3829 (N_3829,N_1483,N_1386);
nand U3830 (N_3830,N_1902,N_2342);
nor U3831 (N_3831,N_679,N_919);
nor U3832 (N_3832,N_154,N_1362);
nor U3833 (N_3833,N_460,N_887);
and U3834 (N_3834,N_690,N_49);
nor U3835 (N_3835,N_187,N_914);
and U3836 (N_3836,N_1450,N_2301);
or U3837 (N_3837,N_73,N_1100);
or U3838 (N_3838,N_1193,N_1670);
xnor U3839 (N_3839,N_1353,N_820);
xor U3840 (N_3840,N_1250,N_498);
xor U3841 (N_3841,N_528,N_1980);
or U3842 (N_3842,N_2443,N_1125);
or U3843 (N_3843,N_2074,N_731);
nand U3844 (N_3844,N_2380,N_1785);
and U3845 (N_3845,N_987,N_2091);
or U3846 (N_3846,N_2400,N_140);
and U3847 (N_3847,N_2135,N_41);
and U3848 (N_3848,N_1761,N_403);
nor U3849 (N_3849,N_108,N_493);
and U3850 (N_3850,N_2276,N_757);
or U3851 (N_3851,N_2353,N_1533);
nor U3852 (N_3852,N_1817,N_148);
and U3853 (N_3853,N_370,N_2118);
or U3854 (N_3854,N_377,N_981);
nor U3855 (N_3855,N_457,N_1550);
and U3856 (N_3856,N_1445,N_1976);
or U3857 (N_3857,N_1755,N_1970);
and U3858 (N_3858,N_2074,N_340);
xor U3859 (N_3859,N_1712,N_1846);
or U3860 (N_3860,N_817,N_1300);
nand U3861 (N_3861,N_480,N_1594);
or U3862 (N_3862,N_1767,N_1869);
nand U3863 (N_3863,N_1344,N_818);
and U3864 (N_3864,N_2417,N_1892);
or U3865 (N_3865,N_1651,N_248);
or U3866 (N_3866,N_518,N_2206);
nor U3867 (N_3867,N_642,N_2159);
or U3868 (N_3868,N_1858,N_1387);
nand U3869 (N_3869,N_1467,N_1300);
nor U3870 (N_3870,N_1223,N_1447);
nor U3871 (N_3871,N_518,N_418);
or U3872 (N_3872,N_2495,N_1427);
nor U3873 (N_3873,N_2270,N_2165);
or U3874 (N_3874,N_2158,N_608);
and U3875 (N_3875,N_382,N_2230);
nor U3876 (N_3876,N_1939,N_1014);
and U3877 (N_3877,N_2437,N_1496);
nor U3878 (N_3878,N_881,N_1594);
and U3879 (N_3879,N_2294,N_342);
and U3880 (N_3880,N_124,N_1103);
and U3881 (N_3881,N_402,N_1639);
or U3882 (N_3882,N_1068,N_1995);
and U3883 (N_3883,N_2391,N_1597);
and U3884 (N_3884,N_1346,N_351);
xnor U3885 (N_3885,N_1387,N_1543);
or U3886 (N_3886,N_2112,N_510);
or U3887 (N_3887,N_1815,N_1830);
and U3888 (N_3888,N_477,N_882);
and U3889 (N_3889,N_946,N_145);
or U3890 (N_3890,N_1495,N_743);
nor U3891 (N_3891,N_794,N_459);
or U3892 (N_3892,N_861,N_235);
and U3893 (N_3893,N_913,N_1573);
xnor U3894 (N_3894,N_1256,N_2252);
and U3895 (N_3895,N_149,N_35);
nand U3896 (N_3896,N_707,N_1503);
nor U3897 (N_3897,N_2193,N_334);
nor U3898 (N_3898,N_418,N_9);
nor U3899 (N_3899,N_2450,N_174);
or U3900 (N_3900,N_63,N_89);
nand U3901 (N_3901,N_953,N_2402);
nor U3902 (N_3902,N_2175,N_1254);
and U3903 (N_3903,N_430,N_2372);
nor U3904 (N_3904,N_863,N_1964);
or U3905 (N_3905,N_516,N_43);
and U3906 (N_3906,N_534,N_1342);
or U3907 (N_3907,N_64,N_2457);
nor U3908 (N_3908,N_1023,N_743);
or U3909 (N_3909,N_2101,N_2068);
nor U3910 (N_3910,N_339,N_2014);
or U3911 (N_3911,N_1019,N_487);
nor U3912 (N_3912,N_796,N_1300);
and U3913 (N_3913,N_1843,N_2361);
nor U3914 (N_3914,N_1880,N_2288);
or U3915 (N_3915,N_1238,N_1514);
and U3916 (N_3916,N_2046,N_1930);
nor U3917 (N_3917,N_1269,N_2243);
and U3918 (N_3918,N_524,N_761);
nand U3919 (N_3919,N_201,N_43);
and U3920 (N_3920,N_591,N_30);
or U3921 (N_3921,N_1672,N_802);
nand U3922 (N_3922,N_2092,N_1836);
nand U3923 (N_3923,N_2330,N_1996);
nand U3924 (N_3924,N_508,N_357);
nor U3925 (N_3925,N_1520,N_1234);
nand U3926 (N_3926,N_1430,N_1301);
nand U3927 (N_3927,N_1420,N_1439);
or U3928 (N_3928,N_1473,N_780);
nor U3929 (N_3929,N_1290,N_537);
nor U3930 (N_3930,N_622,N_984);
or U3931 (N_3931,N_2340,N_692);
nor U3932 (N_3932,N_1051,N_2246);
nor U3933 (N_3933,N_542,N_2013);
nor U3934 (N_3934,N_52,N_2484);
nand U3935 (N_3935,N_1764,N_1013);
nor U3936 (N_3936,N_35,N_214);
or U3937 (N_3937,N_2137,N_1893);
nor U3938 (N_3938,N_2123,N_397);
nor U3939 (N_3939,N_748,N_1217);
and U3940 (N_3940,N_404,N_873);
and U3941 (N_3941,N_509,N_121);
or U3942 (N_3942,N_834,N_2239);
and U3943 (N_3943,N_1519,N_903);
or U3944 (N_3944,N_275,N_888);
or U3945 (N_3945,N_2434,N_1366);
nor U3946 (N_3946,N_1653,N_1540);
xnor U3947 (N_3947,N_743,N_1703);
nand U3948 (N_3948,N_482,N_525);
nor U3949 (N_3949,N_1445,N_655);
and U3950 (N_3950,N_1015,N_2350);
nand U3951 (N_3951,N_861,N_2345);
nor U3952 (N_3952,N_1547,N_2385);
or U3953 (N_3953,N_1228,N_1093);
nand U3954 (N_3954,N_1200,N_120);
and U3955 (N_3955,N_1668,N_992);
nor U3956 (N_3956,N_480,N_869);
nor U3957 (N_3957,N_246,N_1098);
or U3958 (N_3958,N_711,N_1268);
nor U3959 (N_3959,N_462,N_2390);
or U3960 (N_3960,N_1849,N_884);
or U3961 (N_3961,N_1638,N_2235);
or U3962 (N_3962,N_233,N_1810);
or U3963 (N_3963,N_220,N_2173);
or U3964 (N_3964,N_929,N_2027);
nand U3965 (N_3965,N_2006,N_1069);
or U3966 (N_3966,N_1235,N_325);
nor U3967 (N_3967,N_2047,N_662);
nand U3968 (N_3968,N_2183,N_2410);
nor U3969 (N_3969,N_1901,N_454);
and U3970 (N_3970,N_1868,N_210);
or U3971 (N_3971,N_697,N_2055);
or U3972 (N_3972,N_2191,N_460);
and U3973 (N_3973,N_1532,N_2402);
nand U3974 (N_3974,N_1060,N_2458);
nor U3975 (N_3975,N_1035,N_1176);
and U3976 (N_3976,N_2171,N_1656);
nand U3977 (N_3977,N_765,N_1996);
or U3978 (N_3978,N_951,N_2249);
nor U3979 (N_3979,N_26,N_1748);
nand U3980 (N_3980,N_2321,N_187);
and U3981 (N_3981,N_2389,N_546);
nand U3982 (N_3982,N_115,N_574);
nor U3983 (N_3983,N_1653,N_601);
nand U3984 (N_3984,N_2253,N_2097);
nand U3985 (N_3985,N_777,N_2249);
nor U3986 (N_3986,N_1283,N_1970);
nand U3987 (N_3987,N_1317,N_1642);
and U3988 (N_3988,N_609,N_706);
nand U3989 (N_3989,N_123,N_781);
nand U3990 (N_3990,N_1271,N_8);
or U3991 (N_3991,N_1688,N_1620);
and U3992 (N_3992,N_1394,N_1286);
nor U3993 (N_3993,N_2167,N_595);
nand U3994 (N_3994,N_2345,N_309);
nor U3995 (N_3995,N_274,N_1608);
and U3996 (N_3996,N_513,N_1218);
and U3997 (N_3997,N_1959,N_1361);
or U3998 (N_3998,N_1816,N_1241);
or U3999 (N_3999,N_2026,N_1665);
nand U4000 (N_4000,N_1025,N_1761);
nor U4001 (N_4001,N_1259,N_62);
and U4002 (N_4002,N_1928,N_805);
nand U4003 (N_4003,N_744,N_2372);
and U4004 (N_4004,N_1205,N_2190);
or U4005 (N_4005,N_1798,N_585);
nand U4006 (N_4006,N_1516,N_1839);
nor U4007 (N_4007,N_1169,N_1498);
nor U4008 (N_4008,N_485,N_959);
and U4009 (N_4009,N_1052,N_1563);
nand U4010 (N_4010,N_1807,N_1679);
nand U4011 (N_4011,N_1139,N_2199);
or U4012 (N_4012,N_2273,N_1884);
and U4013 (N_4013,N_1704,N_1437);
nand U4014 (N_4014,N_1590,N_2032);
and U4015 (N_4015,N_2190,N_2033);
nor U4016 (N_4016,N_1132,N_2296);
xnor U4017 (N_4017,N_1687,N_999);
nor U4018 (N_4018,N_1822,N_1313);
nand U4019 (N_4019,N_1585,N_971);
nor U4020 (N_4020,N_510,N_263);
and U4021 (N_4021,N_1097,N_1182);
nor U4022 (N_4022,N_1374,N_103);
or U4023 (N_4023,N_219,N_1971);
and U4024 (N_4024,N_1983,N_1939);
nand U4025 (N_4025,N_520,N_2001);
or U4026 (N_4026,N_832,N_94);
nand U4027 (N_4027,N_457,N_528);
nand U4028 (N_4028,N_2374,N_172);
nand U4029 (N_4029,N_131,N_319);
nor U4030 (N_4030,N_1224,N_148);
and U4031 (N_4031,N_952,N_571);
nand U4032 (N_4032,N_218,N_966);
nand U4033 (N_4033,N_1391,N_127);
nand U4034 (N_4034,N_327,N_1657);
and U4035 (N_4035,N_529,N_32);
nor U4036 (N_4036,N_1205,N_528);
nand U4037 (N_4037,N_1290,N_1293);
and U4038 (N_4038,N_1461,N_2467);
or U4039 (N_4039,N_133,N_435);
nor U4040 (N_4040,N_41,N_1476);
xor U4041 (N_4041,N_1909,N_1401);
nor U4042 (N_4042,N_483,N_1958);
and U4043 (N_4043,N_1590,N_2319);
and U4044 (N_4044,N_269,N_2115);
nor U4045 (N_4045,N_1642,N_1859);
nor U4046 (N_4046,N_187,N_1456);
nor U4047 (N_4047,N_1283,N_345);
and U4048 (N_4048,N_2063,N_2159);
nand U4049 (N_4049,N_1140,N_568);
or U4050 (N_4050,N_579,N_1985);
nor U4051 (N_4051,N_258,N_112);
or U4052 (N_4052,N_456,N_1436);
nand U4053 (N_4053,N_2419,N_1386);
nor U4054 (N_4054,N_494,N_760);
and U4055 (N_4055,N_2494,N_2491);
nand U4056 (N_4056,N_2140,N_1328);
nand U4057 (N_4057,N_853,N_2439);
or U4058 (N_4058,N_279,N_74);
nor U4059 (N_4059,N_2349,N_1455);
or U4060 (N_4060,N_1825,N_141);
or U4061 (N_4061,N_95,N_1702);
xor U4062 (N_4062,N_232,N_191);
nor U4063 (N_4063,N_582,N_1472);
nor U4064 (N_4064,N_1474,N_195);
nor U4065 (N_4065,N_1226,N_1301);
nor U4066 (N_4066,N_2109,N_2191);
nor U4067 (N_4067,N_1262,N_1852);
nand U4068 (N_4068,N_813,N_1690);
and U4069 (N_4069,N_633,N_974);
or U4070 (N_4070,N_27,N_544);
nand U4071 (N_4071,N_665,N_1261);
nand U4072 (N_4072,N_36,N_1412);
or U4073 (N_4073,N_937,N_2488);
or U4074 (N_4074,N_377,N_320);
nand U4075 (N_4075,N_1398,N_2348);
nor U4076 (N_4076,N_1962,N_170);
or U4077 (N_4077,N_890,N_618);
nand U4078 (N_4078,N_1892,N_2393);
nand U4079 (N_4079,N_1972,N_538);
and U4080 (N_4080,N_2163,N_806);
nor U4081 (N_4081,N_2171,N_472);
nand U4082 (N_4082,N_2334,N_1404);
and U4083 (N_4083,N_553,N_2482);
nor U4084 (N_4084,N_1544,N_1487);
nor U4085 (N_4085,N_1287,N_1726);
nand U4086 (N_4086,N_1968,N_2427);
or U4087 (N_4087,N_2471,N_2154);
and U4088 (N_4088,N_687,N_1477);
nor U4089 (N_4089,N_2230,N_252);
nor U4090 (N_4090,N_2273,N_1383);
or U4091 (N_4091,N_1300,N_1427);
nand U4092 (N_4092,N_1381,N_1945);
nor U4093 (N_4093,N_628,N_1287);
and U4094 (N_4094,N_79,N_1118);
or U4095 (N_4095,N_1011,N_218);
nand U4096 (N_4096,N_715,N_780);
and U4097 (N_4097,N_839,N_425);
nor U4098 (N_4098,N_479,N_842);
nand U4099 (N_4099,N_539,N_1616);
or U4100 (N_4100,N_541,N_418);
nand U4101 (N_4101,N_1050,N_425);
or U4102 (N_4102,N_2037,N_540);
nand U4103 (N_4103,N_1655,N_622);
or U4104 (N_4104,N_846,N_1730);
nor U4105 (N_4105,N_309,N_264);
nor U4106 (N_4106,N_650,N_1834);
or U4107 (N_4107,N_1020,N_1323);
or U4108 (N_4108,N_549,N_1145);
nor U4109 (N_4109,N_2491,N_2423);
nand U4110 (N_4110,N_724,N_1844);
and U4111 (N_4111,N_822,N_352);
xnor U4112 (N_4112,N_2224,N_1403);
nor U4113 (N_4113,N_1108,N_2115);
nand U4114 (N_4114,N_152,N_732);
and U4115 (N_4115,N_596,N_1377);
and U4116 (N_4116,N_2177,N_1076);
and U4117 (N_4117,N_2129,N_179);
nand U4118 (N_4118,N_1875,N_1729);
xnor U4119 (N_4119,N_2179,N_895);
or U4120 (N_4120,N_1714,N_2206);
nand U4121 (N_4121,N_1137,N_2068);
nand U4122 (N_4122,N_243,N_2283);
and U4123 (N_4123,N_1617,N_1607);
nor U4124 (N_4124,N_1014,N_2238);
nand U4125 (N_4125,N_1959,N_776);
or U4126 (N_4126,N_1674,N_1015);
or U4127 (N_4127,N_2445,N_1581);
nor U4128 (N_4128,N_1242,N_1601);
nor U4129 (N_4129,N_983,N_1435);
and U4130 (N_4130,N_993,N_1005);
and U4131 (N_4131,N_1702,N_376);
nor U4132 (N_4132,N_2369,N_517);
and U4133 (N_4133,N_1817,N_2061);
and U4134 (N_4134,N_989,N_1564);
and U4135 (N_4135,N_1784,N_2376);
and U4136 (N_4136,N_1434,N_2248);
and U4137 (N_4137,N_1052,N_267);
nand U4138 (N_4138,N_764,N_700);
and U4139 (N_4139,N_537,N_1655);
or U4140 (N_4140,N_1694,N_259);
nor U4141 (N_4141,N_2480,N_717);
nor U4142 (N_4142,N_1260,N_336);
nand U4143 (N_4143,N_2075,N_538);
nand U4144 (N_4144,N_1574,N_2476);
nand U4145 (N_4145,N_910,N_879);
nand U4146 (N_4146,N_1167,N_706);
or U4147 (N_4147,N_1843,N_2386);
nand U4148 (N_4148,N_2442,N_2367);
and U4149 (N_4149,N_436,N_208);
nand U4150 (N_4150,N_1316,N_36);
xnor U4151 (N_4151,N_694,N_927);
nor U4152 (N_4152,N_1150,N_1229);
nor U4153 (N_4153,N_24,N_555);
nor U4154 (N_4154,N_721,N_540);
nand U4155 (N_4155,N_1215,N_893);
and U4156 (N_4156,N_1492,N_730);
nand U4157 (N_4157,N_137,N_616);
nor U4158 (N_4158,N_1121,N_1698);
or U4159 (N_4159,N_834,N_421);
or U4160 (N_4160,N_2208,N_796);
nand U4161 (N_4161,N_1079,N_71);
and U4162 (N_4162,N_1729,N_25);
or U4163 (N_4163,N_281,N_285);
nor U4164 (N_4164,N_592,N_639);
and U4165 (N_4165,N_702,N_397);
nand U4166 (N_4166,N_1861,N_638);
nor U4167 (N_4167,N_632,N_2106);
and U4168 (N_4168,N_2211,N_585);
nand U4169 (N_4169,N_381,N_1717);
nor U4170 (N_4170,N_1336,N_1991);
or U4171 (N_4171,N_1932,N_427);
nand U4172 (N_4172,N_1233,N_1410);
and U4173 (N_4173,N_2142,N_992);
nor U4174 (N_4174,N_2130,N_751);
nand U4175 (N_4175,N_925,N_1334);
and U4176 (N_4176,N_36,N_2083);
and U4177 (N_4177,N_889,N_2358);
and U4178 (N_4178,N_2434,N_1681);
nand U4179 (N_4179,N_631,N_1413);
nor U4180 (N_4180,N_1327,N_1980);
nor U4181 (N_4181,N_1382,N_277);
nor U4182 (N_4182,N_1171,N_1097);
nor U4183 (N_4183,N_159,N_1703);
or U4184 (N_4184,N_2309,N_1576);
nand U4185 (N_4185,N_1254,N_1209);
nand U4186 (N_4186,N_969,N_809);
nor U4187 (N_4187,N_716,N_829);
and U4188 (N_4188,N_403,N_929);
and U4189 (N_4189,N_1716,N_1917);
and U4190 (N_4190,N_2392,N_876);
and U4191 (N_4191,N_935,N_2210);
or U4192 (N_4192,N_545,N_1213);
nand U4193 (N_4193,N_1969,N_181);
nand U4194 (N_4194,N_1326,N_1772);
and U4195 (N_4195,N_1267,N_2201);
nand U4196 (N_4196,N_1000,N_1907);
nor U4197 (N_4197,N_495,N_1333);
or U4198 (N_4198,N_1829,N_2162);
nor U4199 (N_4199,N_134,N_2195);
and U4200 (N_4200,N_547,N_1679);
and U4201 (N_4201,N_502,N_682);
nand U4202 (N_4202,N_1638,N_581);
and U4203 (N_4203,N_1363,N_2305);
or U4204 (N_4204,N_926,N_1370);
nand U4205 (N_4205,N_73,N_2125);
or U4206 (N_4206,N_1032,N_661);
or U4207 (N_4207,N_607,N_729);
or U4208 (N_4208,N_876,N_1523);
nor U4209 (N_4209,N_683,N_564);
nand U4210 (N_4210,N_37,N_491);
nand U4211 (N_4211,N_392,N_1861);
and U4212 (N_4212,N_22,N_2016);
or U4213 (N_4213,N_2449,N_535);
nor U4214 (N_4214,N_179,N_1409);
and U4215 (N_4215,N_2037,N_1997);
or U4216 (N_4216,N_908,N_1499);
and U4217 (N_4217,N_1690,N_1253);
or U4218 (N_4218,N_340,N_749);
nor U4219 (N_4219,N_2471,N_2209);
or U4220 (N_4220,N_92,N_4);
nor U4221 (N_4221,N_2086,N_463);
or U4222 (N_4222,N_642,N_865);
nor U4223 (N_4223,N_428,N_2343);
and U4224 (N_4224,N_71,N_838);
nand U4225 (N_4225,N_148,N_2428);
or U4226 (N_4226,N_0,N_2497);
or U4227 (N_4227,N_1176,N_825);
and U4228 (N_4228,N_1892,N_2310);
nand U4229 (N_4229,N_894,N_2453);
nor U4230 (N_4230,N_1387,N_2393);
and U4231 (N_4231,N_1841,N_1850);
nor U4232 (N_4232,N_343,N_164);
nand U4233 (N_4233,N_1412,N_2268);
nand U4234 (N_4234,N_1363,N_1926);
nand U4235 (N_4235,N_674,N_811);
nor U4236 (N_4236,N_1218,N_158);
or U4237 (N_4237,N_389,N_1778);
and U4238 (N_4238,N_425,N_752);
nor U4239 (N_4239,N_787,N_1651);
nor U4240 (N_4240,N_1118,N_918);
xor U4241 (N_4241,N_1018,N_82);
and U4242 (N_4242,N_2306,N_2275);
nor U4243 (N_4243,N_1678,N_1444);
nor U4244 (N_4244,N_1098,N_438);
or U4245 (N_4245,N_1385,N_861);
nand U4246 (N_4246,N_1745,N_1682);
xor U4247 (N_4247,N_1000,N_431);
or U4248 (N_4248,N_2115,N_1630);
and U4249 (N_4249,N_1990,N_48);
and U4250 (N_4250,N_1787,N_2007);
nand U4251 (N_4251,N_1752,N_1220);
nand U4252 (N_4252,N_1884,N_2122);
nor U4253 (N_4253,N_2447,N_1469);
nand U4254 (N_4254,N_1746,N_1497);
and U4255 (N_4255,N_2437,N_1750);
nand U4256 (N_4256,N_1514,N_2461);
and U4257 (N_4257,N_1655,N_1178);
and U4258 (N_4258,N_2414,N_214);
and U4259 (N_4259,N_409,N_1021);
or U4260 (N_4260,N_436,N_1564);
nand U4261 (N_4261,N_2036,N_1316);
xnor U4262 (N_4262,N_1483,N_2123);
and U4263 (N_4263,N_1948,N_2342);
and U4264 (N_4264,N_2198,N_537);
nor U4265 (N_4265,N_294,N_628);
nand U4266 (N_4266,N_485,N_1562);
nor U4267 (N_4267,N_584,N_1681);
or U4268 (N_4268,N_1650,N_2327);
nand U4269 (N_4269,N_2061,N_281);
nand U4270 (N_4270,N_1898,N_1576);
nand U4271 (N_4271,N_142,N_297);
nand U4272 (N_4272,N_2035,N_1257);
xor U4273 (N_4273,N_1146,N_2313);
or U4274 (N_4274,N_516,N_2099);
or U4275 (N_4275,N_2395,N_1303);
or U4276 (N_4276,N_1791,N_408);
nor U4277 (N_4277,N_242,N_2171);
nor U4278 (N_4278,N_1935,N_2118);
and U4279 (N_4279,N_242,N_1055);
nand U4280 (N_4280,N_2312,N_1412);
and U4281 (N_4281,N_1440,N_1317);
nor U4282 (N_4282,N_2198,N_1450);
or U4283 (N_4283,N_612,N_907);
nor U4284 (N_4284,N_2287,N_1883);
and U4285 (N_4285,N_2156,N_440);
or U4286 (N_4286,N_755,N_304);
nor U4287 (N_4287,N_1102,N_2497);
and U4288 (N_4288,N_203,N_735);
nor U4289 (N_4289,N_1740,N_2130);
nor U4290 (N_4290,N_1541,N_1539);
and U4291 (N_4291,N_998,N_2474);
nor U4292 (N_4292,N_280,N_1310);
nor U4293 (N_4293,N_1837,N_2065);
and U4294 (N_4294,N_65,N_2264);
xor U4295 (N_4295,N_2051,N_1106);
or U4296 (N_4296,N_1379,N_421);
nand U4297 (N_4297,N_1643,N_1173);
and U4298 (N_4298,N_1452,N_2426);
and U4299 (N_4299,N_1009,N_1115);
nand U4300 (N_4300,N_1319,N_1392);
or U4301 (N_4301,N_2316,N_2404);
or U4302 (N_4302,N_1636,N_2386);
or U4303 (N_4303,N_1980,N_1338);
and U4304 (N_4304,N_1201,N_857);
or U4305 (N_4305,N_2012,N_2153);
nor U4306 (N_4306,N_2205,N_1503);
nand U4307 (N_4307,N_104,N_1365);
and U4308 (N_4308,N_1439,N_448);
and U4309 (N_4309,N_957,N_1941);
or U4310 (N_4310,N_1125,N_189);
nand U4311 (N_4311,N_2495,N_1254);
and U4312 (N_4312,N_326,N_729);
or U4313 (N_4313,N_535,N_334);
and U4314 (N_4314,N_2477,N_1289);
and U4315 (N_4315,N_1899,N_1242);
and U4316 (N_4316,N_527,N_173);
or U4317 (N_4317,N_953,N_1430);
nor U4318 (N_4318,N_8,N_518);
nand U4319 (N_4319,N_898,N_2457);
or U4320 (N_4320,N_461,N_298);
and U4321 (N_4321,N_1280,N_1389);
nor U4322 (N_4322,N_1321,N_1524);
and U4323 (N_4323,N_2419,N_536);
or U4324 (N_4324,N_1021,N_2299);
nand U4325 (N_4325,N_2216,N_406);
nand U4326 (N_4326,N_462,N_200);
and U4327 (N_4327,N_400,N_1768);
xor U4328 (N_4328,N_1102,N_2165);
nor U4329 (N_4329,N_672,N_530);
or U4330 (N_4330,N_947,N_1821);
and U4331 (N_4331,N_565,N_179);
nor U4332 (N_4332,N_1372,N_1097);
nand U4333 (N_4333,N_2104,N_1910);
and U4334 (N_4334,N_463,N_1988);
and U4335 (N_4335,N_1736,N_1297);
and U4336 (N_4336,N_1568,N_677);
nor U4337 (N_4337,N_282,N_1097);
nor U4338 (N_4338,N_814,N_1585);
nand U4339 (N_4339,N_1441,N_560);
or U4340 (N_4340,N_1608,N_2478);
nand U4341 (N_4341,N_1200,N_1514);
and U4342 (N_4342,N_1583,N_1192);
nor U4343 (N_4343,N_2365,N_2049);
nor U4344 (N_4344,N_1374,N_34);
xor U4345 (N_4345,N_2101,N_1197);
or U4346 (N_4346,N_2195,N_185);
nor U4347 (N_4347,N_13,N_2293);
xor U4348 (N_4348,N_1109,N_934);
nand U4349 (N_4349,N_2010,N_1693);
nor U4350 (N_4350,N_1812,N_1534);
and U4351 (N_4351,N_1358,N_1137);
or U4352 (N_4352,N_1058,N_798);
nand U4353 (N_4353,N_894,N_1019);
nor U4354 (N_4354,N_2298,N_319);
nand U4355 (N_4355,N_2232,N_362);
and U4356 (N_4356,N_269,N_34);
nor U4357 (N_4357,N_1814,N_794);
nand U4358 (N_4358,N_851,N_284);
and U4359 (N_4359,N_1365,N_1023);
nand U4360 (N_4360,N_981,N_2339);
or U4361 (N_4361,N_47,N_819);
or U4362 (N_4362,N_1160,N_290);
nor U4363 (N_4363,N_1077,N_43);
and U4364 (N_4364,N_1778,N_1992);
xor U4365 (N_4365,N_1609,N_780);
or U4366 (N_4366,N_1047,N_2225);
nand U4367 (N_4367,N_475,N_1063);
or U4368 (N_4368,N_892,N_2162);
nand U4369 (N_4369,N_672,N_1181);
and U4370 (N_4370,N_443,N_2176);
or U4371 (N_4371,N_984,N_663);
nand U4372 (N_4372,N_1951,N_1314);
and U4373 (N_4373,N_2478,N_1134);
and U4374 (N_4374,N_1443,N_1458);
nand U4375 (N_4375,N_1405,N_2059);
and U4376 (N_4376,N_222,N_319);
or U4377 (N_4377,N_385,N_821);
nor U4378 (N_4378,N_704,N_1480);
or U4379 (N_4379,N_440,N_1043);
nor U4380 (N_4380,N_1952,N_879);
nand U4381 (N_4381,N_2169,N_2196);
nand U4382 (N_4382,N_382,N_1493);
nor U4383 (N_4383,N_1312,N_945);
and U4384 (N_4384,N_402,N_2294);
or U4385 (N_4385,N_1478,N_693);
and U4386 (N_4386,N_298,N_2318);
and U4387 (N_4387,N_2037,N_599);
and U4388 (N_4388,N_153,N_1804);
nand U4389 (N_4389,N_1774,N_1095);
nand U4390 (N_4390,N_2457,N_2271);
and U4391 (N_4391,N_394,N_303);
nor U4392 (N_4392,N_728,N_1116);
or U4393 (N_4393,N_1222,N_306);
and U4394 (N_4394,N_312,N_2380);
and U4395 (N_4395,N_891,N_1692);
nand U4396 (N_4396,N_696,N_1559);
nand U4397 (N_4397,N_284,N_198);
and U4398 (N_4398,N_2178,N_2119);
nor U4399 (N_4399,N_2052,N_1084);
nand U4400 (N_4400,N_2212,N_1765);
nand U4401 (N_4401,N_1734,N_702);
and U4402 (N_4402,N_296,N_275);
or U4403 (N_4403,N_1368,N_895);
or U4404 (N_4404,N_588,N_838);
nand U4405 (N_4405,N_572,N_2249);
or U4406 (N_4406,N_1937,N_2203);
nor U4407 (N_4407,N_683,N_535);
and U4408 (N_4408,N_1005,N_585);
or U4409 (N_4409,N_1569,N_805);
or U4410 (N_4410,N_2058,N_391);
nor U4411 (N_4411,N_91,N_1372);
and U4412 (N_4412,N_2391,N_1937);
nand U4413 (N_4413,N_2029,N_1551);
or U4414 (N_4414,N_702,N_2169);
and U4415 (N_4415,N_1203,N_1796);
or U4416 (N_4416,N_1950,N_2169);
and U4417 (N_4417,N_1560,N_343);
and U4418 (N_4418,N_2070,N_1908);
or U4419 (N_4419,N_944,N_2127);
nand U4420 (N_4420,N_439,N_617);
or U4421 (N_4421,N_1328,N_2120);
nand U4422 (N_4422,N_1331,N_55);
or U4423 (N_4423,N_420,N_1663);
and U4424 (N_4424,N_1478,N_2089);
and U4425 (N_4425,N_1110,N_121);
and U4426 (N_4426,N_1476,N_2189);
and U4427 (N_4427,N_1741,N_709);
nand U4428 (N_4428,N_2346,N_567);
nand U4429 (N_4429,N_103,N_1427);
nor U4430 (N_4430,N_2,N_411);
nor U4431 (N_4431,N_2013,N_2280);
and U4432 (N_4432,N_1212,N_2170);
nand U4433 (N_4433,N_555,N_1183);
nor U4434 (N_4434,N_718,N_2374);
nand U4435 (N_4435,N_1595,N_1599);
nand U4436 (N_4436,N_822,N_1847);
or U4437 (N_4437,N_1112,N_309);
xnor U4438 (N_4438,N_2185,N_807);
or U4439 (N_4439,N_2443,N_2362);
and U4440 (N_4440,N_210,N_2240);
and U4441 (N_4441,N_1373,N_1186);
or U4442 (N_4442,N_1583,N_1228);
xor U4443 (N_4443,N_1214,N_1422);
and U4444 (N_4444,N_1621,N_449);
or U4445 (N_4445,N_1331,N_169);
and U4446 (N_4446,N_1950,N_283);
nor U4447 (N_4447,N_1300,N_755);
and U4448 (N_4448,N_1779,N_1361);
nor U4449 (N_4449,N_1057,N_2188);
nand U4450 (N_4450,N_2157,N_440);
nand U4451 (N_4451,N_1357,N_2208);
nor U4452 (N_4452,N_786,N_2139);
and U4453 (N_4453,N_594,N_2449);
nor U4454 (N_4454,N_552,N_685);
and U4455 (N_4455,N_1345,N_2021);
nor U4456 (N_4456,N_2078,N_1982);
and U4457 (N_4457,N_1856,N_1597);
and U4458 (N_4458,N_811,N_995);
nand U4459 (N_4459,N_1301,N_115);
xnor U4460 (N_4460,N_1449,N_389);
nand U4461 (N_4461,N_228,N_2465);
and U4462 (N_4462,N_1086,N_809);
nand U4463 (N_4463,N_1831,N_1367);
nand U4464 (N_4464,N_1817,N_1170);
nor U4465 (N_4465,N_648,N_2447);
or U4466 (N_4466,N_2359,N_714);
nand U4467 (N_4467,N_472,N_2144);
or U4468 (N_4468,N_780,N_1536);
and U4469 (N_4469,N_867,N_1051);
and U4470 (N_4470,N_2093,N_1849);
or U4471 (N_4471,N_1579,N_1843);
nor U4472 (N_4472,N_739,N_2231);
and U4473 (N_4473,N_437,N_2053);
nand U4474 (N_4474,N_1490,N_1146);
nand U4475 (N_4475,N_208,N_1708);
and U4476 (N_4476,N_1499,N_803);
or U4477 (N_4477,N_461,N_2241);
and U4478 (N_4478,N_1840,N_605);
or U4479 (N_4479,N_2037,N_918);
nand U4480 (N_4480,N_1989,N_2381);
nand U4481 (N_4481,N_1534,N_2114);
nor U4482 (N_4482,N_2478,N_2276);
nand U4483 (N_4483,N_1735,N_2138);
and U4484 (N_4484,N_592,N_1872);
or U4485 (N_4485,N_489,N_391);
and U4486 (N_4486,N_784,N_1791);
nand U4487 (N_4487,N_858,N_1006);
nand U4488 (N_4488,N_1845,N_1028);
nor U4489 (N_4489,N_2321,N_1377);
or U4490 (N_4490,N_1248,N_1381);
nor U4491 (N_4491,N_402,N_2065);
nor U4492 (N_4492,N_2265,N_1192);
or U4493 (N_4493,N_583,N_328);
or U4494 (N_4494,N_1590,N_1845);
or U4495 (N_4495,N_226,N_191);
or U4496 (N_4496,N_2211,N_778);
nor U4497 (N_4497,N_1983,N_612);
nor U4498 (N_4498,N_2298,N_1690);
nor U4499 (N_4499,N_1600,N_1249);
and U4500 (N_4500,N_200,N_1814);
nor U4501 (N_4501,N_640,N_221);
nor U4502 (N_4502,N_1416,N_1624);
and U4503 (N_4503,N_459,N_1988);
nor U4504 (N_4504,N_2382,N_1912);
or U4505 (N_4505,N_1529,N_807);
and U4506 (N_4506,N_485,N_1127);
nand U4507 (N_4507,N_2046,N_1648);
nor U4508 (N_4508,N_1694,N_70);
or U4509 (N_4509,N_152,N_2465);
nor U4510 (N_4510,N_382,N_1021);
nand U4511 (N_4511,N_375,N_1762);
or U4512 (N_4512,N_557,N_1062);
and U4513 (N_4513,N_989,N_1335);
xor U4514 (N_4514,N_46,N_827);
nor U4515 (N_4515,N_60,N_426);
nand U4516 (N_4516,N_2082,N_2314);
and U4517 (N_4517,N_2068,N_1379);
and U4518 (N_4518,N_224,N_2408);
and U4519 (N_4519,N_1785,N_728);
or U4520 (N_4520,N_1777,N_323);
or U4521 (N_4521,N_773,N_1096);
nand U4522 (N_4522,N_1589,N_1270);
or U4523 (N_4523,N_1975,N_1354);
nand U4524 (N_4524,N_1151,N_2313);
or U4525 (N_4525,N_535,N_309);
nand U4526 (N_4526,N_1187,N_864);
nand U4527 (N_4527,N_280,N_1669);
and U4528 (N_4528,N_118,N_555);
nand U4529 (N_4529,N_1171,N_1804);
nor U4530 (N_4530,N_1435,N_1164);
nor U4531 (N_4531,N_2430,N_1599);
nand U4532 (N_4532,N_1383,N_1120);
nor U4533 (N_4533,N_947,N_2183);
or U4534 (N_4534,N_1746,N_938);
or U4535 (N_4535,N_1503,N_1176);
nand U4536 (N_4536,N_185,N_1145);
nand U4537 (N_4537,N_250,N_2387);
nand U4538 (N_4538,N_1480,N_444);
nor U4539 (N_4539,N_348,N_321);
nand U4540 (N_4540,N_1428,N_328);
nand U4541 (N_4541,N_1159,N_293);
or U4542 (N_4542,N_1543,N_70);
nand U4543 (N_4543,N_2025,N_1014);
nand U4544 (N_4544,N_2250,N_2207);
and U4545 (N_4545,N_816,N_333);
nand U4546 (N_4546,N_2361,N_1485);
nor U4547 (N_4547,N_351,N_2421);
and U4548 (N_4548,N_115,N_453);
and U4549 (N_4549,N_62,N_1341);
and U4550 (N_4550,N_658,N_1448);
and U4551 (N_4551,N_1819,N_2294);
nand U4552 (N_4552,N_663,N_866);
nand U4553 (N_4553,N_138,N_18);
or U4554 (N_4554,N_1265,N_1233);
and U4555 (N_4555,N_478,N_1124);
nor U4556 (N_4556,N_1776,N_2301);
nand U4557 (N_4557,N_1128,N_382);
nor U4558 (N_4558,N_606,N_1608);
nor U4559 (N_4559,N_1868,N_1491);
or U4560 (N_4560,N_547,N_64);
nor U4561 (N_4561,N_1394,N_825);
or U4562 (N_4562,N_638,N_1157);
or U4563 (N_4563,N_1178,N_1739);
or U4564 (N_4564,N_2131,N_1858);
and U4565 (N_4565,N_1292,N_844);
nand U4566 (N_4566,N_1670,N_2043);
xor U4567 (N_4567,N_1877,N_1115);
and U4568 (N_4568,N_2304,N_14);
or U4569 (N_4569,N_338,N_1181);
nor U4570 (N_4570,N_1847,N_1254);
and U4571 (N_4571,N_2332,N_254);
or U4572 (N_4572,N_877,N_459);
nor U4573 (N_4573,N_2311,N_2084);
nand U4574 (N_4574,N_2251,N_2022);
nor U4575 (N_4575,N_475,N_1244);
and U4576 (N_4576,N_2397,N_964);
or U4577 (N_4577,N_25,N_74);
nand U4578 (N_4578,N_539,N_1956);
or U4579 (N_4579,N_2115,N_2062);
nand U4580 (N_4580,N_1519,N_1844);
nor U4581 (N_4581,N_1223,N_2402);
nand U4582 (N_4582,N_2423,N_288);
nor U4583 (N_4583,N_1361,N_1115);
nor U4584 (N_4584,N_392,N_817);
and U4585 (N_4585,N_1316,N_2064);
nor U4586 (N_4586,N_258,N_617);
nand U4587 (N_4587,N_1133,N_386);
nand U4588 (N_4588,N_1116,N_1519);
and U4589 (N_4589,N_1665,N_50);
or U4590 (N_4590,N_703,N_1252);
nand U4591 (N_4591,N_1941,N_650);
nor U4592 (N_4592,N_909,N_919);
and U4593 (N_4593,N_1603,N_629);
nor U4594 (N_4594,N_1162,N_1897);
nor U4595 (N_4595,N_1812,N_1330);
nand U4596 (N_4596,N_728,N_1400);
nor U4597 (N_4597,N_2382,N_572);
and U4598 (N_4598,N_2164,N_612);
or U4599 (N_4599,N_898,N_73);
nor U4600 (N_4600,N_1799,N_1325);
and U4601 (N_4601,N_1089,N_579);
nor U4602 (N_4602,N_1288,N_1794);
nand U4603 (N_4603,N_1902,N_1809);
and U4604 (N_4604,N_868,N_913);
nor U4605 (N_4605,N_1231,N_389);
and U4606 (N_4606,N_1891,N_2410);
and U4607 (N_4607,N_2116,N_2491);
or U4608 (N_4608,N_887,N_552);
and U4609 (N_4609,N_1941,N_325);
xnor U4610 (N_4610,N_1066,N_1295);
nor U4611 (N_4611,N_943,N_2161);
xor U4612 (N_4612,N_2114,N_309);
and U4613 (N_4613,N_1641,N_1476);
or U4614 (N_4614,N_1483,N_796);
and U4615 (N_4615,N_1809,N_2207);
nand U4616 (N_4616,N_2279,N_1392);
nand U4617 (N_4617,N_456,N_350);
and U4618 (N_4618,N_2089,N_153);
and U4619 (N_4619,N_504,N_100);
or U4620 (N_4620,N_1647,N_758);
and U4621 (N_4621,N_2441,N_1080);
or U4622 (N_4622,N_2453,N_977);
nand U4623 (N_4623,N_2276,N_1357);
nand U4624 (N_4624,N_582,N_1844);
and U4625 (N_4625,N_356,N_644);
and U4626 (N_4626,N_1007,N_1033);
or U4627 (N_4627,N_295,N_634);
xor U4628 (N_4628,N_630,N_271);
or U4629 (N_4629,N_178,N_1613);
nand U4630 (N_4630,N_68,N_640);
and U4631 (N_4631,N_1006,N_635);
and U4632 (N_4632,N_1008,N_1359);
or U4633 (N_4633,N_397,N_989);
nand U4634 (N_4634,N_746,N_1661);
nand U4635 (N_4635,N_1499,N_804);
nand U4636 (N_4636,N_296,N_2372);
nand U4637 (N_4637,N_1586,N_1170);
nor U4638 (N_4638,N_1689,N_1114);
or U4639 (N_4639,N_830,N_973);
nor U4640 (N_4640,N_2267,N_2350);
nand U4641 (N_4641,N_669,N_256);
nand U4642 (N_4642,N_1281,N_1071);
nand U4643 (N_4643,N_1549,N_2206);
nand U4644 (N_4644,N_1999,N_1145);
nand U4645 (N_4645,N_1986,N_2387);
nor U4646 (N_4646,N_550,N_1051);
and U4647 (N_4647,N_709,N_2084);
or U4648 (N_4648,N_437,N_388);
or U4649 (N_4649,N_1969,N_1552);
and U4650 (N_4650,N_213,N_2097);
or U4651 (N_4651,N_1204,N_2453);
or U4652 (N_4652,N_556,N_2331);
or U4653 (N_4653,N_1617,N_822);
nand U4654 (N_4654,N_2153,N_461);
nand U4655 (N_4655,N_1415,N_271);
nand U4656 (N_4656,N_1554,N_295);
nor U4657 (N_4657,N_2466,N_1296);
nand U4658 (N_4658,N_191,N_124);
nor U4659 (N_4659,N_197,N_1860);
nor U4660 (N_4660,N_1366,N_1971);
and U4661 (N_4661,N_8,N_863);
nand U4662 (N_4662,N_215,N_815);
nor U4663 (N_4663,N_1086,N_1033);
nand U4664 (N_4664,N_2399,N_343);
and U4665 (N_4665,N_647,N_1360);
nand U4666 (N_4666,N_1690,N_2333);
and U4667 (N_4667,N_1888,N_1508);
nor U4668 (N_4668,N_2119,N_1365);
or U4669 (N_4669,N_2405,N_1953);
and U4670 (N_4670,N_1009,N_245);
or U4671 (N_4671,N_1220,N_1654);
and U4672 (N_4672,N_1437,N_992);
and U4673 (N_4673,N_1268,N_233);
xnor U4674 (N_4674,N_2197,N_2055);
nand U4675 (N_4675,N_749,N_1722);
and U4676 (N_4676,N_996,N_267);
and U4677 (N_4677,N_1192,N_293);
and U4678 (N_4678,N_75,N_1468);
nor U4679 (N_4679,N_1087,N_1892);
or U4680 (N_4680,N_106,N_1410);
nor U4681 (N_4681,N_2498,N_509);
nand U4682 (N_4682,N_1581,N_689);
or U4683 (N_4683,N_823,N_1400);
and U4684 (N_4684,N_740,N_1715);
nand U4685 (N_4685,N_324,N_2049);
xnor U4686 (N_4686,N_1093,N_246);
and U4687 (N_4687,N_1280,N_1763);
nor U4688 (N_4688,N_2099,N_870);
and U4689 (N_4689,N_1576,N_436);
and U4690 (N_4690,N_1411,N_2307);
or U4691 (N_4691,N_608,N_2293);
and U4692 (N_4692,N_311,N_266);
nor U4693 (N_4693,N_1529,N_928);
nand U4694 (N_4694,N_905,N_1426);
nor U4695 (N_4695,N_1152,N_1602);
nor U4696 (N_4696,N_12,N_1972);
or U4697 (N_4697,N_1447,N_1518);
and U4698 (N_4698,N_21,N_2259);
or U4699 (N_4699,N_1432,N_1728);
and U4700 (N_4700,N_1494,N_746);
or U4701 (N_4701,N_1955,N_716);
or U4702 (N_4702,N_519,N_1519);
nor U4703 (N_4703,N_196,N_781);
nor U4704 (N_4704,N_1709,N_1162);
or U4705 (N_4705,N_44,N_1720);
nand U4706 (N_4706,N_1666,N_1533);
nor U4707 (N_4707,N_2435,N_1108);
and U4708 (N_4708,N_2377,N_1729);
nand U4709 (N_4709,N_791,N_824);
xor U4710 (N_4710,N_1704,N_581);
nor U4711 (N_4711,N_2335,N_1871);
and U4712 (N_4712,N_857,N_896);
and U4713 (N_4713,N_2202,N_2346);
or U4714 (N_4714,N_671,N_2044);
nor U4715 (N_4715,N_530,N_188);
nand U4716 (N_4716,N_304,N_529);
and U4717 (N_4717,N_372,N_2005);
or U4718 (N_4718,N_2423,N_2360);
or U4719 (N_4719,N_1860,N_716);
xnor U4720 (N_4720,N_339,N_1809);
or U4721 (N_4721,N_1743,N_2086);
or U4722 (N_4722,N_2086,N_467);
nor U4723 (N_4723,N_1503,N_2390);
or U4724 (N_4724,N_1001,N_2491);
or U4725 (N_4725,N_331,N_912);
nand U4726 (N_4726,N_1166,N_1196);
nand U4727 (N_4727,N_1612,N_2176);
nand U4728 (N_4728,N_217,N_2060);
and U4729 (N_4729,N_1569,N_1059);
nor U4730 (N_4730,N_40,N_2150);
and U4731 (N_4731,N_712,N_1386);
and U4732 (N_4732,N_594,N_1170);
and U4733 (N_4733,N_2030,N_835);
xor U4734 (N_4734,N_2126,N_1020);
nand U4735 (N_4735,N_2261,N_1059);
xnor U4736 (N_4736,N_2035,N_1945);
nor U4737 (N_4737,N_1252,N_2288);
nor U4738 (N_4738,N_453,N_644);
and U4739 (N_4739,N_642,N_498);
and U4740 (N_4740,N_2406,N_1516);
and U4741 (N_4741,N_1883,N_922);
nor U4742 (N_4742,N_1718,N_2255);
nand U4743 (N_4743,N_2321,N_2004);
and U4744 (N_4744,N_1397,N_1905);
nor U4745 (N_4745,N_716,N_198);
and U4746 (N_4746,N_1597,N_2027);
and U4747 (N_4747,N_818,N_1910);
or U4748 (N_4748,N_2473,N_1911);
and U4749 (N_4749,N_850,N_1386);
nor U4750 (N_4750,N_2489,N_607);
or U4751 (N_4751,N_2359,N_1238);
or U4752 (N_4752,N_2348,N_741);
or U4753 (N_4753,N_205,N_1385);
or U4754 (N_4754,N_181,N_22);
and U4755 (N_4755,N_1306,N_282);
or U4756 (N_4756,N_2407,N_1373);
nand U4757 (N_4757,N_866,N_686);
nand U4758 (N_4758,N_385,N_459);
nand U4759 (N_4759,N_1950,N_2073);
nor U4760 (N_4760,N_1640,N_2004);
or U4761 (N_4761,N_1609,N_2303);
and U4762 (N_4762,N_2159,N_2366);
and U4763 (N_4763,N_386,N_2036);
nand U4764 (N_4764,N_739,N_562);
nand U4765 (N_4765,N_997,N_674);
nand U4766 (N_4766,N_808,N_2305);
and U4767 (N_4767,N_376,N_891);
or U4768 (N_4768,N_745,N_1303);
nand U4769 (N_4769,N_88,N_1565);
nand U4770 (N_4770,N_663,N_607);
or U4771 (N_4771,N_2023,N_993);
and U4772 (N_4772,N_1710,N_600);
or U4773 (N_4773,N_2451,N_416);
or U4774 (N_4774,N_1612,N_2030);
and U4775 (N_4775,N_1938,N_2367);
nand U4776 (N_4776,N_1294,N_2193);
and U4777 (N_4777,N_1,N_677);
nand U4778 (N_4778,N_2263,N_2258);
and U4779 (N_4779,N_1432,N_1921);
nor U4780 (N_4780,N_2016,N_1175);
and U4781 (N_4781,N_376,N_2452);
nor U4782 (N_4782,N_406,N_454);
or U4783 (N_4783,N_2082,N_2125);
or U4784 (N_4784,N_505,N_86);
and U4785 (N_4785,N_395,N_2487);
nand U4786 (N_4786,N_2224,N_1707);
and U4787 (N_4787,N_1801,N_326);
or U4788 (N_4788,N_1469,N_1714);
nand U4789 (N_4789,N_1970,N_2302);
or U4790 (N_4790,N_1299,N_1976);
nand U4791 (N_4791,N_143,N_2488);
and U4792 (N_4792,N_558,N_330);
and U4793 (N_4793,N_1564,N_509);
nor U4794 (N_4794,N_2468,N_1476);
nor U4795 (N_4795,N_2033,N_511);
or U4796 (N_4796,N_1657,N_1070);
and U4797 (N_4797,N_1746,N_678);
and U4798 (N_4798,N_1084,N_1916);
nor U4799 (N_4799,N_1857,N_1788);
nand U4800 (N_4800,N_1132,N_957);
and U4801 (N_4801,N_736,N_2084);
nand U4802 (N_4802,N_2073,N_289);
nor U4803 (N_4803,N_265,N_241);
nor U4804 (N_4804,N_930,N_1533);
xor U4805 (N_4805,N_2215,N_1969);
or U4806 (N_4806,N_256,N_1340);
nand U4807 (N_4807,N_793,N_456);
nor U4808 (N_4808,N_2152,N_597);
nand U4809 (N_4809,N_1961,N_686);
nor U4810 (N_4810,N_888,N_1822);
nor U4811 (N_4811,N_1400,N_700);
or U4812 (N_4812,N_859,N_1930);
and U4813 (N_4813,N_1596,N_684);
nand U4814 (N_4814,N_101,N_1081);
nand U4815 (N_4815,N_833,N_183);
nand U4816 (N_4816,N_745,N_685);
and U4817 (N_4817,N_2435,N_2428);
nand U4818 (N_4818,N_1630,N_81);
nand U4819 (N_4819,N_822,N_2352);
nand U4820 (N_4820,N_1972,N_233);
nor U4821 (N_4821,N_372,N_2325);
nand U4822 (N_4822,N_116,N_2421);
nor U4823 (N_4823,N_1513,N_2042);
or U4824 (N_4824,N_1759,N_1121);
or U4825 (N_4825,N_569,N_2095);
nor U4826 (N_4826,N_1663,N_193);
or U4827 (N_4827,N_1041,N_1359);
or U4828 (N_4828,N_1992,N_1352);
xnor U4829 (N_4829,N_911,N_1783);
or U4830 (N_4830,N_1775,N_2262);
nand U4831 (N_4831,N_1891,N_1421);
and U4832 (N_4832,N_354,N_2443);
nor U4833 (N_4833,N_2348,N_1346);
or U4834 (N_4834,N_2438,N_1123);
or U4835 (N_4835,N_1762,N_1198);
nand U4836 (N_4836,N_1834,N_2068);
or U4837 (N_4837,N_1347,N_2020);
or U4838 (N_4838,N_746,N_1715);
nand U4839 (N_4839,N_1084,N_129);
nand U4840 (N_4840,N_541,N_159);
and U4841 (N_4841,N_1798,N_209);
and U4842 (N_4842,N_820,N_198);
and U4843 (N_4843,N_1418,N_342);
nor U4844 (N_4844,N_2063,N_1599);
and U4845 (N_4845,N_378,N_2461);
or U4846 (N_4846,N_1068,N_655);
nand U4847 (N_4847,N_1329,N_378);
and U4848 (N_4848,N_1946,N_426);
nor U4849 (N_4849,N_1770,N_166);
nor U4850 (N_4850,N_2299,N_2161);
and U4851 (N_4851,N_2003,N_828);
or U4852 (N_4852,N_685,N_2217);
nor U4853 (N_4853,N_121,N_490);
and U4854 (N_4854,N_2344,N_1559);
or U4855 (N_4855,N_1517,N_1425);
and U4856 (N_4856,N_1644,N_119);
nor U4857 (N_4857,N_1416,N_2445);
and U4858 (N_4858,N_891,N_900);
or U4859 (N_4859,N_2225,N_895);
and U4860 (N_4860,N_785,N_1086);
nor U4861 (N_4861,N_1832,N_641);
and U4862 (N_4862,N_1954,N_770);
nand U4863 (N_4863,N_720,N_1576);
or U4864 (N_4864,N_224,N_451);
nor U4865 (N_4865,N_106,N_441);
nand U4866 (N_4866,N_1979,N_699);
nor U4867 (N_4867,N_551,N_306);
nand U4868 (N_4868,N_599,N_1788);
or U4869 (N_4869,N_1700,N_1925);
or U4870 (N_4870,N_315,N_1635);
or U4871 (N_4871,N_2018,N_1494);
nor U4872 (N_4872,N_10,N_2110);
nand U4873 (N_4873,N_725,N_2135);
nor U4874 (N_4874,N_50,N_565);
nand U4875 (N_4875,N_2285,N_1565);
nand U4876 (N_4876,N_1301,N_2094);
nand U4877 (N_4877,N_13,N_159);
nand U4878 (N_4878,N_1355,N_671);
or U4879 (N_4879,N_1152,N_1298);
and U4880 (N_4880,N_938,N_410);
nand U4881 (N_4881,N_267,N_1632);
and U4882 (N_4882,N_2368,N_1121);
nand U4883 (N_4883,N_102,N_284);
or U4884 (N_4884,N_1857,N_1826);
or U4885 (N_4885,N_942,N_364);
nand U4886 (N_4886,N_1795,N_847);
or U4887 (N_4887,N_1318,N_1369);
or U4888 (N_4888,N_2313,N_1315);
nand U4889 (N_4889,N_1358,N_16);
or U4890 (N_4890,N_2188,N_265);
and U4891 (N_4891,N_570,N_1271);
and U4892 (N_4892,N_1005,N_869);
nand U4893 (N_4893,N_2080,N_2079);
nand U4894 (N_4894,N_2348,N_1995);
nor U4895 (N_4895,N_1905,N_1434);
or U4896 (N_4896,N_239,N_1355);
and U4897 (N_4897,N_1871,N_2264);
nor U4898 (N_4898,N_1632,N_925);
and U4899 (N_4899,N_741,N_1931);
nand U4900 (N_4900,N_705,N_732);
or U4901 (N_4901,N_1802,N_1491);
and U4902 (N_4902,N_908,N_1897);
or U4903 (N_4903,N_1991,N_1601);
or U4904 (N_4904,N_2343,N_2069);
xor U4905 (N_4905,N_2071,N_1372);
nand U4906 (N_4906,N_1800,N_1431);
nor U4907 (N_4907,N_777,N_143);
and U4908 (N_4908,N_2380,N_1257);
nor U4909 (N_4909,N_2475,N_1051);
xor U4910 (N_4910,N_2288,N_1440);
and U4911 (N_4911,N_2380,N_774);
or U4912 (N_4912,N_651,N_1462);
and U4913 (N_4913,N_2175,N_1291);
and U4914 (N_4914,N_1068,N_982);
nand U4915 (N_4915,N_159,N_88);
and U4916 (N_4916,N_726,N_679);
nand U4917 (N_4917,N_980,N_1562);
xnor U4918 (N_4918,N_124,N_1555);
or U4919 (N_4919,N_952,N_2220);
and U4920 (N_4920,N_1838,N_2248);
or U4921 (N_4921,N_2448,N_2123);
or U4922 (N_4922,N_2270,N_269);
and U4923 (N_4923,N_800,N_1235);
or U4924 (N_4924,N_553,N_1085);
or U4925 (N_4925,N_860,N_1317);
nand U4926 (N_4926,N_1316,N_1100);
nor U4927 (N_4927,N_1986,N_1398);
and U4928 (N_4928,N_1095,N_704);
nor U4929 (N_4929,N_2011,N_717);
or U4930 (N_4930,N_2097,N_1540);
nor U4931 (N_4931,N_1840,N_302);
nand U4932 (N_4932,N_2376,N_1237);
or U4933 (N_4933,N_2462,N_1915);
xor U4934 (N_4934,N_1188,N_2222);
and U4935 (N_4935,N_88,N_107);
nand U4936 (N_4936,N_263,N_1858);
or U4937 (N_4937,N_1507,N_935);
and U4938 (N_4938,N_18,N_1483);
xnor U4939 (N_4939,N_425,N_1501);
and U4940 (N_4940,N_904,N_760);
and U4941 (N_4941,N_2325,N_1151);
and U4942 (N_4942,N_1818,N_1286);
or U4943 (N_4943,N_2303,N_18);
nand U4944 (N_4944,N_1641,N_1942);
nand U4945 (N_4945,N_1185,N_351);
and U4946 (N_4946,N_193,N_1689);
or U4947 (N_4947,N_301,N_2345);
nor U4948 (N_4948,N_1826,N_819);
nor U4949 (N_4949,N_1972,N_160);
or U4950 (N_4950,N_748,N_1720);
and U4951 (N_4951,N_767,N_1970);
nand U4952 (N_4952,N_1331,N_1237);
nor U4953 (N_4953,N_1119,N_1832);
nor U4954 (N_4954,N_2069,N_2173);
and U4955 (N_4955,N_2294,N_908);
or U4956 (N_4956,N_366,N_1732);
or U4957 (N_4957,N_1165,N_1298);
nand U4958 (N_4958,N_2431,N_1550);
nor U4959 (N_4959,N_1442,N_1245);
nand U4960 (N_4960,N_2085,N_1615);
and U4961 (N_4961,N_185,N_163);
nor U4962 (N_4962,N_1453,N_333);
xor U4963 (N_4963,N_1569,N_2074);
nor U4964 (N_4964,N_2389,N_1958);
nor U4965 (N_4965,N_768,N_1271);
and U4966 (N_4966,N_1191,N_594);
nand U4967 (N_4967,N_658,N_363);
nand U4968 (N_4968,N_768,N_166);
or U4969 (N_4969,N_793,N_2324);
and U4970 (N_4970,N_1900,N_18);
nor U4971 (N_4971,N_1829,N_2443);
or U4972 (N_4972,N_1856,N_2285);
nor U4973 (N_4973,N_107,N_847);
nand U4974 (N_4974,N_2028,N_1993);
and U4975 (N_4975,N_1140,N_2219);
nand U4976 (N_4976,N_1717,N_1314);
and U4977 (N_4977,N_1066,N_647);
or U4978 (N_4978,N_511,N_420);
or U4979 (N_4979,N_2249,N_1580);
or U4980 (N_4980,N_1943,N_328);
and U4981 (N_4981,N_1940,N_1150);
nor U4982 (N_4982,N_1234,N_394);
nor U4983 (N_4983,N_2189,N_909);
or U4984 (N_4984,N_750,N_1685);
or U4985 (N_4985,N_1787,N_131);
nand U4986 (N_4986,N_1926,N_441);
and U4987 (N_4987,N_926,N_2468);
or U4988 (N_4988,N_283,N_1479);
nor U4989 (N_4989,N_1616,N_1570);
or U4990 (N_4990,N_934,N_2330);
nand U4991 (N_4991,N_1277,N_284);
nand U4992 (N_4992,N_1748,N_1792);
or U4993 (N_4993,N_1692,N_1952);
or U4994 (N_4994,N_2149,N_2357);
or U4995 (N_4995,N_2300,N_1389);
or U4996 (N_4996,N_2295,N_683);
or U4997 (N_4997,N_1199,N_2464);
nand U4998 (N_4998,N_209,N_1337);
or U4999 (N_4999,N_1285,N_1880);
or UO_0 (O_0,N_3109,N_4349);
nor UO_1 (O_1,N_3757,N_3857);
nor UO_2 (O_2,N_2533,N_2953);
nand UO_3 (O_3,N_3934,N_3259);
or UO_4 (O_4,N_4118,N_4901);
or UO_5 (O_5,N_3189,N_3446);
nor UO_6 (O_6,N_4254,N_4031);
nand UO_7 (O_7,N_3768,N_3111);
and UO_8 (O_8,N_3560,N_3214);
or UO_9 (O_9,N_4823,N_2674);
and UO_10 (O_10,N_4749,N_3213);
nor UO_11 (O_11,N_2597,N_4251);
nand UO_12 (O_12,N_2992,N_2902);
nor UO_13 (O_13,N_3094,N_4745);
and UO_14 (O_14,N_2876,N_3639);
nand UO_15 (O_15,N_4314,N_4259);
or UO_16 (O_16,N_3564,N_3584);
nand UO_17 (O_17,N_2565,N_3566);
or UO_18 (O_18,N_2628,N_4389);
and UO_19 (O_19,N_4830,N_4121);
and UO_20 (O_20,N_4353,N_3902);
xor UO_21 (O_21,N_3979,N_2934);
and UO_22 (O_22,N_3037,N_4980);
or UO_23 (O_23,N_3572,N_4120);
nor UO_24 (O_24,N_4681,N_4036);
nor UO_25 (O_25,N_3855,N_4456);
nand UO_26 (O_26,N_2683,N_3506);
nor UO_27 (O_27,N_4498,N_3157);
nand UO_28 (O_28,N_4674,N_4781);
nor UO_29 (O_29,N_3669,N_2870);
nand UO_30 (O_30,N_3676,N_3479);
and UO_31 (O_31,N_2569,N_3098);
nor UO_32 (O_32,N_3498,N_2756);
nor UO_33 (O_33,N_4257,N_3346);
xnor UO_34 (O_34,N_3627,N_4009);
and UO_35 (O_35,N_3968,N_4045);
and UO_36 (O_36,N_4042,N_3910);
nand UO_37 (O_37,N_3158,N_4923);
nand UO_38 (O_38,N_3725,N_4175);
nand UO_39 (O_39,N_2842,N_4744);
nor UO_40 (O_40,N_4538,N_3394);
nor UO_41 (O_41,N_4184,N_4469);
xnor UO_42 (O_42,N_3672,N_2768);
nand UO_43 (O_43,N_3337,N_4873);
or UO_44 (O_44,N_3699,N_4424);
or UO_45 (O_45,N_3279,N_3803);
nand UO_46 (O_46,N_3173,N_4037);
and UO_47 (O_47,N_2918,N_2723);
and UO_48 (O_48,N_4912,N_3435);
or UO_49 (O_49,N_2670,N_3271);
and UO_50 (O_50,N_4714,N_2727);
nand UO_51 (O_51,N_4577,N_3860);
nand UO_52 (O_52,N_3222,N_2690);
and UO_53 (O_53,N_2894,N_3997);
nor UO_54 (O_54,N_3804,N_2779);
or UO_55 (O_55,N_3796,N_3220);
nand UO_56 (O_56,N_4137,N_3389);
nor UO_57 (O_57,N_4866,N_4084);
or UO_58 (O_58,N_4574,N_4740);
and UO_59 (O_59,N_3495,N_3439);
or UO_60 (O_60,N_4810,N_2998);
nand UO_61 (O_61,N_4330,N_3011);
nor UO_62 (O_62,N_3526,N_4591);
and UO_63 (O_63,N_3053,N_4324);
xnor UO_64 (O_64,N_4971,N_4530);
nand UO_65 (O_65,N_3928,N_3123);
nand UO_66 (O_66,N_3976,N_4156);
nand UO_67 (O_67,N_4652,N_4378);
or UO_68 (O_68,N_4943,N_4559);
and UO_69 (O_69,N_2782,N_2607);
nor UO_70 (O_70,N_3964,N_2958);
and UO_71 (O_71,N_3028,N_3946);
xor UO_72 (O_72,N_3649,N_3800);
nand UO_73 (O_73,N_3689,N_4896);
or UO_74 (O_74,N_3587,N_4826);
nand UO_75 (O_75,N_4524,N_4972);
xnor UO_76 (O_76,N_4179,N_3944);
nor UO_77 (O_77,N_3453,N_4769);
or UO_78 (O_78,N_3146,N_2623);
nor UO_79 (O_79,N_4565,N_4139);
and UO_80 (O_80,N_4091,N_4768);
nor UO_81 (O_81,N_4479,N_4484);
or UO_82 (O_82,N_2844,N_4447);
nand UO_83 (O_83,N_3936,N_3315);
nor UO_84 (O_84,N_2616,N_4004);
or UO_85 (O_85,N_2691,N_3151);
or UO_86 (O_86,N_2729,N_4428);
or UO_87 (O_87,N_4627,N_3846);
nand UO_88 (O_88,N_4271,N_4522);
or UO_89 (O_89,N_2738,N_3207);
nand UO_90 (O_90,N_3361,N_2721);
or UO_91 (O_91,N_4289,N_3142);
nor UO_92 (O_92,N_3283,N_2743);
nand UO_93 (O_93,N_3478,N_2999);
xor UO_94 (O_94,N_3562,N_3040);
nand UO_95 (O_95,N_4857,N_3540);
xor UO_96 (O_96,N_4395,N_4169);
nand UO_97 (O_97,N_2851,N_4193);
nor UO_98 (O_98,N_2830,N_3813);
nand UO_99 (O_99,N_2575,N_4101);
nor UO_100 (O_100,N_3835,N_4216);
or UO_101 (O_101,N_4489,N_3191);
and UO_102 (O_102,N_4820,N_3019);
or UO_103 (O_103,N_3538,N_4317);
nand UO_104 (O_104,N_3014,N_3168);
and UO_105 (O_105,N_3422,N_4816);
nor UO_106 (O_106,N_2875,N_2862);
nor UO_107 (O_107,N_3126,N_2715);
or UO_108 (O_108,N_2922,N_2502);
nand UO_109 (O_109,N_3443,N_4959);
or UO_110 (O_110,N_3785,N_2733);
and UO_111 (O_111,N_3172,N_3635);
or UO_112 (O_112,N_2706,N_2961);
nor UO_113 (O_113,N_3752,N_4159);
nor UO_114 (O_114,N_3074,N_2677);
nand UO_115 (O_115,N_4679,N_2649);
xnor UO_116 (O_116,N_4644,N_4108);
and UO_117 (O_117,N_3680,N_4828);
xor UO_118 (O_118,N_4352,N_2503);
xnor UO_119 (O_119,N_4523,N_4710);
nor UO_120 (O_120,N_3782,N_3243);
nand UO_121 (O_121,N_2976,N_4548);
nand UO_122 (O_122,N_4372,N_4936);
and UO_123 (O_123,N_3115,N_3603);
nor UO_124 (O_124,N_2696,N_4629);
or UO_125 (O_125,N_3728,N_2750);
and UO_126 (O_126,N_4918,N_3240);
and UO_127 (O_127,N_4895,N_2765);
nor UO_128 (O_128,N_3006,N_2567);
nor UO_129 (O_129,N_3816,N_3036);
nor UO_130 (O_130,N_3704,N_3862);
xor UO_131 (O_131,N_4481,N_2773);
and UO_132 (O_132,N_3314,N_2647);
and UO_133 (O_133,N_3853,N_4623);
nor UO_134 (O_134,N_3140,N_2511);
nand UO_135 (O_135,N_2589,N_3553);
or UO_136 (O_136,N_3227,N_3416);
or UO_137 (O_137,N_4829,N_2559);
or UO_138 (O_138,N_3937,N_4541);
and UO_139 (O_139,N_2653,N_2991);
nand UO_140 (O_140,N_3960,N_4669);
nor UO_141 (O_141,N_4991,N_2536);
or UO_142 (O_142,N_4265,N_2679);
nand UO_143 (O_143,N_2563,N_4285);
nor UO_144 (O_144,N_3356,N_3079);
nor UO_145 (O_145,N_4490,N_4474);
and UO_146 (O_146,N_3223,N_4398);
and UO_147 (O_147,N_4527,N_2813);
or UO_148 (O_148,N_4071,N_4181);
nor UO_149 (O_149,N_2913,N_4465);
nor UO_150 (O_150,N_4850,N_4907);
nor UO_151 (O_151,N_2893,N_3848);
and UO_152 (O_152,N_3382,N_3867);
nand UO_153 (O_153,N_4228,N_2771);
and UO_154 (O_154,N_2975,N_4536);
and UO_155 (O_155,N_4645,N_2891);
nand UO_156 (O_156,N_3253,N_4663);
nand UO_157 (O_157,N_3286,N_4468);
or UO_158 (O_158,N_4666,N_3234);
or UO_159 (O_159,N_4255,N_3907);
or UO_160 (O_160,N_2985,N_2711);
nand UO_161 (O_161,N_3693,N_4570);
nor UO_162 (O_162,N_3543,N_3952);
nor UO_163 (O_163,N_3720,N_3657);
or UO_164 (O_164,N_2686,N_2621);
nand UO_165 (O_165,N_4968,N_2957);
nand UO_166 (O_166,N_2896,N_4958);
nand UO_167 (O_167,N_3194,N_4551);
and UO_168 (O_168,N_4420,N_4805);
or UO_169 (O_169,N_4290,N_4041);
or UO_170 (O_170,N_4619,N_2929);
and UO_171 (O_171,N_2701,N_3056);
nor UO_172 (O_172,N_3459,N_3050);
and UO_173 (O_173,N_4162,N_3503);
nor UO_174 (O_174,N_2665,N_4725);
nand UO_175 (O_175,N_2507,N_2518);
nor UO_176 (O_176,N_2553,N_3476);
or UO_177 (O_177,N_2549,N_2906);
or UO_178 (O_178,N_4965,N_4925);
and UO_179 (O_179,N_3177,N_3778);
nor UO_180 (O_180,N_3268,N_4329);
and UO_181 (O_181,N_3201,N_3089);
and UO_182 (O_182,N_2822,N_2501);
nor UO_183 (O_183,N_3822,N_3811);
or UO_184 (O_184,N_4584,N_4607);
and UO_185 (O_185,N_3027,N_3504);
and UO_186 (O_186,N_4438,N_2529);
or UO_187 (O_187,N_3444,N_3861);
nor UO_188 (O_188,N_4864,N_4643);
nor UO_189 (O_189,N_4192,N_3766);
and UO_190 (O_190,N_4273,N_4032);
nor UO_191 (O_191,N_3690,N_4412);
xnor UO_192 (O_192,N_3100,N_2745);
nor UO_193 (O_193,N_4753,N_4222);
nand UO_194 (O_194,N_4564,N_2583);
nor UO_195 (O_195,N_3351,N_4476);
and UO_196 (O_196,N_2714,N_2637);
or UO_197 (O_197,N_4408,N_2718);
nor UO_198 (O_198,N_3180,N_4556);
nand UO_199 (O_199,N_4982,N_4385);
nand UO_200 (O_200,N_4677,N_4478);
nor UO_201 (O_201,N_4340,N_4717);
and UO_202 (O_202,N_4836,N_3262);
or UO_203 (O_203,N_3310,N_2836);
and UO_204 (O_204,N_2989,N_4964);
nor UO_205 (O_205,N_2886,N_3580);
nand UO_206 (O_206,N_3674,N_2702);
nor UO_207 (O_207,N_2633,N_2785);
nor UO_208 (O_208,N_4702,N_2919);
xor UO_209 (O_209,N_2852,N_4076);
nand UO_210 (O_210,N_3149,N_3386);
or UO_211 (O_211,N_3159,N_3773);
nor UO_212 (O_212,N_3001,N_3246);
nand UO_213 (O_213,N_3534,N_2708);
and UO_214 (O_214,N_3380,N_4954);
and UO_215 (O_215,N_3043,N_3398);
or UO_216 (O_216,N_4440,N_2869);
or UO_217 (O_217,N_3633,N_4201);
and UO_218 (O_218,N_3107,N_4086);
nor UO_219 (O_219,N_2551,N_2660);
or UO_220 (O_220,N_3837,N_4834);
or UO_221 (O_221,N_4328,N_4676);
nand UO_222 (O_222,N_3719,N_3113);
or UO_223 (O_223,N_4535,N_2821);
or UO_224 (O_224,N_4592,N_4446);
xor UO_225 (O_225,N_3959,N_3880);
nand UO_226 (O_226,N_4167,N_2560);
nand UO_227 (O_227,N_3329,N_3845);
or UO_228 (O_228,N_4871,N_3638);
nor UO_229 (O_229,N_3806,N_3667);
nand UO_230 (O_230,N_4783,N_3842);
and UO_231 (O_231,N_3808,N_3278);
or UO_232 (O_232,N_2952,N_2645);
nor UO_233 (O_233,N_4305,N_3130);
nor UO_234 (O_234,N_4609,N_3359);
nor UO_235 (O_235,N_3762,N_3396);
or UO_236 (O_236,N_3723,N_3588);
nand UO_237 (O_237,N_4521,N_4161);
nor UO_238 (O_238,N_2736,N_4675);
or UO_239 (O_239,N_3654,N_4747);
nand UO_240 (O_240,N_3895,N_4888);
nand UO_241 (O_241,N_3033,N_3288);
and UO_242 (O_242,N_4132,N_3701);
nand UO_243 (O_243,N_3894,N_4715);
and UO_244 (O_244,N_4779,N_4143);
nand UO_245 (O_245,N_3962,N_2635);
or UO_246 (O_246,N_4734,N_4597);
and UO_247 (O_247,N_3841,N_3708);
and UO_248 (O_248,N_2766,N_4087);
nor UO_249 (O_249,N_2923,N_2856);
or UO_250 (O_250,N_3652,N_4471);
nand UO_251 (O_251,N_3576,N_2781);
and UO_252 (O_252,N_4406,N_2513);
and UO_253 (O_253,N_4660,N_2889);
or UO_254 (O_254,N_4989,N_3664);
nand UO_255 (O_255,N_2930,N_4622);
or UO_256 (O_256,N_4376,N_3397);
or UO_257 (O_257,N_4572,N_4914);
nand UO_258 (O_258,N_2545,N_2587);
or UO_259 (O_259,N_4417,N_4653);
nor UO_260 (O_260,N_4000,N_4932);
and UO_261 (O_261,N_4347,N_3629);
and UO_262 (O_262,N_3912,N_3623);
nand UO_263 (O_263,N_4951,N_4600);
nand UO_264 (O_264,N_4413,N_3174);
nand UO_265 (O_265,N_4432,N_4399);
nor UO_266 (O_266,N_3181,N_4311);
or UO_267 (O_267,N_2546,N_4593);
or UO_268 (O_268,N_4765,N_3204);
or UO_269 (O_269,N_4001,N_4778);
nor UO_270 (O_270,N_3646,N_3301);
nor UO_271 (O_271,N_2601,N_3438);
or UO_272 (O_272,N_4845,N_4291);
nand UO_273 (O_273,N_2979,N_4852);
nor UO_274 (O_274,N_4099,N_2969);
nor UO_275 (O_275,N_4135,N_3509);
nand UO_276 (O_276,N_3292,N_4631);
and UO_277 (O_277,N_3660,N_4690);
or UO_278 (O_278,N_3625,N_4069);
nor UO_279 (O_279,N_4908,N_2861);
nand UO_280 (O_280,N_3618,N_4831);
nor UO_281 (O_281,N_3415,N_2837);
nand UO_282 (O_282,N_3449,N_4142);
xor UO_283 (O_283,N_4557,N_4081);
or UO_284 (O_284,N_3252,N_3843);
or UO_285 (O_285,N_4583,N_2620);
and UO_286 (O_286,N_4343,N_4217);
nand UO_287 (O_287,N_4332,N_2845);
or UO_288 (O_288,N_2624,N_4787);
nor UO_289 (O_289,N_2828,N_3230);
nand UO_290 (O_290,N_3349,N_3484);
nor UO_291 (O_291,N_3103,N_3413);
or UO_292 (O_292,N_4308,N_4310);
or UO_293 (O_293,N_3235,N_3557);
nor UO_294 (O_294,N_2899,N_2539);
nand UO_295 (O_295,N_4602,N_4392);
nor UO_296 (O_296,N_4299,N_3745);
nand UO_297 (O_297,N_3399,N_4851);
or UO_298 (O_298,N_4242,N_4334);
or UO_299 (O_299,N_3695,N_2885);
and UO_300 (O_300,N_2693,N_3076);
and UO_301 (O_301,N_3465,N_3241);
nor UO_302 (O_302,N_3705,N_3090);
or UO_303 (O_303,N_3497,N_4414);
nor UO_304 (O_304,N_4729,N_3748);
nor UO_305 (O_305,N_3573,N_4790);
or UO_306 (O_306,N_3939,N_2746);
or UO_307 (O_307,N_3330,N_4067);
or UO_308 (O_308,N_2866,N_4421);
nor UO_309 (O_309,N_3148,N_2854);
or UO_310 (O_310,N_3215,N_4759);
nand UO_311 (O_311,N_4373,N_3978);
or UO_312 (O_312,N_4919,N_2948);
and UO_313 (O_313,N_4097,N_4292);
nand UO_314 (O_314,N_2940,N_3170);
nor UO_315 (O_315,N_4470,N_4282);
nor UO_316 (O_316,N_4301,N_4287);
nor UO_317 (O_317,N_2949,N_4599);
nor UO_318 (O_318,N_3886,N_4503);
nor UO_319 (O_319,N_3797,N_3706);
nand UO_320 (O_320,N_3350,N_4634);
nand UO_321 (O_321,N_3753,N_4531);
nand UO_322 (O_322,N_3379,N_2943);
xor UO_323 (O_323,N_4213,N_3188);
nand UO_324 (O_324,N_3885,N_4739);
and UO_325 (O_325,N_2688,N_3596);
xnor UO_326 (O_326,N_3993,N_3810);
nor UO_327 (O_327,N_2689,N_4134);
nor UO_328 (O_328,N_4661,N_4322);
or UO_329 (O_329,N_4754,N_4750);
or UO_330 (O_330,N_3044,N_3668);
and UO_331 (O_331,N_2786,N_4230);
and UO_332 (O_332,N_4341,N_2722);
nor UO_333 (O_333,N_2700,N_2770);
nand UO_334 (O_334,N_3833,N_4357);
or UO_335 (O_335,N_3125,N_2788);
nand UO_336 (O_336,N_2598,N_4893);
and UO_337 (O_337,N_2685,N_3141);
nand UO_338 (O_338,N_2627,N_4902);
and UO_339 (O_339,N_3004,N_4294);
xnor UO_340 (O_340,N_3571,N_4534);
and UO_341 (O_341,N_4309,N_3134);
nand UO_342 (O_342,N_2657,N_3717);
and UO_343 (O_343,N_3869,N_3539);
nand UO_344 (O_344,N_4448,N_4359);
nand UO_345 (O_345,N_3600,N_4766);
and UO_346 (O_346,N_4241,N_4415);
nand UO_347 (O_347,N_3777,N_4140);
or UO_348 (O_348,N_4491,N_4727);
nor UO_349 (O_349,N_2936,N_3185);
or UO_350 (O_350,N_4325,N_2803);
and UO_351 (O_351,N_2772,N_3529);
or UO_352 (O_352,N_3331,N_3297);
or UO_353 (O_353,N_4946,N_2680);
nand UO_354 (O_354,N_3392,N_2882);
and UO_355 (O_355,N_2605,N_3303);
nand UO_356 (O_356,N_3954,N_2606);
nor UO_357 (O_357,N_4388,N_2506);
nand UO_358 (O_358,N_4670,N_2871);
and UO_359 (O_359,N_3062,N_3216);
nor UO_360 (O_360,N_2622,N_4764);
nor UO_361 (O_361,N_4165,N_4950);
and UO_362 (O_362,N_4350,N_4070);
or UO_363 (O_363,N_3770,N_3991);
or UO_364 (O_364,N_3073,N_4568);
nand UO_365 (O_365,N_2523,N_4872);
nand UO_366 (O_366,N_4975,N_4967);
or UO_367 (O_367,N_4569,N_4065);
nand UO_368 (O_368,N_3516,N_2543);
nand UO_369 (O_369,N_3041,N_3311);
nand UO_370 (O_370,N_2857,N_3414);
or UO_371 (O_371,N_3075,N_4755);
or UO_372 (O_372,N_3957,N_3608);
nand UO_373 (O_373,N_2780,N_2636);
and UO_374 (O_374,N_4960,N_2776);
or UO_375 (O_375,N_2873,N_3918);
and UO_376 (O_376,N_2824,N_4492);
or UO_377 (O_377,N_4742,N_3160);
and UO_378 (O_378,N_3219,N_3949);
nand UO_379 (O_379,N_3533,N_4898);
nand UO_380 (O_380,N_3656,N_4077);
and UO_381 (O_381,N_3953,N_3555);
and UO_382 (O_382,N_3929,N_4680);
nor UO_383 (O_383,N_3236,N_4539);
xor UO_384 (O_384,N_4684,N_3913);
nor UO_385 (O_385,N_2522,N_3634);
and UO_386 (O_386,N_3265,N_4721);
or UO_387 (O_387,N_4034,N_3823);
and UO_388 (O_388,N_3282,N_4499);
nor UO_389 (O_389,N_4444,N_3686);
nor UO_390 (O_390,N_3611,N_3304);
nand UO_391 (O_391,N_3511,N_4657);
nor UO_392 (O_392,N_3523,N_3077);
nor UO_393 (O_393,N_2667,N_3784);
or UO_394 (O_394,N_4573,N_4855);
nand UO_395 (O_395,N_4029,N_4604);
nor UO_396 (O_396,N_3711,N_3530);
nand UO_397 (O_397,N_4117,N_4174);
nand UO_398 (O_398,N_3924,N_3750);
nand UO_399 (O_399,N_4297,N_4697);
nor UO_400 (O_400,N_2914,N_3992);
nand UO_401 (O_401,N_4921,N_4394);
or UO_402 (O_402,N_3124,N_2682);
or UO_403 (O_403,N_2530,N_4500);
and UO_404 (O_404,N_4033,N_4987);
or UO_405 (O_405,N_4945,N_4164);
or UO_406 (O_406,N_3373,N_4453);
and UO_407 (O_407,N_2911,N_4369);
and UO_408 (O_408,N_2541,N_3316);
or UO_409 (O_409,N_4074,N_2892);
and UO_410 (O_410,N_2832,N_4562);
and UO_411 (O_411,N_3255,N_3898);
nand UO_412 (O_412,N_4701,N_4104);
and UO_413 (O_413,N_4840,N_2654);
and UO_414 (O_414,N_4187,N_4526);
and UO_415 (O_415,N_2652,N_2988);
nor UO_416 (O_416,N_3624,N_2784);
or UO_417 (O_417,N_3513,N_3819);
nand UO_418 (O_418,N_2950,N_2872);
or UO_419 (O_419,N_3905,N_3767);
nor UO_420 (O_420,N_3139,N_3493);
nand UO_421 (O_421,N_3986,N_2568);
nand UO_422 (O_422,N_4374,N_4152);
and UO_423 (O_423,N_3249,N_4948);
nor UO_424 (O_424,N_3769,N_4794);
and UO_425 (O_425,N_3875,N_2809);
or UO_426 (O_426,N_3950,N_3199);
or UO_427 (O_427,N_4694,N_4882);
and UO_428 (O_428,N_3605,N_3293);
nor UO_429 (O_429,N_4223,N_4812);
or UO_430 (O_430,N_2757,N_3710);
xnor UO_431 (O_431,N_2900,N_3696);
and UO_432 (O_432,N_3071,N_4040);
nand UO_433 (O_433,N_4326,N_3369);
or UO_434 (O_434,N_4712,N_3749);
and UO_435 (O_435,N_3556,N_3677);
xor UO_436 (O_436,N_4585,N_4012);
or UO_437 (O_437,N_4028,N_2887);
and UO_438 (O_438,N_2880,N_4126);
and UO_439 (O_439,N_4785,N_3250);
nor UO_440 (O_440,N_4072,N_2777);
and UO_441 (O_441,N_3794,N_4011);
nand UO_442 (O_442,N_3925,N_3287);
nand UO_443 (O_443,N_2825,N_4784);
xor UO_444 (O_444,N_2585,N_4450);
nand UO_445 (O_445,N_3659,N_3532);
or UO_446 (O_446,N_4833,N_4757);
nand UO_447 (O_447,N_3120,N_2846);
or UO_448 (O_448,N_4268,N_4844);
nand UO_449 (O_449,N_3274,N_3171);
nand UO_450 (O_450,N_3179,N_3574);
or UO_451 (O_451,N_4300,N_3615);
and UO_452 (O_452,N_2978,N_4728);
nor UO_453 (O_453,N_4687,N_4335);
or UO_454 (O_454,N_4892,N_3942);
nand UO_455 (O_455,N_3494,N_3802);
and UO_456 (O_456,N_3483,N_4824);
nor UO_457 (O_457,N_4280,N_4947);
nor UO_458 (O_458,N_3195,N_3563);
nor UO_459 (O_459,N_3238,N_4256);
and UO_460 (O_460,N_2564,N_2527);
nor UO_461 (O_461,N_4480,N_4013);
nand UO_462 (O_462,N_4970,N_4400);
nor UO_463 (O_463,N_4689,N_3258);
nand UO_464 (O_464,N_3747,N_4682);
or UO_465 (O_465,N_4780,N_4472);
or UO_466 (O_466,N_3718,N_4506);
or UO_467 (O_467,N_2850,N_3256);
xnor UO_468 (O_468,N_3809,N_2521);
and UO_469 (O_469,N_4402,N_4501);
nor UO_470 (O_470,N_4969,N_3746);
or UO_471 (O_471,N_2713,N_3897);
and UO_472 (O_472,N_4155,N_2731);
nor UO_473 (O_473,N_3482,N_4930);
nand UO_474 (O_474,N_2964,N_4158);
nand UO_475 (O_475,N_3368,N_2816);
and UO_476 (O_476,N_4722,N_2712);
nand UO_477 (O_477,N_4956,N_4560);
or UO_478 (O_478,N_3681,N_4900);
and UO_479 (O_479,N_3095,N_4818);
xor UO_480 (O_480,N_4990,N_3514);
nor UO_481 (O_481,N_3908,N_3110);
or UO_482 (O_482,N_4984,N_4052);
or UO_483 (O_483,N_4664,N_3568);
nor UO_484 (O_484,N_3683,N_3729);
nand UO_485 (O_485,N_4008,N_3850);
or UO_486 (O_486,N_3721,N_3257);
nand UO_487 (O_487,N_2510,N_4723);
nand UO_488 (O_488,N_4460,N_4596);
or UO_489 (O_489,N_2612,N_4377);
and UO_490 (O_490,N_3059,N_3183);
or UO_491 (O_491,N_4207,N_2599);
nand UO_492 (O_492,N_4233,N_2618);
nand UO_493 (O_493,N_4825,N_4316);
nand UO_494 (O_494,N_3881,N_4073);
or UO_495 (O_495,N_3176,N_4598);
and UO_496 (O_496,N_3879,N_3305);
nand UO_497 (O_497,N_4363,N_2890);
nand UO_498 (O_498,N_3945,N_4048);
nor UO_499 (O_499,N_2843,N_4128);
nand UO_500 (O_500,N_3034,N_3010);
nor UO_501 (O_501,N_2739,N_3352);
and UO_502 (O_502,N_4913,N_3921);
nand UO_503 (O_503,N_4811,N_3764);
and UO_504 (O_504,N_3990,N_4808);
or UO_505 (O_505,N_4085,N_3799);
nand UO_506 (O_506,N_3919,N_4038);
and UO_507 (O_507,N_4962,N_4588);
or UO_508 (O_508,N_3313,N_3859);
nor UO_509 (O_509,N_3003,N_4735);
and UO_510 (O_510,N_4166,N_3023);
or UO_511 (O_511,N_4730,N_3628);
nor UO_512 (O_512,N_2796,N_3464);
and UO_513 (O_513,N_4889,N_4708);
nand UO_514 (O_514,N_4905,N_4929);
and UO_515 (O_515,N_4488,N_3295);
nor UO_516 (O_516,N_4151,N_4110);
and UO_517 (O_517,N_3348,N_2810);
or UO_518 (O_518,N_2576,N_4386);
or UO_519 (O_519,N_4094,N_2879);
nor UO_520 (O_520,N_2831,N_2792);
nand UO_521 (O_521,N_4610,N_4046);
or UO_522 (O_522,N_4182,N_2984);
nand UO_523 (O_523,N_4509,N_4275);
nand UO_524 (O_524,N_3858,N_4869);
nand UO_525 (O_525,N_2928,N_2544);
nand UO_526 (O_526,N_3456,N_4274);
nand UO_527 (O_527,N_2858,N_4457);
and UO_528 (O_528,N_3162,N_4655);
nand UO_529 (O_529,N_3772,N_4938);
nor UO_530 (O_530,N_4380,N_3068);
or UO_531 (O_531,N_3412,N_3844);
nand UO_532 (O_532,N_4648,N_3083);
or UO_533 (O_533,N_3760,N_4410);
or UO_534 (O_534,N_3462,N_3707);
nor UO_535 (O_535,N_2793,N_3679);
or UO_536 (O_536,N_3436,N_3994);
xor UO_537 (O_537,N_4988,N_4246);
or UO_538 (O_538,N_3480,N_4693);
or UO_539 (O_539,N_3515,N_4510);
nand UO_540 (O_540,N_4835,N_4917);
or UO_541 (O_541,N_2590,N_3666);
nor UO_542 (O_542,N_4853,N_4147);
nor UO_543 (O_543,N_4191,N_4066);
and UO_544 (O_544,N_4606,N_3864);
nor UO_545 (O_545,N_3739,N_3626);
and UO_546 (O_546,N_3420,N_4848);
nor UO_547 (O_547,N_4995,N_4199);
and UO_548 (O_548,N_4200,N_4931);
nor UO_549 (O_549,N_3008,N_3281);
and UO_550 (O_550,N_4736,N_2909);
xor UO_551 (O_551,N_4007,N_3254);
nor UO_552 (O_552,N_4586,N_4927);
nor UO_553 (O_553,N_3377,N_2797);
nand UO_554 (O_554,N_2631,N_3218);
and UO_555 (O_555,N_4051,N_2658);
or UO_556 (O_556,N_2990,N_3722);
and UO_557 (O_557,N_3671,N_4858);
or UO_558 (O_558,N_3604,N_2942);
nand UO_559 (O_559,N_2877,N_3226);
nand UO_560 (O_560,N_3093,N_3029);
and UO_561 (O_561,N_4552,N_3709);
and UO_562 (O_562,N_2946,N_3759);
nand UO_563 (O_563,N_2791,N_4571);
and UO_564 (O_564,N_4870,N_4049);
nand UO_565 (O_565,N_3082,N_3733);
nor UO_566 (O_566,N_4263,N_3969);
nand UO_567 (O_567,N_2562,N_2848);
and UO_568 (O_568,N_4266,N_4732);
xnor UO_569 (O_569,N_3277,N_4797);
or UO_570 (O_570,N_2932,N_2938);
xor UO_571 (O_571,N_3963,N_4514);
and UO_572 (O_572,N_4146,N_3536);
xor UO_573 (O_573,N_3106,N_4212);
or UO_574 (O_574,N_2581,N_3345);
nor UO_575 (O_575,N_3131,N_3334);
or UO_576 (O_576,N_3712,N_3448);
nand UO_577 (O_577,N_4837,N_3901);
nand UO_578 (O_578,N_3724,N_3353);
or UO_579 (O_579,N_4594,N_3595);
or UO_580 (O_580,N_3341,N_2787);
nor UO_581 (O_581,N_3289,N_4180);
and UO_582 (O_582,N_3013,N_4587);
or UO_583 (O_583,N_4906,N_3112);
or UO_584 (O_584,N_3136,N_3589);
nand UO_585 (O_585,N_3000,N_4150);
nor UO_586 (O_586,N_4418,N_4083);
and UO_587 (O_587,N_3165,N_4079);
nand UO_588 (O_588,N_4994,N_2526);
nand UO_589 (O_589,N_3447,N_4370);
nor UO_590 (O_590,N_3903,N_4261);
nor UO_591 (O_591,N_4115,N_3519);
nor UO_592 (O_592,N_2574,N_3966);
or UO_593 (O_593,N_3088,N_4434);
and UO_594 (O_594,N_4204,N_3632);
nand UO_595 (O_595,N_3205,N_3481);
nand UO_596 (O_596,N_4366,N_3097);
nand UO_597 (O_597,N_2516,N_2997);
nand UO_598 (O_598,N_4237,N_3193);
nand UO_599 (O_599,N_4656,N_3049);
or UO_600 (O_600,N_3882,N_4603);
nand UO_601 (O_601,N_2572,N_4107);
or UO_602 (O_602,N_4665,N_4382);
nand UO_603 (O_603,N_3801,N_2823);
and UO_604 (O_604,N_3224,N_4511);
and UO_605 (O_605,N_3820,N_4519);
and UO_606 (O_606,N_3298,N_4737);
nand UO_607 (O_607,N_3726,N_3432);
nor UO_608 (O_608,N_3367,N_2678);
nor UO_609 (O_609,N_4590,N_4206);
nor UO_610 (O_610,N_4978,N_4941);
nand UO_611 (O_611,N_4553,N_2865);
and UO_612 (O_612,N_2588,N_4337);
nor UO_613 (O_613,N_4801,N_4429);
and UO_614 (O_614,N_3793,N_3610);
and UO_615 (O_615,N_3197,N_3357);
nor UO_616 (O_616,N_2800,N_2659);
nand UO_617 (O_617,N_3598,N_2619);
or UO_618 (O_618,N_3518,N_4177);
nand UO_619 (O_619,N_3663,N_3786);
or UO_620 (O_620,N_3525,N_4496);
nor UO_621 (O_621,N_2986,N_2704);
or UO_622 (O_622,N_2910,N_3388);
and UO_623 (O_623,N_2724,N_3871);
and UO_624 (O_624,N_3554,N_4957);
nand UO_625 (O_625,N_4763,N_4815);
nor UO_626 (O_626,N_3878,N_4057);
or UO_627 (O_627,N_3441,N_2625);
nand UO_628 (O_628,N_3102,N_2901);
nand UO_629 (O_629,N_3319,N_2528);
nand UO_630 (O_630,N_3099,N_3621);
nor UO_631 (O_631,N_3116,N_3487);
or UO_632 (O_632,N_3471,N_4685);
nand UO_633 (O_633,N_2740,N_4993);
nor UO_634 (O_634,N_4579,N_3239);
or UO_635 (O_635,N_3064,N_3932);
and UO_636 (O_636,N_3616,N_4976);
or UO_637 (O_637,N_3870,N_3362);
nand UO_638 (O_638,N_4075,N_3290);
or UO_639 (O_639,N_3940,N_2790);
or UO_640 (O_640,N_3948,N_4832);
or UO_641 (O_641,N_2995,N_4302);
and UO_642 (O_642,N_4056,N_3505);
nor UO_643 (O_643,N_2737,N_3009);
or UO_644 (O_644,N_3891,N_4396);
nor UO_645 (O_645,N_2769,N_3232);
and UO_646 (O_646,N_4449,N_4211);
nand UO_647 (O_647,N_3390,N_4654);
or UO_648 (O_648,N_3055,N_4773);
nand UO_649 (O_649,N_4483,N_3065);
and UO_650 (O_650,N_4138,N_4095);
nand UO_651 (O_651,N_3984,N_2993);
nor UO_652 (O_652,N_2973,N_2959);
nor UO_653 (O_653,N_2802,N_2730);
or UO_654 (O_654,N_3468,N_3958);
and UO_655 (O_655,N_4103,N_3328);
xor UO_656 (O_656,N_4157,N_2808);
nand UO_657 (O_657,N_3385,N_4365);
nor UO_658 (O_658,N_3096,N_3923);
or UO_659 (O_659,N_3938,N_3450);
nand UO_660 (O_660,N_2775,N_3343);
or UO_661 (O_661,N_3400,N_4683);
or UO_662 (O_662,N_3322,N_4630);
and UO_663 (O_663,N_4817,N_3469);
or UO_664 (O_664,N_3426,N_2941);
nor UO_665 (O_665,N_3457,N_3306);
nor UO_666 (O_666,N_3358,N_3569);
or UO_667 (O_667,N_3911,N_4875);
and UO_668 (O_668,N_4841,N_3731);
and UO_669 (O_669,N_4475,N_3597);
and UO_670 (O_670,N_4992,N_4979);
or UO_671 (O_671,N_2806,N_3229);
or UO_672 (O_672,N_4286,N_2532);
nand UO_673 (O_673,N_2707,N_2818);
nand UO_674 (O_674,N_4706,N_3684);
and UO_675 (O_675,N_4215,N_3060);
nand UO_676 (O_676,N_3187,N_3558);
and UO_677 (O_677,N_3166,N_2921);
and UO_678 (O_678,N_3547,N_3424);
nor UO_679 (O_679,N_2874,N_4130);
nor UO_680 (O_680,N_3233,N_4068);
and UO_681 (O_681,N_3323,N_2799);
nor UO_682 (O_682,N_3454,N_3890);
nor UO_683 (O_683,N_2681,N_2687);
nor UO_684 (O_684,N_4716,N_2883);
nand UO_685 (O_685,N_4762,N_4025);
and UO_686 (O_686,N_4983,N_4351);
and UO_687 (O_687,N_4786,N_4847);
nor UO_688 (O_688,N_4462,N_4493);
or UO_689 (O_689,N_3344,N_2591);
nand UO_690 (O_690,N_3977,N_3132);
nand UO_691 (O_691,N_3742,N_3237);
nand UO_692 (O_692,N_3024,N_3933);
nor UO_693 (O_693,N_3788,N_4427);
and UO_694 (O_694,N_3466,N_3018);
nand UO_695 (O_695,N_4822,N_3164);
nand UO_696 (O_696,N_2648,N_4558);
or UO_697 (O_697,N_2935,N_2945);
or UO_698 (O_698,N_3653,N_3461);
nor UO_699 (O_699,N_3418,N_4173);
and UO_700 (O_700,N_4283,N_2726);
and UO_701 (O_701,N_3593,N_4720);
and UO_702 (O_702,N_3128,N_3916);
or UO_703 (O_703,N_2525,N_2644);
and UO_704 (O_704,N_4320,N_3261);
and UO_705 (O_705,N_2717,N_4796);
nor UO_706 (O_706,N_2602,N_3084);
xor UO_707 (O_707,N_3970,N_3192);
nor UO_708 (O_708,N_3548,N_3863);
and UO_709 (O_709,N_4580,N_4422);
and UO_710 (O_710,N_3834,N_3658);
nor UO_711 (O_711,N_4512,N_4319);
nor UO_712 (O_712,N_3403,N_2954);
nand UO_713 (O_713,N_4821,N_2912);
nand UO_714 (O_714,N_4027,N_3080);
and UO_715 (O_715,N_3643,N_4055);
nor UO_716 (O_716,N_4133,N_3081);
nor UO_717 (O_717,N_4356,N_2761);
nor UO_718 (O_718,N_3873,N_3324);
or UO_719 (O_719,N_4023,N_3727);
nor UO_720 (O_720,N_3583,N_2609);
and UO_721 (O_721,N_3865,N_4924);
and UO_722 (O_722,N_3776,N_4868);
and UO_723 (O_723,N_4355,N_3340);
and UO_724 (O_724,N_4567,N_3758);
and UO_725 (O_725,N_4502,N_3965);
or UO_726 (O_726,N_4178,N_4141);
and UO_727 (O_727,N_3428,N_4761);
and UO_728 (O_728,N_2552,N_4795);
xor UO_729 (O_729,N_4883,N_3072);
or UO_730 (O_730,N_3839,N_2519);
nor UO_731 (O_731,N_3531,N_4148);
nor UO_732 (O_732,N_4628,N_3650);
nor UO_733 (O_733,N_4210,N_3002);
nor UO_734 (O_734,N_3821,N_2829);
or UO_735 (O_735,N_4464,N_2753);
nor UO_736 (O_736,N_4249,N_3251);
and UO_737 (O_737,N_4515,N_3202);
or UO_738 (O_738,N_2684,N_4214);
or UO_739 (O_739,N_2666,N_3868);
xnor UO_740 (O_740,N_4642,N_2643);
or UO_741 (O_741,N_4774,N_2694);
nor UO_742 (O_742,N_4315,N_4804);
and UO_743 (O_743,N_3242,N_4986);
or UO_744 (O_744,N_4486,N_3876);
nand UO_745 (O_745,N_2698,N_3020);
or UO_746 (O_746,N_4617,N_4860);
nor UO_747 (O_747,N_4636,N_3528);
and UO_748 (O_748,N_4542,N_4915);
nor UO_749 (O_749,N_3217,N_3620);
nor UO_750 (O_750,N_4017,N_2638);
or UO_751 (O_751,N_2881,N_4696);
nor UO_752 (O_752,N_4445,N_2639);
nor UO_753 (O_753,N_4867,N_2547);
or UO_754 (O_754,N_3685,N_3856);
and UO_755 (O_755,N_3154,N_4433);
nand UO_756 (O_756,N_3551,N_3366);
nor UO_757 (O_757,N_3592,N_4293);
nor UO_758 (O_758,N_2504,N_3066);
or UO_759 (O_759,N_2937,N_3914);
nand UO_760 (O_760,N_4096,N_4381);
nor UO_761 (O_761,N_3736,N_4544);
nor UO_762 (O_762,N_4545,N_4467);
nor UO_763 (O_763,N_3138,N_2672);
nand UO_764 (O_764,N_3781,N_3818);
nor UO_765 (O_765,N_2719,N_3408);
or UO_766 (O_766,N_3026,N_2662);
xnor UO_767 (O_767,N_2982,N_2531);
nand UO_768 (O_768,N_4688,N_4354);
nor UO_769 (O_769,N_4423,N_3694);
and UO_770 (O_770,N_3698,N_3761);
nor UO_771 (O_771,N_4234,N_4089);
nand UO_772 (O_772,N_4198,N_4321);
nand UO_773 (O_773,N_4411,N_3735);
nor UO_774 (O_774,N_4059,N_4375);
and UO_775 (O_775,N_2838,N_3791);
nand UO_776 (O_776,N_3732,N_3317);
xor UO_777 (O_777,N_4119,N_4678);
nor UO_778 (O_778,N_3500,N_3021);
nor UO_779 (O_779,N_3266,N_4806);
nor UO_780 (O_780,N_3789,N_4123);
nand UO_781 (O_781,N_2582,N_4624);
nor UO_782 (O_782,N_2554,N_3636);
or UO_783 (O_783,N_4884,N_3063);
and UO_784 (O_784,N_3614,N_3599);
and UO_785 (O_785,N_3061,N_4595);
nand UO_786 (O_786,N_2634,N_3045);
and UO_787 (O_787,N_3039,N_4303);
nor UO_788 (O_788,N_4934,N_2860);
and UO_789 (O_789,N_3852,N_4813);
and UO_790 (O_790,N_3339,N_2956);
and UO_791 (O_791,N_2570,N_4842);
nor UO_792 (O_792,N_4614,N_3335);
nor UO_793 (O_793,N_3108,N_4168);
nor UO_794 (O_794,N_3499,N_4333);
and UO_795 (O_795,N_2675,N_4899);
or UO_796 (O_796,N_3210,N_4346);
nor UO_797 (O_797,N_3774,N_2655);
nor UO_798 (O_798,N_3887,N_4578);
or UO_799 (O_799,N_4203,N_3825);
or UO_800 (O_800,N_4770,N_4777);
nand UO_801 (O_801,N_4391,N_3645);
and UO_802 (O_802,N_4904,N_2855);
nor UO_803 (O_803,N_4430,N_4473);
nand UO_804 (O_804,N_4190,N_2840);
nand UO_805 (O_805,N_3617,N_4384);
nand UO_806 (O_806,N_2987,N_2725);
xnor UO_807 (O_807,N_3775,N_2661);
and UO_808 (O_808,N_2795,N_3417);
nor UO_809 (O_809,N_4485,N_3433);
and UO_810 (O_810,N_2548,N_3067);
or UO_811 (O_811,N_3275,N_3883);
and UO_812 (O_812,N_4647,N_2925);
and UO_813 (O_813,N_4963,N_4856);
and UO_814 (O_814,N_2981,N_4225);
nor UO_815 (O_815,N_2812,N_3688);
nor UO_816 (O_816,N_4163,N_2804);
nand UO_817 (O_817,N_2540,N_4877);
and UO_818 (O_818,N_2586,N_3186);
nand UO_819 (O_819,N_3017,N_4436);
nor UO_820 (O_820,N_3245,N_4760);
and UO_821 (O_821,N_4974,N_4005);
nor UO_822 (O_822,N_4922,N_4756);
or UO_823 (O_823,N_3524,N_3391);
and UO_824 (O_824,N_3754,N_3147);
or UO_825 (O_825,N_3091,N_4718);
and UO_826 (O_826,N_4487,N_4555);
or UO_827 (O_827,N_3651,N_3485);
nand UO_828 (O_828,N_4903,N_3817);
xor UO_829 (O_829,N_3826,N_2561);
or UO_830 (O_830,N_4463,N_2748);
and UO_831 (O_831,N_4897,N_2705);
nand UO_832 (O_832,N_3931,N_4803);
nor UO_833 (O_833,N_3606,N_3590);
or UO_834 (O_834,N_2580,N_4383);
or UO_835 (O_835,N_4461,N_3458);
and UO_836 (O_836,N_4949,N_3831);
and UO_837 (O_837,N_2710,N_3419);
nand UO_838 (O_838,N_4442,N_4113);
or UO_839 (O_839,N_3365,N_3550);
nand UO_840 (O_840,N_3384,N_2926);
or UO_841 (O_841,N_2920,N_3692);
nand UO_842 (O_842,N_2960,N_4920);
or UO_843 (O_843,N_3273,N_3007);
or UO_844 (O_844,N_3838,N_4149);
and UO_845 (O_845,N_3541,N_3372);
xnor UO_846 (O_846,N_3425,N_2947);
nand UO_847 (O_847,N_4482,N_4846);
nor UO_848 (O_848,N_4220,N_3393);
xnor UO_849 (O_849,N_3030,N_4668);
nor UO_850 (O_850,N_4726,N_4116);
or UO_851 (O_851,N_4626,N_4699);
or UO_852 (O_852,N_2835,N_3807);
nand UO_853 (O_853,N_4387,N_4549);
and UO_854 (O_854,N_3264,N_4575);
nor UO_855 (O_855,N_3877,N_2758);
and UO_856 (O_856,N_4782,N_3122);
or UO_857 (O_857,N_4443,N_2558);
and UO_858 (O_858,N_4295,N_4940);
and UO_859 (O_859,N_4125,N_4707);
nand UO_860 (O_860,N_3198,N_2692);
or UO_861 (O_861,N_4751,N_3888);
nor UO_862 (O_862,N_4100,N_3828);
nand UO_863 (O_863,N_4620,N_4061);
nand UO_864 (O_864,N_3015,N_4238);
nor UO_865 (O_865,N_4264,N_2640);
nor UO_866 (O_866,N_3427,N_4916);
and UO_867 (O_867,N_4533,N_3737);
and UO_868 (O_868,N_4171,N_3490);
nand UO_869 (O_869,N_4528,N_3889);
nor UO_870 (O_870,N_3387,N_4284);
xor UO_871 (O_871,N_3840,N_4189);
nand UO_872 (O_872,N_3522,N_4307);
or UO_873 (O_873,N_4671,N_4205);
nor UO_874 (O_874,N_2884,N_2759);
nor UO_875 (O_875,N_4508,N_2755);
nor UO_876 (O_876,N_4758,N_4646);
nand UO_877 (O_877,N_2847,N_3338);
or UO_878 (O_878,N_4153,N_4044);
xor UO_879 (O_879,N_2839,N_3470);
or UO_880 (O_880,N_3294,N_4367);
nand UO_881 (O_881,N_3900,N_4019);
nor UO_882 (O_882,N_4014,N_4775);
and UO_883 (O_883,N_3655,N_4431);
and UO_884 (O_884,N_3983,N_4306);
nor UO_885 (O_885,N_4933,N_4788);
nor UO_886 (O_886,N_3460,N_4030);
nor UO_887 (O_887,N_3016,N_2534);
nor UO_888 (O_888,N_4439,N_3260);
nand UO_889 (O_889,N_2955,N_3682);
or UO_890 (O_890,N_2614,N_3475);
or UO_891 (O_891,N_2905,N_4186);
nand UO_892 (O_892,N_2827,N_4998);
nor UO_893 (O_893,N_2996,N_2676);
nor UO_894 (O_894,N_4935,N_2555);
or UO_895 (O_895,N_3849,N_3619);
and UO_896 (O_896,N_2610,N_3300);
nand UO_897 (O_897,N_4537,N_2728);
xor UO_898 (O_898,N_4944,N_2641);
or UO_899 (O_899,N_3678,N_3119);
nor UO_900 (O_900,N_4543,N_2584);
nor UO_901 (O_901,N_4724,N_4122);
nor UO_902 (O_902,N_3581,N_4827);
nor UO_903 (O_903,N_3477,N_4741);
nand UO_904 (O_904,N_2815,N_3248);
or UO_905 (O_905,N_4809,N_3225);
nor UO_906 (O_906,N_2977,N_4226);
nand UO_907 (O_907,N_4566,N_3411);
and UO_908 (O_908,N_3702,N_4231);
and UO_909 (O_909,N_2927,N_4719);
and UO_910 (O_910,N_3824,N_3336);
nand UO_911 (O_911,N_3830,N_4368);
nand UO_912 (O_912,N_3127,N_3586);
and UO_913 (O_913,N_3982,N_2751);
nand UO_914 (O_914,N_4793,N_4127);
nor UO_915 (O_915,N_3542,N_4454);
nand UO_916 (O_916,N_4955,N_2579);
and UO_917 (O_917,N_4879,N_4455);
nand UO_918 (O_918,N_3451,N_4641);
nand UO_919 (O_919,N_3401,N_2703);
and UO_920 (O_920,N_4451,N_2538);
or UO_921 (O_921,N_2878,N_3473);
and UO_922 (O_922,N_3405,N_2613);
and UO_923 (O_923,N_4236,N_2833);
nand UO_924 (O_924,N_4673,N_3501);
or UO_925 (O_925,N_4767,N_2592);
and UO_926 (O_926,N_3156,N_3647);
and UO_927 (O_927,N_3570,N_4441);
or UO_928 (O_928,N_3565,N_2963);
nand UO_929 (O_929,N_3145,N_4197);
or UO_930 (O_930,N_2595,N_3703);
nand UO_931 (O_931,N_2767,N_2577);
nor UO_932 (O_932,N_4270,N_4064);
or UO_933 (O_933,N_3276,N_3038);
and UO_934 (O_934,N_2762,N_4218);
or UO_935 (O_935,N_4112,N_4667);
or UO_936 (O_936,N_4863,N_4880);
nand UO_937 (O_937,N_3884,N_3042);
and UO_938 (O_938,N_2604,N_4026);
nand UO_939 (O_939,N_3492,N_3221);
nor UO_940 (O_940,N_4323,N_3263);
nor UO_941 (O_941,N_3247,N_3537);
or UO_942 (O_942,N_3787,N_2798);
nand UO_943 (O_943,N_4221,N_2783);
nand UO_944 (O_944,N_3641,N_3996);
nand UO_945 (O_945,N_3545,N_2778);
and UO_946 (O_946,N_3714,N_4109);
nand UO_947 (O_947,N_3906,N_4358);
nand UO_948 (O_948,N_4267,N_4278);
and UO_949 (O_949,N_3445,N_4966);
nand UO_950 (O_950,N_4731,N_3376);
and UO_951 (O_951,N_2741,N_3951);
or UO_952 (O_952,N_2671,N_4006);
and UO_953 (O_953,N_3284,N_3520);
or UO_954 (O_954,N_4738,N_4202);
and UO_955 (O_955,N_2974,N_3054);
and UO_956 (O_956,N_3577,N_2669);
or UO_957 (O_957,N_4262,N_3035);
or UO_958 (O_958,N_3244,N_3434);
and UO_959 (O_959,N_4426,N_3827);
and UO_960 (O_960,N_3069,N_3904);
or UO_961 (O_961,N_3463,N_3133);
or UO_962 (O_962,N_4576,N_4589);
nor UO_963 (O_963,N_3078,N_2859);
nand UO_964 (O_964,N_3354,N_4494);
or UO_965 (O_965,N_2970,N_3926);
nor UO_966 (O_966,N_4020,N_3612);
or UO_967 (O_967,N_3360,N_3270);
and UO_968 (O_968,N_3406,N_4466);
nor UO_969 (O_969,N_2508,N_4894);
or UO_970 (O_970,N_4973,N_2853);
or UO_971 (O_971,N_3496,N_2515);
nand UO_972 (O_972,N_4111,N_4616);
nor UO_973 (O_973,N_4997,N_4981);
and UO_974 (O_974,N_3544,N_4035);
and UO_975 (O_975,N_2695,N_4686);
or UO_976 (O_976,N_2895,N_3798);
nor UO_977 (O_977,N_4819,N_2514);
or UO_978 (O_978,N_4865,N_2968);
nor UO_979 (O_979,N_3507,N_4659);
and UO_980 (O_980,N_3697,N_3307);
and UO_981 (O_981,N_3691,N_4800);
or UO_982 (O_982,N_3452,N_3579);
and UO_983 (O_983,N_2965,N_4170);
nand UO_984 (O_984,N_3155,N_3231);
or UO_985 (O_985,N_2535,N_3730);
nand UO_986 (O_986,N_3790,N_3561);
nor UO_987 (O_987,N_4339,N_4390);
or UO_988 (O_988,N_3431,N_2632);
and UO_989 (O_989,N_4612,N_3092);
or UO_990 (O_990,N_4649,N_2760);
or UO_991 (O_991,N_4277,N_4563);
and UO_992 (O_992,N_4002,N_2841);
nor UO_993 (O_993,N_3150,N_3987);
and UO_994 (O_994,N_3741,N_4961);
or UO_995 (O_995,N_3375,N_2716);
and UO_996 (O_996,N_3892,N_2903);
and UO_997 (O_997,N_4854,N_4272);
nor UO_998 (O_998,N_4050,N_4043);
and UO_999 (O_999,N_2630,N_3410);
endmodule