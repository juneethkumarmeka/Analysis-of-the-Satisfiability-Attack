module basic_500_3000_500_3_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_387,In_497);
and U1 (N_1,In_127,In_247);
or U2 (N_2,In_408,In_13);
nand U3 (N_3,In_280,In_205);
or U4 (N_4,In_19,In_499);
or U5 (N_5,In_403,In_150);
nand U6 (N_6,In_289,In_466);
nand U7 (N_7,In_250,In_172);
or U8 (N_8,In_154,In_382);
nand U9 (N_9,In_312,In_490);
nor U10 (N_10,In_310,In_0);
nor U11 (N_11,In_314,In_67);
xor U12 (N_12,In_158,In_396);
xnor U13 (N_13,In_422,In_75);
and U14 (N_14,In_462,In_376);
nand U15 (N_15,In_491,In_446);
nand U16 (N_16,In_366,In_121);
and U17 (N_17,In_156,In_231);
nand U18 (N_18,In_225,In_89);
nor U19 (N_19,In_404,In_116);
and U20 (N_20,In_284,In_311);
nand U21 (N_21,In_7,In_394);
nor U22 (N_22,In_61,In_431);
and U23 (N_23,In_409,In_418);
or U24 (N_24,In_174,In_399);
and U25 (N_25,In_458,In_463);
xnor U26 (N_26,In_182,In_465);
or U27 (N_27,In_306,In_370);
or U28 (N_28,In_361,In_270);
or U29 (N_29,In_375,In_371);
nor U30 (N_30,In_5,In_260);
xnor U31 (N_31,In_71,In_115);
xnor U32 (N_32,In_430,In_325);
or U33 (N_33,In_2,In_330);
nand U34 (N_34,In_484,In_288);
nand U35 (N_35,In_91,In_291);
nand U36 (N_36,In_272,In_50);
or U37 (N_37,In_294,In_14);
and U38 (N_38,In_295,In_444);
xor U39 (N_39,In_326,In_334);
nor U40 (N_40,In_1,In_357);
and U41 (N_41,In_238,In_134);
nor U42 (N_42,In_167,In_378);
and U43 (N_43,In_346,In_169);
xor U44 (N_44,In_364,In_384);
or U45 (N_45,In_253,In_34);
or U46 (N_46,In_259,In_307);
or U47 (N_47,In_338,In_128);
nor U48 (N_48,In_398,In_110);
nor U49 (N_49,In_243,In_226);
nor U50 (N_50,In_379,In_38);
nand U51 (N_51,In_482,In_35);
or U52 (N_52,In_57,In_281);
nand U53 (N_53,In_283,In_123);
and U54 (N_54,In_233,In_6);
and U55 (N_55,In_240,In_439);
nor U56 (N_56,In_470,In_406);
nor U57 (N_57,In_39,In_309);
or U58 (N_58,In_54,In_267);
and U59 (N_59,In_15,In_478);
nand U60 (N_60,In_447,In_493);
nand U61 (N_61,In_262,In_227);
nor U62 (N_62,In_355,In_70);
nand U63 (N_63,In_318,In_26);
and U64 (N_64,In_471,In_223);
nand U65 (N_65,In_488,In_323);
nand U66 (N_66,In_148,In_33);
and U67 (N_67,In_461,In_173);
xor U68 (N_68,In_141,In_219);
or U69 (N_69,In_441,In_383);
nand U70 (N_70,In_269,In_159);
and U71 (N_71,In_305,In_130);
nor U72 (N_72,In_152,In_160);
nand U73 (N_73,In_146,In_199);
nand U74 (N_74,In_189,In_339);
and U75 (N_75,In_392,In_393);
nor U76 (N_76,In_153,In_87);
nor U77 (N_77,In_230,In_98);
or U78 (N_78,In_131,In_390);
or U79 (N_79,In_194,In_195);
nand U80 (N_80,In_315,In_443);
xor U81 (N_81,In_356,In_46);
nor U82 (N_82,In_303,In_178);
nor U83 (N_83,In_363,In_229);
nor U84 (N_84,In_273,In_304);
nand U85 (N_85,In_486,In_336);
and U86 (N_86,In_248,In_135);
and U87 (N_87,In_63,In_456);
or U88 (N_88,In_348,In_96);
and U89 (N_89,In_433,In_22);
nor U90 (N_90,In_197,In_36);
and U91 (N_91,In_349,In_391);
nor U92 (N_92,In_145,In_28);
and U93 (N_93,In_165,In_236);
nand U94 (N_94,In_129,In_81);
and U95 (N_95,In_350,In_101);
or U96 (N_96,In_113,In_58);
or U97 (N_97,In_44,In_126);
and U98 (N_98,In_286,In_401);
xor U99 (N_99,In_193,In_221);
nand U100 (N_100,In_388,In_86);
xnor U101 (N_101,In_88,In_29);
or U102 (N_102,In_452,In_78);
xnor U103 (N_103,In_18,In_450);
nor U104 (N_104,In_360,In_457);
nor U105 (N_105,In_100,In_245);
or U106 (N_106,In_414,In_274);
or U107 (N_107,In_285,In_73);
nor U108 (N_108,In_140,In_296);
nand U109 (N_109,In_161,In_410);
or U110 (N_110,In_120,In_164);
or U111 (N_111,In_151,In_359);
nand U112 (N_112,In_454,In_32);
and U113 (N_113,In_125,In_282);
nor U114 (N_114,In_12,In_144);
nand U115 (N_115,In_142,In_251);
and U116 (N_116,In_483,In_157);
or U117 (N_117,In_302,In_438);
and U118 (N_118,In_149,In_464);
or U119 (N_119,In_48,In_90);
nor U120 (N_120,In_133,In_417);
xor U121 (N_121,In_354,In_440);
and U122 (N_122,In_147,In_389);
and U123 (N_123,In_42,In_220);
nor U124 (N_124,In_494,In_292);
and U125 (N_125,In_498,In_427);
or U126 (N_126,In_420,In_56);
and U127 (N_127,In_254,In_474);
and U128 (N_128,In_485,In_411);
or U129 (N_129,In_196,In_400);
nor U130 (N_130,In_137,In_386);
nor U131 (N_131,In_265,In_190);
nand U132 (N_132,In_143,In_343);
nand U133 (N_133,In_426,In_171);
nor U134 (N_134,In_425,In_489);
xor U135 (N_135,In_308,In_424);
and U136 (N_136,In_480,In_341);
or U137 (N_137,In_256,In_94);
or U138 (N_138,In_279,In_469);
nand U139 (N_139,In_210,In_271);
xnor U140 (N_140,In_419,In_316);
nand U141 (N_141,In_217,In_421);
nand U142 (N_142,In_397,In_79);
or U143 (N_143,In_324,In_367);
or U144 (N_144,In_211,In_185);
nand U145 (N_145,In_188,In_442);
nor U146 (N_146,In_429,In_290);
and U147 (N_147,In_170,In_402);
nor U148 (N_148,In_276,In_407);
or U149 (N_149,In_473,In_84);
or U150 (N_150,In_24,In_268);
nor U151 (N_151,In_53,In_132);
xor U152 (N_152,In_155,In_41);
or U153 (N_153,In_76,In_475);
and U154 (N_154,In_64,In_496);
or U155 (N_155,In_369,In_180);
nand U156 (N_156,In_168,In_299);
and U157 (N_157,In_460,In_83);
or U158 (N_158,In_412,In_329);
nor U159 (N_159,In_8,In_202);
nor U160 (N_160,In_106,In_455);
or U161 (N_161,In_432,In_492);
and U162 (N_162,In_213,In_206);
nand U163 (N_163,In_445,In_377);
and U164 (N_164,In_212,In_395);
nand U165 (N_165,In_416,In_112);
nor U166 (N_166,In_275,In_104);
xor U167 (N_167,In_21,In_82);
or U168 (N_168,In_413,In_244);
nand U169 (N_169,In_317,In_380);
and U170 (N_170,In_263,In_52);
nor U171 (N_171,In_252,In_72);
nor U172 (N_172,In_246,In_301);
or U173 (N_173,In_31,In_293);
nor U174 (N_174,In_374,In_258);
xnor U175 (N_175,In_179,In_477);
nor U176 (N_176,In_333,In_122);
or U177 (N_177,In_103,In_365);
and U178 (N_178,In_97,In_342);
nand U179 (N_179,In_467,In_49);
or U180 (N_180,In_249,In_228);
or U181 (N_181,In_320,In_40);
nor U182 (N_182,In_203,In_319);
nand U183 (N_183,In_11,In_321);
nand U184 (N_184,In_136,In_65);
and U185 (N_185,In_479,In_93);
or U186 (N_186,In_487,In_472);
or U187 (N_187,In_214,In_17);
nand U188 (N_188,In_80,In_138);
nor U189 (N_189,In_218,In_232);
and U190 (N_190,In_453,In_47);
or U191 (N_191,In_449,In_241);
and U192 (N_192,In_184,In_51);
xor U193 (N_193,In_266,In_175);
nor U194 (N_194,In_68,In_448);
and U195 (N_195,In_166,In_278);
and U196 (N_196,In_85,In_4);
xnor U197 (N_197,In_340,In_468);
and U198 (N_198,In_327,In_9);
or U199 (N_199,In_224,In_344);
xnor U200 (N_200,In_322,In_124);
and U201 (N_201,In_105,In_222);
or U202 (N_202,In_216,In_111);
and U203 (N_203,In_92,In_451);
and U204 (N_204,In_313,In_37);
or U205 (N_205,In_25,In_200);
xor U206 (N_206,In_353,In_331);
or U207 (N_207,In_352,In_255);
xor U208 (N_208,In_423,In_55);
nor U209 (N_209,In_235,In_69);
nand U210 (N_210,In_74,In_300);
and U211 (N_211,In_114,In_119);
nor U212 (N_212,In_207,In_345);
nor U213 (N_213,In_237,In_204);
xor U214 (N_214,In_20,In_437);
and U215 (N_215,In_62,In_381);
or U216 (N_216,In_27,In_95);
nand U217 (N_217,In_436,In_362);
and U218 (N_218,In_332,In_77);
xnor U219 (N_219,In_162,In_10);
or U220 (N_220,In_107,In_139);
nand U221 (N_221,In_385,In_234);
or U222 (N_222,In_335,In_261);
or U223 (N_223,In_459,In_23);
nand U224 (N_224,In_347,In_109);
nor U225 (N_225,In_30,In_43);
xor U226 (N_226,In_287,In_215);
nor U227 (N_227,In_208,In_264);
xnor U228 (N_228,In_177,In_66);
nor U229 (N_229,In_434,In_45);
or U230 (N_230,In_351,In_373);
and U231 (N_231,In_328,In_3);
nor U232 (N_232,In_186,In_476);
nand U233 (N_233,In_118,In_192);
and U234 (N_234,In_372,In_358);
xnor U235 (N_235,In_99,In_209);
and U236 (N_236,In_187,In_257);
nor U237 (N_237,In_428,In_117);
xor U238 (N_238,In_239,In_108);
nand U239 (N_239,In_298,In_198);
and U240 (N_240,In_415,In_176);
or U241 (N_241,In_337,In_191);
and U242 (N_242,In_481,In_102);
nor U243 (N_243,In_242,In_368);
xor U244 (N_244,In_201,In_405);
and U245 (N_245,In_163,In_435);
nor U246 (N_246,In_181,In_297);
xnor U247 (N_247,In_59,In_183);
and U248 (N_248,In_495,In_277);
nor U249 (N_249,In_16,In_60);
nor U250 (N_250,In_367,In_11);
nand U251 (N_251,In_470,In_218);
or U252 (N_252,In_271,In_52);
and U253 (N_253,In_479,In_154);
xnor U254 (N_254,In_2,In_302);
nor U255 (N_255,In_89,In_320);
and U256 (N_256,In_176,In_171);
nand U257 (N_257,In_354,In_2);
and U258 (N_258,In_240,In_341);
nand U259 (N_259,In_136,In_154);
xor U260 (N_260,In_33,In_62);
nor U261 (N_261,In_225,In_161);
or U262 (N_262,In_448,In_384);
nor U263 (N_263,In_393,In_176);
or U264 (N_264,In_262,In_35);
or U265 (N_265,In_70,In_68);
nor U266 (N_266,In_12,In_123);
or U267 (N_267,In_246,In_51);
nor U268 (N_268,In_255,In_17);
and U269 (N_269,In_42,In_231);
nand U270 (N_270,In_39,In_4);
nor U271 (N_271,In_471,In_33);
nor U272 (N_272,In_200,In_240);
and U273 (N_273,In_68,In_154);
nor U274 (N_274,In_196,In_269);
nand U275 (N_275,In_262,In_410);
or U276 (N_276,In_41,In_184);
nand U277 (N_277,In_63,In_381);
and U278 (N_278,In_424,In_198);
nor U279 (N_279,In_392,In_245);
xor U280 (N_280,In_72,In_54);
and U281 (N_281,In_420,In_94);
and U282 (N_282,In_375,In_212);
nand U283 (N_283,In_337,In_213);
xnor U284 (N_284,In_418,In_142);
or U285 (N_285,In_255,In_76);
and U286 (N_286,In_469,In_21);
nor U287 (N_287,In_305,In_330);
nand U288 (N_288,In_243,In_198);
nand U289 (N_289,In_411,In_217);
xnor U290 (N_290,In_243,In_49);
nor U291 (N_291,In_43,In_479);
nor U292 (N_292,In_360,In_312);
nand U293 (N_293,In_230,In_433);
nor U294 (N_294,In_317,In_196);
nor U295 (N_295,In_413,In_361);
and U296 (N_296,In_373,In_387);
nor U297 (N_297,In_0,In_28);
or U298 (N_298,In_123,In_1);
nor U299 (N_299,In_323,In_141);
or U300 (N_300,In_370,In_422);
nor U301 (N_301,In_9,In_3);
or U302 (N_302,In_57,In_265);
nand U303 (N_303,In_269,In_77);
or U304 (N_304,In_20,In_142);
or U305 (N_305,In_460,In_419);
or U306 (N_306,In_341,In_247);
nand U307 (N_307,In_23,In_246);
nor U308 (N_308,In_371,In_7);
xnor U309 (N_309,In_259,In_400);
xnor U310 (N_310,In_30,In_161);
or U311 (N_311,In_412,In_440);
nor U312 (N_312,In_107,In_96);
or U313 (N_313,In_282,In_327);
nor U314 (N_314,In_381,In_436);
and U315 (N_315,In_426,In_103);
or U316 (N_316,In_370,In_221);
and U317 (N_317,In_26,In_113);
or U318 (N_318,In_403,In_239);
or U319 (N_319,In_158,In_487);
nor U320 (N_320,In_227,In_213);
nor U321 (N_321,In_63,In_318);
nor U322 (N_322,In_127,In_353);
or U323 (N_323,In_99,In_387);
or U324 (N_324,In_381,In_149);
or U325 (N_325,In_432,In_276);
and U326 (N_326,In_25,In_243);
xnor U327 (N_327,In_492,In_53);
or U328 (N_328,In_185,In_468);
nor U329 (N_329,In_384,In_348);
nand U330 (N_330,In_236,In_354);
nor U331 (N_331,In_60,In_77);
and U332 (N_332,In_329,In_377);
and U333 (N_333,In_178,In_69);
and U334 (N_334,In_34,In_128);
nor U335 (N_335,In_52,In_162);
and U336 (N_336,In_231,In_99);
and U337 (N_337,In_403,In_23);
nand U338 (N_338,In_124,In_166);
or U339 (N_339,In_386,In_123);
nor U340 (N_340,In_266,In_452);
nand U341 (N_341,In_69,In_244);
nand U342 (N_342,In_219,In_16);
and U343 (N_343,In_228,In_285);
or U344 (N_344,In_154,In_441);
xnor U345 (N_345,In_309,In_236);
or U346 (N_346,In_358,In_279);
nand U347 (N_347,In_278,In_73);
nor U348 (N_348,In_62,In_47);
nor U349 (N_349,In_238,In_2);
and U350 (N_350,In_474,In_21);
nand U351 (N_351,In_385,In_291);
or U352 (N_352,In_168,In_93);
nor U353 (N_353,In_349,In_159);
nand U354 (N_354,In_136,In_138);
xnor U355 (N_355,In_262,In_408);
xor U356 (N_356,In_153,In_437);
and U357 (N_357,In_190,In_444);
nand U358 (N_358,In_248,In_357);
nor U359 (N_359,In_187,In_169);
or U360 (N_360,In_65,In_302);
xor U361 (N_361,In_353,In_490);
xnor U362 (N_362,In_16,In_194);
nor U363 (N_363,In_353,In_383);
xnor U364 (N_364,In_422,In_459);
nand U365 (N_365,In_44,In_284);
nand U366 (N_366,In_280,In_46);
or U367 (N_367,In_479,In_306);
and U368 (N_368,In_229,In_124);
or U369 (N_369,In_110,In_369);
nand U370 (N_370,In_282,In_212);
and U371 (N_371,In_143,In_320);
and U372 (N_372,In_228,In_241);
xnor U373 (N_373,In_445,In_149);
and U374 (N_374,In_477,In_457);
and U375 (N_375,In_200,In_157);
nand U376 (N_376,In_243,In_182);
nand U377 (N_377,In_440,In_459);
nand U378 (N_378,In_440,In_453);
and U379 (N_379,In_294,In_112);
and U380 (N_380,In_457,In_353);
nor U381 (N_381,In_282,In_438);
and U382 (N_382,In_403,In_443);
or U383 (N_383,In_307,In_352);
xnor U384 (N_384,In_271,In_269);
nand U385 (N_385,In_459,In_217);
xnor U386 (N_386,In_22,In_479);
nor U387 (N_387,In_72,In_468);
nand U388 (N_388,In_225,In_203);
or U389 (N_389,In_417,In_254);
nand U390 (N_390,In_371,In_466);
or U391 (N_391,In_330,In_389);
and U392 (N_392,In_413,In_393);
nand U393 (N_393,In_70,In_100);
nor U394 (N_394,In_240,In_97);
or U395 (N_395,In_154,In_266);
xor U396 (N_396,In_435,In_82);
or U397 (N_397,In_286,In_344);
xor U398 (N_398,In_82,In_76);
and U399 (N_399,In_454,In_128);
or U400 (N_400,In_204,In_492);
or U401 (N_401,In_397,In_413);
nor U402 (N_402,In_257,In_453);
nor U403 (N_403,In_307,In_383);
and U404 (N_404,In_233,In_390);
nor U405 (N_405,In_150,In_493);
nand U406 (N_406,In_378,In_25);
nor U407 (N_407,In_303,In_174);
and U408 (N_408,In_334,In_266);
nand U409 (N_409,In_75,In_44);
and U410 (N_410,In_378,In_227);
or U411 (N_411,In_254,In_161);
nand U412 (N_412,In_486,In_315);
or U413 (N_413,In_185,In_327);
nand U414 (N_414,In_173,In_66);
and U415 (N_415,In_490,In_360);
and U416 (N_416,In_405,In_141);
or U417 (N_417,In_174,In_305);
nand U418 (N_418,In_109,In_28);
and U419 (N_419,In_171,In_369);
xnor U420 (N_420,In_438,In_57);
nor U421 (N_421,In_240,In_457);
nand U422 (N_422,In_305,In_206);
nand U423 (N_423,In_96,In_111);
and U424 (N_424,In_478,In_266);
nand U425 (N_425,In_340,In_249);
and U426 (N_426,In_29,In_309);
nor U427 (N_427,In_409,In_315);
nand U428 (N_428,In_57,In_107);
xnor U429 (N_429,In_181,In_312);
nand U430 (N_430,In_99,In_168);
nor U431 (N_431,In_189,In_99);
nand U432 (N_432,In_68,In_308);
or U433 (N_433,In_449,In_49);
nor U434 (N_434,In_224,In_314);
or U435 (N_435,In_170,In_325);
nand U436 (N_436,In_303,In_386);
or U437 (N_437,In_431,In_148);
xnor U438 (N_438,In_482,In_364);
nand U439 (N_439,In_104,In_18);
nor U440 (N_440,In_119,In_497);
nand U441 (N_441,In_243,In_93);
and U442 (N_442,In_168,In_243);
and U443 (N_443,In_190,In_168);
or U444 (N_444,In_106,In_497);
xor U445 (N_445,In_29,In_371);
nand U446 (N_446,In_478,In_364);
nand U447 (N_447,In_408,In_256);
nand U448 (N_448,In_77,In_225);
or U449 (N_449,In_311,In_467);
nand U450 (N_450,In_385,In_78);
and U451 (N_451,In_448,In_227);
or U452 (N_452,In_32,In_380);
and U453 (N_453,In_108,In_311);
and U454 (N_454,In_105,In_120);
nand U455 (N_455,In_389,In_176);
nand U456 (N_456,In_16,In_344);
xor U457 (N_457,In_186,In_375);
or U458 (N_458,In_56,In_439);
and U459 (N_459,In_122,In_6);
or U460 (N_460,In_384,In_290);
and U461 (N_461,In_306,In_39);
nor U462 (N_462,In_319,In_404);
nand U463 (N_463,In_9,In_172);
nor U464 (N_464,In_132,In_458);
and U465 (N_465,In_33,In_340);
nand U466 (N_466,In_74,In_33);
nor U467 (N_467,In_489,In_27);
xor U468 (N_468,In_62,In_438);
nor U469 (N_469,In_223,In_53);
nand U470 (N_470,In_260,In_60);
or U471 (N_471,In_50,In_192);
nor U472 (N_472,In_491,In_396);
and U473 (N_473,In_410,In_338);
and U474 (N_474,In_112,In_400);
nor U475 (N_475,In_369,In_35);
or U476 (N_476,In_342,In_391);
nand U477 (N_477,In_393,In_301);
or U478 (N_478,In_216,In_255);
or U479 (N_479,In_126,In_393);
and U480 (N_480,In_88,In_470);
or U481 (N_481,In_200,In_0);
xnor U482 (N_482,In_25,In_33);
nor U483 (N_483,In_463,In_245);
or U484 (N_484,In_95,In_303);
nand U485 (N_485,In_111,In_484);
xnor U486 (N_486,In_321,In_291);
nand U487 (N_487,In_87,In_78);
nand U488 (N_488,In_260,In_121);
and U489 (N_489,In_353,In_18);
or U490 (N_490,In_161,In_483);
and U491 (N_491,In_92,In_455);
and U492 (N_492,In_51,In_401);
nand U493 (N_493,In_66,In_175);
nor U494 (N_494,In_120,In_1);
or U495 (N_495,In_494,In_33);
or U496 (N_496,In_403,In_282);
and U497 (N_497,In_258,In_342);
or U498 (N_498,In_45,In_298);
nor U499 (N_499,In_41,In_92);
nor U500 (N_500,In_43,In_35);
or U501 (N_501,In_49,In_480);
and U502 (N_502,In_295,In_91);
or U503 (N_503,In_199,In_98);
nor U504 (N_504,In_288,In_180);
or U505 (N_505,In_82,In_490);
or U506 (N_506,In_496,In_182);
nand U507 (N_507,In_164,In_45);
nor U508 (N_508,In_428,In_257);
nand U509 (N_509,In_428,In_407);
nor U510 (N_510,In_89,In_60);
nand U511 (N_511,In_475,In_134);
nand U512 (N_512,In_6,In_293);
and U513 (N_513,In_493,In_191);
xnor U514 (N_514,In_20,In_311);
or U515 (N_515,In_10,In_105);
and U516 (N_516,In_281,In_307);
and U517 (N_517,In_129,In_494);
nand U518 (N_518,In_308,In_359);
and U519 (N_519,In_429,In_89);
nand U520 (N_520,In_397,In_447);
nor U521 (N_521,In_363,In_379);
or U522 (N_522,In_22,In_361);
nor U523 (N_523,In_184,In_442);
nand U524 (N_524,In_367,In_125);
nor U525 (N_525,In_171,In_74);
xor U526 (N_526,In_239,In_241);
xor U527 (N_527,In_361,In_215);
xnor U528 (N_528,In_256,In_148);
and U529 (N_529,In_369,In_231);
nand U530 (N_530,In_355,In_322);
and U531 (N_531,In_77,In_12);
nor U532 (N_532,In_337,In_112);
or U533 (N_533,In_372,In_192);
and U534 (N_534,In_241,In_386);
nand U535 (N_535,In_284,In_456);
nand U536 (N_536,In_195,In_497);
nand U537 (N_537,In_436,In_301);
or U538 (N_538,In_60,In_24);
and U539 (N_539,In_261,In_405);
nand U540 (N_540,In_201,In_213);
or U541 (N_541,In_50,In_282);
or U542 (N_542,In_224,In_465);
and U543 (N_543,In_493,In_412);
or U544 (N_544,In_233,In_487);
nor U545 (N_545,In_443,In_474);
or U546 (N_546,In_161,In_387);
nor U547 (N_547,In_26,In_98);
and U548 (N_548,In_488,In_123);
nor U549 (N_549,In_387,In_124);
or U550 (N_550,In_430,In_197);
nand U551 (N_551,In_33,In_258);
nor U552 (N_552,In_286,In_276);
or U553 (N_553,In_340,In_260);
nand U554 (N_554,In_107,In_317);
xor U555 (N_555,In_112,In_83);
nor U556 (N_556,In_235,In_271);
or U557 (N_557,In_144,In_46);
nor U558 (N_558,In_362,In_200);
nor U559 (N_559,In_12,In_364);
nor U560 (N_560,In_157,In_321);
xor U561 (N_561,In_367,In_282);
nand U562 (N_562,In_464,In_302);
and U563 (N_563,In_368,In_92);
nor U564 (N_564,In_419,In_462);
nand U565 (N_565,In_11,In_1);
and U566 (N_566,In_77,In_96);
and U567 (N_567,In_418,In_28);
nor U568 (N_568,In_434,In_366);
and U569 (N_569,In_443,In_272);
or U570 (N_570,In_324,In_195);
nor U571 (N_571,In_158,In_315);
nand U572 (N_572,In_46,In_85);
nor U573 (N_573,In_195,In_320);
and U574 (N_574,In_138,In_5);
nor U575 (N_575,In_412,In_118);
xor U576 (N_576,In_36,In_252);
or U577 (N_577,In_210,In_113);
xor U578 (N_578,In_349,In_445);
nand U579 (N_579,In_14,In_378);
and U580 (N_580,In_419,In_56);
and U581 (N_581,In_348,In_400);
and U582 (N_582,In_478,In_27);
nor U583 (N_583,In_218,In_349);
nor U584 (N_584,In_433,In_361);
nand U585 (N_585,In_89,In_210);
and U586 (N_586,In_305,In_196);
nand U587 (N_587,In_255,In_48);
nor U588 (N_588,In_225,In_437);
nor U589 (N_589,In_211,In_317);
nor U590 (N_590,In_333,In_47);
and U591 (N_591,In_358,In_87);
and U592 (N_592,In_483,In_397);
nor U593 (N_593,In_150,In_193);
or U594 (N_594,In_363,In_317);
and U595 (N_595,In_148,In_149);
and U596 (N_596,In_70,In_203);
or U597 (N_597,In_462,In_31);
and U598 (N_598,In_149,In_117);
and U599 (N_599,In_428,In_210);
or U600 (N_600,In_391,In_90);
nor U601 (N_601,In_103,In_490);
or U602 (N_602,In_319,In_15);
and U603 (N_603,In_212,In_494);
and U604 (N_604,In_311,In_87);
or U605 (N_605,In_106,In_453);
nor U606 (N_606,In_249,In_238);
nor U607 (N_607,In_71,In_63);
nand U608 (N_608,In_374,In_128);
and U609 (N_609,In_459,In_396);
nor U610 (N_610,In_183,In_485);
nand U611 (N_611,In_353,In_157);
xnor U612 (N_612,In_235,In_463);
nand U613 (N_613,In_305,In_497);
nor U614 (N_614,In_240,In_172);
nor U615 (N_615,In_74,In_428);
and U616 (N_616,In_453,In_174);
nand U617 (N_617,In_442,In_2);
nor U618 (N_618,In_67,In_453);
nor U619 (N_619,In_256,In_129);
nand U620 (N_620,In_425,In_363);
and U621 (N_621,In_185,In_476);
nand U622 (N_622,In_43,In_131);
nor U623 (N_623,In_173,In_246);
and U624 (N_624,In_128,In_300);
or U625 (N_625,In_1,In_27);
or U626 (N_626,In_278,In_150);
nor U627 (N_627,In_173,In_462);
xor U628 (N_628,In_192,In_291);
nor U629 (N_629,In_413,In_202);
nand U630 (N_630,In_109,In_71);
nand U631 (N_631,In_436,In_470);
nand U632 (N_632,In_109,In_5);
nand U633 (N_633,In_21,In_303);
xnor U634 (N_634,In_118,In_411);
or U635 (N_635,In_102,In_307);
nor U636 (N_636,In_312,In_442);
xor U637 (N_637,In_47,In_66);
nor U638 (N_638,In_301,In_137);
or U639 (N_639,In_482,In_294);
xor U640 (N_640,In_169,In_192);
nor U641 (N_641,In_46,In_49);
or U642 (N_642,In_85,In_202);
and U643 (N_643,In_304,In_119);
nand U644 (N_644,In_447,In_257);
or U645 (N_645,In_113,In_388);
and U646 (N_646,In_257,In_133);
xor U647 (N_647,In_149,In_108);
and U648 (N_648,In_181,In_51);
nor U649 (N_649,In_33,In_235);
nor U650 (N_650,In_309,In_172);
nand U651 (N_651,In_127,In_235);
or U652 (N_652,In_143,In_11);
and U653 (N_653,In_45,In_397);
nor U654 (N_654,In_141,In_284);
or U655 (N_655,In_380,In_290);
or U656 (N_656,In_41,In_192);
or U657 (N_657,In_336,In_368);
nand U658 (N_658,In_298,In_495);
xnor U659 (N_659,In_314,In_372);
nand U660 (N_660,In_497,In_67);
or U661 (N_661,In_168,In_321);
or U662 (N_662,In_434,In_286);
nor U663 (N_663,In_484,In_355);
nor U664 (N_664,In_266,In_362);
or U665 (N_665,In_125,In_404);
or U666 (N_666,In_13,In_86);
nand U667 (N_667,In_167,In_291);
nor U668 (N_668,In_486,In_98);
xnor U669 (N_669,In_327,In_147);
nand U670 (N_670,In_432,In_275);
nand U671 (N_671,In_153,In_107);
and U672 (N_672,In_273,In_311);
nand U673 (N_673,In_399,In_480);
nand U674 (N_674,In_248,In_306);
xnor U675 (N_675,In_199,In_97);
and U676 (N_676,In_0,In_295);
or U677 (N_677,In_497,In_193);
nor U678 (N_678,In_401,In_400);
nor U679 (N_679,In_151,In_15);
nor U680 (N_680,In_25,In_485);
nand U681 (N_681,In_149,In_52);
or U682 (N_682,In_388,In_333);
nand U683 (N_683,In_56,In_92);
xnor U684 (N_684,In_228,In_404);
and U685 (N_685,In_15,In_330);
or U686 (N_686,In_338,In_22);
and U687 (N_687,In_219,In_93);
and U688 (N_688,In_113,In_104);
and U689 (N_689,In_296,In_95);
nor U690 (N_690,In_170,In_348);
nand U691 (N_691,In_365,In_126);
nand U692 (N_692,In_244,In_366);
nand U693 (N_693,In_121,In_153);
xnor U694 (N_694,In_208,In_26);
nand U695 (N_695,In_62,In_353);
and U696 (N_696,In_351,In_454);
or U697 (N_697,In_234,In_167);
nand U698 (N_698,In_405,In_15);
or U699 (N_699,In_359,In_34);
xor U700 (N_700,In_267,In_174);
or U701 (N_701,In_235,In_335);
nor U702 (N_702,In_413,In_203);
nand U703 (N_703,In_402,In_335);
xor U704 (N_704,In_376,In_120);
and U705 (N_705,In_490,In_324);
nand U706 (N_706,In_471,In_300);
nor U707 (N_707,In_12,In_221);
xor U708 (N_708,In_478,In_120);
nor U709 (N_709,In_155,In_221);
and U710 (N_710,In_99,In_171);
nand U711 (N_711,In_491,In_435);
and U712 (N_712,In_455,In_224);
nand U713 (N_713,In_60,In_177);
or U714 (N_714,In_128,In_122);
xor U715 (N_715,In_293,In_303);
and U716 (N_716,In_165,In_83);
or U717 (N_717,In_115,In_420);
nand U718 (N_718,In_249,In_73);
and U719 (N_719,In_381,In_469);
and U720 (N_720,In_241,In_86);
nor U721 (N_721,In_232,In_410);
and U722 (N_722,In_402,In_499);
and U723 (N_723,In_436,In_39);
or U724 (N_724,In_29,In_292);
nand U725 (N_725,In_451,In_411);
or U726 (N_726,In_187,In_303);
nor U727 (N_727,In_211,In_250);
nor U728 (N_728,In_68,In_460);
xor U729 (N_729,In_345,In_123);
and U730 (N_730,In_299,In_162);
and U731 (N_731,In_395,In_0);
nor U732 (N_732,In_492,In_375);
and U733 (N_733,In_148,In_416);
nand U734 (N_734,In_94,In_434);
nand U735 (N_735,In_321,In_251);
xor U736 (N_736,In_311,In_205);
nand U737 (N_737,In_196,In_365);
and U738 (N_738,In_231,In_343);
and U739 (N_739,In_338,In_370);
or U740 (N_740,In_154,In_289);
nand U741 (N_741,In_403,In_161);
and U742 (N_742,In_101,In_77);
nor U743 (N_743,In_481,In_226);
and U744 (N_744,In_217,In_287);
nand U745 (N_745,In_116,In_255);
or U746 (N_746,In_141,In_103);
or U747 (N_747,In_164,In_110);
and U748 (N_748,In_319,In_78);
nor U749 (N_749,In_425,In_127);
or U750 (N_750,In_182,In_352);
and U751 (N_751,In_171,In_373);
or U752 (N_752,In_426,In_288);
nor U753 (N_753,In_270,In_311);
xnor U754 (N_754,In_153,In_474);
and U755 (N_755,In_199,In_279);
nand U756 (N_756,In_139,In_313);
or U757 (N_757,In_282,In_400);
nor U758 (N_758,In_124,In_33);
or U759 (N_759,In_297,In_264);
and U760 (N_760,In_67,In_20);
and U761 (N_761,In_81,In_31);
and U762 (N_762,In_233,In_110);
or U763 (N_763,In_373,In_24);
or U764 (N_764,In_263,In_423);
xnor U765 (N_765,In_11,In_310);
or U766 (N_766,In_42,In_185);
or U767 (N_767,In_202,In_264);
or U768 (N_768,In_107,In_128);
nor U769 (N_769,In_379,In_193);
or U770 (N_770,In_244,In_408);
nand U771 (N_771,In_478,In_128);
or U772 (N_772,In_345,In_367);
nand U773 (N_773,In_19,In_422);
nand U774 (N_774,In_383,In_295);
nand U775 (N_775,In_498,In_137);
and U776 (N_776,In_136,In_207);
nand U777 (N_777,In_495,In_104);
nand U778 (N_778,In_342,In_425);
or U779 (N_779,In_15,In_216);
or U780 (N_780,In_457,In_165);
and U781 (N_781,In_318,In_335);
and U782 (N_782,In_455,In_260);
nor U783 (N_783,In_390,In_173);
or U784 (N_784,In_76,In_134);
or U785 (N_785,In_309,In_276);
xnor U786 (N_786,In_499,In_454);
nand U787 (N_787,In_391,In_398);
xor U788 (N_788,In_55,In_335);
and U789 (N_789,In_432,In_337);
and U790 (N_790,In_31,In_143);
nor U791 (N_791,In_391,In_176);
or U792 (N_792,In_168,In_173);
nand U793 (N_793,In_379,In_49);
nand U794 (N_794,In_228,In_128);
nand U795 (N_795,In_210,In_346);
nand U796 (N_796,In_287,In_326);
or U797 (N_797,In_125,In_63);
nand U798 (N_798,In_100,In_265);
and U799 (N_799,In_320,In_420);
and U800 (N_800,In_108,In_480);
and U801 (N_801,In_167,In_268);
nor U802 (N_802,In_237,In_477);
nor U803 (N_803,In_435,In_94);
nand U804 (N_804,In_226,In_29);
nand U805 (N_805,In_342,In_406);
or U806 (N_806,In_117,In_112);
or U807 (N_807,In_207,In_303);
and U808 (N_808,In_418,In_170);
and U809 (N_809,In_160,In_224);
or U810 (N_810,In_186,In_233);
nand U811 (N_811,In_250,In_168);
or U812 (N_812,In_378,In_398);
nor U813 (N_813,In_33,In_16);
or U814 (N_814,In_238,In_439);
nand U815 (N_815,In_2,In_417);
and U816 (N_816,In_118,In_341);
or U817 (N_817,In_192,In_297);
xor U818 (N_818,In_402,In_277);
nor U819 (N_819,In_192,In_465);
or U820 (N_820,In_470,In_407);
nor U821 (N_821,In_24,In_439);
nand U822 (N_822,In_332,In_114);
xnor U823 (N_823,In_296,In_337);
xor U824 (N_824,In_163,In_489);
xnor U825 (N_825,In_307,In_76);
or U826 (N_826,In_33,In_32);
and U827 (N_827,In_216,In_457);
nor U828 (N_828,In_47,In_127);
or U829 (N_829,In_259,In_208);
and U830 (N_830,In_246,In_6);
or U831 (N_831,In_379,In_300);
xnor U832 (N_832,In_261,In_387);
nor U833 (N_833,In_208,In_263);
nor U834 (N_834,In_108,In_374);
or U835 (N_835,In_393,In_297);
nand U836 (N_836,In_474,In_498);
nand U837 (N_837,In_291,In_193);
and U838 (N_838,In_421,In_227);
nand U839 (N_839,In_145,In_8);
xnor U840 (N_840,In_101,In_96);
nand U841 (N_841,In_309,In_165);
nand U842 (N_842,In_148,In_116);
nor U843 (N_843,In_262,In_314);
nor U844 (N_844,In_432,In_439);
nand U845 (N_845,In_200,In_85);
or U846 (N_846,In_476,In_73);
nand U847 (N_847,In_421,In_446);
and U848 (N_848,In_39,In_292);
or U849 (N_849,In_28,In_270);
xnor U850 (N_850,In_332,In_107);
nand U851 (N_851,In_317,In_187);
nand U852 (N_852,In_226,In_44);
nand U853 (N_853,In_216,In_408);
nor U854 (N_854,In_180,In_236);
and U855 (N_855,In_365,In_482);
or U856 (N_856,In_141,In_340);
and U857 (N_857,In_269,In_15);
and U858 (N_858,In_118,In_410);
xnor U859 (N_859,In_54,In_299);
nor U860 (N_860,In_161,In_221);
nand U861 (N_861,In_472,In_363);
or U862 (N_862,In_181,In_269);
or U863 (N_863,In_71,In_12);
nand U864 (N_864,In_271,In_39);
or U865 (N_865,In_382,In_110);
and U866 (N_866,In_195,In_149);
or U867 (N_867,In_182,In_317);
nand U868 (N_868,In_285,In_137);
and U869 (N_869,In_432,In_26);
nand U870 (N_870,In_315,In_222);
nand U871 (N_871,In_178,In_471);
or U872 (N_872,In_465,In_76);
xnor U873 (N_873,In_200,In_327);
nand U874 (N_874,In_238,In_455);
and U875 (N_875,In_279,In_179);
nor U876 (N_876,In_317,In_479);
nand U877 (N_877,In_247,In_389);
or U878 (N_878,In_466,In_134);
xnor U879 (N_879,In_110,In_192);
xor U880 (N_880,In_449,In_441);
nand U881 (N_881,In_369,In_114);
and U882 (N_882,In_319,In_399);
nand U883 (N_883,In_268,In_63);
nor U884 (N_884,In_311,In_340);
and U885 (N_885,In_154,In_113);
nand U886 (N_886,In_250,In_388);
and U887 (N_887,In_459,In_298);
or U888 (N_888,In_440,In_32);
or U889 (N_889,In_4,In_299);
and U890 (N_890,In_370,In_393);
nor U891 (N_891,In_180,In_139);
nand U892 (N_892,In_64,In_183);
nand U893 (N_893,In_270,In_307);
and U894 (N_894,In_434,In_193);
and U895 (N_895,In_484,In_99);
and U896 (N_896,In_74,In_350);
xor U897 (N_897,In_414,In_457);
and U898 (N_898,In_315,In_79);
nor U899 (N_899,In_25,In_161);
and U900 (N_900,In_262,In_413);
and U901 (N_901,In_318,In_184);
nand U902 (N_902,In_10,In_454);
and U903 (N_903,In_474,In_236);
and U904 (N_904,In_139,In_164);
nand U905 (N_905,In_63,In_351);
nor U906 (N_906,In_21,In_271);
xor U907 (N_907,In_254,In_366);
and U908 (N_908,In_114,In_165);
or U909 (N_909,In_246,In_43);
nand U910 (N_910,In_148,In_187);
and U911 (N_911,In_35,In_107);
or U912 (N_912,In_171,In_5);
or U913 (N_913,In_439,In_415);
nand U914 (N_914,In_404,In_202);
nand U915 (N_915,In_332,In_185);
nand U916 (N_916,In_237,In_228);
or U917 (N_917,In_448,In_117);
nor U918 (N_918,In_301,In_112);
or U919 (N_919,In_137,In_368);
xor U920 (N_920,In_220,In_401);
nor U921 (N_921,In_396,In_363);
and U922 (N_922,In_474,In_83);
or U923 (N_923,In_90,In_341);
nand U924 (N_924,In_487,In_325);
nand U925 (N_925,In_426,In_393);
or U926 (N_926,In_275,In_39);
nand U927 (N_927,In_270,In_320);
xnor U928 (N_928,In_80,In_19);
xnor U929 (N_929,In_321,In_105);
nand U930 (N_930,In_8,In_251);
nand U931 (N_931,In_62,In_264);
and U932 (N_932,In_451,In_176);
nor U933 (N_933,In_105,In_366);
xor U934 (N_934,In_387,In_347);
nand U935 (N_935,In_213,In_118);
nand U936 (N_936,In_58,In_83);
nor U937 (N_937,In_53,In_384);
or U938 (N_938,In_122,In_65);
or U939 (N_939,In_7,In_70);
nand U940 (N_940,In_428,In_470);
nand U941 (N_941,In_228,In_296);
nor U942 (N_942,In_458,In_377);
and U943 (N_943,In_32,In_316);
or U944 (N_944,In_236,In_499);
or U945 (N_945,In_123,In_24);
nand U946 (N_946,In_359,In_481);
and U947 (N_947,In_299,In_91);
or U948 (N_948,In_325,In_82);
nor U949 (N_949,In_237,In_167);
nor U950 (N_950,In_35,In_144);
and U951 (N_951,In_296,In_215);
or U952 (N_952,In_233,In_184);
xnor U953 (N_953,In_65,In_53);
nand U954 (N_954,In_145,In_160);
and U955 (N_955,In_91,In_383);
nand U956 (N_956,In_376,In_67);
or U957 (N_957,In_16,In_463);
xnor U958 (N_958,In_21,In_405);
nor U959 (N_959,In_100,In_10);
or U960 (N_960,In_227,In_152);
and U961 (N_961,In_173,In_8);
or U962 (N_962,In_140,In_312);
nand U963 (N_963,In_487,In_409);
nor U964 (N_964,In_226,In_403);
xnor U965 (N_965,In_9,In_428);
nor U966 (N_966,In_104,In_37);
and U967 (N_967,In_385,In_67);
nand U968 (N_968,In_245,In_371);
nand U969 (N_969,In_486,In_365);
nor U970 (N_970,In_436,In_337);
nor U971 (N_971,In_133,In_213);
nor U972 (N_972,In_201,In_152);
nand U973 (N_973,In_402,In_328);
and U974 (N_974,In_205,In_164);
and U975 (N_975,In_296,In_459);
or U976 (N_976,In_383,In_186);
nor U977 (N_977,In_28,In_427);
nand U978 (N_978,In_333,In_177);
nor U979 (N_979,In_302,In_198);
and U980 (N_980,In_52,In_93);
nand U981 (N_981,In_72,In_197);
or U982 (N_982,In_112,In_262);
nand U983 (N_983,In_206,In_360);
or U984 (N_984,In_455,In_291);
nor U985 (N_985,In_11,In_393);
or U986 (N_986,In_144,In_74);
nand U987 (N_987,In_177,In_362);
nor U988 (N_988,In_211,In_107);
and U989 (N_989,In_52,In_76);
nor U990 (N_990,In_139,In_468);
and U991 (N_991,In_394,In_490);
nor U992 (N_992,In_176,In_66);
nand U993 (N_993,In_376,In_272);
and U994 (N_994,In_288,In_73);
xor U995 (N_995,In_190,In_109);
or U996 (N_996,In_492,In_105);
nand U997 (N_997,In_334,In_335);
nor U998 (N_998,In_296,In_117);
or U999 (N_999,In_472,In_111);
and U1000 (N_1000,N_761,N_843);
or U1001 (N_1001,N_307,N_694);
nor U1002 (N_1002,N_447,N_911);
nor U1003 (N_1003,N_591,N_786);
xor U1004 (N_1004,N_808,N_268);
nor U1005 (N_1005,N_396,N_580);
nor U1006 (N_1006,N_673,N_466);
nand U1007 (N_1007,N_951,N_215);
nand U1008 (N_1008,N_169,N_946);
xor U1009 (N_1009,N_674,N_490);
nand U1010 (N_1010,N_770,N_563);
and U1011 (N_1011,N_882,N_343);
nor U1012 (N_1012,N_96,N_857);
nor U1013 (N_1013,N_572,N_149);
or U1014 (N_1014,N_944,N_986);
or U1015 (N_1015,N_354,N_245);
nor U1016 (N_1016,N_531,N_285);
nor U1017 (N_1017,N_616,N_665);
or U1018 (N_1018,N_769,N_739);
or U1019 (N_1019,N_908,N_655);
or U1020 (N_1020,N_461,N_899);
and U1021 (N_1021,N_732,N_237);
xnor U1022 (N_1022,N_416,N_874);
nor U1023 (N_1023,N_481,N_925);
or U1024 (N_1024,N_265,N_181);
nand U1025 (N_1025,N_984,N_450);
nor U1026 (N_1026,N_782,N_733);
and U1027 (N_1027,N_541,N_240);
xnor U1028 (N_1028,N_127,N_637);
or U1029 (N_1029,N_208,N_816);
nor U1030 (N_1030,N_428,N_949);
xor U1031 (N_1031,N_669,N_205);
and U1032 (N_1032,N_690,N_195);
nor U1033 (N_1033,N_876,N_627);
xor U1034 (N_1034,N_787,N_287);
or U1035 (N_1035,N_869,N_864);
or U1036 (N_1036,N_35,N_862);
nor U1037 (N_1037,N_401,N_160);
nand U1038 (N_1038,N_484,N_507);
nor U1039 (N_1039,N_46,N_192);
nor U1040 (N_1040,N_757,N_508);
or U1041 (N_1041,N_676,N_894);
nor U1042 (N_1042,N_523,N_742);
and U1043 (N_1043,N_480,N_686);
nand U1044 (N_1044,N_41,N_184);
nand U1045 (N_1045,N_996,N_498);
or U1046 (N_1046,N_547,N_55);
nor U1047 (N_1047,N_311,N_140);
or U1048 (N_1048,N_34,N_652);
or U1049 (N_1049,N_972,N_110);
nor U1050 (N_1050,N_200,N_985);
or U1051 (N_1051,N_934,N_749);
nand U1052 (N_1052,N_705,N_227);
or U1053 (N_1053,N_796,N_333);
or U1054 (N_1054,N_682,N_472);
nand U1055 (N_1055,N_483,N_358);
and U1056 (N_1056,N_385,N_706);
nand U1057 (N_1057,N_317,N_859);
and U1058 (N_1058,N_282,N_83);
and U1059 (N_1059,N_931,N_136);
nand U1060 (N_1060,N_535,N_218);
nor U1061 (N_1061,N_768,N_820);
and U1062 (N_1062,N_479,N_458);
xnor U1063 (N_1063,N_660,N_444);
nor U1064 (N_1064,N_856,N_722);
xnor U1065 (N_1065,N_922,N_106);
xor U1066 (N_1066,N_153,N_687);
and U1067 (N_1067,N_314,N_38);
nor U1068 (N_1068,N_391,N_395);
or U1069 (N_1069,N_14,N_131);
nand U1070 (N_1070,N_842,N_460);
nand U1071 (N_1071,N_981,N_210);
nand U1072 (N_1072,N_113,N_568);
or U1073 (N_1073,N_390,N_664);
and U1074 (N_1074,N_18,N_893);
or U1075 (N_1075,N_817,N_79);
or U1076 (N_1076,N_873,N_709);
nand U1077 (N_1077,N_906,N_696);
nand U1078 (N_1078,N_763,N_67);
and U1079 (N_1079,N_593,N_90);
or U1080 (N_1080,N_239,N_810);
and U1081 (N_1081,N_740,N_69);
nand U1082 (N_1082,N_948,N_501);
or U1083 (N_1083,N_302,N_585);
and U1084 (N_1084,N_289,N_767);
nor U1085 (N_1085,N_328,N_513);
nor U1086 (N_1086,N_361,N_849);
and U1087 (N_1087,N_952,N_646);
or U1088 (N_1088,N_117,N_21);
or U1089 (N_1089,N_191,N_525);
and U1090 (N_1090,N_725,N_273);
nand U1091 (N_1091,N_154,N_607);
or U1092 (N_1092,N_233,N_737);
or U1093 (N_1093,N_558,N_392);
nand U1094 (N_1094,N_97,N_403);
xor U1095 (N_1095,N_771,N_956);
or U1096 (N_1096,N_592,N_267);
and U1097 (N_1097,N_526,N_965);
nand U1098 (N_1098,N_425,N_429);
nand U1099 (N_1099,N_663,N_270);
and U1100 (N_1100,N_601,N_647);
or U1101 (N_1101,N_721,N_728);
and U1102 (N_1102,N_53,N_835);
and U1103 (N_1103,N_983,N_916);
xnor U1104 (N_1104,N_603,N_921);
xor U1105 (N_1105,N_649,N_362);
nand U1106 (N_1106,N_129,N_549);
and U1107 (N_1107,N_22,N_836);
and U1108 (N_1108,N_299,N_860);
and U1109 (N_1109,N_754,N_870);
or U1110 (N_1110,N_798,N_125);
nand U1111 (N_1111,N_834,N_953);
nand U1112 (N_1112,N_630,N_368);
or U1113 (N_1113,N_274,N_126);
xnor U1114 (N_1114,N_731,N_297);
nand U1115 (N_1115,N_756,N_567);
nor U1116 (N_1116,N_747,N_412);
nand U1117 (N_1117,N_793,N_847);
nor U1118 (N_1118,N_506,N_10);
or U1119 (N_1119,N_524,N_77);
nor U1120 (N_1120,N_625,N_180);
nand U1121 (N_1121,N_222,N_61);
or U1122 (N_1122,N_42,N_701);
nand U1123 (N_1123,N_24,N_130);
xor U1124 (N_1124,N_310,N_621);
and U1125 (N_1125,N_794,N_379);
nor U1126 (N_1126,N_552,N_642);
nand U1127 (N_1127,N_107,N_597);
nand U1128 (N_1128,N_219,N_84);
and U1129 (N_1129,N_813,N_528);
or U1130 (N_1130,N_296,N_471);
or U1131 (N_1131,N_809,N_364);
nand U1132 (N_1132,N_389,N_324);
nor U1133 (N_1133,N_777,N_305);
nand U1134 (N_1134,N_714,N_692);
or U1135 (N_1135,N_464,N_811);
or U1136 (N_1136,N_631,N_868);
nand U1137 (N_1137,N_662,N_653);
or U1138 (N_1138,N_897,N_402);
xor U1139 (N_1139,N_539,N_25);
or U1140 (N_1140,N_773,N_475);
and U1141 (N_1141,N_927,N_459);
and U1142 (N_1142,N_691,N_930);
xor U1143 (N_1143,N_774,N_75);
or U1144 (N_1144,N_954,N_881);
xnor U1145 (N_1145,N_968,N_420);
nor U1146 (N_1146,N_202,N_807);
or U1147 (N_1147,N_224,N_561);
and U1148 (N_1148,N_86,N_648);
or U1149 (N_1149,N_684,N_183);
nand U1150 (N_1150,N_998,N_293);
xor U1151 (N_1151,N_196,N_203);
xor U1152 (N_1152,N_765,N_212);
nor U1153 (N_1153,N_111,N_557);
or U1154 (N_1154,N_712,N_979);
nand U1155 (N_1155,N_907,N_91);
and U1156 (N_1156,N_244,N_342);
nand U1157 (N_1157,N_58,N_841);
nand U1158 (N_1158,N_966,N_468);
nand U1159 (N_1159,N_858,N_292);
nand U1160 (N_1160,N_964,N_485);
and U1161 (N_1161,N_16,N_905);
nand U1162 (N_1162,N_880,N_672);
or U1163 (N_1163,N_729,N_29);
or U1164 (N_1164,N_40,N_26);
and U1165 (N_1165,N_915,N_330);
and U1166 (N_1166,N_456,N_277);
nor U1167 (N_1167,N_409,N_230);
or U1168 (N_1168,N_666,N_904);
or U1169 (N_1169,N_453,N_31);
nor U1170 (N_1170,N_123,N_114);
nand U1171 (N_1171,N_321,N_940);
nand U1172 (N_1172,N_279,N_411);
nand U1173 (N_1173,N_863,N_800);
and U1174 (N_1174,N_942,N_433);
nor U1175 (N_1175,N_231,N_667);
and U1176 (N_1176,N_249,N_823);
or U1177 (N_1177,N_346,N_65);
xor U1178 (N_1178,N_118,N_382);
and U1179 (N_1179,N_848,N_896);
xor U1180 (N_1180,N_325,N_708);
xor U1181 (N_1181,N_137,N_251);
nor U1182 (N_1182,N_300,N_148);
nor U1183 (N_1183,N_989,N_442);
nand U1184 (N_1184,N_0,N_750);
and U1185 (N_1185,N_15,N_675);
xor U1186 (N_1186,N_753,N_586);
nor U1187 (N_1187,N_766,N_815);
and U1188 (N_1188,N_536,N_37);
and U1189 (N_1189,N_23,N_242);
xor U1190 (N_1190,N_758,N_936);
and U1191 (N_1191,N_308,N_133);
xor U1192 (N_1192,N_688,N_166);
and U1193 (N_1193,N_776,N_824);
or U1194 (N_1194,N_730,N_469);
nor U1195 (N_1195,N_397,N_867);
and U1196 (N_1196,N_805,N_959);
or U1197 (N_1197,N_295,N_910);
nor U1198 (N_1198,N_494,N_168);
or U1199 (N_1199,N_564,N_879);
and U1200 (N_1200,N_748,N_359);
nor U1201 (N_1201,N_509,N_194);
nor U1202 (N_1202,N_167,N_441);
nor U1203 (N_1203,N_598,N_71);
nor U1204 (N_1204,N_2,N_262);
or U1205 (N_1205,N_252,N_121);
nor U1206 (N_1206,N_845,N_398);
nor U1207 (N_1207,N_545,N_670);
nand U1208 (N_1208,N_155,N_829);
nor U1209 (N_1209,N_298,N_421);
and U1210 (N_1210,N_413,N_958);
and U1211 (N_1211,N_306,N_13);
nand U1212 (N_1212,N_573,N_241);
or U1213 (N_1213,N_8,N_290);
xnor U1214 (N_1214,N_799,N_538);
nand U1215 (N_1215,N_932,N_473);
nor U1216 (N_1216,N_978,N_57);
nor U1217 (N_1217,N_929,N_68);
or U1218 (N_1218,N_540,N_375);
or U1219 (N_1219,N_831,N_370);
nor U1220 (N_1220,N_211,N_717);
or U1221 (N_1221,N_724,N_284);
or U1222 (N_1222,N_641,N_253);
nor U1223 (N_1223,N_496,N_451);
or U1224 (N_1224,N_937,N_263);
nor U1225 (N_1225,N_974,N_178);
nand U1226 (N_1226,N_999,N_44);
nor U1227 (N_1227,N_527,N_920);
nor U1228 (N_1228,N_632,N_336);
nor U1229 (N_1229,N_566,N_759);
nor U1230 (N_1230,N_103,N_47);
nor U1231 (N_1231,N_264,N_246);
or U1232 (N_1232,N_720,N_119);
and U1233 (N_1233,N_519,N_833);
and U1234 (N_1234,N_120,N_376);
nor U1235 (N_1235,N_806,N_434);
and U1236 (N_1236,N_872,N_229);
and U1237 (N_1237,N_578,N_33);
xor U1238 (N_1238,N_973,N_762);
nand U1239 (N_1239,N_259,N_991);
nand U1240 (N_1240,N_344,N_455);
or U1241 (N_1241,N_515,N_656);
nor U1242 (N_1242,N_746,N_488);
or U1243 (N_1243,N_751,N_101);
xnor U1244 (N_1244,N_695,N_579);
nor U1245 (N_1245,N_380,N_723);
nand U1246 (N_1246,N_193,N_410);
xnor U1247 (N_1247,N_883,N_518);
or U1248 (N_1248,N_530,N_839);
and U1249 (N_1249,N_960,N_657);
nor U1250 (N_1250,N_182,N_316);
nor U1251 (N_1251,N_581,N_559);
nor U1252 (N_1252,N_514,N_755);
nand U1253 (N_1253,N_349,N_788);
nand U1254 (N_1254,N_112,N_924);
or U1255 (N_1255,N_726,N_877);
nor U1256 (N_1256,N_574,N_704);
nand U1257 (N_1257,N_304,N_280);
or U1258 (N_1258,N_606,N_78);
and U1259 (N_1259,N_64,N_997);
nand U1260 (N_1260,N_365,N_885);
or U1261 (N_1261,N_529,N_784);
or U1262 (N_1262,N_443,N_415);
xor U1263 (N_1263,N_257,N_889);
and U1264 (N_1264,N_512,N_914);
and U1265 (N_1265,N_94,N_571);
nand U1266 (N_1266,N_52,N_624);
nand U1267 (N_1267,N_59,N_6);
nor U1268 (N_1268,N_727,N_73);
or U1269 (N_1269,N_935,N_462);
nor U1270 (N_1270,N_609,N_143);
or U1271 (N_1271,N_644,N_837);
nor U1272 (N_1272,N_772,N_801);
or U1273 (N_1273,N_497,N_291);
and U1274 (N_1274,N_618,N_283);
or U1275 (N_1275,N_735,N_825);
and U1276 (N_1276,N_335,N_790);
nor U1277 (N_1277,N_478,N_795);
and U1278 (N_1278,N_66,N_711);
nand U1279 (N_1279,N_340,N_173);
or U1280 (N_1280,N_95,N_108);
nand U1281 (N_1281,N_892,N_629);
nor U1282 (N_1282,N_636,N_791);
and U1283 (N_1283,N_171,N_671);
nand U1284 (N_1284,N_532,N_188);
and U1285 (N_1285,N_158,N_923);
nor U1286 (N_1286,N_439,N_661);
nand U1287 (N_1287,N_286,N_312);
xnor U1288 (N_1288,N_353,N_634);
or U1289 (N_1289,N_596,N_901);
nand U1290 (N_1290,N_615,N_743);
nand U1291 (N_1291,N_332,N_778);
or U1292 (N_1292,N_957,N_165);
or U1293 (N_1293,N_427,N_247);
nand U1294 (N_1294,N_5,N_134);
or U1295 (N_1295,N_393,N_124);
nand U1296 (N_1296,N_738,N_424);
and U1297 (N_1297,N_174,N_620);
and U1298 (N_1298,N_463,N_432);
nand U1299 (N_1299,N_161,N_20);
xor U1300 (N_1300,N_363,N_792);
or U1301 (N_1301,N_994,N_221);
xor U1302 (N_1302,N_760,N_151);
nand U1303 (N_1303,N_577,N_635);
nand U1304 (N_1304,N_12,N_565);
and U1305 (N_1305,N_736,N_407);
nand U1306 (N_1306,N_617,N_614);
nor U1307 (N_1307,N_685,N_27);
nand U1308 (N_1308,N_371,N_39);
nor U1309 (N_1309,N_803,N_159);
nand U1310 (N_1310,N_697,N_802);
or U1311 (N_1311,N_832,N_553);
nand U1312 (N_1312,N_322,N_377);
or U1313 (N_1313,N_853,N_323);
nand U1314 (N_1314,N_476,N_900);
and U1315 (N_1315,N_105,N_628);
nor U1316 (N_1316,N_56,N_678);
nor U1317 (N_1317,N_139,N_214);
xnor U1318 (N_1318,N_967,N_320);
nor U1319 (N_1319,N_982,N_612);
and U1320 (N_1320,N_157,N_437);
nand U1321 (N_1321,N_309,N_318);
nor U1322 (N_1322,N_588,N_374);
and U1323 (N_1323,N_838,N_594);
or U1324 (N_1324,N_830,N_152);
nor U1325 (N_1325,N_1,N_85);
nor U1326 (N_1326,N_446,N_186);
or U1327 (N_1327,N_608,N_903);
nand U1328 (N_1328,N_457,N_797);
or U1329 (N_1329,N_569,N_339);
or U1330 (N_1330,N_223,N_185);
xor U1331 (N_1331,N_404,N_719);
or U1332 (N_1332,N_645,N_595);
or U1333 (N_1333,N_560,N_217);
and U1334 (N_1334,N_266,N_633);
nand U1335 (N_1335,N_367,N_199);
and U1336 (N_1336,N_659,N_871);
xnor U1337 (N_1337,N_775,N_570);
and U1338 (N_1338,N_502,N_236);
nor U1339 (N_1339,N_668,N_987);
xnor U1340 (N_1340,N_132,N_818);
and U1341 (N_1341,N_980,N_700);
nand U1342 (N_1342,N_116,N_543);
nor U1343 (N_1343,N_933,N_255);
nor U1344 (N_1344,N_477,N_74);
and U1345 (N_1345,N_431,N_970);
or U1346 (N_1346,N_804,N_715);
xnor U1347 (N_1347,N_550,N_950);
nand U1348 (N_1348,N_11,N_898);
and U1349 (N_1349,N_164,N_408);
nand U1350 (N_1350,N_517,N_76);
nor U1351 (N_1351,N_82,N_917);
nand U1352 (N_1352,N_172,N_941);
or U1353 (N_1353,N_610,N_963);
nand U1354 (N_1354,N_331,N_258);
nor U1355 (N_1355,N_969,N_313);
or U1356 (N_1356,N_104,N_521);
nand U1357 (N_1357,N_426,N_378);
or U1358 (N_1358,N_551,N_142);
xor U1359 (N_1359,N_487,N_147);
and U1360 (N_1360,N_63,N_689);
nand U1361 (N_1361,N_926,N_643);
and U1362 (N_1362,N_851,N_405);
and U1363 (N_1363,N_220,N_45);
nor U1364 (N_1364,N_288,N_844);
and U1365 (N_1365,N_341,N_28);
nor U1366 (N_1366,N_294,N_888);
or U1367 (N_1367,N_781,N_315);
or U1368 (N_1368,N_135,N_582);
or U1369 (N_1369,N_734,N_785);
or U1370 (N_1370,N_520,N_533);
nor U1371 (N_1371,N_840,N_373);
nor U1372 (N_1372,N_658,N_387);
nand U1373 (N_1373,N_122,N_913);
nand U1374 (N_1374,N_522,N_576);
nor U1375 (N_1375,N_326,N_886);
and U1376 (N_1376,N_890,N_698);
or U1377 (N_1377,N_962,N_400);
or U1378 (N_1378,N_206,N_875);
or U1379 (N_1379,N_861,N_360);
nor U1380 (N_1380,N_445,N_470);
or U1381 (N_1381,N_977,N_228);
nand U1382 (N_1382,N_542,N_355);
nor U1383 (N_1383,N_454,N_436);
or U1384 (N_1384,N_43,N_912);
nor U1385 (N_1385,N_943,N_235);
nor U1386 (N_1386,N_232,N_744);
nand U1387 (N_1387,N_613,N_546);
or U1388 (N_1388,N_993,N_537);
or U1389 (N_1389,N_419,N_72);
or U1390 (N_1390,N_81,N_971);
nor U1391 (N_1391,N_583,N_197);
or U1392 (N_1392,N_226,N_49);
nand U1393 (N_1393,N_482,N_812);
and U1394 (N_1394,N_144,N_699);
nand U1395 (N_1395,N_414,N_866);
nor U1396 (N_1396,N_878,N_681);
nand U1397 (N_1397,N_819,N_189);
and U1398 (N_1398,N_826,N_789);
nor U1399 (N_1399,N_179,N_955);
and U1400 (N_1400,N_677,N_256);
or U1401 (N_1401,N_62,N_128);
nor U1402 (N_1402,N_187,N_510);
and U1403 (N_1403,N_89,N_7);
nand U1404 (N_1404,N_887,N_99);
nand U1405 (N_1405,N_347,N_350);
nand U1406 (N_1406,N_975,N_156);
xnor U1407 (N_1407,N_209,N_599);
and U1408 (N_1408,N_170,N_327);
nand U1409 (N_1409,N_163,N_418);
xnor U1410 (N_1410,N_87,N_345);
and U1411 (N_1411,N_109,N_718);
nor U1412 (N_1412,N_357,N_177);
and U1413 (N_1413,N_17,N_175);
and U1414 (N_1414,N_384,N_319);
xnor U1415 (N_1415,N_752,N_115);
and U1416 (N_1416,N_50,N_474);
and U1417 (N_1417,N_261,N_48);
nor U1418 (N_1418,N_271,N_422);
nand U1419 (N_1419,N_976,N_430);
or U1420 (N_1420,N_276,N_141);
nand U1421 (N_1421,N_351,N_366);
or U1422 (N_1422,N_92,N_440);
or U1423 (N_1423,N_909,N_650);
and U1424 (N_1424,N_988,N_138);
xnor U1425 (N_1425,N_556,N_814);
and U1426 (N_1426,N_348,N_945);
nor U1427 (N_1427,N_654,N_369);
and U1428 (N_1428,N_865,N_895);
and U1429 (N_1429,N_503,N_716);
or U1430 (N_1430,N_250,N_990);
and U1431 (N_1431,N_448,N_939);
or U1432 (N_1432,N_902,N_70);
nand U1433 (N_1433,N_102,N_198);
nand U1434 (N_1434,N_640,N_201);
nand U1435 (N_1435,N_854,N_828);
or U1436 (N_1436,N_381,N_32);
or U1437 (N_1437,N_683,N_780);
nor U1438 (N_1438,N_891,N_590);
or U1439 (N_1439,N_467,N_275);
and U1440 (N_1440,N_822,N_622);
and U1441 (N_1441,N_19,N_741);
xor U1442 (N_1442,N_548,N_465);
nor U1443 (N_1443,N_176,N_534);
nand U1444 (N_1444,N_544,N_204);
and U1445 (N_1445,N_855,N_504);
xor U1446 (N_1446,N_54,N_500);
xor U1447 (N_1447,N_386,N_638);
nand U1448 (N_1448,N_51,N_555);
nor U1449 (N_1449,N_938,N_713);
and U1450 (N_1450,N_611,N_619);
or U1451 (N_1451,N_562,N_961);
or U1452 (N_1452,N_639,N_352);
or U1453 (N_1453,N_225,N_98);
and U1454 (N_1454,N_388,N_850);
nor U1455 (N_1455,N_575,N_919);
nand U1456 (N_1456,N_150,N_489);
or U1457 (N_1457,N_764,N_783);
nand U1458 (N_1458,N_213,N_254);
and U1459 (N_1459,N_435,N_329);
nor U1460 (N_1460,N_707,N_584);
and U1461 (N_1461,N_372,N_623);
or U1462 (N_1462,N_60,N_337);
nand U1463 (N_1463,N_383,N_3);
nand U1464 (N_1464,N_602,N_693);
and U1465 (N_1465,N_884,N_626);
or U1466 (N_1466,N_452,N_928);
nor U1467 (N_1467,N_100,N_449);
and U1468 (N_1468,N_260,N_93);
nand U1469 (N_1469,N_281,N_238);
nand U1470 (N_1470,N_234,N_486);
nor U1471 (N_1471,N_162,N_495);
or U1472 (N_1472,N_992,N_821);
nor U1473 (N_1473,N_146,N_846);
and U1474 (N_1474,N_827,N_947);
and U1475 (N_1475,N_417,N_600);
nor U1476 (N_1476,N_30,N_88);
nand U1477 (N_1477,N_438,N_703);
or U1478 (N_1478,N_356,N_492);
nor U1479 (N_1479,N_248,N_852);
or U1480 (N_1480,N_511,N_4);
nor U1481 (N_1481,N_589,N_190);
nand U1482 (N_1482,N_499,N_207);
xor U1483 (N_1483,N_301,N_36);
nor U1484 (N_1484,N_679,N_491);
nor U1485 (N_1485,N_9,N_710);
nand U1486 (N_1486,N_702,N_651);
or U1487 (N_1487,N_406,N_272);
and U1488 (N_1488,N_303,N_80);
or U1489 (N_1489,N_680,N_145);
nand U1490 (N_1490,N_216,N_605);
or U1491 (N_1491,N_278,N_243);
nand U1492 (N_1492,N_516,N_338);
nor U1493 (N_1493,N_918,N_587);
and U1494 (N_1494,N_493,N_399);
nor U1495 (N_1495,N_423,N_269);
nor U1496 (N_1496,N_505,N_745);
nand U1497 (N_1497,N_779,N_394);
nor U1498 (N_1498,N_995,N_554);
and U1499 (N_1499,N_604,N_334);
or U1500 (N_1500,N_33,N_175);
nor U1501 (N_1501,N_240,N_890);
nand U1502 (N_1502,N_137,N_401);
or U1503 (N_1503,N_957,N_487);
nor U1504 (N_1504,N_722,N_989);
nor U1505 (N_1505,N_456,N_691);
nor U1506 (N_1506,N_908,N_136);
and U1507 (N_1507,N_906,N_228);
xnor U1508 (N_1508,N_661,N_450);
xnor U1509 (N_1509,N_970,N_84);
nor U1510 (N_1510,N_222,N_612);
nand U1511 (N_1511,N_668,N_70);
xor U1512 (N_1512,N_474,N_903);
or U1513 (N_1513,N_84,N_942);
xnor U1514 (N_1514,N_23,N_950);
nand U1515 (N_1515,N_761,N_571);
nor U1516 (N_1516,N_552,N_988);
and U1517 (N_1517,N_650,N_445);
nand U1518 (N_1518,N_562,N_546);
nor U1519 (N_1519,N_989,N_980);
nand U1520 (N_1520,N_716,N_186);
and U1521 (N_1521,N_807,N_296);
nor U1522 (N_1522,N_957,N_988);
nand U1523 (N_1523,N_237,N_423);
and U1524 (N_1524,N_439,N_758);
or U1525 (N_1525,N_996,N_50);
xor U1526 (N_1526,N_848,N_504);
xnor U1527 (N_1527,N_336,N_770);
and U1528 (N_1528,N_847,N_77);
nor U1529 (N_1529,N_531,N_545);
nor U1530 (N_1530,N_366,N_336);
and U1531 (N_1531,N_416,N_98);
xor U1532 (N_1532,N_922,N_689);
xor U1533 (N_1533,N_550,N_330);
and U1534 (N_1534,N_361,N_193);
nor U1535 (N_1535,N_231,N_596);
nor U1536 (N_1536,N_796,N_52);
nor U1537 (N_1537,N_623,N_834);
nor U1538 (N_1538,N_954,N_114);
or U1539 (N_1539,N_618,N_950);
nor U1540 (N_1540,N_954,N_290);
xnor U1541 (N_1541,N_510,N_816);
or U1542 (N_1542,N_65,N_770);
or U1543 (N_1543,N_596,N_238);
nand U1544 (N_1544,N_907,N_256);
nor U1545 (N_1545,N_142,N_945);
or U1546 (N_1546,N_572,N_469);
nand U1547 (N_1547,N_146,N_214);
and U1548 (N_1548,N_693,N_697);
or U1549 (N_1549,N_222,N_561);
nor U1550 (N_1550,N_301,N_163);
nor U1551 (N_1551,N_353,N_780);
nand U1552 (N_1552,N_52,N_871);
and U1553 (N_1553,N_996,N_383);
and U1554 (N_1554,N_720,N_607);
nand U1555 (N_1555,N_106,N_508);
nor U1556 (N_1556,N_23,N_715);
and U1557 (N_1557,N_808,N_338);
and U1558 (N_1558,N_788,N_397);
nor U1559 (N_1559,N_186,N_838);
or U1560 (N_1560,N_515,N_870);
and U1561 (N_1561,N_366,N_836);
nor U1562 (N_1562,N_130,N_112);
nand U1563 (N_1563,N_80,N_951);
or U1564 (N_1564,N_564,N_263);
nor U1565 (N_1565,N_707,N_867);
xor U1566 (N_1566,N_998,N_645);
and U1567 (N_1567,N_626,N_791);
or U1568 (N_1568,N_943,N_858);
nor U1569 (N_1569,N_226,N_253);
xor U1570 (N_1570,N_875,N_266);
and U1571 (N_1571,N_17,N_672);
or U1572 (N_1572,N_169,N_595);
nor U1573 (N_1573,N_134,N_633);
or U1574 (N_1574,N_394,N_575);
nand U1575 (N_1575,N_334,N_459);
nand U1576 (N_1576,N_460,N_701);
nand U1577 (N_1577,N_123,N_661);
or U1578 (N_1578,N_535,N_786);
and U1579 (N_1579,N_248,N_996);
or U1580 (N_1580,N_807,N_597);
nand U1581 (N_1581,N_199,N_490);
xnor U1582 (N_1582,N_641,N_985);
nor U1583 (N_1583,N_331,N_617);
and U1584 (N_1584,N_487,N_306);
nor U1585 (N_1585,N_513,N_564);
nand U1586 (N_1586,N_598,N_891);
nand U1587 (N_1587,N_733,N_199);
and U1588 (N_1588,N_104,N_149);
or U1589 (N_1589,N_4,N_589);
xnor U1590 (N_1590,N_291,N_821);
nand U1591 (N_1591,N_677,N_316);
nand U1592 (N_1592,N_901,N_679);
nand U1593 (N_1593,N_992,N_381);
xor U1594 (N_1594,N_404,N_303);
and U1595 (N_1595,N_855,N_702);
or U1596 (N_1596,N_906,N_643);
nor U1597 (N_1597,N_571,N_974);
nand U1598 (N_1598,N_9,N_584);
and U1599 (N_1599,N_420,N_888);
nor U1600 (N_1600,N_285,N_304);
and U1601 (N_1601,N_227,N_931);
or U1602 (N_1602,N_44,N_400);
or U1603 (N_1603,N_881,N_594);
nand U1604 (N_1604,N_648,N_131);
or U1605 (N_1605,N_749,N_944);
nand U1606 (N_1606,N_968,N_221);
nor U1607 (N_1607,N_45,N_180);
nand U1608 (N_1608,N_395,N_406);
nand U1609 (N_1609,N_222,N_229);
nand U1610 (N_1610,N_651,N_82);
nor U1611 (N_1611,N_770,N_417);
nand U1612 (N_1612,N_866,N_166);
xor U1613 (N_1613,N_506,N_931);
and U1614 (N_1614,N_343,N_862);
xor U1615 (N_1615,N_892,N_835);
nand U1616 (N_1616,N_353,N_704);
and U1617 (N_1617,N_471,N_941);
and U1618 (N_1618,N_800,N_64);
nor U1619 (N_1619,N_971,N_515);
or U1620 (N_1620,N_259,N_151);
nand U1621 (N_1621,N_637,N_627);
or U1622 (N_1622,N_575,N_607);
nor U1623 (N_1623,N_216,N_844);
nor U1624 (N_1624,N_725,N_179);
or U1625 (N_1625,N_734,N_520);
xor U1626 (N_1626,N_258,N_388);
xnor U1627 (N_1627,N_805,N_414);
nor U1628 (N_1628,N_88,N_302);
nand U1629 (N_1629,N_897,N_958);
nor U1630 (N_1630,N_417,N_783);
and U1631 (N_1631,N_785,N_35);
or U1632 (N_1632,N_199,N_286);
nand U1633 (N_1633,N_835,N_198);
nand U1634 (N_1634,N_679,N_854);
or U1635 (N_1635,N_824,N_386);
and U1636 (N_1636,N_554,N_548);
nand U1637 (N_1637,N_993,N_896);
xor U1638 (N_1638,N_192,N_881);
nor U1639 (N_1639,N_655,N_555);
nor U1640 (N_1640,N_316,N_148);
nor U1641 (N_1641,N_587,N_969);
xor U1642 (N_1642,N_161,N_248);
nor U1643 (N_1643,N_463,N_229);
and U1644 (N_1644,N_650,N_90);
or U1645 (N_1645,N_856,N_151);
and U1646 (N_1646,N_333,N_850);
or U1647 (N_1647,N_474,N_836);
or U1648 (N_1648,N_49,N_277);
or U1649 (N_1649,N_905,N_801);
nor U1650 (N_1650,N_25,N_687);
nor U1651 (N_1651,N_392,N_373);
nor U1652 (N_1652,N_530,N_714);
nor U1653 (N_1653,N_780,N_68);
and U1654 (N_1654,N_789,N_815);
and U1655 (N_1655,N_278,N_838);
xor U1656 (N_1656,N_923,N_62);
nor U1657 (N_1657,N_38,N_565);
nor U1658 (N_1658,N_674,N_719);
or U1659 (N_1659,N_381,N_67);
and U1660 (N_1660,N_295,N_959);
xor U1661 (N_1661,N_638,N_565);
nor U1662 (N_1662,N_163,N_219);
and U1663 (N_1663,N_886,N_57);
xor U1664 (N_1664,N_691,N_375);
nor U1665 (N_1665,N_779,N_527);
xnor U1666 (N_1666,N_423,N_70);
nor U1667 (N_1667,N_391,N_238);
or U1668 (N_1668,N_436,N_346);
nand U1669 (N_1669,N_20,N_295);
and U1670 (N_1670,N_62,N_785);
nand U1671 (N_1671,N_347,N_297);
xor U1672 (N_1672,N_759,N_552);
nand U1673 (N_1673,N_66,N_321);
or U1674 (N_1674,N_6,N_216);
or U1675 (N_1675,N_854,N_372);
xnor U1676 (N_1676,N_129,N_925);
nor U1677 (N_1677,N_223,N_633);
and U1678 (N_1678,N_55,N_986);
and U1679 (N_1679,N_286,N_186);
and U1680 (N_1680,N_10,N_478);
and U1681 (N_1681,N_513,N_847);
and U1682 (N_1682,N_456,N_270);
and U1683 (N_1683,N_834,N_140);
and U1684 (N_1684,N_767,N_875);
or U1685 (N_1685,N_205,N_850);
or U1686 (N_1686,N_128,N_351);
and U1687 (N_1687,N_215,N_757);
or U1688 (N_1688,N_141,N_948);
or U1689 (N_1689,N_791,N_409);
nor U1690 (N_1690,N_302,N_578);
nor U1691 (N_1691,N_600,N_497);
or U1692 (N_1692,N_188,N_774);
nor U1693 (N_1693,N_646,N_106);
nor U1694 (N_1694,N_33,N_98);
and U1695 (N_1695,N_836,N_111);
or U1696 (N_1696,N_64,N_916);
nand U1697 (N_1697,N_7,N_910);
nor U1698 (N_1698,N_297,N_650);
or U1699 (N_1699,N_574,N_597);
nand U1700 (N_1700,N_424,N_867);
and U1701 (N_1701,N_168,N_487);
or U1702 (N_1702,N_310,N_263);
xnor U1703 (N_1703,N_953,N_145);
or U1704 (N_1704,N_879,N_39);
or U1705 (N_1705,N_78,N_507);
nor U1706 (N_1706,N_914,N_192);
or U1707 (N_1707,N_885,N_105);
nand U1708 (N_1708,N_964,N_451);
xnor U1709 (N_1709,N_258,N_779);
or U1710 (N_1710,N_880,N_7);
nand U1711 (N_1711,N_533,N_400);
or U1712 (N_1712,N_498,N_812);
and U1713 (N_1713,N_281,N_783);
or U1714 (N_1714,N_933,N_590);
nand U1715 (N_1715,N_860,N_102);
nor U1716 (N_1716,N_770,N_574);
and U1717 (N_1717,N_806,N_67);
and U1718 (N_1718,N_681,N_668);
and U1719 (N_1719,N_40,N_534);
nand U1720 (N_1720,N_146,N_762);
or U1721 (N_1721,N_649,N_786);
and U1722 (N_1722,N_628,N_99);
and U1723 (N_1723,N_147,N_669);
and U1724 (N_1724,N_231,N_465);
nor U1725 (N_1725,N_12,N_132);
nor U1726 (N_1726,N_348,N_13);
or U1727 (N_1727,N_459,N_617);
nor U1728 (N_1728,N_175,N_68);
nor U1729 (N_1729,N_28,N_460);
nor U1730 (N_1730,N_457,N_261);
and U1731 (N_1731,N_478,N_422);
xor U1732 (N_1732,N_805,N_913);
nor U1733 (N_1733,N_228,N_808);
nand U1734 (N_1734,N_211,N_436);
and U1735 (N_1735,N_856,N_64);
xnor U1736 (N_1736,N_238,N_272);
nor U1737 (N_1737,N_518,N_109);
nand U1738 (N_1738,N_545,N_53);
nor U1739 (N_1739,N_114,N_262);
xnor U1740 (N_1740,N_367,N_181);
nor U1741 (N_1741,N_441,N_316);
nor U1742 (N_1742,N_555,N_715);
nand U1743 (N_1743,N_22,N_615);
xnor U1744 (N_1744,N_629,N_585);
xor U1745 (N_1745,N_371,N_598);
and U1746 (N_1746,N_374,N_162);
nor U1747 (N_1747,N_166,N_889);
or U1748 (N_1748,N_898,N_327);
nor U1749 (N_1749,N_673,N_841);
and U1750 (N_1750,N_694,N_416);
nor U1751 (N_1751,N_48,N_436);
xnor U1752 (N_1752,N_658,N_8);
or U1753 (N_1753,N_853,N_768);
and U1754 (N_1754,N_787,N_384);
or U1755 (N_1755,N_398,N_486);
xnor U1756 (N_1756,N_201,N_86);
nor U1757 (N_1757,N_940,N_837);
nor U1758 (N_1758,N_244,N_42);
nor U1759 (N_1759,N_111,N_760);
nand U1760 (N_1760,N_701,N_947);
and U1761 (N_1761,N_228,N_918);
or U1762 (N_1762,N_829,N_770);
nor U1763 (N_1763,N_363,N_961);
nand U1764 (N_1764,N_936,N_398);
and U1765 (N_1765,N_206,N_158);
and U1766 (N_1766,N_543,N_962);
xor U1767 (N_1767,N_53,N_773);
xor U1768 (N_1768,N_527,N_361);
nand U1769 (N_1769,N_927,N_776);
nor U1770 (N_1770,N_142,N_538);
or U1771 (N_1771,N_809,N_501);
nand U1772 (N_1772,N_143,N_41);
nand U1773 (N_1773,N_146,N_481);
nand U1774 (N_1774,N_920,N_217);
or U1775 (N_1775,N_466,N_766);
nand U1776 (N_1776,N_299,N_476);
and U1777 (N_1777,N_120,N_806);
nand U1778 (N_1778,N_141,N_855);
xnor U1779 (N_1779,N_941,N_38);
or U1780 (N_1780,N_498,N_676);
nand U1781 (N_1781,N_906,N_588);
xnor U1782 (N_1782,N_683,N_701);
nand U1783 (N_1783,N_794,N_24);
or U1784 (N_1784,N_726,N_847);
and U1785 (N_1785,N_914,N_221);
nand U1786 (N_1786,N_460,N_440);
or U1787 (N_1787,N_542,N_866);
nor U1788 (N_1788,N_137,N_997);
and U1789 (N_1789,N_369,N_71);
nor U1790 (N_1790,N_298,N_916);
and U1791 (N_1791,N_677,N_878);
or U1792 (N_1792,N_594,N_181);
and U1793 (N_1793,N_699,N_360);
nor U1794 (N_1794,N_354,N_366);
or U1795 (N_1795,N_16,N_224);
or U1796 (N_1796,N_945,N_527);
nor U1797 (N_1797,N_217,N_36);
or U1798 (N_1798,N_604,N_883);
nand U1799 (N_1799,N_6,N_345);
or U1800 (N_1800,N_174,N_298);
and U1801 (N_1801,N_644,N_686);
or U1802 (N_1802,N_555,N_299);
nor U1803 (N_1803,N_492,N_454);
xor U1804 (N_1804,N_807,N_627);
and U1805 (N_1805,N_884,N_83);
xor U1806 (N_1806,N_653,N_249);
and U1807 (N_1807,N_877,N_403);
nor U1808 (N_1808,N_796,N_523);
or U1809 (N_1809,N_155,N_895);
or U1810 (N_1810,N_695,N_341);
nand U1811 (N_1811,N_88,N_180);
nor U1812 (N_1812,N_343,N_48);
xor U1813 (N_1813,N_321,N_56);
nor U1814 (N_1814,N_910,N_114);
or U1815 (N_1815,N_621,N_423);
and U1816 (N_1816,N_595,N_818);
xnor U1817 (N_1817,N_974,N_119);
and U1818 (N_1818,N_265,N_114);
nor U1819 (N_1819,N_316,N_63);
nand U1820 (N_1820,N_455,N_380);
and U1821 (N_1821,N_166,N_767);
and U1822 (N_1822,N_409,N_498);
nor U1823 (N_1823,N_751,N_23);
or U1824 (N_1824,N_332,N_339);
nand U1825 (N_1825,N_57,N_435);
and U1826 (N_1826,N_269,N_496);
or U1827 (N_1827,N_652,N_647);
nand U1828 (N_1828,N_938,N_372);
or U1829 (N_1829,N_279,N_886);
or U1830 (N_1830,N_293,N_218);
or U1831 (N_1831,N_540,N_458);
or U1832 (N_1832,N_119,N_810);
or U1833 (N_1833,N_600,N_626);
and U1834 (N_1834,N_507,N_601);
or U1835 (N_1835,N_655,N_152);
nand U1836 (N_1836,N_875,N_481);
or U1837 (N_1837,N_28,N_681);
or U1838 (N_1838,N_256,N_527);
nand U1839 (N_1839,N_814,N_674);
xor U1840 (N_1840,N_990,N_692);
nand U1841 (N_1841,N_853,N_137);
or U1842 (N_1842,N_560,N_162);
xnor U1843 (N_1843,N_70,N_592);
and U1844 (N_1844,N_608,N_69);
and U1845 (N_1845,N_384,N_267);
and U1846 (N_1846,N_351,N_35);
and U1847 (N_1847,N_384,N_1);
or U1848 (N_1848,N_944,N_861);
nor U1849 (N_1849,N_478,N_959);
or U1850 (N_1850,N_444,N_170);
or U1851 (N_1851,N_219,N_808);
or U1852 (N_1852,N_64,N_439);
nor U1853 (N_1853,N_821,N_549);
nand U1854 (N_1854,N_381,N_851);
nor U1855 (N_1855,N_361,N_186);
xnor U1856 (N_1856,N_628,N_298);
nand U1857 (N_1857,N_878,N_672);
or U1858 (N_1858,N_682,N_436);
nand U1859 (N_1859,N_968,N_902);
or U1860 (N_1860,N_907,N_576);
xor U1861 (N_1861,N_14,N_52);
xnor U1862 (N_1862,N_374,N_947);
nand U1863 (N_1863,N_76,N_886);
or U1864 (N_1864,N_471,N_195);
nand U1865 (N_1865,N_593,N_332);
nor U1866 (N_1866,N_849,N_98);
nor U1867 (N_1867,N_11,N_785);
or U1868 (N_1868,N_670,N_480);
nor U1869 (N_1869,N_961,N_970);
xor U1870 (N_1870,N_510,N_16);
nand U1871 (N_1871,N_176,N_604);
and U1872 (N_1872,N_378,N_986);
or U1873 (N_1873,N_182,N_946);
or U1874 (N_1874,N_632,N_217);
xor U1875 (N_1875,N_654,N_238);
nand U1876 (N_1876,N_584,N_588);
and U1877 (N_1877,N_125,N_566);
nand U1878 (N_1878,N_855,N_727);
nor U1879 (N_1879,N_680,N_739);
nor U1880 (N_1880,N_854,N_395);
xor U1881 (N_1881,N_980,N_898);
xnor U1882 (N_1882,N_408,N_520);
and U1883 (N_1883,N_370,N_459);
nor U1884 (N_1884,N_408,N_586);
nand U1885 (N_1885,N_757,N_117);
or U1886 (N_1886,N_715,N_850);
or U1887 (N_1887,N_517,N_396);
nor U1888 (N_1888,N_360,N_192);
and U1889 (N_1889,N_205,N_619);
nor U1890 (N_1890,N_817,N_29);
nor U1891 (N_1891,N_92,N_115);
nor U1892 (N_1892,N_608,N_843);
nor U1893 (N_1893,N_919,N_316);
nor U1894 (N_1894,N_527,N_30);
nand U1895 (N_1895,N_595,N_492);
nand U1896 (N_1896,N_375,N_84);
xor U1897 (N_1897,N_761,N_126);
xor U1898 (N_1898,N_833,N_82);
nand U1899 (N_1899,N_660,N_79);
and U1900 (N_1900,N_248,N_592);
nor U1901 (N_1901,N_703,N_802);
nand U1902 (N_1902,N_288,N_394);
or U1903 (N_1903,N_891,N_867);
or U1904 (N_1904,N_625,N_391);
xor U1905 (N_1905,N_529,N_294);
and U1906 (N_1906,N_820,N_991);
or U1907 (N_1907,N_541,N_966);
nor U1908 (N_1908,N_754,N_48);
nor U1909 (N_1909,N_887,N_468);
and U1910 (N_1910,N_156,N_795);
nand U1911 (N_1911,N_545,N_522);
and U1912 (N_1912,N_656,N_240);
xnor U1913 (N_1913,N_530,N_558);
nand U1914 (N_1914,N_823,N_572);
and U1915 (N_1915,N_757,N_307);
and U1916 (N_1916,N_626,N_176);
nor U1917 (N_1917,N_305,N_10);
nor U1918 (N_1918,N_822,N_248);
or U1919 (N_1919,N_346,N_384);
or U1920 (N_1920,N_715,N_535);
and U1921 (N_1921,N_878,N_462);
xor U1922 (N_1922,N_947,N_972);
and U1923 (N_1923,N_250,N_450);
nand U1924 (N_1924,N_861,N_835);
nor U1925 (N_1925,N_726,N_793);
nor U1926 (N_1926,N_612,N_359);
nor U1927 (N_1927,N_209,N_714);
nor U1928 (N_1928,N_460,N_754);
or U1929 (N_1929,N_411,N_741);
xnor U1930 (N_1930,N_162,N_935);
nand U1931 (N_1931,N_370,N_148);
nor U1932 (N_1932,N_249,N_64);
nor U1933 (N_1933,N_7,N_296);
nor U1934 (N_1934,N_752,N_640);
or U1935 (N_1935,N_63,N_846);
nand U1936 (N_1936,N_905,N_528);
nand U1937 (N_1937,N_378,N_616);
nor U1938 (N_1938,N_148,N_374);
nor U1939 (N_1939,N_426,N_526);
or U1940 (N_1940,N_234,N_326);
xor U1941 (N_1941,N_264,N_468);
nand U1942 (N_1942,N_795,N_712);
xor U1943 (N_1943,N_851,N_926);
or U1944 (N_1944,N_651,N_10);
nor U1945 (N_1945,N_318,N_757);
nand U1946 (N_1946,N_3,N_47);
nor U1947 (N_1947,N_850,N_500);
nand U1948 (N_1948,N_705,N_530);
nand U1949 (N_1949,N_314,N_441);
and U1950 (N_1950,N_582,N_208);
xor U1951 (N_1951,N_954,N_884);
or U1952 (N_1952,N_310,N_307);
and U1953 (N_1953,N_110,N_407);
nand U1954 (N_1954,N_560,N_721);
nor U1955 (N_1955,N_758,N_935);
nor U1956 (N_1956,N_122,N_915);
or U1957 (N_1957,N_575,N_159);
nand U1958 (N_1958,N_285,N_163);
nand U1959 (N_1959,N_769,N_218);
and U1960 (N_1960,N_106,N_607);
or U1961 (N_1961,N_291,N_958);
and U1962 (N_1962,N_397,N_315);
nor U1963 (N_1963,N_632,N_7);
and U1964 (N_1964,N_99,N_805);
or U1965 (N_1965,N_344,N_551);
xnor U1966 (N_1966,N_354,N_385);
nor U1967 (N_1967,N_926,N_407);
nand U1968 (N_1968,N_211,N_577);
and U1969 (N_1969,N_566,N_589);
and U1970 (N_1970,N_521,N_649);
and U1971 (N_1971,N_561,N_828);
and U1972 (N_1972,N_423,N_788);
nand U1973 (N_1973,N_762,N_654);
nor U1974 (N_1974,N_857,N_929);
and U1975 (N_1975,N_67,N_962);
and U1976 (N_1976,N_315,N_171);
nor U1977 (N_1977,N_628,N_138);
xnor U1978 (N_1978,N_861,N_100);
nand U1979 (N_1979,N_941,N_210);
or U1980 (N_1980,N_507,N_320);
nor U1981 (N_1981,N_328,N_872);
nand U1982 (N_1982,N_270,N_273);
or U1983 (N_1983,N_35,N_358);
or U1984 (N_1984,N_285,N_985);
nor U1985 (N_1985,N_386,N_534);
nand U1986 (N_1986,N_936,N_261);
and U1987 (N_1987,N_200,N_793);
xor U1988 (N_1988,N_374,N_655);
nor U1989 (N_1989,N_956,N_752);
nor U1990 (N_1990,N_98,N_375);
nand U1991 (N_1991,N_130,N_502);
and U1992 (N_1992,N_841,N_696);
or U1993 (N_1993,N_992,N_835);
or U1994 (N_1994,N_90,N_413);
nand U1995 (N_1995,N_90,N_403);
or U1996 (N_1996,N_223,N_802);
nor U1997 (N_1997,N_728,N_85);
or U1998 (N_1998,N_814,N_368);
nor U1999 (N_1999,N_465,N_773);
nor U2000 (N_2000,N_1225,N_1533);
or U2001 (N_2001,N_1781,N_1964);
nand U2002 (N_2002,N_1978,N_1896);
xnor U2003 (N_2003,N_1329,N_1232);
and U2004 (N_2004,N_1555,N_1854);
xor U2005 (N_2005,N_1079,N_1181);
or U2006 (N_2006,N_1989,N_1217);
and U2007 (N_2007,N_1594,N_1447);
or U2008 (N_2008,N_1012,N_1548);
nand U2009 (N_2009,N_1497,N_1113);
nor U2010 (N_2010,N_1114,N_1644);
nand U2011 (N_2011,N_1492,N_1299);
or U2012 (N_2012,N_1008,N_1064);
nor U2013 (N_2013,N_1277,N_1146);
nand U2014 (N_2014,N_1154,N_1233);
and U2015 (N_2015,N_1442,N_1776);
nand U2016 (N_2016,N_1968,N_1386);
and U2017 (N_2017,N_1619,N_1509);
nand U2018 (N_2018,N_1482,N_1946);
or U2019 (N_2019,N_1957,N_1748);
nor U2020 (N_2020,N_1549,N_1613);
and U2021 (N_2021,N_1705,N_1280);
nor U2022 (N_2022,N_1566,N_1629);
and U2023 (N_2023,N_1024,N_1481);
xor U2024 (N_2024,N_1410,N_1027);
nand U2025 (N_2025,N_1556,N_1580);
nor U2026 (N_2026,N_1675,N_1536);
and U2027 (N_2027,N_1044,N_1059);
xnor U2028 (N_2028,N_1137,N_1955);
xor U2029 (N_2029,N_1042,N_1342);
or U2030 (N_2030,N_1473,N_1278);
and U2031 (N_2031,N_1956,N_1170);
nor U2032 (N_2032,N_1128,N_1071);
nand U2033 (N_2033,N_1805,N_1456);
nand U2034 (N_2034,N_1332,N_1680);
nand U2035 (N_2035,N_1035,N_1863);
or U2036 (N_2036,N_1296,N_1301);
or U2037 (N_2037,N_1838,N_1763);
nand U2038 (N_2038,N_1298,N_1377);
nand U2039 (N_2039,N_1685,N_1450);
nand U2040 (N_2040,N_1275,N_1972);
nor U2041 (N_2041,N_1733,N_1801);
and U2042 (N_2042,N_1292,N_1785);
nand U2043 (N_2043,N_1303,N_1740);
nand U2044 (N_2044,N_1798,N_1971);
and U2045 (N_2045,N_1373,N_1922);
and U2046 (N_2046,N_1226,N_1392);
and U2047 (N_2047,N_1938,N_1975);
nand U2048 (N_2048,N_1411,N_1300);
or U2049 (N_2049,N_1631,N_1932);
or U2050 (N_2050,N_1845,N_1165);
and U2051 (N_2051,N_1322,N_1852);
nand U2052 (N_2052,N_1016,N_1717);
xnor U2053 (N_2053,N_1351,N_1078);
nor U2054 (N_2054,N_1976,N_1129);
nor U2055 (N_2055,N_1356,N_1090);
or U2056 (N_2056,N_1849,N_1985);
xnor U2057 (N_2057,N_1446,N_1229);
or U2058 (N_2058,N_1219,N_1311);
or U2059 (N_2059,N_1507,N_1230);
nand U2060 (N_2060,N_1454,N_1074);
xor U2061 (N_2061,N_1856,N_1187);
and U2062 (N_2062,N_1252,N_1179);
or U2063 (N_2063,N_1043,N_1244);
and U2064 (N_2064,N_1799,N_1169);
nand U2065 (N_2065,N_1716,N_1937);
or U2066 (N_2066,N_1660,N_1818);
xor U2067 (N_2067,N_1242,N_1766);
nor U2068 (N_2068,N_1816,N_1337);
and U2069 (N_2069,N_1315,N_1485);
nor U2070 (N_2070,N_1729,N_1056);
and U2071 (N_2071,N_1634,N_1222);
nor U2072 (N_2072,N_1495,N_1089);
nor U2073 (N_2073,N_1098,N_1115);
xor U2074 (N_2074,N_1671,N_1757);
and U2075 (N_2075,N_1006,N_1822);
or U2076 (N_2076,N_1531,N_1681);
and U2077 (N_2077,N_1665,N_1568);
nor U2078 (N_2078,N_1095,N_1684);
nor U2079 (N_2079,N_1397,N_1084);
nand U2080 (N_2080,N_1258,N_1504);
and U2081 (N_2081,N_1574,N_1324);
nand U2082 (N_2082,N_1737,N_1775);
nor U2083 (N_2083,N_1100,N_1867);
or U2084 (N_2084,N_1520,N_1344);
nand U2085 (N_2085,N_1573,N_1182);
or U2086 (N_2086,N_1515,N_1360);
or U2087 (N_2087,N_1037,N_1579);
or U2088 (N_2088,N_1449,N_1167);
nand U2089 (N_2089,N_1657,N_1065);
and U2090 (N_2090,N_1532,N_1758);
and U2091 (N_2091,N_1802,N_1599);
nand U2092 (N_2092,N_1439,N_1490);
or U2093 (N_2093,N_1527,N_1227);
nand U2094 (N_2094,N_1718,N_1508);
or U2095 (N_2095,N_1910,N_1357);
nor U2096 (N_2096,N_1340,N_1279);
or U2097 (N_2097,N_1807,N_1476);
or U2098 (N_2098,N_1792,N_1944);
nor U2099 (N_2099,N_1372,N_1993);
xnor U2100 (N_2100,N_1068,N_1239);
nand U2101 (N_2101,N_1370,N_1109);
or U2102 (N_2102,N_1518,N_1567);
nand U2103 (N_2103,N_1274,N_1502);
nor U2104 (N_2104,N_1418,N_1614);
nor U2105 (N_2105,N_1917,N_1948);
nand U2106 (N_2106,N_1713,N_1941);
or U2107 (N_2107,N_1840,N_1711);
and U2108 (N_2108,N_1820,N_1092);
and U2109 (N_2109,N_1047,N_1029);
and U2110 (N_2110,N_1281,N_1431);
nor U2111 (N_2111,N_1590,N_1814);
nor U2112 (N_2112,N_1891,N_1694);
and U2113 (N_2113,N_1604,N_1404);
nor U2114 (N_2114,N_1622,N_1212);
and U2115 (N_2115,N_1345,N_1709);
and U2116 (N_2116,N_1554,N_1769);
and U2117 (N_2117,N_1843,N_1487);
nand U2118 (N_2118,N_1734,N_1139);
nor U2119 (N_2119,N_1609,N_1125);
or U2120 (N_2120,N_1969,N_1815);
or U2121 (N_2121,N_1529,N_1148);
or U2122 (N_2122,N_1381,N_1672);
and U2123 (N_2123,N_1894,N_1829);
or U2124 (N_2124,N_1736,N_1326);
and U2125 (N_2125,N_1004,N_1984);
nor U2126 (N_2126,N_1382,N_1460);
and U2127 (N_2127,N_1997,N_1073);
or U2128 (N_2128,N_1297,N_1739);
nor U2129 (N_2129,N_1517,N_1288);
nor U2130 (N_2130,N_1379,N_1451);
or U2131 (N_2131,N_1367,N_1659);
or U2132 (N_2132,N_1996,N_1582);
and U2133 (N_2133,N_1666,N_1184);
and U2134 (N_2134,N_1328,N_1869);
xnor U2135 (N_2135,N_1704,N_1905);
nand U2136 (N_2136,N_1986,N_1846);
nand U2137 (N_2137,N_1995,N_1848);
xnor U2138 (N_2138,N_1510,N_1223);
or U2139 (N_2139,N_1821,N_1803);
and U2140 (N_2140,N_1019,N_1506);
and U2141 (N_2141,N_1907,N_1817);
or U2142 (N_2142,N_1319,N_1791);
nor U2143 (N_2143,N_1427,N_1144);
nor U2144 (N_2144,N_1724,N_1082);
nor U2145 (N_2145,N_1403,N_1908);
or U2146 (N_2146,N_1116,N_1876);
or U2147 (N_2147,N_1358,N_1428);
and U2148 (N_2148,N_1276,N_1147);
and U2149 (N_2149,N_1257,N_1687);
nor U2150 (N_2150,N_1149,N_1827);
nor U2151 (N_2151,N_1467,N_1088);
nand U2152 (N_2152,N_1835,N_1118);
nand U2153 (N_2153,N_1131,N_1871);
nor U2154 (N_2154,N_1172,N_1690);
or U2155 (N_2155,N_1134,N_1009);
or U2156 (N_2156,N_1909,N_1030);
nand U2157 (N_2157,N_1330,N_1857);
nor U2158 (N_2158,N_1415,N_1263);
or U2159 (N_2159,N_1828,N_1437);
nand U2160 (N_2160,N_1346,N_1879);
nor U2161 (N_2161,N_1648,N_1316);
nand U2162 (N_2162,N_1645,N_1156);
and U2163 (N_2163,N_1112,N_1207);
or U2164 (N_2164,N_1958,N_1707);
or U2165 (N_2165,N_1695,N_1094);
nor U2166 (N_2166,N_1168,N_1773);
xnor U2167 (N_2167,N_1587,N_1458);
or U2168 (N_2168,N_1284,N_1669);
and U2169 (N_2169,N_1562,N_1140);
nand U2170 (N_2170,N_1954,N_1878);
and U2171 (N_2171,N_1860,N_1236);
nor U2172 (N_2172,N_1152,N_1347);
or U2173 (N_2173,N_1783,N_1979);
or U2174 (N_2174,N_1870,N_1466);
nand U2175 (N_2175,N_1173,N_1676);
nor U2176 (N_2176,N_1935,N_1294);
and U2177 (N_2177,N_1363,N_1689);
and U2178 (N_2178,N_1738,N_1438);
nor U2179 (N_2179,N_1753,N_1399);
and U2180 (N_2180,N_1433,N_1457);
nor U2181 (N_2181,N_1183,N_1304);
or U2182 (N_2182,N_1265,N_1010);
and U2183 (N_2183,N_1243,N_1699);
nand U2184 (N_2184,N_1559,N_1111);
xor U2185 (N_2185,N_1143,N_1673);
or U2186 (N_2186,N_1563,N_1962);
or U2187 (N_2187,N_1352,N_1591);
nor U2188 (N_2188,N_1534,N_1110);
nand U2189 (N_2189,N_1824,N_1444);
or U2190 (N_2190,N_1528,N_1105);
nand U2191 (N_2191,N_1949,N_1474);
or U2192 (N_2192,N_1331,N_1176);
or U2193 (N_2193,N_1916,N_1234);
nor U2194 (N_2194,N_1538,N_1691);
or U2195 (N_2195,N_1639,N_1371);
or U2196 (N_2196,N_1180,N_1395);
or U2197 (N_2197,N_1677,N_1161);
nor U2198 (N_2198,N_1866,N_1637);
and U2199 (N_2199,N_1786,N_1884);
or U2200 (N_2200,N_1470,N_1120);
nor U2201 (N_2201,N_1570,N_1195);
nand U2202 (N_2202,N_1099,N_1076);
or U2203 (N_2203,N_1790,N_1742);
nand U2204 (N_2204,N_1145,N_1751);
nand U2205 (N_2205,N_1026,N_1141);
nand U2206 (N_2206,N_1961,N_1063);
nor U2207 (N_2207,N_1777,N_1543);
nand U2208 (N_2208,N_1939,N_1286);
nand U2209 (N_2209,N_1545,N_1999);
nand U2210 (N_2210,N_1066,N_1264);
or U2211 (N_2211,N_1069,N_1809);
nand U2212 (N_2212,N_1633,N_1539);
or U2213 (N_2213,N_1755,N_1812);
nor U2214 (N_2214,N_1260,N_1889);
and U2215 (N_2215,N_1551,N_1833);
or U2216 (N_2216,N_1374,N_1654);
nor U2217 (N_2217,N_1421,N_1934);
or U2218 (N_2218,N_1423,N_1540);
and U2219 (N_2219,N_1463,N_1583);
and U2220 (N_2220,N_1133,N_1417);
nand U2221 (N_2221,N_1192,N_1953);
nor U2222 (N_2222,N_1213,N_1875);
nand U2223 (N_2223,N_1384,N_1643);
or U2224 (N_2224,N_1607,N_1560);
or U2225 (N_2225,N_1202,N_1664);
or U2226 (N_2226,N_1117,N_1919);
nand U2227 (N_2227,N_1537,N_1214);
and U2228 (N_2228,N_1253,N_1618);
and U2229 (N_2229,N_1892,N_1434);
or U2230 (N_2230,N_1692,N_1250);
and U2231 (N_2231,N_1220,N_1308);
or U2232 (N_2232,N_1475,N_1398);
and U2233 (N_2233,N_1904,N_1965);
nor U2234 (N_2234,N_1756,N_1620);
and U2235 (N_2235,N_1526,N_1422);
nand U2236 (N_2236,N_1174,N_1661);
nor U2237 (N_2237,N_1931,N_1942);
and U2238 (N_2238,N_1132,N_1096);
or U2239 (N_2239,N_1282,N_1290);
and U2240 (N_2240,N_1477,N_1067);
or U2241 (N_2241,N_1462,N_1858);
nor U2242 (N_2242,N_1647,N_1310);
nand U2243 (N_2243,N_1578,N_1032);
nor U2244 (N_2244,N_1868,N_1940);
and U2245 (N_2245,N_1393,N_1834);
or U2246 (N_2246,N_1569,N_1261);
xor U2247 (N_2247,N_1760,N_1901);
nor U2248 (N_2248,N_1649,N_1636);
or U2249 (N_2249,N_1072,N_1899);
or U2250 (N_2250,N_1697,N_1658);
and U2251 (N_2251,N_1336,N_1036);
nand U2252 (N_2252,N_1679,N_1499);
or U2253 (N_2253,N_1101,N_1542);
and U2254 (N_2254,N_1627,N_1761);
and U2255 (N_2255,N_1511,N_1977);
and U2256 (N_2256,N_1991,N_1708);
or U2257 (N_2257,N_1200,N_1855);
or U2258 (N_2258,N_1898,N_1126);
and U2259 (N_2259,N_1391,N_1205);
nand U2260 (N_2260,N_1780,N_1959);
nor U2261 (N_2261,N_1831,N_1254);
xor U2262 (N_2262,N_1194,N_1541);
or U2263 (N_2263,N_1459,N_1103);
or U2264 (N_2264,N_1893,N_1522);
nor U2265 (N_2265,N_1887,N_1124);
and U2266 (N_2266,N_1231,N_1602);
nand U2267 (N_2267,N_1060,N_1847);
xnor U2268 (N_2268,N_1033,N_1926);
nor U2269 (N_2269,N_1859,N_1000);
nand U2270 (N_2270,N_1535,N_1603);
and U2271 (N_2271,N_1521,N_1389);
nand U2272 (N_2272,N_1686,N_1023);
nand U2273 (N_2273,N_1193,N_1334);
or U2274 (N_2274,N_1662,N_1874);
and U2275 (N_2275,N_1663,N_1218);
nor U2276 (N_2276,N_1455,N_1880);
nor U2277 (N_2277,N_1429,N_1960);
nor U2278 (N_2278,N_1104,N_1045);
or U2279 (N_2279,N_1199,N_1617);
and U2280 (N_2280,N_1696,N_1771);
nor U2281 (N_2281,N_1266,N_1469);
nand U2282 (N_2282,N_1754,N_1974);
and U2283 (N_2283,N_1653,N_1851);
nor U2284 (N_2284,N_1318,N_1872);
or U2285 (N_2285,N_1178,N_1610);
nor U2286 (N_2286,N_1918,N_1712);
nand U2287 (N_2287,N_1714,N_1080);
nand U2288 (N_2288,N_1632,N_1572);
or U2289 (N_2289,N_1430,N_1700);
xor U2290 (N_2290,N_1952,N_1682);
and U2291 (N_2291,N_1106,N_1701);
or U2292 (N_2292,N_1362,N_1906);
xnor U2293 (N_2293,N_1123,N_1920);
nand U2294 (N_2294,N_1841,N_1598);
nor U2295 (N_2295,N_1380,N_1861);
nor U2296 (N_2296,N_1107,N_1557);
nor U2297 (N_2297,N_1493,N_1408);
and U2298 (N_2298,N_1121,N_1216);
and U2299 (N_2299,N_1921,N_1013);
and U2300 (N_2300,N_1268,N_1038);
nand U2301 (N_2301,N_1383,N_1836);
nor U2302 (N_2302,N_1628,N_1837);
nand U2303 (N_2303,N_1048,N_1640);
nand U2304 (N_2304,N_1083,N_1503);
nand U2305 (N_2305,N_1001,N_1782);
nand U2306 (N_2306,N_1787,N_1626);
and U2307 (N_2307,N_1524,N_1097);
nor U2308 (N_2308,N_1577,N_1093);
nor U2309 (N_2309,N_1523,N_1445);
nor U2310 (N_2310,N_1638,N_1588);
and U2311 (N_2311,N_1895,N_1414);
xor U2312 (N_2312,N_1723,N_1987);
xnor U2313 (N_2313,N_1491,N_1890);
nor U2314 (N_2314,N_1811,N_1865);
or U2315 (N_2315,N_1175,N_1850);
nor U2316 (N_2316,N_1720,N_1102);
nand U2317 (N_2317,N_1902,N_1994);
or U2318 (N_2318,N_1122,N_1269);
or U2319 (N_2319,N_1656,N_1262);
and U2320 (N_2320,N_1164,N_1930);
or U2321 (N_2321,N_1668,N_1519);
nor U2322 (N_2322,N_1784,N_1018);
xnor U2323 (N_2323,N_1287,N_1353);
and U2324 (N_2324,N_1550,N_1436);
nand U2325 (N_2325,N_1435,N_1224);
nand U2326 (N_2326,N_1589,N_1070);
nand U2327 (N_2327,N_1015,N_1153);
nand U2328 (N_2328,N_1270,N_1407);
or U2329 (N_2329,N_1320,N_1945);
nand U2330 (N_2330,N_1611,N_1947);
or U2331 (N_2331,N_1388,N_1593);
xnor U2332 (N_2332,N_1259,N_1888);
nor U2333 (N_2333,N_1484,N_1251);
nor U2334 (N_2334,N_1249,N_1196);
and U2335 (N_2335,N_1272,N_1981);
and U2336 (N_2336,N_1553,N_1630);
nand U2337 (N_2337,N_1592,N_1789);
nand U2338 (N_2338,N_1206,N_1349);
or U2339 (N_2339,N_1793,N_1237);
nor U2340 (N_2340,N_1702,N_1291);
nand U2341 (N_2341,N_1341,N_1642);
and U2342 (N_2342,N_1443,N_1565);
or U2343 (N_2343,N_1943,N_1394);
and U2344 (N_2344,N_1483,N_1983);
and U2345 (N_2345,N_1882,N_1797);
and U2346 (N_2346,N_1440,N_1478);
or U2347 (N_2347,N_1054,N_1744);
or U2348 (N_2348,N_1051,N_1151);
or U2349 (N_2349,N_1335,N_1615);
xor U2350 (N_2350,N_1077,N_1188);
nand U2351 (N_2351,N_1448,N_1359);
xnor U2352 (N_2352,N_1601,N_1075);
and U2353 (N_2353,N_1750,N_1584);
and U2354 (N_2354,N_1703,N_1215);
nor U2355 (N_2355,N_1652,N_1385);
or U2356 (N_2356,N_1914,N_1544);
nand U2357 (N_2357,N_1881,N_1108);
and U2358 (N_2358,N_1325,N_1135);
or U2359 (N_2359,N_1973,N_1516);
and U2360 (N_2360,N_1496,N_1832);
and U2361 (N_2361,N_1885,N_1488);
or U2362 (N_2362,N_1119,N_1929);
and U2363 (N_2363,N_1606,N_1586);
nand U2364 (N_2364,N_1350,N_1501);
nor U2365 (N_2365,N_1525,N_1749);
and U2366 (N_2366,N_1728,N_1623);
or U2367 (N_2367,N_1877,N_1616);
nor U2368 (N_2368,N_1479,N_1364);
nand U2369 (N_2369,N_1788,N_1683);
and U2370 (N_2370,N_1376,N_1897);
xor U2371 (N_2371,N_1765,N_1810);
or U2372 (N_2372,N_1752,N_1409);
nor U2373 (N_2373,N_1267,N_1052);
and U2374 (N_2374,N_1348,N_1767);
xnor U2375 (N_2375,N_1864,N_1412);
nand U2376 (N_2376,N_1950,N_1369);
xnor U2377 (N_2377,N_1091,N_1285);
nor U2378 (N_2378,N_1406,N_1354);
nand U2379 (N_2379,N_1513,N_1162);
nand U2380 (N_2380,N_1245,N_1317);
and U2381 (N_2381,N_1823,N_1800);
and U2382 (N_2382,N_1323,N_1839);
or U2383 (N_2383,N_1034,N_1053);
xnor U2384 (N_2384,N_1339,N_1039);
nor U2385 (N_2385,N_1400,N_1585);
and U2386 (N_2386,N_1710,N_1171);
and U2387 (N_2387,N_1365,N_1913);
or U2388 (N_2388,N_1951,N_1651);
and U2389 (N_2389,N_1333,N_1600);
and U2390 (N_2390,N_1413,N_1925);
nand U2391 (N_2391,N_1461,N_1197);
nor U2392 (N_2392,N_1612,N_1057);
and U2393 (N_2393,N_1608,N_1204);
or U2394 (N_2394,N_1210,N_1726);
nand U2395 (N_2395,N_1127,N_1240);
nand U2396 (N_2396,N_1228,N_1361);
and U2397 (N_2397,N_1923,N_1970);
nand U2398 (N_2398,N_1201,N_1667);
or U2399 (N_2399,N_1514,N_1830);
nor U2400 (N_2400,N_1424,N_1903);
nor U2401 (N_2401,N_1031,N_1988);
or U2402 (N_2402,N_1159,N_1605);
nor U2403 (N_2403,N_1779,N_1924);
nor U2404 (N_2404,N_1419,N_1058);
nor U2405 (N_2405,N_1747,N_1998);
and U2406 (N_2406,N_1853,N_1595);
or U2407 (N_2407,N_1558,N_1722);
or U2408 (N_2408,N_1883,N_1990);
xnor U2409 (N_2409,N_1017,N_1862);
or U2410 (N_2410,N_1933,N_1808);
nor U2411 (N_2411,N_1007,N_1186);
nor U2412 (N_2412,N_1211,N_1338);
nor U2413 (N_2413,N_1795,N_1900);
nor U2414 (N_2414,N_1238,N_1177);
xnor U2415 (N_2415,N_1575,N_1471);
nand U2416 (N_2416,N_1635,N_1844);
nand U2417 (N_2417,N_1625,N_1731);
or U2418 (N_2418,N_1256,N_1725);
nand U2419 (N_2419,N_1040,N_1313);
and U2420 (N_2420,N_1321,N_1759);
and U2421 (N_2421,N_1688,N_1087);
nand U2422 (N_2422,N_1003,N_1806);
or U2423 (N_2423,N_1650,N_1198);
nor U2424 (N_2424,N_1561,N_1886);
and U2425 (N_2425,N_1813,N_1396);
nand U2426 (N_2426,N_1378,N_1086);
nand U2427 (N_2427,N_1764,N_1770);
xnor U2428 (N_2428,N_1293,N_1375);
nor U2429 (N_2429,N_1826,N_1745);
or U2430 (N_2430,N_1307,N_1735);
nor U2431 (N_2431,N_1646,N_1721);
xor U2432 (N_2432,N_1505,N_1746);
nor U2433 (N_2433,N_1130,N_1772);
and U2434 (N_2434,N_1005,N_1028);
xor U2435 (N_2435,N_1425,N_1796);
nand U2436 (N_2436,N_1390,N_1730);
or U2437 (N_2437,N_1670,N_1401);
or U2438 (N_2438,N_1283,N_1498);
xnor U2439 (N_2439,N_1221,N_1842);
and U2440 (N_2440,N_1085,N_1982);
nor U2441 (N_2441,N_1530,N_1050);
and U2442 (N_2442,N_1355,N_1157);
nor U2443 (N_2443,N_1912,N_1967);
or U2444 (N_2444,N_1190,N_1472);
or U2445 (N_2445,N_1387,N_1046);
nand U2446 (N_2446,N_1873,N_1774);
and U2447 (N_2447,N_1166,N_1727);
nor U2448 (N_2448,N_1295,N_1185);
or U2449 (N_2449,N_1247,N_1289);
xor U2450 (N_2450,N_1208,N_1235);
or U2451 (N_2451,N_1189,N_1255);
or U2452 (N_2452,N_1138,N_1564);
nor U2453 (N_2453,N_1025,N_1191);
nor U2454 (N_2454,N_1494,N_1416);
xor U2455 (N_2455,N_1055,N_1719);
and U2456 (N_2456,N_1405,N_1486);
nor U2457 (N_2457,N_1241,N_1426);
or U2458 (N_2458,N_1762,N_1020);
or U2459 (N_2459,N_1306,N_1480);
nor U2460 (N_2460,N_1049,N_1155);
and U2461 (N_2461,N_1366,N_1273);
nor U2462 (N_2462,N_1819,N_1576);
nand U2463 (N_2463,N_1512,N_1963);
xor U2464 (N_2464,N_1022,N_1547);
and U2465 (N_2465,N_1966,N_1209);
xnor U2466 (N_2466,N_1041,N_1248);
and U2467 (N_2467,N_1011,N_1021);
or U2468 (N_2468,N_1402,N_1160);
xnor U2469 (N_2469,N_1597,N_1621);
and U2470 (N_2470,N_1992,N_1150);
nor U2471 (N_2471,N_1203,N_1698);
xor U2472 (N_2472,N_1641,N_1980);
nor U2473 (N_2473,N_1136,N_1743);
and U2474 (N_2474,N_1302,N_1465);
xor U2475 (N_2475,N_1768,N_1732);
nor U2476 (N_2476,N_1778,N_1596);
nor U2477 (N_2477,N_1014,N_1706);
nand U2478 (N_2478,N_1581,N_1928);
or U2479 (N_2479,N_1062,N_1343);
nor U2480 (N_2480,N_1489,N_1142);
and U2481 (N_2481,N_1081,N_1678);
or U2482 (N_2482,N_1552,N_1002);
nand U2483 (N_2483,N_1794,N_1804);
and U2484 (N_2484,N_1693,N_1314);
and U2485 (N_2485,N_1655,N_1741);
nand U2486 (N_2486,N_1453,N_1911);
nor U2487 (N_2487,N_1441,N_1927);
xnor U2488 (N_2488,N_1246,N_1464);
nor U2489 (N_2489,N_1500,N_1825);
and U2490 (N_2490,N_1624,N_1674);
nor U2491 (N_2491,N_1915,N_1432);
nor U2492 (N_2492,N_1061,N_1312);
or U2493 (N_2493,N_1468,N_1305);
nor U2494 (N_2494,N_1368,N_1936);
and U2495 (N_2495,N_1571,N_1158);
and U2496 (N_2496,N_1452,N_1715);
nor U2497 (N_2497,N_1420,N_1309);
xnor U2498 (N_2498,N_1271,N_1163);
and U2499 (N_2499,N_1546,N_1327);
or U2500 (N_2500,N_1542,N_1339);
nor U2501 (N_2501,N_1496,N_1912);
nor U2502 (N_2502,N_1359,N_1881);
or U2503 (N_2503,N_1620,N_1021);
and U2504 (N_2504,N_1396,N_1368);
nand U2505 (N_2505,N_1950,N_1647);
or U2506 (N_2506,N_1904,N_1917);
and U2507 (N_2507,N_1290,N_1034);
nor U2508 (N_2508,N_1633,N_1993);
xor U2509 (N_2509,N_1459,N_1415);
nor U2510 (N_2510,N_1863,N_1286);
nor U2511 (N_2511,N_1777,N_1027);
or U2512 (N_2512,N_1979,N_1923);
nand U2513 (N_2513,N_1473,N_1993);
nand U2514 (N_2514,N_1113,N_1940);
nand U2515 (N_2515,N_1798,N_1932);
and U2516 (N_2516,N_1981,N_1991);
and U2517 (N_2517,N_1376,N_1371);
nand U2518 (N_2518,N_1921,N_1100);
xor U2519 (N_2519,N_1970,N_1230);
nor U2520 (N_2520,N_1981,N_1613);
nand U2521 (N_2521,N_1618,N_1572);
and U2522 (N_2522,N_1195,N_1861);
or U2523 (N_2523,N_1896,N_1654);
or U2524 (N_2524,N_1611,N_1240);
nor U2525 (N_2525,N_1323,N_1473);
and U2526 (N_2526,N_1267,N_1526);
or U2527 (N_2527,N_1351,N_1772);
or U2528 (N_2528,N_1668,N_1780);
or U2529 (N_2529,N_1024,N_1673);
nor U2530 (N_2530,N_1900,N_1698);
nand U2531 (N_2531,N_1546,N_1804);
and U2532 (N_2532,N_1330,N_1299);
and U2533 (N_2533,N_1220,N_1339);
and U2534 (N_2534,N_1132,N_1965);
nand U2535 (N_2535,N_1836,N_1160);
and U2536 (N_2536,N_1910,N_1675);
or U2537 (N_2537,N_1605,N_1756);
nand U2538 (N_2538,N_1572,N_1359);
and U2539 (N_2539,N_1282,N_1222);
nor U2540 (N_2540,N_1249,N_1687);
nor U2541 (N_2541,N_1161,N_1329);
or U2542 (N_2542,N_1223,N_1687);
nor U2543 (N_2543,N_1175,N_1226);
nand U2544 (N_2544,N_1123,N_1462);
nand U2545 (N_2545,N_1550,N_1117);
or U2546 (N_2546,N_1420,N_1108);
nand U2547 (N_2547,N_1953,N_1537);
or U2548 (N_2548,N_1709,N_1504);
and U2549 (N_2549,N_1660,N_1486);
xnor U2550 (N_2550,N_1708,N_1119);
and U2551 (N_2551,N_1561,N_1755);
and U2552 (N_2552,N_1008,N_1748);
nor U2553 (N_2553,N_1513,N_1171);
nand U2554 (N_2554,N_1198,N_1161);
nor U2555 (N_2555,N_1558,N_1673);
or U2556 (N_2556,N_1766,N_1577);
nor U2557 (N_2557,N_1301,N_1044);
nand U2558 (N_2558,N_1536,N_1508);
or U2559 (N_2559,N_1899,N_1651);
xnor U2560 (N_2560,N_1082,N_1988);
and U2561 (N_2561,N_1613,N_1468);
nor U2562 (N_2562,N_1110,N_1137);
or U2563 (N_2563,N_1429,N_1272);
or U2564 (N_2564,N_1586,N_1155);
xnor U2565 (N_2565,N_1409,N_1617);
nor U2566 (N_2566,N_1072,N_1623);
and U2567 (N_2567,N_1719,N_1844);
nand U2568 (N_2568,N_1107,N_1588);
and U2569 (N_2569,N_1083,N_1710);
xor U2570 (N_2570,N_1102,N_1395);
or U2571 (N_2571,N_1548,N_1021);
and U2572 (N_2572,N_1245,N_1535);
nor U2573 (N_2573,N_1762,N_1810);
and U2574 (N_2574,N_1038,N_1042);
and U2575 (N_2575,N_1673,N_1123);
nor U2576 (N_2576,N_1331,N_1567);
and U2577 (N_2577,N_1808,N_1344);
nor U2578 (N_2578,N_1125,N_1990);
nor U2579 (N_2579,N_1666,N_1878);
or U2580 (N_2580,N_1377,N_1528);
and U2581 (N_2581,N_1858,N_1661);
nand U2582 (N_2582,N_1262,N_1060);
or U2583 (N_2583,N_1828,N_1740);
nand U2584 (N_2584,N_1134,N_1115);
nor U2585 (N_2585,N_1296,N_1161);
and U2586 (N_2586,N_1699,N_1803);
and U2587 (N_2587,N_1601,N_1692);
and U2588 (N_2588,N_1357,N_1774);
nand U2589 (N_2589,N_1218,N_1215);
or U2590 (N_2590,N_1033,N_1100);
nand U2591 (N_2591,N_1495,N_1075);
nor U2592 (N_2592,N_1517,N_1490);
or U2593 (N_2593,N_1314,N_1925);
and U2594 (N_2594,N_1206,N_1850);
nand U2595 (N_2595,N_1227,N_1795);
nand U2596 (N_2596,N_1483,N_1562);
xor U2597 (N_2597,N_1678,N_1590);
and U2598 (N_2598,N_1894,N_1091);
nand U2599 (N_2599,N_1411,N_1795);
nor U2600 (N_2600,N_1564,N_1800);
nand U2601 (N_2601,N_1743,N_1127);
nor U2602 (N_2602,N_1155,N_1323);
nor U2603 (N_2603,N_1681,N_1307);
nand U2604 (N_2604,N_1595,N_1863);
xnor U2605 (N_2605,N_1986,N_1679);
or U2606 (N_2606,N_1476,N_1591);
xnor U2607 (N_2607,N_1101,N_1058);
and U2608 (N_2608,N_1293,N_1813);
nand U2609 (N_2609,N_1102,N_1532);
or U2610 (N_2610,N_1718,N_1300);
and U2611 (N_2611,N_1094,N_1372);
nor U2612 (N_2612,N_1296,N_1260);
nor U2613 (N_2613,N_1855,N_1494);
nor U2614 (N_2614,N_1554,N_1271);
and U2615 (N_2615,N_1624,N_1867);
and U2616 (N_2616,N_1011,N_1534);
or U2617 (N_2617,N_1309,N_1978);
xor U2618 (N_2618,N_1674,N_1938);
xor U2619 (N_2619,N_1678,N_1380);
or U2620 (N_2620,N_1556,N_1510);
xnor U2621 (N_2621,N_1960,N_1344);
nand U2622 (N_2622,N_1008,N_1833);
or U2623 (N_2623,N_1704,N_1363);
or U2624 (N_2624,N_1628,N_1840);
or U2625 (N_2625,N_1307,N_1559);
and U2626 (N_2626,N_1039,N_1763);
nor U2627 (N_2627,N_1243,N_1942);
or U2628 (N_2628,N_1195,N_1785);
nor U2629 (N_2629,N_1773,N_1470);
nand U2630 (N_2630,N_1841,N_1789);
or U2631 (N_2631,N_1794,N_1599);
nand U2632 (N_2632,N_1864,N_1653);
xor U2633 (N_2633,N_1778,N_1241);
and U2634 (N_2634,N_1399,N_1444);
nand U2635 (N_2635,N_1007,N_1682);
nor U2636 (N_2636,N_1769,N_1610);
xnor U2637 (N_2637,N_1139,N_1674);
xnor U2638 (N_2638,N_1493,N_1702);
xnor U2639 (N_2639,N_1553,N_1080);
nor U2640 (N_2640,N_1658,N_1052);
and U2641 (N_2641,N_1304,N_1429);
and U2642 (N_2642,N_1375,N_1629);
nor U2643 (N_2643,N_1641,N_1441);
or U2644 (N_2644,N_1522,N_1496);
nand U2645 (N_2645,N_1789,N_1999);
nor U2646 (N_2646,N_1078,N_1833);
or U2647 (N_2647,N_1277,N_1754);
and U2648 (N_2648,N_1806,N_1613);
and U2649 (N_2649,N_1227,N_1584);
nand U2650 (N_2650,N_1304,N_1959);
xnor U2651 (N_2651,N_1883,N_1537);
nand U2652 (N_2652,N_1636,N_1962);
and U2653 (N_2653,N_1925,N_1146);
nor U2654 (N_2654,N_1710,N_1584);
or U2655 (N_2655,N_1623,N_1420);
nor U2656 (N_2656,N_1961,N_1997);
nand U2657 (N_2657,N_1526,N_1614);
nor U2658 (N_2658,N_1384,N_1525);
nand U2659 (N_2659,N_1555,N_1646);
nand U2660 (N_2660,N_1274,N_1489);
nor U2661 (N_2661,N_1049,N_1041);
and U2662 (N_2662,N_1206,N_1941);
or U2663 (N_2663,N_1349,N_1012);
nand U2664 (N_2664,N_1931,N_1507);
or U2665 (N_2665,N_1724,N_1256);
nor U2666 (N_2666,N_1631,N_1905);
and U2667 (N_2667,N_1106,N_1308);
xnor U2668 (N_2668,N_1488,N_1270);
nand U2669 (N_2669,N_1257,N_1230);
nand U2670 (N_2670,N_1056,N_1182);
nor U2671 (N_2671,N_1475,N_1779);
nand U2672 (N_2672,N_1734,N_1951);
xor U2673 (N_2673,N_1085,N_1677);
nor U2674 (N_2674,N_1754,N_1420);
nor U2675 (N_2675,N_1632,N_1188);
nand U2676 (N_2676,N_1551,N_1108);
nor U2677 (N_2677,N_1773,N_1191);
nand U2678 (N_2678,N_1727,N_1495);
and U2679 (N_2679,N_1183,N_1857);
or U2680 (N_2680,N_1261,N_1132);
or U2681 (N_2681,N_1716,N_1919);
nor U2682 (N_2682,N_1278,N_1331);
nor U2683 (N_2683,N_1264,N_1750);
nor U2684 (N_2684,N_1282,N_1839);
nand U2685 (N_2685,N_1645,N_1065);
nand U2686 (N_2686,N_1080,N_1742);
or U2687 (N_2687,N_1770,N_1407);
and U2688 (N_2688,N_1102,N_1205);
xnor U2689 (N_2689,N_1521,N_1218);
or U2690 (N_2690,N_1170,N_1763);
nor U2691 (N_2691,N_1593,N_1461);
and U2692 (N_2692,N_1393,N_1804);
xor U2693 (N_2693,N_1204,N_1851);
xor U2694 (N_2694,N_1442,N_1962);
nand U2695 (N_2695,N_1640,N_1542);
xnor U2696 (N_2696,N_1727,N_1056);
nor U2697 (N_2697,N_1226,N_1099);
or U2698 (N_2698,N_1221,N_1678);
nor U2699 (N_2699,N_1438,N_1725);
or U2700 (N_2700,N_1760,N_1963);
and U2701 (N_2701,N_1771,N_1542);
nor U2702 (N_2702,N_1810,N_1153);
nor U2703 (N_2703,N_1749,N_1935);
and U2704 (N_2704,N_1333,N_1864);
and U2705 (N_2705,N_1137,N_1951);
xnor U2706 (N_2706,N_1654,N_1274);
and U2707 (N_2707,N_1648,N_1364);
nand U2708 (N_2708,N_1459,N_1396);
and U2709 (N_2709,N_1267,N_1343);
and U2710 (N_2710,N_1762,N_1677);
and U2711 (N_2711,N_1876,N_1274);
or U2712 (N_2712,N_1995,N_1809);
xnor U2713 (N_2713,N_1751,N_1247);
and U2714 (N_2714,N_1289,N_1835);
xnor U2715 (N_2715,N_1637,N_1817);
xor U2716 (N_2716,N_1639,N_1483);
nand U2717 (N_2717,N_1032,N_1352);
nand U2718 (N_2718,N_1001,N_1972);
nor U2719 (N_2719,N_1460,N_1907);
and U2720 (N_2720,N_1567,N_1115);
nand U2721 (N_2721,N_1634,N_1040);
nand U2722 (N_2722,N_1246,N_1625);
or U2723 (N_2723,N_1192,N_1080);
xor U2724 (N_2724,N_1710,N_1030);
or U2725 (N_2725,N_1995,N_1861);
nor U2726 (N_2726,N_1751,N_1435);
nor U2727 (N_2727,N_1176,N_1606);
and U2728 (N_2728,N_1201,N_1645);
nand U2729 (N_2729,N_1639,N_1761);
or U2730 (N_2730,N_1467,N_1289);
nor U2731 (N_2731,N_1735,N_1514);
nand U2732 (N_2732,N_1008,N_1865);
or U2733 (N_2733,N_1492,N_1482);
nor U2734 (N_2734,N_1238,N_1703);
nand U2735 (N_2735,N_1280,N_1213);
nand U2736 (N_2736,N_1053,N_1059);
and U2737 (N_2737,N_1429,N_1290);
or U2738 (N_2738,N_1572,N_1380);
xor U2739 (N_2739,N_1253,N_1735);
nor U2740 (N_2740,N_1175,N_1105);
nor U2741 (N_2741,N_1447,N_1764);
nor U2742 (N_2742,N_1482,N_1231);
nor U2743 (N_2743,N_1717,N_1879);
nand U2744 (N_2744,N_1386,N_1115);
and U2745 (N_2745,N_1505,N_1469);
xor U2746 (N_2746,N_1173,N_1348);
and U2747 (N_2747,N_1187,N_1173);
or U2748 (N_2748,N_1714,N_1962);
or U2749 (N_2749,N_1785,N_1137);
xnor U2750 (N_2750,N_1089,N_1376);
and U2751 (N_2751,N_1497,N_1996);
or U2752 (N_2752,N_1170,N_1023);
nor U2753 (N_2753,N_1646,N_1386);
nand U2754 (N_2754,N_1061,N_1454);
nand U2755 (N_2755,N_1714,N_1220);
nand U2756 (N_2756,N_1775,N_1631);
or U2757 (N_2757,N_1635,N_1357);
nor U2758 (N_2758,N_1564,N_1729);
or U2759 (N_2759,N_1983,N_1168);
nor U2760 (N_2760,N_1517,N_1931);
or U2761 (N_2761,N_1972,N_1517);
nand U2762 (N_2762,N_1943,N_1062);
xor U2763 (N_2763,N_1424,N_1632);
xnor U2764 (N_2764,N_1460,N_1326);
or U2765 (N_2765,N_1015,N_1510);
or U2766 (N_2766,N_1438,N_1647);
and U2767 (N_2767,N_1015,N_1214);
nor U2768 (N_2768,N_1034,N_1830);
nand U2769 (N_2769,N_1605,N_1965);
or U2770 (N_2770,N_1339,N_1577);
nand U2771 (N_2771,N_1034,N_1703);
or U2772 (N_2772,N_1920,N_1555);
nor U2773 (N_2773,N_1917,N_1027);
xnor U2774 (N_2774,N_1390,N_1908);
and U2775 (N_2775,N_1858,N_1640);
or U2776 (N_2776,N_1256,N_1362);
xor U2777 (N_2777,N_1942,N_1714);
and U2778 (N_2778,N_1378,N_1963);
or U2779 (N_2779,N_1764,N_1479);
and U2780 (N_2780,N_1288,N_1970);
xor U2781 (N_2781,N_1797,N_1529);
nand U2782 (N_2782,N_1308,N_1021);
nor U2783 (N_2783,N_1338,N_1060);
nor U2784 (N_2784,N_1456,N_1300);
or U2785 (N_2785,N_1726,N_1190);
nand U2786 (N_2786,N_1904,N_1853);
xnor U2787 (N_2787,N_1974,N_1235);
or U2788 (N_2788,N_1411,N_1366);
or U2789 (N_2789,N_1017,N_1933);
nor U2790 (N_2790,N_1412,N_1321);
and U2791 (N_2791,N_1134,N_1421);
nor U2792 (N_2792,N_1918,N_1869);
nor U2793 (N_2793,N_1537,N_1694);
or U2794 (N_2794,N_1637,N_1106);
or U2795 (N_2795,N_1030,N_1596);
and U2796 (N_2796,N_1014,N_1728);
and U2797 (N_2797,N_1871,N_1970);
and U2798 (N_2798,N_1495,N_1424);
or U2799 (N_2799,N_1266,N_1738);
nand U2800 (N_2800,N_1047,N_1669);
and U2801 (N_2801,N_1838,N_1064);
nor U2802 (N_2802,N_1301,N_1157);
nor U2803 (N_2803,N_1734,N_1336);
xor U2804 (N_2804,N_1062,N_1349);
nor U2805 (N_2805,N_1943,N_1423);
xnor U2806 (N_2806,N_1462,N_1334);
and U2807 (N_2807,N_1175,N_1290);
nor U2808 (N_2808,N_1738,N_1071);
nor U2809 (N_2809,N_1769,N_1943);
nand U2810 (N_2810,N_1730,N_1136);
nand U2811 (N_2811,N_1131,N_1107);
and U2812 (N_2812,N_1443,N_1738);
or U2813 (N_2813,N_1876,N_1546);
nor U2814 (N_2814,N_1366,N_1430);
nor U2815 (N_2815,N_1489,N_1153);
nand U2816 (N_2816,N_1444,N_1002);
nor U2817 (N_2817,N_1771,N_1772);
nand U2818 (N_2818,N_1567,N_1465);
nand U2819 (N_2819,N_1627,N_1390);
or U2820 (N_2820,N_1419,N_1823);
and U2821 (N_2821,N_1105,N_1751);
nand U2822 (N_2822,N_1879,N_1392);
nand U2823 (N_2823,N_1648,N_1476);
nand U2824 (N_2824,N_1655,N_1037);
or U2825 (N_2825,N_1198,N_1170);
or U2826 (N_2826,N_1835,N_1651);
and U2827 (N_2827,N_1669,N_1966);
xnor U2828 (N_2828,N_1029,N_1489);
nor U2829 (N_2829,N_1046,N_1339);
nand U2830 (N_2830,N_1664,N_1557);
nand U2831 (N_2831,N_1005,N_1927);
and U2832 (N_2832,N_1608,N_1513);
and U2833 (N_2833,N_1667,N_1228);
xor U2834 (N_2834,N_1229,N_1672);
and U2835 (N_2835,N_1064,N_1876);
nand U2836 (N_2836,N_1954,N_1017);
or U2837 (N_2837,N_1002,N_1725);
nor U2838 (N_2838,N_1311,N_1814);
nand U2839 (N_2839,N_1012,N_1766);
nand U2840 (N_2840,N_1787,N_1340);
or U2841 (N_2841,N_1200,N_1353);
or U2842 (N_2842,N_1081,N_1228);
and U2843 (N_2843,N_1595,N_1746);
and U2844 (N_2844,N_1977,N_1411);
and U2845 (N_2845,N_1654,N_1724);
nor U2846 (N_2846,N_1064,N_1801);
nor U2847 (N_2847,N_1103,N_1457);
nor U2848 (N_2848,N_1802,N_1896);
xnor U2849 (N_2849,N_1520,N_1087);
and U2850 (N_2850,N_1871,N_1845);
nor U2851 (N_2851,N_1771,N_1310);
and U2852 (N_2852,N_1471,N_1743);
nand U2853 (N_2853,N_1803,N_1998);
nor U2854 (N_2854,N_1659,N_1240);
xor U2855 (N_2855,N_1153,N_1905);
or U2856 (N_2856,N_1452,N_1871);
xnor U2857 (N_2857,N_1188,N_1054);
nand U2858 (N_2858,N_1718,N_1088);
and U2859 (N_2859,N_1155,N_1660);
and U2860 (N_2860,N_1637,N_1352);
xnor U2861 (N_2861,N_1376,N_1161);
or U2862 (N_2862,N_1117,N_1831);
nand U2863 (N_2863,N_1015,N_1068);
or U2864 (N_2864,N_1354,N_1933);
or U2865 (N_2865,N_1324,N_1393);
nor U2866 (N_2866,N_1791,N_1881);
nand U2867 (N_2867,N_1145,N_1897);
and U2868 (N_2868,N_1985,N_1966);
nand U2869 (N_2869,N_1122,N_1089);
and U2870 (N_2870,N_1594,N_1592);
or U2871 (N_2871,N_1607,N_1860);
and U2872 (N_2872,N_1668,N_1069);
and U2873 (N_2873,N_1968,N_1464);
nand U2874 (N_2874,N_1341,N_1474);
nand U2875 (N_2875,N_1065,N_1938);
nor U2876 (N_2876,N_1698,N_1117);
and U2877 (N_2877,N_1001,N_1952);
nor U2878 (N_2878,N_1073,N_1335);
nand U2879 (N_2879,N_1258,N_1355);
nor U2880 (N_2880,N_1680,N_1492);
and U2881 (N_2881,N_1192,N_1368);
xor U2882 (N_2882,N_1140,N_1888);
nor U2883 (N_2883,N_1068,N_1834);
nor U2884 (N_2884,N_1117,N_1304);
nand U2885 (N_2885,N_1372,N_1654);
nand U2886 (N_2886,N_1536,N_1270);
nor U2887 (N_2887,N_1179,N_1999);
and U2888 (N_2888,N_1485,N_1754);
xor U2889 (N_2889,N_1687,N_1693);
or U2890 (N_2890,N_1401,N_1814);
nand U2891 (N_2891,N_1140,N_1518);
nor U2892 (N_2892,N_1346,N_1970);
and U2893 (N_2893,N_1367,N_1138);
xor U2894 (N_2894,N_1917,N_1077);
nor U2895 (N_2895,N_1152,N_1517);
nor U2896 (N_2896,N_1551,N_1421);
or U2897 (N_2897,N_1575,N_1819);
nand U2898 (N_2898,N_1803,N_1519);
nand U2899 (N_2899,N_1409,N_1112);
xnor U2900 (N_2900,N_1604,N_1713);
xor U2901 (N_2901,N_1695,N_1763);
nand U2902 (N_2902,N_1583,N_1386);
and U2903 (N_2903,N_1513,N_1919);
or U2904 (N_2904,N_1144,N_1180);
xnor U2905 (N_2905,N_1439,N_1748);
and U2906 (N_2906,N_1026,N_1659);
and U2907 (N_2907,N_1533,N_1491);
and U2908 (N_2908,N_1426,N_1568);
nand U2909 (N_2909,N_1776,N_1543);
and U2910 (N_2910,N_1263,N_1806);
or U2911 (N_2911,N_1882,N_1935);
nand U2912 (N_2912,N_1987,N_1321);
or U2913 (N_2913,N_1203,N_1480);
xor U2914 (N_2914,N_1571,N_1906);
and U2915 (N_2915,N_1146,N_1406);
or U2916 (N_2916,N_1338,N_1931);
or U2917 (N_2917,N_1167,N_1762);
or U2918 (N_2918,N_1051,N_1121);
nor U2919 (N_2919,N_1157,N_1030);
nor U2920 (N_2920,N_1306,N_1302);
nor U2921 (N_2921,N_1846,N_1481);
and U2922 (N_2922,N_1526,N_1326);
nand U2923 (N_2923,N_1742,N_1287);
nor U2924 (N_2924,N_1288,N_1698);
nand U2925 (N_2925,N_1873,N_1712);
nand U2926 (N_2926,N_1039,N_1786);
nor U2927 (N_2927,N_1572,N_1065);
nand U2928 (N_2928,N_1413,N_1214);
nand U2929 (N_2929,N_1557,N_1212);
nor U2930 (N_2930,N_1709,N_1195);
nand U2931 (N_2931,N_1720,N_1408);
xor U2932 (N_2932,N_1056,N_1328);
or U2933 (N_2933,N_1520,N_1378);
nor U2934 (N_2934,N_1314,N_1315);
nor U2935 (N_2935,N_1351,N_1956);
or U2936 (N_2936,N_1067,N_1338);
or U2937 (N_2937,N_1066,N_1171);
nor U2938 (N_2938,N_1487,N_1068);
and U2939 (N_2939,N_1062,N_1444);
or U2940 (N_2940,N_1452,N_1301);
nand U2941 (N_2941,N_1877,N_1438);
nand U2942 (N_2942,N_1354,N_1292);
xor U2943 (N_2943,N_1412,N_1516);
nor U2944 (N_2944,N_1920,N_1403);
or U2945 (N_2945,N_1128,N_1383);
nand U2946 (N_2946,N_1404,N_1656);
and U2947 (N_2947,N_1604,N_1217);
or U2948 (N_2948,N_1347,N_1817);
or U2949 (N_2949,N_1527,N_1049);
and U2950 (N_2950,N_1434,N_1597);
nand U2951 (N_2951,N_1661,N_1257);
nor U2952 (N_2952,N_1438,N_1357);
nand U2953 (N_2953,N_1925,N_1027);
and U2954 (N_2954,N_1178,N_1572);
nand U2955 (N_2955,N_1342,N_1347);
or U2956 (N_2956,N_1081,N_1854);
or U2957 (N_2957,N_1026,N_1718);
nor U2958 (N_2958,N_1160,N_1222);
xor U2959 (N_2959,N_1781,N_1324);
and U2960 (N_2960,N_1386,N_1125);
nor U2961 (N_2961,N_1964,N_1037);
nand U2962 (N_2962,N_1124,N_1813);
and U2963 (N_2963,N_1505,N_1574);
or U2964 (N_2964,N_1893,N_1668);
or U2965 (N_2965,N_1757,N_1699);
nand U2966 (N_2966,N_1473,N_1134);
nor U2967 (N_2967,N_1111,N_1866);
nand U2968 (N_2968,N_1762,N_1836);
or U2969 (N_2969,N_1865,N_1890);
nor U2970 (N_2970,N_1461,N_1823);
or U2971 (N_2971,N_1075,N_1457);
nand U2972 (N_2972,N_1281,N_1447);
nor U2973 (N_2973,N_1016,N_1421);
nor U2974 (N_2974,N_1636,N_1566);
nor U2975 (N_2975,N_1103,N_1748);
or U2976 (N_2976,N_1442,N_1302);
and U2977 (N_2977,N_1416,N_1094);
nor U2978 (N_2978,N_1300,N_1391);
or U2979 (N_2979,N_1350,N_1943);
nor U2980 (N_2980,N_1506,N_1223);
xnor U2981 (N_2981,N_1296,N_1798);
nor U2982 (N_2982,N_1188,N_1945);
or U2983 (N_2983,N_1613,N_1234);
nor U2984 (N_2984,N_1171,N_1916);
nand U2985 (N_2985,N_1519,N_1897);
nand U2986 (N_2986,N_1649,N_1042);
and U2987 (N_2987,N_1819,N_1441);
and U2988 (N_2988,N_1283,N_1286);
nor U2989 (N_2989,N_1120,N_1186);
nor U2990 (N_2990,N_1104,N_1744);
nor U2991 (N_2991,N_1418,N_1928);
nand U2992 (N_2992,N_1057,N_1288);
nand U2993 (N_2993,N_1000,N_1824);
nor U2994 (N_2994,N_1972,N_1292);
nand U2995 (N_2995,N_1121,N_1579);
nor U2996 (N_2996,N_1693,N_1769);
nor U2997 (N_2997,N_1584,N_1359);
nand U2998 (N_2998,N_1896,N_1606);
and U2999 (N_2999,N_1501,N_1896);
nand UO_0 (O_0,N_2618,N_2180);
and UO_1 (O_1,N_2605,N_2110);
nand UO_2 (O_2,N_2268,N_2823);
nor UO_3 (O_3,N_2368,N_2416);
xor UO_4 (O_4,N_2280,N_2303);
and UO_5 (O_5,N_2253,N_2164);
nand UO_6 (O_6,N_2767,N_2496);
or UO_7 (O_7,N_2924,N_2410);
or UO_8 (O_8,N_2327,N_2464);
nand UO_9 (O_9,N_2182,N_2324);
or UO_10 (O_10,N_2075,N_2377);
and UO_11 (O_11,N_2925,N_2214);
xor UO_12 (O_12,N_2521,N_2523);
nand UO_13 (O_13,N_2020,N_2814);
and UO_14 (O_14,N_2504,N_2449);
nor UO_15 (O_15,N_2536,N_2511);
and UO_16 (O_16,N_2367,N_2480);
nor UO_17 (O_17,N_2503,N_2465);
nand UO_18 (O_18,N_2989,N_2635);
or UO_19 (O_19,N_2561,N_2019);
or UO_20 (O_20,N_2260,N_2205);
and UO_21 (O_21,N_2195,N_2749);
and UO_22 (O_22,N_2971,N_2026);
nand UO_23 (O_23,N_2699,N_2228);
and UO_24 (O_24,N_2724,N_2422);
or UO_25 (O_25,N_2546,N_2983);
nand UO_26 (O_26,N_2350,N_2168);
nor UO_27 (O_27,N_2805,N_2097);
nand UO_28 (O_28,N_2352,N_2151);
nand UO_29 (O_29,N_2117,N_2959);
or UO_30 (O_30,N_2236,N_2219);
or UO_31 (O_31,N_2815,N_2131);
or UO_32 (O_32,N_2152,N_2122);
nor UO_33 (O_33,N_2656,N_2990);
nand UO_34 (O_34,N_2044,N_2506);
xnor UO_35 (O_35,N_2165,N_2060);
xnor UO_36 (O_36,N_2949,N_2556);
nor UO_37 (O_37,N_2756,N_2525);
xor UO_38 (O_38,N_2757,N_2322);
or UO_39 (O_39,N_2156,N_2966);
or UO_40 (O_40,N_2808,N_2944);
and UO_41 (O_41,N_2065,N_2601);
nor UO_42 (O_42,N_2970,N_2568);
or UO_43 (O_43,N_2050,N_2126);
nor UO_44 (O_44,N_2101,N_2302);
or UO_45 (O_45,N_2285,N_2574);
or UO_46 (O_46,N_2399,N_2084);
nor UO_47 (O_47,N_2271,N_2957);
nand UO_48 (O_48,N_2333,N_2658);
xnor UO_49 (O_49,N_2366,N_2866);
xnor UO_50 (O_50,N_2630,N_2755);
nand UO_51 (O_51,N_2922,N_2081);
or UO_52 (O_52,N_2754,N_2598);
nand UO_53 (O_53,N_2397,N_2441);
nand UO_54 (O_54,N_2783,N_2670);
xor UO_55 (O_55,N_2437,N_2940);
and UO_56 (O_56,N_2137,N_2894);
xor UO_57 (O_57,N_2284,N_2715);
and UO_58 (O_58,N_2633,N_2514);
or UO_59 (O_59,N_2313,N_2812);
and UO_60 (O_60,N_2336,N_2896);
and UO_61 (O_61,N_2223,N_2432);
xor UO_62 (O_62,N_2181,N_2495);
or UO_63 (O_63,N_2096,N_2744);
nor UO_64 (O_64,N_2762,N_2042);
and UO_65 (O_65,N_2301,N_2672);
nand UO_66 (O_66,N_2578,N_2479);
nor UO_67 (O_67,N_2895,N_2588);
nor UO_68 (O_68,N_2877,N_2120);
or UO_69 (O_69,N_2270,N_2674);
nor UO_70 (O_70,N_2735,N_2745);
nand UO_71 (O_71,N_2087,N_2770);
and UO_72 (O_72,N_2551,N_2030);
or UO_73 (O_73,N_2473,N_2834);
and UO_74 (O_74,N_2104,N_2747);
xor UO_75 (O_75,N_2321,N_2887);
or UO_76 (O_76,N_2429,N_2171);
xnor UO_77 (O_77,N_2736,N_2472);
nor UO_78 (O_78,N_2974,N_2945);
nor UO_79 (O_79,N_2290,N_2776);
nand UO_80 (O_80,N_2991,N_2451);
nor UO_81 (O_81,N_2162,N_2337);
and UO_82 (O_82,N_2055,N_2821);
nand UO_83 (O_83,N_2047,N_2712);
or UO_84 (O_84,N_2232,N_2936);
and UO_85 (O_85,N_2490,N_2130);
nand UO_86 (O_86,N_2817,N_2294);
xnor UO_87 (O_87,N_2438,N_2882);
or UO_88 (O_88,N_2099,N_2641);
and UO_89 (O_89,N_2984,N_2912);
nor UO_90 (O_90,N_2826,N_2828);
xor UO_91 (O_91,N_2436,N_2299);
and UO_92 (O_92,N_2811,N_2994);
and UO_93 (O_93,N_2406,N_2142);
and UO_94 (O_94,N_2502,N_2937);
nand UO_95 (O_95,N_2952,N_2540);
nor UO_96 (O_96,N_2686,N_2381);
or UO_97 (O_97,N_2080,N_2548);
or UO_98 (O_98,N_2893,N_2390);
nand UO_99 (O_99,N_2376,N_2530);
or UO_100 (O_100,N_2249,N_2146);
and UO_101 (O_101,N_2680,N_2709);
nand UO_102 (O_102,N_2565,N_2610);
nand UO_103 (O_103,N_2741,N_2296);
nor UO_104 (O_104,N_2233,N_2589);
or UO_105 (O_105,N_2033,N_2380);
or UO_106 (O_106,N_2230,N_2391);
or UO_107 (O_107,N_2604,N_2393);
nand UO_108 (O_108,N_2418,N_2558);
nor UO_109 (O_109,N_2003,N_2849);
and UO_110 (O_110,N_2183,N_2807);
xor UO_111 (O_111,N_2961,N_2595);
nand UO_112 (O_112,N_2631,N_2076);
or UO_113 (O_113,N_2953,N_2694);
nor UO_114 (O_114,N_2430,N_2403);
nor UO_115 (O_115,N_2824,N_2577);
or UO_116 (O_116,N_2964,N_2489);
nor UO_117 (O_117,N_2640,N_2873);
xnor UO_118 (O_118,N_2078,N_2455);
or UO_119 (O_119,N_2790,N_2948);
xor UO_120 (O_120,N_2501,N_2043);
nand UO_121 (O_121,N_2174,N_2123);
nor UO_122 (O_122,N_2813,N_2795);
or UO_123 (O_123,N_2201,N_2031);
and UO_124 (O_124,N_2022,N_2338);
and UO_125 (O_125,N_2484,N_2655);
and UO_126 (O_126,N_2668,N_2660);
or UO_127 (O_127,N_2014,N_2213);
or UO_128 (O_128,N_2073,N_2037);
nor UO_129 (O_129,N_2196,N_2899);
xor UO_130 (O_130,N_2144,N_2478);
and UO_131 (O_131,N_2404,N_2837);
nand UO_132 (O_132,N_2408,N_2133);
or UO_133 (O_133,N_2600,N_2951);
and UO_134 (O_134,N_2444,N_2319);
nand UO_135 (O_135,N_2323,N_2697);
nand UO_136 (O_136,N_2759,N_2531);
nor UO_137 (O_137,N_2586,N_2217);
nor UO_138 (O_138,N_2287,N_2279);
nor UO_139 (O_139,N_2066,N_2474);
or UO_140 (O_140,N_2510,N_2785);
and UO_141 (O_141,N_2909,N_2200);
or UO_142 (O_142,N_2650,N_2845);
nor UO_143 (O_143,N_2061,N_2910);
nand UO_144 (O_144,N_2728,N_2879);
nor UO_145 (O_145,N_2861,N_2161);
and UO_146 (O_146,N_2252,N_2127);
or UO_147 (O_147,N_2960,N_2685);
nor UO_148 (O_148,N_2798,N_2209);
xor UO_149 (O_149,N_2291,N_2278);
or UO_150 (O_150,N_2256,N_2802);
xnor UO_151 (O_151,N_2638,N_2039);
or UO_152 (O_152,N_2569,N_2636);
and UO_153 (O_153,N_2431,N_2599);
xor UO_154 (O_154,N_2965,N_2816);
nand UO_155 (O_155,N_2515,N_2713);
or UO_156 (O_156,N_2538,N_2651);
nand UO_157 (O_157,N_2372,N_2726);
or UO_158 (O_158,N_2809,N_2138);
or UO_159 (O_159,N_2239,N_2447);
and UO_160 (O_160,N_2926,N_2150);
and UO_161 (O_161,N_2778,N_2696);
nor UO_162 (O_162,N_2539,N_2850);
nor UO_163 (O_163,N_2663,N_2797);
nand UO_164 (O_164,N_2513,N_2286);
or UO_165 (O_165,N_2257,N_2178);
nand UO_166 (O_166,N_2360,N_2402);
or UO_167 (O_167,N_2742,N_2840);
nor UO_168 (O_168,N_2801,N_2227);
or UO_169 (O_169,N_2224,N_2093);
xnor UO_170 (O_170,N_2722,N_2235);
or UO_171 (O_171,N_2344,N_2012);
xnor UO_172 (O_172,N_2036,N_2520);
nand UO_173 (O_173,N_2976,N_2916);
and UO_174 (O_174,N_2838,N_2481);
nand UO_175 (O_175,N_2897,N_2023);
xnor UO_176 (O_176,N_2424,N_2560);
and UO_177 (O_177,N_2312,N_2269);
or UO_178 (O_178,N_2194,N_2774);
nand UO_179 (O_179,N_2892,N_2332);
and UO_180 (O_180,N_2220,N_2335);
or UO_181 (O_181,N_2086,N_2679);
or UO_182 (O_182,N_2267,N_2004);
nand UO_183 (O_183,N_2967,N_2508);
nand UO_184 (O_184,N_2624,N_2107);
or UO_185 (O_185,N_2609,N_2932);
and UO_186 (O_186,N_2264,N_2914);
and UO_187 (O_187,N_2109,N_2891);
nand UO_188 (O_188,N_2639,N_2248);
and UO_189 (O_189,N_2623,N_2833);
nor UO_190 (O_190,N_2225,N_2751);
and UO_191 (O_191,N_2943,N_2884);
nor UO_192 (O_192,N_2906,N_2564);
and UO_193 (O_193,N_2659,N_2572);
and UO_194 (O_194,N_2516,N_2292);
or UO_195 (O_195,N_2015,N_2996);
and UO_196 (O_196,N_2677,N_2032);
nand UO_197 (O_197,N_2664,N_2450);
or UO_198 (O_198,N_2160,N_2326);
and UO_199 (O_199,N_2750,N_2761);
nor UO_200 (O_200,N_2029,N_2646);
nor UO_201 (O_201,N_2512,N_2730);
and UO_202 (O_202,N_2100,N_2018);
nand UO_203 (O_203,N_2708,N_2027);
nor UO_204 (O_204,N_2051,N_2777);
and UO_205 (O_205,N_2293,N_2606);
nor UO_206 (O_206,N_2218,N_2198);
or UO_207 (O_207,N_2112,N_2671);
or UO_208 (O_208,N_2727,N_2216);
or UO_209 (O_209,N_2375,N_2373);
nand UO_210 (O_210,N_2276,N_2579);
and UO_211 (O_211,N_2973,N_2505);
nor UO_212 (O_212,N_2718,N_2766);
or UO_213 (O_213,N_2364,N_2246);
nor UO_214 (O_214,N_2869,N_2839);
or UO_215 (O_215,N_2038,N_2662);
xnor UO_216 (O_216,N_2445,N_2184);
and UO_217 (O_217,N_2460,N_2192);
or UO_218 (O_218,N_2389,N_2820);
or UO_219 (O_219,N_2534,N_2085);
nand UO_220 (O_220,N_2596,N_2204);
nand UO_221 (O_221,N_2421,N_2673);
and UO_222 (O_222,N_2986,N_2314);
xor UO_223 (O_223,N_2582,N_2584);
nand UO_224 (O_224,N_2443,N_2440);
and UO_225 (O_225,N_2494,N_2028);
xnor UO_226 (O_226,N_2315,N_2265);
nand UO_227 (O_227,N_2738,N_2466);
nand UO_228 (O_228,N_2143,N_2691);
and UO_229 (O_229,N_2346,N_2193);
nor UO_230 (O_230,N_2625,N_2509);
nand UO_231 (O_231,N_2847,N_2522);
or UO_232 (O_232,N_2435,N_2468);
or UO_233 (O_233,N_2304,N_2862);
and UO_234 (O_234,N_2108,N_2931);
nand UO_235 (O_235,N_2005,N_2475);
nand UO_236 (O_236,N_2999,N_2258);
nand UO_237 (O_237,N_2234,N_2665);
xnor UO_238 (O_238,N_2134,N_2563);
nor UO_239 (O_239,N_2024,N_2423);
nand UO_240 (O_240,N_2409,N_2394);
nor UO_241 (O_241,N_2836,N_2958);
xor UO_242 (O_242,N_2116,N_2800);
nand UO_243 (O_243,N_2706,N_2016);
nor UO_244 (O_244,N_2827,N_2825);
or UO_245 (O_245,N_2477,N_2388);
or UO_246 (O_246,N_2345,N_2469);
xnor UO_247 (O_247,N_2251,N_2067);
and UO_248 (O_248,N_2806,N_2591);
nor UO_249 (O_249,N_2056,N_2607);
nand UO_250 (O_250,N_2173,N_2634);
or UO_251 (O_251,N_2359,N_2698);
and UO_252 (O_252,N_2172,N_2678);
nor UO_253 (O_253,N_2632,N_2654);
xnor UO_254 (O_254,N_2954,N_2542);
xor UO_255 (O_255,N_2581,N_2157);
xor UO_256 (O_256,N_2835,N_2125);
nand UO_257 (O_257,N_2769,N_2357);
nand UO_258 (O_258,N_2689,N_2541);
and UO_259 (O_259,N_2907,N_2872);
and UO_260 (O_260,N_2851,N_2476);
xnor UO_261 (O_261,N_2487,N_2457);
nand UO_262 (O_262,N_2692,N_2620);
xor UO_263 (O_263,N_2118,N_2488);
nor UO_264 (O_264,N_2830,N_2237);
or UO_265 (O_265,N_2935,N_2009);
or UO_266 (O_266,N_2946,N_2622);
or UO_267 (O_267,N_2255,N_2119);
nand UO_268 (O_268,N_2412,N_2210);
or UO_269 (O_269,N_2493,N_2064);
nand UO_270 (O_270,N_2463,N_2764);
or UO_271 (O_271,N_2446,N_2780);
nor UO_272 (O_272,N_2102,N_2401);
nand UO_273 (O_273,N_2997,N_2950);
nand UO_274 (O_274,N_2177,N_2361);
nand UO_275 (O_275,N_2203,N_2842);
and UO_276 (O_276,N_2452,N_2746);
and UO_277 (O_277,N_2095,N_2619);
nand UO_278 (O_278,N_2356,N_2865);
nor UO_279 (O_279,N_2433,N_2537);
and UO_280 (O_280,N_2517,N_2331);
and UO_281 (O_281,N_2998,N_2771);
xnor UO_282 (O_282,N_2580,N_2170);
nand UO_283 (O_283,N_2308,N_2804);
and UO_284 (O_284,N_2329,N_2720);
nor UO_285 (O_285,N_2995,N_2855);
nor UO_286 (O_286,N_2316,N_2062);
nand UO_287 (O_287,N_2587,N_2583);
and UO_288 (O_288,N_2492,N_2046);
nor UO_289 (O_289,N_2860,N_2590);
nor UO_290 (O_290,N_2454,N_2867);
or UO_291 (O_291,N_2661,N_2021);
nand UO_292 (O_292,N_2254,N_2486);
nor UO_293 (O_293,N_2532,N_2467);
nor UO_294 (O_294,N_2417,N_2442);
nor UO_295 (O_295,N_2272,N_2566);
xor UO_296 (O_296,N_2787,N_2900);
nor UO_297 (O_297,N_2049,N_2334);
nand UO_298 (O_298,N_2262,N_2621);
nor UO_299 (O_299,N_2310,N_2148);
or UO_300 (O_300,N_2981,N_2841);
xor UO_301 (O_301,N_2616,N_2765);
nor UO_302 (O_302,N_2339,N_2094);
nor UO_303 (O_303,N_2881,N_2667);
nor UO_304 (O_304,N_2202,N_2351);
or UO_305 (O_305,N_2384,N_2544);
nor UO_306 (O_306,N_2535,N_2325);
nor UO_307 (O_307,N_2886,N_2491);
nor UO_308 (O_308,N_2643,N_2693);
xnor UO_309 (O_309,N_2968,N_2413);
and UO_310 (O_310,N_2374,N_2889);
nor UO_311 (O_311,N_2753,N_2627);
nor UO_312 (O_312,N_2238,N_2611);
and UO_313 (O_313,N_2462,N_2186);
and UO_314 (O_314,N_2576,N_2796);
nor UO_315 (O_315,N_2245,N_2675);
nand UO_316 (O_316,N_2034,N_2006);
or UO_317 (O_317,N_2992,N_2642);
nor UO_318 (O_318,N_2387,N_2169);
nand UO_319 (O_319,N_2309,N_2711);
xor UO_320 (O_320,N_2121,N_2939);
nand UO_321 (O_321,N_2306,N_2602);
nor UO_322 (O_322,N_2365,N_2972);
xnor UO_323 (O_323,N_2105,N_2407);
nor UO_324 (O_324,N_2676,N_2092);
nand UO_325 (O_325,N_2420,N_2760);
or UO_326 (O_326,N_2371,N_2215);
nand UO_327 (O_327,N_2550,N_2300);
nor UO_328 (O_328,N_2190,N_2608);
nand UO_329 (O_329,N_2603,N_2637);
or UO_330 (O_330,N_2348,N_2305);
nor UO_331 (O_331,N_2930,N_2045);
xor UO_332 (O_332,N_2552,N_2434);
xor UO_333 (O_333,N_2054,N_2275);
or UO_334 (O_334,N_2002,N_2941);
or UO_335 (O_335,N_2079,N_2427);
nor UO_336 (O_336,N_2775,N_2231);
xnor UO_337 (O_337,N_2793,N_2135);
nand UO_338 (O_338,N_2528,N_2261);
and UO_339 (O_339,N_2593,N_2363);
and UO_340 (O_340,N_2854,N_2132);
nand UO_341 (O_341,N_2396,N_2773);
nand UO_342 (O_342,N_2281,N_2197);
and UO_343 (O_343,N_2189,N_2555);
or UO_344 (O_344,N_2657,N_2282);
or UO_345 (O_345,N_2519,N_2058);
nand UO_346 (O_346,N_2784,N_2263);
or UO_347 (O_347,N_2048,N_2880);
xnor UO_348 (O_348,N_2547,N_2977);
nand UO_349 (O_349,N_2707,N_2859);
and UO_350 (O_350,N_2928,N_2848);
or UO_351 (O_351,N_2752,N_2179);
nand UO_352 (O_352,N_2781,N_2794);
or UO_353 (O_353,N_2063,N_2008);
nand UO_354 (O_354,N_2947,N_2905);
nand UO_355 (O_355,N_2035,N_2113);
nor UO_356 (O_356,N_2355,N_2353);
and UO_357 (O_357,N_2311,N_2690);
nor UO_358 (O_358,N_2340,N_2297);
nor UO_359 (O_359,N_2386,N_2057);
or UO_360 (O_360,N_2259,N_2459);
nand UO_361 (O_361,N_2072,N_2846);
or UO_362 (O_362,N_2111,N_2498);
or UO_363 (O_363,N_2158,N_2853);
or UO_364 (O_364,N_2740,N_2725);
and UO_365 (O_365,N_2653,N_2714);
nand UO_366 (O_366,N_2342,N_2874);
or UO_367 (O_367,N_2549,N_2307);
nand UO_368 (O_368,N_2975,N_2649);
nand UO_369 (O_369,N_2684,N_2571);
and UO_370 (O_370,N_2898,N_2832);
or UO_371 (O_371,N_2803,N_2383);
nor UO_372 (O_372,N_2226,N_2758);
nor UO_373 (O_373,N_2128,N_2149);
xnor UO_374 (O_374,N_2938,N_2732);
or UO_375 (O_375,N_2915,N_2933);
or UO_376 (O_376,N_2320,N_2969);
nand UO_377 (O_377,N_2318,N_2956);
xnor UO_378 (O_378,N_2426,N_2629);
nand UO_379 (O_379,N_2083,N_2382);
xnor UO_380 (O_380,N_2266,N_2920);
nor UO_381 (O_381,N_2734,N_2557);
and UO_382 (O_382,N_2704,N_2000);
nand UO_383 (O_383,N_2191,N_2013);
nand UO_384 (O_384,N_2592,N_2145);
nor UO_385 (O_385,N_2929,N_2358);
or UO_386 (O_386,N_2917,N_2461);
nand UO_387 (O_387,N_2703,N_2074);
or UO_388 (O_388,N_2883,N_2980);
nor UO_389 (O_389,N_2717,N_2543);
nand UO_390 (O_390,N_2103,N_2985);
nand UO_391 (O_391,N_2283,N_2695);
and UO_392 (O_392,N_2818,N_2669);
nor UO_393 (O_393,N_2878,N_2385);
or UO_394 (O_394,N_2106,N_2347);
xor UO_395 (O_395,N_2617,N_2328);
nor UO_396 (O_396,N_2567,N_2615);
or UO_397 (O_397,N_2153,N_2700);
or UO_398 (O_398,N_2955,N_2763);
nor UO_399 (O_399,N_2369,N_2439);
nand UO_400 (O_400,N_2507,N_2229);
or UO_401 (O_401,N_2856,N_2483);
nor UO_402 (O_402,N_2918,N_2139);
xor UO_403 (O_403,N_2124,N_2533);
and UO_404 (O_404,N_2902,N_2743);
xnor UO_405 (O_405,N_2362,N_2088);
nor UO_406 (O_406,N_2570,N_2978);
and UO_407 (O_407,N_2244,N_2831);
and UO_408 (O_408,N_2829,N_2559);
or UO_409 (O_409,N_2870,N_2482);
or UO_410 (O_410,N_2001,N_2871);
nor UO_411 (O_411,N_2868,N_2527);
xnor UO_412 (O_412,N_2748,N_2702);
nand UO_413 (O_413,N_2876,N_2011);
xor UO_414 (O_414,N_2628,N_2415);
nor UO_415 (O_415,N_2163,N_2059);
nand UO_416 (O_416,N_2167,N_2129);
and UO_417 (O_417,N_2666,N_2370);
or UO_418 (O_418,N_2212,N_2927);
xnor UO_419 (O_419,N_2518,N_2068);
and UO_420 (O_420,N_2988,N_2411);
nor UO_421 (O_421,N_2626,N_2987);
nor UO_422 (O_422,N_2553,N_2500);
xnor UO_423 (O_423,N_2010,N_2354);
xor UO_424 (O_424,N_2993,N_2791);
nor UO_425 (O_425,N_2136,N_2979);
and UO_426 (O_426,N_2400,N_2207);
nor UO_427 (O_427,N_2017,N_2526);
nand UO_428 (O_428,N_2792,N_2395);
xor UO_429 (O_429,N_2497,N_2458);
nor UO_430 (O_430,N_2141,N_2456);
or UO_431 (O_431,N_2779,N_2863);
and UO_432 (O_432,N_2140,N_2901);
xnor UO_433 (O_433,N_2211,N_2890);
and UO_434 (O_434,N_2683,N_2295);
and UO_435 (O_435,N_2904,N_2185);
nor UO_436 (O_436,N_2962,N_2188);
nor UO_437 (O_437,N_2612,N_2982);
xnor UO_438 (O_438,N_2090,N_2716);
nand UO_439 (O_439,N_2739,N_2040);
or UO_440 (O_440,N_2647,N_2575);
and UO_441 (O_441,N_2274,N_2701);
xor UO_442 (O_442,N_2378,N_2597);
or UO_443 (O_443,N_2705,N_2819);
nor UO_444 (O_444,N_2379,N_2199);
xor UO_445 (O_445,N_2903,N_2154);
or UO_446 (O_446,N_2070,N_2098);
xnor UO_447 (O_447,N_2562,N_2222);
nand UO_448 (O_448,N_2688,N_2242);
nor UO_449 (O_449,N_2864,N_2942);
nand UO_450 (O_450,N_2768,N_2573);
or UO_451 (O_451,N_2919,N_2052);
nor UO_452 (O_452,N_2614,N_2613);
or UO_453 (O_453,N_2448,N_2250);
nor UO_454 (O_454,N_2398,N_2007);
or UO_455 (O_455,N_2414,N_2789);
or UO_456 (O_456,N_2524,N_2392);
xnor UO_457 (O_457,N_2077,N_2529);
and UO_458 (O_458,N_2843,N_2545);
nand UO_459 (O_459,N_2786,N_2913);
nand UO_460 (O_460,N_2240,N_2221);
nor UO_461 (O_461,N_2857,N_2428);
or UO_462 (O_462,N_2349,N_2343);
nand UO_463 (O_463,N_2710,N_2934);
or UO_464 (O_464,N_2298,N_2485);
nor UO_465 (O_465,N_2288,N_2471);
nand UO_466 (O_466,N_2115,N_2822);
or UO_467 (O_467,N_2921,N_2788);
or UO_468 (O_468,N_2648,N_2175);
or UO_469 (O_469,N_2810,N_2844);
nor UO_470 (O_470,N_2645,N_2554);
nor UO_471 (O_471,N_2723,N_2071);
nand UO_472 (O_472,N_2594,N_2682);
nand UO_473 (O_473,N_2114,N_2089);
and UO_474 (O_474,N_2852,N_2888);
nor UO_475 (O_475,N_2858,N_2963);
and UO_476 (O_476,N_2166,N_2585);
nand UO_477 (O_477,N_2499,N_2147);
nand UO_478 (O_478,N_2082,N_2721);
or UO_479 (O_479,N_2875,N_2923);
or UO_480 (O_480,N_2731,N_2317);
xnor UO_481 (O_481,N_2729,N_2733);
or UO_482 (O_482,N_2644,N_2799);
nand UO_483 (O_483,N_2885,N_2025);
xor UO_484 (O_484,N_2453,N_2405);
xor UO_485 (O_485,N_2155,N_2187);
and UO_486 (O_486,N_2425,N_2681);
or UO_487 (O_487,N_2687,N_2341);
nand UO_488 (O_488,N_2911,N_2719);
and UO_489 (O_489,N_2243,N_2289);
or UO_490 (O_490,N_2782,N_2247);
nand UO_491 (O_491,N_2091,N_2277);
and UO_492 (O_492,N_2208,N_2330);
xnor UO_493 (O_493,N_2241,N_2273);
nand UO_494 (O_494,N_2470,N_2737);
xor UO_495 (O_495,N_2176,N_2053);
nor UO_496 (O_496,N_2069,N_2419);
and UO_497 (O_497,N_2041,N_2772);
and UO_498 (O_498,N_2206,N_2652);
or UO_499 (O_499,N_2908,N_2159);
endmodule